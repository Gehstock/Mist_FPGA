library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity VICTORY_ROM_PGM_0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of VICTORY_ROM_PGM_0 is
	type rom is array(0 to  10239) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"31",X"00",X"44",X"C3",X"40",X"02",X"00",X"FF",X"FF",X"FF",X"FF",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"24",X"52",X"22",X"75",X"0D",X"01",X"69",X"02",X"21",X"B0",X"0D",X"36",X"00",X"11",
		X"B1",X"0D",X"ED",X"B0",X"21",X"00",X"00",X"22",X"69",X"0D",X"22",X"6B",X"0D",X"22",X"61",X"0D",
		X"22",X"63",X"0D",X"DD",X"36",X"F5",X"00",X"3A",X"C9",X"33",X"20",X"4C",X"45",X"56",X"45",X"4C",
		X"20",X"4D",X"41",X"54",X"52",X"49",X"58",X"20",X"50",X"52",X"4F",X"54",X"45",X"43",X"54",X"49",
		X"4F",X"4E",X"52",X"30",X"51",X"1A",X"FE",X"2F",X"20",X"F2",X"3E",X"0D",X"12",X"13",X"3E",X"01",
		X"32",X"86",X"0D",X"1A",X"13",X"21",X"F5",X"E5",X"21",X"00",X"40",X"34",X"AF",X"32",X"01",X"70",
		X"3C",X"32",X"01",X"70",X"3A",X"00",X"78",X"E1",X"F1",X"C9",X"21",X"F5",X"C5",X"D5",X"E5",X"DD",
		X"E5",X"FD",X"E5",X"3A",X"00",X"78",X"CD",X"22",X"01",X"AF",X"32",X"01",X"70",X"3E",X"01",X"32",
		X"01",X"70",X"21",X"00",X"40",X"7E",X"BE",X"28",X"FD",X"3A",X"00",X"70",X"CB",X"5F",X"3E",X"01",
		X"28",X"04",X"3A",X"09",X"40",X"2F",X"32",X"06",X"70",X"32",X"07",X"70",X"21",X"4E",X"40",X"11",
		X"00",X"58",X"01",X"80",X"00",X"ED",X"B0",X"DD",X"21",X"2C",X"40",X"3A",X"00",X"60",X"CD",X"21",
		X"13",X"3A",X"00",X"68",X"CD",X"21",X"13",X"3A",X"00",X"70",X"CD",X"21",X"13",X"DD",X"21",X"B8",
		X"1B",X"CD",X"31",X"13",X"11",X"D4",X"1B",X"28",X"08",X"CD",X"31",X"13",X"11",X"DC",X"1B",X"20",
		X"29",X"3A",X"00",X"68",X"07",X"07",X"07",X"E6",X"06",X"6F",X"26",X"00",X"19",X"3A",X"14",X"40",
		X"86",X"27",X"32",X"14",X"40",X"23",X"3A",X"15",X"40",X"8E",X"27",X"30",X"02",X"3E",X"99",X"32",
		X"15",X"40",X"CD",X"3A",X"12",X"3E",X"14",X"32",X"0D",X"40",X"3E",X"01",X"21",X"0D",X"40",X"35",
		X"F2",X"15",X"01",X"34",X"AF",X"32",X"03",X"60",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"F1",
		X"C9",X"21",X"DD",X"21",X"20",X"42",X"3A",X"09",X"40",X"FE",X"02",X"CA",X"5F",X"01",X"DD",X"CB",
		X"00",X"46",X"C2",X"64",X"01",X"DD",X"CB",X"00",X"4E",X"C4",X"9F",X"01",X"DD",X"CB",X"00",X"66",
		X"C4",X"E3",X"01",X"DD",X"CB",X"00",X"6E",X"C4",X"00",X"02",X"DD",X"CB",X"00",X"76",X"C4",X"22",
		X"02",X"DD",X"CB",X"00",X"56",X"C4",X"B3",X"01",X"DD",X"CB",X"00",X"5E",X"C4",X"C6",X"01",X"DD",
		X"CB",X"01",X"46",X"C9",X"3A",X"47",X"01",X"2A",X"22",X"42",X"7E",X"32",X"00",X"78",X"FE",X"FF",
		X"CA",X"99",X"01",X"3E",X"01",X"32",X"06",X"68",X"32",X"07",X"68",X"DD",X"7E",X"04",X"B7",X"28",
		X"08",X"3A",X"35",X"01",X"DD",X"35",X"04",X"18",X"C8",X"23",X"7E",X"DD",X"77",X"04",X"3E",X"FF",
		X"32",X"00",X"78",X"23",X"22",X"22",X"42",X"18",X"B8",X"DD",X"CB",X"00",X"86",X"18",X"B2",X"DD",
		X"7E",X"05",X"FE",X"FF",X"32",X"00",X"78",X"28",X"04",X"DD",X"35",X"05",X"C9",X"DD",X"CB",X"00",
		X"8E",X"C9",X"21",X"3E",X"01",X"32",X"03",X"68",X"DD",X"35",X"06",X"F0",X"AF",X"32",X"03",X"68",
		X"DD",X"CB",X"00",X"96",X"C9",X"21",X"DD",X"7E",X"07",X"B7",X"28",X"0D",X"2F",X"E6",X"02",X"CD",
		X"58",X"13",X"32",X"05",X"68",X"DD",X"35",X"07",X"C9",X"DD",X"CB",X"00",X"9E",X"AF",X"32",X"05",
		X"68",X"C9",X"21",X"DD",X"7E",X"08",X"B7",X"28",X"0D",X"2F",X"E6",X"07",X"87",X"87",X"87",X"32",
		X"00",X"78",X"DD",X"35",X"08",X"C9",X"3E",X"FF",X"32",X"00",X"78",X"DD",X"CB",X"00",X"A6",X"C9",
		X"DD",X"7E",X"09",X"FE",X"80",X"28",X"10",X"C6",X"04",X"DD",X"77",X"09",X"ED",X"44",X"C6",X"40",
		X"CD",X"53",X"13",X"32",X"00",X"78",X"C9",X"3E",X"FF",X"32",X"00",X"78",X"DD",X"CB",X"00",X"AE",
		X"C9",X"21",X"DD",X"7E",X"0A",X"FE",X"FF",X"CA",X"35",X"02",X"DD",X"34",X"0A",X"E6",X"1F",X"87",
		X"87",X"32",X"00",X"78",X"C9",X"3E",X"FF",X"32",X"00",X"78",X"DD",X"CB",X"00",X"B6",X"C9",X"21",
		X"31",X"00",X"44",X"CD",X"AA",X"02",X"CD",X"A4",X"10",X"DD",X"21",X"00",X"50",X"0E",X"10",X"06",
		X"10",X"78",X"C6",X"02",X"E6",X"FC",X"FE",X"08",X"28",X"10",X"DD",X"36",X"00",X"68",X"DD",X"36",
		X"01",X"69",X"DD",X"36",X"20",X"6A",X"DD",X"36",X"21",X"6B",X"DD",X"23",X"DD",X"23",X"10",X"E1",
		X"11",X"20",X"00",X"DD",X"19",X"CD",X"7B",X"00",X"0D",X"20",X"D4",X"21",X"64",X"00",X"CD",X"A0",
		X"03",X"DD",X"21",X"00",X"18",X"CD",X"7B",X"11",X"21",X"64",X"00",X"CD",X"A0",X"03",X"18",X"01",
		X"21",X"31",X"00",X"44",X"AF",X"32",X"09",X"40",X"21",X"D2",X"18",X"AF",X"86",X"2C",X"20",X"FC",
		X"08",X"CD",X"C2",X"02",X"CD",X"81",X"03",X"18",X"E8",X"21",X"21",X"00",X"40",X"11",X"01",X"40",
		X"01",X"2F",X"02",X"36",X"00",X"ED",X"B0",X"21",X"32",X"40",X"22",X"26",X"40",X"CD",X"A4",X"10",
		X"C9",X"21",X"CD",X"A4",X"10",X"DD",X"21",X"FB",X"53",X"06",X"20",X"11",X"E0",X"FF",X"DD",X"36",
		X"FF",X"90",X"DD",X"36",X"00",X"90",X"DD",X"36",X"01",X"90",X"DD",X"36",X"02",X"90",X"DD",X"19",
		X"10",X"EC",X"18",X"01",X"21",X"21",X"64",X"00",X"CD",X"A0",X"03",X"DD",X"21",X"84",X"40",X"FD",
		X"21",X"FB",X"53",X"21",X"32",X"1A",X"01",X"10",X"C0",X"18",X"01",X"21",X"78",X"E6",X"07",X"20",
		X"13",X"0D",X"FA",X"14",X"03",X"7E",X"2B",X"FD",X"77",X"01",X"7E",X"2B",X"FD",X"77",X"00",X"11",
		X"20",X"00",X"FD",X"19",X"DD",X"34",X"00",X"DD",X"34",X"02",X"C5",X"E5",X"DD",X"E5",X"21",X"01",
		X"00",X"CD",X"A0",X"03",X"DD",X"E1",X"E1",X"C1",X"10",X"D2",X"DD",X"21",X"89",X"19",X"DD",X"6E",
		X"00",X"DD",X"7E",X"01",X"FE",X"FF",X"CA",X"54",X"03",X"E6",X"03",X"C6",X"50",X"67",X"DD",X"7E",
		X"01",X"CB",X"3F",X"CB",X"3F",X"C6",X"90",X"77",X"21",X"01",X"00",X"CD",X"A0",X"03",X"DD",X"23",
		X"DD",X"23",X"18",X"DA",X"21",X"32",X"00",X"CD",X"A0",X"03",X"DD",X"21",X"74",X"03",X"CD",X"7B",
		X"11",X"21",X"64",X"00",X"CD",X"A0",X"03",X"DD",X"21",X"61",X"18",X"CD",X"7B",X"11",X"21",X"F4",
		X"01",X"C3",X"A0",X"03",X"E5",X"51",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"24",X"FF",X"FF",
		X"21",X"3E",X"02",X"32",X"09",X"40",X"21",X"76",X"1A",X"22",X"0E",X"40",X"21",X"A0",X"0F",X"22",
		X"2A",X"40",X"21",X"42",X"40",X"22",X"26",X"40",X"CD",X"12",X"05",X"CD",X"CA",X"04",X"C9",X"21",
		X"CD",X"7B",X"00",X"3A",X"15",X"40",X"B7",X"C2",X"B1",X"03",X"2B",X"7C",X"B5",X"20",X"F1",X"C9",
		X"21",X"31",X"00",X"44",X"CD",X"A4",X"10",X"DD",X"21",X"23",X"18",X"CD",X"7B",X"11",X"CD",X"7B",
		X"00",X"3A",X"15",X"40",X"FE",X"01",X"28",X"07",X"DD",X"21",X"4E",X"18",X"CD",X"7B",X"11",X"DD",
		X"21",X"BC",X"1B",X"CD",X"31",X"13",X"01",X"99",X"01",X"28",X"08",X"CD",X"31",X"13",X"01",X"98",
		X"02",X"20",X"DB",X"3A",X"15",X"40",X"B8",X"38",X"D5",X"81",X"27",X"32",X"15",X"40",X"78",X"3D",
		X"32",X"0A",X"40",X"C3",X"F7",X"03",X"21",X"21",X"5C",X"1A",X"11",X"32",X"40",X"01",X"10",X"00",
		X"ED",X"B0",X"3A",X"00",X"70",X"CB",X"57",X"28",X"08",X"3E",X"02",X"32",X"39",X"40",X"32",X"41",
		X"40",X"AF",X"32",X"09",X"40",X"3A",X"09",X"40",X"B7",X"DD",X"21",X"32",X"40",X"28",X"04",X"DD",
		X"21",X"3A",X"40",X"DD",X"22",X"26",X"40",X"DD",X"7E",X"07",X"B7",X"CA",X"8A",X"04",X"DD",X"6E",
		X"04",X"DD",X"66",X"05",X"22",X"0E",X"40",X"DD",X"E5",X"CD",X"A4",X"10",X"3A",X"09",X"40",X"DD",
		X"21",X"56",X"19",X"B7",X"28",X"04",X"DD",X"21",X"65",X"19",X"CD",X"7B",X"11",X"DD",X"2A",X"26",
		X"40",X"CD",X"A6",X"12",X"DD",X"E1",X"CD",X"12",X"05",X"AF",X"21",X"E4",X"1B",X"CD",X"F5",X"10",
		X"CD",X"CA",X"04",X"CD",X"7B",X"00",X"3A",X"20",X"42",X"CB",X"47",X"20",X"F6",X"DD",X"2A",X"26",
		X"40",X"DD",X"35",X"07",X"FA",X"8A",X"04",X"3A",X"0A",X"40",X"B7",X"CA",X"15",X"04",X"3A",X"09",
		X"40",X"EE",X"01",X"32",X"09",X"40",X"C3",X"15",X"04",X"21",X"DD",X"21",X"BA",X"04",X"CD",X"7B",
		X"11",X"06",X"64",X"CD",X"7B",X"00",X"10",X"FB",X"DD",X"2A",X"26",X"40",X"DD",X"CB",X"07",X"7E",
		X"28",X"04",X"DD",X"36",X"07",X"00",X"3A",X"0A",X"40",X"B7",X"3A",X"39",X"40",X"21",X"41",X"40",
		X"28",X"01",X"B6",X"B7",X"CA",X"91",X"02",X"C3",X"77",X"04",X"90",X"50",X"47",X"41",X"4D",X"45",
		X"20",X"4F",X"56",X"45",X"52",X"5B",X"24",X"FF",X"FF",X"21",X"2A",X"1E",X"40",X"23",X"22",X"1E",
		X"40",X"3A",X"09",X"40",X"FE",X"02",X"20",X"0A",X"2A",X"2A",X"40",X"2B",X"22",X"2A",X"40",X"CB",
		X"7C",X"C0",X"CD",X"7B",X"00",X"CD",X"8C",X"09",X"CD",X"DF",X"05",X"CD",X"31",X"0B",X"CD",X"95",
		X"0F",X"CD",X"25",X"09",X"CD",X"0E",X"0C",X"CD",X"EF",X"0E",X"CD",X"3A",X"0A",X"CD",X"3B",X"07",
		X"CD",X"23",X"10",X"20",X"C5",X"CD",X"57",X"10",X"3A",X"06",X"40",X"FE",X"FF",X"C2",X"CA",X"04",
		X"C9",X"21",X"21",X"35",X"1A",X"11",X"F6",X"41",X"01",X"20",X"00",X"ED",X"B0",X"CD",X"A4",X"10",
		X"3E",X"01",X"32",X"04",X"70",X"21",X"00",X"04",X"22",X"16",X"40",X"3E",X"80",X"32",X"01",X"40",
		X"CD",X"F6",X"09",X"21",X"D3",X"40",X"06",X"0A",X"11",X"08",X"00",X"36",X"FF",X"19",X"10",X"FB",
		X"21",X"56",X"1A",X"11",X"CE",X"40",X"01",X"08",X"00",X"ED",X"B0",X"21",X"D3",X"41",X"06",X"06",
		X"11",X"06",X"00",X"36",X"FF",X"19",X"10",X"FB",X"21",X"23",X"41",X"11",X"09",X"00",X"06",X"14",
		X"36",X"FF",X"19",X"10",X"FB",X"DD",X"21",X"E0",X"53",X"06",X"20",X"11",X"E0",X"FF",X"DD",X"36",
		X"04",X"90",X"DD",X"36",X"05",X"2B",X"0E",X"90",X"78",X"E6",X"07",X"20",X"02",X"0E",X"97",X"DD",
		X"71",X"1C",X"DD",X"36",X"1D",X"90",X"DD",X"36",X"1E",X"90",X"DD",X"19",X"10",X"E0",X"DD",X"21",
		X"D4",X"05",X"CD",X"7B",X"11",X"3E",X"95",X"21",X"A1",X"53",X"11",X"41",X"50",X"06",X"03",X"77",
		X"12",X"23",X"13",X"10",X"FA",X"3E",X"9A",X"32",X"04",X"52",X"3E",X"98",X"32",X"E4",X"51",X"AF",
		X"32",X"05",X"40",X"32",X"06",X"40",X"32",X"08",X"40",X"32",X"0B",X"40",X"3E",X"B8",X"32",X"07",
		X"40",X"21",X"00",X"00",X"22",X"12",X"40",X"06",X"20",X"C5",X"CD",X"E1",X"06",X"C1",X"10",X"F9",
		X"CD",X"F6",X"09",X"C9",X"25",X"52",X"52",X"41",X"44",X"41",X"52",X"24",X"FF",X"FF",X"21",X"3A",
		X"1E",X"40",X"2F",X"E6",X"03",X"CC",X"F4",X"05",X"CD",X"90",X"06",X"3A",X"1E",X"40",X"E6",X"01",
		X"CC",X"E1",X"06",X"C9",X"3A",X"06",X"40",X"B7",X"C0",X"CD",X"76",X"06",X"21",X"23",X"52",X"06",
		X"04",X"FD",X"21",X"0F",X"1A",X"11",X"F6",X"41",X"0E",X"08",X"AF",X"EB",X"B6",X"23",X"0D",X"20",
		X"FB",X"EB",X"B7",X"28",X"04",X"FD",X"7E",X"00",X"77",X"FD",X"23",X"D5",X"11",X"E0",X"FF",X"19",
		X"D1",X"10",X"E5",X"DD",X"21",X"CE",X"40",X"06",X"0A",X"DD",X"7E",X"05",X"FE",X"FF",X"CA",X"6C",
		X"06",X"DD",X"5E",X"00",X"DD",X"56",X"01",X"CB",X"3A",X"CB",X"1B",X"7B",X"E6",X"E0",X"5F",X"21",
		X"E1",X"53",X"B7",X"ED",X"52",X"DD",X"7E",X"02",X"FE",X"8C",X"30",X"06",X"2C",X"FE",X"46",X"30",
		X"01",X"2C",X"DD",X"7E",X"05",X"B7",X"0E",X"0D",X"28",X"02",X"0E",X"0C",X"FE",X"58",X"20",X"02",
		X"0E",X"42",X"7E",X"FE",X"95",X"28",X"05",X"FE",X"10",X"38",X"01",X"71",X"11",X"08",X"00",X"DD",
		X"19",X"05",X"C2",X"29",X"06",X"C9",X"DD",X"21",X"81",X"53",X"06",X"1A",X"11",X"E0",X"FF",X"DD",
		X"36",X"00",X"90",X"DD",X"36",X"01",X"90",X"DD",X"36",X"02",X"90",X"DD",X"19",X"10",X"F0",X"C9",
		X"21",X"8E",X"40",X"06",X"20",X"36",X"00",X"23",X"10",X"FB",X"FD",X"21",X"8E",X"40",X"0E",X"08",
		X"06",X"0A",X"DD",X"21",X"CE",X"40",X"DD",X"7E",X"05",X"FE",X"FF",X"CA",X"D7",X"06",X"CD",X"67",
		X"13",X"C2",X"D7",X"06",X"7D",X"D6",X"08",X"FD",X"77",X"00",X"3E",X"F8",X"DD",X"96",X"02",X"FD",
		X"77",X"03",X"DD",X"7E",X"04",X"FD",X"77",X"01",X"DD",X"7E",X"03",X"C6",X"05",X"FD",X"77",X"02",
		X"11",X"04",X"00",X"FD",X"19",X"0D",X"C8",X"11",X"08",X"00",X"DD",X"19",X"05",X"C2",X"A6",X"06",
		X"C9",X"2A",X"16",X"40",X"3A",X"07",X"40",X"C6",X"08",X"32",X"07",X"40",X"CD",X"4E",X"13",X"19",
		X"CD",X"9B",X"13",X"3A",X"1E",X"40",X"E6",X"0F",X"CC",X"F6",X"09",X"3A",X"09",X"40",X"FE",X"02",
		X"28",X"19",X"B7",X"21",X"A0",X"53",X"28",X"03",X"21",X"40",X"51",X"3A",X"1E",X"40",X"CB",X"67",
		X"3E",X"0F",X"28",X"03",X"3A",X"09",X"40",X"3C",X"77",X"18",X"10",X"21",X"00",X"00",X"22",X"42",
		X"40",X"22",X"44",X"40",X"3A",X"15",X"40",X"B7",X"C2",X"B1",X"03",X"2A",X"12",X"40",X"7C",X"B5",
		X"C8",X"CD",X"9B",X"13",X"21",X"00",X"00",X"22",X"12",X"40",X"C9",X"3A",X"06",X"40",X"CB",X"7F",
		X"C0",X"3A",X"09",X"40",X"FE",X"02",X"CA",X"D3",X"07",X"B7",X"DD",X"21",X"C0",X"1B",X"28",X"04",
		X"DD",X"21",X"C8",X"1B",X"DD",X"E5",X"FD",X"21",X"D4",X"40",X"CD",X"9D",X"07",X"FD",X"23",X"DD",
		X"E1",X"11",X"04",X"00",X"DD",X"19",X"CD",X"9D",X"07",X"CD",X"81",X"07",X"3A",X"09",X"40",X"B7",
		X"DD",X"21",X"D0",X"1B",X"28",X"04",X"DD",X"21",X"D2",X"1B",X"CD",X"31",X"13",X"CC",X"65",X"08",
		X"C9",X"3A",X"CF",X"40",X"B7",X"20",X"08",X"3A",X"D4",X"40",X"CB",X"7F",X"C8",X"18",X"09",X"FE",
		X"07",X"C0",X"3A",X"D4",X"40",X"CB",X"7F",X"C0",X"AF",X"32",X"D4",X"40",X"C9",X"3A",X"1E",X"40",
		X"E6",X"03",X"C0",X"CD",X"31",X"13",X"20",X"10",X"FD",X"7E",X"00",X"FE",X"08",X"C8",X"FD",X"CB",
		X"00",X"7E",X"20",X"1A",X"FD",X"34",X"00",X"C9",X"CD",X"31",X"13",X"20",X"11",X"FD",X"7E",X"00",
		X"FE",X"F8",X"C8",X"B7",X"28",X"04",X"CB",X"7F",X"28",X"04",X"FD",X"35",X"00",X"C9",X"AF",X"FD",
		X"77",X"00",X"C9",X"CD",X"C2",X"15",X"FE",X"32",X"0E",X"0A",X"D2",X"53",X"08",X"DD",X"21",X"D6",
		X"40",X"06",X"09",X"0E",X"FF",X"DD",X"7E",X"05",X"FE",X"FF",X"CA",X"3F",X"08",X"FE",X"58",X"CA",
		X"3F",X"08",X"C5",X"DD",X"7E",X"06",X"CD",X"4E",X"13",X"EB",X"29",X"29",X"29",X"29",X"DD",X"5E",
		X"00",X"DD",X"56",X"01",X"19",X"ED",X"5B",X"CE",X"40",X"CD",X"08",X"09",X"47",X"B7",X"20",X"01",
		X"4F",X"59",X"D5",X"DD",X"7E",X"07",X"87",X"87",X"87",X"DD",X"86",X"02",X"6F",X"26",X"00",X"ED",
		X"5B",X"D0",X"40",X"54",X"CD",X"08",X"09",X"B7",X"20",X"01",X"4F",X"D1",X"51",X"80",X"C1",X"B9",
		X"30",X"0D",X"FE",X"0A",X"30",X"04",X"CB",X"2B",X"CB",X"2A",X"ED",X"53",X"D4",X"40",X"4F",X"11",
		X"08",X"00",X"DD",X"19",X"05",X"C2",X"E5",X"07",X"79",X"FE",X"FF",X"20",X"06",X"21",X"00",X"00",
		X"22",X"D4",X"40",X"CD",X"C2",X"15",X"FE",X"50",X"D2",X"61",X"08",X"79",X"FE",X"08",X"DC",X"65",
		X"08",X"CD",X"81",X"07",X"C9",X"DD",X"21",X"D2",X"41",X"06",X"06",X"11",X"06",X"00",X"DD",X"7E",
		X"01",X"FE",X"FF",X"28",X"05",X"DD",X"19",X"10",X"F5",X"C9",X"3E",X"03",X"CD",X"F5",X"10",X"DD",
		X"E5",X"2A",X"16",X"40",X"11",X"00",X"04",X"19",X"CB",X"3C",X"CB",X"1D",X"CD",X"C2",X"15",X"E6",
		X"60",X"C6",X"10",X"5F",X"16",X"00",X"19",X"E5",X"11",X"1C",X"00",X"01",X"0C",X"02",X"D9",X"D1",
		X"2A",X"CE",X"40",X"CD",X"08",X"09",X"69",X"ED",X"43",X"10",X"40",X"E5",X"DD",X"77",X"02",X"11",
		X"1C",X"00",X"2A",X"D0",X"40",X"CD",X"08",X"09",X"E1",X"26",X"08",X"DD",X"77",X"04",X"DD",X"BE",
		X"02",X"30",X"02",X"DD",X"7E",X"02",X"3C",X"DD",X"77",X"05",X"DD",X"36",X"03",X"00",X"D9",X"DD",
		X"7E",X"04",X"DD",X"BE",X"02",X"38",X"10",X"DD",X"7E",X"04",X"CB",X"3F",X"DD",X"BE",X"02",X"0E",
		X"34",X"30",X"02",X"0E",X"35",X"18",X"02",X"0E",X"36",X"3A",X"10",X"40",X"CB",X"7F",X"79",X"28",
		X"02",X"C6",X"04",X"4F",X"CD",X"4B",X"15",X"2A",X"24",X"40",X"DD",X"E1",X"DD",X"75",X"00",X"DD",
		X"74",X"01",X"C8",X"DD",X"36",X"01",X"FF",X"C9",X"B7",X"ED",X"52",X"4C",X"F2",X"14",X"09",X"19",
		X"EB",X"B7",X"ED",X"52",X"29",X"29",X"29",X"29",X"29",X"00",X"CB",X"11",X"9F",X"87",X"3C",X"87",
		X"87",X"87",X"4F",X"7C",X"C9",X"DD",X"21",X"CE",X"40",X"06",X"0A",X"AF",X"32",X"08",X"40",X"DD",
		X"7E",X"05",X"FE",X"FF",X"CA",X"47",X"09",X"21",X"08",X"40",X"34",X"3A",X"1E",X"40",X"90",X"E6",
		X"01",X"C2",X"47",X"09",X"CD",X"51",X"09",X"11",X"08",X"00",X"DD",X"19",X"05",X"C2",X"2F",X"09",
		X"C9",X"DD",X"7E",X"06",X"CD",X"4E",X"13",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"19",X"7C",X"E6",
		X"07",X"67",X"DD",X"75",X"00",X"DD",X"74",X"01",X"DD",X"7E",X"07",X"CD",X"4E",X"13",X"DD",X"6E",
		X"02",X"26",X"00",X"19",X"DD",X"7E",X"05",X"B7",X"20",X"09",X"7D",X"FE",X"C8",X"30",X"08",X"FE",
		X"38",X"38",X"04",X"DD",X"75",X"02",X"C9",X"DD",X"36",X"07",X"00",X"C9",X"21",X"0B",X"40",X"7E",
		X"B7",X"CA",X"98",X"09",X"35",X"CD",X"F6",X"09",X"3A",X"06",X"40",X"CB",X"7F",X"C0",X"2A",X"16",
		X"40",X"11",X"00",X"FC",X"19",X"29",X"29",X"29",X"29",X"7C",X"32",X"56",X"40",X"2A",X"16",X"40",
		X"CB",X"3C",X"CB",X"1D",X"7D",X"ED",X"44",X"32",X"0C",X"40",X"DD",X"21",X"CE",X"40",X"CD",X"67",
		X"13",X"11",X"3C",X"00",X"B7",X"ED",X"52",X"38",X"08",X"19",X"11",X"C4",X"00",X"B7",X"ED",X"52",
		X"D8",X"ED",X"5B",X"16",X"40",X"4D",X"19",X"22",X"16",X"40",X"3A",X"01",X"40",X"91",X"32",X"01",
		X"40",X"2A",X"16",X"40",X"11",X"70",X"00",X"CB",X"79",X"28",X"03",X"11",X"90",X"FF",X"19",X"CD",
		X"9B",X"13",X"CD",X"F6",X"09",X"C9",X"21",X"57",X"40",X"36",X"05",X"23",X"23",X"23",X"3A",X"0B",
		X"40",X"E6",X"07",X"4F",X"DD",X"E5",X"DD",X"2A",X"26",X"40",X"DD",X"7E",X"06",X"32",X"51",X"40",
		X"32",X"53",X"40",X"32",X"55",X"40",X"DD",X"E1",X"06",X"19",X"3A",X"01",X"40",X"81",X"77",X"23",
		X"71",X"23",X"10",X"FA",X"3E",X"05",X"06",X"04",X"21",X"85",X"40",X"77",X"23",X"23",X"10",X"FB",
		X"3A",X"0C",X"40",X"32",X"86",X"40",X"32",X"88",X"40",X"C9",X"3A",X"1E",X"40",X"E6",X"0F",X"C0",
		X"DD",X"2A",X"0E",X"40",X"CD",X"4C",X"0A",X"DD",X"22",X"0E",X"40",X"C9",X"DD",X"7E",X"00",X"FE",
		X"01",X"CA",X"6B",X"0A",X"FE",X"02",X"CA",X"7D",X"0A",X"FE",X"03",X"CA",X"DD",X"0A",X"FE",X"04",
		X"CA",X"ED",X"0A",X"FE",X"05",X"CA",X"25",X"0B",X"DD",X"23",X"C9",X"21",X"05",X"40",X"DD",X"7E",
		X"01",X"BE",X"28",X"02",X"34",X"C9",X"DD",X"23",X"DD",X"23",X"36",X"00",X"C9",X"DD",X"7E",X"05",
		X"B7",X"20",X"17",X"3A",X"CF",X"40",X"FE",X"04",X"3E",X"FF",X"38",X"02",X"3E",X"01",X"FD",X"2A",
		X"26",X"40",X"DD",X"CB",X"06",X"46",X"28",X"02",X"ED",X"44",X"32",X"04",X"40",X"CB",X"7F",X"DD",
		X"7E",X"06",X"28",X"02",X"ED",X"44",X"6F",X"26",X"00",X"29",X"29",X"29",X"DD",X"5E",X"07",X"DD",
		X"4E",X"02",X"DD",X"46",X"01",X"D9",X"2A",X"04",X"40",X"FD",X"2A",X"26",X"40",X"FD",X"7E",X"06",
		X"FE",X"03",X"38",X"02",X"3E",X"02",X"DD",X"86",X"03",X"47",X"04",X"05",X"28",X"03",X"29",X"18",
		X"FA",X"26",X"00",X"D9",X"CD",X"37",X"15",X"11",X"08",X"00",X"DD",X"19",X"C9",X"2A",X"0E",X"40",
		X"FD",X"2A",X"26",X"40",X"FD",X"75",X"04",X"FD",X"74",X"05",X"DD",X"23",X"C9",X"DD",X"21",X"76",
		X"1A",X"FD",X"2A",X"26",X"40",X"FD",X"34",X"06",X"DD",X"E5",X"CD",X"A4",X"10",X"DD",X"21",X"0D",
		X"0B",X"CD",X"7B",X"11",X"CD",X"A6",X"12",X"CD",X"1D",X"05",X"DD",X"E1",X"C9",X"82",X"53",X"54",
		X"45",X"4D",X"50",X"4F",X"52",X"41",X"52",X"59",X"20",X"43",X"45",X"41",X"53",X"45",X"46",X"49",
		X"52",X"45",X"24",X"FF",X"FF",X"3A",X"08",X"40",X"DD",X"BE",X"01",X"D0",X"DD",X"23",X"DD",X"23",
		X"C9",X"CD",X"38",X"0B",X"CD",X"64",X"0B",X"C9",X"DD",X"21",X"1E",X"41",X"06",X"14",X"78",X"90",
		X"CD",X"99",X"0B",X"20",X"17",X"DD",X"7E",X"05",X"FE",X"FF",X"28",X"10",X"DD",X"7E",X"08",X"FE",
		X"FF",X"28",X"09",X"CD",X"F3",X"0B",X"20",X"04",X"DD",X"7E",X"08",X"77",X"11",X"09",X"00",X"DD",
		X"19",X"10",X"DB",X"C9",X"DD",X"21",X"1E",X"41",X"06",X"14",X"78",X"CD",X"99",X"0B",X"20",X"21",
		X"DD",X"7E",X"05",X"FE",X"FF",X"28",X"1A",X"CD",X"A9",X"0B",X"DD",X"7E",X"05",X"3C",X"28",X"11",
		X"CD",X"F3",X"0B",X"20",X"0C",X"7E",X"DD",X"77",X"08",X"DD",X"7E",X"04",X"FE",X"FF",X"28",X"01",
		X"77",X"11",X"09",X"00",X"DD",X"19",X"10",X"D2",X"C9",X"4F",X"DD",X"7E",X"05",X"E6",X"7E",X"FE",
		X"02",X"C8",X"3A",X"1E",X"40",X"91",X"E6",X"03",X"C9",X"DD",X"7E",X"05",X"E6",X"7F",X"FE",X"02",
		X"28",X"0F",X"FE",X"03",X"C8",X"FE",X"04",X"28",X"10",X"FE",X"05",X"28",X"11",X"CD",X"51",X"09",
		X"C9",X"CD",X"51",X"09",X"DD",X"36",X"05",X"03",X"C9",X"DD",X"36",X"05",X"FF",X"C9",X"DD",X"36",
		X"06",X"00",X"DD",X"36",X"07",X"00",X"DD",X"7E",X"03",X"FE",X"10",X"28",X"0E",X"DD",X"34",X"03",
		X"E6",X"0C",X"C6",X"E0",X"DD",X"77",X"04",X"CD",X"5E",X"14",X"C9",X"DD",X"36",X"05",X"04",X"CD",
		X"7C",X"14",X"C9",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"CD",X"AE",X"15",X"C0",X"DD",X"7E",X"02",
		X"ED",X"44",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"5F",X"16",X"50",X"19",X"AF",X"C9",X"DD",X"21",
		X"CE",X"40",X"06",X"0A",X"DD",X"7E",X"05",X"C5",X"CD",X"24",X"0C",X"C1",X"11",X"08",X"00",X"DD",
		X"19",X"10",X"F1",X"C9",X"FE",X"FF",X"C8",X"B7",X"CA",X"4A",X"0C",X"FE",X"01",X"CA",X"4F",X"0C",
		X"FE",X"02",X"CA",X"6A",X"0C",X"FE",X"03",X"CA",X"B4",X"0C",X"FE",X"04",X"CA",X"D3",X"0C",X"FE",
		X"05",X"CA",X"31",X"0D",X"FE",X"58",X"CA",X"D2",X"0D",X"C9",X"DD",X"36",X"03",X"00",X"C9",X"CD",
		X"FA",X"0D",X"CD",X"C2",X"15",X"FE",X"01",X"21",X"13",X"1C",X"3E",X"00",X"DC",X"F5",X"10",X"CD",
		X"C2",X"15",X"FE",X"1E",X"DC",X"49",X"0E",X"C3",X"2E",X"0E",X"CD",X"C2",X"15",X"FE",X"01",X"3E",
		X"00",X"21",X"23",X"1C",X"DC",X"F5",X"10",X"DD",X"36",X"03",X"02",X"CD",X"FA",X"0D",X"CD",X"C2",
		X"15",X"FE",X"02",X"30",X"14",X"DD",X"7E",X"06",X"CD",X"53",X"13",X"4F",X"DD",X"7E",X"01",X"FE",
		X"04",X"79",X"38",X"02",X"ED",X"44",X"DD",X"77",X"06",X"FD",X"2A",X"26",X"40",X"FD",X"7E",X"06",
		X"0E",X"02",X"38",X"08",X"FE",X"02",X"0E",X"08",X"38",X"02",X"0E",X"14",X"CD",X"C2",X"15",X"B9",
		X"D0",X"C3",X"3A",X"0E",X"DD",X"36",X"03",X"02",X"CD",X"FA",X"0D",X"CD",X"C2",X"15",X"FE",X"01",
		X"21",X"33",X"1C",X"3E",X"00",X"DC",X"F5",X"10",X"CD",X"C2",X"15",X"FE",X"1E",X"DC",X"49",X"0E",
		X"C3",X"3A",X"0E",X"3E",X"06",X"CD",X"F5",X"10",X"CD",X"FA",X"0D",X"DD",X"6E",X"00",X"DD",X"66",
		X"01",X"CD",X"7B",X"13",X"B7",X"28",X"04",X"DD",X"36",X"07",X"FC",X"C6",X"30",X"DD",X"BE",X"02",
		X"D8",X"DD",X"36",X"06",X"00",X"DD",X"36",X"07",X"04",X"DD",X"36",X"05",X"58",X"DD",X"6E",X"00",
		X"DD",X"66",X"01",X"11",X"C0",X"FF",X"19",X"06",X"10",X"C5",X"E5",X"CD",X"7B",X"13",X"7D",X"B4",
		X"28",X"10",X"7E",X"CB",X"3F",X"D6",X"02",X"CB",X"7F",X"28",X"01",X"AF",X"77",X"E1",X"E5",X"CD",
		X"9B",X"13",X"E1",X"11",X"08",X"00",X"19",X"C1",X"10",X"DF",X"C9",X"3E",X"15",X"32",X"15",X"40",
		X"C9",X"3E",X"04",X"CD",X"F5",X"10",X"CD",X"FA",X"0D",X"CD",X"C2",X"15",X"E6",X"1F",X"20",X"2E",
		X"FD",X"2A",X"26",X"40",X"FD",X"7E",X"06",X"FE",X"03",X"0E",X"02",X"30",X"01",X"4F",X"0C",X"0C",
		X"0C",X"DD",X"7E",X"01",X"FE",X"04",X"30",X"0B",X"DD",X"7E",X"06",X"B9",X"28",X"10",X"DD",X"34",
		X"06",X"18",X"0B",X"DD",X"7E",X"06",X"ED",X"44",X"B9",X"28",X"03",X"DD",X"35",X"06",X"CD",X"C2",
		X"15",X"E6",X"28",X"DC",X"49",X"0E",X"2A",X"12",X"40",X"7C",X"B5",X"C0",X"FD",X"2A",X"26",X"40",
		X"FD",X"7E",X"06",X"FE",X"01",X"0E",X"28",X"38",X"08",X"0E",X"50",X"FE",X"02",X"38",X"02",X"0E",
		X"78",X"CD",X"C2",X"15",X"B9",X"D0",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"E5",X"CD",X"7B",X"13",
		X"7D",X"B4",X"28",X"27",X"7E",X"B7",X"28",X"23",X"3D",X"30",X"02",X"3E",X"00",X"77",X"E1",X"22",
		X"12",X"40",X"3E",X"0A",X"32",X"0B",X"40",X"CD",X"F3",X"0B",X"C0",X"2C",X"7D",X"E6",X"1F",X"FE",
		X"1A",X"D0",X"7E",X"FE",X"90",X"C0",X"36",X"95",X"23",X"18",X"F7",X"E1",X"C9",X"DD",X"36",X"05",
		X"FF",X"C9",X"DD",X"36",X"07",X"FF",X"DD",X"7E",X"02",X"FE",X"1E",X"38",X"18",X"DD",X"7E",X"03",
		X"FE",X"20",X"28",X"11",X"E6",X"03",X"C6",X"3C",X"DD",X"77",X"04",X"CD",X"C2",X"15",X"E6",X"01",
		X"C0",X"DD",X"34",X"03",X"C9",X"DD",X"36",X"05",X"FF",X"C9",X"3A",X"1E",X"40",X"3C",X"E6",X"07",
		X"C0",X"DD",X"7E",X"05",X"FE",X"01",X"DD",X"7E",X"06",X"28",X"01",X"2F",X"E6",X"80",X"4F",X"DD",
		X"7E",X"04",X"E6",X"7F",X"B1",X"DD",X"77",X"04",X"DD",X"7E",X"01",X"B7",X"20",X"08",X"DD",X"7E",
		X"00",X"FE",X"3F",X"DA",X"2A",X"0E",X"CD",X"78",X"0E",X"C9",X"E1",X"C3",X"CD",X"0D",X"DD",X"6E",
		X"00",X"DD",X"66",X"01",X"CD",X"7B",X"13",X"FE",X"03",X"D8",X"DD",X"6E",X"00",X"DD",X"66",X"01",
		X"CD",X"7B",X"13",X"B7",X"C8",X"CD",X"CD",X"0E",X"C9",X"2A",X"CE",X"40",X"DD",X"5E",X"00",X"DD",
		X"56",X"01",X"CD",X"08",X"09",X"FE",X"08",X"D0",X"3A",X"D0",X"40",X"DD",X"BE",X"02",X"38",X"0C",
		X"DD",X"7E",X"02",X"FE",X"3C",X"38",X"05",X"DD",X"36",X"07",X"FD",X"C9",X"DD",X"7E",X"02",X"FE",
		X"BE",X"30",X"ED",X"DD",X"36",X"07",X"03",X"C9",X"DD",X"7E",X"01",X"FE",X"04",X"30",X"05",X"3E",
		X"08",X"DD",X"96",X"01",X"FE",X"04",X"28",X"21",X"FE",X"05",X"28",X"30",X"DD",X"7E",X"05",X"FE",
		X"01",X"28",X"11",X"FE",X"04",X"28",X"0D",X"3A",X"1E",X"40",X"CB",X"77",X"3E",X"01",X"28",X"02",
		X"3E",X"FF",X"18",X"01",X"AF",X"DD",X"77",X"07",X"C9",X"DD",X"7E",X"02",X"FE",X"50",X"38",X"DC",
		X"DD",X"7E",X"06",X"CD",X"53",X"13",X"ED",X"44",X"DD",X"77",X"07",X"C9",X"CD",X"C2",X"15",X"E6",
		X"3F",X"C6",X"80",X"DD",X"BE",X"02",X"38",X"C4",X"DD",X"36",X"07",X"01",X"C9",X"DD",X"7E",X"02",
		X"FE",X"C8",X"D0",X"3E",X"01",X"CD",X"F5",X"10",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"DD",X"5E",
		X"02",X"16",X"00",X"01",X"3C",X"01",X"D9",X"21",X"00",X"F8",X"D9",X"CD",X"57",X"15",X"C9",X"DD",
		X"21",X"D2",X"41",X"06",X"06",X"DD",X"7E",X"01",X"FE",X"FF",X"CA",X"46",X"0F",X"DD",X"6E",X"00",
		X"DD",X"66",X"01",X"E5",X"FD",X"E1",X"FD",X"7E",X"05",X"FE",X"03",X"C2",X"46",X"0F",X"DD",X"35",
		X"05",X"CA",X"33",X"0F",X"DD",X"7E",X"02",X"DD",X"BE",X"04",X"38",X"05",X"CD",X"4E",X"0F",X"18",
		X"03",X"CD",X"6E",X"0F",X"0E",X"01",X"CD",X"60",X"13",X"CD",X"BB",X"14",X"CD",X"60",X"13",X"20",
		X"02",X"18",X"13",X"FD",X"36",X"05",X"05",X"DD",X"36",X"01",X"FF",X"CD",X"60",X"13",X"0E",X"03",
		X"CD",X"BB",X"14",X"CD",X"60",X"13",X"11",X"06",X"00",X"DD",X"19",X"10",X"A8",X"C9",X"FD",X"36",
		X"07",X"00",X"FD",X"36",X"05",X"02",X"DD",X"7E",X"03",X"DD",X"86",X"04",X"DD",X"96",X"02",X"30",
		X"07",X"DD",X"86",X"02",X"DD",X"77",X"03",X"C9",X"FD",X"36",X"07",X"08",X"18",X"F6",X"FD",X"36",
		X"06",X"00",X"FD",X"36",X"05",X"02",X"DD",X"7E",X"03",X"DD",X"86",X"02",X"DD",X"96",X"04",X"30",
		X"05",X"DD",X"86",X"04",X"18",X"DE",X"0E",X"08",X"FD",X"CB",X"04",X"56",X"20",X"02",X"0E",X"F8",
		X"FD",X"71",X"06",X"18",X"CF",X"DD",X"21",X"1E",X"41",X"06",X"14",X"DD",X"7E",X"05",X"C5",X"DD",
		X"E5",X"CD",X"AF",X"0F",X"DD",X"E1",X"C1",X"11",X"09",X"00",X"DD",X"19",X"10",X"ED",X"C9",X"FE",
		X"FF",X"C8",X"FE",X"01",X"28",X"01",X"C9",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"CD",X"7B",X"13",
		X"87",X"87",X"87",X"C6",X"40",X"DD",X"BE",X"02",X"D8",X"DD",X"36",X"05",X"FF",X"CD",X"F3",X"0B",
		X"20",X"02",X"36",X"10",X"3E",X"1E",X"32",X"0B",X"40",X"3E",X"02",X"CD",X"F5",X"10",X"DD",X"6E",
		X"00",X"DD",X"66",X"01",X"11",X"F0",X"FF",X"19",X"0E",X"00",X"CD",X"01",X"10",X"0E",X"01",X"CD",
		X"01",X"10",X"0E",X"02",X"CD",X"01",X"10",X"0E",X"01",X"CD",X"01",X"10",X"0E",X"00",X"CD",X"01",
		X"10",X"E5",X"22",X"1C",X"40",X"D5",X"C5",X"CD",X"7B",X"13",X"C1",X"7D",X"B4",X"28",X"07",X"7E",
		X"91",X"30",X"02",X"3E",X"00",X"77",X"2A",X"1C",X"40",X"CD",X"9B",X"13",X"D1",X"E1",X"11",X"08",
		X"00",X"19",X"C9",X"3A",X"06",X"40",X"B7",X"C2",X"55",X"10",X"CD",X"C2",X"15",X"E6",X"0F",X"C0",
		X"3A",X"1F",X"40",X"CB",X"47",X"21",X"F6",X"41",X"11",X"01",X"00",X"20",X"06",X"21",X"15",X"42",
		X"11",X"FF",X"FF",X"01",X"00",X"20",X"7E",X"B7",X"20",X"05",X"19",X"10",X"F9",X"AF",X"C9",X"22",
		X"28",X"40",X"F6",X"FF",X"C9",X"AF",X"C9",X"3E",X"FF",X"32",X"0B",X"40",X"21",X"06",X"40",X"34",
		X"F2",X"95",X"10",X"3E",X"FF",X"32",X"D3",X"40",X"AF",X"32",X"0B",X"40",X"CD",X"F6",X"09",X"2A",
		X"16",X"40",X"7C",X"FE",X"04",X"20",X"04",X"7D",X"FE",X"08",X"D8",X"3E",X"80",X"32",X"06",X"40",
		X"F5",X"3E",X"00",X"21",X"43",X"1C",X"CD",X"F5",X"10",X"F1",X"21",X"FC",X"FF",X"30",X"03",X"21",
		X"04",X"00",X"C3",X"D1",X"09",X"7E",X"FE",X"01",X"C0",X"CD",X"76",X"06",X"DD",X"21",X"74",X"19",
		X"CD",X"7B",X"11",X"C9",X"CD",X"7B",X"00",X"06",X"04",X"21",X"00",X"50",X"36",X"10",X"2C",X"20",
		X"FB",X"24",X"10",X"F8",X"21",X"00",X"00",X"22",X"20",X"42",X"3E",X"FF",X"32",X"00",X"78",X"AF",
		X"32",X"03",X"68",X"32",X"05",X"68",X"32",X"04",X"70",X"32",X"0C",X"40",X"21",X"4E",X"40",X"06",
		X"80",X"36",X"00",X"23",X"10",X"FB",X"AF",X"32",X"01",X"40",X"3E",X"07",X"32",X"4F",X"40",X"32",
		X"8D",X"40",X"DD",X"21",X"D2",X"18",X"CD",X"7B",X"11",X"CD",X"F0",X"11",X"C9",X"3E",X"F2",X"C6",
		X"23",X"FD",X"77",X"0C",X"C9",X"DD",X"E5",X"CD",X"FD",X"10",X"DD",X"E1",X"C9",X"DD",X"21",X"20",
		X"42",X"FE",X"00",X"CA",X"25",X"11",X"FE",X"01",X"CA",X"36",X"11",X"FE",X"02",X"CA",X"44",X"11",
		X"FE",X"03",X"CA",X"4D",X"11",X"FE",X"04",X"CA",X"56",X"11",X"FE",X"05",X"CA",X"64",X"11",X"FE",
		X"06",X"CA",X"6D",X"11",X"C9",X"DD",X"CB",X"00",X"46",X"C0",X"22",X"22",X"42",X"DD",X"36",X"04",
		X"14",X"DD",X"CB",X"00",X"C6",X"C9",X"DD",X"CB",X"00",X"4E",X"C0",X"DD",X"CB",X"00",X"CE",X"DD",
		X"36",X"05",X"50",X"C9",X"DD",X"CB",X"00",X"D6",X"DD",X"36",X"06",X"78",X"C9",X"DD",X"CB",X"00",
		X"DE",X"DD",X"36",X"07",X"14",X"C9",X"DD",X"CB",X"00",X"66",X"C0",X"DD",X"36",X"08",X"80",X"DD",
		X"CB",X"00",X"E6",X"C9",X"DD",X"36",X"09",X"00",X"DD",X"CB",X"00",X"EE",X"C9",X"DD",X"CB",X"00",
		X"76",X"C0",X"DD",X"36",X"0A",X"00",X"DD",X"CB",X"00",X"F6",X"C9",X"DD",X"6E",X"00",X"DD",X"66",
		X"01",X"DD",X"23",X"DD",X"23",X"11",X"E0",X"FF",X"24",X"C8",X"25",X"DD",X"7E",X"00",X"FE",X"80",
		X"D2",X"B2",X"11",X"DD",X"23",X"FE",X"20",X"0E",X"10",X"28",X"03",X"D6",X"30",X"4F",X"71",X"19",
		X"7C",X"E6",X"03",X"C6",X"50",X"67",X"DD",X"7E",X"00",X"FE",X"24",X"20",X"DE",X"DD",X"23",X"C3",
		X"7B",X"11",X"DD",X"23",X"D6",X"B0",X"87",X"87",X"4F",X"C6",X"02",X"77",X"23",X"3C",X"77",X"2B",
		X"19",X"23",X"D6",X"02",X"77",X"2B",X"18",X"D6",X"7E",X"1F",X"1F",X"1F",X"1F",X"CD",X"D8",X"11",
		X"7E",X"CD",X"D8",X"11",X"2B",X"10",X"F1",X"C9",X"11",X"E0",X"FF",X"FD",X"19",X"E6",X"0F",X"FE",
		X"0A",X"38",X"02",X"C6",X"07",X"B7",X"20",X"02",X"0D",X"F0",X"0E",X"FF",X"FD",X"77",X"20",X"C9",
		X"21",X"34",X"40",X"01",X"01",X"03",X"FD",X"21",X"40",X"53",X"CD",X"C8",X"11",X"21",X"4C",X"40",
		X"01",X"01",X"03",X"FD",X"21",X"20",X"52",X"CD",X"C8",X"11",X"21",X"3C",X"40",X"01",X"01",X"03",
		X"FD",X"21",X"E0",X"50",X"CD",X"C8",X"11",X"DD",X"2A",X"26",X"40",X"21",X"DF",X"51",X"DD",X"7E",
		X"07",X"3D",X"06",X"05",X"11",X"C0",X"FF",X"3D",X"FA",X"31",X"12",X"36",X"2C",X"05",X"19",X"18",
		X"F6",X"05",X"FA",X"3A",X"12",X"36",X"10",X"19",X"18",X"F7",X"21",X"15",X"40",X"01",X"FF",X"01",
		X"FD",X"21",X"7F",X"52",X"CD",X"C8",X"11",X"7E",X"FE",X"50",X"3E",X"10",X"38",X"02",X"3E",X"2D",
		X"FD",X"77",X"00",X"C9",X"DD",X"E5",X"FD",X"E5",X"E5",X"D5",X"C5",X"6F",X"26",X"00",X"29",X"11",
		X"16",X"42",X"19",X"7E",X"23",X"4E",X"2A",X"26",X"40",X"86",X"27",X"77",X"23",X"79",X"8E",X"27",
		X"77",X"23",X"06",X"02",X"3E",X"00",X"8E",X"27",X"77",X"23",X"10",X"F8",X"CD",X"8A",X"12",X"CD",
		X"F0",X"11",X"C1",X"D1",X"E1",X"FD",X"E1",X"DD",X"E1",X"C9",X"2A",X"26",X"40",X"23",X"23",X"23",
		X"11",X"4D",X"40",X"06",X"04",X"1A",X"BE",X"20",X"05",X"2B",X"1B",X"10",X"F8",X"C9",X"D0",X"7E",
		X"12",X"2B",X"1B",X"10",X"FA",X"C9",X"DD",X"E5",X"DD",X"21",X"F7",X"18",X"CD",X"7B",X"11",X"21",
		X"6C",X"1A",X"11",X"16",X"42",X"01",X"0A",X"00",X"ED",X"B0",X"DD",X"2A",X"26",X"40",X"DD",X"4E",
		X"06",X"06",X"05",X"FD",X"21",X"4A",X"51",X"DD",X"21",X"16",X"42",X"FD",X"E5",X"C5",X"DD",X"6E",
		X"00",X"DD",X"66",X"01",X"41",X"05",X"FA",X"EB",X"12",X"7D",X"87",X"27",X"6F",X"7C",X"8F",X"27",
		X"67",X"38",X"0E",X"DD",X"75",X"00",X"DD",X"74",X"01",X"18",X"EA",X"DD",X"75",X"00",X"DD",X"74",
		X"01",X"DD",X"E5",X"E1",X"23",X"01",X"00",X"02",X"CD",X"C8",X"11",X"C1",X"FD",X"E1",X"FD",X"23",
		X"FD",X"23",X"FD",X"23",X"DD",X"23",X"DD",X"23",X"10",X"C1",X"06",X"C8",X"CD",X"7B",X"00",X"78",
		X"CB",X"3F",X"CB",X"3F",X"E6",X"04",X"32",X"53",X"40",X"32",X"55",X"40",X"10",X"EE",X"DD",X"E1",
		X"C9",X"2F",X"4F",X"2F",X"DD",X"A6",X"03",X"DD",X"71",X"03",X"2F",X"DD",X"77",X"00",X"DD",X"23",
		X"C9",X"DD",X"CB",X"00",X"7E",X"21",X"2C",X"40",X"20",X"03",X"21",X"2F",X"40",X"DD",X"5E",X"00",
		X"16",X"00",X"CB",X"BB",X"19",X"7E",X"DD",X"A6",X"01",X"DD",X"23",X"DD",X"23",X"C9",X"5F",X"17",
		X"9F",X"57",X"C9",X"B7",X"F0",X"ED",X"44",X"C9",X"B7",X"C8",X"3E",X"01",X"F0",X"3E",X"FF",X"C9",
		X"DD",X"E5",X"FD",X"E3",X"DD",X"E1",X"C9",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"ED",X"5B",X"16",
		X"40",X"B7",X"ED",X"52",X"11",X"80",X"00",X"19",X"7C",X"B7",X"C9",X"11",X"80",X"FC",X"19",X"7C",
		X"B7",X"20",X"14",X"CB",X"3C",X"CB",X"1D",X"CB",X"3C",X"CB",X"1D",X"CB",X"3C",X"CB",X"1D",X"11",
		X"F6",X"41",X"19",X"F6",X"FF",X"7E",X"C9",X"AF",X"6F",X"67",X"C9",X"CD",X"AE",X"15",X"C0",X"11",
		X"1A",X"50",X"19",X"22",X"1A",X"40",X"E5",X"06",X"15",X"36",X"90",X"2B",X"10",X"FB",X"2A",X"18",
		X"40",X"11",X"F8",X"FF",X"19",X"CD",X"7B",X"13",X"4F",X"C5",X"2A",X"18",X"40",X"11",X"08",X"00",
		X"19",X"CD",X"7B",X"13",X"C1",X"47",X"C5",X"2A",X"18",X"40",X"CD",X"7B",X"13",X"C1",X"E1",X"5F",
		X"B7",X"28",X"08",X"E6",X"7F",X"36",X"10",X"2B",X"3D",X"20",X"FA",X"7B",X"B1",X"B0",X"28",X"11",
		X"79",X"93",X"CD",X"55",X"14",X"87",X"87",X"57",X"78",X"93",X"CD",X"55",X"14",X"B2",X"C6",X"80",
		X"77",X"2A",X"1A",X"40",X"3A",X"18",X"40",X"E6",X"38",X"3E",X"97",X"28",X"02",X"3E",X"90",X"23",
		X"77",X"23",X"23",X"23",X"36",X"90",X"2A",X"16",X"40",X"11",X"00",X"04",X"19",X"CB",X"3C",X"CB",
		X"1D",X"EB",X"2A",X"18",X"40",X"B7",X"ED",X"52",X"5D",X"54",X"7C",X"B7",X"01",X"33",X"1A",X"20",
		X"13",X"CB",X"7D",X"C2",X"34",X"14",X"7D",X"1F",X"1F",X"E6",X"1E",X"6F",X"26",X"00",X"01",X"13",
		X"1A",X"09",X"44",X"4D",X"3A",X"18",X"40",X"2F",X"2A",X"16",X"40",X"CB",X"3C",X"CB",X"1D",X"85",
		X"C6",X"80",X"E6",X"F8",X"6F",X"26",X"00",X"29",X"29",X"11",X"1C",X"50",X"19",X"EB",X"60",X"69",
		X"ED",X"A0",X"ED",X"A0",X"C9",X"3E",X"01",X"C8",X"3E",X"02",X"D0",X"3E",X"00",X"C9",X"DD",X"E5",
		X"4F",X"CD",X"70",X"14",X"C2",X"B3",X"14",X"CD",X"8D",X"14",X"20",X"01",X"71",X"0C",X"18",X"F7",
		X"C5",X"CD",X"F3",X"0B",X"C1",X"C0",X"DD",X"21",X"B6",X"14",X"AF",X"C9",X"DD",X"E5",X"CD",X"70",
		X"14",X"20",X"30",X"CD",X"8D",X"14",X"20",X"02",X"36",X"90",X"0C",X"18",X"F6",X"DD",X"7E",X"00",
		X"FE",X"80",X"28",X"1E",X"DD",X"23",X"D5",X"CD",X"4E",X"13",X"19",X"D1",X"7C",X"E6",X"03",X"C6",
		X"50",X"67",X"7E",X"FE",X"90",X"C8",X"FE",X"34",X"D8",X"FE",X"3C",X"38",X"03",X"FE",X"E0",X"D8",
		X"BF",X"C9",X"E1",X"DD",X"E1",X"C9",X"00",X"01",X"1F",X"01",X"80",X"FD",X"E5",X"C5",X"06",X"09",
		X"FD",X"21",X"D6",X"40",X"1E",X"00",X"D5",X"FD",X"7E",X"05",X"FE",X"FF",X"CA",X"29",X"15",X"DD",
		X"6E",X"00",X"DD",X"66",X"01",X"FD",X"5E",X"00",X"FD",X"56",X"01",X"C5",X"CD",X"08",X"09",X"C1",
		X"B9",X"D2",X"29",X"15",X"DD",X"6E",X"02",X"26",X"00",X"FD",X"5E",X"02",X"54",X"C5",X"CD",X"08",
		X"09",X"C1",X"B9",X"30",X"34",X"D1",X"1C",X"D5",X"FD",X"36",X"03",X"00",X"FD",X"7E",X"05",X"FD",
		X"36",X"05",X"58",X"FE",X"01",X"1E",X"01",X"28",X"17",X"1D",X"FE",X"02",X"28",X"12",X"FE",X"03",
		X"1E",X"02",X"28",X"0C",X"1C",X"FE",X"04",X"28",X"07",X"1C",X"FE",X"05",X"28",X"02",X"18",X"09",
		X"7B",X"CD",X"54",X"12",X"3E",X"05",X"CD",X"F5",X"10",X"11",X"08",X"00",X"FD",X"19",X"D1",X"10",
		X"95",X"7B",X"B7",X"C1",X"FD",X"E1",X"C9",X"DD",X"E5",X"D5",X"C5",X"DD",X"21",X"D6",X"40",X"06",
		X"09",X"11",X"08",X"00",X"CD",X"71",X"15",X"DD",X"E1",X"AF",X"C9",X"DD",X"E5",X"D5",X"C5",X"DD",
		X"21",X"1E",X"41",X"06",X"0A",X"18",X"0A",X"DD",X"E5",X"D5",X"C5",X"DD",X"21",X"78",X"41",X"06",
		X"0A",X"11",X"09",X"00",X"CD",X"71",X"15",X"D9",X"DD",X"36",X"08",X"FF",X"D9",X"DD",X"E1",X"AF",
		X"C9",X"E3",X"22",X"20",X"40",X"DD",X"7E",X"05",X"FE",X"FF",X"28",X"0C",X"DD",X"19",X"10",X"F5",
		X"E1",X"C1",X"D1",X"DD",X"E1",X"F6",X"FF",X"C9",X"E1",X"C1",X"D1",X"DD",X"22",X"24",X"40",X"DD",
		X"75",X"00",X"DD",X"74",X"01",X"DD",X"73",X"02",X"DD",X"36",X"03",X"00",X"DD",X"71",X"04",X"DD",
		X"70",X"05",X"D9",X"DD",X"75",X"06",X"DD",X"74",X"07",X"D9",X"2A",X"20",X"40",X"E9",X"22",X"18",
		X"40",X"CD",X"6D",X"13",X"C0",X"3A",X"18",X"40",X"2F",X"E6",X"F8",X"6F",X"26",X"00",X"29",X"29",
		X"AF",X"C9",X"E5",X"ED",X"5F",X"2A",X"22",X"40",X"8C",X"CE",X"91",X"8E",X"67",X"8D",X"CE",X"BB",
		X"0F",X"6F",X"22",X"22",X"40",X"E1",X"C9",X"09",X"24",X"80",X"20",X"00",X"48",X"44",X"89",X"02",
		X"40",X"44",X"48",X"00",X"08",X"04",X"22",X"10",X"12",X"00",X"84",X"24",X"92",X"01",X"10",X"92",
		X"40",X"80",X"00",X"01",X"00",X"88",X"81",X"21",X"24",X"80",X"91",X"24",X"08",X"09",X"20",X"20",
		X"08",X"48",X"20",X"04",X"89",X"01",X"20",X"08",X"04",X"90",X"12",X"21",X"11",X"20",X"40",X"12",
		X"41",X"12",X"41",X"00",X"40",X"48",X"40",X"48",X"80",X"02",X"10",X"00",X"92",X"42",X"10",X"44",
		X"40",X"40",X"42",X"49",X"04",X"88",X"92",X"40",X"12",X"01",X"00",X"24",X"91",X"01",X"10",X"00",
		X"80",X"09",X"24",X"48",X"42",X"44",X"21",X"08",X"84",X"80",X"42",X"10",X"80",X"90",X"00",X"01",
		X"20",X"00",X"04",X"48",X"80",X"92",X"49",X"24",X"90",X"24",X"00",X"00",X"00",X"08",X"92",X"24",
		X"22",X"04",X"89",X"24",X"10",X"91",X"01",X"20",X"82",X"44",X"91",X"00",X"88",X"11",X"10",X"84",
		X"82",X"24",X"82",X"08",X"92",X"22",X"48",X"01",X"08",X"49",X"10",X"88",X"48",X"42",X"49",X"24",
		X"92",X"10",X"49",X"24",X"44",X"80",X"84",X"11",X"01",X"02",X"10",X"48",X"40",X"92",X"22",X"04",
		X"00",X"80",X"04",X"04",X"04",X"41",X"01",X"09",X"09",X"24",X"00",X"40",X"11",X"20",X"01",X"02",
		X"21",X"02",X"10",X"80",X"20",X"84",X"20",X"20",X"02",X"21",X"10",X"82",X"21",X"04",X"48",X"42",
		X"21",X"08",X"44",X"00",X"00",X"00",X"00",X"02",X"00",X"48",X"08",X"11",X"04",X"88",X"49",X"10",
		X"49",X"20",X"04",X"40",X"00",X"20",X"10",X"90",X"01",X"20",X"02",X"21",X"09",X"20",X"84",X"24",
		X"90",X"20",X"01",X"02",X"20",X"42",X"10",X"09",X"20",X"80",X"40",X"41",X"08",X"89",X"08",X"90",
		X"20",X"88",X"00",X"92",X"04",X"24",X"04",X"21",X"04",X"90",X"92",X"42",X"49",X"09",X"04",X"01",
		X"00",X"22",X"40",X"88",X"80",X"00",X"84",X"00",X"88",X"10",X"88",X"24",X"22",X"11",X"09",X"22",
		X"12",X"12",X"04",X"00",X"24",X"92",X"49",X"24",X"82",X"49",X"21",X"20",X"40",X"01",X"09",X"11",
		X"12",X"21",X"00",X"82",X"44",X"80",X"80",X"24",X"02",X"02",X"42",X"08",X"10",X"12",X"08",X"42",
		X"12",X"24",X"81",X"04",X"92",X"22",X"49",X"04",X"80",X"90",X"24",X"10",X"84",X"01",X"02",X"04",
		X"00",X"00",X"00",X"00",X"00",X"08",X"84",X"20",X"10",X"02",X"00",X"00",X"20",X"24",X"80",X"80",
		X"00",X"92",X"04",X"00",X"21",X"11",X"04",X"92",X"02",X"44",X"80",X"81",X"10",X"82",X"12",X"10",
		X"91",X"24",X"84",X"92",X"24",X"80",X"49",X"24",X"49",X"24",X"92",X"24",X"22",X"12",X"41",X"24",
		X"24",X"92",X"49",X"20",X"08",X"11",X"04",X"20",X"10",X"10",X"81",X"08",X"40",X"08",X"49",X"20",
		X"91",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"49",X"24",X"20",X"01",X"00",X"01",X"02",X"40",X"84",
		X"11",X"01",X"22",X"48",X"02",X"09",X"00",X"40",X"12",X"12",X"01",X"00",X"84",X"20",X"40",X"40",
		X"42",X"48",X"10",X"00",X"08",X"41",X"11",X"01",X"04",X"42",X"49",X"12",X"41",X"04",X"00",X"09",
		X"24",X"20",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"40",X"02",X"10",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AF",X"52",X"5B",X"56",X"49",X"43",X"54",X"4F",X"52",X"59",X"5B",X"24",X"11",X"53",X"43",X"4F",
		X"4D",X"53",X"4F",X"46",X"54",X"20",X"31",X"39",X"38",X"32",X"20",X"20",X"20",X"47",X"32",X"30",
		X"24",X"FF",X"FF",X"08",X"53",X"50",X"52",X"45",X"53",X"53",X"20",X"50",X"4C",X"41",X"59",X"20",
		X"42",X"55",X"54",X"54",X"4F",X"4E",X"5B",X"24",X"AC",X"52",X"4F",X"4E",X"45",X"20",X"50",X"4C",
		X"41",X"59",X"45",X"52",X"24",X"4E",X"52",X"4F",X"4E",X"4C",X"59",X"24",X"FF",X"FF",X"0E",X"53",
		X"4F",X"52",X"20",X"54",X"57",X"4F",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"53",X"24",X"FF",
		X"FF",X"4E",X"53",X"44",X"45",X"46",X"45",X"4E",X"44",X"20",X"54",X"48",X"45",X"20",X"49",X"53",
		X"4C",X"41",X"4E",X"44",X"20",X"46",X"52",X"4F",X"4D",X"24",X"D0",X"52",X"54",X"48",X"45",X"20",
		X"41",X"54",X"54",X"41",X"43",X"4B",X"49",X"4E",X"47",X"24",X"D2",X"52",X"45",X"4E",X"45",X"4D",
		X"59",X"20",X"41",X"49",X"52",X"46",X"4F",X"52",X"43",X"45",X"24",X"35",X"53",X"43",X"4F",X"4D",
		X"53",X"4F",X"46",X"54",X"20",X"31",X"39",X"38",X"32",X"20",X"20",X"20",X"47",X"32",X"30",X"24",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"A0",X"53",X"31",X"5B",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"48",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"32",X"5B",X"24",X"7F",X"53",X"43",X"52",X"45",X"44",
		X"49",X"54",X"53",X"5B",X"24",X"FF",X"FF",X"86",X"53",X"53",X"43",X"4F",X"52",X"45",X"53",X"20",
		X"4E",X"4F",X"57",X"20",X"53",X"45",X"54",X"20",X"41",X"54",X"5B",X"24",X"68",X"52",X"45",X"4E",
		X"45",X"4D",X"59",X"20",X"20",X"20",X"20",X"20",X"20",X"56",X"41",X"4C",X"55",X"45",X"24",X"8A",
		X"52",X"43",X"4F",X"50",X"54",X"45",X"52",X"53",X"24",X"8D",X"52",X"46",X"49",X"47",X"48",X"54",
		X"45",X"52",X"53",X"24",X"90",X"52",X"42",X"4F",X"4D",X"42",X"45",X"52",X"53",X"24",X"93",X"52",
		X"4D",X"49",X"53",X"53",X"49",X"4C",X"45",X"53",X"24",X"96",X"52",X"53",X"4B",X"49",X"4D",X"4D",
		X"45",X"52",X"53",X"24",X"FF",X"FF",X"42",X"52",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"4F",
		X"4E",X"45",X"24",X"FF",X"FF",X"43",X"52",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"54",X"57",
		X"4F",X"24",X"FF",X"FF",X"02",X"53",X"49",X"53",X"4C",X"41",X"4E",X"44",X"20",X"44",X"45",X"53",
		X"54",X"52",X"4F",X"59",X"45",X"44",X"24",X"FF",X"FF",X"A3",X"03",X"A4",X"03",X"A5",X"03",X"A6",
		X"03",X"A7",X"03",X"A8",X"13",X"88",X"0B",X"89",X"13",X"69",X"0B",X"6A",X"13",X"4A",X"0F",X"49",
		X"07",X"29",X"0F",X"28",X"07",X"08",X"0F",X"07",X"03",X"06",X"03",X"05",X"03",X"04",X"03",X"03",
		X"03",X"C7",X"02",X"C8",X"02",X"C9",X"02",X"CA",X"02",X"47",X"0A",X"67",X"02",X"87",X"06",X"88",
		X"02",X"89",X"02",X"8A",X"12",X"6A",X"02",X"4A",X"0E",X"C7",X"01",X"E7",X"01",X"07",X"02",X"E8",
		X"01",X"E9",X"01",X"EA",X"01",X"47",X"09",X"67",X"01",X"87",X"05",X"88",X"01",X"89",X"01",X"8A",
		X"11",X"6A",X"01",X"4A",X"0D",X"49",X"01",X"48",X"01",X"C7",X"08",X"E7",X"00",X"07",X"01",X"08",
		X"01",X"09",X"01",X"0A",X"01",X"E9",X"00",X"C8",X"00",X"EA",X"10",X"C9",X"0C",X"CA",X"08",X"47",
		X"04",X"48",X"0C",X"68",X"00",X"69",X"00",X"6A",X"00",X"87",X"08",X"88",X"10",X"FF",X"FF",X"82",
		X"8A",X"89",X"84",X"90",X"54",X"57",X"55",X"90",X"56",X"90",X"90",X"90",X"90",X"90",X"4F",X"53",
		X"50",X"90",X"51",X"90",X"52",X"90",X"90",X"90",X"90",X"90",X"54",X"57",X"55",X"90",X"56",X"90",
		X"90",X"90",X"90",X"90",X"90",X"01",X"02",X"03",X"03",X"04",X"03",X"02",X"01",X"01",X"02",X"01",
		X"02",X"03",X"04",X"05",X"04",X"03",X"02",X"02",X"03",X"02",X"01",X"01",X"02",X"03",X"04",X"03",
		X"02",X"01",X"01",X"02",X"01",X"00",X"00",X"04",X"80",X"00",X"16",X"00",X"00",X"00",X"00",X"00",
		X"76",X"1A",X"00",X"03",X"00",X"00",X"00",X"00",X"76",X"1A",X"00",X"03",X"23",X"05",X"54",X"09",
		X"42",X"13",X"00",X"18",X"00",X"24",X"03",X"02",X"02",X"1B",X"01",X"00",X"FF",X"B4",X"6E",X"02",
		X"02",X"1B",X"01",X"00",X"FF",X"AF",X"8C",X"02",X"02",X"1B",X"01",X"00",X"FF",X"AA",X"50",X"05",
		X"03",X"02",X"02",X"1B",X"01",X"00",X"01",X"A0",X"6E",X"02",X"02",X"1B",X"01",X"00",X"01",X"AF",
		X"8C",X"05",X"03",X"02",X"02",X"1B",X"01",X"00",X"01",X"B4",X"50",X"05",X"02",X"03",X"01",X"05",
		X"02",X"01",X"18",X"02",X"00",X"00",X"0C",X"6E",X"02",X"01",X"18",X"02",X"00",X"00",X"0C",X"B4",
		X"01",X"0A",X"02",X"01",X"18",X"01",X"00",X"00",X"14",X"80",X"02",X"01",X"18",X"01",X"00",X"00",
		X"10",X"50",X"05",X"03",X"02",X"01",X"18",X"01",X"00",X"00",X"14",X"80",X"02",X"01",X"18",X"01",
		X"00",X"00",X"12",X"C8",X"02",X"01",X"18",X"01",X"00",X"00",X"10",X"C8",X"02",X"01",X"18",X"01",
		X"00",X"00",X"0E",X"80",X"05",X"02",X"03",X"02",X"03",X"1D",X"01",X"00",X"01",X"0C",X"50",X"02",
		X"03",X"1D",X"01",X"00",X"01",X"12",X"5A",X"02",X"03",X"1D",X"01",X"00",X"01",X"0E",X"C8",X"02",
		X"03",X"1D",X"02",X"00",X"01",X"16",X"C8",X"05",X"03",X"02",X"03",X"1D",X"01",X"00",X"01",X"1E",
		X"64",X"02",X"03",X"1D",X"01",X"00",X"01",X"1A",X"64",X"05",X"02",X"03",X"02",X"04",X"1C",X"01",
		X"00",X"01",X"0C",X"32",X"02",X"04",X"1C",X"01",X"00",X"01",X"0C",X"C8",X"05",X"02",X"02",X"04",
		X"1C",X"01",X"00",X"FF",X"0C",X"80",X"02",X"04",X"1C",X"01",X"00",X"FF",X"0D",X"50",X"02",X"04",
		X"1C",X"01",X"00",X"FF",X"0D",X"C8",X"05",X"02",X"02",X"04",X"1C",X"02",X"00",X"FF",X"0D",X"32",
		X"05",X"02",X"02",X"04",X"1C",X"01",X"00",X"01",X"10",X"32",X"01",X"05",X"02",X"04",X"1C",X"01",
		X"00",X"FF",X"10",X"C8",X"05",X"03",X"02",X"04",X"1C",X"02",X"00",X"01",X"10",X"80",X"05",X"02",
		X"03",X"02",X"05",X"1E",X"01",X"00",X"FF",X"64",X"80",X"02",X"05",X"1E",X"01",X"00",X"FF",X"96",
		X"B4",X"02",X"05",X"1E",X"01",X"00",X"FF",X"5A",X"B4",X"02",X"05",X"1E",X"01",X"00",X"FF",X"10",
		X"80",X"05",X"03",X"02",X"05",X"1E",X"01",X"00",X"FF",X"20",X"80",X"02",X"05",X"1E",X"01",X"00",
		X"01",X"20",X"80",X"01",X"14",X"05",X"02",X"04",X"80",X"01",X"81",X"20",X"81",X"01",X"81",X"02",
		X"00",X"08",X"00",X"04",X"00",X"80",X"00",X"20",X"01",X"08",X"01",X"04",X"00",X"40",X"00",X"02",
		X"80",X"10",X"81",X"10",X"50",X"00",X"00",X"01",X"50",X"00",X"00",X"01",X"00",X"03",X"00",X"06",
		X"00",X"03",X"00",X"06",X"FE",X"0A",X"90",X"0A",X"7C",X"0A",X"58",X"0A",X"20",X"0A",X"58",X"0A",
		X"7C",X"0A",X"90",X"0A",X"7C",X"0A",X"58",X"14",X"20",X"14",X"FE",X"0A",X"90",X"0A",X"7C",X"0A",
		X"58",X"0A",X"20",X"0A",X"58",X"0A",X"7C",X"0A",X"90",X"0A",X"7C",X"0A",X"58",X"14",X"90",X"FF",
		X"FF",X"FF",X"FF",X"FE",X"10",X"80",X"10",X"58",X"10",X"38",X"10",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FE",X"0A",X"40",X"0A",X"20",X"0A",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FE",X"08",X"90",X"08",X"20",X"08",X"90",X"08",X"20",X"08",X"90",X"08",X"20",
		X"08",X"FF",X"FF",X"FE",X"08",X"9C",X"0A",X"90",X"0A",X"80",X"0A",X"7C",X"0A",X"80",X"0A",X"90",
		X"1E",X"20",X"1E",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C9",X"CD",X"4C",X"1B",X"5E",X"23",
		X"56",X"EB",X"C9",X"78",X"FE",X"05",X"D2",X"7D",X"1B",X"D5",X"CD",X"3E",X"1B",X"D1",X"B7",X"3E",
		X"2D",X"CA",X"79",X"18",X"7E",X"B7",X"F2",X"79",X"18",X"2F",X"C3",X"79",X"18",X"F5",X"7E",X"B7",
		X"FA",X"8B",X"1B",X"CD",X"79",X"18",X"3E",X"3D",X"C3",X"91",X"1B",X"2F",X"CD",X"79",X"18",X"3E",
		X"27",X"CD",X"79",X"18",X"F1",X"C2",X"A8",X"1B",X"7E",X"B7",X"21",X"C1",X"21",X"FA",X"A3",X"1B",
		X"21",X"F1",X"21",X"7E",X"CD",X"C1",X"18",X"C9",X"D5",X"CD",X"5B",X"1B",X"CD",X"23",X"19",X"D1",
		X"C9",X"CD",X"D1",X"18",X"CD",X"77",X"18",X"06",X"00",X"C5",X"E5",X"CD",X"63",X"1B",X"E1",X"C1",
		X"04",X"23",X"78",X"FE",X"0B",X"D0",X"FE",X"05",X"DA",X"B9",X"1B",X"CD",X"77",X"18",X"C3",X"B9",
		X"1B",X"11",X"35",X"1D",X"21",X"2A",X"1D",X"CD",X"B1",X"1B",X"11",X"45",X"1D",X"21",X"3A",X"1D",
		X"CD",X"B1",X"1B",X"CD",X"77",X"18",X"CD",X"20",X"1F",X"F5",X"D5",X"C5",X"CD",X"D6",X"13",X"D2",
		X"19",X"1C",X"2A",X"F6",X"21",X"22",X"0C",X"00",X"21",X"10",X"00",X"36",X"FF",X"CD",X"06",X"00",
		X"C3",X"63",X"1C",X"0E",X"00",X"FE",X"CB",X"CA",X"12",X"1C",X"FE",X"DD",X"D8",X"E6",X"CF",X"FE",
		X"CD",X"C0",X"23",X"7E",X"4F",X"CD",X"C1",X"18",X"C9",X"2B",X"22",X"66",X"21",X"2A",X"F6",X"21",
		X"7E",X"CD",X"C1",X"18",X"7E",X"CD",X"03",X"1C",X"23",X"CD",X"3A",X"19",X"DA",X"63",X"1C",X"F5",
		X"CD",X"77",X"18",X"F1",X"B3",X"CA",X"4A",X"1C",X"5E",X"23",X"56",X"79",X"FE",X"36",X"C2",X"44",
		X"1C",X"7A",X"53",X"5F",X"CD",X"EA",X"18",X"C3",X"63",X"1C",X"7E",X"CD",X"C1",X"18",X"2A",X"F6",
		X"21",X"7E",X"E6",X"C7",X"FE",X"00",X"C2",X"63",X"1C",X"23",X"5E",X"16",X"00",X"2B",X"19",X"EB",
		X"CD",X"EA",X"18",X"2A",X"F6",X"21",X"7E",X"47",X"E6",X"C0",X"FE",X"80",X"C2",X"7A",X"1C",X"78",
		X"E6",X"07",X"FE",X"06",X"C2",X"26",X"1D",X"C3",X"A7",X"1C",X"FE",X"40",X"C2",X"97",X"1C",X"78",
		X"FE",X"76",X"CA",X"26",X"1D",X"E6",X"07",X"FE",X"06",X"CA",X"B3",X"1C",X"78",X"E6",X"38",X"FE",
		X"30",X"C2",X"26",X"1D",X"C3",X"B3",X"1C",X"78",X"FE",X"36",X"CA",X"B3",X"1C",X"FE",X"34",X"CA",
		X"A7",X"1C",X"FE",X"35",X"C2",X"B9",X"1C",X"3E",X"3D",X"CD",X"79",X"18",X"2A",X"F4",X"21",X"7E",
		X"CD",X"C1",X"18",X"2A",X"F4",X"21",X"C3",X"CC",X"1C",X"E6",X"E7",X"FE",X"02",X"C2",X"E0",X"1C",
		X"78",X"E6",X"10",X"2A",X"EC",X"21",X"C2",X"CC",X"1C",X"2A",X"EE",X"21",X"3A",X"4A",X"21",X"B7",
		X"C2",X"26",X"1D",X"EB",X"CD",X"F3",X"20",X"CA",X"26",X"1D",X"CD",X"F9",X"18",X"C3",X"26",X"1D",
		X"78",X"FE",X"CB",X"C2",X"F4",X"1C",X"2A",X"AE",X"21",X"7E",X"E6",X"07",X"FE",X"06",X"C2",X"26",
		X"1D",X"C3",X"B3",X"1C",X"E6",X"DD",X"FE",X"DD",X"C2",X"26",X"1D",X"2A",X"AE",X"21",X"7E",X"FE",
		X"39",X"CA",X"26",X"1D",X"FE",X"34",X"DA",X"26",X"1D",X"FE",X"CC",X"CA",X"26",X"1D",X"23",X"5E",
		X"16",X"00",X"78",X"FE",X"DD",X"CA",X"1F",X"1D",X"FD",X"E5",X"E1",X"19",X"C3",X"CC",X"1C",X"DD",
		X"E5",X"E1",X"19",X"C3",X"CC",X"1C",X"C1",X"D1",X"F1",X"C9",X"43",X"5A",X"4D",X"45",X"49",X"41",
		X"42",X"44",X"48",X"53",X"50",X"F6",X"F4",X"FC",X"FA",X"FE",X"BC",X"A5",X"B2",X"BA",X"B6",X"BE",
		X"BD",X"BB",X"B7",X"58",X"59",X"C6",X"C4",X"C2",X"C0",X"BE",X"01",X"07",X"08",X"03",X"05",X"21",
		X"00",X"00",X"22",X"54",X"21",X"AF",X"32",X"53",X"21",X"C9",X"F3",X"22",X"F4",X"21",X"E1",X"2B",
		X"22",X"F6",X"21",X"F5",X"21",X"02",X"00",X"39",X"F1",X"31",X"F4",X"21",X"E5",X"F5",X"C5",X"D5",
		X"21",X"00",X"00",X"39",X"31",X"C2",X"21",X"08",X"F5",X"08",X"D9",X"C5",X"D5",X"E5",X"D9",X"DD",
		X"E5",X"FD",X"E5",X"F9",X"00",X"00",X"00",X"FB",X"2A",X"F6",X"21",X"7E",X"FE",X"FF",X"F5",X"E5",
		X"3A",X"20",X"21",X"32",X"44",X"21",X"21",X"40",X"21",X"0E",X"08",X"E5",X"7E",X"B7",X"CA",X"A8",
		X"1D",X"23",X"5E",X"23",X"56",X"23",X"7E",X"12",X"E1",X"11",X"FC",X"FF",X"19",X"0D",X"C2",X"9B",
		X"1D",X"CD",X"FD",X"1E",X"21",X"56",X"21",X"7E",X"36",X"00",X"B7",X"CA",X"CB",X"1D",X"3D",X"47",
		X"23",X"5E",X"23",X"56",X"23",X"7E",X"12",X"78",X"C3",X"BA",X"1D",X"E1",X"F1",X"CA",X"EF",X"1D",
		X"23",X"22",X"F6",X"21",X"EB",X"21",X"B5",X"0E",X"4E",X"23",X"46",X"CD",X"17",X"11",X"DA",X"EF",
		X"1D",X"CD",X"4F",X"1D",X"2A",X"51",X"21",X"EB",X"3E",X"82",X"B7",X"37",X"C3",X"55",X"11",X"3A",
		X"23",X"21",X"B7",X"C2",X"94",X"1E",X"21",X"24",X"21",X"0E",X"08",X"E5",X"7E",X"B7",X"CA",X"51",
		X"1E",X"23",X"7E",X"23",X"56",X"2A",X"F6",X"21",X"BD",X"C2",X"51",X"1E",X"7A",X"BC",X"C2",X"51",
		X"1E",X"E1",X"7E",X"3D",X"C2",X"1F",X"1E",X"F5",X"3D",X"32",X"23",X"21",X"C3",X"36",X"1E",X"77",
		X"F5",X"CD",X"CA",X"1E",X"FE",X"02",X"CA",X"36",X"1E",X"3A",X"4A",X"21",X"B7",X"CA",X"36",X"1E",
		X"CD",X"20",X"1F",X"C3",X"55",X"11",X"CD",X"D1",X"18",X"F1",X"3C",X"CD",X"C1",X"18",X"21",X"C3",
		X"1E",X"CD",X"86",X"18",X"2A",X"F6",X"21",X"EB",X"CD",X"EA",X"18",X"CD",X"D1",X"1B",X"C3",X"55",
		X"11",X"E1",X"11",X"04",X"00",X"19",X"0D",X"C2",X"FB",X"1D",X"CD",X"DB",X"18",X"C2",X"94",X"1E",
		X"CD",X"CA",X"1E",X"CA",X"7C",X"1E",X"3D",X"C2",X"70",X"1E",X"CD",X"20",X"1F",X"C3",X"55",X"11",
		X"2A",X"F6",X"21",X"CD",X"0C",X"19",X"CD",X"D1",X"1B",X"C3",X"55",X"11",X"3A",X"44",X"21",X"B7",
		X"CA",X"94",X"1E",X"2A",X"48",X"21",X"4D",X"44",X"2A",X"46",X"21",X"EB",X"3A",X"45",X"21",X"B7",
		X"37",X"C3",X"55",X"11",X"CD",X"D1",X"18",X"CD",X"FD",X"1E",X"21",X"00",X"00",X"22",X"4F",X"21",
		X"CD",X"4F",X"1D",X"32",X"23",X"21",X"3E",X"2A",X"CD",X"79",X"18",X"2A",X"F6",X"21",X"CD",X"D6",
		X"13",X"D2",X"B7",X"1E",X"22",X"0C",X"00",X"CD",X"E9",X"18",X"2A",X"F4",X"21",X"22",X"64",X"21",
		X"C3",X"16",X"0F",X"20",X"50",X"41",X"53",X"53",X"20",X"00",X"21",X"53",X"21",X"7E",X"B7",X"C8",
		X"E5",X"2A",X"54",X"21",X"2B",X"22",X"54",X"21",X"7C",X"B5",X"E1",X"C2",X"E3",X"1E",X"77",X"3D",
		X"32",X"23",X"21",X"7E",X"B7",X"C9",X"11",X"13",X"00",X"21",X"CD",X"20",X"7E",X"A0",X"23",X"BE",
		X"23",X"CA",X"F9",X"1E",X"14",X"1D",X"C2",X"EC",X"1E",X"5A",X"16",X"00",X"C9",X"3A",X"20",X"21",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",
		X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F0",X"B0",X"B0",X"B0",X"F8",X"B8",X"B8",X"B8",X"F8");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
