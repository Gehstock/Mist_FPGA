library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_C1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_C1 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"0F",X"EC",X"28",X"F2",X"FE",X"1F",X"08",X"72",X"2A",X"F2",X"FE",X"1F",X"08",X"80",X"2B",X"F2",
		X"FE",X"1F",X"08",X"8E",X"2C",X"F2",X"FE",X"1F",X"08",X"9C",X"2D",X"F2",X"FE",X"1F",X"08",X"AA",
		X"2E",X"F2",X"FE",X"1F",X"08",X"B8",X"2F",X"F2",X"FE",X"1F",X"08",X"C6",X"30",X"F2",X"FE",X"1F",
		X"08",X"D4",X"31",X"F2",X"FE",X"1F",X"08",X"E2",X"32",X"F2",X"FE",X"1F",X"08",X"FA",X"29",X"88",
		X"FF",X"5F",X"0A",X"84",X"74",X"64",X"64",X"34",X"24",X"14",X"04",X"3C",X"2C",X"1C",X"0C",X"6C",
		X"7C",X"8C",X"9C",X"70",X"71",X"72",X"73",X"33",X"34",X"35",X"36",X"57",X"58",X"59",X"5A",X"3C",
		X"3D",X"3E",X"3F",X"71",X"72",X"73",X"74",X"3B",X"4B",X"5B",X"6B",X"25",X"15",X"05",X"05",X"8C",
		X"8D",X"8E",X"8F",X"70",X"71",X"72",X"73",X"0A",X"1A",X"2A",X"3A",X"37",X"47",X"57",X"67",X"8C",
		X"8D",X"8E",X"8F",X"70",X"71",X"72",X"73",X"34",X"35",X"36",X"37",X"48",X"49",X"4A",X"4B",X"7C",
		X"7D",X"7E",X"7F",X"53",X"54",X"55",X"56",X"46",X"47",X"48",X"49",X"39",X"3A",X"3B",X"3C",X"7C",
		X"7D",X"7E",X"7F",X"80",X"81",X"82",X"83",X"36",X"46",X"56",X"66",X"39",X"3A",X"3B",X"3C",X"7C",
		X"7D",X"7E",X"7F",X"70",X"71",X"72",X"73",X"28",X"38",X"48",X"58",X"0B",X"1B",X"2B",X"3B",X"6C",
		X"6D",X"6E",X"6F",X"60",X"61",X"62",X"63",X"98",X"88",X"78",X"68",X"49",X"4A",X"4B",X"4C",X"6C",
		X"6D",X"6E",X"6F",X"90",X"91",X"92",X"93",X"04",X"14",X"24",X"34",X"49",X"4A",X"4B",X"4C",X"7C",
		X"7D",X"7E",X"7F",X"96",X"A6",X"B6",X"C6",X"D6",X"00",X"00",X"00",X"00",X"3F",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"95",X"FB",X"33",X"33",X"33",X"33",
		X"22",X"22",X"22",X"22",X"22",X"22",X"33",X"34",X"44",X"D9",X"A2",X"33",X"33",X"32",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"23",X"34",X"44",X"5E",X"A2",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"33",X"44",X"5E",X"A2",X"22",X"21",X"12",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"33",X"55",X"5E",X"A2",X"11",X"1F",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"44",X"55",X"5E",X"A1",X"10",X"16",X"65",X"55",X"55",X"55",X"D9",X"11",X"1F",
		X"B4",X"55",X"55",X"55",X"5E",X"A1",X"00",X"07",X"66",X"66",X"55",X"56",X"6D",X"91",X"FB",X"44",
		X"55",X"55",X"55",X"6E",X"A1",X"00",X"07",X"77",X"66",X"66",X"66",X"66",X"EF",X"B4",X"44",X"55",
		X"66",X"66",X"6E",X"D9",X"10",X"07",X"77",X"76",X"66",X"66",X"66",X"EB",X"34",X"45",X"56",X"66",
		X"66",X"6E",X"1D",X"90",X"07",X"77",X"77",X"77",X"77",X"7F",X"B3",X"34",X"45",X"67",X"77",X"77",
		X"6E",X"3F",X"CC",X"CC",X"CC",X"10",X"77",X"77",X"FB",X"33",X"33",X"44",X"88",X"88",X"88",X"8B",
		X"FB",X"22",X"22",X"22",X"10",X"00",X"7F",X"B2",X"22",X"22",X"22",X"33",X"34",X"44",X"D9",X"A2",
		X"22",X"22",X"22",X"11",X"10",X"FA",X"22",X"22",X"22",X"22",X"23",X"33",X"44",X"5E",X"A2",X"22",
		X"22",X"21",X"11",X"0F",X"BA",X"22",X"22",X"22",X"22",X"22",X"33",X"44",X"5E",X"A2",X"21",X"11",
		X"11",X"00",X"FB",X"5D",X"92",X"22",X"22",X"22",X"22",X"23",X"44",X"5E",X"A1",X"10",X"00",X"10",
		X"0F",X"B5",X"55",X"D9",X"11",X"11",X"11",X"11",X"24",X"44",X"5E",X"A1",X"11",X"10",X"DC",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"B5",X"54",X"4E",X"A1",X"00",X"07",X"65",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"4E",X"A1",X"00",X"07",X"65",X"56",X"65",X"66",
		X"66",X"66",X"66",X"66",X"66",X"65",X"55",X"5E",X"A1",X"00",X"76",X"66",X"66",X"66",X"66",X"66",
		X"66",X"66",X"66",X"66",X"66",X"55",X"5E",X"A1",X"00",X"77",X"66",X"66",X"66",X"66",X"66",X"66",
		X"66",X"66",X"66",X"66",X"65",X"5E",X"A1",X"00",X"77",X"76",X"66",X"66",X"66",X"66",X"66",X"66",
		X"66",X"66",X"66",X"65",X"5E",X"A1",X"00",X"77",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"66",X"66",X"66",X"6E",X"D9",X"00",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"77",X"77",X"FB",X"1D",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"B7",X"3F",X"CC",X"CC",X"CC",X"CC",X"95",X"3F",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"95",X"FB",X"33",X"34",X"44",X"45",X"D9",X"FB",X"22",X"22",X"22",X"23",X"33",X"34",X"45",X"D9",
		X"A2",X"23",X"33",X"44",X"44",X"5E",X"B2",X"22",X"22",X"22",X"22",X"33",X"34",X"45",X"5E",X"A2",
		X"22",X"33",X"44",X"44",X"5E",X"22",X"22",X"22",X"22",X"22",X"23",X"34",X"55",X"5E",X"A2",X"22",
		X"23",X"34",X"44",X"5E",X"22",X"22",X"22",X"12",X"22",X"12",X"34",X"55",X"5E",X"A2",X"11",X"12",
		X"34",X"44",X"4E",X"11",X"11",X"11",X"F8",X"88",X"88",X"45",X"55",X"5E",X"A1",X"11",X"0E",X"34",
		X"44",X"5E",X"11",X"11",X"17",X"A1",X"FB",X"44",X"55",X"55",X"5E",X"A1",X"11",X"7E",X"34",X"44",
		X"5E",X"11",X"11",X"07",X"D8",X"B4",X"44",X"55",X"55",X"6E",X"A1",X"10",X"7E",X"34",X"44",X"5E",
		X"11",X"10",X"07",X"7A",X"34",X"44",X"55",X"56",X"6E",X"A1",X"00",X"0E",X"33",X"44",X"5E",X"91",
		X"00",X"00",X"7A",X"33",X"44",X"55",X"66",X"FB",X"A0",X"00",X"0E",X"33",X"33",X"4E",X"D9",X"00",
		X"77",X"7A",X"33",X"34",X"56",X"6F",X"B7",X"A0",X"00",X"0E",X"33",X"33",X"3D",X"8B",X"10",X"77",
		X"7A",X"33",X"34",X"4C",X"CC",X"95",X"A0",X"00",X"0E",X"33",X"33",X"33",X"21",X"00",X"07",X"7A",
		X"23",X"33",X"34",X"44",X"D9",X"A1",X"00",X"7E",X"22",X"22",X"22",X"21",X"00",X"00",X"7A",X"22",
		X"33",X"34",X"44",X"5E",X"A1",X"00",X"7E",X"22",X"22",X"22",X"11",X"00",X"00",X"7A",X"22",X"23",
		X"34",X"44",X"4E",X"A1",X"00",X"7D",X"91",X"22",X"21",X"11",X"00",X"00",X"FC",X"92",X"22",X"34",
		X"44",X"4E",X"A1",X"00",X"07",X"D9",X"11",X"11",X"11",X"00",X"0F",X"B5",X"D9",X"22",X"34",X"44",
		X"4E",X"A1",X"00",X"07",X"7D",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"44",X"44",X"4E",
		X"3F",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"95",X"FB",
		X"44",X"45",X"55",X"56",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"D9",X"A4",X"44",
		X"45",X"55",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"6E",X"A3",X"44",X"45",
		X"55",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"6E",X"A3",X"44",X"44",X"5F",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"97",X"77",X"7E",X"A3",X"33",X"44",X"4D",X"9F",
		X"B3",X"33",X"33",X"33",X"33",X"3D",X"9F",X"B0",X"07",X"7E",X"D9",X"33",X"34",X"44",X"DB",X"22",
		X"22",X"22",X"33",X"33",X"33",X"DB",X"10",X"07",X"7E",X"0D",X"93",X"33",X"44",X"42",X"22",X"22",
		X"22",X"22",X"33",X"32",X"21",X"10",X"00",X"7E",X"01",X"D9",X"33",X"34",X"12",X"22",X"22",X"22",
		X"22",X"22",X"22",X"11",X"10",X"00",X"0E",X"00",X"1D",X"93",X"33",X"11",X"11",X"1F",X"88",X"89",
		X"22",X"21",X"11",X"10",X"00",X"7E",X"00",X"01",X"E1",X"13",X"11",X"11",X"4A",X"11",X"1D",X"92",
		X"11",X"11",X"10",X"07",X"FB",X"00",X"0F",X"B1",X"13",X"33",X"33",X"3D",X"93",X"33",X"D8",X"88",
		X"88",X"88",X"88",X"B7",X"00",X"FB",X"11",X"10",X"33",X"33",X"33",X"DC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"95",X"0F",X"B1",X"11",X"07",X"22",X"23",X"22",X"22",X"22",X"22",X"22",X"33",X"34",
		X"44",X"D9",X"FB",X"11",X"10",X"07",X"F9",X"22",X"22",X"22",X"22",X"22",X"22",X"23",X"34",X"44",
		X"5E",X"A1",X"11",X"00",X"0F",X"BD",X"92",X"22",X"22",X"22",X"22",X"22",X"22",X"34",X"44",X"5E",
		X"A1",X"10",X"00",X"FB",X"55",X"D9",X"11",X"11",X"11",X"11",X"11",X"22",X"24",X"44",X"5E",X"A1",
		X"00",X"00",X"6C",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"B4",X"44",X"4E",X"3F",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"9F",X"CC",X"CC",X"CC",X"95",X"FB",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"33",X"34",X"DB",X"23",X"33",X"34",X"D9",X"A2",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"23",X"33",X"32",X"22",X"33",X"34",X"4E",X"A2",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"23",X"22",X"22",X"23",X"34",X"5E",X"A2",X"22",X"12",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"11",X"12",X"45",X"5E",X"A1",X"11",X"11",X"FC",X"CC",X"CC",X"CC",
		X"CC",X"C9",X"33",X"33",X"33",X"F4",X"55",X"5E",X"A1",X"11",X"1F",X"B4",X"44",X"45",X"55",X"56",
		X"6D",X"88",X"88",X"88",X"B5",X"55",X"5E",X"A1",X"11",X"0E",X"34",X"44",X"45",X"55",X"56",X"66",
		X"66",X"66",X"66",X"56",X"66",X"6E",X"A1",X"10",X"0E",X"34",X"44",X"45",X"56",X"66",X"66",X"66",
		X"66",X"66",X"66",X"66",X"6E",X"A1",X"00",X"0E",X"33",X"44",X"45",X"66",X"66",X"66",X"66",X"66",
		X"66",X"66",X"66",X"6E",X"A0",X"00",X"0E",X"33",X"34",X"45",X"89",X"77",X"77",X"66",X"66",X"66",
		X"66",X"66",X"FB",X"A0",X"00",X"0E",X"33",X"33",X"4E",X"4D",X"97",X"77",X"77",X"77",X"77",X"77",
		X"7F",X"B7",X"A0",X"00",X"0E",X"22",X"23",X"33",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"95",X"A0",X"00",X"0E",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"23",X"33",X"44",X"44",X"D9",
		X"A0",X"00",X"0E",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"33",X"34",X"44",X"5E",X"A0",
		X"00",X"0D",X"92",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"23",X"34",X"45",X"5E",X"A0",X"00",
		X"76",X"D9",X"11",X"11",X"11",X"11",X"11",X"11",X"22",X"22",X"34",X"55",X"5E",X"A0",X"00",X"07",
		X"6D",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"45",X"55",X"5E",X"3F",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"95",X"43",X"FC",X"CC",X"CC",X"CC",X"CC",X"CC",X"95",X"FB",X"22",X"23",X"33",X"34",
		X"45",X"D9",X"3F",X"B2",X"23",X"33",X"33",X"44",X"44",X"D9",X"A2",X"22",X"22",X"33",X"34",X"44",
		X"5D",X"8B",X"22",X"22",X"33",X"33",X"44",X"44",X"5E",X"A2",X"22",X"22",X"23",X"34",X"44",X"55",
		X"E2",X"22",X"22",X"23",X"33",X"44",X"44",X"5E",X"A1",X"11",X"11",X"12",X"34",X"44",X"55",X"E2",
		X"22",X"22",X"22",X"33",X"44",X"44",X"5E",X"A1",X"11",X"11",X"FC",X"94",X"44",X"45",X"E1",X"11",
		X"11",X"1F",X"93",X"44",X"44",X"5E",X"A1",X"11",X"17",X"D9",X"A4",X"44",X"45",X"E1",X"11",X"11",
		X"1A",X"D9",X"34",X"44",X"5E",X"A1",X"11",X"07",X"7D",X"A3",X"44",X"45",X"E1",X"11",X"10",X"7D",
		X"9A",X"44",X"44",X"5E",X"D9",X"00",X"07",X"76",X"A3",X"34",X"45",X"E9",X"11",X"00",X"77",X"DA",
		X"44",X"44",X"5E",X"2A",X"00",X"00",X"76",X"A3",X"33",X"45",X"AD",X"90",X"00",X"07",X"6A",X"44",
		X"44",X"5E",X"FB",X"10",X"00",X"7E",X"23",X"33",X"35",X"A4",X"E0",X"00",X"07",X"7A",X"44",X"44",
		X"5E",X"A1",X"10",X"00",X"7E",X"23",X"33",X"33",X"D8",X"B1",X"10",X"07",X"7A",X"44",X"44",X"5E",
		X"A1",X"10",X"00",X"7A",X"23",X"33",X"33",X"32",X"11",X"00",X"07",X"7A",X"44",X"44",X"5E",X"A1",
		X"10",X"00",X"7A",X"22",X"22",X"22",X"22",X"11",X"00",X"07",X"7A",X"44",X"45",X"5E",X"A1",X"00",
		X"00",X"7A",X"22",X"22",X"22",X"21",X"11",X"00",X"07",X"7A",X"44",X"55",X"5E",X"A1",X"00",X"00",
		X"7D",X"92",X"22",X"22",X"11",X"10",X"00",X"07",X"FB",X"45",X"55",X"5E",X"A1",X"00",X"00",X"76",
		X"D9",X"11",X"11",X"11",X"10",X"00",X"0F",X"B4",X"55",X"55",X"5E",X"A1",X"00",X"00",X"77",X"6D",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CB",X"55",X"55",X"55",X"5E",X"23",X"FC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"95",X"44",X"3F",X"CC",X"CC",X"CC",X"CC",X"95",X"3F",X"B2",X"22",X"23",X"33",X"44",X"44",
		X"D9",X"53",X"FB",X"33",X"33",X"34",X"45",X"D9",X"2A",X"22",X"22",X"22",X"33",X"34",X"44",X"4D",
		X"9F",X"B3",X"23",X"33",X"34",X"44",X"5E",X"2A",X"22",X"22",X"22",X"23",X"33",X"34",X"44",X"DA",
		X"22",X"22",X"33",X"34",X"44",X"5E",X"2A",X"22",X"11",X"11",X"22",X"33",X"34",X"44",X"4A",X"22",
		X"22",X"23",X"34",X"44",X"5E",X"2A",X"11",X"11",X"10",X"EA",X"23",X"34",X"44",X"4A",X"22",X"22",
		X"22",X"34",X"44",X"5E",X"2A",X"11",X"11",X"07",X"7D",X"92",X"34",X"44",X"4A",X"11",X"11",X"1E",
		X"44",X"44",X"4E",X"1D",X"91",X"10",X"07",X"77",X"D9",X"33",X"44",X"4A",X"11",X"11",X"0E",X"44",
		X"44",X"4E",X"11",X"D9",X"00",X"07",X"77",X"7E",X"33",X"44",X"4A",X"11",X"10",X"0E",X"44",X"44",
		X"4E",X"11",X"1D",X"90",X"07",X"77",X"7E",X"33",X"34",X"4A",X"11",X"00",X"0E",X"44",X"44",X"4E",
		X"13",X"41",X"D9",X"07",X"77",X"7E",X"33",X"34",X"4A",X"10",X"00",X"0E",X"44",X"44",X"4E",X"3F",
		X"CC",X"CB",X"10",X"77",X"7E",X"33",X"33",X"4B",X"10",X"00",X"0E",X"44",X"44",X"4E",X"FB",X"22",
		X"22",X"10",X"01",X"1E",X"22",X"22",X"32",X"10",X"00",X"0E",X"44",X"44",X"4E",X"A2",X"22",X"21",
		X"10",X"00",X"7E",X"22",X"22",X"21",X"10",X"00",X"0E",X"44",X"44",X"4E",X"A2",X"21",X"11",X"00",
		X"00",X"0E",X"22",X"22",X"11",X"00",X"00",X"0E",X"44",X"54",X"4E",X"A2",X"11",X"11",X"00",X"00",
		X"FC",X"92",X"21",X"11",X"00",X"00",X"FB",X"55",X"44",X"4E",X"A1",X"11",X"11",X"00",X"0F",X"B1",
		X"D9",X"11",X"11",X"00",X"0F",X"B5",X"55",X"44",X"4E",X"A0",X"00",X"0D",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"CB",X"55",X"55",X"44",X"4E",X"3F",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"93",X"FC",X"CC",X"CC",X"CC",X"CC",X"95",X"FB",X"22",X"22",X"22",X"23",X"33",X"34",X"44",X"D8",
		X"B2",X"23",X"33",X"34",X"44",X"D9",X"A2",X"22",X"22",X"22",X"22",X"33",X"34",X"44",X"5E",X"22",
		X"22",X"33",X"34",X"44",X"4E",X"A2",X"22",X"22",X"22",X"22",X"23",X"34",X"45",X"5E",X"22",X"22",
		X"23",X"34",X"44",X"4E",X"A2",X"22",X"11",X"11",X"11",X"22",X"34",X"55",X"5E",X"22",X"22",X"22");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
