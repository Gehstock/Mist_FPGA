library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity obj_7t is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of obj_7t is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"07",X"00",X"00",X"00",X"00",X"0C",X"1E",X"1C",X"1F",X"0F",X"06",X"00",X"00",X"00",X"00",
		X"0C",X"18",X"1C",X"18",X"00",X"00",X"00",X"04",X"0E",X"3E",X"7C",X"3D",X"00",X"00",X"00",X"00",
		X"30",X"60",X"60",X"60",X"00",X"00",X"01",X"03",X"17",X"37",X"37",X"0A",X"00",X"00",X"00",X"00",
		X"78",X"38",X"00",X"00",X"00",X"00",X"00",X"24",X"7E",X"7E",X"3C",X"0D",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"1C",X"08",X"08",X"00",X"00",X"0D",X"1F",X"07",X"07",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"30",X"18",X"08",X"03",X"07",X"07",X"07",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"3C",X"00",X"00",X"00",X"1E",X"3E",X"78",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"40",X"70",X"38",X"10",X"04",X"0E",X"3E",X"7C",X"39",X"00",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0E",
		X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"EE",X"FE",X"FE",X"7D",X"33",X"00",X"03",X"02",X"00",
		X"00",X"02",X"08",X"00",X"00",X"00",X"04",X"EE",X"FE",X"FE",X"7D",X"33",X"00",X"03",X"02",X"00",
		X"10",X"80",X"20",X"00",X"00",X"00",X"04",X"EE",X"EE",X"FE",X"7D",X"33",X"00",X"03",X"02",X"00",
		X"78",X"00",X"00",X"00",X"00",X"18",X"1D",X"FE",X"7D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"78",X"00",X"00",X"00",X"3D",X"FC",X"39",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"20",X"20",X"C2",X"01",X"02",X"09",X"09",X"18",X"18",X"38",X"10",X"03",X"03",X"00",
		X"10",X"10",X"20",X"20",X"C2",X"01",X"02",X"29",X"79",X"78",X"38",X"18",X"00",X"03",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"06",X"47",X"E0",X"C0",X"C0",X"40",X"04",X"0E",X"0E",X"3E",X"3E",X"3E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"1F",X"3E",X"1C",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"0E",X"0F",X"0F",X"07",X"06",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"3F",X"7F",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"7F",X"3F",
		X"00",X"00",X"18",X"38",X"3C",X"7F",X"7F",X"7F",X"7F",X"3F",X"3F",X"1F",X"1F",X"0F",X"07",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"38",X"3E",X"7F",X"7F",X"7F",X"7F",X"3F",X"3F",X"1F",X"1F",X"0F",X"07",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",X"00",X"00",X"00",
		X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",X"FE",X"7E",X"7E",X"3E",X"1E",X"06",X"00",X"00",X"00",X"00",
		X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",X"FE",X"7E",X"7E",X"3E",X"1E",X"06",X"00",X"00",X"00",X"00",
		X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",X"FE",X"7E",X"7E",X"3E",X"1E",X"06",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"FC",X"FC",X"FC",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FC",X"FC",X"FC",
		X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",X"FE",X"7E",X"3E",X"7E",X"FE",X"FE",X"FC",X"FC",X"FC",X"FC",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",X"FE",X"7E",X"7E",X"3E",X"1E",X"06",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"00",X"00",X"00",X"00",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"00",X"00",X"00",X"00",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"7C",X"3E",X"0E",X"00",X"00",X"00",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FF",X"FF",X"FC",X"FC",X"FC",X"7C",X"3E",X"0E",X"00",X"00",X"00",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"7E",X"FE",X"FC",X"FC",X"FC",X"7C",X"3E",X"0E",X"00",X"00",X"00",
		X"1E",X"7E",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"7C",X"3E",X"0E",X"00",X"00",X"00",
		X"1E",X"7E",X"FC",X"FC",X"FC",X"7E",X"FE",X"FC",X"FC",X"FC",X"7C",X"3E",X"0E",X"00",X"00",X"00",
		X"3E",X"7E",X"FC",X"FC",X"7C",X"3E",X"0E",X"00",X"00",X"FC",X"7C",X"3E",X"0E",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"0E",X"0E",X"0E",X"FE",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"0E",X"0E",X"0E",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"00",X"00",X"00",X"00",X"06",X"1E",X"3E",X"7E",X"7E",X"FE",X"FE",X"FE",X"FC",X"FC",X"FC",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"07",X"1F",X"1F",X"3B",X"3F",X"3F",X"1F",X"1C",X"3F",X"38",X"73",X"F3",X"DB",X"49",X"07",
		X"03",X"07",X"1F",X"1F",X"3B",X"BF",X"FF",X"EF",X"7C",X"7F",X"38",X"13",X"03",X"1B",X"09",X"07",
		X"07",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"1F",X"3F",X"3F",X"3F",X"1F",X"1F",X"4F",X"FF",X"FF",X"FF",X"03",X"03",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"FF",X"FF",X"00",X"FF",X"FF",X"00",X"FF",X"FF",X"00",
		X"0D",X"0D",X"1D",X"39",X"FB",X"E3",X"0F",X"FE",X"F8",X"03",X"FF",X"FE",X"00",X"FF",X"FF",X"00",
		X"0D",X"0D",X"0D",X"0D",X"0D",X"0D",X"0D",X"0D",X"0D",X"0D",X"0D",X"0D",X"0D",X"0D",X"0D",X"0D",
		X"00",X"09",X"06",X"09",X"10",X"29",X"06",X"29",X"70",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"06",X"09",X"10",X"29",X"06",X"29",X"30",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"3F",X"61",X"D2",X"0C",X"52",X"21",X"12",X"0C",X"12",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"1C",X"3F",X"61",X"D2",X"0C",X"52",X"21",X"12",X"0C",X"12",X"00",X"00",X"00",X"00",X"00",
		X"18",X"3F",X"61",X"D2",X"0C",X"52",X"21",X"12",X"0C",X"12",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E1",X"C1",X"3F",X"61",X"D2",X"0C",X"52",X"21",X"12",X"0C",X"12",X"00",X"00",X"00",X"00",X"00",
		X"C1",X"BF",X"61",X"D2",X"0C",X"52",X"21",X"12",X"0C",X"12",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"1C",X"1E",X"1F",X"0C",X"08",X"01",X"02",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"11",X"1C",X"1F",X"0C",X"08",X"01",X"02",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0E",X"0F",X"0E",X"04",X"00",X"01",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"3F",X"0F",X"0F",X"04",X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"07",X"07",X"0F",X"09",X"02",X"02",X"04",X"00",X"00",X"00",X"01",X"01",X"00",
		X"00",X"01",X"0A",X"04",X"04",X"04",X"0A",X"01",X"00",X"01",X"F0",X"F8",X"F8",X"00",X"08",X"00",
		X"00",X"01",X"0A",X"04",X"04",X"04",X"0A",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"06",X"09",X"10",X"29",X"06",X"09",X"70",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"06",X"09",X"10",X"29",X"06",X"09",X"70",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"06",X"09",X"10",X"29",X"06",X"09",X"70",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"08",X"09",X"0A",X"0D",X"08",X"0D",X"06",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"00",X"01",X"02",X"02",X"09",X"0E",X"06",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"05",X"02",X"02",X"01",X"06",X"06",X"03",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"0A",X"04",X"04",X"04",X"0A",X"01",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"01",X"0A",X"04",X"04",X"04",X"0A",X"01",X"00",X"01",X"00",X"00",
		X"00",X"00",X"00",X"01",X"0A",X"04",X"04",X"04",X"0A",X"01",X"00",X"01",X"00",X"00",X"00",X"00",
		X"00",X"1F",X"10",X"0A",X"04",X"02",X"01",X"01",X"02",X"04",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"20",X"11",X"0A",X"04",X"02",X"03",X"01",X"02",X"04",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"41",X"23",X"16",X"0C",X"0E",X"13",X"03",X"0F",X"16",X"05",X"01",X"02",X"00",X"00",X"00",
		X"00",X"08",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"21",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"08",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"3F",X"0F",X"33",X"1C",X"0E",X"08",X"00",X"00",X"C0",X"F0",X"FC",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"BF",X"DF",X"07",X"00",X"03",X"01",X"00",X"80",X"C0",X"E0",X"F8",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"3E",X"1C",X"08",X"10",X"20",X"40",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"1F",X"0F",X"80",X"60",X"18",X"07",X"00",X"80",X"E0",X"F8",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"1F",X"07",X"80",X"60",X"18",X"07",X"00",X"80",X"E0",X"F8",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C0",X"80",X"00",X"7F",X"00",X"00",X"80",X"C0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"1F",X"11",X"11",X"01",X"00",X"10",X"11",X"F1",X"F1",
		X"FF",X"FF",X"FF",X"1F",X"11",X"11",X"01",X"01",X"10",X"10",X"11",X"F1",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F1",X"F1",X"10",X"10",X"01",X"01",X"11",X"11",X"1F",X"1F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"06",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"3F",X"4F",X"33",X"3C",X"0E",X"00",X"00",X"00",X"C0",X"F0",X"FC",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"BF",X"DF",X"67",X"00",X"07",X"03",X"00",X"80",X"C0",X"E0",X"F8",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"7E",X"3C",X"00",X"00",X"00",X"00",X"00",
		X"03",X"0C",X"11",X"27",X"2D",X"49",X"51",X"50",X"50",X"50",X"50",X"28",X"24",X"13",X"0C",X"07",
		X"00",X"20",X"21",X"62",X"65",X"75",X"5D",X"49",X"42",X"6E",X"2C",X"37",X"1B",X"0C",X"07",X"00",
		X"03",X"0C",X"13",X"14",X"28",X"28",X"28",X"2C",X"13",X"0C",X"07",X"80",X"00",X"01",X"0F",X"03",
		X"00",X"00",X"03",X"0C",X"11",X"15",X"2A",X"29",X"28",X"28",X"14",X"17",X"08",X"07",X"00",X"00",
		X"00",X"00",X"08",X"00",X"11",X"1B",X"1E",X"15",X"11",X"0A",X"0D",X"06",X"03",X"00",X"00",X"00",
		X"00",X"00",X"03",X"04",X"0B",X"0A",X"0A",X"0B",X"04",X"03",X"00",X"00",X"04",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"02",X"05",X"02",X"03",X"02",X"05",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0D",X"06",X"05",X"02",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"05",X"05",X"02",X"01",X"00",X"00",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"08",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"07",X"0F",X"0F",X"0E",X"0E",X"0E",X"0E",X"0F",X"07",X"03",X"00",X"00",X"00",X"00",
		X"00",X"03",X"07",X"07",X"0F",X"0F",X"07",X"07",X"07",X"03",X"03",X"01",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"03",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"3F",X"30",X"00",X"00",X"00",X"00",X"05",X"03",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"0C",X"08",X"08",X"02",X"00",X"00",X"00",X"02",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"0C",X"08",X"08",X"02",X"00",X"00",X"00",X"02",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"07",X"2C",X"08",X"08",X"02",X"00",X"00",X"00",X"02",X"02",X"00",X"00",X"00",
		X"00",X"00",X"42",X"02",X"0A",X"0A",X"08",X"02",X"00",X"00",X"00",X"00",X"01",X"03",X"04",X"08",
		X"00",X"00",X"02",X"02",X"0A",X"0A",X"08",X"02",X"00",X"00",X"00",X"00",X"01",X"03",X"04",X"08",
		X"00",X"00",X"02",X"22",X"0A",X"0A",X"08",X"02",X"00",X"00",X"00",X"00",X"01",X"03",X"04",X"08",
		X"00",X"0A",X"01",X"01",X"04",X"08",X"08",X"0B",X"04",X"00",X"02",X"02",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"01",X"01",X"04",X"08",X"08",X"0B",X"04",X"00",X"02",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"3C",X"63",X"D4",X"09",X"49",X"36",X"09",X"09",X"16",X"09",X"00",X"00",X"00",X"00",X"00",
		X"00",X"18",X"3E",X"6B",X"08",X"14",X"08",X"08",X"02",X"00",X"01",X"03",X"03",X"03",X"03",X"01",
		X"00",X"01",X"3B",X"07",X"06",X"02",X"00",X"00",X"00",X"00",X"24",X"0E",X"0E",X"0E",X"0E",X"04",
		X"00",X"03",X"17",X"0F",X"04",X"00",X"00",X"00",X"00",X"40",X"10",X"38",X"38",X"38",X"38",X"10",
		X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"0F",X"0C",X"18",X"1F",X"19",X"1F",X"19",X"14",X"1B",X"0C",X"07",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"3F",X"00",X"00",X"00",X"00",
		X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"FF",X"FF",X"07",X"00",X"F8",X"FF",X"C7",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"FF",X"FF",X"F0",X"00",X"0F",X"FF",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",
		X"FF",X"FF",X"FE",X"00",X"01",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"02",X"02",X"02",X"00",X"02",X"00",X"00",X"00",X"02",X"01",X"03",X"04",X"08",
		X"00",X"00",X"03",X"04",X"04",X"05",X"06",X"06",X"02",X"00",X"00",X"01",X"01",X"01",X"00",X"00",
		X"00",X"00",X"03",X"04",X"04",X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"04",X"04",X"05",X"06",X"06",X"02",X"00",X"00",X"01",X"01",X"01",X"00",X"00",
		X"00",X"F3",X"74",X"1C",X"0F",X"50",X"70",X"3C",X"03",X"01",X"01",X"19",X"3F",X"3E",X"3E",X"1C",
		X"78",X"3B",X"14",X"0C",X"4F",X"70",X"30",X"1C",X"13",X"71",X"F1",X"F1",X"EB",X"70",X"00",X"00",
		X"00",X"F3",X"74",X"1C",X"0F",X"70",X"F0",X"FC",X"F3",X"71",X"01",X"01",X"0B",X"30",X"00",X"00",
		X"E7",X"68",X"BF",X"D7",X"79",X"3C",X"33",X"31",X"41",X"01",X"0B",X"30",X"00",X"00",X"00",X"00",
		X"41",X"E1",X"F1",X"73",X"3C",X"10",X"10",X"0F",X"18",X"14",X"0B",X"18",X"18",X"10",X"00",X"00",
		X"41",X"E1",X"F1",X"73",X"3C",X"10",X"10",X"0F",X"18",X"64",X"E3",X"00",X"00",X"00",X"00",X"00",
		X"00",X"1F",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"02",X"05",X"01",X"00",X"00",X"00",X"00",
		X"00",X"1F",X"00",X"00",X"00",X"00",X"0F",X"0E",X"0E",X"0E",X"05",X"01",X"00",X"00",X"00",X"00",
		X"00",X"1F",X"00",X"3F",X"1A",X"1D",X"0F",X"0E",X"0E",X"0E",X"05",X"01",X"00",X"00",X"00",X"00",
		X"3F",X"7F",X"3F",X"3A",X"1D",X"1F",X"0F",X"0E",X"0E",X"0E",X"07",X"03",X"03",X"03",X"01",X"01",
		X"00",X"1F",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"1F",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"0F",X"1F",X"3F",X"3F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"3F",X"3F",X"1F",X"0F",X"03",
		X"03",X"0F",X"1F",X"3F",X"3F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"3F",X"1F",X"0F",X"03",
		X"03",X"0F",X"1F",X"3F",X"3F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"3F",X"3F",X"1F",X"0F",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"07",X"0F",X"0F",X"0E",X"0E",X"0E",X"0E",X"0F",X"07",X"03",X"00",X"00",X"00",
		X"00",X"00",X"03",X"07",X"07",X"0F",X"0F",X"07",X"07",X"07",X"03",X"03",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"03",X"03",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"04",X"0B",X"16",X"14",X"00",X"14",X"16",X"0B",X"04",X"03",X"00",X"00",X"00",
		X"07",X"0F",X"18",X"37",X"6C",X"68",X"68",X"00",X"68",X"68",X"6C",X"37",X"18",X"0F",X"07",X"00",
		X"00",X"07",X"0F",X"1F",X"3C",X"38",X"38",X"39",X"38",X"38",X"3C",X"1F",X"0F",X"07",X"00",X"00",
		X"00",X"00",X"00",X"07",X"0F",X"0E",X"0C",X"0D",X"0C",X"0E",X"0F",X"07",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"02",X"02",X"02",X"00",X"04",X"00",
		X"00",X"00",X"00",X"00",X"03",X"06",X"06",X"04",X"04",X"00",X"02",X"01",X"01",X"02",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"02",X"04",X"04",X"04",X"0C",X"0C",X"0C",X"0C",X"14",
		X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"02",X"04",X"04",X"04",X"0C",X"0C",X"0C",X"0C",X"14",
		X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"02",X"04",X"04",X"04",X"0C",X"0C",X"0C",X"0C",X"14",
		X"00",X"09",X"06",X"09",X"10",X"09",X"06",X"09",X"70",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"25",X"22",X"12",X"15",X"08",X"05",X"02",X"01",X"00",X"00",X"00",X"00",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"42",X"02",X"02",X"21",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"28",X"20",X"00",X"03",X"06",X"04",X"06",X"05",X"00",X"00",X"00",X"00",
		X"00",X"06",X"00",X"00",X"00",X"00",X"07",X"04",X"00",X"03",X"04",X"04",X"02",X"01",X"02",X"00",
		X"00",X"00",X"00",X"10",X"0D",X"12",X"22",X"25",X"18",X"25",X"02",X"04",X"18",X"00",X"00",X"00",
		X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"00",X"01",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"06",X"07",X"03",X"00",X"00",X"00",X"0A",X"00",
		X"00",X"00",X"00",X"00",X"03",X"00",X"02",X"03",X"03",X"21",X"10",X"00",X"04",X"02",X"02",X"00",
		X"00",X"02",X"04",X"00",X"15",X"20",X"20",X"01",X"02",X"02",X"02",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"73",X"7C",X"F0",X"F0",X"CF",X"18",X"14",X"0B",X"18",X"18",X"10",X"00",X"00",
		X"0E",X"1F",X"1F",X"1F",X"02",X"0A",X"35",X"74",X"02",X"02",X"01",X"00",X"00",X"01",X"01",X"01",
		X"01",X"01",X"01",X"00",X"00",X"01",X"02",X"02",X"74",X"35",X"0A",X"02",X"0F",X"1F",X"1F",X"0E",
		X"00",X"00",X"08",X"0C",X"0C",X"05",X"0A",X"0C",X"67",X"F8",X"F8",X"7E",X"39",X"00",X"00",X"00",
		X"00",X"31",X"79",X"7A",X"7B",X"7C",X"32",X"11",X"11",X"08",X"08",X"1C",X"26",X"03",X"00",X"00",
		X"00",X"00",X"03",X"26",X"1C",X"08",X"08",X"11",X"11",X"32",X"3C",X"3B",X"3E",X"3D",X"19",X"00",
		X"0D",X"06",X"0E",X"06",X"06",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3B",X"3D",X"1D",X"1D",X"1F",X"0F",X"0E",X"0F",X"07",X"06",X"07",X"05",X"01",X"01",X"00",X"00",
		X"0D",X"06",X"06",X"02",X"02",X"03",X"01",X"01",X"03",X"03",X"03",X"0A",X"00",X"01",X"11",X"0E",
		X"3D",X"0D",X"06",X"06",X"03",X"03",X"02",X"00",X"00",X"00",X"00",X"40",X"20",X"32",X"00",X"00",
		X"07",X"00",X"00",X"00",X"00",X"02",X"00",X"20",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"1C",X"00",X"00",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"10",X"17",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1C",X"10",X"00",X"00",
		X"10",X"10",X"10",X"17",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1C",X"10",X"00",X"00",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"00",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"1E",X"3E",X"7E",X"7E",X"FE",X"FE",X"FE",X"FC",X"FC",X"FC",X"FC",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",X"00",X"00",
		X"80",X"00",X"00",X"FF",X"26",X"04",X"55",X"55",X"55",X"55",X"55",X"56",X"FF",X"00",X"00",X"80",
		X"FF",X"FF",X"FF",X"80",X"00",X"00",X"FF",X"26",X"05",X"55",X"55",X"56",X"FF",X"00",X"00",X"80",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"00",X"00",X"04",X"55",X"54",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
