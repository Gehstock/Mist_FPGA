library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ZIGZAG_1H is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ZIGZAG_1H is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",X"00",X"02",X"02",X"FE",X"FE",X"42",X"02",X"00",X"00",
		X"62",X"F2",X"BA",X"9A",X"9E",X"CE",X"46",X"00",X"8C",X"DE",X"F2",X"B2",X"92",X"86",X"04",X"00",
		X"08",X"FE",X"FE",X"C8",X"68",X"38",X"18",X"00",X"1C",X"BE",X"A2",X"A2",X"A2",X"E6",X"E4",X"00",
		X"0C",X"9E",X"92",X"92",X"D2",X"7E",X"3C",X"00",X"C0",X"E0",X"B0",X"9E",X"8E",X"C0",X"C0",X"00",
		X"0C",X"6E",X"9A",X"9A",X"B2",X"F2",X"6C",X"00",X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",X"00",
		X"C0",X"80",X"80",X"C0",X"C0",X"80",X"80",X"C0",X"03",X"01",X"01",X"03",X"03",X"01",X"01",X"03",
		X"FF",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",
		X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",X"44",X"C6",X"82",X"82",X"C6",X"7C",X"38",X"00",
		X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",X"82",X"92",X"92",X"92",X"FE",X"FE",X"00",X"00",
		X"80",X"90",X"90",X"90",X"90",X"FE",X"FE",X"00",X"9E",X"9E",X"92",X"82",X"C6",X"7C",X"38",X"00",
		X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",X"82",X"82",X"FE",X"FE",X"82",X"82",X"00",X"00",
		X"FC",X"FE",X"02",X"02",X"02",X"06",X"04",X"00",X"82",X"C6",X"6E",X"3C",X"18",X"FE",X"FE",X"00",
		X"02",X"02",X"02",X"02",X"FE",X"FE",X"00",X"00",X"FE",X"FE",X"70",X"38",X"70",X"FE",X"FE",X"00",
		X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",X"00",
		X"70",X"F8",X"88",X"88",X"88",X"FE",X"FE",X"00",X"7A",X"FC",X"8E",X"8A",X"82",X"FE",X"7C",X"00",
		X"72",X"F6",X"9E",X"8C",X"88",X"FE",X"FE",X"00",X"0C",X"5E",X"D2",X"92",X"92",X"F6",X"64",X"00",
		X"80",X"80",X"FE",X"FE",X"80",X"80",X"00",X"00",X"FC",X"FE",X"02",X"02",X"02",X"FE",X"FC",X"00",
		X"F0",X"F8",X"1C",X"0E",X"1C",X"F8",X"F0",X"00",X"F8",X"FE",X"1C",X"38",X"1C",X"FE",X"F8",X"00",
		X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",X"C0",X"F0",X"1E",X"1E",X"F0",X"C0",X"00",X"00",
		X"C2",X"E2",X"F2",X"BA",X"9E",X"8E",X"86",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"9B",X"FF",X"FF",X"9B",X"01",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"1F",X"1F",X"3F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"3F",X"1F",X"1F",X"3F",
		X"0F",X"07",X"07",X"0F",X"0F",X"1F",X"BF",X"FF",X"FF",X"BF",X"1F",X"0F",X"0F",X"07",X"07",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"80",X"D9",X"FF",X"FF",X"D9",X"80",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"F8",X"F8",X"FC",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"FC",X"F8",X"F8",X"FC",
		X"F0",X"E0",X"E0",X"F0",X"F0",X"F8",X"FD",X"FF",X"FF",X"FD",X"F8",X"F0",X"F0",X"E0",X"E0",X"F0",
		X"C0",X"80",X"80",X"C0",X"C0",X"80",X"C0",X"E0",X"03",X"01",X"01",X"03",X"03",X"01",X"03",X"07",
		X"C0",X"E0",X"F9",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"07",X"9F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"80",X"C0",X"E0",X"F9",X"FF",X"FF",X"FF",X"03",X"01",X"03",X"07",X"9F",X"FF",X"FF",X"FF",
		X"E0",X"C0",X"80",X"C0",X"C0",X"80",X"80",X"C0",X"07",X"03",X"01",X"03",X"03",X"01",X"01",X"03",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F9",X"E0",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"9F",X"07",X"03",
		X"FF",X"FF",X"FF",X"F9",X"E0",X"C0",X"80",X"C0",X"FF",X"FF",X"FF",X"9F",X"07",X"03",X"01",X"03",
		X"C0",X"80",X"80",X"C0",X"C0",X"E0",X"F9",X"FF",X"03",X"01",X"01",X"03",X"03",X"07",X"9F",X"FF",
		X"FF",X"F9",X"E0",X"C0",X"C0",X"80",X"80",X"C0",X"FF",X"9F",X"07",X"03",X"03",X"01",X"01",X"03",
		X"C0",X"80",X"80",X"C0",X"C0",X"80",X"80",X"C0",X"03",X"01",X"01",X"03",X"03",X"01",X"01",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"FF",X"FF",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"60",X"30",X"18",X"0C",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"40",X"60",X"C0",X"80",X"C0",X"C0",
		X"0F",X"3B",X"10",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"05",X"07",X"27",X"3F",X"00",X"00",X"00",X"00",X"08",X"D8",X"E0",X"C0",
		X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"05",X"02",X"07",X"2F",X"3B",X"00",X"00",X"00",X"88",X"C8",X"F0",X"C0",X"C0",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"13",X"1F",X"00",X"00",X"00",X"00",X"40",X"40",X"E4",X"FC",
		X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"E0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"38",X"70",X"F7",X"FF",X"00",X"00",X"FC",X"20",X"70",X"E0",X"FC",X"F0",
		X"F7",X"70",X"38",X"00",X"00",X"00",X"00",X"00",X"FC",X"E0",X"70",X"20",X"FC",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"0C",X"7F",X"00",X"00",X"00",X"18",X"08",X"1C",X"FE",X"F8",
		X"0C",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"1C",X"08",X"18",X"00",X"00",X"00",X"00",
		X"02",X"07",X"07",X"0F",X"0F",X"0F",X"1F",X"18",X"00",X"00",X"00",X"80",X"80",X"80",X"C0",X"C0",
		X"17",X"37",X"38",X"3F",X"70",X"7F",X"7F",X"00",X"40",X"60",X"E0",X"E0",X"70",X"F0",X"F0",X"00",
		X"02",X"02",X"07",X"07",X"0F",X"0F",X"1F",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"00",
		X"C3",X"FF",X"FF",X"7E",X"00",X"00",X"C3",X"C3",X"00",X"00",X"7E",X"FF",X"FF",X"C3",X"C3",X"C3",
		X"00",X"01",X"03",X"07",X"03",X"07",X"0F",X"3F",X"80",X"80",X"D8",X"F8",X"F8",X"F0",X"F0",X"F0",
		X"1F",X"1F",X"1F",X"0F",X"03",X"07",X"07",X"01",X"F8",X"F8",X"F0",X"E0",X"F8",X"FC",X"78",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"90",
		X"07",X"02",X"02",X"08",X"00",X"00",X"00",X"00",X"C0",X"80",X"A0",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"24",X"04",X"4E",X"27",X"00",X"00",X"20",X"40",X"11",X"80",X"A4",X"C8",
		X"07",X"03",X"25",X"00",X"08",X"00",X"00",X"00",X"C0",X"20",X"90",X"A0",X"20",X"50",X"00",X"00",
		X"00",X"00",X"42",X"20",X"04",X"0F",X"E7",X"3F",X"00",X"20",X"44",X"C8",X"80",X"80",X"D0",X"EC",
		X"07",X"07",X"0D",X"1D",X"29",X"42",X"01",X"00",X"C0",X"A0",X"B0",X"88",X"44",X"20",X"10",X"08",
		X"3C",X"62",X"95",X"A5",X"A5",X"99",X"42",X"3F",X"C0",X"20",X"20",X"20",X"C0",X"00",X"C0",X"20",
		X"0A",X"0A",X"0E",X"00",X"00",X"0F",X"04",X"00",X"20",X"20",X"40",X"00",X"20",X"E0",X"20",X"00",
		X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"C0",X"20",X"20",X"C0",X"00",X"C0",X"20",X"20",
		X"07",X"00",X"06",X"09",X"08",X"08",X"04",X"00",X"C0",X"00",X"20",X"20",X"A0",X"60",X"20",X"00",
		X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"C0",X"20",X"20",X"C0",X"00",X"C0",X"20",X"20",
		X"07",X"00",X"08",X"0D",X"0B",X"09",X"08",X"00",X"C0",X"00",X"C0",X"20",X"20",X"20",X"20",X"00",
		X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"C0",X"20",X"20",X"C0",X"00",X"C0",X"20",X"20",
		X"07",X"00",X"06",X"09",X"09",X"09",X"06",X"00",X"C0",X"00",X"C0",X"20",X"20",X"20",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"07",X"08",X"08",X"07",X"00",X"00",X"00",X"00",X"C0",X"20",X"20",X"C0",
		X"00",X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"00",X"C0",X"20",X"20",X"C0",X"00",X"C0",X"20",
		X"08",X"07",X"00",X"00",X"0F",X"04",X"00",X"00",X"20",X"C0",X"00",X"20",X"E0",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"07",X"00",X"06",X"09",X"08",X"08",X"04",X"20",X"C0",X"00",X"20",X"20",X"A0",X"60",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"07",X"00",X"00",X"0F",X"40",X"20",X"10",X"20",X"C0",X"00",X"40",X"E0",X"40",X"40",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"07",X"00",X"06",X"09",X"09",X"09",X"06",X"20",X"C0",X"00",X"C0",X"20",X"20",X"20",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"07",X"00",X"00",X"09",X"09",X"09",X"07",X"20",X"C0",X"00",X"C0",X"20",X"20",X"20",X"C0",
		X"00",X"00",X"0F",X"04",X"00",X"00",X"00",X"00",X"00",X"20",X"E0",X"20",X"00",X"00",X"00",X"00",
		X"08",X"07",X"00",X"06",X"09",X"08",X"08",X"04",X"20",X"C0",X"00",X"20",X"20",X"A0",X"60",X"20",
		X"00",X"0C",X"0B",X"09",X"00",X"00",X"00",X"00",X"00",X"C0",X"20",X"20",X"20",X"40",X"00",X"00",
		X"FE",X"FC",X"F1",X"C1",X"80",X"AD",X"B7",X"9F",X"0F",X"E3",X"09",X"81",X"01",X"61",X"F1",X"F9",
		X"C7",X"F0",X"F6",X"EF",X"ED",X"E3",X"F8",X"FF",X"31",X"B1",X"F3",X"E1",X"E1",X"B9",X"79",X"03",
		X"00",X"00",X"01",X"01",X"00",X"2D",X"37",X"1F",X"00",X"E0",X"08",X"80",X"00",X"60",X"F0",X"F8",
		X"07",X"00",X"06",X"0F",X"0D",X"03",X"00",X"00",X"30",X"B0",X"F2",X"E0",X"E0",X"B8",X"78",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"05",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"78",
		X"0B",X"06",X"01",X"00",X"00",X"00",X"00",X"00",X"86",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"08",X"0C",X"06",X"3A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"0E",X"1C",X"38",X"10",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"07",X"00",X"00",X"18",X"10",X"1C",X"0E",X"06",X"32",
		X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CE",X"02",X"0E",X"1E",X"1C",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"8C",X"8C",X"58",X"58",X"30",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"30",X"58",X"58",X"8C",X"8C",X"00",X"00",
		X"00",X"00",X"00",X"03",X"06",X"06",X"03",X"01",X"00",X"00",X"00",X"E0",X"C0",X"C0",X"E0",X"C0",
		X"01",X"03",X"06",X"06",X"03",X"00",X"00",X"00",X"C0",X"E0",X"30",X"30",X"E0",X"00",X"00",X"00",
		X"00",X"00",X"20",X"20",X"10",X"18",X"0C",X"0E",X"00",X"00",X"00",X"20",X"20",X"64",X"CC",X"7C",
		X"04",X"0C",X"0C",X"04",X"00",X"00",X"00",X"00",X"3C",X"38",X"3C",X"3C",X"0C",X"38",X"00",X"00",
		X"00",X"00",X"00",X"03",X"07",X"07",X"07",X"02",X"00",X"00",X"38",X"E0",X"E0",X"E4",X"EC",X"40",
		X"02",X"07",X"07",X"07",X"03",X"00",X"00",X"00",X"40",X"EC",X"E4",X"E0",X"E0",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"0D",X"02",X"04",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"02",X"62",X"27",X"10",X"E6",X"92",X"0C",X"68",X"20",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"61",X"13",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"12",X"04",X"F1",X"52",X"31",X"36",X"05",X"04",X"C0",X"20",X"A0",X"20",X"20",X"40",X"40",X"80",
		X"05",X"04",X"02",X"01",X"00",X"01",X"01",X"01",X"C0",X"40",X"40",X"40",X"C0",X"C0",X"FC",X"8A",
		X"01",X"06",X"08",X"00",X"00",X"00",X"00",X"00",X"72",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"02",X"00",X"78",X"20",X"20",X"10",X"10",X"20",X"20",
		X"13",X"0F",X"E3",X"00",X"00",X"00",X"00",X"00",X"70",X"D0",X"10",X"0C",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"04",X"04",X"1C",X"00",X"00",X"00",X"00",X"04",X"B4",X"FC",X"FC",
		X"1C",X"0D",X"0F",X"07",X"03",X"00",X"00",X"00",X"C0",X"C4",X"94",X"9C",X"8C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"09",X"09",X"39",X"00",X"00",X"00",X"00",X"00",X"7C",X"FC",X"F4",
		X"39",X"1B",X"1F",X"0F",X"07",X"00",X"00",X"00",X"F4",X"3C",X"1C",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"02",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"40",X"20",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"40",X"40",X"20",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"02",X"02",X"40",X"40",X"80",X"80",X"00",X"00",X"00",X"00",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"40",X"40",X"20",X"20",
		X"00",X"00",X"00",X"00",X"01",X"01",X"02",X"02",X"40",X"40",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"40",X"40",X"20",X"20",
		X"00",X"00",X"00",X"00",X"01",X"01",X"02",X"02",X"40",X"40",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"18",X"04",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"0C",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"30",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"0C",X"03",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0C",
		X"30",X"0C",X"03",X"00",X"00",X"00",X"00",X"00",X"30",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"FE",X"38",X"10",X"10",X"00",X"3C",
		X"3C",X"3F",X"3F",X"39",X"0F",X"0F",X"00",X"00",X"08",X"08",X"08",X"20",X"20",X"60",X"60",X"00",
		X"00",X"00",X"00",X"30",X"0C",X"00",X"00",X"00",X"00",X"00",X"38",X"0C",X"00",X"00",X"00",X"38",
		X"3E",X"3F",X"37",X"3B",X"3F",X"1F",X"00",X"00",X"0C",X"04",X"00",X"20",X"20",X"60",X"60",X"00",
		X"00",X"0C",X"0C",X"06",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"7C",X"F7",X"C3",X"77",X"1E",X"00",X"01",X"21",X"20",X"20",X"20",X"E0",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"12",X"00",X"00",X"00",X"00",X"00",X"01",
		X"3E",X"7E",X"F3",X"F3",X"CF",X"CF",X"7E",X"38",X"01",X"00",X"30",X"30",X"70",X"70",X"70",X"00",
		X"00",X"01",X"06",X"0A",X"16",X"1F",X"0E",X"0C",X"00",X"80",X"00",X"00",X"04",X"84",X"C0",X"40",
		X"0E",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"C0",X"C4",X"CC",X"E0",X"60",X"10",X"70",X"00",
		X"06",X"00",X"0E",X"1E",X"36",X"2F",X"3F",X"1E",X"00",X"08",X"0C",X"00",X"00",X"C0",X"E0",X"E2",
		X"1C",X"0E",X"07",X"03",X"00",X"00",X"00",X"00",X"66",X"E6",X"E0",X"F0",X"3C",X"12",X"06",X"00",
		X"00",X"30",X"10",X"78",X"FE",X"EF",X"C7",X"6E",X"00",X"03",X"03",X"03",X"00",X"80",X"C0",X"E3",
		X"7E",X"38",X"1E",X"0E",X"07",X"03",X"00",X"00",X"F3",X"37",X"F7",X"E0",X"EC",X"F6",X"36",X"06",
		X"00",X"00",X"00",X"00",X"78",X"FE",X"DF",X"8F",X"00",X"00",X"01",X"01",X"01",X"00",X"80",X"E0",
		X"DC",X"F8",X"78",X"3C",X"3C",X"1F",X"0F",X"07",X"F1",X"F1",X"39",X"39",X"F8",X"F0",X"E0",X"9C",
		X"00",X"00",X"00",X"08",X"00",X"08",X"00",X"00",X"00",X"00",X"84",X"1C",X"80",X"10",X"18",X"0C",
		X"00",X"0E",X"1F",X"19",X"09",X"07",X"00",X"00",X"04",X"40",X"70",X"78",X"70",X"38",X"30",X"00",
		X"00",X"00",X"00",X"02",X"04",X"02",X"04",X"02",X"00",X"00",X"00",X"38",X"18",X"0C",X"04",X"00",
		X"00",X"00",X"0E",X"1F",X"13",X"09",X"07",X"00",X"38",X"18",X"0C",X"64",X"C0",X"60",X"00",X"00",
		X"00",X"0F",X"1F",X"19",X"1F",X"1F",X"19",X"1F",X"00",X"84",X"C4",X"C4",X"9C",X"84",X"C0",X"C4",
		X"1F",X"1F",X"0F",X"06",X"06",X"00",X"00",X"00",X"C4",X"9C",X"04",X"20",X"20",X"E0",X"00",X"00",
		X"00",X"3E",X"7F",X"67",X"7E",X"7E",X"67",X"7F",X"00",X"00",X"40",X"60",X"30",X"00",X"00",X"40",
		X"7F",X"7E",X"3C",X"18",X"18",X"00",X"00",X"00",X"60",X"30",X"00",X"80",X"80",X"E0",X"00",X"00",
		X"00",X"00",X"30",X"1C",X"17",X"09",X"07",X"00",X"00",X"00",X"F8",X"CC",X"64",X"24",X"24",X"68",
		X"00",X"07",X"09",X"17",X"1C",X"30",X"00",X"00",X"68",X"2C",X"24",X"64",X"CC",X"F8",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"09",X"33",X"3C",X"00",X"00",X"00",X"3C",X"24",X"24",X"6C",X"68",X"C8",
		X"00",X"3C",X"33",X"09",X"0F",X"00",X"00",X"00",X"C8",X"68",X"6C",X"24",X"24",X"3C",X"00",X"00",
		X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"C0",X"20",X"20",X"C0",X"00",X"C0",X"20",X"20",
		X"07",X"00",X"06",X"09",X"08",X"08",X"04",X"00",X"C0",X"00",X"20",X"20",X"A0",X"60",X"20",X"00",
		X"00",X"01",X"03",X"07",X"03",X"07",X"0F",X"3F",X"80",X"80",X"D8",X"F8",X"F8",X"F0",X"F0",X"F0",
		X"1F",X"1F",X"1F",X"0F",X"03",X"07",X"07",X"01",X"F8",X"F8",X"F0",X"E0",X"F8",X"FC",X"78",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"1F",X"04",X"0E",X"0C",X"3E",X"30",X"60",
		X"00",X"00",X"01",X"01",X"01",X"03",X"02",X"02",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",
		X"0D",X"08",X"00",X"00",X"00",X"00",X"00",X"07",X"FC",X"FD",X"7B",X"76",X"EF",X"77",X"7B",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3D",X"18",X"1E",X"1E",X"3D",X"7D",X"0E",X"07",
		X"00",X"00",X"08",X"08",X"38",X"1C",X"2F",X"07",X"00",X"08",X"0C",X"1E",X"18",X"1B",X"93",X"E7",
		X"01",X"00",X"19",X"06",X"00",X"00",X"11",X"1F",X"FE",X"BE",X"F0",X"EF",X"F0",X"FC",X"FD",X"F1",
		X"07",X"08",X"08",X"08",X"07",X"00",X"09",X"0A",X"C0",X"20",X"20",X"20",X"C0",X"00",X"C0",X"20",
		X"0A",X"0A",X"0E",X"00",X"00",X"0F",X"04",X"00",X"20",X"20",X"40",X"00",X"20",X"E0",X"20",X"00",
		X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"C0",X"20",X"20",X"C0",X"00",X"C0",X"20",X"20",
		X"07",X"00",X"06",X"09",X"08",X"08",X"04",X"00",X"C0",X"00",X"20",X"20",X"A0",X"60",X"20",X"00",
		X"00",X"00",X"00",X"0A",X"0E",X"03",X"00",X"00",X"04",X"60",X"88",X"F8",X"F8",X"1C",X"0C",X"04",
		X"00",X"00",X"00",X"00",X"06",X"01",X"00",X"00",X"00",X"00",X"66",X"0C",X"7C",X"98",X"70",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"0C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"12",X"04",X"04",X"02",X"00",X"02",X"00",
		X"00",X"00",X"00",X"00",X"07",X"08",X"08",X"07",X"00",X"00",X"00",X"00",X"C0",X"20",X"20",X"C0",
		X"00",X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"00",X"C0",X"20",X"20",X"C0",X"00",X"C0",X"20",
		X"08",X"07",X"00",X"00",X"0F",X"04",X"00",X"00",X"20",X"C0",X"00",X"20",X"E0",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"07",X"00",X"06",X"09",X"08",X"08",X"04",X"20",X"C0",X"00",X"20",X"20",X"A0",X"60",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"07",X"00",X"00",X"0F",X"04",X"02",X"01",X"20",X"C0",X"00",X"40",X"E0",X"40",X"40",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"07",X"00",X"06",X"09",X"09",X"09",X"06",X"20",X"C0",X"00",X"C0",X"20",X"20",X"20",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"07",X"00",X"00",X"09",X"09",X"09",X"07",X"20",X"C0",X"00",X"C0",X"20",X"20",X"20",X"C0",
		X"00",X"00",X"0F",X"04",X"00",X"00",X"00",X"00",X"00",X"20",X"E0",X"20",X"00",X"00",X"00",X"00",
		X"08",X"07",X"00",X"06",X"09",X"08",X"08",X"04",X"20",X"C0",X"00",X"20",X"20",X"A0",X"60",X"20",
		X"00",X"0C",X"0B",X"09",X"00",X"00",X"00",X"00",X"00",X"C0",X"20",X"20",X"20",X"40",X"00",X"00",
		X"FE",X"FC",X"F1",X"C1",X"80",X"AD",X"B7",X"9F",X"0F",X"E3",X"09",X"81",X"01",X"61",X"F1",X"F9",
		X"C7",X"F0",X"F6",X"EF",X"ED",X"E3",X"F8",X"FF",X"31",X"B1",X"F3",X"E1",X"E1",X"B9",X"79",X"03",
		X"00",X"00",X"01",X"01",X"00",X"2D",X"37",X"1F",X"00",X"E0",X"08",X"80",X"00",X"60",X"F0",X"F8",
		X"07",X"00",X"06",X"0F",X"0D",X"03",X"00",X"00",X"30",X"B0",X"F2",X"E0",X"E0",X"B8",X"78",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"05",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"78",
		X"0B",X"06",X"01",X"00",X"00",X"00",X"00",X"00",X"86",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"08",X"0C",X"06",X"3A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"0E",X"1C",X"38",X"10",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"07",X"00",X"00",X"18",X"10",X"1C",X"0E",X"06",X"32",
		X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CE",X"02",X"0E",X"1E",X"1C",X"10",X"00",X"00",
		X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"C0",X"20",X"20",X"C0",X"00",X"C0",X"20",X"20",
		X"07",X"00",X"08",X"0D",X"0B",X"09",X"08",X"00",X"C0",X"00",X"C0",X"20",X"20",X"20",X"40",X"00",
		X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"C0",X"20",X"20",X"C0",X"00",X"C0",X"20",X"20",
		X"07",X"00",X"00",X"0F",X"04",X"02",X"01",X"00",X"C0",X"00",X"40",X"E0",X"40",X"40",X"40",X"C0",
		X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"C0",X"20",X"20",X"C0",X"00",X"C0",X"20",X"20",
		X"07",X"00",X"09",X"0A",X"0A",X"0A",X"0E",X"00",X"C0",X"00",X"C0",X"20",X"20",X"20",X"40",X"00",
		X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"C0",X"20",X"20",X"C0",X"00",X"C0",X"20",X"20",
		X"07",X"00",X"07",X"08",X"08",X"07",X"00",X"0F",X"C0",X"00",X"C0",X"20",X"20",X"C0",X"00",X"E0",
		X"00",X"00",X"03",X"0F",X"1F",X"00",X"00",X"20",X"00",X"00",X"80",X"E0",X"F0",X"18",X"18",X"38",
		X"63",X"C7",X"FF",X"C7",X"62",X"2E",X"00",X"00",X"C0",X"80",X"98",X"F4",X"1C",X"04",X"00",X"00",
		X"00",X"01",X"03",X"07",X"0F",X"00",X"00",X"00",X"70",X"FC",X"26",X"30",X"38",X"2C",X"2C",X"3C",
		X"01",X"03",X"03",X"03",X"01",X"07",X"00",X"00",X"C8",X"C0",X"FC",X"FC",X"08",X"38",X"00",X"00",
		X"00",X"00",X"01",X"08",X"18",X"18",X"38",X"38",X"70",X"F8",X"AC",X"20",X"24",X"74",X"FC",X"F0",
		X"38",X"18",X"19",X"0F",X"07",X"00",X"00",X"00",X"F0",X"90",X"10",X"78",X"28",X"1C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"18",X"38",X"78",X"00",X"00",X"00",X"00",X"00",X"04",X"74",X"FC",
		X"78",X"F8",X"FF",X"D9",X"4F",X"67",X"20",X"00",X"F0",X"F0",X"34",X"34",X"3C",X"30",X"00",X"00",
		X"00",X"00",X"03",X"0F",X"1F",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"F0",X"18",X"18",X"38",
		X"13",X"37",X"7F",X"37",X"12",X"0E",X"00",X"00",X"C0",X"80",X"98",X"F4",X"1C",X"04",X"00",X"00",
		X"00",X"00",X"01",X"07",X"0F",X"00",X"00",X"00",X"00",X"00",X"C0",X"F0",X"F8",X"0C",X"0C",X"1C",
		X"07",X"0F",X"1F",X"0F",X"05",X"07",X"00",X"00",X"F0",X"E0",X"E4",X"F8",X"08",X"38",X"00",X"00",
		X"00",X"00",X"00",X"08",X"18",X"18",X"38",X"38",X"00",X"20",X"70",X"F8",X"24",X"74",X"FC",X"F0",
		X"38",X"18",X"19",X"0F",X"07",X"00",X"00",X"00",X"F0",X"90",X"10",X"38",X"28",X"1C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"18",X"18",X"38",X"00",X"00",X"00",X"20",X"70",X"FC",X"F4",X"FC",
		X"38",X"38",X"18",X"18",X"0F",X"07",X"00",X"00",X"F0",X"F0",X"F4",X"94",X"1C",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"60",X"E6",
		X"11",X"31",X"31",X"71",X"71",X"73",X"3E",X"1C",X"FC",X"FC",X"F8",X"F0",X"E0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"30",X"33",X"13",X"1A",X"1E",X"1E",
		X"02",X"06",X"06",X"0E",X"0E",X"0E",X"07",X"03",X"3C",X"3C",X"3C",X"38",X"20",X"70",X"C0",X"80",
		X"00",X"01",X"01",X"00",X"00",X"01",X"01",X"01",X"00",X"20",X"B0",X"90",X"F0",X"F0",X"F8",X"F8",
		X"00",X"00",X"00",X"00",X"03",X"01",X"00",X"00",X"F0",X"18",X"0C",X"0C",X"FC",X"F8",X"70",X"00",
		X"00",X"00",X"00",X"08",X"04",X"02",X"00",X"1C",X"00",X"00",X"80",X"88",X"90",X"20",X"00",X"1C",
		X"00",X"02",X"04",X"08",X"00",X"00",X"00",X"00",X"00",X"20",X"90",X"88",X"80",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
