library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity prom_ic24 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of prom_ic24 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"10",X"38",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"00",X"00",X"44",X"10",X"10",X"40",X"00",X"00",X"00",X"00",X"00",X"08",X"40",X"00",X"90",X"94",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"80",X"40",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"80",X"C0",X"64",X"32",X"19",X"0F",X"07",X"07",X"0D",X"19",X"32",X"64",X"C0",X"80",X"00",
		X"80",X"20",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"40",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"05",X"0A",X"14",X"28",X"40",X"80",X"00",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",
		X"18",X"1B",X"03",X"00",X"08",X"08",X"01",X"00",X"00",X"00",X"02",X"01",X"21",X"04",X"41",X"41",
		X"04",X"00",X"15",X"00",X"44",X"28",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"01",
		X"07",X"0D",X"18",X"30",X"60",X"C8",X"D0",X"E0",X"E0",X"D0",X"C8",X"60",X"30",X"18",X"0D",X"07",
		X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"05",
		X"02",X"04",X"08",X"10",X"28",X"50",X"A0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"77",X"00",X"77",X"00",X"77",
		X"77",X"00",X"77",X"00",X"77",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",
		X"0F",X"F8",X"00",X"77",X"07",X"70",X"07",X"70",X"70",X"07",X"70",X"07",X"77",X"00",X"F8",X"0F",
		X"F0",X"1F",X"00",X"77",X"07",X"77",X"00",X"70",X"70",X"00",X"77",X"07",X"77",X"00",X"1F",X"F0",
		X"20",X"20",X"20",X"20",X"F0",X"F0",X"F0",X"F0",X"02",X"02",X"02",X"02",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"18",X"7E",X"7E",X"18",X"18",X"00",
		X"01",X"03",X"01",X"01",X"07",X"03",X"01",X"03",X"1F",X"03",X"1F",X"0F",X"07",X"1F",X"03",X"0F",
		X"7F",X"0F",X"7F",X"3F",X"0F",X"7F",X"1F",X"3F",X"FF",X"3F",X"7F",X"FF",X"3F",X"FF",X"3F",X"7F",
		X"00",X"0E",X"00",X"0E",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"0E",X"00",X"0E",X"00",X"0E",
		X"0E",X"00",X"0E",X"00",X"0E",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"0E",X"00",X"0E",X"00",
		X"0F",X"F8",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"F8",X"0F",
		X"F0",X"1F",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"1F",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"20",X"20",X"20",X"20",X"0F",X"0F",X"0F",X"0F",X"02",X"02",X"02",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"18",X"00",X"00",X"18",X"18",X"00",
		X"FF",X"FF",X"7E",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"7E",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",
		X"60",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"60",
		X"00",X"60",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"00",
		X"00",X"60",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"00",X"00",
		X"07",X"0C",X"38",X"60",X"C6",X"6C",X"38",X"00",X"00",X"38",X"6C",X"C6",X"60",X"38",X"0C",X"07",
		X"07",X"1C",X"70",X"C0",X"80",X"D8",X"70",X"00",X"00",X"70",X"D8",X"80",X"C0",X"70",X"1C",X"07",
		X"07",X"1C",X"70",X"C0",X"80",X"C0",X"60",X"00",X"00",X"60",X"C0",X"80",X"C0",X"70",X"1C",X"07",
		X"07",X"3C",X"60",X"C0",X"80",X"80",X"80",X"00",X"00",X"80",X"80",X"80",X"C0",X"60",X"3C",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"10",X"00",X"00",X"00",
		X"10",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",
		X"00",X"38",X"44",X"9A",X"82",X"9A",X"44",X"38",X"44",X"9A",X"82",X"9A",X"44",X"38",X"00",X"00",
		X"82",X"9A",X"44",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"44",X"9A",
		X"44",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"44",X"9A",X"82",X"9A",
		X"3C",X"42",X"99",X"81",X"81",X"99",X"42",X"3C",X"99",X"81",X"81",X"99",X"42",X"3C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"42",X"81",X"99",X"42",X"3C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"3C",X"42",X"99",X"81",X"42",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"3C",X"42",X"99",X"81",X"81",X"99",X"01",X"31",X"32",X"02",X"8C",X"70",X"00",X"00",
		X"00",X"00",X"00",X"70",X"8C",X"02",X"32",X"31",X"04",X"04",X"02",X"02",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"02",X"02",X"04",X"01",X"31",X"32",X"02",X"04",X"08",X"F0",X"00",
		X"00",X"00",X"F0",X"08",X"04",X"02",X"32",X"31",X"08",X"08",X"04",X"1C",X"02",X"01",X"00",X"00",
		X"00",X"00",X"00",X"01",X"02",X"1C",X"04",X"08",X"80",X"30",X"30",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"30",X"01",X"00",X"20",X"3C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"3C",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"20",X"30",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"70",X"60",
		X"03",X"60",X"70",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1E",X"70",X"60",
		X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"B0",X"80",X"B0",
		X"70",X"1E",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"1E",X"70",X"01",X"03",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"B0",X"80",X"B0",X"B0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"60",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"1E",X"31",X"63",X"07",X"33",X"31",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"B0",X"80",X"B0",X"B0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"01",X"03",X"01",X"70",X"1E",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"1E",
		X"00",X"60",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"60",
		X"0F",X"07",X"03",X"18",X"F0",X"60",X"C0",X"00",X"00",X"00",X"C0",X"60",X"F0",X"18",X"03",X"07",
		X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"00",X"60",
		X"02",X"18",X"F8",X"30",X"E0",X"00",X"00",X"00",X"E0",X"30",X"F8",X"18",X"02",X"06",X"0E",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"00",X"60",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"F0",X"20",X"E0",X"00",X"00",X"00",X"00",
		X"38",X"18",X"02",X"06",X"06",X"06",X"02",X"18",X"00",X"00",X"00",X"00",X"00",X"E0",X"20",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"00",X"60",X"60",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"06",X"0E",X"06",X"02",X"E8",X"38",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"38",X"E8",X"80",X"B0",X"30",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"B0",X"03",X"01",X"60",X"3E",X"60",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"60",X"3E",X"60",X"01",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
