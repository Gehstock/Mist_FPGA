library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_1L is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_1L is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"CD",X"05",X"22",X"3A",X"8D",X"80",X"FE",X"00",X"20",X"0A",X"3A",X"28",X"80",X"CB",X"57",X"20",
		X"03",X"CD",X"C0",X"20",X"3A",X"53",X"84",X"E6",X"03",X"FE",X"03",X"28",X"17",X"3A",X"A7",X"81",
		X"B7",X"FE",X"14",X"38",X"15",X"3E",X"00",X"32",X"A7",X"81",X"3E",X"03",X"32",X"53",X"84",X"3E",
		X"1B",X"CD",X"FC",X"00",X"CD",X"4B",X"23",X"CD",X"C9",X"00",X"3A",X"00",X"89",X"CB",X"47",X"28",
		X"06",X"CD",X"33",X"25",X"CD",X"C9",X"00",X"3A",X"60",X"84",X"FE",X"00",X"28",X"17",X"3D",X"32",
		X"60",X"84",X"FE",X"00",X"20",X"0F",X"21",X"00",X"00",X"22",X"08",X"85",X"22",X"0A",X"85",X"22",
		X"0C",X"85",X"22",X"0E",X"85",X"3A",X"02",X"89",X"FE",X"FF",X"28",X"16",X"3A",X"13",X"89",X"FE",
		X"00",X"28",X"3C",X"3D",X"32",X"13",X"89",X"FE",X"00",X"20",X"34",X"3A",X"0C",X"89",X"FE",X"02",
		X"20",X"0A",X"CD",X"36",X"60",X"3A",X"02",X"89",X"FE",X"FF",X"28",X"23",X"21",X"00",X"00",X"22",
		X"10",X"85",X"22",X"12",X"85",X"22",X"14",X"85",X"22",X"16",X"85",X"3A",X"0C",X"89",X"FE",X"03",
		X"20",X"08",X"3E",X"01",X"32",X"80",X"80",X"32",X"77",X"80",X"3E",X"00",X"32",X"0C",X"89",X"3A",
		X"8D",X"80",X"FE",X"00",X"CA",X"C3",X"00",X"3A",X"28",X"80",X"CB",X"57",X"C2",X"C3",X"00",X"C9",
		X"3A",X"28",X"80",X"CB",X"57",X"C2",X"75",X"21",X"DD",X"21",X"A2",X"81",X"FD",X"21",X"80",X"84",
		X"3A",X"A2",X"81",X"FE",X"00",X"CA",X"5D",X"21",X"FD",X"CB",X"00",X"76",X"C2",X"4B",X"21",X"3A",
		X"02",X"85",X"16",X"00",X"5F",X"21",X"08",X"00",X"19",X"54",X"5D",X"26",X"00",X"FD",X"6E",X"01",
		X"01",X"08",X"00",X"09",X"B7",X"ED",X"52",X"CD",X"F0",X"1F",X"11",X"0A",X"00",X"B7",X"ED",X"52",
		X"D2",X"4B",X"21",X"3A",X"03",X"85",X"16",X"00",X"5F",X"21",X"08",X"00",X"19",X"54",X"5D",X"26",
		X"00",X"FD",X"6E",X"02",X"01",X"08",X"00",X"09",X"B7",X"ED",X"52",X"CD",X"F0",X"1F",X"11",X"08",
		X"00",X"B7",X"ED",X"52",X"D2",X"4B",X"21",X"CD",X"76",X"21",X"3A",X"53",X"84",X"E6",X"03",X"FE",
		X"03",X"28",X"0A",X"3A",X"28",X"80",X"CB",X"7F",X"20",X"03",X"CD",X"06",X"29",X"CD",X"CF",X"22",
		X"3A",X"A2",X"81",X"FE",X"00",X"CA",X"5D",X"21",X"C3",X"75",X"21",X"FD",X"7E",X"00",X"E6",X"3F",
		X"FE",X"17",X"CA",X"75",X"21",X"11",X"05",X"00",X"FD",X"19",X"C3",X"D8",X"20",X"3A",X"70",X"80",
		X"FE",X"00",X"28",X"0A",X"3E",X"01",X"32",X"74",X"80",X"32",X"77",X"80",X"18",X"07",X"3E",X"01",
		X"32",X"78",X"80",X"18",X"00",X"C9",X"C5",X"DD",X"E5",X"FD",X"E5",X"FD",X"36",X"04",X"00",X"01",
		X"00",X"01",X"3E",X"19",X"FD",X"CB",X"00",X"7E",X"28",X"10",X"01",X"00",X"02",X"3A",X"AB",X"81",
		X"3C",X"32",X"AB",X"81",X"FD",X"36",X"04",X"01",X"3E",X"18",X"CD",X"FC",X"00",X"CD",X"E4",X"00",
		X"FD",X"46",X"01",X"FD",X"4E",X"02",X"CD",X"DE",X"00",X"E5",X"DD",X"E1",X"DD",X"36",X"00",X"86",
		X"DD",X"36",X"01",X"87",X"11",X"E0",X"FF",X"DD",X"19",X"DD",X"36",X"00",X"84",X"DD",X"36",X"01",
		X"85",X"FD",X"CB",X"00",X"F6",X"FD",X"36",X"03",X"01",X"3A",X"A2",X"81",X"FE",X"00",X"28",X"01",
		X"3D",X"32",X"A2",X"81",X"3A",X"A7",X"81",X"3C",X"FD",X"CB",X"00",X"7E",X"28",X"0C",X"3C",X"4F",
		X"FD",X"CB",X"00",X"BE",X"3E",X"00",X"32",X"A6",X"81",X"79",X"4F",X"3A",X"53",X"84",X"E6",X"03",
		X"FE",X"03",X"28",X"0B",X"3A",X"28",X"80",X"CB",X"7F",X"20",X"04",X"79",X"32",X"A7",X"81",X"FD",
		X"E1",X"DD",X"E1",X"C1",X"C9",X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",X"DD",X"21",X"80",X"84",
		X"DD",X"7E",X"00",X"FE",X"FF",X"CA",X"C7",X"22",X"DD",X"CB",X"00",X"76",X"CA",X"BC",X"22",X"DD",
		X"7E",X"03",X"FE",X"00",X"CA",X"BC",X"22",X"DD",X"7E",X"03",X"3C",X"DD",X"77",X"03",X"FE",X"05",
		X"C2",X"57",X"22",X"DD",X"46",X"01",X"DD",X"4E",X"02",X"CD",X"DE",X"00",X"E5",X"FD",X"E1",X"FD",
		X"36",X"00",X"8A",X"FD",X"36",X"01",X"8B",X"11",X"E0",X"FF",X"FD",X"19",X"FD",X"36",X"00",X"88",
		X"FD",X"36",X"01",X"89",X"C3",X"BC",X"22",X"FE",X"09",X"C2",X"80",X"22",X"DD",X"46",X"01",X"DD",
		X"4E",X"02",X"CD",X"DE",X"00",X"E5",X"FD",X"E1",X"FD",X"36",X"00",X"8E",X"FD",X"36",X"01",X"8F",
		X"11",X"E0",X"FF",X"FD",X"19",X"FD",X"36",X"00",X"8C",X"FD",X"36",X"01",X"8D",X"C3",X"BC",X"22",
		X"FE",X"0D",X"DA",X"BC",X"22",X"DD",X"46",X"01",X"DD",X"4E",X"02",X"CD",X"DE",X"00",X"E5",X"FD",
		X"E1",X"FD",X"36",X"00",X"00",X"FD",X"36",X"01",X"00",X"11",X"E0",X"FF",X"FD",X"19",X"FD",X"36",
		X"00",X"00",X"FD",X"36",X"01",X"00",X"11",X"00",X"04",X"19",X"36",X"0A",X"23",X"36",X"0A",X"11",
		X"E0",X"FF",X"19",X"36",X"0A",X"2B",X"36",X"0A",X"DD",X"36",X"03",X"00",X"CD",X"2D",X"60",X"11",
		X"05",X"00",X"DD",X"19",X"C3",X"10",X"22",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"C9",X"C5",
		X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",X"3A",X"A2",X"81",X"FE",X"00",X"CA",X"43",X"23",X"3A",X"A6",
		X"81",X"FE",X"01",X"CA",X"43",X"23",X"3E",X"01",X"32",X"A6",X"81",X"FD",X"7E",X"00",X"FE",X"FF",
		X"20",X"04",X"FD",X"21",X"80",X"84",X"FD",X"CB",X"00",X"76",X"28",X"07",X"11",X"05",X"00",X"FD",
		X"19",X"18",X"E8",X"FD",X"CB",X"00",X"FE",X"FD",X"46",X"01",X"FD",X"4E",X"02",X"CD",X"DE",X"00",
		X"E5",X"DD",X"E1",X"11",X"00",X"04",X"19",X"3A",X"A4",X"85",X"47",X"70",X"3A",X"A2",X"85",X"DD",
		X"77",X"00",X"23",X"DD",X"23",X"70",X"3A",X"A3",X"85",X"DD",X"77",X"00",X"11",X"DF",X"FF",X"19",
		X"DD",X"19",X"70",X"3A",X"A0",X"85",X"DD",X"77",X"00",X"23",X"DD",X"23",X"70",X"3A",X"A1",X"85",
		X"DD",X"77",X"00",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"C9",X"3A",X"28",X"80",X"CB",X"57",
		X"C0",X"3A",X"8E",X"80",X"FE",X"00",X"C0",X"DD",X"21",X"53",X"84",X"3A",X"53",X"84",X"E6",X"03",
		X"FE",X"03",X"C2",X"46",X"24",X"DD",X"CB",X"00",X"56",X"20",X"2D",X"21",X"00",X"00",X"22",X"0C",
		X"85",X"22",X"0E",X"85",X"DD",X"CB",X"00",X"D6",X"DD",X"36",X"02",X"3D",X"DD",X"36",X"03",X"0E",
		X"DD",X"36",X"04",X"78",X"DD",X"36",X"05",X"78",X"DD",X"36",X"0C",X"01",X"DD",X"36",X"0D",X"00",
		X"3E",X"00",X"32",X"58",X"88",X"CD",X"A9",X"24",X"CD",X"47",X"24",X"FE",X"00",X"C2",X"01",X"24",
		X"DD",X"46",X"04",X"DD",X"4E",X"05",X"DD",X"36",X"01",X"00",X"FD",X"E5",X"FD",X"21",X"08",X"85",
		X"CD",X"F2",X"5F",X"FD",X"E1",X"FE",X"00",X"CA",X"DB",X"23",X"4F",X"E6",X"0C",X"28",X"09",X"2A",
		X"5D",X"84",X"CD",X"F3",X"1F",X"22",X"5D",X"84",X"3E",X"1C",X"CD",X"FC",X"00",X"79",X"E6",X"03",
		X"28",X"09",X"2A",X"5B",X"84",X"CD",X"F3",X"1F",X"22",X"5B",X"84",X"3A",X"53",X"84",X"E6",X"C0",
		X"FE",X"C0",X"20",X"1A",X"DD",X"CB",X"00",X"BE",X"DD",X"CB",X"00",X"B6",X"3A",X"5F",X"84",X"3C",
		X"FE",X"07",X"28",X"04",X"38",X"02",X"3E",X"01",X"32",X"5F",X"84",X"CD",X"A9",X"24",X"C3",X"38",
		X"24",X"3E",X"1A",X"CD",X"FC",X"00",X"3A",X"28",X"80",X"CB",X"FF",X"32",X"28",X"80",X"21",X"2C",
		X"01",X"22",X"36",X"80",X"21",X"00",X"00",X"22",X"53",X"84",X"22",X"55",X"84",X"CD",X"10",X"25",
		X"DD",X"66",X"0C",X"DD",X"36",X"0C",X"00",X"7C",X"21",X"00",X"00",X"FD",X"21",X"08",X"85",X"CD",
		X"F3",X"00",X"DD",X"36",X"0D",X"1E",X"18",X"03",X"CD",X"F3",X"2C",X"DD",X"21",X"54",X"84",X"FD",
		X"21",X"08",X"85",X"CD",X"24",X"2D",X"C9",X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",X"3A",X"8D",
		X"80",X"FE",X"00",X"20",X"4A",X"3A",X"28",X"80",X"CB",X"57",X"20",X"43",X"11",X"00",X"00",X"3A",
		X"02",X"85",X"5F",X"21",X"08",X"00",X"19",X"EB",X"01",X"00",X"00",X"DD",X"4E",X"04",X"21",X"08",
		X"00",X"09",X"ED",X"52",X"CD",X"F0",X"1F",X"7D",X"FE",X"0A",X"D2",X"9F",X"24",X"11",X"00",X"00",
		X"3A",X"03",X"85",X"5F",X"21",X"0A",X"00",X"19",X"EB",X"01",X"00",X"00",X"DD",X"4E",X"05",X"21",
		X"08",X"00",X"09",X"ED",X"52",X"CD",X"F0",X"1F",X"7D",X"FE",X"0A",X"28",X"04",X"38",X"02",X"3E",
		X"00",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"C9",X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",
		X"FD",X"21",X"00",X"88",X"11",X"0A",X"00",X"FD",X"7E",X"00",X"E6",X"7F",X"FE",X"0E",X"28",X"04",
		X"FD",X"19",X"18",X"F3",X"21",X"48",X"0D",X"3A",X"5F",X"84",X"FE",X"00",X"28",X"0F",X"3D",X"21",
		X"9E",X"0D",X"11",X"12",X"00",X"FE",X"00",X"28",X"04",X"19",X"3D",X"18",X"F8",X"FD",X"75",X"01",
		X"FD",X"74",X"02",X"E5",X"DD",X"E1",X"06",X"07",X"FD",X"21",X"E2",X"8C",X"78",X"FE",X"00",X"28",
		X"17",X"DD",X"7E",X"00",X"FD",X"77",X"00",X"DD",X"7E",X"01",X"FD",X"77",X"01",X"DD",X"23",X"DD",
		X"23",X"FD",X"23",X"FD",X"23",X"05",X"18",X"E4",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"C9",
		X"C5",X"FD",X"E5",X"3A",X"5F",X"84",X"3D",X"FD",X"21",X"7E",X"2F",X"FE",X"00",X"28",X"07",X"FD",
		X"23",X"FD",X"23",X"3D",X"18",X"F5",X"FD",X"46",X"01",X"FD",X"4E",X"00",X"CD",X"E4",X"00",X"FD",
		X"E1",X"C1",X"C9",X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",X"DD",X"21",X"00",X"89",X"DD",X"CB",
		X"00",X"4E",X"20",X"06",X"CD",X"27",X"27",X"CD",X"00",X"28",X"DD",X"7E",X"11",X"FE",X"00",X"C2",
		X"95",X"26",X"DD",X"CB",X"00",X"7E",X"C2",X"E6",X"26",X"DD",X"CB",X"00",X"56",X"C2",X"9E",X"25",
		X"CD",X"C4",X"27",X"FE",X"00",X"C2",X"33",X"26",X"DD",X"36",X"03",X"0C",X"DD",X"36",X"0D",X"FF",
		X"DD",X"36",X"0E",X"03",X"DD",X"36",X"0F",X"00",X"DD",X"CB",X"00",X"D6",X"DD",X"36",X"07",X"00",
		X"DD",X"36",X"0A",X"00",X"DD",X"36",X"0B",X"00",X"21",X"AA",X"00",X"22",X"08",X"89",X"3A",X"2B",
		X"80",X"CB",X"47",X"28",X"06",X"21",X"56",X"FF",X"22",X"08",X"89",X"C3",X"1F",X"27",X"DD",X"46",
		X"04",X"DD",X"4E",X"05",X"DD",X"36",X"01",X"01",X"FD",X"E5",X"FD",X"21",X"10",X"85",X"CD",X"F2",
		X"5F",X"FD",X"E1",X"47",X"DD",X"4E",X"10",X"DD",X"36",X"10",X"00",X"E6",X"03",X"FE",X"00",X"28",
		X"01",X"0C",X"78",X"2A",X"0A",X"89",X"11",X"0A",X"00",X"19",X"22",X"0A",X"89",X"CB",X"57",X"CA",
		X"2B",X"26",X"ED",X"5B",X"0A",X"89",X"21",X"00",X"00",X"DD",X"71",X"10",X"22",X"0A",X"89",X"7B",
		X"FE",X"46",X"38",X"11",X"3E",X"1D",X"CD",X"FC",X"00",X"DD",X"36",X"0D",X"10",X"DD",X"36",X"0E",
		X"01",X"DD",X"36",X"0F",X"00",X"3A",X"0D",X"89",X"FE",X"FF",X"28",X"0C",X"FE",X"00",X"20",X"08",
		X"DD",X"36",X"0D",X"FF",X"DD",X"36",X"0E",X"03",X"78",X"E6",X"03",X"FE",X"00",X"28",X"24",X"3E",
		X"1D",X"CD",X"FC",X"00",X"2A",X"08",X"89",X"CD",X"F3",X"1F",X"22",X"08",X"89",X"DD",X"36",X"0D",
		X"10",X"DD",X"36",X"0E",X"01",X"DD",X"36",X"0F",X"00",X"18",X"08",X"DD",X"36",X"0D",X"FF",X"DD",
		X"36",X"0E",X"03",X"3A",X"10",X"89",X"FE",X"03",X"D2",X"C9",X"26",X"DD",X"46",X"04",X"DD",X"4E",
		X"05",X"CD",X"47",X"24",X"FE",X"00",X"CA",X"19",X"27",X"3A",X"0C",X"89",X"FE",X"02",X"20",X"05",
		X"3E",X"01",X"32",X"88",X"80",X"3A",X"0C",X"89",X"FE",X"03",X"3E",X"1E",X"20",X"0C",X"3E",X"01",
		X"CD",X"FC",X"00",X"3E",X"01",X"32",X"8E",X"80",X"3E",X"28",X"CD",X"FC",X"00",X"DD",X"36",X"11",
		X"10",X"DD",X"36",X"02",X"AD",X"DD",X"36",X"03",X"2B",X"3A",X"04",X"89",X"D6",X"08",X"32",X"04",
		X"89",X"3A",X"05",X"89",X"D6",X"08",X"32",X"05",X"89",X"21",X"00",X"00",X"22",X"08",X"89",X"22",
		X"0A",X"89",X"C3",X"1C",X"27",X"DD",X"35",X"11",X"DD",X"7E",X"11",X"FE",X"00",X"20",X"7D",X"3A",
		X"04",X"89",X"C6",X"08",X"32",X"04",X"89",X"3A",X"05",X"89",X"C6",X"08",X"32",X"05",X"89",X"DD",
		X"36",X"13",X"1E",X"3A",X"0C",X"89",X"3D",X"FD",X"21",X"10",X"85",X"21",X"01",X"00",X"CD",X"F3",
		X"00",X"CD",X"89",X"28",X"CD",X"FC",X"28",X"18",X"53",X"DD",X"CB",X"00",X"FE",X"DD",X"36",X"12",
		X"05",X"DD",X"36",X"0D",X"05",X"DD",X"36",X"0E",X"05",X"DD",X"36",X"0F",X"00",X"21",X"00",X"00",
		X"22",X"08",X"89",X"22",X"0A",X"89",X"DD",X"46",X"04",X"DD",X"4E",X"05",X"CD",X"47",X"24",X"FE",
		X"00",X"C2",X"49",X"26",X"CD",X"C4",X"27",X"FE",X"00",X"20",X"21",X"3A",X"12",X"89",X"FE",X"10",
		X"30",X"12",X"DD",X"34",X"12",X"3A",X"12",X"89",X"32",X"0D",X"89",X"32",X"0E",X"89",X"DD",X"36",
		X"0F",X"00",X"18",X"08",X"CD",X"A7",X"28",X"18",X"03",X"CD",X"C4",X"27",X"CD",X"3C",X"28",X"FD",
		X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"C9",X"E5",X"21",X"00",X"00",X"22",X"14",X"85",X"22",X"16",
		X"85",X"DD",X"CB",X"00",X"C6",X"DD",X"CB",X"00",X"CE",X"DD",X"36",X"03",X"1C",X"21",X"00",X"00",
		X"22",X"06",X"89",X"22",X"0A",X"89",X"21",X"80",X"FF",X"22",X"0A",X"89",X"DD",X"36",X"0D",X"20",
		X"DD",X"36",X"0E",X"01",X"DD",X"36",X"0F",X"00",X"DD",X"36",X"10",X"00",X"DD",X"36",X"11",X"00",
		X"DD",X"36",X"12",X"00",X"DD",X"36",X"13",X"00",X"CD",X"C9",X"00",X"3A",X"25",X"80",X"FE",X"AA",
		X"20",X"1F",X"3A",X"70",X"80",X"FE",X"00",X"28",X"18",X"3A",X"14",X"80",X"CB",X"7F",X"28",X"07",
		X"3A",X"24",X"80",X"CB",X"67",X"28",X"0A",X"DD",X"36",X"02",X"14",X"DD",X"36",X"0C",X"03",X"18",
		X"2E",X"3A",X"14",X"80",X"CB",X"7F",X"28",X"09",X"3A",X"B3",X"81",X"FE",X"3C",X"38",X"18",X"18",
		X"07",X"3A",X"B3",X"81",X"FE",X"28",X"38",X"0F",X"3E",X"00",X"32",X"B3",X"81",X"DD",X"36",X"02",
		X"10",X"DD",X"36",X"0C",X"02",X"18",X"08",X"DD",X"36",X"02",X"0C",X"DD",X"36",X"0C",X"01",X"CD",
		X"F0",X"3F",X"E1",X"C9",X"E5",X"3A",X"0D",X"89",X"FE",X"FF",X"28",X"08",X"FE",X"00",X"CA",X"FE",
		X"27",X"DD",X"35",X"0D",X"DD",X"34",X"0F",X"3A",X"0E",X"89",X"DD",X"BE",X"0F",X"28",X"03",X"D2",
		X"FC",X"27",X"3A",X"02",X"89",X"E6",X"03",X"FE",X"03",X"20",X"0A",X"DD",X"CB",X"02",X"86",X"DD",
		X"CB",X"02",X"8E",X"18",X"03",X"DD",X"34",X"02",X"DD",X"36",X"0F",X"00",X"3E",X"01",X"E1",X"C9",
		X"D5",X"E5",X"FD",X"E5",X"FD",X"21",X"00",X"88",X"11",X"0A",X"00",X"FD",X"7E",X"00",X"E6",X"7F",
		X"FE",X"0C",X"28",X"04",X"FD",X"19",X"18",X"F3",X"21",X"C4",X"0E",X"3A",X"0C",X"89",X"FE",X"00",
		X"28",X"0F",X"3D",X"21",X"D4",X"0E",X"11",X"12",X"00",X"FE",X"00",X"28",X"04",X"19",X"3D",X"18",
		X"F8",X"FD",X"75",X"01",X"FD",X"74",X"02",X"FD",X"E1",X"E1",X"D1",X"C9",X"D5",X"E5",X"3A",X"8D",
		X"80",X"FE",X"00",X"20",X"29",X"2A",X"0A",X"89",X"7C",X"B5",X"20",X"11",X"DD",X"66",X"04",X"DD",
		X"6E",X"06",X"ED",X"5B",X"08",X"89",X"19",X"DD",X"74",X"04",X"DD",X"75",X"06",X"DD",X"66",X"05",
		X"DD",X"6E",X"07",X"ED",X"5B",X"0A",X"89",X"19",X"DD",X"74",X"05",X"DD",X"75",X"07",X"3A",X"02",
		X"89",X"32",X"10",X"85",X"3A",X"03",X"89",X"32",X"11",X"85",X"3A",X"04",X"89",X"32",X"12",X"85",
		X"3A",X"05",X"89",X"32",X"13",X"85",X"E1",X"D1",X"C9",X"CD",X"C1",X"28",X"3A",X"0C",X"89",X"FE",
		X"01",X"20",X"0B",X"3A",X"AC",X"81",X"FE",X"04",X"30",X"04",X"3C",X"32",X"AC",X"81",X"3E",X"00",
		X"32",X"00",X"89",X"32",X"10",X"89",X"C9",X"E5",X"3E",X"00",X"32",X"00",X"89",X"32",X"10",X"89",
		X"21",X"00",X"00",X"22",X"02",X"89",X"22",X"06",X"89",X"22",X"08",X"89",X"22",X"0A",X"89",X"E1",
		X"C9",X"C5",X"FD",X"E5",X"3A",X"0C",X"89",X"3D",X"FD",X"21",X"8C",X"2F",X"FE",X"00",X"28",X"07",
		X"FD",X"23",X"FD",X"23",X"3D",X"18",X"F5",X"FD",X"46",X"01",X"FD",X"4E",X"00",X"CD",X"E4",X"00",
		X"FD",X"E1",X"C1",X"C9",X"C5",X"D5",X"E5",X"21",X"EA",X"2D",X"11",X"14",X"89",X"01",X"68",X"00",
		X"ED",X"B0",X"CD",X"CF",X"00",X"CA",X"2D",X"10",X"E1",X"D1",X"C1",X"C9",X"CD",X"10",X"29",X"CD",
		X"CF",X"00",X"CE",X"2D",X"02",X"C9",X"CD",X"50",X"29",X"CD",X"CF",X"00",X"D2",X"2D",X"0C",X"C9",
		X"D5",X"E5",X"FD",X"E5",X"FD",X"21",X"52",X"2E",X"3A",X"AC",X"81",X"11",X"08",X"00",X"FE",X"00",
		X"28",X"05",X"FD",X"19",X"3D",X"18",X"F7",X"FD",X"66",X"01",X"FD",X"6E",X"00",X"22",X"26",X"89",
		X"FD",X"66",X"03",X"FD",X"6E",X"02",X"22",X"28",X"89",X"FD",X"66",X"05",X"FD",X"6E",X"04",X"22",
		X"2E",X"89",X"FD",X"66",X"07",X"FD",X"6E",X"06",X"22",X"30",X"89",X"FD",X"E1",X"E1",X"D1",X"C9",
		X"D5",X"E5",X"FD",X"E5",X"21",X"24",X"24",X"22",X"36",X"89",X"22",X"3C",X"89",X"22",X"42",X"89",
		X"22",X"48",X"89",X"22",X"4E",X"89",X"22",X"54",X"89",X"22",X"5A",X"89",X"22",X"60",X"89",X"22",
		X"66",X"89",X"22",X"6C",X"89",X"22",X"72",X"89",X"22",X"78",X"89",X"FD",X"21",X"7A",X"2E",X"3A",
		X"A7",X"81",X"CB",X"3F",X"11",X"04",X"00",X"FE",X"00",X"28",X"0A",X"FD",X"19",X"3D",X"FE",X"00",
		X"28",X"03",X"FD",X"19",X"3D",X"FD",X"66",X"01",X"FD",X"6E",X"00",X"22",X"36",X"89",X"22",X"3C",
		X"89",X"FD",X"66",X"03",X"FD",X"6E",X"02",X"22",X"42",X"89",X"22",X"48",X"89",X"FE",X"00",X"CA",
		X"18",X"2A",X"FD",X"21",X"86",X"2E",X"3D",X"FE",X"00",X"28",X"11",X"FD",X"19",X"3D",X"FE",X"00",
		X"28",X"0A",X"FD",X"19",X"3D",X"FE",X"00",X"28",X"03",X"FD",X"19",X"3D",X"FD",X"66",X"01",X"FD",
		X"6E",X"00",X"22",X"4E",X"89",X"22",X"54",X"89",X"FD",X"66",X"03",X"FD",X"6E",X"02",X"22",X"5A",
		X"89",X"22",X"60",X"89",X"FE",X"00",X"CA",X"18",X"2A",X"FD",X"21",X"96",X"2E",X"3D",X"28",X"10",
		X"FD",X"19",X"3D",X"FE",X"00",X"28",X"09",X"FD",X"19",X"3D",X"FE",X"00",X"28",X"02",X"FD",X"19",
		X"FD",X"66",X"01",X"FD",X"6E",X"00",X"22",X"66",X"89",X"22",X"6C",X"89",X"FD",X"66",X"03",X"FD",
		X"6E",X"02",X"22",X"72",X"89",X"22",X"78",X"89",X"FD",X"E1",X"E1",X"D1",X"C9",X"DD",X"7E",X"10",
		X"FE",X"00",X"28",X"06",X"DD",X"35",X"10",X"C3",X"A9",X"2A",X"2A",X"5C",X"82",X"B7",X"CB",X"2C",
		X"CB",X"1D",X"DD",X"CB",X"09",X"7E",X"28",X"03",X"CD",X"F3",X"1F",X"DD",X"74",X"09",X"DD",X"75",
		X"08",X"2A",X"5C",X"82",X"DD",X"CB",X"0B",X"7E",X"28",X"03",X"CD",X"F3",X"1F",X"DD",X"74",X"0B",
		X"DD",X"75",X"0A",X"DD",X"46",X"04",X"DD",X"4E",X"05",X"CD",X"F2",X"5F",X"FE",X"00",X"CA",X"94",
		X"2A",X"DD",X"36",X"10",X"01",X"4F",X"E6",X"0C",X"FE",X"00",X"28",X"0F",X"DD",X"66",X"0B",X"DD",
		X"6E",X"0A",X"CD",X"F3",X"1F",X"DD",X"74",X"0B",X"DD",X"75",X"0A",X"79",X"E6",X"03",X"FE",X"00",
		X"28",X"0F",X"DD",X"66",X"09",X"DD",X"6E",X"08",X"CD",X"F3",X"1F",X"DD",X"74",X"09",X"DD",X"75",
		X"08",X"C3",X"A9",X"2A",X"21",X"6E",X"2F",X"CD",X"10",X"2B",X"FD",X"74",X"00",X"FD",X"75",X"01",
		X"CD",X"AA",X"2A",X"CD",X"F3",X"2C",X"CD",X"89",X"2B",X"C9",X"C5",X"D5",X"E5",X"21",X"A6",X"2E",
		X"DD",X"7E",X"01",X"FE",X"02",X"28",X"18",X"21",X"CE",X"2E",X"FE",X"03",X"28",X"11",X"21",X"F6",
		X"2E",X"FE",X"04",X"28",X"0A",X"21",X"1E",X"2F",X"FE",X"05",X"28",X"03",X"21",X"46",X"2F",X"DD",
		X"CB",X"09",X"7E",X"20",X"04",X"11",X"14",X"00",X"19",X"DD",X"34",X"11",X"DD",X"4E",X"11",X"7E",
		X"B9",X"28",X"02",X"30",X"27",X"23",X"54",X"5D",X"DD",X"34",X"12",X"DD",X"34",X"12",X"06",X"00",
		X"DD",X"4E",X"12",X"09",X"7E",X"FE",X"FF",X"20",X"07",X"DD",X"36",X"12",X"00",X"62",X"6B",X"7E",
		X"DD",X"77",X"02",X"23",X"7E",X"DD",X"77",X"03",X"DD",X"36",X"11",X"00",X"E1",X"D1",X"C1",X"C9",
		X"D5",X"11",X"00",X"00",X"DD",X"7E",X"08",X"DD",X"B6",X"09",X"20",X"07",X"DD",X"CB",X"0B",X"7E",
		X"C2",X"83",X"2B",X"23",X"23",X"DD",X"CB",X"09",X"7E",X"20",X"07",X"DD",X"CB",X"0B",X"7E",X"C2",
		X"83",X"2B",X"23",X"23",X"DD",X"7E",X"0A",X"DD",X"B6",X"0B",X"20",X"07",X"DD",X"CB",X"09",X"7E",
		X"CA",X"83",X"2B",X"23",X"23",X"DD",X"CB",X"09",X"7E",X"20",X"07",X"DD",X"CB",X"0B",X"7E",X"CA",
		X"83",X"2B",X"23",X"23",X"DD",X"7E",X"08",X"DD",X"B6",X"09",X"20",X"07",X"DD",X"CB",X"0B",X"7E",
		X"CA",X"83",X"2B",X"23",X"23",X"DD",X"CB",X"09",X"7E",X"28",X"06",X"DD",X"CB",X"0B",X"7E",X"20",
		X"12",X"23",X"23",X"DD",X"7E",X"0A",X"DD",X"B6",X"0B",X"20",X"06",X"DD",X"CB",X"09",X"7E",X"20",
		X"02",X"23",X"23",X"56",X"23",X"5E",X"EB",X"D1",X"C9",X"C5",X"DD",X"7E",X"04",X"FD",X"77",X"02",
		X"DD",X"7E",X"01",X"0E",X"04",X"CB",X"4F",X"28",X"02",X"0E",X"FC",X"DD",X"7E",X"05",X"81",X"FD",
		X"77",X"03",X"C1",X"C9",X"2A",X"60",X"82",X"DD",X"75",X"0C",X"DD",X"74",X"0D",X"DD",X"75",X"0E",
		X"DD",X"74",X"0F",X"DD",X"7E",X"01",X"FE",X"04",X"20",X"1C",X"DD",X"36",X"0C",X"00",X"DD",X"36",
		X"0D",X"00",X"2A",X"5C",X"82",X"DD",X"CB",X"09",X"7E",X"28",X"03",X"CD",X"F3",X"1F",X"DD",X"74",
		X"09",X"DD",X"75",X"08",X"18",X"19",X"3A",X"02",X"85",X"47",X"DD",X"7E",X"04",X"90",X"38",X"0F",
		X"DD",X"66",X"0D",X"DD",X"6E",X"0C",X"CD",X"F3",X"1F",X"DD",X"74",X"0D",X"DD",X"75",X"0C",X"DD",
		X"7E",X"01",X"FE",X"03",X"20",X"1C",X"DD",X"36",X"0E",X"00",X"DD",X"36",X"0F",X"00",X"2A",X"5C",
		X"82",X"DD",X"CB",X"0B",X"7E",X"28",X"03",X"CD",X"F3",X"1F",X"DD",X"74",X"0B",X"DD",X"75",X"0A",
		X"18",X"19",X"3A",X"03",X"85",X"47",X"DD",X"7E",X"05",X"90",X"38",X"0F",X"DD",X"66",X"0F",X"DD",
		X"6E",X"0E",X"CD",X"F3",X"1F",X"DD",X"74",X"0F",X"DD",X"75",X"0E",X"DD",X"46",X"04",X"DD",X"4E",
		X"05",X"CD",X"F2",X"5F",X"FE",X"00",X"CA",X"79",X"2C",X"DD",X"36",X"10",X"01",X"4F",X"E6",X"0C",
		X"FE",X"00",X"28",X"17",X"DD",X"66",X"0B",X"DD",X"6E",X"0A",X"CD",X"F3",X"1F",X"DD",X"74",X"0B",
		X"DD",X"75",X"0A",X"DD",X"36",X"0E",X"00",X"DD",X"36",X"0F",X"00",X"79",X"E6",X"03",X"FE",X"00",
		X"28",X"17",X"DD",X"66",X"09",X"DD",X"6E",X"08",X"CD",X"F3",X"1F",X"DD",X"74",X"09",X"DD",X"75",
		X"08",X"DD",X"36",X"0C",X"00",X"DD",X"36",X"0D",X"00",X"CD",X"92",X"2C",X"CD",X"F3",X"2C",X"21",
		X"6E",X"2F",X"CD",X"10",X"2B",X"FD",X"74",X"00",X"FD",X"75",X"01",X"CD",X"AA",X"2A",X"CD",X"89",
		X"2B",X"C9",X"C5",X"D5",X"E5",X"DD",X"7E",X"01",X"FE",X"04",X"28",X"26",X"DD",X"66",X"09",X"DD",
		X"6E",X"08",X"DD",X"56",X"0D",X"DD",X"5E",X"0C",X"19",X"44",X"4D",X"CD",X"F0",X"1F",X"ED",X"5B",
		X"5C",X"82",X"ED",X"52",X"7C",X"B5",X"28",X"04",X"CB",X"7C",X"28",X"06",X"DD",X"70",X"09",X"DD",
		X"71",X"08",X"DD",X"7E",X"01",X"FE",X"03",X"28",X"26",X"DD",X"66",X"0B",X"DD",X"6E",X"0A",X"DD",
		X"56",X"0F",X"DD",X"5E",X"0E",X"19",X"44",X"4D",X"CD",X"F0",X"1F",X"ED",X"5B",X"5C",X"82",X"ED",
		X"52",X"7C",X"B5",X"28",X"04",X"CB",X"7C",X"28",X"06",X"DD",X"70",X"0B",X"DD",X"71",X"0A",X"D1",
		X"E1",X"C1",X"C9",X"3A",X"8D",X"80",X"FE",X"00",X"C0",X"E5",X"D5",X"DD",X"66",X"04",X"DD",X"6E",
		X"06",X"DD",X"56",X"09",X"DD",X"5E",X"08",X"19",X"DD",X"74",X"04",X"DD",X"75",X"06",X"DD",X"66",
		X"05",X"DD",X"6E",X"07",X"DD",X"56",X"0B",X"DD",X"5E",X"0A",X"19",X"DD",X"74",X"05",X"DD",X"75",
		X"07",X"D1",X"E1",X"C9",X"DD",X"7E",X"01",X"FD",X"77",X"00",X"DD",X"7E",X"02",X"FD",X"77",X"01",
		X"DD",X"7E",X"03",X"FD",X"77",X"02",X"DD",X"7E",X"04",X"FD",X"77",X"03",X"C9",X"DD",X"46",X"04",
		X"DD",X"4E",X"05",X"CD",X"F2",X"5F",X"FE",X"00",X"CA",X"B4",X"2D",X"4F",X"16",X"00",X"DD",X"5E",
		X"04",X"3A",X"02",X"85",X"26",X"00",X"6F",X"B7",X"ED",X"52",X"3A",X"64",X"82",X"54",X"5D",X"FE",
		X"00",X"28",X"04",X"19",X"3D",X"18",X"F8",X"CB",X"7C",X"28",X"04",X"CB",X"49",X"20",X"08",X"CB",
		X"7C",X"20",X"07",X"CB",X"41",X"28",X"03",X"CD",X"F3",X"1F",X"DD",X"75",X"08",X"DD",X"74",X"09",
		X"16",X"00",X"DD",X"5E",X"05",X"3A",X"03",X"85",X"26",X"00",X"6F",X"B7",X"ED",X"52",X"3A",X"64",
		X"82",X"54",X"5D",X"FE",X"00",X"28",X"04",X"19",X"3D",X"18",X"F8",X"CB",X"7C",X"28",X"04",X"CB",
		X"59",X"20",X"08",X"CB",X"7C",X"20",X"07",X"CB",X"51",X"28",X"03",X"CD",X"F3",X"1F",X"DD",X"75",
		X"0A",X"DD",X"74",X"0B",X"CD",X"F3",X"2C",X"21",X"6E",X"2F",X"CD",X"10",X"2B",X"FD",X"74",X"00",
		X"FD",X"75",X"01",X"CD",X"AA",X"2A",X"CD",X"89",X"2B",X"C9",X"14",X"89",X"1C",X"89",X"24",X"89",
		X"2C",X"89",X"34",X"89",X"3A",X"89",X"40",X"89",X"46",X"89",X"4C",X"89",X"52",X"89",X"58",X"89",
		X"5E",X"89",X"64",X"89",X"6A",X"89",X"70",X"89",X"76",X"89",X"00",X"0E",X"C2",X"0E",X"C0",X"0E",
		X"FF",X"FF",X"01",X"0E",X"C3",X"0E",X"C1",X"0E",X"FF",X"FF",X"00",X"10",X"C6",X"0E",X"C4",X"0E",
		X"FF",X"FF",X"01",X"10",X"C7",X"0E",X"C5",X"0E",X"FF",X"FF",X"00",X"0D",X"E4",X"0E",X"FF",X"FF",
		X"01",X"0D",X"E4",X"0E",X"FF",X"FF",X"00",X"12",X"D8",X"0E",X"FF",X"FF",X"01",X"12",X"D8",X"0E",
		X"FF",X"FF",X"00",X"0C",X"00",X"0E",X"FF",X"FF",X"01",X"0C",X"00",X"0E",X"FF",X"FF",X"00",X"13",
		X"00",X"0E",X"FF",X"FF",X"01",X"13",X"00",X"0E",X"FF",X"FF",X"00",X"0B",X"00",X"0E",X"FF",X"FF",
		X"01",X"0B",X"00",X"0E",X"FF",X"FF",X"00",X"14",X"00",X"0E",X"FF",X"FF",X"01",X"14",X"00",X"0E",
		X"FF",X"FF",X"C6",X"0E",X"C4",X"0E",X"C7",X"0E",X"C5",X"0E",X"CA",X"0E",X"C8",X"0E",X"CB",X"0E",
		X"C9",X"0E",X"CE",X"0E",X"CC",X"0E",X"CF",X"0E",X"CD",X"0E",X"D2",X"0E",X"D0",X"0E",X"D3",X"0E",
		X"D1",X"0E",X"D6",X"0E",X"D4",X"0E",X"D7",X"0E",X"D5",X"0E",X"E4",X"0E",X"D8",X"0E",X"E5",X"0E",
		X"D9",X"0E",X"E6",X"0E",X"DA",X"0E",X"E8",X"0E",X"DC",X"0E",X"E9",X"0E",X"DD",X"0E",X"EA",X"0E",
		X"DE",X"0E",X"EB",X"0E",X"DF",X"0E",X"EC",X"0E",X"E0",X"0E",X"ED",X"0E",X"E1",X"0E",X"EE",X"0E",
		X"E2",X"0E",X"EF",X"0E",X"E3",X"0E",X"07",X"50",X"04",X"51",X"04",X"52",X"04",X"53",X"04",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"50",X"84",X"51",X"84",X"52",
		X"84",X"53",X"84",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"02",X"67",
		X"04",X"68",X"04",X"69",X"04",X"6A",X"04",X"6B",X"04",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"02",X"67",X"04",X"68",X"04",X"69",X"04",X"6A",X"04",X"6B",X"04",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"54",X"04",X"55",X"04",X"56",X"04",X"57",X"04",X"58",
		X"04",X"59",X"04",X"5A",X"04",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"5A",X"04",X"59",X"04",X"58",
		X"04",X"57",X"04",X"56",X"04",X"55",X"04",X"54",X"04",X"FF",X"FF",X"FF",X"FF",X"FF",X"06",X"38",
		X"04",X"39",X"04",X"3A",X"04",X"3B",X"04",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"06",X"38",X"84",X"39",X"84",X"3A",X"84",X"3B",X"84",X"FF",X"FF",X"39",X"04",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"06",X"60",X"04",X"61",X"04",X"62",X"04",X"63",X"04",X"64",
		X"04",X"65",X"04",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"06",X"65",X"04",X"64",X"04",X"63",
		X"04",X"62",X"04",X"61",X"04",X"60",X"04",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"02",X"00",X"03",X"00",X"05",X"00",X"08",X"00",X"12",X"00",X"20",X"00",X"10",X"00",X"30",
		X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C3",X"E4",X"28",X"C3",X"FC",X"28",X"C3",X"06",X"29",X"C3",X"05",X"22",X"C3",X"FF",X"FF",X"00",
		X"C3",X"1D",X"2A",X"C3",X"A4",X"2B",X"C3",X"3D",X"2D",X"C3",X"A9",X"24",X"00",X"00",X"00",X"00",
		X"3A",X"88",X"80",X"FE",X"03",X"CA",X"83",X"30",X"3A",X"8E",X"80",X"B7",X"C2",X"83",X"30",X"CD",
		X"8F",X"3C",X"3A",X"28",X"80",X"CB",X"7F",X"C2",X"3A",X"30",X"3A",X"8D",X"80",X"B7",X"C2",X"3A",
		X"30",X"CD",X"83",X"31",X"CD",X"1A",X"32",X"CD",X"5A",X"33",X"3E",X"01",X"CD",X"81",X"3D",X"C4",
		X"44",X"3D",X"3E",X"20",X"CD",X"81",X"3D",X"C4",X"C8",X"3C",X"DD",X"21",X"78",X"82",X"FD",X"21",
		X"18",X"85",X"11",X"19",X"00",X"06",X"09",X"0E",X"00",X"C5",X"D5",X"DD",X"7E",X"00",X"B7",X"CA",
		X"5E",X"30",X"1F",X"0C",X"D2",X"52",X"30",X"21",X"86",X"30",X"79",X"CD",X"EA",X"00",X"D1",X"C1",
		X"DD",X"19",X"D5",X"11",X"08",X"00",X"FD",X"19",X"D1",X"10",X"DE",X"CD",X"00",X"60",X"3A",X"8D",
		X"80",X"B7",X"CA",X"83",X"30",X"3A",X"28",X"80",X"CB",X"57",X"C2",X"83",X"30",X"3E",X"00",X"32",
		X"4B",X"82",X"C9",X"C3",X"C3",X"00",X"81",X"31",X"98",X"30",X"81",X"31",X"EF",X"30",X"81",X"31",
		X"81",X"31",X"35",X"31",X"81",X"31",X"81",X"31",X"DD",X"7E",X"01",X"21",X"CF",X"30",X"CD",X"EA",
		X"00",X"DD",X"7E",X"01",X"FE",X"0C",X"D2",X"CE",X"30",X"DD",X"7E",X"01",X"FE",X"01",X"CA",X"CE",
		X"30",X"DD",X"7E",X"01",X"FE",X"08",X"CA",X"CE",X"30",X"DD",X"7E",X"01",X"FE",X"07",X"CA",X"CE",
		X"30",X"3A",X"4A",X"82",X"B7",X"C2",X"CE",X"30",X"21",X"BB",X"3D",X"CD",X"07",X"36",X"C9",X"81",
		X"31",X"1C",X"32",X"73",X"32",X"81",X"31",X"10",X"33",X"81",X"31",X"81",X"31",X"1D",X"33",X"66",
		X"32",X"81",X"31",X"81",X"31",X"81",X"31",X"CE",X"39",X"1F",X"3A",X"C0",X"3A",X"81",X"31",X"00",
		X"DD",X"7E",X"01",X"21",X"15",X"31",X"CD",X"EA",X"00",X"DD",X"7E",X"01",X"FE",X"0C",X"D2",X"14",
		X"31",X"CD",X"CB",X"34",X"CD",X"32",X"3B",X"3A",X"4A",X"82",X"B7",X"C2",X"14",X"31",X"21",X"C3",
		X"3D",X"CD",X"07",X"36",X"C9",X"81",X"31",X"81",X"31",X"E2",X"33",X"63",X"34",X"81",X"31",X"81",
		X"31",X"81",X"31",X"81",X"31",X"81",X"31",X"81",X"31",X"81",X"31",X"81",X"31",X"CE",X"39",X"1F",
		X"3A",X"C0",X"3A",X"81",X"31",X"00",X"DD",X"7E",X"01",X"21",X"61",X"31",X"CD",X"EA",X"00",X"DD",
		X"7E",X"01",X"FE",X"0C",X"30",X"1A",X"3A",X"4A",X"82",X"B7",X"C2",X"60",X"31",X"DD",X"7E",X"13",
		X"B7",X"CA",X"5A",X"31",X"DD",X"35",X"13",X"C3",X"60",X"31",X"21",X"C7",X"3D",X"CD",X"07",X"36",
		X"C9",X"81",X"31",X"6B",X"35",X"F2",X"35",X"F9",X"35",X"F9",X"35",X"F9",X"35",X"00",X"36",X"81",
		X"31",X"81",X"31",X"81",X"31",X"81",X"31",X"81",X"31",X"CE",X"39",X"1F",X"3A",X"C0",X"3A",X"81",
		X"31",X"00",X"C9",X"21",X"D2",X"80",X"7E",X"23",X"BE",X"CA",X"19",X"32",X"2A",X"DA",X"80",X"2B",
		X"22",X"DA",X"80",X"7D",X"B4",X"C2",X"19",X"32",X"3A",X"D3",X"80",X"3C",X"32",X"D3",X"80",X"2A",
		X"D4",X"80",X"22",X"DA",X"80",X"DD",X"21",X"AA",X"82",X"06",X"07",X"CD",X"B7",X"38",X"B7",X"C2",
		X"19",X"32",X"21",X"CF",X"3D",X"CD",X"67",X"38",X"3A",X"2B",X"80",X"D6",X"78",X"38",X"09",X"DD",
		X"7E",X"04",X"FE",X"78",X"30",X"EC",X"18",X"07",X"DD",X"7E",X"04",X"FE",X"78",X"38",X"E3",X"DD",
		X"7E",X"04",X"C6",X"F8",X"DD",X"77",X"04",X"DD",X"7E",X"05",X"C6",X"F8",X"DD",X"77",X"05",X"DD",
		X"36",X"00",X"01",X"DD",X"36",X"01",X"01",X"DD",X"36",X"03",X"0F",X"DD",X"CB",X"03",X"EE",X"21",
		X"80",X"00",X"DD",X"75",X"08",X"DD",X"74",X"09",X"DD",X"36",X"0E",X"10",X"DD",X"36",X"0F",X"00",
		X"DD",X"36",X"14",X"01",X"2A",X"D6",X"80",X"DD",X"75",X"16",X"DD",X"74",X"17",X"3A",X"8D",X"80",
		X"B7",X"C2",X"19",X"32",X"3E",X"15",X"CD",X"FC",X"00",X"C9",X"00",X"C9",X"00",X"DD",X"35",X"14",
		X"C2",X"65",X"32",X"DD",X"36",X"14",X"06",X"21",X"73",X"3E",X"01",X"01",X"00",X"DD",X"7E",X"10",
		X"CD",X"F6",X"00",X"7E",X"FE",X"FF",X"CA",X"41",X"32",X"DD",X"77",X"02",X"DD",X"34",X"10",X"18",
		X"24",X"DD",X"36",X"02",X"04",X"DD",X"36",X"03",X"04",X"DD",X"36",X"10",X"00",X"DD",X"36",X"14",
		X"1E",X"DD",X"36",X"01",X"08",X"DD",X"7E",X"04",X"C6",X"08",X"DD",X"77",X"04",X"DD",X"7E",X"05",
		X"C6",X"08",X"DD",X"77",X"05",X"C9",X"DD",X"35",X"14",X"C2",X"6F",X"32",X"CD",X"AF",X"3B",X"CD",
		X"D6",X"32",X"C9",X"DD",X"6E",X"16",X"DD",X"66",X"17",X"7C",X"B5",X"CA",X"85",X"32",X"2B",X"DD",
		X"75",X"16",X"DD",X"74",X"17",X"CD",X"33",X"36",X"DD",X"7E",X"01",X"FE",X"02",X"C2",X"93",X"32",
		X"CD",X"09",X"60",X"CD",X"D6",X"32",X"CD",X"28",X"37",X"DD",X"7E",X"05",X"FE",X"D0",X"DA",X"D5",
		X"32",X"DD",X"36",X"01",X"07",X"DD",X"36",X"02",X"BC",X"DD",X"36",X"03",X"0F",X"DD",X"7E",X"04",
		X"C6",X"F8",X"DD",X"77",X"04",X"DD",X"7E",X"05",X"C6",X"F8",X"DD",X"77",X"05",X"DD",X"CB",X"03",
		X"EE",X"DD",X"36",X"10",X"00",X"DD",X"36",X"14",X"01",X"3A",X"8D",X"80",X"B7",X"C2",X"D5",X"32",
		X"3E",X"2D",X"CD",X"FC",X"00",X"C9",X"3A",X"4B",X"82",X"B7",X"C2",X"0F",X"33",X"3A",X"28",X"80",
		X"CB",X"7F",X"CA",X"0F",X"33",X"DD",X"E5",X"DD",X"E5",X"E1",X"11",X"E1",X"00",X"DD",X"19",X"DD",
		X"E5",X"D1",X"01",X"19",X"00",X"ED",X"B0",X"DD",X"E1",X"DD",X"36",X"01",X"0E",X"3E",X"22",X"DD",
		X"36",X"03",X"0B",X"DD",X"36",X"02",X"3F",X"FD",X"36",X"04",X"00",X"FD",X"36",X"05",X"00",X"C9",
		X"CD",X"03",X"60",X"CD",X"A9",X"36",X"CD",X"D6",X"32",X"CD",X"7A",X"37",X"C9",X"DD",X"35",X"14",
		X"C2",X"59",X"33",X"DD",X"36",X"14",X"06",X"21",X"73",X"3E",X"01",X"01",X"00",X"DD",X"7E",X"10",
		X"CD",X"F6",X"00",X"7E",X"FE",X"FF",X"CA",X"41",X"33",X"DD",X"77",X"02",X"DD",X"34",X"10",X"18",
		X"18",X"DD",X"36",X"00",X"20",X"DD",X"36",X"01",X"01",X"DD",X"7E",X"04",X"C6",X"08",X"DD",X"77",
		X"04",X"DD",X"7E",X"05",X"C6",X"08",X"DD",X"77",X"05",X"C9",X"21",X"C0",X"80",X"7E",X"23",X"BE",
		X"CA",X"E1",X"33",X"47",X"C5",X"DD",X"21",X"78",X"82",X"06",X"02",X"CD",X"B7",X"38",X"B7",X"C2",
		X"DE",X"33",X"DD",X"36",X"00",X"04",X"DD",X"36",X"01",X"02",X"DD",X"36",X"02",X"29",X"DD",X"36",
		X"03",X"84",X"DD",X"36",X"0D",X"01",X"DD",X"36",X"0E",X"00",X"DD",X"36",X"12",X"01",X"21",X"4F",
		X"3E",X"CD",X"70",X"38",X"3A",X"2B",X"80",X"D6",X"78",X"38",X"09",X"DD",X"7E",X"04",X"FE",X"78",
		X"30",X"EC",X"18",X"07",X"DD",X"7E",X"04",X"FE",X"78",X"38",X"E3",X"C1",X"C5",X"05",X"C2",X"C2",
		X"33",X"2A",X"4C",X"82",X"DD",X"5E",X"04",X"DD",X"56",X"05",X"B7",X"ED",X"52",X"CA",X"8E",X"33",
		X"18",X"09",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"22",X"4C",X"82",X"21",X"C4",X"80",X"CD",X"87",
		X"38",X"3A",X"C1",X"80",X"3C",X"32",X"C1",X"80",X"3A",X"C8",X"80",X"DD",X"77",X"16",X"C1",X"10",
		X"83",X"C9",X"DD",X"7E",X"18",X"B7",X"C2",X"59",X"34",X"DD",X"36",X"18",X"01",X"CD",X"1D",X"3C",
		X"B7",X"C2",X"59",X"34",X"DD",X"35",X"12",X"C2",X"59",X"34",X"DD",X"36",X"12",X"03",X"2A",X"C4",
		X"80",X"DD",X"75",X"08",X"DD",X"74",X"09",X"DD",X"75",X"0A",X"DD",X"74",X"0B",X"DD",X"7E",X"11",
		X"DD",X"77",X"10",X"3A",X"C2",X"80",X"32",X"6C",X"84",X"32",X"6D",X"84",X"32",X"6E",X"84",X"32",
		X"6F",X"84",X"21",X"6C",X"84",X"CD",X"9E",X"38",X"CD",X"06",X"60",X"B7",X"C3",X"34",X"34",X"CD",
		X"DC",X"38",X"18",X"0E",X"CD",X"1C",X"39",X"DD",X"70",X"11",X"7A",X"BB",X"D2",X"42",X"34",X"DD",
		X"71",X"11",X"CD",X"FC",X"3B",X"CD",X"84",X"39",X"B7",X"CA",X"4F",X"34",X"CD",X"0D",X"37",X"CD",
		X"06",X"3B",X"DD",X"7E",X"0F",X"B7",X"C2",X"5F",X"34",X"CD",X"09",X"60",X"CD",X"7A",X"3B",X"CD",
		X"D6",X"32",X"C9",X"DD",X"35",X"12",X"C2",X"C7",X"34",X"DD",X"7E",X"13",X"DD",X"77",X"12",X"DD",
		X"6E",X"14",X"DD",X"66",X"15",X"7E",X"FE",X"FF",X"CA",X"87",X"34",X"DD",X"77",X"02",X"23",X"DD",
		X"75",X"14",X"DD",X"74",X"15",X"18",X"40",X"23",X"3E",X"04",X"B6",X"DD",X"77",X"03",X"23",X"7E",
		X"DD",X"77",X"02",X"DD",X"36",X"0D",X"06",X"DD",X"36",X"0E",X"00",X"DD",X"36",X"12",X"03",X"DD",
		X"36",X"13",X"00",X"DD",X"36",X"14",X"00",X"DD",X"36",X"15",X"00",X"DD",X"36",X"01",X"02",X"DD",
		X"7E",X"0F",X"B7",X"CA",X"C7",X"34",X"DD",X"7E",X"17",X"DD",X"77",X"11",X"DD",X"36",X"17",X"00",
		X"CD",X"CB",X"34",X"DD",X"36",X"0F",X"00",X"CD",X"D6",X"32",X"C9",X"DD",X"7E",X"10",X"DD",X"BE",
		X"11",X"CA",X"F0",X"34",X"21",X"F1",X"34",X"01",X"08",X"00",X"DD",X"7E",X"10",X"CD",X"F6",X"00",
		X"DD",X"7E",X"11",X"CD",X"EA",X"00",X"DD",X"7E",X"11",X"DD",X"77",X"10",X"DD",X"36",X"01",X"03",
		X"C9",X"81",X"31",X"11",X"35",X"16",X"35",X"1B",X"35",X"20",X"35",X"81",X"31",X"25",X"35",X"2A",
		X"35",X"2F",X"35",X"34",X"35",X"81",X"31",X"39",X"35",X"3E",X"35",X"43",X"35",X"48",X"35",X"81",
		X"31",X"21",X"78",X"3E",X"18",X"37",X"21",X"7F",X"3E",X"18",X"32",X"21",X"86",X"3E",X"18",X"2D",
		X"21",X"8D",X"3E",X"18",X"28",X"21",X"94",X"3E",X"18",X"23",X"21",X"9B",X"3E",X"18",X"1E",X"21",
		X"A2",X"3E",X"18",X"19",X"21",X"A9",X"3E",X"18",X"14",X"21",X"B0",X"3E",X"18",X"0F",X"21",X"B7",
		X"3E",X"18",X"0A",X"21",X"BE",X"3E",X"18",X"05",X"21",X"C5",X"3E",X"18",X"00",X"DD",X"7E",X"03",
		X"E6",X"0F",X"B6",X"DD",X"77",X"03",X"23",X"7E",X"DD",X"77",X"02",X"23",X"DD",X"75",X"14",X"DD",
		X"74",X"15",X"DD",X"36",X"12",X"06",X"DD",X"36",X"13",X"06",X"C9",X"3A",X"B0",X"81",X"21",X"68",
		X"82",X"01",X"01",X"00",X"CD",X"F6",X"00",X"7E",X"E6",X"0F",X"F5",X"C6",X"02",X"DD",X"77",X"01",
		X"F1",X"21",X"D2",X"3E",X"01",X"02",X"00",X"CD",X"F6",X"00",X"7E",X"DD",X"77",X"03",X"23",X"7E",
		X"DD",X"77",X"02",X"DD",X"E5",X"06",X"13",X"DD",X"36",X"06",X"00",X"DD",X"23",X"10",X"F8",X"DD",
		X"E1",X"DD",X"36",X"13",X"1E",X"3E",X"01",X"32",X"77",X"82",X"3A",X"B0",X"81",X"3C",X"32",X"B0",
		X"81",X"3A",X"B0",X"81",X"FE",X"08",X"DA",X"BE",X"35",X"3E",X"00",X"32",X"B0",X"81",X"DD",X"36",
		X"0A",X"0A",X"DD",X"7E",X"01",X"FE",X"04",X"C2",X"D3",X"35",X"2A",X"5C",X"82",X"DD",X"75",X"0A",
		X"DD",X"74",X"0B",X"DD",X"7E",X"01",X"FE",X"02",X"C2",X"F1",X"35",X"FD",X"36",X"00",X"69",X"FD",
		X"36",X"01",X"45",X"DD",X"7E",X"04",X"FD",X"77",X"02",X"DD",X"7E",X"05",X"C6",X"FC",X"FD",X"77",
		X"03",X"C9",X"CD",X"F0",X"2F",X"CD",X"D6",X"32",X"C9",X"CD",X"F3",X"2F",X"CD",X"D6",X"32",X"C9",
		X"CD",X"F6",X"2F",X"CD",X"D6",X"32",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3A",
		X"8D",X"80",X"B7",X"C2",X"32",X"36",X"3A",X"28",X"80",X"CB",X"7F",X"C2",X"32",X"36",X"CD",X"9E",
		X"38",X"CD",X"06",X"60",X"B7",X"CA",X"32",X"36",X"21",X"28",X"80",X"CB",X"D6",X"3E",X"01",X"32",
		X"4B",X"82",X"C9",X"DD",X"46",X"04",X"DD",X"4E",X"05",X"78",X"E6",X"07",X"C2",X"A8",X"36",X"CD",
		X"00",X"38",X"B7",X"CA",X"A8",X"36",X"DD",X"7E",X"11",X"3C",X"E6",X"01",X"DD",X"77",X"11",X"AF",
		X"B1",X"C2",X"A8",X"36",X"DD",X"7E",X"16",X"DD",X"B6",X"17",X"C2",X"A8",X"36",X"2A",X"D6",X"80",
		X"DD",X"75",X"16",X"DD",X"74",X"17",X"DD",X"36",X"01",X"04",X"DD",X"36",X"08",X"00",X"DD",X"36",
		X"09",X"00",X"21",X"80",X"00",X"DD",X"75",X"0A",X"DD",X"74",X"0B",X"DD",X"36",X"10",X"00",X"DD",
		X"7E",X"11",X"B7",X"C2",X"90",X"36",X"DD",X"7E",X"04",X"D6",X"08",X"DD",X"77",X"04",X"18",X"08",
		X"DD",X"7E",X"04",X"C6",X"08",X"DD",X"77",X"04",X"DD",X"36",X"14",X"01",X"3A",X"8D",X"80",X"B7",
		X"C2",X"A8",X"36",X"3E",X"16",X"CD",X"FC",X"00",X"C9",X"DD",X"7E",X"04",X"C6",X"08",X"47",X"DD",
		X"7E",X"05",X"C6",X"14",X"4F",X"CD",X"DE",X"00",X"7E",X"CD",X"D6",X"5F",X"B7",X"CA",X"04",X"37",
		X"DD",X"36",X"0A",X"00",X"DD",X"36",X"0B",X"00",X"21",X"80",X"00",X"DD",X"75",X"08",X"DD",X"74",
		X"09",X"DD",X"36",X"0E",X"10",X"DD",X"36",X"0F",X"00",X"DD",X"36",X"10",X"00",X"DD",X"36",X"14",
		X"06",X"DD",X"36",X"15",X"00",X"DD",X"7E",X"05",X"E6",X"F8",X"C6",X"08",X"DD",X"77",X"05",X"DD",
		X"36",X"01",X"02",X"3A",X"8D",X"80",X"B7",X"C2",X"04",X"37",X"3E",X"17",X"CD",X"FC",X"00",X"3E",
		X"96",X"CD",X"FC",X"00",X"C9",X"11",X"F5",X"3E",X"CD",X"6B",X"39",X"B7",X"C9",X"21",X"57",X"3E",
		X"DD",X"7E",X"10",X"01",X"04",X"00",X"CD",X"F6",X"00",X"7E",X"DD",X"77",X"11",X"E5",X"CD",X"84",
		X"39",X"E1",X"23",X"B7",X"C2",X"19",X"37",X"C9",X"DD",X"7E",X"12",X"DD",X"BE",X"11",X"C2",X"4F",
		X"37",X"DD",X"35",X"14",X"C2",X"61",X"37",X"DD",X"36",X"14",X"06",X"CD",X"62",X"37",X"DD",X"34",
		X"10",X"DD",X"7E",X"10",X"FE",X"04",X"DA",X"61",X"37",X"DD",X"36",X"10",X"00",X"18",X"12",X"DD",
		X"7E",X"11",X"DD",X"77",X"12",X"DD",X"36",X"10",X"00",X"DD",X"36",X"14",X"06",X"DD",X"36",X"02",
		X"04",X"C9",X"DD",X"7E",X"11",X"B7",X"21",X"6F",X"3E",X"C2",X"6F",X"37",X"21",X"6B",X"3E",X"DD",
		X"5E",X"10",X"16",X"00",X"19",X"7E",X"DD",X"77",X"02",X"C9",X"DD",X"35",X"14",X"20",X"1A",X"DD",
		X"36",X"14",X"04",X"21",X"67",X"3E",X"DD",X"4E",X"10",X"06",X"00",X"09",X"7E",X"DD",X"77",X"02",
		X"DD",X"7E",X"10",X"3C",X"E6",X"03",X"DD",X"77",X"10",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"21",X"9F",X"3D",X"CD",X"30",X"38",X"CD",X"DE",X"00",X"7E",X"CD",X"D6",X"5F",X"B7",X"C2",X"26",
		X"38",X"21",X"97",X"3D",X"CD",X"30",X"38",X"CD",X"DE",X"00",X"7E",X"CD",X"D6",X"5F",X"B7",X"CA",
		X"2B",X"38",X"AF",X"C3",X"2F",X"38",X"0E",X"01",X"C3",X"2D",X"38",X"0E",X"00",X"3E",X"01",X"C9",
		X"DD",X"7E",X"11",X"E5",X"21",X"3A",X"38",X"C3",X"EA",X"00",X"42",X"38",X"47",X"38",X"4F",X"38",
		X"57",X"38",X"E1",X"CD",X"5B",X"38",X"C9",X"E1",X"CD",X"9B",X"38",X"CD",X"5B",X"38",X"C9",X"E1",
		X"CD",X"99",X"38",X"CD",X"5B",X"38",X"C9",X"E1",X"CD",X"97",X"38",X"DD",X"7E",X"04",X"86",X"47",
		X"23",X"DD",X"7E",X"05",X"86",X"4F",X"C9",X"01",X"08",X"00",X"3A",X"A1",X"81",X"CD",X"F6",X"00",
		X"CD",X"C9",X"00",X"3A",X"25",X"80",X"E6",X"03",X"87",X"16",X"00",X"5F",X"19",X"7E",X"DD",X"77",
		X"05",X"23",X"7E",X"DD",X"77",X"04",X"C9",X"5E",X"23",X"56",X"DD",X"73",X"08",X"DD",X"72",X"09",
		X"DD",X"73",X"0A",X"DD",X"72",X"0B",X"C9",X"23",X"23",X"23",X"23",X"23",X"23",X"C9",X"3A",X"2B",
		X"80",X"C6",X"08",X"47",X"3A",X"2C",X"80",X"C6",X"08",X"4F",X"DD",X"7E",X"04",X"C6",X"08",X"57",
		X"DD",X"7E",X"05",X"C6",X"08",X"5F",X"C9",X"11",X"19",X"00",X"AF",X"DD",X"B6",X"00",X"CA",X"CA",
		X"38",X"DD",X"19",X"10",X"F5",X"3E",X"01",X"C3",X"CC",X"38",X"3E",X"00",X"C9",X"DD",X"E5",X"06",
		X"19",X"DD",X"36",X"00",X"00",X"DD",X"23",X"10",X"F8",X"DD",X"E1",X"C9",X"CD",X"C9",X"00",X"3A",
		X"25",X"80",X"E6",X"03",X"21",X"EA",X"38",X"C3",X"EA",X"00",X"1B",X"39",X"F2",X"38",X"1B",X"39",
		X"08",X"39",X"DD",X"7E",X"11",X"FE",X"02",X"D2",X"01",X"39",X"DD",X"36",X"11",X"02",X"C3",X"1B",
		X"39",X"DD",X"36",X"11",X"00",X"C3",X"1B",X"39",X"DD",X"7E",X"11",X"FE",X"02",X"D2",X"17",X"39",
		X"DD",X"36",X"11",X"03",X"C3",X"1B",X"39",X"DD",X"36",X"11",X"01",X"C9",X"3A",X"2B",X"80",X"C6",
		X"08",X"6F",X"26",X"00",X"DD",X"7E",X"04",X"C6",X"08",X"5F",X"16",X"00",X"B7",X"ED",X"52",X"22",
		X"50",X"82",X"3A",X"2C",X"80",X"C6",X"08",X"6F",X"26",X"00",X"DD",X"7E",X"05",X"C6",X"08",X"5F",
		X"16",X"00",X"B7",X"ED",X"52",X"22",X"52",X"82",X"2A",X"50",X"82",X"7D",X"57",X"06",X"00",X"CB",
		X"7C",X"F2",X"59",X"39",X"ED",X"44",X"57",X"06",X"01",X"2A",X"52",X"82",X"7D",X"5F",X"0E",X"03",
		X"CB",X"7C",X"F2",X"6A",X"39",X"ED",X"44",X"5F",X"0E",X"02",X"C9",X"C5",X"E5",X"D5",X"E1",X"47",
		X"7E",X"23",X"FE",X"FF",X"CA",X"7F",X"39",X"B8",X"C2",X"70",X"39",X"AF",X"C3",X"81",X"39",X"3E",
		X"01",X"E1",X"C1",X"C9",X"21",X"AF",X"3D",X"CD",X"30",X"38",X"CD",X"DE",X"00",X"06",X"04",X"CD",
		X"A8",X"39",X"7E",X"C5",X"E5",X"CD",X"D6",X"5F",X"E1",X"C1",X"B7",X"C2",X"A5",X"39",X"10",X"EF",
		X"3E",X"00",X"C3",X"A7",X"39",X"3E",X"01",X"C9",X"E5",X"21",X"B0",X"39",X"78",X"C3",X"EA",X"00",
		X"CC",X"39",X"BA",X"39",X"BF",X"39",X"C7",X"39",X"CC",X"39",X"E1",X"23",X"C3",X"CD",X"39",X"E1",
		X"11",X"1F",X"00",X"19",X"C3",X"CD",X"39",X"E1",X"23",X"C3",X"CD",X"39",X"E1",X"C9",X"3A",X"49",
		X"82",X"FE",X"02",X"D2",X"DC",X"39",X"DD",X"35",X"14",X"C2",X"1E",X"3A",X"FD",X"36",X"04",X"00",
		X"FD",X"36",X"05",X"00",X"FD",X"36",X"06",X"00",X"FD",X"36",X"07",X"00",X"DD",X"7E",X"00",X"FE",
		X"01",X"C2",X"FE",X"39",X"3A",X"D3",X"80",X"3D",X"32",X"D3",X"80",X"C3",X"0D",X"3A",X"DD",X"7E",
		X"00",X"FE",X"20",X"CA",X"F4",X"39",X"3A",X"C1",X"80",X"3D",X"32",X"C1",X"80",X"CD",X"CD",X"38",
		X"3A",X"49",X"82",X"B7",X"CA",X"1E",X"3A",X"3A",X"49",X"82",X"3D",X"32",X"49",X"82",X"C9",X"DD",
		X"35",X"14",X"C2",X"81",X"3A",X"DD",X"7E",X"15",X"DD",X"77",X"14",X"21",X"DC",X"3E",X"16",X"00",
		X"DD",X"5E",X"10",X"19",X"7E",X"FE",X"FF",X"C2",X"7B",X"3A",X"DD",X"CB",X"03",X"AE",X"DD",X"7E",
		X"04",X"C6",X"08",X"DD",X"77",X"04",X"DD",X"7E",X"05",X"C6",X"08",X"DD",X"77",X"05",X"3A",X"47",
		X"82",X"21",X"03",X"00",X"CD",X"F3",X"00",X"CD",X"F1",X"3A",X"3A",X"47",X"82",X"FE",X"06",X"D2",
		X"69",X"3A",X"3A",X"47",X"82",X"3C",X"32",X"47",X"82",X"DD",X"36",X"14",X"1E",X"DD",X"36",X"01",
		X"0C",X"3A",X"49",X"82",X"3C",X"32",X"49",X"82",X"C3",X"81",X"3A",X"DD",X"77",X"02",X"DD",X"34",
		X"10",X"C9",X"21",X"CB",X"3D",X"CD",X"9E",X"38",X"CD",X"06",X"60",X"B7",X"CA",X"BF",X"3A",X"3E",
		X"2C",X"CD",X"FC",X"00",X"3A",X"B3",X"81",X"3C",X"32",X"B3",X"81",X"DD",X"36",X"10",X"00",X"DD",
		X"36",X"14",X"01",X"DD",X"36",X"15",X"04",X"DD",X"36",X"03",X"2D",X"DD",X"36",X"01",X"0D",X"DD",
		X"7E",X"04",X"C6",X"F8",X"DD",X"77",X"04",X"DD",X"7E",X"05",X"C6",X"F8",X"DD",X"77",X"05",X"C9",
		X"3A",X"28",X"80",X"CB",X"77",X"CA",X"CF",X"3A",X"DD",X"36",X"02",X"00",X"C3",X"D3",X"3A",X"DD",
		X"36",X"02",X"3F",X"3A",X"28",X"80",X"CB",X"7F",X"CA",X"E1",X"3A",X"CD",X"82",X"3A",X"C3",X"F0",
		X"3A",X"DD",X"E5",X"DD",X"E5",X"D1",X"E1",X"01",X"E1",X"00",X"09",X"01",X"19",X"00",X"ED",X"B0",
		X"C9",X"3A",X"47",X"82",X"01",X"02",X"00",X"21",X"01",X"3F",X"CD",X"F6",X"00",X"7E",X"4F",X"23",
		X"7E",X"47",X"CD",X"E4",X"00",X"C9",X"DD",X"35",X"16",X"C2",X"31",X"3B",X"3A",X"C8",X"80",X"DD",
		X"77",X"16",X"DD",X"7E",X"11",X"DD",X"77",X"17",X"CD",X"C9",X"00",X"3A",X"25",X"80",X"E6",X"03",
		X"DD",X"BE",X"10",X"28",X"F3",X"DD",X"BE",X"11",X"28",X"EE",X"DD",X"77",X"11",X"DD",X"36",X"0F",
		X"01",X"C9",X"3A",X"CC",X"80",X"3D",X"32",X"CC",X"80",X"C2",X"79",X"3B",X"3A",X"C6",X"80",X"32",
		X"CC",X"80",X"2A",X"C4",X"80",X"11",X"08",X"00",X"19",X"E5",X"11",X"00",X"02",X"B7",X"ED",X"52",
		X"E1",X"DA",X"55",X"3B",X"EB",X"22",X"C4",X"80",X"3A",X"4F",X"82",X"3D",X"32",X"4F",X"82",X"3A",
		X"C8",X"80",X"67",X"3A",X"C9",X"80",X"6F",X"7C",X"FE",X"18",X"D2",X"79",X"3B",X"11",X"20",X"00",
		X"19",X"7C",X"32",X"C8",X"80",X"7D",X"32",X"C9",X"80",X"C9",X"DD",X"35",X"0D",X"C2",X"AE",X"3B",
		X"DD",X"36",X"0D",X"06",X"21",X"CC",X"3E",X"DD",X"7E",X"11",X"FE",X"02",X"DA",X"92",X"3B",X"21",
		X"CF",X"3E",X"DD",X"7E",X"0E",X"01",X"01",X"00",X"CD",X"F6",X"00",X"7E",X"DD",X"77",X"02",X"DD",
		X"34",X"0E",X"DD",X"7E",X"0E",X"FE",X"03",X"DA",X"AE",X"3B",X"DD",X"36",X"0E",X"00",X"C9",X"DD",
		X"7E",X"04",X"C6",X"08",X"47",X"DD",X"7E",X"05",X"C6",X"14",X"4F",X"CD",X"DE",X"00",X"7E",X"CD",
		X"D6",X"5F",X"B7",X"C2",X"F3",X"3B",X"2A",X"D6",X"80",X"DD",X"75",X"16",X"DD",X"74",X"17",X"DD",
		X"36",X"08",X"00",X"DD",X"36",X"09",X"00",X"21",X"80",X"00",X"DD",X"75",X"0A",X"DD",X"74",X"0B",
		X"DD",X"36",X"10",X"00",X"DD",X"36",X"14",X"01",X"DD",X"36",X"01",X"04",X"3E",X"16",X"CD",X"FC",
		X"00",X"18",X"08",X"DD",X"36",X"14",X"06",X"DD",X"36",X"01",X"02",X"C9",X"DD",X"5E",X"10",X"16",
		X"00",X"21",X"11",X"3F",X"19",X"7E",X"DD",X"BE",X"11",X"C2",X"1C",X"3C",X"DD",X"7E",X"11",X"FE",
		X"02",X"D2",X"19",X"3C",X"DD",X"71",X"11",X"18",X"03",X"DD",X"70",X"11",X"C9",X"DD",X"7E",X"04",
		X"C6",X"08",X"E6",X"0F",X"11",X"88",X"3C",X"CD",X"6B",X"39",X"B7",X"20",X"54",X"DD",X"7E",X"05",
		X"C6",X"08",X"E6",X"0F",X"11",X"88",X"3C",X"CD",X"6B",X"39",X"B7",X"20",X"44",X"DD",X"7E",X"0C",
		X"B7",X"20",X"42",X"DD",X"36",X"0C",X"01",X"DD",X"7E",X"04",X"3C",X"E6",X"0F",X"FE",X"08",X"30",
		X"0D",X"3E",X"F0",X"DD",X"34",X"04",X"DD",X"A6",X"04",X"DD",X"77",X"04",X"18",X"04",X"3E",X"F8",
		X"18",X"F1",X"DD",X"7E",X"05",X"3C",X"E6",X"0F",X"FE",X"08",X"30",X"0D",X"3E",X"F0",X"DD",X"34",
		X"05",X"DD",X"A6",X"05",X"DD",X"77",X"05",X"18",X"04",X"3E",X"F8",X"18",X"F1",X"3E",X"00",X"18",
		X"06",X"DD",X"36",X"0C",X"00",X"3E",X"01",X"C9",X"0F",X"00",X"01",X"07",X"08",X"09",X"FF",X"3A",
		X"28",X"80",X"CB",X"7F",X"C2",X"C2",X"3C",X"DD",X"21",X"78",X"82",X"11",X"19",X"00",X"06",X"09",
		X"DD",X"7E",X"01",X"FE",X"0C",X"D2",X"C2",X"3C",X"DD",X"19",X"10",X"F4",X"3E",X"00",X"32",X"47",
		X"82",X"3A",X"4A",X"82",X"B7",X"CA",X"C7",X"3C",X"3A",X"4A",X"82",X"3D",X"32",X"4A",X"82",X"C3",
		X"C7",X"3C",X"3E",X"1E",X"32",X"4A",X"82",X"C9",X"2A",X"70",X"82",X"2B",X"22",X"70",X"82",X"7C",
		X"B5",X"C2",X"F3",X"3C",X"2A",X"5E",X"82",X"22",X"70",X"82",X"2A",X"5C",X"82",X"11",X"04",X"00",
		X"19",X"22",X"5C",X"82",X"01",X"40",X"04",X"B7",X"ED",X"42",X"DA",X"F3",X"3C",X"21",X"40",X"04",
		X"22",X"5C",X"82",X"2A",X"72",X"82",X"2B",X"22",X"72",X"82",X"7C",X"B5",X"C2",X"1C",X"3D",X"2A",
		X"62",X"82",X"22",X"72",X"82",X"2A",X"60",X"82",X"11",X"02",X"00",X"19",X"22",X"60",X"82",X"01",
		X"80",X"00",X"B7",X"ED",X"42",X"DA",X"1C",X"3D",X"ED",X"43",X"74",X"82",X"2A",X"74",X"82",X"2B",
		X"22",X"74",X"82",X"7C",X"B5",X"C2",X"43",X"3D",X"2A",X"66",X"82",X"22",X"74",X"82",X"3A",X"64",
		X"82",X"FE",X"0A",X"D2",X"3E",X"3D",X"C6",X"01",X"32",X"64",X"82",X"C3",X"43",X"3D",X"3E",X"0A",
		X"32",X"64",X"82",X"C9",X"2A",X"DC",X"80",X"2B",X"22",X"DC",X"80",X"7C",X"B5",X"C2",X"80",X"3D",
		X"2A",X"D8",X"80",X"22",X"DC",X"80",X"11",X"10",X"00",X"2A",X"D4",X"80",X"B7",X"ED",X"52",X"CA",
		X"65",X"3D",X"F2",X"68",X"3D",X"21",X"18",X"00",X"22",X"D4",X"80",X"2A",X"D6",X"80",X"11",X"10",
		X"00",X"B7",X"ED",X"52",X"CA",X"7A",X"3D",X"F2",X"7D",X"3D",X"21",X"01",X"00",X"22",X"D6",X"80",
		X"C9",X"21",X"78",X"82",X"11",X"19",X"00",X"06",X"09",X"BE",X"CA",X"93",X"3D",X"19",X"10",X"F9",
		X"AF",X"18",X"02",X"3E",X"01",X"B7",X"C9",X"0C",X"14",X"04",X"14",X"00",X"00",X"00",X"00",X"14",
		X"0C",X"FC",X"0C",X"00",X"00",X"00",X"00",X"10",X"14",X"00",X"14",X"10",X"FC",X"00",X"FC",X"1C",
		X"04",X"FC",X"04",X"0C",X"F4",X"0C",X"14",X"08",X"08",X"40",X"00",X"08",X"08",X"08",X"08",X"08",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"0C",X"0C",X"0C",X"0C",X"48",
		X"48",X"30",X"A8",X"48",X"48",X"30",X"A8",X"30",X"60",X"30",X"A0",X"30",X"60",X"30",X"A0",X"48",
		X"30",X"60",X"A8",X"48",X"30",X"60",X"A8",X"48",X"48",X"48",X"C0",X"48",X"48",X"48",X"C0",X"48",
		X"48",X"48",X"A8",X"48",X"48",X"48",X"A8",X"30",X"30",X"30",X"C0",X"30",X"30",X"30",X"C0",X"60",
		X"48",X"60",X"A8",X"60",X"48",X"60",X"A8",X"30",X"30",X"30",X"C0",X"30",X"30",X"30",X"C0",X"30",
		X"48",X"30",X"90",X"30",X"48",X"30",X"90",X"30",X"48",X"30",X"A8",X"30",X"48",X"30",X"A8",X"48",
		X"60",X"48",X"A8",X"48",X"60",X"48",X"A8",X"48",X"30",X"48",X"C0",X"48",X"30",X"48",X"C0",X"30",
		X"60",X"30",X"A8",X"30",X"60",X"30",X"A8",X"18",X"60",X"78",X"A8",X"18",X"60",X"78",X"A8",X"48",
		X"30",X"30",X"C0",X"48",X"30",X"30",X"C0",X"18",X"60",X"18",X"A8",X"18",X"60",X"18",X"A8",X"18",
		X"D8",X"18",X"18",X"D8",X"18",X"D8",X"D8",X"00",X"02",X"03",X"01",X"01",X"03",X"02",X"00",X"02",
		X"01",X"00",X"03",X"03",X"00",X"01",X"02",X"04",X"05",X"04",X"05",X"06",X"07",X"08",X"07",X"09",
		X"0A",X"0B",X"0A",X"BC",X"BD",X"BE",X"BF",X"FF",X"00",X"30",X"2D",X"2F",X"FF",X"00",X"29",X"00",
		X"30",X"2D",X"2E",X"FF",X"00",X"2C",X"00",X"30",X"2D",X"2E",X"FF",X"00",X"2C",X"80",X"30",X"2D",
		X"2F",X"FF",X"80",X"29",X"80",X"30",X"2D",X"2E",X"FF",X"00",X"2C",X"80",X"30",X"2D",X"2E",X"FF",
		X"00",X"2C",X"80",X"2F",X"29",X"2A",X"FF",X"80",X"2B",X"00",X"2F",X"29",X"2A",X"FF",X"00",X"2B",
		X"00",X"2C",X"2D",X"2E",X"FF",X"00",X"2D",X"80",X"2F",X"29",X"2A",X"FF",X"80",X"2B",X"00",X"2F",
		X"29",X"2A",X"FF",X"00",X"2B",X"00",X"2C",X"2D",X"2E",X"FF",X"00",X"2D",X"29",X"2A",X"2B",X"2C",
		X"2D",X"2E",X"04",X"50",X"04",X"34",X"04",X"54",X"04",X"38",X"04",X"60",X"A0",X"A1",X"A2",X"A3",
		X"FF",X"00",X"01",X"02",X"03",X"04",X"05",X"80",X"81",X"82",X"83",X"90",X"91",X"92",X"93",X"FF",
		X"80",X"81",X"82",X"83",X"FF",X"60",X"61",X"62",X"63",X"66",X"67",X"68",X"69",X"6A",X"A0",X"A2",
		X"FF",X"00",X"01",X"00",X"02",X"00",X"03",X"00",X"05",X"00",X"08",X"00",X"12",X"00",X"20",X"00",
		X"00",X"01",X"00",X"03",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3A",X"03",X"B0",X"FD",X"7E",X"03",X"C3",X"98",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3A",X"03",X"B0",X"FD",X"7E",X"03",X"C3",X"D8",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3A",X"03",X"B0",X"3A",X"00",X"B0",X"E6",X"10",X"C2",X"39",X"05",X"2B",X"7C",X"B5",X"C3",X"2A",
		X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"21",X"CF",X"3D",X"C3",X"67",X"38",X"C3",X"81",X"31",X"C3",X"81",X"31",X"C3",X"81",X"31",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
