library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity wacko_sp_bits_4 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of wacko_sp_bits_4 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"E0",X"00",X"90",X"EE",X"E0",X"00",X"90",X"9E",X"00",X"00",X"90",X"33",X"E0",X"00",
		X"99",X"99",X"90",X"00",X"39",X"9A",X"99",X"00",X"33",X"A9",X"AA",X"00",X"39",X"F9",X"FA",X"00",
		X"3B",X"FF",X"FF",X"00",X"9B",X"FF",X"F9",X"00",X"93",X"99",X"99",X"00",X"93",X"33",X"33",X"00",
		X"09",X"33",X"33",X"00",X"09",X"99",X"33",X"00",X"00",X"49",X"33",X"00",X"99",X"94",X"33",X"00",
		X"39",X"4B",X"33",X"00",X"39",X"B3",X"33",X"00",X"33",X"3B",X"33",X"00",X"93",X"3B",X"99",X"00",
		X"99",X"39",X"09",X"00",X"09",X"33",X"09",X"00",X"00",X"93",X"99",X"00",X"90",X"33",X"33",X"00",
		X"99",X"33",X"99",X"00",X"39",X"33",X"09",X"00",X"39",X"39",X"09",X"00",X"33",X"39",X"99",X"00",
		X"39",X"33",X"33",X"00",X"39",X"33",X"93",X"00",X"99",X"33",X"99",X"00",X"99",X"99",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"00",X"00",
		X"00",X"92",X"99",X"00",X"00",X"99",X"22",X"00",X"00",X"92",X"22",X"00",X"00",X"22",X"29",X"00",
		X"99",X"29",X"29",X"90",X"22",X"29",X"29",X"90",X"99",X"29",X"22",X"90",X"94",X"22",X"29",X"90",
		X"99",X"22",X"29",X"90",X"DD",X"29",X"22",X"90",X"22",X"99",X"92",X"90",X"99",X"59",X"92",X"90",
		X"99",X"59",X"92",X"00",X"99",X"99",X"92",X"00",X"99",X"99",X"92",X"00",X"99",X"99",X"92",X"00",
		X"95",X"99",X"22",X"00",X"99",X"22",X"22",X"00",X"DD",X"29",X"22",X"00",X"29",X"22",X"22",X"00",
		X"22",X"99",X"22",X"90",X"99",X"99",X"92",X"90",X"99",X"92",X"92",X"90",X"99",X"22",X"22",X"00",
		X"92",X"22",X"22",X"00",X"92",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",
		X"00",X"09",X"00",X"00",X"00",X"9D",X"00",X"00",X"00",X"9D",X"00",X"00",X"00",X"9D",X"99",X"00",
		X"00",X"99",X"22",X"00",X"00",X"92",X"22",X"00",X"00",X"22",X"29",X"00",X"99",X"29",X"29",X"90",
		X"22",X"29",X"29",X"90",X"99",X"29",X"22",X"90",X"99",X"22",X"29",X"90",X"99",X"22",X"29",X"90",
		X"DD",X"29",X"22",X"90",X"22",X"99",X"92",X"90",X"99",X"59",X"92",X"90",X"99",X"59",X"92",X"00",
		X"99",X"99",X"92",X"00",X"22",X"92",X"92",X"00",X"22",X"22",X"92",X"00",X"29",X"22",X"22",X"00",
		X"99",X"22",X"22",X"00",X"99",X"92",X"22",X"00",X"99",X"99",X"22",X"00",X"99",X"DD",X"22",X"90",
		X"29",X"22",X"92",X"90",X"29",X"22",X"92",X"90",X"99",X"22",X"22",X"00",X"92",X"22",X"22",X"00",
		X"92",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",
		X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"99",X"00",X"22",X"22",X"9A",X"00",
		X"99",X"22",X"99",X"00",X"9A",X"22",X"99",X"00",X"99",X"22",X"22",X"00",X"99",X"22",X"22",X"00",
		X"22",X"22",X"22",X"00",X"99",X"22",X"22",X"00",X"22",X"99",X"22",X"00",X"22",X"9D",X"22",X"00",
		X"99",X"9D",X"22",X"00",X"00",X"99",X"22",X"00",X"99",X"00",X"29",X"00",X"29",X"00",X"29",X"00",
		X"22",X"00",X"29",X"00",X"22",X"00",X"29",X"00",X"22",X"00",X"29",X"00",X"22",X"00",X"29",X"00",
		X"22",X"00",X"99",X"00",X"99",X"00",X"22",X"00",X"90",X"00",X"29",X"00",X"90",X"00",X"99",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"09",X"99",X"90",
		X"00",X"09",X"22",X"90",X"00",X"99",X"22",X"90",X"00",X"92",X"22",X"90",X"00",X"99",X"99",X"90",
		X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"99",X"22",X"92",X"00",
		X"9A",X"92",X"92",X"00",X"99",X"99",X"92",X"00",X"99",X"22",X"92",X"00",X"22",X"92",X"29",X"00",
		X"99",X"92",X"99",X"00",X"29",X"22",X"92",X"90",X"99",X"22",X"92",X"99",X"92",X"22",X"92",X"29",
		X"22",X"22",X"99",X"29",X"22",X"22",X"09",X"29",X"22",X"19",X"00",X"29",X"22",X"00",X"99",X"99",
		X"22",X"00",X"22",X"90",X"22",X"00",X"22",X"00",X"29",X"00",X"22",X"00",X"29",X"00",X"22",X"00",
		X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",
		X"92",X"00",X"92",X"00",X"99",X"00",X"99",X"90",X"99",X"00",X"09",X"99",X"99",X"00",X"09",X"29",
		X"22",X"00",X"00",X"29",X"22",X"00",X"00",X"29",X"22",X"00",X"00",X"99",X"99",X"00",X"00",X"00",
		X"00",X"00",X"90",X"90",X"00",X"00",X"99",X"90",X"00",X"09",X"BB",X"90",X"00",X"99",X"BB",X"90",
		X"00",X"99",X"BB",X"90",X"00",X"99",X"BB",X"00",X"99",X"BB",X"BB",X"00",X"9B",X"BB",X"BB",X"00",
		X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"9B",X"00",X"BB",X"99",X"99",X"00",X"BB",X"95",X"99",X"00",
		X"99",X"95",X"99",X"00",X"99",X"95",X"99",X"00",X"94",X"99",X"99",X"00",X"44",X"BB",X"99",X"00",
		X"4B",X"BB",X"BB",X"00",X"9B",X"BB",X"BB",X"00",X"BB",X"99",X"BB",X"00",X"99",X"9B",X"BB",X"00",
		X"00",X"9B",X"BB",X"00",X"00",X"9B",X"BB",X"00",X"00",X"9B",X"B9",X"00",X"00",X"99",X"99",X"00",
		X"00",X"77",X"9B",X"00",X"09",X"77",X"BB",X"00",X"99",X"77",X"BB",X"00",X"9B",X"99",X"BB",X"00",
		X"BB",X"11",X"BB",X"00",X"B9",X"77",X"BB",X"00",X"99",X"99",X"BB",X"00",X"97",X"11",X"BB",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"90",X"00",X"00",X"99",X"90",X"00",X"09",X"BB",X"90",
		X"00",X"99",X"BB",X"90",X"00",X"99",X"BB",X"90",X"00",X"99",X"BB",X"00",X"99",X"BB",X"BB",X"00",
		X"9B",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",
		X"BB",X"99",X"9B",X"00",X"99",X"95",X"99",X"00",X"99",X"95",X"99",X"00",X"99",X"99",X"99",X"00",
		X"44",X"99",X"99",X"00",X"B4",X"BB",X"99",X"00",X"9B",X"BB",X"BB",X"00",X"BB",X"99",X"BB",X"00",
		X"99",X"9B",X"BB",X"00",X"00",X"9B",X"BB",X"00",X"00",X"9B",X"BB",X"00",X"00",X"9B",X"99",X"00",
		X"00",X"99",X"9B",X"00",X"00",X"77",X"BB",X"00",X"09",X"77",X"BB",X"00",X"99",X"77",X"BB",X"00",
		X"9B",X"99",X"BB",X"00",X"BB",X"11",X"BB",X"00",X"B9",X"77",X"BB",X"00",X"99",X"99",X"BB",X"00",
		X"97",X"77",X"BB",X"09",X"99",X"99",X"BB",X"9B",X"11",X"11",X"BB",X"9B",X"77",X"77",X"BB",X"9B",
		X"77",X"77",X"BB",X"BB",X"99",X"77",X"BB",X"B9",X"11",X"17",X"BB",X"B9",X"77",X"79",X"BB",X"B9",
		X"77",X"99",X"BB",X"19",X"99",X"9B",X"BB",X"B9",X"11",X"B9",X"BB",X"B9",X"77",X"B9",X"B9",X"B9",
		X"77",X"B9",X"B9",X"B9",X"77",X"BB",X"B9",X"B9",X"99",X"9B",X"BB",X"99",X"91",X"9B",X"9B",X"90",
		X"99",X"99",X"9B",X"90",X"B9",X"79",X"99",X"00",X"B9",X"79",X"BB",X"00",X"BB",X"99",X"BB",X"00",
		X"99",X"00",X"99",X"00",X"BB",X"00",X"BB",X"99",X"BB",X"00",X"B9",X"B9",X"BB",X"00",X"B9",X"B9",
		X"99",X"00",X"B9",X"B9",X"BB",X"00",X"BB",X"B9",X"BB",X"00",X"BB",X"B9",X"BB",X"00",X"BB",X"99",
		X"BB",X"00",X"99",X"90",X"BB",X"00",X"00",X"90",X"B9",X"00",X"09",X"90",X"99",X"00",X"09",X"90",
		X"97",X"11",X"BB",X"00",X"97",X"77",X"BB",X"09",X"99",X"99",X"BB",X"9B",X"1B",X"B9",X"BB",X"BB",
		X"9B",X"BB",X"BB",X"BB",X"99",X"BB",X"BB",X"BB",X"99",X"BB",X"B9",X"B9",X"11",X"BB",X"99",X"B9",
		X"77",X"B9",X"B9",X"B9",X"77",X"99",X"99",X"B9",X"99",X"9B",X"90",X"B9",X"11",X"BB",X"90",X"B9",
		X"77",X"BB",X"00",X"B9",X"77",X"BB",X"00",X"B9",X"77",X"BB",X"90",X"B9",X"99",X"9B",X"99",X"99",
		X"91",X"9B",X"BB",X"90",X"99",X"99",X"BB",X"90",X"09",X"79",X"BB",X"00",X"09",X"79",X"BB",X"00",
		X"00",X"99",X"BB",X"00",X"00",X"B9",X"99",X"00",X"00",X"B9",X"90",X"00",X"00",X"B9",X"00",X"00",
		X"00",X"B9",X"00",X"00",X"99",X"B9",X"00",X"00",X"BB",X"99",X"00",X"00",X"BB",X"BB",X"00",X"00",
		X"99",X"BB",X"00",X"00",X"9B",X"BB",X"00",X"00",X"9B",X"BB",X"00",X"00",X"99",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"66",X"00",X"00",
		X"09",X"66",X"99",X"00",X"09",X"66",X"69",X"00",X"99",X"66",X"69",X"00",X"96",X"66",X"99",X"00",
		X"66",X"66",X"66",X"00",X"69",X"99",X"66",X"00",X"99",X"E9",X"66",X"00",X"9E",X"99",X"69",X"00",
		X"9E",X"E9",X"69",X"00",X"EE",X"E9",X"99",X"00",X"EE",X"E9",X"96",X"00",X"EE",X"EE",X"96",X"00",
		X"EE",X"EE",X"96",X"00",X"EE",X"CC",X"66",X"00",X"EE",X"C9",X"66",X"00",X"99",X"99",X"66",X"00",
		X"C9",X"99",X"66",X"00",X"CC",X"99",X"66",X"00",X"CC",X"99",X"66",X"00",X"CC",X"99",X"66",X"00",
		X"CC",X"99",X"66",X"00",X"99",X"99",X"66",X"00",X"99",X"9C",X"66",X"00",X"99",X"CC",X"66",X"00",
		X"99",X"C9",X"66",X"00",X"99",X"99",X"66",X"00",X"CC",X"DD",X"66",X"00",X"99",X"66",X"66",X"00",
		X"00",X"99",X"00",X"00",X"09",X"66",X"00",X"00",X"09",X"66",X"00",X"00",X"09",X"66",X"00",X"00",
		X"99",X"66",X"90",X"00",X"66",X"66",X"99",X"00",X"66",X"66",X"66",X"00",X"69",X"99",X"66",X"00",
		X"99",X"E9",X"66",X"00",X"9E",X"99",X"69",X"00",X"9E",X"E9",X"69",X"00",X"EE",X"E9",X"99",X"00",
		X"EE",X"E9",X"96",X"00",X"EE",X"EE",X"96",X"00",X"EE",X"EE",X"96",X"00",X"EE",X"CC",X"66",X"00",
		X"EE",X"C9",X"66",X"00",X"99",X"99",X"66",X"00",X"C9",X"99",X"66",X"00",X"CC",X"99",X"66",X"00",
		X"CC",X"99",X"66",X"00",X"CC",X"99",X"66",X"00",X"CC",X"9C",X"66",X"00",X"99",X"CC",X"66",X"00",
		X"99",X"CC",X"66",X"00",X"99",X"CC",X"66",X"00",X"99",X"C9",X"66",X"00",X"CC",X"99",X"66",X"00",
		X"99",X"DD",X"66",X"00",X"6D",X"66",X"66",X"00",X"66",X"66",X"66",X"00",X"66",X"66",X"66",X"00",
		X"66",X"66",X"66",X"00",X"66",X"66",X"66",X"00",X"66",X"66",X"66",X"90",X"66",X"66",X"66",X"90",
		X"66",X"66",X"96",X"90",X"66",X"66",X"96",X"90",X"99",X"66",X"66",X"90",X"95",X"66",X"66",X"90",
		X"95",X"99",X"66",X"90",X"95",X"DD",X"66",X"90",X"95",X"DD",X"66",X"90",X"95",X"DD",X"66",X"90",
		X"99",X"99",X"96",X"90",X"66",X"66",X"96",X"90",X"66",X"66",X"96",X"90",X"D6",X"66",X"96",X"90",
		X"9D",X"66",X"96",X"90",X"9D",X"66",X"96",X"90",X"96",X"69",X"96",X"90",X"96",X"99",X"96",X"90",
		X"66",X"99",X"96",X"90",X"66",X"9D",X"99",X"90",X"66",X"99",X"9C",X"90",X"66",X"09",X"99",X"90",
		X"66",X"09",X"99",X"00",X"69",X"09",X"99",X"00",X"69",X"09",X"99",X"90",X"99",X"99",X"99",X"99",
		X"90",X"99",X"09",X"C9",X"90",X"97",X"09",X"99",X"90",X"77",X"09",X"C9",X"90",X"99",X"09",X"99",
		X"66",X"66",X"66",X"00",X"66",X"66",X"66",X"00",X"66",X"66",X"96",X"00",X"66",X"66",X"96",X"00",
		X"99",X"66",X"66",X"00",X"95",X"66",X"66",X"00",X"95",X"99",X"66",X"00",X"95",X"DD",X"66",X"00",
		X"95",X"DD",X"66",X"00",X"95",X"DD",X"66",X"00",X"99",X"99",X"66",X"00",X"66",X"66",X"66",X"00",
		X"66",X"66",X"66",X"00",X"66",X"66",X"66",X"00",X"96",X"66",X"66",X"00",X"99",X"66",X"66",X"00",
		X"D9",X"66",X"66",X"00",X"99",X"66",X"66",X"00",X"C9",X"66",X"66",X"00",X"C9",X"66",X"99",X"00",
		X"C9",X"66",X"CC",X"00",X"C9",X"66",X"CC",X"00",X"99",X"66",X"CC",X"00",X"97",X"66",X"9C",X"00",
		X"77",X"99",X"9C",X"00",X"77",X"77",X"CC",X"00",X"79",X"77",X"CC",X"00",X"99",X"77",X"CC",X"00",
		X"77",X"99",X"CC",X"00",X"77",X"00",X"CC",X"00",X"99",X"00",X"C9",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9B",X"00",X"00",
		X"00",X"E9",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"9E",X"00",X"00",X"99",X"9E",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"9E",X"00",X"00",X"9E",X"99",X"00",X"09",X"EE",X"99",X"00",
		X"09",X"99",X"99",X"00",X"09",X"99",X"E9",X"00",X"99",X"99",X"9E",X"00",X"99",X"99",X"9B",X"00",
		X"E9",X"99",X"99",X"00",X"E9",X"99",X"E9",X"00",X"E9",X"9E",X"EE",X"00",X"9E",X"E9",X"E9",X"00",
		X"99",X"99",X"E9",X"00",X"99",X"9E",X"E9",X"00",X"EE",X"9E",X"E9",X"00",X"EE",X"EE",X"9B",X"00",
		X"99",X"E9",X"9E",X"00",X"9E",X"E9",X"9B",X"00",X"9E",X"99",X"9B",X"00",X"EE",X"EE",X"E9",X"00",
		X"00",X"99",X"00",X"00",X"00",X"9B",X"00",X"00",X"00",X"E9",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"9E",X"00",X"00",X"99",X"9E",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"9E",X"00",
		X"00",X"9E",X"99",X"00",X"09",X"EE",X"99",X"00",X"09",X"99",X"99",X"00",X"09",X"99",X"E9",X"00",
		X"99",X"99",X"9E",X"00",X"99",X"99",X"9B",X"00",X"E9",X"99",X"99",X"00",X"E9",X"99",X"99",X"00",
		X"E9",X"99",X"9E",X"00",X"9E",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"9E",X"99",X"00",
		X"EE",X"9E",X"E9",X"00",X"EE",X"EE",X"9B",X"00",X"99",X"E9",X"9E",X"00",X"9E",X"E9",X"9B",X"00",
		X"9E",X"99",X"9B",X"00",X"EE",X"E9",X"E9",X"00",X"EE",X"EE",X"E9",X"00",X"EE",X"EE",X"E9",X"00",
		X"9E",X"99",X"E9",X"00",X"9E",X"BE",X"E9",X"00",X"99",X"9B",X"E9",X"00",X"EE",X"9B",X"EE",X"00",
		X"E9",X"99",X"E4",X"00",X"99",X"E9",X"EE",X"00",X"99",X"E9",X"9E",X"00",X"E9",X"9E",X"9E",X"00",
		X"E9",X"99",X"9E",X"00",X"9E",X"E9",X"EE",X"00",X"99",X"99",X"E9",X"00",X"99",X"99",X"99",X"00",
		X"E9",X"9E",X"9E",X"00",X"E9",X"9E",X"99",X"00",X"99",X"99",X"E9",X"00",X"9E",X"9B",X"EE",X"00",
		X"9E",X"99",X"E9",X"00",X"99",X"09",X"E9",X"00",X"E9",X"09",X"99",X"00",X"E9",X"09",X"E9",X"00",
		X"99",X"00",X"99",X"00",X"E9",X"00",X"9B",X"00",X"E9",X"00",X"9B",X"00",X"9E",X"00",X"9B",X"00",
		X"9E",X"09",X"99",X"00",X"94",X"99",X"E9",X"00",X"99",X"9E",X"99",X"00",X"E9",X"99",X"EE",X"00",
		X"EE",X"E9",X"EE",X"00",X"99",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"9E",X"E9",X"00",X"9E",X"9E",X"E9",X"00",X"9E",X"99",X"E9",X"00",X"9E",X"BE",X"E9",X"00",
		X"99",X"9B",X"E9",X"00",X"EE",X"99",X"E9",X"00",X"E9",X"99",X"E9",X"00",X"99",X"99",X"99",X"00",
		X"99",X"EE",X"99",X"00",X"E9",X"9E",X"99",X"00",X"E9",X"99",X"9B",X"00",X"9E",X"E9",X"9E",X"00",
		X"99",X"99",X"B9",X"00",X"E9",X"99",X"99",X"00",X"E9",X"9E",X"9E",X"00",X"99",X"9E",X"9E",X"00",
		X"E9",X"99",X"99",X"00",X"EE",X"9E",X"99",X"00",X"EE",X"99",X"9E",X"00",X"E9",X"09",X"9E",X"00",
		X"99",X"00",X"99",X"00",X"E9",X"00",X"9E",X"00",X"E9",X"00",X"EE",X"00",X"E9",X"00",X"E9",X"90",
		X"B9",X"00",X"E9",X"90",X"99",X"00",X"99",X"99",X"BB",X"00",X"99",X"E9",X"9E",X"00",X"E9",X"E9",
		X"99",X"00",X"EE",X"99",X"9B",X"90",X"9E",X"90",X"9E",X"90",X"9E",X"00",X"99",X"90",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"09",X"99",X"90",X"00",X"09",X"99",X"90",X"00",X"09",X"97",X"99",
		X"99",X"09",X"77",X"97",X"99",X"49",X"99",X"97",X"94",X"49",X"99",X"99",X"44",X"49",X"99",X"90",
		X"49",X"04",X"99",X"00",X"99",X"04",X"79",X"00",X"77",X"00",X"77",X"00",X"79",X"40",X"99",X"00",
		X"79",X"90",X"E9",X"00",X"99",X"94",X"EE",X"00",X"99",X"99",X"7E",X"00",X"99",X"79",X"77",X"00",
		X"94",X"79",X"77",X"00",X"94",X"77",X"77",X"00",X"99",X"77",X"77",X"00",X"99",X"77",X"77",X"00",
		X"77",X"77",X"77",X"00",X"99",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",
		X"09",X"77",X"77",X"00",X"99",X"77",X"77",X"00",X"97",X"77",X"77",X"00",X"77",X"97",X"79",X"00",
		X"77",X"99",X"99",X"00",X"99",X"44",X"97",X"00",X"94",X"99",X"77",X"00",X"44",X"49",X"77",X"00",
		X"00",X"00",X"09",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"93",X"00",X"00",X"99",X"99",X"09",
		X"00",X"79",X"77",X"00",X"99",X"79",X"99",X"00",X"77",X"99",X"9F",X"00",X"97",X"09",X"99",X"00",
		X"97",X"00",X"99",X"00",X"97",X"00",X"79",X"00",X"97",X"00",X"77",X"00",X"79",X"00",X"77",X"00",
		X"99",X"00",X"99",X"00",X"99",X"40",X"E7",X"00",X"F9",X"90",X"77",X"00",X"99",X"94",X"77",X"00",
		X"97",X"99",X"77",X"00",X"77",X"79",X"77",X"00",X"77",X"79",X"77",X"00",X"99",X"79",X"77",X"00",
		X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",
		X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"99",X"77",X"77",X"00",X"97",X"97",X"79",X"00",
		X"77",X"99",X"99",X"00",X"99",X"44",X"97",X"00",X"94",X"99",X"77",X"00",X"44",X"49",X"77",X"00",
		X"44",X"49",X"77",X"00",X"99",X"99",X"77",X"00",X"11",X"91",X"77",X"00",X"91",X"99",X"77",X"00",
		X"91",X"19",X"77",X"00",X"99",X"99",X"77",X"00",X"91",X"94",X"77",X"00",X"91",X"99",X"77",X"00",
		X"99",X"19",X"77",X"00",X"94",X"99",X"97",X"00",X"94",X"91",X"97",X"00",X"94",X"99",X"97",X"00",
		X"94",X"19",X"97",X"00",X"99",X"99",X"99",X"00",X"91",X"44",X"99",X"00",X"91",X"44",X"99",X"00",
		X"91",X"99",X"99",X"00",X"99",X"11",X"09",X"00",X"91",X"19",X"00",X"00",X"91",X"99",X"00",X"09",
		X"91",X"19",X"00",X"09",X"99",X"19",X"00",X"99",X"94",X"99",X"00",X"97",X"99",X"97",X"00",X"97",
		X"79",X"97",X"00",X"77",X"79",X"97",X"99",X"77",X"79",X"99",X"77",X"77",X"79",X"19",X"77",X"77",
		X"77",X"19",X"77",X"79",X"97",X"99",X"77",X"99",X"99",X"44",X"97",X"90",X"09",X"99",X"99",X"00",
		X"44",X"49",X"77",X"00",X"99",X"99",X"77",X"00",X"11",X"91",X"77",X"00",X"91",X"99",X"77",X"00",
		X"91",X"19",X"77",X"00",X"99",X"99",X"77",X"00",X"91",X"94",X"77",X"00",X"91",X"99",X"97",X"00",
		X"99",X"19",X"97",X"00",X"94",X"99",X"97",X"90",X"94",X"91",X"99",X"90",X"94",X"99",X"E9",X"99",
		X"94",X"19",X"79",X"79",X"99",X"99",X"79",X"79",X"91",X"44",X"99",X"99",X"91",X"44",X"90",X"00",
		X"91",X"99",X"90",X"99",X"99",X"11",X"00",X"79",X"91",X"19",X"00",X"79",X"91",X"99",X"00",X"79",
		X"91",X"19",X"00",X"79",X"99",X"19",X"00",X"79",X"94",X"99",X"99",X"99",X"99",X"97",X"77",X"00",
		X"79",X"97",X"77",X"00",X"79",X"97",X"77",X"00",X"79",X"99",X"77",X"00",X"79",X"19",X"77",X"00",
		X"97",X"19",X"77",X"00",X"99",X"99",X"79",X"00",X"09",X"44",X"90",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"29",X"00",X"90",X"99",X"29",X"99",
		X"99",X"99",X"29",X"99",X"99",X"99",X"29",X"90",X"99",X"99",X"29",X"00",X"99",X"99",X"29",X"90",
		X"99",X"92",X"99",X"99",X"99",X"92",X"29",X"90",X"99",X"92",X"99",X"00",X"99",X"29",X"99",X"09",
		X"99",X"29",X"99",X"99",X"99",X"29",X"99",X"99",X"99",X"29",X"99",X"99",X"99",X"22",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"90",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"22",X"99",X"00",X"99",X"22",X"99",X"00",
		X"99",X"22",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"29",X"00",
		X"90",X"99",X"29",X"00",X"99",X"99",X"29",X"00",X"99",X"99",X"29",X"00",X"99",X"99",X"29",X"90",
		X"99",X"92",X"99",X"99",X"99",X"92",X"29",X"90",X"99",X"92",X"99",X"00",X"99",X"29",X"99",X"00",
		X"99",X"29",X"99",X"00",X"99",X"29",X"99",X"99",X"99",X"29",X"99",X"99",X"99",X"22",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"90",
		X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"00",X"99",X"22",X"99",X"00",X"99",X"22",X"99",X"00",
		X"99",X"22",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"90",
		X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"29",X"99",X"99",X"99",X"22",
		X"99",X"99",X"D9",X"22",X"99",X"99",X"D9",X"22",X"99",X"99",X"D9",X"29",X"99",X"99",X"99",X"99",
		X"99",X"99",X"9D",X"90",X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"09",X"99",X"99",X"00",X"09",X"99",X"99",X"00",X"09",X"99",X"99",X"90",
		X"09",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"92",X"99",X"00",
		X"99",X"22",X"99",X"00",X"99",X"22",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"92",X"9D",X"00",X"99",X"99",X"D9",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"95",X"00",X"00",
		X"00",X"95",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"90",X"E9",X"00",X"00",X"99",X"EE",X"09",X"00",X"39",X"EE",X"99",X"00",X"39",X"99",X"93",X"00",
		X"33",X"9F",X"33",X"00",X"39",X"99",X"33",X"00",X"99",X"F9",X"39",X"00",X"99",X"F9",X"99",X"00",
		X"93",X"9F",X"99",X"00",X"39",X"9F",X"39",X"00",X"99",X"99",X"93",X"00",X"93",X"33",X"93",X"00",
		X"99",X"33",X"99",X"00",X"09",X"33",X"99",X"00",X"09",X"33",X"90",X"00",X"00",X"33",X"99",X"00",
		X"00",X"33",X"39",X"00",X"90",X"39",X"33",X"00",X"99",X"99",X"93",X"00",X"39",X"9B",X"99",X"00",
		X"33",X"33",X"93",X"00",X"99",X"33",X"33",X"00",X"00",X"99",X"39",X"00",X"00",X"99",X"99",X"00",
		X"00",X"33",X"00",X"00",X"99",X"33",X"00",X"00",X"33",X"39",X"00",X"00",X"93",X"99",X"00",X"00",
		X"93",X"99",X"90",X"00",X"99",X"00",X"99",X"00",X"09",X"00",X"39",X"00",X"09",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",
		X"99",X"00",X"99",X"00",X"D9",X"00",X"9D",X"00",X"9D",X"00",X"D9",X"00",X"9D",X"00",X"D9",X"90",
		X"99",X"00",X"99",X"90",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"DD",X"99",X"99",X"99",X"DD",X"99",X"99",
		X"99",X"DD",X"99",X"99",X"99",X"DD",X"99",X"99",X"09",X"99",X"99",X"99",X"09",X"99",X"99",X"09",
		X"09",X"99",X"09",X"09",X"00",X"99",X"09",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"09",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"D9",X"99",X"9D",X"00",X"9D",X"99",X"D9",X"00",
		X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"99",X"99",X"DD",X"99",X"99",
		X"99",X"DD",X"99",X"99",X"99",X"DD",X"99",X"99",X"99",X"DD",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"00",X"09",X"09",X"00",X"00",X"09",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",
		X"90",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"DD",X"99",X"99",X"00",X"DD",X"99",X"D9",X"00",X"9D",X"DD",X"D9",X"00",X"99",X"DD",X"99",X"00",
		X"99",X"DD",X"99",X"00",X"99",X"DD",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"09",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"AA",X"00",X"00",X"00",X"AF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"AA",X"0A",X"00",X"00",X"FF",X"AF",X"00",X"00",X"AA",X"AF",X"00",X"00",X"AF",X"FF",X"00",
		X"00",X"AF",X"FF",X"00",X"00",X"FF",X"AF",X"00",X"00",X"FF",X"AF",X"00",X"AA",X"FA",X"AA",X"00",
		X"FF",X"AA",X"FA",X"00",X"FF",X"AF",X"FF",X"A0",X"FF",X"FF",X"FF",X"A0",X"FF",X"FF",X"FF",X"A0",
		X"AF",X"AA",X"AF",X"00",X"AF",X"AF",X"AF",X"00",X"AF",X"AF",X"FF",X"00",X"FF",X"FF",X"AF",X"A0",
		X"FF",X"AA",X"AF",X"A0",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FA",X"00",X"AF",X"FF",X"FF",X"00",
		X"AF",X"FA",X"FF",X"00",X"AA",X"FA",X"FF",X"00",X"AA",X"FF",X"FA",X"00",X"FA",X"FF",X"AA",X"00",
		X"FA",X"AA",X"FF",X"00",X"AA",X"FA",X"FF",X"00",X"00",X"AA",X"FA",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"AA",X"00",
		X"FA",X"00",X"FF",X"A0",X"AA",X"00",X"FF",X"AA",X"A0",X"00",X"FF",X"FA",X"A0",X"00",X"FF",X"AA",
		X"00",X"00",X"FF",X"A0",X"00",X"00",X"AF",X"A0",X"00",X"AA",X"AA",X"A0",X"00",X"FF",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"FA",X"00",X"00",X"00",X"FA",X"00",X"00",X"00",X"A0",X"00",X"00",X"AA",X"00",X"00",X"00",
		X"FA",X"00",X"00",X"00",X"FA",X"00",X"00",X"00",X"AF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"AF",X"00",X"00",X"00",X"FF",X"00",X"0A",X"00",X"FF",X"00",X"0A",X"00",
		X"FF",X"00",X"0A",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"A0",X"00",X"00",X"00",X"A0",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",
		X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"00",X"F3",X"F0",X"33",X"00",
		X"F0",X"F0",X"00",X"00",X"FF",X"F0",X"FF",X"AA",X"F3",X"F0",X"33",X"00",X"F0",X"F0",X"00",X"00",
		X"F0",X"30",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",
		X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"0A",X"00",X"00",
		X"00",X"0A",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"0A",X"A0",X"A0",X"00",X"0A",X"A0",X"00",
		X"00",X"00",X"0A",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"FF",X"90",X"00",
		X"00",X"FF",X"90",X"00",X"00",X"F9",X"99",X"00",X"00",X"F9",X"59",X"00",X"00",X"99",X"59",X"00",
		X"00",X"9F",X"59",X"00",X"00",X"99",X"55",X"00",X"00",X"F9",X"F5",X"00",X"00",X"FF",X"F5",X"00",
		X"00",X"FF",X"F5",X"00",X"00",X"FF",X"F5",X"00",X"00",X"FF",X"F5",X"00",X"00",X"FF",X"F5",X"00",
		X"00",X"FF",X"F5",X"00",X"00",X"FF",X"F5",X"00",X"00",X"FF",X"F5",X"00",X"00",X"FF",X"59",X"00",
		X"00",X"FF",X"59",X"00",X"00",X"9F",X"59",X"00",X"00",X"9F",X"99",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"99",X"00",X"99",X"00",
		X"55",X"00",X"55",X"00",X"99",X"00",X"99",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"99",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"9F",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"F9",X"99",X"00",X"00",X"F9",X"59",X"00",X"00",X"99",X"59",X"00",
		X"00",X"9F",X"59",X"00",X"00",X"99",X"55",X"00",X"00",X"F9",X"F5",X"00",X"00",X"F9",X"95",X"00",
		X"00",X"99",X"99",X"00",X"00",X"9F",X"F5",X"00",X"00",X"99",X"F5",X"00",X"00",X"F9",X"F5",X"00",
		X"00",X"99",X"F5",X"00",X"00",X"9F",X"F5",X"00",X"00",X"FF",X"F5",X"00",X"00",X"FF",X"59",X"00",
		X"00",X"FF",X"59",X"00",X"00",X"9F",X"59",X"00",X"00",X"9F",X"99",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"99",X"00",X"99",X"00",
		X"55",X"00",X"55",X"00",X"99",X"00",X"99",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"99",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"9F",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"59",X"00",X"00",X"99",X"59",X"00",
		X"00",X"9F",X"99",X"00",X"00",X"99",X"95",X"00",X"00",X"F9",X"F5",X"00",X"00",X"F9",X"95",X"00",
		X"00",X"99",X"99",X"00",X"00",X"9F",X"F5",X"00",X"00",X"99",X"F5",X"00",X"00",X"F9",X"F9",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"95",X"00",X"00",X"FF",X"95",X"00",X"00",X"99",X"59",X"00",
		X"00",X"99",X"59",X"00",X"00",X"9F",X"99",X"00",X"00",X"9F",X"99",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"99",X"00",X"99",X"00",
		X"55",X"00",X"55",X"00",X"99",X"00",X"99",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"99",X"00",
		X"99",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",
		X"9F",X"09",X"00",X"00",X"9F",X"99",X"60",X"00",X"F9",X"99",X"93",X"90",X"99",X"29",X"90",X"90",
		X"00",X"99",X"93",X"90",X"00",X"99",X"A0",X"90",X"00",X"99",X"9A",X"00",X"02",X"99",X"94",X"00",
		X"00",X"99",X"9A",X"00",X"10",X"99",X"97",X"00",X"00",X"99",X"9A",X"50",X"00",X"99",X"A0",X"00",
		X"04",X"99",X"A0",X"00",X"90",X"99",X"30",X"00",X"F9",X"99",X"44",X"90",X"F9",X"9E",X"00",X"90",
		X"FF",X"0E",X"00",X"90",X"F9",X"0E",X"00",X"00",X"F9",X"0E",X"00",X"00",X"99",X"00",X"00",X"00",
		X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",
		X"03",X"50",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"09",X"00",X"09",X"00",X"09",X"90",X"09",X"00",X"00",X"99",X"09",X"00",
		X"90",X"94",X"09",X"00",X"99",X"94",X"99",X"00",X"A9",X"94",X"95",X"00",X"AA",X"44",X"55",X"00",
		X"AA",X"94",X"59",X"90",X"3A",X"A9",X"99",X"90",X"33",X"9A",X"AA",X"99",X"AA",X"AA",X"A3",X"A9",
		X"33",X"99",X"A3",X"39",X"3A",X"99",X"AA",X"A9",X"A5",X"44",X"9A",X"A9",X"33",X"44",X"99",X"59",
		X"3A",X"99",X"49",X"A9",X"3A",X"9F",X"49",X"39",X"A9",X"9F",X"49",X"A9",X"99",X"9F",X"49",X"39",
		X"90",X"9F",X"99",X"A9",X"90",X"9A",X"99",X"A9",X"00",X"99",X"90",X"A9",X"00",X"94",X"90",X"A9",
		X"00",X"49",X"99",X"39",X"00",X"99",X"59",X"A9",X"00",X"90",X"95",X"39",X"09",X"99",X"99",X"A9",
		X"09",X"59",X"59",X"A9",X"09",X"99",X"99",X"A9",X"00",X"00",X"59",X"A9",X"00",X"00",X"99",X"99",
		X"09",X"00",X"99",X"00",X"09",X"00",X"A9",X"00",X"09",X"90",X"A9",X"00",X"00",X"99",X"39",X"00",
		X"00",X"94",X"39",X"00",X"00",X"94",X"99",X"00",X"00",X"94",X"95",X"00",X"00",X"44",X"55",X"00",
		X"00",X"94",X"59",X"00",X"00",X"A9",X"99",X"00",X"00",X"9A",X"33",X"00",X"00",X"AA",X"AA",X"00",
		X"00",X"99",X"AA",X"00",X"00",X"99",X"A3",X"00",X"00",X"44",X"9A",X"00",X"00",X"44",X"99",X"00",
		X"00",X"99",X"49",X"00",X"00",X"9F",X"49",X"00",X"00",X"9F",X"49",X"00",X"00",X"9F",X"49",X"00",
		X"00",X"9F",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"93",X"00",X"00",X"94",X"9A",X"00",
		X"00",X"49",X"99",X"00",X"00",X"99",X"59",X"00",X"00",X"90",X"95",X"00",X"00",X"99",X"59",X"00",
		X"00",X"59",X"59",X"00",X"09",X"99",X"99",X"00",X"09",X"00",X"A9",X"00",X"09",X"00",X"9A",X"00",
		X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"09",X"00",X"00",X"99",X"09",X"00",
		X"00",X"94",X"99",X"00",X"00",X"94",X"99",X"00",X"00",X"94",X"95",X"00",X"00",X"44",X"55",X"00",
		X"00",X"94",X"A9",X"00",X"00",X"A9",X"99",X"00",X"00",X"AA",X"33",X"00",X"00",X"AA",X"AA",X"00",
		X"09",X"99",X"3A",X"00",X"09",X"99",X"A3",X"00",X"09",X"44",X"9A",X"00",X"09",X"44",X"99",X"00",
		X"09",X"99",X"49",X"00",X"09",X"9F",X"49",X"00",X"09",X"9F",X"49",X"00",X"99",X"9F",X"49",X"00",
		X"9A",X"9A",X"99",X"00",X"9A",X"99",X"99",X"00",X"9A",X"99",X"9A",X"00",X"9A",X"94",X"9A",X"00",
		X"9A",X"49",X"99",X"00",X"9A",X"99",X"59",X"00",X"9A",X"90",X"95",X"00",X"99",X"99",X"59",X"00",
		X"09",X"59",X"59",X"00",X"00",X"99",X"99",X"00",X"00",X"90",X"99",X"00",X"00",X"90",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"44",X"90",X"00",
		X"99",X"99",X"49",X"00",X"94",X"22",X"44",X"00",X"44",X"99",X"94",X"00",X"44",X"99",X"99",X"00",
		X"15",X"99",X"95",X"99",X"55",X"99",X"55",X"19",X"51",X"99",X"15",X"E9",X"11",X"17",X"11",X"99",
		X"91",X"77",X"11",X"90",X"EE",X"77",X"EE",X"00",X"99",X"77",X"EE",X"00",X"09",X"99",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"44",X"90",X"00",
		X"99",X"99",X"49",X"00",X"94",X"22",X"44",X"00",X"44",X"99",X"94",X"00",X"44",X"99",X"29",X"00",
		X"17",X"99",X"97",X"99",X"77",X"99",X"77",X"19",X"71",X"99",X"17",X"E9",X"11",X"15",X"11",X"99",
		X"91",X"55",X"11",X"90",X"EE",X"55",X"EE",X"00",X"99",X"55",X"EE",X"00",X"09",X"99",X"99",X"00",
		X"90",X"E0",X"00",X"00",X"90",X"EE",X"00",X"00",X"90",X"99",X"00",X"00",X"90",X"FF",X"90",X"00",
		X"99",X"F4",X"F9",X"00",X"39",X"FF",X"4F",X"00",X"33",X"FF",X"FF",X"00",X"39",X"99",X"FF",X"00",
		X"3B",X"99",X"F4",X"00",X"9B",X"FF",X"FF",X"00",X"93",X"FF",X"99",X"00",X"93",X"99",X"33",X"00",
		X"09",X"33",X"33",X"07",X"09",X"99",X"33",X"00",X"00",X"99",X"33",X"00",X"00",X"9F",X"33",X"00",
		X"50",X"99",X"33",X"00",X"00",X"33",X"33",X"00",X"00",X"3B",X"33",X"50",X"10",X"3B",X"99",X"00",
		X"11",X"39",X"99",X"00",X"A1",X"33",X"99",X"07",X"99",X"33",X"94",X"40",X"14",X"43",X"79",X"00",
		X"95",X"49",X"95",X"00",X"57",X"B5",X"54",X"50",X"71",X"45",X"11",X"45",X"49",X"17",X"A1",X"00",
		X"04",X"59",X"59",X"00",X"11",X"9A",X"55",X"00",X"05",X"0A",X"10",X"40",X"00",X"00",X"11",X"04",
		X"00",X"0E",X"E0",X"00",X"90",X"EE",X"E0",X"00",X"90",X"9E",X"00",X"00",X"90",X"33",X"E0",X"00",
		X"99",X"99",X"90",X"00",X"39",X"9A",X"99",X"00",X"33",X"AF",X"A3",X"00",X"39",X"FF",X"FF",X"00",
		X"3B",X"99",X"FF",X"00",X"9B",X"99",X"F9",X"00",X"93",X"FF",X"99",X"00",X"93",X"99",X"33",X"00",
		X"09",X"33",X"33",X"00",X"09",X"93",X"33",X"00",X"00",X"99",X"33",X"00",X"00",X"B9",X"33",X"00",
		X"00",X"3B",X"33",X"00",X"00",X"33",X"33",X"00",X"00",X"3B",X"33",X"00",X"00",X"3B",X"99",X"00",
		X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"09",X"33",X"90",X"00",X"99",X"33",X"99",X"00",
		X"33",X"33",X"39",X"00",X"39",X"93",X"99",X"00",X"99",X"93",X"93",X"00",X"09",X"19",X"33",X"00",
		X"00",X"39",X"33",X"00",X"00",X"39",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"90",X"90",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"FF",X"90",X"00",
		X"00",X"FF",X"90",X"00",X"00",X"FF",X"99",X"00",X"00",X"FF",X"59",X"00",X"00",X"FF",X"59",X"00",
		X"00",X"FF",X"59",X"00",X"00",X"FF",X"55",X"00",X"00",X"FF",X"F5",X"00",X"00",X"FF",X"F5",X"00",
		X"00",X"FF",X"F5",X"00",X"00",X"FF",X"F5",X"00",X"00",X"FF",X"F5",X"00",X"00",X"FF",X"F5",X"00",
		X"00",X"FF",X"F5",X"00",X"00",X"FF",X"F5",X"00",X"00",X"FF",X"F5",X"00",X"00",X"FF",X"59",X"00",
		X"00",X"FF",X"59",X"00",X"00",X"9F",X"59",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"99",X"00",X"99",X"00",
		X"55",X"00",X"55",X"00",X"99",X"00",X"99",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"90",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"09",X"99",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"90",X"99",X"00",X"00",X"90",X"49",X"00",X"00",X"99",X"49",X"00",
		X"09",X"BB",X"99",X"90",X"09",X"BB",X"9B",X"90",X"99",X"BB",X"BB",X"90",X"99",X"BB",X"B9",X"90",
		X"11",X"99",X"B9",X"90",X"E1",X"99",X"BB",X"00",X"EE",X"99",X"99",X"00",X"1E",X"99",X"59",X"00",
		X"1E",X"99",X"99",X"00",X"11",X"B9",X"99",X"99",X"11",X"BB",X"9B",X"B1",X"11",X"9B",X"BB",X"99",
		X"11",X"99",X"99",X"B9",X"11",X"BB",X"90",X"91",X"99",X"BB",X"90",X"99",X"9B",X"BB",X"90",X"90",
		X"BB",X"BB",X"90",X"00",X"9B",X"BB",X"90",X"00",X"9B",X"1B",X"99",X"00",X"99",X"9B",X"99",X"19",
		X"90",X"B9",X"9B",X"B9",X"90",X"B9",X"9B",X"19",X"90",X"BB",X"9B",X"B9",X"00",X"BB",X"99",X"99",
		X"00",X"BB",X"09",X"90",X"00",X"BB",X"09",X"00",X"00",X"9B",X"09",X"00",X"00",X"99",X"00",X"00",
		X"99",X"00",X"00",X"00",X"9E",X"00",X"99",X"00",X"99",X"00",X"39",X"00",X"19",X"99",X"39",X"00",
		X"11",X"BB",X"99",X"90",X"E1",X"BB",X"9B",X"90",X"EE",X"BB",X"BB",X"90",X"EE",X"BB",X"B9",X"90",
		X"1E",X"B9",X"B9",X"90",X"11",X"99",X"BB",X"00",X"11",X"99",X"99",X"00",X"11",X"99",X"59",X"90",
		X"11",X"B9",X"99",X"90",X"11",X"BB",X"BB",X"99",X"99",X"9B",X"99",X"B9",X"BB",X"99",X"BB",X"B9",
		X"B9",X"BB",X"BB",X"99",X"BB",X"BB",X"99",X"00",X"9B",X"BB",X"99",X"00",X"09",X"BB",X"90",X"00",
		X"00",X"BB",X"90",X"00",X"00",X"BB",X"90",X"00",X"00",X"1B",X"99",X"00",X"00",X"9B",X"99",X"19",
		X"00",X"B9",X"9B",X"B9",X"00",X"B9",X"9B",X"19",X"00",X"BB",X"9B",X"B9",X"00",X"BB",X"99",X"99",
		X"00",X"BB",X"09",X"90",X"00",X"BB",X"00",X"00",X"00",X"9B",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"90",X"00",
		X"00",X"66",X"99",X"00",X"99",X"66",X"69",X"00",X"99",X"66",X"99",X"00",X"EE",X"96",X"99",X"00",
		X"9E",X"99",X"96",X"00",X"49",X"E9",X"96",X"00",X"49",X"EC",X"96",X"00",X"99",X"E9",X"96",X"00",
		X"99",X"C9",X"96",X"00",X"CC",X"CC",X"96",X"00",X"CC",X"99",X"96",X"00",X"9C",X"C9",X"96",X"00",
		X"99",X"C9",X"99",X"00",X"99",X"C9",X"99",X"00",X"CC",X"C9",X"99",X"00",X"CC",X"99",X"66",X"00",
		X"9C",X"96",X"66",X"00",X"99",X"69",X"66",X"00",X"66",X"69",X"69",X"00",X"66",X"99",X"99",X"00",
		X"96",X"96",X"90",X"00",X"99",X"99",X"90",X"00",X"C9",X"CC",X"90",X"00",X"99",X"CC",X"90",X"00",
		X"00",X"99",X"99",X"00",X"00",X"97",X"79",X"00",X"00",X"97",X"79",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"90",X"00",
		X"09",X"66",X"99",X"00",X"99",X"66",X"69",X"00",X"EE",X"96",X"96",X"00",X"99",X"99",X"96",X"00",
		X"49",X"E9",X"96",X"00",X"49",X"EC",X"96",X"00",X"99",X"E9",X"96",X"00",X"99",X"C9",X"96",X"00",
		X"CC",X"CC",X"96",X"00",X"CC",X"99",X"96",X"00",X"9C",X"C9",X"96",X"00",X"99",X"C9",X"96",X"00",
		X"99",X"C9",X"96",X"00",X"99",X"C9",X"99",X"00",X"CC",X"99",X"99",X"00",X"9C",X"99",X"99",X"00",
		X"99",X"66",X"96",X"00",X"00",X"66",X"96",X"00",X"00",X"69",X"96",X"00",X"00",X"69",X"96",X"00",
		X"09",X"99",X"96",X"99",X"09",X"90",X"96",X"79",X"09",X"90",X"96",X"79",X"99",X"00",X"96",X"79",
		X"77",X"00",X"96",X"79",X"77",X"00",X"99",X"79",X"99",X"00",X"00",X"79",X"00",X"00",X"00",X"99",
		X"00",X"99",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"9E",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"99",X"99",X"99",X"00",X"9E",X"99",X"E9",X"00",X"9E",X"99",X"E9",X"99",X"BB",X"9E",X"EE",X"E9",
		X"BB",X"99",X"EE",X"99",X"99",X"99",X"E9",X"00",X"E9",X"99",X"99",X"90",X"E9",X"99",X"EE",X"90",
		X"E9",X"99",X"EE",X"90",X"EB",X"99",X"99",X"90",X"9B",X"99",X"9E",X"90",X"99",X"E9",X"9E",X"90",
		X"99",X"E9",X"99",X"00",X"99",X"E9",X"99",X"00",X"99",X"9E",X"90",X"00",X"9E",X"9E",X"99",X"00",
		X"9E",X"99",X"E9",X"00",X"99",X"09",X"E9",X"00",X"EE",X"09",X"EE",X"00",X"99",X"09",X"E9",X"00",
		X"E9",X"09",X"99",X"00",X"E9",X"00",X"9E",X"00",X"99",X"00",X"99",X"00",X"00",X"00",X"90",X"00",
		X"00",X"99",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"9E",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"09",X"99",X"99",X"00",X"99",X"99",X"E9",X"00",X"E9",X"99",X"EE",X"00",X"E9",X"9E",X"99",X"00",
		X"E9",X"99",X"E9",X"00",X"E9",X"99",X"E1",X"00",X"99",X"99",X"E9",X"90",X"E9",X"99",X"99",X"90",
		X"99",X"99",X"E9",X"99",X"9E",X"99",X"99",X"E9",X"9E",X"99",X"9E",X"E9",X"99",X"E9",X"99",X"99",
		X"9B",X"E9",X"90",X"99",X"9B",X"E9",X"90",X"E9",X"9B",X"9E",X"99",X"99",X"9E",X"9E",X"E9",X"90",
		X"9E",X"99",X"99",X"90",X"99",X"00",X"9B",X"00",X"49",X"00",X"EB",X"00",X"49",X"00",X"99",X"00",
		X"99",X"00",X"E9",X"00",X"9E",X"00",X"E9",X"90",X"9B",X"00",X"99",X"90",X"99",X"00",X"09",X"90",
		X"99",X"00",X"99",X"00",X"77",X"00",X"77",X"00",X"97",X"00",X"77",X"00",X"99",X"00",X"99",X"90",
		X"99",X"99",X"9F",X"99",X"97",X"79",X"99",X"79",X"77",X"79",X"99",X"79",X"77",X"79",X"99",X"99",
		X"79",X"77",X"77",X"90",X"99",X"77",X"99",X"00",X"97",X"77",X"99",X"00",X"77",X"77",X"77",X"00",
		X"77",X"77",X"77",X"90",X"77",X"77",X"77",X"99",X"77",X"99",X"97",X"79",X"97",X"94",X"97",X"79",
		X"94",X"94",X"97",X"79",X"94",X"94",X"97",X"79",X"9A",X"99",X"97",X"79",X"99",X"19",X"97",X"79",
		X"90",X"99",X"99",X"49",X"00",X"91",X"77",X"49",X"00",X"99",X"77",X"A9",X"00",X"91",X"97",X"99",
		X"00",X"91",X"99",X"90",X"00",X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"90",
		X"00",X"00",X"97",X"90",X"00",X"00",X"77",X"90",X"00",X"00",X"77",X"90",X"00",X"00",X"99",X"90",
		X"99",X"00",X"99",X"00",X"77",X"00",X"77",X"00",X"97",X"00",X"77",X"00",X"99",X"00",X"99",X"90",
		X"99",X"99",X"9F",X"99",X"99",X"79",X"99",X"79",X"99",X"79",X"99",X"79",X"49",X"79",X"49",X"99",
		X"97",X"77",X"49",X"90",X"77",X"77",X"97",X"00",X"99",X"77",X"77",X"00",X"09",X"77",X"99",X"00",
		X"99",X"77",X"77",X"00",X"97",X"77",X"77",X"00",X"97",X"99",X"77",X"00",X"97",X"94",X"77",X"00",
		X"77",X"94",X"77",X"00",X"77",X"94",X"77",X"00",X"77",X"99",X"77",X"00",X"77",X"19",X"79",X"90",
		X"77",X"99",X"49",X"90",X"77",X"91",X"49",X"90",X"77",X"99",X"79",X"99",X"77",X"91",X"79",X"99",
		X"77",X"99",X"A9",X"99",X"99",X"00",X"99",X"79",X"09",X"00",X"09",X"99",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"79",X"00",X"00",X"00",X"79",X"00",X"00",X"00",X"99",
		X"99",X"00",X"00",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"22",X"99",X"00",X"99",X"22",X"29",X"00",X"99",X"92",X"29",X"00",X"99",X"99",X"29",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"95",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"95",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"DD",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"90",X"00",X"99",X"99",X"90",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"00",X"09",X"99",X"00",
		X"00",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"90",X"29",X"00",X"99",X"99",X"29",X"00",
		X"99",X"22",X"29",X"00",X"09",X"92",X"22",X"00",X"09",X"99",X"92",X"00",X"99",X"99",X"92",X"00",
		X"99",X"49",X"29",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"90",X"99",X"59",X"99",X"90",
		X"09",X"99",X"99",X"90",X"09",X"99",X"99",X"90",X"99",X"99",X"99",X"90",X"99",X"59",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"9D",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"09",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"22",X"D9",X"00",X"00",X"29",X"D9",X"00",
		X"00",X"29",X"D9",X"00",X"09",X"29",X"D9",X"00",X"49",X"22",X"D9",X"99",X"92",X"22",X"D9",X"29",
		X"99",X"99",X"D9",X"29",X"09",X"95",X"99",X"99",X"00",X"99",X"99",X"90",X"99",X"99",X"22",X"90",
		X"92",X"99",X"2A",X"90",X"99",X"99",X"22",X"99",X"29",X"59",X"29",X"D9",X"A2",X"99",X"99",X"D9",
		X"99",X"22",X"9D",X"D9",X"99",X"99",X"9D",X"D9",X"DD",X"92",X"9D",X"90",X"DD",X"22",X"D2",X"00",
		X"D2",X"22",X"DD",X"00",X"2D",X"2A",X"DD",X"00",X"DD",X"22",X"D9",X"00",X"DD",X"22",X"99",X"00",
		X"9D",X"22",X"90",X"00",X"99",X"22",X"99",X"00",X"00",X"99",X"22",X"00",X"00",X"00",X"22",X"00",
		X"00",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"92",X"00",X"09",X"00",X"99",X"00",X"09",X"00",
		X"00",X"00",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"22",X"D9",X"00",X"00",X"29",X"D9",X"00",
		X"00",X"29",X"D9",X"00",X"09",X"29",X"D9",X"00",X"99",X"22",X"D9",X"00",X"92",X"22",X"D9",X"00",
		X"99",X"99",X"99",X"00",X"09",X"95",X"00",X"00",X"00",X"99",X"90",X"00",X"99",X"99",X"99",X"00",
		X"92",X"95",X"D9",X"00",X"99",X"99",X"D9",X"00",X"09",X"22",X"DD",X"00",X"00",X"99",X"2D",X"00",
		X"00",X"DD",X"DD",X"00",X"00",X"A2",X"DD",X"00",X"00",X"99",X"DD",X"00",X"00",X"92",X"D2",X"00",
		X"00",X"92",X"2D",X"00",X"00",X"99",X"DD",X"00",X"00",X"29",X"DD",X"00",X"00",X"D9",X"DD",X"00",
		X"00",X"99",X"DD",X"00",X"00",X"29",X"99",X"00",X"00",X"29",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"0E",X"E0",X"00",X"90",X"EE",X"E0",X"00",X"90",X"9E",X"00",X"00",X"90",X"33",X"E0",X"00",
		X"99",X"99",X"90",X"00",X"39",X"9F",X"99",X"00",X"33",X"FF",X"93",X"00",X"39",X"FF",X"93",X"00",
		X"3B",X"AF",X"93",X"00",X"9B",X"9A",X"93",X"00",X"93",X"99",X"39",X"00",X"93",X"33",X"33",X"00",
		X"09",X"33",X"33",X"00",X"09",X"99",X"33",X"00",X"00",X"93",X"33",X"00",X"00",X"99",X"33",X"00",
		X"00",X"39",X"33",X"00",X"00",X"33",X"33",X"00",X"00",X"3B",X"33",X"00",X"00",X"3B",X"99",X"00",
		X"00",X"39",X"99",X"00",X"99",X"33",X"44",X"00",X"94",X"33",X"94",X"00",X"44",X"93",X"99",X"00",
		X"15",X"99",X"95",X"99",X"55",X"B9",X"55",X"19",X"51",X"99",X"15",X"E9",X"11",X"17",X"11",X"99",
		X"91",X"77",X"11",X"90",X"EE",X"77",X"EE",X"00",X"99",X"77",X"EE",X"00",X"09",X"99",X"99",X"00",
		X"00",X"EE",X"E0",X"00",X"00",X"9E",X"00",X"00",X"90",X"E3",X"00",X"00",X"99",X"99",X"99",X"00",
		X"39",X"9F",X"39",X"00",X"33",X"F9",X"93",X"00",X"39",X"F9",X"93",X"00",X"3B",X"A9",X"93",X"00",
		X"9B",X"9F",X"93",X"00",X"93",X"99",X"39",X"00",X"93",X"33",X"33",X"00",X"09",X"33",X"33",X"00",
		X"09",X"99",X"33",X"00",X"00",X"93",X"33",X"00",X"00",X"99",X"33",X"00",X"00",X"99",X"33",X"00",
		X"00",X"33",X"33",X"00",X"00",X"33",X"33",X"00",X"00",X"3B",X"99",X"00",X"00",X"39",X"00",X"00",
		X"00",X"33",X"99",X"00",X"99",X"33",X"44",X"00",X"94",X"33",X"94",X"00",X"44",X"93",X"99",X"00",
		X"17",X"99",X"97",X"99",X"77",X"B9",X"77",X"19",X"71",X"99",X"17",X"E9",X"11",X"15",X"11",X"99",
		X"91",X"55",X"11",X"90",X"EE",X"55",X"EE",X"00",X"99",X"55",X"EE",X"00",X"09",X"99",X"99",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"9F",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"9A",X"99",X"00",X"00",X"9A",X"59",X"00",X"00",X"99",X"59",X"00",
		X"00",X"9F",X"99",X"00",X"00",X"99",X"95",X"00",X"00",X"F9",X"95",X"00",X"00",X"F9",X"95",X"00",
		X"00",X"99",X"99",X"00",X"00",X"94",X"F5",X"00",X"00",X"99",X"F5",X"00",X"00",X"F9",X"F9",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"95",X"00",X"00",X"F9",X"95",X"00",X"00",X"99",X"59",X"00",
		X"00",X"94",X"59",X"00",X"00",X"99",X"99",X"00",X"00",X"9F",X"99",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"99",X"00",X"99",X"00",
		X"55",X"00",X"55",X"00",X"99",X"00",X"99",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"99",X"00",
		X"99",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",
		X"9F",X"04",X"00",X"00",X"9F",X"94",X"60",X"00",X"F9",X"94",X"A3",X"90",X"99",X"29",X"90",X"90",
		X"00",X"94",X"93",X"90",X"00",X"99",X"A0",X"90",X"00",X"4A",X"9A",X"00",X"02",X"94",X"94",X"00",
		X"00",X"94",X"9A",X"00",X"10",X"99",X"97",X"00",X"00",X"49",X"9A",X"50",X"00",X"99",X"A0",X"00",
		X"04",X"9A",X"A0",X"00",X"90",X"4A",X"30",X"00",X"F9",X"49",X"44",X"90",X"F9",X"9A",X"00",X"90",
		X"FF",X"0E",X"00",X"90",X"F9",X"0E",X"00",X"00",X"F9",X"0E",X"00",X"00",X"99",X"00",X"00",X"00",
		X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",
		X"03",X"50",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
