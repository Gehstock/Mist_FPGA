library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity obj3 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of obj3 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"01",X"10",X"47",X"10",X"F0",X"0F",
		X"00",X"F0",X"1F",X"F1",X"1F",X"F1",X"F1",X"1F",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"0F",X"1E",X"10",X"47",X"10",X"01",X"00",
		X"D3",X"1F",X"F1",X"F1",X"1F",X"F1",X"1F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"21",X"12",X"21",X"9E",X"10",X"F0",X"0F",
		X"F1",X"2E",X"F1",X"2E",X"F1",X"F1",X"0F",X"69",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",
		X"03",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"0F",X"00",X"23",X"00",X"00",X"00",
		X"1F",X"F0",X"F0",X"0F",X"F0",X"0F",X"07",X"00",X"00",X"88",X"88",X"88",X"88",X"88",X"C4",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"31",X"52",X"3C",X"E1",X"96",X"78",X"70",X"61",
		X"00",X"88",X"88",X"88",X"C4",X"E2",X"2E",X"97",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"00",X"01",X"00",X"00",X"00",X"1E",X"0F",X"07",X"0F",X"06",X"00",X"11",X"00",
		X"1F",X"3C",X"F0",X"F0",X"C3",X"3C",X"01",X"00",X"00",X"88",X"88",X"CC",X"F3",X"86",X"08",X"00",
		X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"11",X"22",X"62",X"A6",X"79",X"D2",X"B4",X"78",X"61",
		X"00",X"00",X"00",X"00",X"88",X"C4",X"2E",X"5B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"43",X"87",X"0F",X"03",X"03",X"04",X"00",X"00",
		X"96",X"3C",X"78",X"69",X"12",X"44",X"00",X"00",X"88",X"C4",X"7B",X"C3",X"86",X"0C",X"00",X"00",
		X"22",X"13",X"12",X"34",X"25",X"21",X"12",X"12",X"00",X"00",X"88",X"EE",X"F1",X"E1",X"C3",X"C3",
		X"00",X"00",X"00",X"00",X"88",X"6E",X"3D",X"B4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",
		X"44",X"01",X"01",X"00",X"01",X"00",X"00",X"00",X"1E",X"0F",X"0F",X"0B",X"06",X"04",X"00",X"00",
		X"78",X"E1",X"A1",X"12",X"44",X"00",X"00",X"00",X"79",X"D2",X"A4",X"84",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"44",X"73",X"16",X"16",X"16",X"00",X"00",X"00",X"00",X"EE",X"79",X"69",X"69",
		X"00",X"00",X"00",X"00",X"CC",X"3F",X"B4",X"B4",X"00",X"00",X"00",X"00",X"00",X"55",X"FA",X"5A",
		X"12",X"01",X"11",X"00",X"00",X"00",X"00",X"00",X"69",X"07",X"07",X"07",X"04",X"05",X"01",X"00",
		X"3C",X"78",X"49",X"49",X"59",X"00",X"00",X"00",X"5A",X"5A",X"A4",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"88",X"7F",X"2D",X"2D",X"2D",X"00",X"00",X"00",X"00",X"FF",X"C3",X"D2",X"D2",
		X"00",X"00",X"00",X"00",X"FF",X"69",X"69",X"69",X"00",X"00",X"00",X"22",X"EC",X"A4",X"A4",X"A4",
		X"25",X"01",X"11",X"00",X"00",X"00",X"00",X"00",X"C3",X"07",X"07",X"06",X"02",X"02",X"00",X"00",
		X"69",X"49",X"59",X"48",X"08",X"08",X"00",X"00",X"84",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"AA",X"F5",X"A5",X"A5",X"00",X"00",X"00",X"33",X"CF",X"D2",X"D2",X"C3",
		X"00",X"00",X"00",X"77",X"E9",X"69",X"69",X"69",X"00",X"00",X"22",X"EC",X"86",X"86",X"86",X"84",
		X"A5",X"52",X"00",X"00",X"00",X"00",X"00",X"00",X"E1",X"29",X"29",X"A9",X"00",X"00",X"00",X"00",
		X"0E",X"0E",X"0E",X"02",X"0A",X"08",X"00",X"00",X"08",X"88",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"00",X"11",X"67",X"CB",X"D2",
		X"00",X"00",X"11",X"77",X"F8",X"78",X"3C",X"3C",X"88",X"8C",X"84",X"C2",X"4A",X"48",X"84",X"84",
		X"E9",X"B4",X"52",X"12",X"00",X"00",X"00",X"00",X"E1",X"78",X"78",X"84",X"22",X"00",X"00",X"00",
		X"87",X"0F",X"0F",X"0D",X"06",X"02",X"00",X"00",X"22",X"08",X"08",X"00",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"23",X"56",X"CB",
		X"23",X"23",X"74",X"DA",X"E1",X"78",X"3C",X"87",X"00",X"08",X"0C",X"84",X"80",X"08",X"44",X"00",
		X"11",X"76",X"52",X"21",X"10",X"00",X"00",X"00",X"E1",X"78",X"B4",X"C2",X"11",X"00",X"00",X"00",
		X"0F",X"0F",X"86",X"42",X"01",X"00",X"00",X"00",X"08",X"08",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"32",X"74",X"47",X"9E",
		X"C8",X"A4",X"C3",X"78",X"96",X"E1",X"C0",X"68",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",
		X"00",X"11",X"11",X"33",X"FC",X"16",X"01",X"00",X"8F",X"C3",X"F0",X"F0",X"3C",X"C3",X"08",X"00",
		X"87",X"0F",X"0E",X"0F",X"06",X"00",X"88",X"00",X"00",X"08",X"0C",X"00",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"74",X"23",X"74",X"23",X"74",X"74",X"8F",X"BC",
		X"C0",X"2C",X"C2",X"2C",X"C3",X"C0",X"78",X"0F",X"00",X"00",X"00",X"00",X"88",X"00",X"80",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"47",X"F8",X"F8",X"8F",X"F8",X"8F",X"87",X"00",
		X"0F",X"87",X"87",X"08",X"A6",X"08",X"00",X"00",X"06",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"07",
		X"00",X"08",X"08",X"0C",X"0C",X"0E",X"0E",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"66",X"44",X"44",X"77",X"33",X"00",
		X"00",X"66",X"FF",X"99",X"99",X"BB",X"22",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"08",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"11",X"10",X"30",
		X"00",X"00",X"00",X"00",X"FF",X"EE",X"E0",X"C0",X"00",X"00",X"00",X"00",X"08",X"08",X"40",X"40",
		X"20",X"20",X"11",X"11",X"00",X"00",X"00",X"00",X"30",X"07",X"07",X"0F",X"00",X"00",X"00",X"00",
		X"C0",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"11",X"11",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"10",X"30",X"00",X"00",X"00",X"00",X"FF",X"EE",X"E0",X"C0",
		X"00",X"00",X"00",X"00",X"08",X"08",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"11",X"10",X"30",
		X"30",X"07",X"07",X"0F",X"00",X"00",X"00",X"00",X"C0",X"08",X"08",X"00",X"00",X"00",X"00",X"00",
		X"20",X"20",X"11",X"11",X"00",X"00",X"00",X"00",X"30",X"07",X"07",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"EE",X"E0",X"C0",X"00",X"00",X"00",X"00",X"08",X"08",X"40",X"40",
		X"00",X"00",X"00",X"00",X"00",X"11",X"10",X"30",X"00",X"00",X"00",X"00",X"FF",X"EE",X"E0",X"C0",
		X"C0",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"11",X"11",X"00",X"00",X"00",X"00",
		X"30",X"07",X"07",X"0F",X"00",X"00",X"00",X"00",X"C0",X"08",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"EE",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"77",X"70",X"F0",
		X"00",X"00",X"00",X"00",X"CE",X"8A",X"90",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"81",X"45",X"47",X"00",X"00",X"00",X"00",X"F0",X"0E",X"0E",X"0C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"81",X"45",X"47",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"33",X"77",X"70",X"F0",X"00",X"00",X"00",X"00",X"CE",X"8A",X"90",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"77",X"70",X"F0",
		X"F0",X"0E",X"0E",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"81",X"45",X"47",X"00",X"00",X"00",X"00",X"F0",X"0E",X"0C",X"0C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"CE",X"8A",X"90",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"33",X"77",X"70",X"F0",X"00",X"00",X"00",X"00",X"CE",X"8A",X"90",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"81",X"45",X"47",X"00",X"00",X"00",X"00",
		X"F0",X"0E",X"0E",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"CE",X"8A",X"90",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"10",X"30",X"00",X"00",X"00",X"00",X"FF",X"EE",X"E0",X"C0",
		X"00",X"00",X"00",X"00",X"08",X"08",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"11",X"10",X"30",
		X"30",X"07",X"07",X"0F",X"00",X"00",X"00",X"00",X"C0",X"08",X"08",X"00",X"00",X"00",X"00",X"00",
		X"20",X"20",X"11",X"11",X"00",X"00",X"00",X"00",X"30",X"07",X"07",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"EE",X"E0",X"C0",X"00",X"00",X"00",X"00",X"08",X"08",X"40",X"40",
		X"00",X"00",X"00",X"00",X"00",X"11",X"10",X"30",X"00",X"00",X"00",X"00",X"FF",X"EE",X"E0",X"C0",
		X"C0",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"11",X"11",X"00",X"00",X"00",X"00",
		X"30",X"07",X"07",X"0F",X"00",X"00",X"00",X"00",X"C0",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"08",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"11",X"10",X"30",
		X"00",X"00",X"00",X"00",X"FF",X"EE",X"E0",X"C0",X"00",X"00",X"00",X"00",X"08",X"08",X"40",X"40",
		X"20",X"20",X"11",X"11",X"00",X"00",X"00",X"00",X"30",X"07",X"07",X"0F",X"00",X"00",X"00",X"00",
		X"C0",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"11",X"11",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"08",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"20",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"33",X"77",X"70",X"F0",X"00",X"00",X"00",X"00",X"CE",X"8A",X"90",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"77",X"70",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"81",X"45",X"47",X"00",X"00",X"00",X"00",X"F0",X"0E",X"0E",X"0C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"CE",X"8A",X"90",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"33",X"77",X"70",X"F0",X"00",X"00",X"00",X"00",X"CE",X"8A",X"90",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"81",X"45",X"47",X"00",X"00",X"00",X"00",
		X"F0",X"0E",X"0E",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"77",X"70",X"F0",
		X"00",X"00",X"00",X"00",X"CE",X"8A",X"90",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"81",X"45",X"47",X"00",X"00",X"00",X"00",X"F0",X"0E",X"0E",X"0C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"81",X"45",X"47",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"33",X"77",X"70",X"F0",X"00",X"00",X"00",X"00",X"CE",X"8A",X"90",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"77",X"70",X"F0",
		X"F0",X"0E",X"0E",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"81",X"45",X"47",X"00",X"00",X"00",X"00",X"F0",X"0E",X"0E",X"0C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"CE",X"8A",X"90",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"33",X"77",X"70",X"F0",X"00",X"00",X"00",X"00",X"CE",X"8A",X"90",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"81",X"45",X"47",X"00",X"00",X"00",X"00",
		X"F0",X"0E",X"0E",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"77",X"70",X"F0",
		X"00",X"00",X"00",X"00",X"CE",X"8A",X"90",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"81",X"45",X"47",X"00",X"00",X"00",X"00",X"F0",X"0E",X"0E",X"0C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"81",X"45",X"47",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"23",X"30",X"30",X"0F",
		X"00",X"00",X"03",X"70",X"0F",X"F0",X"C3",X"0E",X"00",X"00",X"0C",X"80",X"88",X"00",X"0C",X"00",
		X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"0F",X"30",X"30",X"23",X"00",X"00",X"00",
		X"05",X"0E",X"C3",X"F0",X"0F",X"70",X"03",X"00",X"00",X"00",X"0C",X"00",X"88",X"80",X"0C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"33",X"77",X"77",X"77",X"77",
		X"00",X"0F",X"0F",X"EE",X"EE",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"70",X"70",X"70",X"70",X"30",X"03",X"01",
		X"C0",X"00",X"00",X"C0",X"E0",X"E0",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"77",X"77",X"FF",X"FF",X"77",
		X"0C",X"0C",X"CC",X"CC",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"60",X"70",X"70",X"70",X"30",X"01",X"00",
		X"80",X"00",X"40",X"E0",X"E0",X"C3",X"0F",X"0C",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"00",
		X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"01",X"07",X"0F",X"3F",X"FF",X"FF",X"EE",X"FF",
		X"00",X"08",X"88",X"88",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"10",X"30",X"30",X"10",X"00",X"00",X"00",
		X"88",X"80",X"F0",X"F0",X"F0",X"C3",X"07",X"00",X"00",X"00",X"80",X"C2",X"0E",X"0C",X"08",X"00",
		X"00",X"00",X"01",X"03",X"03",X"11",X"11",X"11",X"04",X"0E",X"2E",X"7F",X"FF",X"EE",X"EE",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"54",X"30",X"10",X"00",X"00",X"00",X"00",
		X"90",X"F0",X"F0",X"F0",X"E1",X"01",X"00",X"00",X"80",X"C2",X"87",X"0E",X"0C",X"08",X"00",X"00",
		X"00",X"01",X"03",X"07",X"17",X"17",X"37",X"33",X"00",X"08",X"88",X"CC",X"CC",X"CC",X"CC",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C2",
		X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"DC",X"10",X"00",X"00",X"00",X"00",X"00",
		X"B0",X"F0",X"F0",X"F0",X"01",X"00",X"00",X"00",X"87",X"86",X"0E",X"0C",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"06",X"06",X"17",X"3F",X"3F",X"00",X"00",X"00",X"00",X"00",X"88",X"CC",X"98",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"C3",X"C3",
		X"37",X"33",X"11",X"00",X"00",X"00",X"00",X"00",X"DC",X"EE",X"FE",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"60",X"00",X"00",X"00",X"00",X"86",X"86",X"86",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"17",X"17",X"17",X"00",X"00",X"00",X"00",X"00",X"88",X"CC",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"90",X"00",X"00",X"00",X"00",X"03",X"C3",X"C3",X"C3",
		X"17",X"13",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"70",X"F0",X"70",X"00",X"00",X"00",X"00",X"00",X"C3",X"C2",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"47",X"70",X"70",X"F0",
		X"00",X"00",X"00",X"F0",X"1F",X"F0",X"F0",X"C0",X"00",X"00",X"00",X"80",X"88",X"00",X"00",X"00",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"F0",X"70",X"70",X"47",X"00",X"00",X"00",
		X"80",X"C0",X"F0",X"F0",X"1F",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"07",X"F8",X"F0",X"70",
		X"00",X"00",X"70",X"B7",X"68",X"E0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"F0",X"70",X"30",X"23",X"00",X"00",X"00",
		X"80",X"F0",X"F0",X"C3",X"3C",X"00",X"00",X"00",X"00",X"80",X"80",X"CC",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"10",X"30",X"43",X"3C",X"F0",X"F0",X"E0",
		X"80",X"C4",X"C8",X"C0",X"C0",X"80",X"80",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"D0",X"F0",X"F0",X"10",X"11",X"00",X"00",X"00",
		X"F0",X"E1",X"87",X"3C",X"00",X"00",X"00",X"00",X"C4",X"E8",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"11",X"00",X"10",X"31",X"53",X"96",X"3C",X"78",X"F0",
		X"00",X"00",X"88",X"80",X"C0",X"80",X"90",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C4",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"D0",X"70",X"B0",X"00",X"00",X"00",X"00",
		X"F0",X"E1",X"C3",X"96",X"8C",X"00",X"00",X"00",X"EC",X"48",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"71",X"72",X"96",X"B4",X"3C",X"78",
		X"00",X"00",X"00",X"00",X"80",X"00",X"90",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"E2",X"F4",
		X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"60",X"70",X"70",X"40",X"00",X"00",X"00",
		X"70",X"F0",X"E1",X"E1",X"22",X"00",X"00",X"00",X"68",X"48",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"10",X"10",X"10",X"01",X"01",X"00",X"00",X"88",X"E8",X"68",X"68",X"E0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"30",X"F0",X"E1",X"00",X"00",X"00",X"00",X"C8",X"C8",X"48",X"80",
		X"01",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"70",X"30",X"20",X"00",X"00",X"00",
		X"E1",X"E1",X"E1",X"62",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"00",X"00",X"00",X"88",X"E8",X"68",X"78",X"78",
		X"00",X"00",X"00",X"00",X"30",X"30",X"70",X"F0",X"00",X"00",X"00",X"C8",X"C8",X"48",X"48",X"48",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"78",X"78",X"F8",X"10",X"00",X"00",X"00",X"00",
		X"70",X"70",X"F0",X"C0",X"80",X"00",X"00",X"00",X"08",X"08",X"88",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"77",X"EF",X"E1",X"00",X"00",X"00",X"00",X"00",X"CC",X"0F",X"00",
		X"0F",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"11",X"00",X"00",X"00",X"00",X"00",
		X"02",X"0F",X"EF",X"77",X"00",X"00",X"00",X"00",X"0C",X"00",X"0F",X"CC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"23",
		X"00",X"00",X"00",X"00",X"77",X"CF",X"8F",X"0E",X"00",X"00",X"00",X"00",X"8E",X"08",X"00",X"0C",
		X"11",X"01",X"0F",X"00",X"00",X"00",X"00",X"00",X"87",X"0F",X"48",X"00",X"00",X"00",X"00",X"00",
		X"03",X"2F",X"FF",X"00",X"00",X"00",X"00",X"00",X"03",X"0C",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"32",
		X"00",X"00",X"00",X"33",X"47",X"CE",X"8E",X"0B",X"00",X"00",X"00",X"0C",X"00",X"04",X"09",X"06",
		X"00",X"00",X"00",X"03",X"06",X"00",X"00",X"00",X"61",X"C3",X"0F",X"0C",X"00",X"00",X"00",X"00",
		X"07",X"7F",X"FF",X"00",X"00",X"00",X"00",X"00",X"6E",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"33",X"23",X"23",
		X"00",X"01",X"CE",X"8C",X"0D",X"0C",X"0B",X"07",X"00",X"00",X"00",X"00",X"02",X"04",X"4C",X"CC",
		X"00",X"00",X"10",X"00",X"01",X"02",X"00",X"00",X"47",X"8F",X"0F",X"0E",X"40",X"00",X"00",X"00",
		X"3F",X"6E",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"23",X"23",X"67",X"67",X"46",
		X"04",X"08",X"0A",X"04",X"09",X"0F",X"37",X"6E",X"00",X"00",X"08",X"08",X"88",X"88",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"43",X"07",X"97",X"2C",X"08",X"08",X"00",X"00",
		X"4C",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"46",X"46",X"47",X"67",X"46",X"46",
		X"00",X"01",X"09",X"1B",X"17",X"1F",X"3F",X"6E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"43",X"16",X"17",X"04",X"04",X"04",
		X"4C",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"46",X"46",X"47",X"76",X"76",X"32",
		X"02",X"02",X"1B",X"1B",X"17",X"3F",X"37",X"26",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"32",X"11",X"11",X"11",X"10",X"00",X"00",X"00",
		X"2E",X"0C",X"0C",X"0C",X"48",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"23",X"30",X"30",X"0F",
		X"00",X"00",X"03",X"70",X"0F",X"F0",X"C3",X"0E",X"00",X"00",X"0C",X"80",X"88",X"00",X"0C",X"00",
		X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"0F",X"30",X"30",X"23",X"00",X"00",X"00",
		X"05",X"0E",X"C3",X"F0",X"0F",X"70",X"03",X"00",X"00",X"00",X"0C",X"00",X"88",X"80",X"0C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"21",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"48",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"84",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"0F",
		X"00",X"00",X"08",X"08",X"08",X"08",X"0C",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"03",X"01",X"01",X"01",X"01",X"00",X"00",
		X"0F",X"0C",X"08",X"08",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"10",X"10",X"30",X"70",X"E1",
		X"00",X"80",X"80",X"80",X"80",X"C0",X"E0",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E1",X"70",X"30",X"10",X"10",X"10",X"10",X"00",
		X"78",X"E0",X"C0",X"80",X"80",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"11",X"11",X"33",X"77",X"EF",
		X"00",X"88",X"88",X"88",X"88",X"CC",X"EE",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",
		X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EF",X"77",X"33",X"11",X"11",X"11",X"11",X"00",
		X"7F",X"EE",X"CC",X"88",X"88",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"10",X"10",X"30",X"F0",X"F0",
		X"80",X"80",X"80",X"80",X"C0",X"C0",X"E0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"70",X"30",X"30",X"10",X"10",X"10",X"10",
		X"F0",X"F0",X"C0",X"80",X"80",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"40",X"00",X"00",
		X"00",X"00",X"00",X"08",X"00",X"40",X"00",X"20",X"00",X"01",X"00",X"80",X"00",X"10",X"00",X"40",
		X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"08",X"20",X"00",X"00",X"00",X"80",
		X"80",X"10",X"20",X"00",X"80",X"20",X"00",X"A2",X"50",X"00",X"11",X"80",X"AA",X"55",X"88",X"BB",
		X"00",X"08",X"00",X"10",X"00",X"80",X"00",X"20",X"00",X"00",X"00",X"01",X"00",X"20",X"00",X"40",
		X"00",X"00",X"00",X"00",X"01",X"20",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A0",X"00",X"88",X"10",X"55",X"AA",X"11",X"DD",X"10",X"80",X"40",X"00",X"10",X"40",X"00",X"54",
		X"00",X"00",X"01",X"40",X"00",X"00",X"00",X"10",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"01",
		X"04",X"00",X"00",X"10",X"00",X"00",X"00",X"01",X"40",X"00",X"10",X"00",X"00",X"10",X"40",X"00",
		X"A2",X"00",X"80",X"10",X"40",X"20",X"00",X"80",X"55",X"99",X"44",X"BB",X"00",X"51",X"00",X"90",
		X"00",X"00",X"00",X"00",X"00",X"02",X"04",X"00",X"00",X"00",X"40",X"08",X"00",X"00",X"00",X"00",
		X"00",X"10",X"00",X"02",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"01",
		X"AA",X"99",X"22",X"DD",X"00",X"A8",X"00",X"90",X"54",X"00",X"10",X"80",X"20",X"40",X"00",X"10",
		X"20",X"00",X"80",X"00",X"00",X"80",X"20",X"00",X"02",X"00",X"00",X"80",X"00",X"00",X"00",X"08",
		X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"08",X"00",X"80",X"00",X"04",X"00",X"02",X"00",X"00",
		X"00",X"00",X"20",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"11",
		X"00",X"00",X"00",X"10",X"00",X"04",X"00",X"22",X"00",X"00",X"11",X"00",X"00",X"00",X"40",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"08",X"20",X"00",X"00",X"00",X"22",
		X"00",X"54",X"00",X"01",X"08",X"22",X"00",X"04",X"44",X"00",X"10",X"80",X"00",X"45",X"08",X"91",
		X"00",X"00",X"88",X"00",X"00",X"00",X"20",X"08",X"00",X"00",X"00",X"80",X"00",X"02",X"00",X"44",
		X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"00",X"80",X"10",X"00",X"2A",X"01",X"98",X"00",X"A2",X"00",X"08",X"01",X"44",X"00",X"02",
		X"00",X"00",X"01",X"40",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",
		X"22",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"01",X"00",X"20",X"00",X"00",X"11",X"04",X"00",
		X"20",X"00",X"88",X"10",X"41",X"00",X"44",X"00",X"15",X"00",X"44",X"12",X"00",X"44",X"01",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"80",X"00",X"00",X"00",X"00",
		X"00",X"10",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"01",X"00",X"00",
		X"8A",X"00",X"22",X"84",X"00",X"22",X"08",X"01",X"40",X"00",X"11",X"80",X"28",X"00",X"22",X"00",
		X"08",X"00",X"40",X"00",X"00",X"88",X"02",X"00",X"44",X"00",X"00",X"00",X"80",X"00",X"00",X"00",
		X"00",X"88",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"80",X"00",X"04",X"00",X"00",X"00",X"00",
		X"88",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"30",X"70",
		X"00",X"00",X"00",X"00",X"00",X"88",X"CC",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"13",X"03",
		X"00",X"00",X"00",X"00",X"00",X"22",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"12",X"04",X"00",X"00",X"00",X"00",X"00",
		X"C4",X"C0",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"F0",
		X"00",X"00",X"00",X"00",X"88",X"88",X"CC",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"03",X"01",X"01",X"00",X"00",X"00",X"00",
		X"F0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"40",X"66",X"10",X"22",X"44",X"20",X"00",X"10",X"00",X"04",X"54",X"A8",X"A7",X"5C",X"B1",
		X"04",X"08",X"46",X"28",X"27",X"A8",X"41",X"3A",X"00",X"00",X"44",X"00",X"51",X"0A",X"00",X"41",
		X"15",X"22",X"02",X"00",X"02",X"11",X"40",X"00",X"46",X"49",X"B9",X"32",X"0A",X"A8",X"00",X"22",
		X"A1",X"15",X"0A",X"51",X"A8",X"04",X"22",X"80",X"8A",X"04",X"A2",X"19",X"02",X"48",X"00",X"01",
		X"00",X"00",X"00",X"22",X"01",X"00",X"00",X"00",X"10",X"00",X"00",X"11",X"00",X"00",X"41",X"08",
		X"00",X"00",X"00",X"00",X"80",X"02",X"00",X"8A",X"11",X"00",X"00",X"80",X"00",X"00",X"00",X"81",
		X"91",X"00",X"00",X"00",X"00",X"20",X"00",X"08",X"14",X"02",X"00",X"98",X"00",X"00",X"00",X"00",
		X"09",X"40",X"88",X"01",X"00",X"80",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"11",X"00",X"90",X"31",X"63",
		X"00",X"00",X"00",X"00",X"22",X"88",X"C4",X"6C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"81",
		X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"65",X"33",X"10",X"44",X"00",X"00",X"00",X"00",
		X"6A",X"C4",X"98",X"00",X"88",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"01",X"32",X"65",
		X"00",X"00",X"00",X"00",X"00",X"88",X"C0",X"AF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5B",X"32",X"01",X"00",X"00",X"00",X"00",X"00",
		X"E4",X"8C",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"0A",X"12",X"10",
		X"00",X"04",X"00",X"08",X"04",X"03",X"00",X"81",X"00",X"80",X"08",X"00",X"00",X"00",X"28",X"26",
		X"20",X"01",X"00",X"00",X"00",X"14",X"82",X"12",X"00",X"00",X"14",X"82",X"10",X"24",X"90",X"24",
		X"4A",X"70",X"54",X"F9",X"30",X"1A",X"30",X"F2",X"D0",X"EB",X"F1",X"B4",X"F2",X"F9",X"F4",X"FB",
		X"00",X"00",X"00",X"04",X"00",X"04",X"04",X"20",X"00",X"00",X"00",X"80",X"08",X"01",X"42",X"00",
		X"00",X"00",X"14",X"80",X"48",X"00",X"01",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",
		X"04",X"70",X"C6",X"B4",X"5A",X"FB",X"F4",X"FD",X"94",X"40",X"A0",X"79",X"B4",X"68",X"E9",X"F5",
		X"00",X"20",X"8F",X"82",X"E8",X"80",X"05",X"82",X"40",X"08",X"90",X"02",X"00",X"80",X"00",X"00",
		X"00",X"00",X"00",X"02",X"01",X"20",X"04",X"20",X"20",X"00",X"00",X"5C",X"71",X"85",X"13",X"00",
		X"21",X"10",X"F9",X"D6",X"50",X"B3",X"45",X"B8",X"FA",X"F5",X"F0",X"F5",X"F0",X"C2",X"AA",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"10",X"11",X"01",X"02",X"10",X"42",X"80",
		X"A1",X"C8",X"14",X"80",X"09",X"00",X"00",X"00",X"32",X"A3",X"68",X"82",X"04",X"31",X"01",X"10",
		X"FA",X"F5",X"F0",X"FA",X"F0",X"E5",X"F0",X"FA",X"F2",X"E5",X"E8",X"C2",X"F9",X"A1",X"52",X"BC",
		X"60",X"3A",X"14",X"A0",X"21",X"80",X"44",X"C8",X"00",X"02",X"18",X"08",X"00",X"00",X"48",X"10",
		X"C2",X"45",X"92",X"6C",X"81",X"50",X"04",X"40",X"85",X"50",X"20",X"84",X"24",X"21",X"10",X"04",
		X"04",X"B8",X"06",X"42",X"21",X"10",X"00",X"80",X"00",X"00",X"00",X"08",X"80",X"48",X"20",X"00",
		X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"80",X"00",X"00",X"40",X"20",X"40",
		X"01",X"08",X"00",X"10",X"80",X"00",X"00",X"20",X"00",X"00",X"40",X"10",X"00",X"40",X"00",X"80",
		X"40",X"20",X"00",X"10",X"00",X"10",X"00",X"28",X"40",X"A0",X"00",X"40",X"A0",X"40",X"90",X"40",
		X"80",X"20",X"80",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"00",X"00",X"00",X"A0",X"00",X"10",X"00",X"80",X"00",X"40",X"00",X"90",X"20",X"10",
		X"00",X"01",X"20",X"00",X"00",X"20",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",
		X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",
		X"10",X"40",X"00",X"A0",X"40",X"80",X"00",X"A0",X"00",X"00",X"80",X"80",X"00",X"C0",X"00",X"40",
		X"28",X"00",X"10",X"00",X"10",X"00",X"20",X"40",X"40",X"90",X"40",X"A0",X"40",X"00",X"A0",X"40",
		X"00",X"00",X"00",X"00",X"00",X"80",X"20",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"40",X"20",X"40",X"00",X"00",X"80",X"00",X"40",
		X"20",X"00",X"00",X"80",X"10",X"00",X"08",X"01",X"80",X"00",X"40",X"00",X"10",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"40",X"90",X"00",X"20",X"10",X"40",X"00",X"30",X"80",X"20",
		X"20",X"90",X"20",X"50",X"00",X"20",X"00",X"90",X"40",X"00",X"80",X"01",X"40",X"80",X"00",X"20",
		X"20",X"80",X"10",X"40",X"00",X"A0",X"00",X"00",X"D0",X"00",X"50",X"60",X"80",X"40",X"00",X"80",
		X"20",X"50",X"00",X"00",X"40",X"00",X"20",X"01",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",
		X"00",X"08",X"00",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0E",X"01",
		X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"01",
		X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"01",X"00",X"00",X"01",X"01",X"00",X"05",
		X"1C",X"2D",X"58",X"93",X"59",X"B3",X"62",X"95",X"2C",X"C5",X"62",X"DD",X"44",X"99",X"44",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"81",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"02",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"82",X"9C",X"A8",X"55",X"AA",X"11",X"22",X"11",X"0B",X"61",X"0A",X"61",X"B0",X"46",X"BA",X"45",
		X"08",X"00",X"00",X"00",X"00",X"08",X"00",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1A",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"51",X"2A",X"51",X"39",X"52",X"06",X"1E",X"08",X"44",X"AA",X"CC",X"22",X"55",X"F5",X"18",X"25",
		X"00",X"04",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"04",X"00",X"00",X"00",X"00",X"00",
		X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"11",X"77",X"DD",X"AA",X"50",X"21",X"4A",X"A9",X"54",X"A8",X"42",X"A1",X"14",X"A1",X"05",
		X"08",X"00",X"08",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",
		X"00",X"08",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",
		X"0C",X"04",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"08",X"00",X"01",X"00",
		X"04",X"00",X"00",X"20",X"00",X"00",X"02",X"41",X"01",X"00",X"40",X"10",X"04",X"00",X"10",X"20",
		X"08",X"04",X"10",X"00",X"00",X"02",X"00",X"00",X"08",X"20",X"20",X"00",X"08",X"10",X"00",X"80",
		X"00",X"40",X"11",X"00",X"44",X"00",X"00",X"88",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"00",X"00",X"01",X"02",X"00",X"00",X"00",X"01",X"00",X"00",X"01",X"40",X"80",X"00",
		X"08",X"00",X"00",X"00",X"00",X"00",X"04",X"08",X"00",X"00",X"00",X"04",X"08",X"00",X"00",X"00",
		X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"10",X"22",X"00",X"00",X"00",
		X"00",X"80",X"01",X"04",X"20",X"00",X"01",X"82",X"09",X"02",X"00",X"00",X"00",X"03",X"00",X"00",
		X"18",X"04",X"00",X"00",X"01",X"00",X"04",X"08",X"20",X"00",X"00",X"20",X"08",X"00",X"00",X"00",
		X"00",X"00",X"88",X"00",X"00",X"11",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"51",X"00",
		X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"08",X"00",X"01",X"02",X"00",X"00",X"00",X"00",
		X"00",X"10",X"00",X"01",X"00",X"00",X"04",X"08",X"00",X"20",X"00",X"00",X"00",X"00",X"02",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"11",X"00",X"00",X"88",X"00",X"20",X"10",
		X"00",X"00",X"40",X"00",X"18",X"00",X"02",X"02",X"00",X"00",X"00",X"04",X"02",X"00",X"00",X"00",
		X"80",X"00",X"02",X"09",X"00",X"00",X"02",X"00",X"00",X"02",X"01",X"00",X"00",X"00",X"02",X"02",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"08",X"00",X"00",X"00",
		X"00",X"00",X"04",X"02",X"01",X"00",X"00",X"03",X"01",X"01",X"01",X"12",X"1E",X"59",X"F3",X"F7",
		X"00",X"08",X"00",X"08",X"87",X"CA",X"ED",X"FE",X"00",X"00",X"04",X"08",X"00",X"00",X"00",X"0B",
		X"0F",X"01",X"00",X"00",X"01",X"00",X"04",X"00",X"F7",X"7B",X"14",X"0F",X"01",X"01",X"00",X"00",
		X"FC",X"D8",X"A1",X"0C",X"08",X"00",X"08",X"08",X"0C",X"08",X"00",X"08",X"04",X"00",X"00",X"00",
		X"08",X"06",X"03",X"03",X"00",X"01",X"10",X"03",X"00",X"00",X"03",X"68",X"D1",X"F3",X"B3",X"73",
		X"08",X"08",X"C2",X"74",X"DC",X"FF",X"FF",X"EE",X"01",X"06",X"0C",X"08",X"80",X"84",X"40",X"8A",
		X"00",X"01",X"00",X"01",X"01",X"07",X"06",X"08",X"E6",X"51",X"59",X"1A",X"3C",X"00",X"00",X"00",
		X"FF",X"FF",X"A8",X"D4",X"25",X"4A",X"08",X"00",X"84",X"40",X"C0",X"08",X"0C",X"04",X"00",X"01",
		X"00",X"00",X"01",X"03",X"03",X"11",X"11",X"11",X"04",X"0E",X"2E",X"7F",X"FF",X"EE",X"EE",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"54",X"30",X"10",X"00",X"00",X"00",X"00",
		X"90",X"F0",X"F0",X"F0",X"E1",X"01",X"00",X"00",X"80",X"C2",X"87",X"0E",X"0C",X"08",X"00",X"00",
		X"00",X"01",X"03",X"07",X"17",X"17",X"37",X"33",X"00",X"08",X"88",X"CC",X"CC",X"CC",X"CC",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C2",
		X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"DC",X"10",X"00",X"00",X"00",X"00",X"00",
		X"B0",X"F0",X"F0",X"F0",X"01",X"00",X"00",X"00",X"87",X"86",X"0E",X"0C",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"CC",X"88",
		X"00",X"00",X"00",X"00",X"00",X"EE",X"11",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"CC",X"88",
		X"00",X"00",X"00",X"00",X"00",X"EE",X"11",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"77",X"CC",X"88",X"77",X"00",X"06",
		X"EE",X"00",X"EE",X"11",X"33",X"EE",X"00",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"68",X"14",X"00",X"00",X"00",X"00",X"00",
		X"F1",X"49",X"C7",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"77",X"CC",X"88",X"77",X"00",X"46",
		X"EE",X"00",X"EE",X"11",X"33",X"EE",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"76",X"00",X"00",X"F0",X"00",X"00",
		X"11",X"11",X"EE",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"03",X"06",X"0C",X"00",X"00",
		X"03",X"06",X"0C",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"03",X"06",X"06",X"0C",X"08",X"09",
		X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"0F",X"03",X"02",X"02",X"02",X"02",X"02",X"01",X"03",X"03",X"06",X"04",X"04",X"04",X"04",
		X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"02",X"02",X"02",X"01",X"01",X"01",X"00",X"07",X"07",X"06",X"05",X"01",X"02",X"0E",X"08",
		X"0E",X"01",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"0C",
		X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"07",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"01",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"0F",X"03",X"00",
		X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",
		X"00",X"00",X"00",X"0E",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"0F",X"01",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"0C",X"04",X"06",X"02",X"03",X"01",X"01",
		X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",
		X"0C",X"06",X"03",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"08",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"00",X"07",X"07",X"03",X"00",X"00",X"00",X"00",
		X"0E",X"0E",X"03",X"0F",X"01",X"00",X"00",X"00",X"0D",X"0C",X"06",X"02",X"00",X"00",X"00",X"00",
		X"08",X"04",X"04",X"04",X"06",X"02",X"02",X"01",X"00",X"07",X"0C",X"0C",X"0C",X"06",X"06",X"03",
		X"00",X"0F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"03",X"0F",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"03",X"0C",X"00",X"03",X"01",
		X"03",X"06",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"03",X"00",X"00",X"00",
		X"00",X"00",X"07",X"0F",X"08",X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"03",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"0C",X"00",X"00",X"00",X"07",X"06",X"03",X"01",X"00",
		X"00",X"00",X"00",X"01",X"0E",X"00",X"00",X"00",X"00",X"00",X"03",X"0C",X"00",X"00",X"00",X"00",
		X"04",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"00",X"00",X"01",X"07",X"0C",X"00",X"00",X"03",X"06",X"0C",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"32",
		X"00",X"00",X"00",X"33",X"47",X"CE",X"8E",X"0B",X"00",X"00",X"00",X"0C",X"00",X"04",X"09",X"06",
		X"00",X"00",X"00",X"03",X"06",X"00",X"00",X"00",X"61",X"C3",X"0F",X"0C",X"00",X"00",X"00",X"00",
		X"07",X"7F",X"FF",X"00",X"00",X"00",X"00",X"00",X"6E",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"33",X"23",X"23",
		X"00",X"01",X"CE",X"8C",X"0D",X"0C",X"0B",X"07",X"00",X"00",X"00",X"00",X"02",X"04",X"4C",X"CC",
		X"00",X"00",X"10",X"00",X"01",X"02",X"00",X"00",X"47",X"8F",X"0F",X"0E",X"40",X"00",X"00",X"00",
		X"3F",X"6E",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"23",X"23",X"67",X"67",X"46",
		X"04",X"08",X"0A",X"04",X"09",X"0F",X"37",X"6E",X"00",X"00",X"08",X"08",X"88",X"88",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"43",X"07",X"97",X"2C",X"08",X"08",X"00",X"00",
		X"4C",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"CC",X"88",
		X"00",X"00",X"00",X"00",X"00",X"EE",X"11",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"46",X"46",X"47",X"76",X"76",X"32",
		X"02",X"02",X"1B",X"1B",X"17",X"3F",X"37",X"26",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"32",X"11",X"11",X"11",X"10",X"00",X"00",X"00",
		X"2E",X"0C",X"0C",X"0C",X"48",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"77",X"88",X"88",X"77",X"00",X"06",
		X"EE",X"00",X"EE",X"11",X"11",X"EE",X"00",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"68",X"14",X"00",X"46",X"99",X"99",X"74",
		X"F1",X"49",X"C7",X"00",X"EE",X"11",X"11",X"E2",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
