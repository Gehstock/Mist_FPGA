library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity journey_bg_bits_2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of journey_bg_bits_2 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"AA",X"42",X"AA",X"52",X"AA",X"52",X"AA",X"54",X"AA",X"00",X"2A",X"00",X"2A",X"AA",X"2A",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"2A",X"AA",X"2A",X"AA",X"0A",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"56",X"AA",X"56",X"AA",X"5A",X"AA",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"5A",X"55",X"5A",X"55",X"6A",X"55",X"6A",X"55",X"AA",
		X"80",X"0A",X"A0",X"0A",X"A8",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"82",X"0A",X"82",X"0A",X"82",X"0A",X"82",X"0A",X"82",X"0A",X"82",X"0A",X"82",X"0A",X"82",X"0A",
		X"A8",X"2A",X"A0",X"2A",X"A0",X"0A",X"80",X"0A",X"82",X"0A",X"82",X"0A",X"82",X"0A",X"82",X"0A",
		X"C5",X"55",X"C5",X"55",X"C5",X"55",X"C5",X"55",X"C5",X"54",X"05",X"40",X"05",X"00",X"00",X"2A",
		X"05",X"4A",X"05",X"42",X"C5",X"42",X"C5",X"50",X"C5",X"50",X"C5",X"54",X"C5",X"54",X"C5",X"55",
		X"0A",X"AA",X"02",X"AA",X"02",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"2A",X"05",X"2A",X"05",X"0A",
		X"5A",X"AA",X"6A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"0A",X"AA",
		X"D5",X"AA",X"D5",X"AA",X"D6",X"AA",X"5A",X"AA",X"6A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",
		X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"56",X"D5",X"5A",X"D5",X"6A",
		X"F6",X"6A",X"F6",X"A5",X"F6",X"55",X"F5",X"55",X"F5",X"55",X"F5",X"55",X"F5",X"55",X"F5",X"55",
		X"F6",X"66",X"F6",X"66",X"F6",X"66",X"F6",X"66",X"F6",X"66",X"F6",X"66",X"F6",X"6A",X"F6",X"6A",
		X"00",X"4F",X"01",X"43",X"35",X"43",X"D6",X"43",X"95",X"40",X"55",X"60",X"55",X"A8",X"5A",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"03",X"00",X"03",X"00",X"0F",X"00",X"0F",
		X"AA",X"00",X"8A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"2A",X"00",X"58",X"00",X"58",X"00",
		X"0B",X"55",X"AA",X"D5",X"AA",X"00",X"56",X"00",X"56",X"00",X"56",X"00",X"5A",X"00",X"6A",X"00",
		X"05",X"57",X"05",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"01",X"55",
		X"5F",X"FF",X"57",X"FF",X"57",X"FF",X"55",X"FF",X"55",X"7F",X"15",X"7F",X"15",X"5F",X"05",X"5F",
		X"FF",X"FE",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"7F",X"FF",X"5F",X"FF",
		X"65",X"96",X"E5",X"96",X"F5",X"96",X"FD",X"96",X"FF",X"96",X"FF",X"D6",X"FF",X"D6",X"FF",X"F6",
		X"65",X"96",X"65",X"96",X"65",X"96",X"65",X"96",X"65",X"96",X"65",X"96",X"65",X"96",X"65",X"96",
		X"55",X"55",X"55",X"55",X"15",X"55",X"00",X"25",X"00",X"A2",X"AA",X"A6",X"AA",X"96",X"6A",X"96",
		X"56",X"C0",X"95",X"F0",X"95",X"7C",X"95",X"6F",X"A5",X"56",X"E9",X"55",X"FD",X"55",X"FF",X"D5",
		X"05",X"00",X"14",X"00",X"50",X"00",X"50",X"55",X"51",X"55",X"55",X"BC",X"55",X"F0",X"55",X"C0",
		X"55",X"55",X"55",X"56",X"55",X"5A",X"56",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"55",X"01",X"55",
		X"00",X"00",X"00",X"00",X"A0",X"0A",X"AA",X"AA",X"A5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"00",X"54",X"00",X"50",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"01",X"00",X"55",X"00",X"55",X"01",X"50",X"05",X"50",X"15",X"40",X"55",X"40",
		X"01",X"5F",X"01",X"57",X"00",X"57",X"00",X"55",X"00",X"15",X"00",X"15",X"00",X"05",X"00",X"05",
		X"57",X"FF",X"57",X"FF",X"57",X"FF",X"56",X"FF",X"55",X"FF",X"15",X"7F",X"05",X"7F",X"05",X"6F",
		X"FF",X"59",X"FF",X"59",X"FF",X"D9",X"FF",X"D9",X"7F",X"F9",X"7F",X"FD",X"6F",X"FD",X"5F",X"FF",
		X"96",X"A1",X"D6",X"A0",X"D6",X"A0",X"F6",X"A8",X"F6",X"6A",X"FE",X"5A",X"FE",X"5A",X"FE",X"59",
		X"FF",X"FF",X"55",X"56",X"55",X"5A",X"55",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"5F",X"AA",X"5F",X"AA",X"5F",X"AA",X"5A",X"AA",X"A9",X"56",X"55",X"FF",X"57",X"FF",X"7F",X"FF",
		X"55",X"54",X"55",X"55",X"55",X"55",X"5F",X"55",X"5F",X"D5",X"5F",X"FD",X"5F",X"FF",X"5F",X"EA",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"AA",X"AA",X"00",X"00",X"15",X"40",X"55",X"50",
		X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",X"02",X"AA",X"AA",X"A5",X"A5",X"55",X"55",X"55",
		X"00",X"05",X"00",X"15",X"00",X"55",X"05",X"55",X"15",X"55",X"55",X"55",X"55",X"40",X"54",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"55",X"50",
		X"55",X"57",X"55",X"57",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"FF",X"55",X"FF",X"55",X"7F",X"55",X"7F",X"55",X"7F",X"55",X"6F",X"55",X"5F",X"55",X"5F",
		X"FF",X"57",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"05",X"55",X"14",X"01",X"10",X"01",X"10",X"01",X"10",X"01",X"11",X"55",X"11",X"55",X"00",X"00",
		X"00",X"00",X"00",X"01",X"15",X"55",X"15",X"55",X"10",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"41",X"11",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"55",X"10",X"55",X"00",X"00",
		X"11",X"55",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"01",X"10",X"05",X"10",X"05",X"00",X"00",
		X"00",X"40",X"15",X"55",X"00",X"40",X"00",X"40",X"00",X"40",X"05",X"40",X"05",X"40",X"00",X"00",
		X"10",X"55",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"11",X"45",X"11",X"45",X"00",X"00",
		X"10",X"55",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"11",X"55",X"11",X"55",X"00",X"00",
		X"14",X"00",X"11",X"00",X"11",X"40",X"10",X"55",X"10",X"15",X"10",X"00",X"10",X"00",X"00",X"00",
		X"15",X"55",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"11",X"55",X"11",X"55",X"00",X"00",
		X"15",X"55",X"15",X"55",X"10",X"40",X"10",X"40",X"10",X"40",X"10",X"40",X"11",X"40",X"00",X"00",
		X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",X"FF",X"F9",X"FF",X"D5",
		X"FA",X"95",X"F9",X"55",X"F5",X"55",X"D5",X"55",X"55",X"56",X"55",X"6A",X"57",X"EA",X"5F",X"EA",
		X"AA",X"99",X"AA",X"A5",X"EA",X"95",X"EA",X"95",X"EA",X"AA",X"FA",X"A0",X"FA",X"A0",X"FA",X"A1",
		X"55",X"55",X"55",X"54",X"55",X"40",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"01",X"55",X"15",X"55",
		X"55",X"40",X"50",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"95",X"55",X"A5",X"55",X"A9",X"55",X"AA",X"95",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"15",X"55",X"15",X"55",X"10",X"40",X"10",X"40",X"10",X"40",X"11",X"55",X"11",X"55",X"00",X"00",
		X"15",X"15",X"11",X"51",X"10",X"41",X"10",X"41",X"10",X"41",X"11",X"55",X"11",X"55",X"00",X"00",
		X"10",X"05",X"10",X"05",X"10",X"05",X"10",X"05",X"10",X"05",X"11",X"55",X"11",X"54",X"00",X"00",
		X"05",X"54",X"14",X"05",X"10",X"01",X"10",X"01",X"10",X"01",X"11",X"55",X"11",X"55",X"00",X"00",
		X"10",X"01",X"10",X"01",X"10",X"41",X"10",X"41",X"10",X"41",X"11",X"55",X"11",X"55",X"00",X"00",
		X"10",X"00",X"10",X"00",X"10",X"40",X"10",X"40",X"10",X"40",X"11",X"55",X"11",X"55",X"00",X"00",
		X"10",X"55",X"10",X"41",X"10",X"41",X"10",X"01",X"10",X"01",X"11",X"55",X"11",X"54",X"00",X"00",
		X"15",X"55",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"05",X"55",X"05",X"55",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"01",X"15",X"55",X"15",X"55",X"10",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"05",X"55",X"05",X"55",X"00",X"01",X"00",X"01",X"00",X"05",X"00",X"05",X"00",X"00",
		X"14",X"01",X"05",X"05",X"01",X"54",X"00",X"50",X"00",X"10",X"05",X"55",X"05",X"55",X"00",X"00",
		X"00",X"05",X"00",X"05",X"00",X"01",X"00",X"01",X"00",X"01",X"05",X"55",X"05",X"55",X"00",X"00",
		X"15",X"55",X"05",X"00",X"01",X"50",X"01",X"50",X"05",X"00",X"15",X"55",X"15",X"55",X"00",X"00",
		X"15",X"55",X"00",X"15",X"01",X"50",X"15",X"00",X"10",X"00",X"11",X"55",X"11",X"55",X"00",X"00",
		X"15",X"55",X"10",X"01",X"10",X"01",X"10",X"01",X"10",X"01",X"11",X"55",X"11",X"55",X"00",X"00",
		X"15",X"40",X"10",X"40",X"10",X"40",X"10",X"40",X"10",X"40",X"11",X"55",X"11",X"55",X"00",X"00",
		X"15",X"55",X"10",X"14",X"10",X"15",X"10",X"01",X"10",X"01",X"11",X"55",X"11",X"55",X"00",X"00",
		X"15",X"45",X"10",X"55",X"10",X"50",X"10",X"40",X"10",X"40",X"11",X"55",X"11",X"55",X"00",X"00",
		X"10",X"55",X"10",X"55",X"10",X"41",X"10",X"41",X"10",X"41",X"11",X"45",X"11",X"45",X"00",X"00",
		X"00",X"00",X"10",X"00",X"10",X"00",X"15",X"55",X"15",X"55",X"10",X"00",X"10",X"00",X"00",X"00",
		X"15",X"55",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"05",X"55",X"05",X"55",X"00",X"00",
		X"15",X"50",X"00",X"14",X"00",X"05",X"00",X"15",X"00",X"54",X"05",X"50",X"05",X"40",X"00",X"00",
		X"15",X"55",X"00",X"14",X"01",X"50",X"01",X"50",X"00",X"14",X"05",X"55",X"05",X"55",X"00",X"00",
		X"14",X"05",X"05",X"14",X"01",X"50",X"00",X"40",X"01",X"50",X"05",X"14",X"00",X"05",X"00",X"00",
		X"14",X"00",X"05",X"00",X"01",X"40",X"00",X"55",X"01",X"55",X"05",X"40",X"05",X"00",X"00",X"00",
		X"10",X"01",X"11",X"01",X"11",X"41",X"10",X"41",X"10",X"51",X"10",X"15",X"10",X"05",X"00",X"00",
		X"FD",X"55",X"F5",X"5F",X"D5",X"7F",X"55",X"5F",X"55",X"5F",X"65",X"7F",X"A5",X"7F",X"95",X"5F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F5",X"FF",X"D5",X"FF",X"55",
		X"00",X"AA",X"AA",X"AA",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"15",X"05",X"55",X"55",X"55",X"55",X"55",X"55",X"40",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"40",X"50",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"15",X"40",X"15",X"54",X"15",
		X"55",X"56",X"00",X"16",X"00",X"1A",X"01",X"5A",X"55",X"AA",X"56",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"57",X"FF",X"55",X"FF",X"55",X"7F",X"55",X"5F",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",
		X"00",X"00",X"00",X"02",X"02",X"AA",X"AA",X"AB",X"AB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"54",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"50",X"00",X"00",
		X"75",X"55",X"75",X"55",X"75",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"55",X"55",X"55",X"55",
		X"D5",X"55",X"D5",X"55",X"F5",X"55",X"75",X"55",X"75",X"55",X"75",X"55",X"75",X"55",X"75",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"55",X"55",X"55",
		X"95",X"00",X"A5",X"40",X"A9",X"55",X"AA",X"55",X"AA",X"95",X"AA",X"A5",X"AA",X"AA",X"AA",X"AA",
		X"55",X"55",X"55",X"55",X"15",X"55",X"05",X"55",X"01",X"55",X"40",X"55",X"50",X"15",X"94",X"05",
		X"0F",X"FF",X"3F",X"FF",X"3F",X"FF",X"57",X"FF",X"55",X"FF",X"55",X"5F",X"55",X"57",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"2A",X"AA",X"AA",X"AA",X"AA",X"AF",X"AF",X"FF",X"5F",X"FF",
		X"01",X"54",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"5F",X"FF",X"57",X"FD",X"55",X"F5",X"55",X"55",X"55",X"55",X"15",X"55",X"15",X"55",X"05",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"F5",X"5F",X"7F",X"FF",X"7F",X"FF",
		X"55",X"5F",X"55",X"57",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"55",X"57",X"55",
		X"00",X"55",X"01",X"55",X"05",X"55",X"15",X"D5",X"57",X"F5",X"5F",X"FD",X"5F",X"FF",X"7F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"15",
		X"02",X"A9",X"2A",X"55",X"A9",X"41",X"A5",X"01",X"A4",X"01",X"94",X"00",X"54",X"00",X"55",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",
		X"40",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"05",
		X"54",X"05",X"54",X"05",X"54",X"15",X"50",X"15",X"50",X"15",X"50",X"15",X"40",X"15",X"40",X"15",
		X"55",X"50",X"55",X"50",X"55",X"40",X"55",X"40",X"55",X"40",X"55",X"40",X"55",X"01",X"55",X"01",
		X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",
		X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"2A",X"0A",X"AA",X"2A",X"AA",X"AA",X"80",X"00",X"0A",
		X"40",X"00",X"40",X"00",X"54",X"00",X"55",X"00",X"55",X"40",X"55",X"50",X"55",X"55",X"55",X"55",
		X"55",X"40",X"55",X"00",X"54",X"00",X"50",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"55",X"54",X"55",X"50",X"55",X"50",X"55",X"40",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"AA",X"A0",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"0A",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"00",X"54",X"00",X"54",X"00",X"55",X"00",X"55",X"40",X"55",X"50",X"55",X"54",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"55",X"50",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"05",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"5F",X"55",X"57",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A8",X"00",X"AA",X"80",
		X"05",X"55",X"00",X"55",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"80",X"00",X"A0",X"00",X"AA",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"55",X"55",X"55",X"55",X"15",X"55",X"01",X"55",X"00",X"55",X"00",X"15",X"00",X"05",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"A8",X"00",X"AA",X"00",X"AA",X"80",
		X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"55",X"05",X"55",X"01",X"55",X"00",X"55",X"00",X"15",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"80",X"AA",X"A0",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"A0",X"00",X"A0",X"00",X"AA",X"00",X"AA",X"80",
		X"15",X"55",X"15",X"55",X"05",X"55",X"05",X"55",X"01",X"55",X"00",X"55",X"00",X"55",X"00",X"15",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"A8",X"00",X"A8",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"80",X"AA",X"80",X"AA",X"A0",X"AA",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"A0",X"00",
		X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",
		X"00",X"55",X"00",X"55",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",
		X"01",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",
		X"05",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"01",X"55",
		X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",
		X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"80",X"AA",X"80",
		X"A8",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"00",
		X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"15",X"54",X"50",X"05",X"44",X"11",X"44",X"11",X"44",X"11",X"45",X"51",X"50",X"05",X"15",X"54",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"D5",X"55",X"B5",X"55",X"AD",X"55",X"B5",X"55",X"AF",X"55",X"AA",X"D5",X"AA",X"BF",
		X"55",X"57",X"55",X"5E",X"55",X"7A",X"55",X"5E",X"57",X"DE",X"5E",X"BA",X"7A",X"A2",X"EA",X"AA",
		X"AA",X"AA",X"5A",X"AA",X"55",X"AA",X"55",X"6A",X"55",X"5A",X"55",X"56",X"55",X"56",X"55",X"55",
		X"EA",X"FB",X"BB",X"AE",X"AE",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AB",X"AA",X"AE",X"AA",X"BA",X"AA",X"EA",X"AA",X"BA",X"AA",X"BA",X"AB",X"EA",X"BE",X"AA",
		X"EA",X"AA",X"BA",X"AA",X"AE",X"AA",X"AB",X"AA",X"AE",X"AA",X"BA",X"AA",X"EA",X"AA",X"EA",X"AA",
		X"EA",X"AA",X"AE",X"AA",X"AB",X"AA",X"AE",X"AA",X"BA",X"AA",X"EA",X"AA",X"BA",X"AA",X"BA",X"AA",
		X"EA",X"AA",X"BA",X"AA",X"AA",X"AA",X"AE",X"AA",X"AB",X"AA",X"AA",X"EA",X"AA",X"AE",X"AA",X"AB",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"90",X"AA",X"40",X"AA",X"40",X"A9",X"00",X"A4",X"00",X"90",X"00",X"40",X"00",X"40",X"00",
		X"A9",X"00",X"A9",X"00",X"A9",X"00",X"A9",X"00",X"A9",X"00",X"A9",X"00",X"A9",X"00",X"A9",X"00",
		X"AA",X"40",X"AA",X"40",X"AA",X"40",X"AA",X"40",X"A9",X"00",X"A9",X"00",X"A9",X"00",X"A9",X"00",
		X"AA",X"A4",X"AA",X"A4",X"AA",X"A4",X"AA",X"A4",X"AA",X"A4",X"AA",X"A4",X"AA",X"90",X"AA",X"90",
		X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",
		X"AA",X"A4",X"AA",X"A4",X"AA",X"A9",X"AA",X"A9",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"A4",X"AA",X"A4",X"AA",X"90",X"AA",X"90",X"AA",X"90",X"AA",X"90",X"AA",X"90",X"AA",X"A4",
		X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",X"A4",X"AA",X"A4",X"AA",X"A4",X"AA",X"A4",
		X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"A9",X"00",X"AA",X"40",X"AA",X"40",X"AA",X"90",X"AA",X"90",X"AA",X"A4",X"AA",X"A4",X"AA",X"A9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"90",X"00",X"A4",X"00",
		X"AA",X"90",X"AA",X"90",X"AA",X"90",X"AA",X"90",X"AA",X"90",X"AA",X"90",X"AA",X"90",X"AA",X"90",
		X"A4",X"00",X"A4",X"00",X"A4",X"00",X"A9",X"00",X"A9",X"00",X"A9",X"00",X"A9",X"00",X"A9",X"00",
		X"A9",X"00",X"A4",X"00",X"A4",X"00",X"90",X"00",X"90",X"00",X"A4",X"00",X"A4",X"00",X"A4",X"00",
		X"AA",X"90",X"AA",X"90",X"AA",X"90",X"AA",X"90",X"AA",X"90",X"AA",X"90",X"AA",X"90",X"AA",X"90",
		X"AA",X"A4",X"AA",X"A4",X"AA",X"A4",X"AA",X"A4",X"AA",X"A4",X"AA",X"A4",X"AA",X"A4",X"AA",X"A4",
		X"A4",X"00",X"A4",X"00",X"A4",X"00",X"A9",X"00",X"A9",X"00",X"A9",X"00",X"AA",X"40",X"AA",X"90",
		X"AA",X"A4",X"AA",X"A4",X"AA",X"A4",X"AA",X"A4",X"AA",X"90",X"AA",X"90",X"AA",X"40",X"AA",X"40",
		X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"E0",X"00",X"E0",X"00",X"F0",X"00",X"B0",X"00",
		X"B8",X"00",X"B8",X"00",X"B8",X"00",X"BE",X"00",X"AE",X"00",X"AE",X"00",X"AF",X"80",X"AB",X"80",
		X"AB",X"A0",X"AB",X"A0",X"AB",X"E0",X"AA",X"E8",X"AA",X"FA",X"AA",X"BA",X"AA",X"BE",X"AA",X"AE",
		X"AA",X"AF",X"AA",X"AB",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"05",X"00",X"01",X"04",X"05",X"40",X"01",X"40",X"01",X"51",X"01",X"10",X"01",X"55",
		X"00",X"55",X"00",X"44",X"01",X"17",X"00",X"01",X"00",X"05",X"00",X"01",X"00",X"10",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",
		X"A0",X"00",X"E0",X"00",X"FA",X"00",X"BA",X"80",X"BE",X"A0",X"AF",X"A8",X"AB",X"EA",X"AA",X"FA",
		X"40",X"00",X"40",X"01",X"50",X"40",X"55",X"05",X"11",X"45",X"45",X"50",X"54",X"55",X"54",X"D1",
		X"45",X"54",X"55",X"05",X"04",X"45",X"00",X"51",X"04",X"00",X"00",X"04",X"00",X"00",X"00",X"00",
		X"01",X"DF",X"00",X"77",X"01",X"1D",X"01",X"47",X"00",X"11",X"00",X"44",X"00",X"00",X"00",X"43",
		X"11",X"55",X"05",X"51",X"51",X"14",X"55",X"74",X"C5",X"10",X"54",X"54",X"45",X"40",X"4C",X"50",
		X"55",X"50",X"54",X"40",X"04",X"00",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"BE",X"AA",X"AF",X"AA",X"AB",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"00",X"AA",X"A8",X"FA",X"AA",X"BE",X"AA",X"AF",X"EA",X"AA",X"FF",X"AA",X"AB",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"A8",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FF",X"AA",X"AF",X"FF",
		X"A8",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"AA",X"A0",X"AA",X"80",X"AA",X"80",X"AA",X"00",X"AA",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"A0",
		X"AA",X"00",X"A8",X"00",X"A0",X"00",X"80",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"A0",X"AA",X"80",
		X"AA",X"AA",X"AA",X"A0",X"AA",X"00",X"A0",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"00",X"03",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00",X"0C",X"00",X"0C",X"00",X"0C",
		X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"30",
		X"0C",X"30",X"0C",X"30",X"03",X"30",X"03",X"C0",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",
		X"30",X"03",X"30",X"03",X"30",X"C3",X"30",X"0C",X"33",X"0C",X"30",X"0C",X"30",X"0C",X"0C",X"30",
		X"30",X"00",X"30",X"00",X"30",X"C0",X"30",X"00",X"33",X"00",X"30",X"00",X"30",X"00",X"30",X"00",
		X"03",X"00",X"0C",X"00",X"0C",X"30",X"0C",X"00",X"0C",X"C0",X"0C",X"00",X"0C",X"00",X"30",X"00",
		X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"03",X"30",X"03",X"00",X"03",X"00",X"03",X"00",
		X"00",X"03",X"00",X"03",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"30",X"00",X"30",X"00",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"30",X"00",X"0F",X"00",X"00",X"FF",X"00",X"00",
		X"30",X"03",X"C0",X"00",X"CC",X"00",X"C0",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C3",X"00",X"C3",X"03",X"03",X"03",X"03",X"03",X"03",X"0C",X"03",X"0C",X"03",X"0C",X"03",
		X"0C",X"00",X"0C",X"03",X"30",X"03",X"30",X"03",X"30",X"0F",X"30",X"0F",X"C0",X"33",X"C0",X"33",
		X"00",X"03",X"00",X"0F",X"0C",X"33",X"00",X"33",X"30",X"C3",X"00",X"C3",X"03",X"03",X"03",X"03",
		X"0C",X"00",X"0C",X"00",X"30",X"30",X"30",X"00",X"C3",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",
		X"00",X"0C",X"00",X"30",X"00",X"30",X"00",X"C0",X"00",X"C0",X"03",X"30",X"03",X"00",X"0C",X"00",
		X"03",X"00",X"0C",X"00",X"30",X"00",X"30",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"0C",X"03",X"00",X"0C",X"30",X"30",X"00",X"30",X"00",X"C0",X"00",X"C0",
		X"00",X"3F",X"00",X"3F",X"0C",X"3F",X"00",X"0F",X"30",X"0F",X"00",X"0F",X"00",X"03",X"00",X"03",
		X"00",X"FF",X"00",X"FF",X"0C",X"FF",X"00",X"FF",X"30",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"0D",X"FF",X"0D",X"FF",X"0D",X"FF",X"03",X"FF",X"33",X"FF",X"03",X"FF",X"03",X"FF",X"03",X"FF",
		X"F5",X"FF",X"F5",X"FF",X"FD",X"FF",X"F5",X"FF",X"F5",X"FF",X"3D",X"FF",X"3D",X"FF",X"0D",X"FF",
		X"D5",X"FF",X"D5",X"FF",X"FD",X"FF",X"F5",X"FF",X"F5",X"FF",X"F5",X"FF",X"F5",X"FF",X"F5",X"FF",
		X"F5",X"7F",X"F5",X"7F",X"FD",X"7F",X"D5",X"7F",X"F5",X"7F",X"D5",X"FF",X"D5",X"FF",X"D5",X"FF",
		X"FC",X"D7",X"FF",X"5F",X"FF",X"5F",X"FD",X"5F",X"FD",X"5F",X"FD",X"5F",X"F5",X"5F",X"F5",X"5F",
		X"FF",X"1A",X"FC",X"09",X"FC",X"0A",X"FC",X"05",X"3C",X"01",X"FC",X"01",X"FC",X"0F",X"FC",X"37",
		X"F5",X"55",X"FD",X"55",X"FD",X"55",X"FD",X"55",X"FD",X"55",X"FD",X"55",X"FD",X"55",X"FD",X"D6",
		X"3F",X"55",X"3D",X"55",X"3D",X"55",X"35",X"55",X"35",X"55",X"D5",X"55",X"D5",X"55",X"F5",X"55",
		X"03",X"FD",X"03",X"F5",X"0F",X"F5",X"0F",X"F5",X"3F",X"D5",X"0F",X"D5",X"0F",X"D5",X"3F",X"55",
		X"03",X"0F",X"0C",X"3F",X"0C",X"3F",X"30",X"3F",X"30",X"FF",X"C3",X"FF",X"C0",X"FF",X"00",X"FD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",X"00",X"0F",X"00",X"3F",X"00",X"CF",
		X"00",X"FF",X"00",X"3F",X"00",X"3F",X"00",X"0F",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"3F",X"FF",X"3F",X"FF",X"0F",X"FF",X"0F",X"FF",X"03",X"FF",X"00",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"15",X"FF",X"15",X"FF",X"55",X"FF",X"D5",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"94",X"00",X"90",X"00",X"90",X"00",X"7C",X"00",X"FC",X"01",X"FC",X"01",X"FF",X"05",X"FF",X"05",
		X"55",X"AA",X"55",X"AA",X"55",X"6A",X"55",X"4A",X"A9",X"4A",X"99",X"42",X"A9",X"02",X"A4",X"00",
		X"56",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"56",X"AA",X"56",X"AA",
		X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"56",X"AA",X"56",X"AA",X"56",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"AA",X"5A",X"AA",X"5A",X"AA",
		X"00",X"AA",X"00",X"AA",X"02",X"AA",X"02",X"AA",X"0A",X"AA",X"0A",X"AA",X"2A",X"AA",X"2A",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"0A",X"00",X"0A",X"00",X"2A",X"00",X"2A",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"FC",X"0F",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"D5",X"FF",X"D5",X"FF",X"D5",X"FF",X"F5",X"FF",X"F5",X"FF",X"F5",X"FF",X"FD",X"FF",X"FF",
		X"55",X"6A",X"55",X"5A",X"55",X"56",X"F5",X"56",X"FD",X"55",X"FD",X"55",X"FF",X"55",X"FF",X"55",
		X"AA",X"AA",X"2A",X"AA",X"2A",X"AA",X"5A",X"AA",X"56",X"AA",X"56",X"AA",X"55",X"AA",X"55",X"6A",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"02",X"AA",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"0A",X"00",X"2A",X"00",X"AA",
		X"FE",X"A0",X"FE",X"A0",X"FE",X"80",X"FA",X"00",X"E8",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",X"FF",X"AA",X"FF",X"A8",
		X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",
		X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F7",X"D7",X"FF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"5D",X"5D",X"5D",X"7D",X"5D",X"7D",X"5D",X"75",X"5D",X"F5",X"5D",X"F5",X"7D",X"F5",X"75",X"D7",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"6A",X"AA",X"56",X"AA",X"57",X"6A",
		X"00",X"AA",X"02",X"AA",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"2A",
		X"FC",X"00",X"F8",X"00",X"F0",X"00",X"E0",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"FA",X"AA",X"EA",X"AB",X"EA",X"AB",X"E8",X"AF",X"88",X"AF",X"00",X"BE",X"00",X"BC",X"00",
		X"AA",X"BF",X"AA",X"BF",X"AA",X"BF",X"AA",X"FE",X"AA",X"FE",X"AA",X"FE",X"AA",X"FA",X"AA",X"FA",
		X"EA",X"AB",X"EA",X"AB",X"EA",X"AF",X"AA",X"AF",X"AA",X"AF",X"AA",X"AF",X"AA",X"BF",X"AA",X"BF",
		X"FF",X"EA",X"FF",X"EA",X"FF",X"AA",X"FF",X"AA",X"FE",X"AA",X"FE",X"AA",X"FA",X"AA",X"FA",X"AB",
		X"5F",X"7F",X"7D",X"7D",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FA",X"FF",X"EA",X"FF",X"EA",
		X"55",X"6A",X"75",X"FA",X"75",X"F7",X"F5",X"D7",X"F7",X"D7",X"D7",X"D7",X"D7",X"5F",X"D7",X"5F",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AB",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"BF",X"AA",X"BF",X"AA",X"BF",X"AA",X"BF",X"AA",X"BF",X"AA",X"FF",X"AA",X"AB",X"AA",X"AB",
		X"AA",X"FF",X"AA",X"FF",X"AA",X"BF",X"AA",X"BF",X"AA",X"BF",X"AA",X"BF",X"AA",X"BF",X"AA",X"BF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"03",X"FE",X"BF",X"FE",X"AB",X"FE",
		X"01",X"55",X"01",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AE",X"FE",X"8F",X"FA",X"03",X"FA",X"03",X"FA",X"00",X"FA",X"00",X"FD",X"00",X"5F",X"00",X"55",
		X"FF",X"BF",X"FF",X"BF",X"FE",X"BF",X"FE",X"FF",X"FE",X"FE",X"BE",X"FE",X"BE",X"FE",X"AE",X"FE",
		X"FE",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",
		X"BF",X"FE",X"BF",X"FE",X"BF",X"FE",X"FF",X"FE",X"FF",X"FF",X"FA",X"FF",X"FA",X"FF",X"FE",X"FF",
		X"55",X"A0",X"5A",X"A0",X"AA",X"80",X"AA",X"E8",X"AB",X"E8",X"AB",X"F8",X"AF",X"FA",X"AF",X"FA",
		X"BF",X"A5",X"AF",X"55",X"ED",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"55",X"55",X"55",X"59",
		X"FE",X"AA",X"FE",X"AA",X"FE",X"AA",X"FE",X"AA",X"FE",X"AA",X"FE",X"AA",X"FE",X"AA",X"FE",X"AA",
		X"FE",X"AA",X"BE",X"AA",X"AA",X"AA",X"BE",X"AA",X"BF",X"AA",X"BF",X"AA",X"FF",X"AA",X"FE",X"AA",
		X"FF",X"F6",X"FE",X"56",X"FE",X"6A",X"FE",X"AA",X"FE",X"AA",X"FE",X"AA",X"FA",X"AA",X"FA",X"AA",
		X"BF",X"F6",X"BF",X"F6",X"BF",X"F6",X"BF",X"F6",X"BF",X"F6",X"FF",X"F6",X"FF",X"F6",X"FF",X"F6",
		X"AF",X"F6",X"AF",X"F6",X"BF",X"F6",X"BF",X"F6",X"BF",X"F6",X"BF",X"F6",X"BF",X"F6",X"BF",X"F6",
		X"AF",X"FA",X"AF",X"FA",X"AF",X"FA",X"AF",X"FA",X"AF",X"EA",X"AF",X"F6",X"AF",X"F6",X"AF",X"F6",
		X"FF",X"DA",X"FF",X"DA",X"FF",X"DA",X"BF",X"EA",X"BF",X"FA",X"AF",X"FA",X"AF",X"FA",X"AF",X"FA",
		X"FF",X"6A",X"FF",X"5A",X"FF",X"DA",X"FF",X"DA",X"FF",X"DA",X"FF",X"DA",X"FF",X"DA",X"FF",X"DA",
		X"AA",X"95",X"AA",X"95",X"EA",X"A5",X"D6",X"A5",X"F5",X"A9",X"FD",X"A9",X"FD",X"69",X"FF",X"69",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"A0",X"15",X"A5",X"55",X"A5",X"55",X"A9",X"55",
		X"54",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"95",X"00",X"54",X"00",X"54",X"00",X"54",X"00",X"5C",X"00",X"7C",X"00",X"F4",X"00",X"54",X"00",
		X"95",X"00",X"95",X"00",X"95",X"00",X"95",X"00",X"95",X"00",X"95",X"00",X"95",X"00",X"95",X"00",
		X"95",X"00",X"A5",X"00",X"E5",X"00",X"E5",X"00",X"E5",X"00",X"E5",X"00",X"E5",X"00",X"A5",X"00",
		X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"90",X"00",X"94",X"00",X"95",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"FF",X"AA",X"FE",X"A8",X"3E",X"A0",X"3F",X"A0",X"0F",X"80",X"0F",X"80",X"03",X"00",X"00",
		X"5F",X"EF",X"5F",X"EF",X"6B",X"AF",X"6B",X"AF",X"6B",X"BF",X"6B",X"BF",X"AB",X"BF",X"AB",X"FF",
		X"97",X"AF",X"97",X"EF",X"97",X"EF",X"97",X"EF",X"5F",X"EF",X"5F",X"EF",X"5F",X"EF",X"5F",X"EF",
		X"A5",X"7B",X"A5",X"7A",X"A5",X"7E",X"A5",X"FE",X"95",X"FE",X"95",X"FF",X"95",X"FF",X"96",X"BF",
		X"A9",X"55",X"A9",X"55",X"A9",X"54",X"A9",X"54",X"A9",X"50",X"A9",X"5C",X"A5",X"5F",X"A5",X"5B",
		X"AA",X"55",X"AA",X"55",X"AA",X"55",X"A9",X"55",X"A9",X"55",X"A9",X"55",X"A9",X"55",X"A9",X"55",
		X"AA",X"50",X"AA",X"50",X"AA",X"50",X"AA",X"50",X"AA",X"54",X"AA",X"54",X"AA",X"54",X"AA",X"55",
		X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"50",X"AA",X"40",X"AA",X"40",
		X"A4",X"04",X"A5",X"00",X"A9",X"00",X"A9",X"40",X"A9",X"41",X"AA",X"55",X"AA",X"55",X"AA",X"55",
		X"55",X"00",X"54",X"01",X"54",X"04",X"51",X"44",X"51",X"54",X"90",X"54",X"90",X"54",X"A4",X"14",
		X"55",X"50",X"55",X"40",X"55",X"40",X"55",X"40",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"50",X"00",
		X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BD",X"54",X"BD",X"54",X"FD",X"50",X"F5",X"40",X"F5",X"40",X"D5",X"00",X"D5",X"00",X"D5",X"00",
		X"EF",X"54",X"EF",X"54",X"EF",X"54",X"EF",X"54",X"AD",X"54",X"BD",X"54",X"BD",X"54",X"BD",X"54",
		X"AF",X"00",X"EF",X"00",X"EF",X"00",X"EF",X"00",X"EF",X"00",X"EF",X"00",X"EF",X"00",X"EF",X"40",
		X"F0",X"00",X"F0",X"00",X"F0",X"00",X"FC",X"00",X"BC",X"00",X"BC",X"00",X"BC",X"00",X"BF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",
		X"14",X"00",X"54",X"00",X"50",X"00",X"50",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"00",X"00",
		X"00",X"10",X"00",X"40",X"00",X"40",X"01",X"40",X"01",X"00",X"05",X"00",X"05",X"00",X"14",X"00",
		X"01",X"00",X"04",X"00",X"54",X"00",X"54",X"00",X"54",X"00",X"54",X"00",X"54",X"10",X"10",X"10",
		X"00",X"00",X"10",X"00",X"10",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"2A",X"00",X"0A",X"00",X"0A",X"00",X"02",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"AA",X"0A",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"2A",
		X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"0A",X"AA",X"0A",X"AA",
		X"0A",X"AA",X"02",X"AA",X"02",X"AA",X"00",X"AA",X"00",X"2A",X"00",X"0A",X"00",X"02",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"2A",X"AA",X"2A",X"AA",
		X"2A",X"AA",X"0A",X"AA",X"02",X"AA",X"00",X"2A",X"00",X"0A",X"00",X"02",X"00",X"00",X"00",X"00",
		X"0A",X"AA",X"02",X"AA",X"00",X"AA",X"00",X"2A",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"0A",X"AA",X"00",X"AA",
		X"AA",X"80",X"AA",X"80",X"AA",X"00",X"AA",X"00",X"A8",X"00",X"A0",X"00",X"80",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"A8",X"AA",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"80",X"00",
		X"00",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"AA",X"AA",
		X"02",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",
		X"AA",X"00",X"AA",X"80",X"AA",X"A0",X"AA",X"A8",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"80",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"00",X"AA",X"00",
		X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"82",X"AA",X"00",X"AA",X"00",X"2A",X"00",X"0A",X"00",X"02",X"00",X"00",
		X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"A0",X"00",X"A8",X"00",
		X"02",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"2A",X"00",X"0A",
		X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",
		X"02",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",
		X"A8",X"0A",X"A8",X"0A",X"A8",X"0A",X"A0",X"0A",X"A0",X"0A",X"80",X"2A",X"80",X"2A",X"00",X"AA",
		X"AA",X"80",X"AA",X"80",X"AA",X"00",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"02",
		X"AA",X"02",X"AA",X"02",X"AA",X"02",X"A8",X"02",X"A8",X"02",X"A8",X"0A",X"A0",X"0A",X"A0",X"0A",
		X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"02",X"AA",X"02",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"02",X"AA",X"0A",X"AA",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"A0",X"AA",X"80",X"AA",X"00",
		X"A8",X"00",X"A0",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"00",X"0A",X"00",X"2A",X"00",X"AA",X"02",X"AA",X"0A",X"AA",X"2A",X"AA",
		X"AA",X"00",X"AA",X"00",X"A8",X"00",X"A8",X"00",X"A0",X"00",X"A0",X"00",X"80",X"00",X"00",X"00",
		X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"00",X"AA",X"00",X"AA",X"00",
		X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AE",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"BA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"0A",X"AA",X"0A",X"AA",X"2A",X"AA",X"AA",X"AA",
		X"00",X"2A",X"00",X"2A",X"00",X"2A",X"00",X"2A",X"00",X"2A",X"00",X"AA",X"00",X"AA",X"00",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",
		X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"95",X"55",X"95",X"55",X"A5",X"55",
		X"7F",X"33",X"57",X"CF",X"5F",X"FF",X"6B",X"FF",X"5A",X"AA",X"AA",X"AA",X"56",X"AA",X"55",X"FF",
		X"D5",X"55",X"FD",X"55",X"55",X"55",X"95",X"55",X"A9",X"55",X"95",X"55",X"55",X"56",X"F5",X"56",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"2A",X"AA",X"0A",X"AA",X"0A",X"AA",X"02",X"AA",X"00",X"AA",
		X"A9",X"55",X"AA",X"55",X"AA",X"95",X"AA",X"A5",X"AA",X"A9",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"5F",X"FF",X"7F",X"FF",X"5F",X"FF",X"56",X"AA",X"55",X"AA",X"95",X"69",X"A9",X"59",X"AA",X"AA",
		X"FD",X"56",X"F5",X"5A",X"D5",X"5A",X"55",X"6A",X"55",X"6A",X"56",X"AA",X"6A",X"AA",X"AA",X"AA",
		X"00",X"0A",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"2A",X"AA",X"02",X"AA",X"00",X"2A",X"00",X"0A",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"0A",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"A0",X"00",X"A0",X"00",X"A8",X"00",X"AA",X"00",
		X"AA",X"A0",X"AA",X"A8",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"A8",X"00",X"AA",X"80",X"AA",X"A0",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"0A",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"CA",X"FF",X"F2",X"FF",X"FC",X"FF",X"FC",X"AA",X"FC",X"AA",X"BC",X"AA",X"BC",X"AA",X"BC",
		X"F2",X"AA",X"F2",X"AA",X"F2",X"AA",X"F2",X"AA",X"F2",X"AA",X"F2",X"BF",X"B2",X"BF",X"A2",X"BF",
		X"AF",X"FF",X"BF",X"FF",X"FF",X"FF",X"FC",X"AA",X"F2",X"AA",X"F2",X"AA",X"F2",X"AA",X"F2",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"BF",X"AA",X"BF",X"AA",X"BF",X"AA",X"BF",
		X"F2",X"AA",X"F2",X"AA",X"F2",X"AA",X"F2",X"AA",X"F2",X"BF",X"F2",X"BF",X"F2",X"BF",X"F2",X"BF",
		X"AF",X"CA",X"AF",X"CA",X"AF",X"CA",X"AF",X"CA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",
		X"FA",X"AF",X"FE",X"BF",X"FF",X"FF",X"FF",X"FF",X"AF",X"F2",X"AF",X"CA",X"AF",X"CA",X"AF",X"CA",
		X"FF",X"FF",X"FF",X"CA",X"F2",X"AA",X"F2",X"AA",X"F2",X"BF",X"F2",X"BF",X"F2",X"BF",X"F2",X"BF",
		X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"BF",X"AF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AF",X"FF",X"FF",X"FF",X"FF",X"F2",X"FC",X"AA",
		X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"2A",X"CA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"F2",X"AA",X"F2",X"AA",X"F2",X"AA",X"F2",X"AA",X"F2",X"AA",X"F2",X"AA",X"F2",X"AA",X"F2",X"AA",
		X"AF",X"2A",X"AF",X"2A",X"AF",X"2A",X"AF",X"2A",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AF",X"2A",X"AF",X"2A",X"AF",X"2A",X"AF",X"2A",X"AF",X"2A",X"AF",X"2A",X"AF",X"2A",
		X"AA",X"BC",X"AA",X"BC",X"AA",X"BC",X"AA",X"BC",X"AA",X"BC",X"AA",X"BC",X"AA",X"BC",X"AA",X"BC",
		X"02",X"04",X"23",X"14",X"FB",X"50",X"EB",X"40",X"FB",X"50",X"23",X"14",X"02",X"04",X"00",X"00",
		X"FF",X"FF",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",
		X"AA",X"EA",X"AA",X"FA",X"AA",X"BA",X"AA",X"BE",X"AA",X"AE",X"AA",X"AF",X"AA",X"AA",X"AA",X"AA",
		X"AE",X"AA",X"AE",X"AA",X"AE",X"AA",X"AE",X"AA",X"AF",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"EA",
		X"AA",X"FA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"EB",X"EA",X"FF",X"AA",X"AA",X"AA",
		X"AA",X"BA",X"AA",X"BA",X"AA",X"BA",X"AA",X"BA",X"AA",X"BA",X"AA",X"BA",X"AA",X"BA",X"AA",X"BA",
		X"00",X"C0",X"00",X"C0",X"00",X"EA",X"AA",X"FA",X"AA",X"BA",X"AA",X"BA",X"AA",X"FF",X"FF",X"FA",
		X"0C",X"00",X"0F",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"C0",X"00",X"C0",
		X"30",X"04",X"31",X"44",X"31",X"11",X"30",X"10",X"30",X"71",X"30",X"04",X"3C",X"10",X"0C",X"00",
		X"10",X"00",X"01",X"04",X"11",X"10",X"00",X"41",X"C4",X"30",X"C4",X"44",X"C1",X"10",X"F0",X"00",
		X"10",X"0F",X"10",X"43",X"41",X"13",X"04",X"43",X"13",X"13",X"44",X"03",X"01",X"10",X"50",X"00",
		X"00",X"C1",X"10",X"F0",X"00",X"30",X"44",X"30",X"13",X"3C",X"41",X"0C",X"10",X"4C",X"00",X"4C",
		X"4F",X"01",X"0F",X"C0",X"43",X"C4",X"13",X"C0",X"03",X"CC",X"10",X"C1",X"44",X"C4",X"00",X"C0",
		X"00",X"00",X"3C",X"30",X"3C",X"00",X"3C",X"00",X"3F",X"04",X"3F",X"30",X"0F",X"00",X"0F",X"04",
		X"30",X"00",X"31",X"30",X"30",X"00",X"31",X"10",X"30",X"04",X"03",X"10",X"00",X"00",X"00",X"04",
		X"3C",X"00",X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"10",X"31",X"00",X"30",X"00",
		X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",
		X"59",X"AA",X"D5",X"AA",X"B5",X"9A",X"AD",X"56",X"B5",X"56",X"AF",X"55",X"AA",X"D5",X"AA",X"BF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"AA",X"95",X"AA",X"96",X"AA",X"6A",X"AA",
		X"A6",X"97",X"A6",X"5E",X"95",X"7A",X"55",X"5E",X"57",X"DE",X"5E",X"BA",X"7A",X"AA",X"EA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"9A",X"AA",X"96",X"AA",X"66",X"AA",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"F2",X"FF",X"F2",X"FF",X"F2",X"FF",X"F2",X"FF",
		X"AF",X"FF",X"BF",X"FF",X"BC",X"AA",X"FC",X"AA",X"FC",X"AA",X"FC",X"AA",X"FC",X"AA",X"F2",X"AA",
		X"FF",X"FC",X"FF",X"FC",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",
		X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
