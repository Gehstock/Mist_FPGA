library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity rome is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of rome is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"A7",X"32",X"48",X"20",X"FC",X"41",X"18",X"78",X"91",X"C8",X"44",X"4D",X"6F",X"9F",X"67",X"CD",
		X"41",X"18",X"EB",X"3E",X"11",X"21",X"00",X"00",X"E5",X"19",X"D2",X"1E",X"18",X"E3",X"E1",X"F5",
		X"79",X"17",X"4F",X"78",X"17",X"47",X"7D",X"17",X"6F",X"7C",X"17",X"67",X"F1",X"3D",X"C2",X"18",
		X"18",X"AF",X"7C",X"1F",X"57",X"7D",X"1F",X"5F",X"3A",X"48",X"20",X"A7",X"79",X"F0",X"2F",X"3C",
		X"C9",X"7C",X"2F",X"67",X"7D",X"2F",X"6F",X"23",X"C9",X"11",X"4A",X"20",X"1A",X"3D",X"CA",X"66",
		X"18",X"12",X"F6",X"30",X"21",X"29",X"20",X"77",X"11",X"B0",X"3E",X"3E",X"01",X"CD",X"30",X"01",
		X"3E",X"1E",X"32",X"25",X"20",X"C9",X"AF",X"32",X"57",X"20",X"32",X"58",X"20",X"32",X"27",X"20",
		X"CD",X"79",X"18",X"FA",X"60",X"18",X"C3",X"10",X"19",X"21",X"86",X"20",X"11",X"0B",X"00",X"19",
		X"7E",X"A7",X"F8",X"7D",X"FE",X"B2",X"C2",X"7F",X"18",X"C9",X"21",X"55",X"20",X"7E",X"A7",X"11",
		X"5E",X"20",X"C2",X"98",X"18",X"11",X"70",X"20",X"23",X"34",X"4E",X"06",X"00",X"21",X"7C",X"19",
		X"09",X"7E",X"EB",X"56",X"2B",X"5E",X"2B",X"77",X"2B",X"1F",X"3E",X"47",X"DA",X"B0",X"18",X"3D",
		X"B6",X"77",X"21",X"22",X"1A",X"09",X"09",X"7E",X"23",X"66",X"6F",X"E9",X"3E",X"0F",X"32",X"24",
		X"20",X"CD",X"D9",X"11",X"D6",X"04",X"FE",X"25",X"D2",X"CD",X"18",X"C6",X"07",X"57",X"EB",X"22",
		X"4E",X"20",X"EB",X"3A",X"09",X"20",X"E6",X"1C",X"4F",X"06",X"00",X"21",X"2E",X"1E",X"09",X"3E",
		X"04",X"C3",X"30",X"01",X"21",X"C8",X"1D",X"3A",X"55",X"20",X"A7",X"CA",X"F1",X"18",X"21",X"E0",
		X"1D",X"CD",X"82",X"1C",X"3E",X"0A",X"32",X"24",X"20",X"2A",X"4E",X"20",X"EB",X"3E",X"0F",X"C3",
		X"6E",X"1B",X"3E",X"0F",X"32",X"24",X"20",X"2A",X"4E",X"20",X"EB",X"3E",X"10",X"C3",X"6E",X"1B",
		X"AF",X"32",X"23",X"20",X"2A",X"0F",X"20",X"22",X"06",X"20",X"C9",X"2A",X"06",X"20",X"23",X"22",
		X"06",X"20",X"C9",X"AF",X"32",X"57",X"20",X"32",X"58",X"20",X"32",X"27",X"20",X"32",X"25",X"20",
		X"CD",X"79",X"18",X"FA",X"4D",X"19",X"3A",X"06",X"20",X"D6",X"67",X"C2",X"4D",X"19",X"32",X"0A",
		X"20",X"21",X"91",X"1A",X"22",X"06",X"20",X"21",X"F6",X"1D",X"C3",X"87",X"1C",X"3E",X"01",X"32",
		X"08",X"20",X"C9",X"8A",X"1B",X"68",X"1B",X"81",X"1B",X"8B",X"1B",X"9D",X"1B",X"A6",X"1B",X"B2",
		X"1B",X"49",X"12",X"11",X"1C",X"24",X"1C",X"5C",X"1C",X"6F",X"1C",X"2B",X"1D",X"48",X"1D",X"7B",
		X"1C",X"7F",X"1C",X"A0",X"80",X"60",X"30",X"0E",X"74",X"74",X"78",X"78",X"7A",X"B0",X"C0",X"D0",
		X"D1",X"58",X"71",X"8F",X"A8",X"FF",X"80",X"50",X"0E",X"9E",X"5E",X"2E",X"0D",X"2A",X"0C",X"30",
		X"0B",X"38",X"12",X"2A",X"13",X"30",X"14",X"38",X"15",X"00",X"12",X"00",X"11",X"00",X"0F",X"00",
		X"0E",X"00",X"00",X"00",X"15",X"01",X"12",X"01",X"11",X"00",X"0F",X"00",X"0E",X"01",X"00",X"00",
		X"BC",X"15",X"BC",X"15",X"BC",X"15",X"BC",X"15",X"BC",X"15",X"BC",X"15",X"BC",X"15",X"D5",X"15",
		X"C5",X"15",X"C5",X"15",X"C5",X"15",X"C5",X"15",X"C5",X"15",X"C5",X"15",X"C5",X"15",X"61",X"16",
		X"06",X"06",X"1A",X"15",X"06",X"FE",X"1A",X"04",X"06",X"00",X"1A",X"09",X"06",X"FA",X"1A",X"FE",
		X"06",X"04",X"1A",X"11",X"06",X"FC",X"1A",X"02",X"06",X"02",X"1A",X"0E",X"FA",X"06",X"FC",X"15",
		X"FA",X"FE",X"FC",X"04",X"FA",X"00",X"FC",X"09",X"FA",X"FA",X"FC",X"FE",X"FA",X"04",X"FC",X"11",
		X"FA",X"FC",X"FC",X"02",X"FA",X"02",X"FC",X"0E",X"E4",X"0A",X"0B",X"38",X"00",X"0B",X"0C",X"30",
		X"17",X"0B",X"0D",X"2A",X"E4",X"0A",X"14",X"38",X"00",X"0B",X"13",X"30",X"17",X"0B",X"12",X"2A",
		X"08",X"09",X"0A",X"09",X"BC",X"18",X"E4",X"18",X"02",X"19",X"8A",X"1B",X"00",X"00",X"00",X"01",
		X"01",X"00",X"01",X"01",X"01",X"02",X"02",X"01",X"02",X"02",X"02",X"03",X"03",X"02",X"03",X"03",
		X"03",X"04",X"04",X"03",X"04",X"04",X"00",X"02",X"FE",X"00",X"02",X"FE",X"00",X"01",X"FF",X"00",
		X"01",X"FF",X"00",X"00",X"FE",X"02",X"00",X"06",X"FA",X"00",X"FF",X"01",X"00",X"FF",X"01",X"00",
		X"01",X"40",X"03",X"42",X"05",X"44",X"06",X"45",X"07",X"46",X"A8",X"E8",X"AA",X"E8",X"AC",X"E8",
		X"AD",X"E8",X"AE",X"E8",X"05",X"02",X"05",X"06",X"09",X"06",X"01",X"0A",X"19",X"01",X"04",X"17",
		X"05",X"06",X"15",X"07",X"02",X"13",X"03",X"03",X"11",X"02",X"07",X"0F",X"06",X"05",X"01",X"04",
		X"01",X"06",X"01",X"11",X"20",X"06",X"00",X"44",X"20",X"04",X"0A",X"AE",X"1A",X"02",X"0E",X"00",
		X"24",X"03",X"1E",X"00",X"02",X"07",X"00",X"24",X"03",X"1E",X"00",X"05",X"9D",X"1A",X"0E",X"08",
		X"0A",X"02",X"09",X"00",X"28",X"03",X"3C",X"00",X"02",X"11",X"00",X"30",X"03",X"3C",X"00",X"02",
		X"0A",X"00",X"3C",X"03",X"3C",X"00",X"08",X"0A",X"09",X"5F",X"20",X"00",X"10",X"08",X"32",X"80",
		X"09",X"71",X"20",X"00",X"10",X"DE",X"36",X"88",X"04",X"00",X"AE",X"1A",X"06",X"01",X"28",X"20",
		X"03",X"5A",X"00",X"0D",X"05",X"E0",X"1A",X"08",X"0F",X"95",X"1C",X"08",X"10",X"9C",X"1D",X"0B",
		X"11",X"20",X"FB",X"1A",X"02",X"12",X"00",X"2C",X"05",X"FF",X"1A",X"02",X"13",X"00",X"30",X"03",
		X"69",X"00",X"08",X"06",X"01",X"44",X"20",X"0A",X"07",X"09",X"5F",X"20",X"01",X"B0",X"01",X"38",
		X"80",X"0B",X"11",X"20",X"26",X"1B",X"06",X"84",X"5B",X"20",X"06",X"35",X"5C",X"20",X"06",X"1E",
		X"28",X"20",X"06",X"50",X"27",X"20",X"09",X"71",X"20",X"01",X"B0",X"DE",X"34",X"88",X"02",X"0B",
		X"A0",X"34",X"03",X"1E",X"00",X"02",X"0C",X"A0",X"34",X"03",X"0F",X"00",X"02",X"08",X"A0",X"34",
		X"02",X"0D",X"A2",X"3E",X"0B",X"47",X"20",X"52",X"1B",X"0C",X"09",X"83",X"20",X"00",X"B0",X"74",
		X"01",X"80",X"06",X"01",X"58",X"20",X"06",X"01",X"57",X"20",X"0B",X"11",X"20",X"63",X"1B",X"06",
		X"00",X"57",X"20",X"04",X"00",X"02",X"1B",X"00",X"1A",X"13",X"CD",X"8B",X"1C",X"EB",X"4F",X"21",
		X"4E",X"1E",X"7E",X"23",X"A7",X"F2",X"72",X"1B",X"0D",X"C2",X"72",X"1B",X"E6",X"7F",X"C3",X"30",
		X"01",X"EB",X"7E",X"32",X"23",X"20",X"23",X"22",X"06",X"20",X"C9",X"EB",X"7E",X"32",X"22",X"20",
		X"23",X"5E",X"23",X"56",X"23",X"22",X"06",X"20",X"EB",X"22",X"0F",X"20",X"C9",X"EB",X"5E",X"23",
		X"56",X"EB",X"22",X"06",X"20",X"C9",X"EB",X"7E",X"23",X"5E",X"23",X"56",X"23",X"22",X"06",X"20",
		X"12",X"C9",X"21",X"0D",X"20",X"7E",X"23",X"B6",X"FE",X"04",X"F2",X"BE",X"1B",X"AF",X"32",X"47",
		X"20",X"21",X"AF",X"0D",X"11",X"0D",X"3A",X"CD",X"F7",X"1B",X"21",X"14",X"1A",X"3A",X"0D",X"20",
		X"CD",X"D9",X"1B",X"21",X"08",X"1A",X"3A",X"0E",X"20",X"A7",X"C8",X"FE",X"03",X"FA",X"E2",X"1B",
		X"3E",X"03",X"F5",X"5E",X"23",X"56",X"23",X"D5",X"5E",X"23",X"56",X"23",X"E3",X"CD",X"F7",X"1B",
		X"E1",X"F1",X"3D",X"C2",X"E2",X"1B",X"C9",X"4E",X"23",X"46",X"23",X"EB",X"C5",X"E5",X"1A",X"13",
		X"77",X"23",X"0D",X"C2",X"FE",X"1B",X"E1",X"01",X"20",X"00",X"09",X"C1",X"05",X"C2",X"FC",X"1B",
		X"C9",X"EB",X"5E",X"23",X"56",X"23",X"0E",X"05",X"7E",X"23",X"12",X"1B",X"0D",X"C2",X"18",X"1C",
		X"22",X"06",X"20",X"C9",X"11",X"0D",X"20",X"01",X"29",X"20",X"CD",X"44",X"1C",X"13",X"CD",X"44",
		X"1C",X"11",X"00",X"24",X"21",X"29",X"20",X"3E",X"02",X"CD",X"30",X"01",X"11",X"1E",X"24",X"3E",
		X"02",X"C3",X"30",X"01",X"1A",X"1F",X"1F",X"1F",X"1F",X"E6",X"0F",X"C2",X"50",X"1C",X"3E",X"10",
		X"C6",X"30",X"02",X"03",X"1A",X"E6",X"0F",X"C6",X"30",X"02",X"03",X"C9",X"EB",X"4E",X"23",X"46",
		X"23",X"5E",X"23",X"56",X"23",X"0A",X"A7",X"C2",X"6B",X"1C",X"EB",X"22",X"06",X"20",X"C9",X"21",
		X"0D",X"3A",X"11",X"BD",X"20",X"01",X"06",X"24",X"C3",X"FC",X"1B",X"CD",X"8B",X"1C",X"E9",X"CD",
		X"8B",X"1C",X"3A",X"0A",X"20",X"A7",X"C8",X"22",X"00",X"20",X"C9",X"EB",X"5E",X"23",X"56",X"23",
		X"22",X"06",X"20",X"EB",X"C9",X"3A",X"12",X"20",X"0E",X"05",X"FE",X"04",X"D2",X"B0",X"1C",X"3D",
		X"07",X"07",X"47",X"DB",X"02",X"E6",X"03",X"B0",X"4F",X"06",X"00",X"21",X"17",X"1D",X"09",X"4E",
		X"11",X"00",X"28",X"11",X"00",X"28",X"04",X"79",X"A7",X"1F",X"4F",X"D2",X"CE",X"1C",X"C5",X"D5",
		X"78",X"CD",X"6E",X"1B",X"E1",X"11",X"00",X"02",X"19",X"EB",X"C1",X"C3",X"B6",X"1C",X"C2",X"B6",
		X"1C",X"D3",X"04",X"DB",X"02",X"2F",X"E6",X"A0",X"CA",X"D1",X"1C",X"07",X"E6",X"01",X"4F",X"DB",
		X"02",X"07",X"E6",X"06",X"B1",X"4F",X"06",X"00",X"21",X"23",X"1D",X"09",X"46",X"21",X"12",X"20",
		X"7E",X"90",X"FA",X"D1",X"1C",X"F3",X"7E",X"90",X"77",X"79",X"E6",X"01",X"3D",X"32",X"11",X"20",
		X"3D",X"32",X"0A",X"20",X"DB",X"02",X"E6",X"0C",X"07",X"07",X"C6",X"64",X"32",X"08",X"20",X"AF",
		X"32",X"0D",X"20",X"32",X"0E",X"20",X"C9",X"2B",X"05",X"08",X"08",X"05",X"05",X"33",X"05",X"05",
		X"05",X"2B",X"05",X"01",X"02",X"01",X"01",X"02",X"04",X"02",X"02",X"3A",X"49",X"20",X"A7",X"C0",
		X"3E",X"01",X"CD",X"C2",X"17",X"32",X"71",X"20",X"21",X"6E",X"20",X"7E",X"E6",X"0F",X"B0",X"77",
		X"2B",X"7E",X"F6",X"42",X"77",X"C3",X"61",X"16",X"3A",X"12",X"20",X"A7",X"C2",X"D1",X"16",X"C9",
		X"00",X"00",X"3F",X"13",X"1D",X"16",X"33",X"18",X"3F",X"1A",X"05",X"1D",X"01",X"1F",X"39",X"20",
		X"27",X"22",X"11",X"24",X"35",X"25",X"13",X"27",X"2B",X"28",X"3F",X"29",X"0F",X"2B",X"19",X"2C",
		X"1F",X"2D",X"21",X"2E",X"21",X"2F",X"1D",X"30",X"15",X"31",X"09",X"32",X"3B",X"32",X"29",X"33",
		X"17",X"34",X"3F",X"34",X"27",X"35",X"0D",X"36",X"31",X"36",X"11",X"37",X"31",X"37",X"0F",X"38",
		X"2B",X"38",X"05",X"39",X"1D",X"39",X"35",X"39",X"0B",X"3A",X"21",X"3A",X"84",X"06",X"14",X"02",
		X"12",X"03",X"11",X"01",X"0F",X"0A",X"11",X"01",X"08",X"01",X"08",X"04",X"0D",X"01",X"0D",X"01",
		X"0D",X"03",X"0D",X"01",X"0C",X"02",X"0D",X"0A",X"0F",X"00",X"84",X"01",X"15",X"02",X"00",X"02",
		X"0E",X"01",X"11",X"03",X"10",X"03",X"0C",X"00",X"84",X"04",X"0F",X"03",X"0F",X"01",X"0F",X"04",
		X"0F",X"03",X"12",X"01",X"11",X"03",X"11",X"01",X"0F",X"03",X"0F",X"01",X"0E",X"08",X"0F",X"00",
		X"84",X"02",X"08",X"01",X"0D",X"01",X"0D",X"02",X"11",X"0A",X"14",X"01",X"14",X"01",X"14",X"02",
		X"11",X"02",X"0D",X"0A",X"11",X"00",X"86",X"03",X"0A",X"01",X"0A",X"06",X"0F",X"03",X"0A",X"01",
		X"0F",X"06",X"13",X"03",X"0A",X"01",X"0F",X"02",X"13",X"03",X"0A",X"01",X"0F",X"02",X"13",X"03",
		X"0A",X"01",X"0F",X"06",X"13",X"03",X"0F",X"01",X"13",X"04",X"16",X"02",X"13",X"02",X"0F",X"06",
		X"0A",X"03",X"0A",X"01",X"0A",X"06",X"0F",X"00",X"40",X"40",X"40",X"40",X"40",X"40",X"55",X"47",
		X"48",X"5B",X"50",X"4F",X"57",X"5B",X"5A",X"41",X"50",X"5B",X"57",X"41",X"4D",X"5B",X"42",X"41",
		X"4D",X"5B",X"54",X"48",X"55",X"44",X"55",X"4D",X"46",X"5B",X"41",X"52",X"47",X"5B",X"8D",X"27",
		X"54",X"4F",X"40",X"53",X"54",X"41",X"52",X"54",X"40",X"47",X"41",X"4D",X"45",X"95",X"2B",X"50",
		X"52",X"45",X"53",X"53",X"40",X"31",X"40",X"50",X"4C",X"41",X"59",X"45",X"52",X"40",X"42",X"55",
		X"54",X"54",X"4F",X"4E",X"9A",X"2D",X"50",X"52",X"45",X"53",X"53",X"40",X"31",X"40",X"4F",X"52",
		X"40",X"32",X"40",X"50",X"4C",X"41",X"59",X"45",X"52",X"40",X"42",X"55",X"54",X"54",X"4F",X"4E",
		X"92",X"29",X"49",X"4E",X"53",X"45",X"52",X"54",X"40",X"31",X"40",X"4D",X"4F",X"52",X"45",X"40",
		X"43",X"4F",X"49",X"4E",X"93",X"2A",X"49",X"4E",X"53",X"45",X"52",X"54",X"40",X"32",X"40",X"4D",
		X"4F",X"52",X"45",X"40",X"43",X"4F",X"49",X"4E",X"53",X"93",X"2A",X"46",X"4F",X"52",X"40",X"54",
		X"57",X"4F",X"40",X"50",X"4C",X"41",X"59",X"45",X"52",X"40",X"47",X"41",X"4D",X"45",X"89",X"89",
		X"24",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"89",X"25",X"42",X"4F",X"4F",X"54",
		X"40",X"48",X"49",X"4C",X"4C",X"8B",X"26",X"49",X"4E",X"53",X"45",X"52",X"54",X"40",X"43",X"4F",
		X"49",X"4E",X"40",X"89",X"24",X"47",X"45",X"54",X"40",X"52",X"45",X"41",X"44",X"59",X"89",X"24",
		X"40",X"40",X"44",X"52",X"41",X"57",X"5B",X"40",X"40",X"8C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",
		X"20",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"89",X"24",X"47",X"41",X"4D",X"45",X"40",X"4F",X"56",
		X"45",X"52",X"87",X"53",X"48",X"4F",X"54",X"13",X"4D",X"45",X"5B",X"87",X"40",X"40",X"40",X"40",
		X"13",X"40",X"40",X"40",X"9A",X"27",X"54",X"57",X"4F",X"40",X"50",X"4C",X"41",X"59",X"45",X"52",
		X"40",X"4F",X"52",X"1D",X"53",X"49",X"4E",X"47",X"4C",X"45",X"40",X"50",X"4C",X"41",X"59",X"45",
		X"52",X"B2",X"2A",X"55",X"53",X"45",X"40",X"50",X"4C",X"41",X"59",X"45",X"52",X"40",X"31",X"40",
		X"48",X"41",X"4E",X"44",X"4C",X"45",X"53",X"28",X"43",X"4F",X"4D",X"50",X"55",X"54",X"45",X"52",
		X"40",X"43",X"4F",X"4E",X"54",X"52",X"4F",X"4C",X"53",X"40",X"4F",X"54",X"48",X"45",X"52",X"40",
		X"43",X"4F",X"57",X"42",X"4F",X"59",X"99",X"2D",X"4D",X"41",X"59",X"40",X"54",X"48",X"45",X"40",
		X"42",X"45",X"54",X"54",X"45",X"52",X"40",X"43",X"4F",X"57",X"42",X"4F",X"59",X"40",X"57",X"49",
		X"4E",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
