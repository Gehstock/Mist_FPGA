library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_6P is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_6P is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"CC",X"FF",X"EE",X"EE",X"EE",X"FF",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"00",X"00",
		X"FF",X"CC",X"FF",X"EE",X"EE",X"EE",X"FF",X"CC",X"EE",X"EE",X"FF",X"EE",X"FF",X"CC",X"00",X"00",
		X"77",X"CC",X"FF",X"EE",X"FF",X"EE",X"EE",X"00",X"FF",X"EE",X"FF",X"EE",X"77",X"CC",X"00",X"00",
		X"FF",X"CC",X"FF",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"FF",X"EE",X"FF",X"CC",X"00",X"00",
		X"FF",X"EE",X"FF",X"EE",X"EE",X"00",X"FF",X"CC",X"EE",X"00",X"FF",X"EE",X"FF",X"EE",X"00",X"00",
		X"FF",X"EE",X"FF",X"EE",X"EE",X"00",X"FF",X"CC",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"00",X"00",
		X"77",X"CC",X"FF",X"EE",X"FF",X"EE",X"EE",X"00",X"EE",X"EE",X"FF",X"EE",X"77",X"EE",X"00",X"00",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"FF",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"00",X"00",
		X"33",X"CC",X"33",X"CC",X"33",X"CC",X"33",X"CC",X"33",X"CC",X"33",X"CC",X"33",X"CC",X"00",X"00",
		X"00",X"EE",X"00",X"EE",X"00",X"EE",X"66",X"EE",X"66",X"EE",X"77",X"EE",X"33",X"CC",X"00",X"00",
		X"EE",X"EE",X"EE",X"EE",X"FF",X"CC",X"FF",X"88",X"FF",X"CC",X"EE",X"EE",X"EE",X"EE",X"00",X"00",
		X"EE",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"FF",X"EE",X"FF",X"EE",X"00",X"00",
		X"EE",X"EE",X"FE",X"EE",X"FF",X"EE",X"FF",X"EE",X"FF",X"EE",X"FD",X"E6",X"DD",X"66",X"00",X"00",
		X"EE",X"66",X"FF",X"66",X"FF",X"EE",X"FF",X"EE",X"FF",X"EE",X"DD",X"EE",X"CC",X"EE",X"00",X"00",
		X"77",X"CC",X"FF",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"FF",X"EE",X"77",X"CC",X"00",X"00",
		X"FF",X"CC",X"FF",X"EE",X"EE",X"EE",X"FF",X"CC",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"00",X"00",
		X"77",X"CC",X"FF",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"FF",X"EE",X"77",X"CC",X"00",X"EE",
		X"FF",X"CC",X"FF",X"EE",X"EE",X"EE",X"FF",X"C8",X"FF",X"CC",X"EE",X"EE",X"EE",X"EE",X"00",X"00",
		X"77",X"EE",X"FF",X"EE",X"EE",X"00",X"FF",X"EE",X"00",X"EE",X"FF",X"EE",X"FF",X"CC",X"00",X"00",
		X"FF",X"EE",X"FF",X"EE",X"33",X"88",X"33",X"88",X"33",X"88",X"33",X"88",X"33",X"88",X"00",X"00",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"FF",X"EE",X"FF",X"EE",X"77",X"CC",X"00",X"00",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"66",X"CC",X"77",X"CC",X"33",X"88",X"33",X"88",X"00",X"00",
		X"DD",X"66",X"FD",X"E6",X"FF",X"EE",X"FF",X"EE",X"FF",X"EE",X"FE",X"EE",X"EE",X"EE",X"00",X"00",
		X"EC",X"E6",X"FE",X"EE",X"F7",X"EC",X"73",X"C8",X"F7",X"EC",X"FE",X"EE",X"EC",X"E6",X"00",X"00",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"77",X"CC",X"33",X"88",X"33",X"88",X"33",X"88",X"00",X"00",
		X"FF",X"EE",X"FF",X"EE",X"11",X"EE",X"77",X"CC",X"FF",X"00",X"FF",X"EE",X"FF",X"EE",X"00",X"00",
		X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"00",X"33",X"00",X"77",X"00",X"FF",X"11",X"FF",X"33",X"FF",X"77",X"FF",X"FF",X"FF",
		X"88",X"00",X"CC",X"00",X"EE",X"00",X"FF",X"00",X"FF",X"88",X"FF",X"CC",X"FF",X"EE",X"FF",X"FF",
		X"FF",X"FF",X"77",X"FF",X"33",X"FF",X"11",X"FF",X"00",X"FF",X"00",X"77",X"00",X"33",X"00",X"11",
		X"FF",X"FF",X"FF",X"EE",X"FF",X"CC",X"FF",X"88",X"FF",X"00",X"EE",X"00",X"CC",X"00",X"88",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"33",X"00",X"33",X"00",X"33",X"00",X"11",X"00",X"11",X"00",X"00",X"00",X"33",X"00",X"00",X"00",
		X"00",X"00",X"22",X"88",X"22",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"88",X"22",X"88",X"FF",X"EE",X"22",X"88",X"FF",X"EE",X"22",X"88",X"22",X"88",X"00",X"00",
		X"11",X"00",X"F7",X"EC",X"D9",X"00",X"F7",X"EC",X"11",X"62",X"F7",X"EC",X"11",X"00",X"00",X"00",
		X"E4",X"22",X"AA",X"44",X"E4",X"88",X"11",X"00",X"22",X"E4",X"44",X"AA",X"88",X"E4",X"00",X"00",
		X"72",X"00",X"55",X"00",X"22",X"00",X"75",X"00",X"98",X"AA",X"C8",X"C4",X"77",X"AA",X"00",X"00",
		X"11",X"88",X"10",X"88",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"88",X"11",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"11",X"00",X"00",X"88",X"00",X"00",
		X"11",X"00",X"00",X"88",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"88",X"11",X"00",X"00",X"00",
		X"00",X"00",X"11",X"00",X"55",X"44",X"22",X"88",X"22",X"88",X"55",X"44",X"11",X"00",X"00",X"00",
		X"00",X"00",X"11",X"00",X"11",X"00",X"77",X"CC",X"11",X"00",X"11",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"88",X"00",X"88",X"11",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"33",X"00",X"00",X"00",
		X"00",X"11",X"00",X"32",X"00",X"64",X"00",X"C8",X"11",X"80",X"32",X"00",X"64",X"00",X"C8",X"00",
		X"33",X"88",X"66",X"CC",X"CC",X"66",X"CC",X"66",X"CC",X"66",X"66",X"CC",X"33",X"88",X"00",X"00",
		X"11",X"88",X"33",X"88",X"77",X"88",X"11",X"88",X"11",X"88",X"11",X"88",X"77",X"EE",X"00",X"00",
		X"77",X"CC",X"CC",X"66",X"00",X"EE",X"33",X"CC",X"77",X"88",X"EE",X"00",X"FF",X"EE",X"00",X"00",
		X"77",X"EE",X"00",X"CC",X"11",X"88",X"33",X"CC",X"00",X"66",X"CC",X"66",X"77",X"CC",X"00",X"00",
		X"11",X"CC",X"33",X"CC",X"66",X"CC",X"CC",X"CC",X"FF",X"EE",X"00",X"CC",X"00",X"CC",X"00",X"00",
		X"FF",X"CC",X"CC",X"00",X"FF",X"CC",X"00",X"66",X"00",X"66",X"CC",X"66",X"77",X"CC",X"00",X"00",
		X"33",X"CC",X"66",X"00",X"CC",X"00",X"FF",X"CC",X"CC",X"66",X"CC",X"66",X"77",X"CC",X"00",X"00",
		X"FF",X"EE",X"CC",X"66",X"00",X"CC",X"11",X"88",X"33",X"00",X"33",X"00",X"33",X"00",X"00",X"00",
		X"77",X"CC",X"CC",X"66",X"CC",X"66",X"77",X"CC",X"CC",X"66",X"CC",X"66",X"77",X"CC",X"00",X"00",
		X"77",X"CC",X"CC",X"66",X"CC",X"66",X"77",X"EE",X"00",X"66",X"00",X"CC",X"77",X"88",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"88",X"11",X"88",X"00",X"00",X"11",X"88",X"11",X"88",X"00",X"00",
		X"11",X"00",X"33",X"00",X"77",X"EE",X"FF",X"EE",X"77",X"EE",X"33",X"00",X"11",X"00",X"00",X"00",
		X"00",X"44",X"00",X"88",X"11",X"00",X"22",X"00",X"11",X"00",X"00",X"88",X"00",X"44",X"00",X"00",
		X"00",X"00",X"00",X"00",X"77",X"CC",X"00",X"00",X"77",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"00",X"11",X"00",X"00",X"88",X"00",X"44",X"00",X"88",X"11",X"00",X"22",X"00",X"00",X"00",
		X"33",X"CC",X"66",X"66",X"66",X"66",X"00",X"CC",X"11",X"88",X"11",X"88",X"00",X"00",X"11",X"88",
		X"33",X"CC",X"44",X"22",X"99",X"99",X"AA",X"11",X"AA",X"11",X"99",X"99",X"44",X"22",X"33",X"CC",
		X"33",X"88",X"66",X"CC",X"CC",X"66",X"CC",X"66",X"FF",X"EE",X"CC",X"66",X"CC",X"66",X"00",X"00",
		X"FF",X"CC",X"CC",X"66",X"CC",X"66",X"FF",X"CC",X"CC",X"66",X"CC",X"66",X"FF",X"CC",X"00",X"00",
		X"77",X"CC",X"CC",X"66",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"66",X"77",X"CC",X"00",X"00",
		X"FF",X"88",X"CC",X"CC",X"CC",X"66",X"CC",X"66",X"CC",X"66",X"CC",X"CC",X"FF",X"88",X"00",X"00",
		X"FF",X"EE",X"CC",X"00",X"CC",X"00",X"FF",X"88",X"CC",X"00",X"CC",X"00",X"FF",X"EE",X"00",X"00",
		X"FF",X"EE",X"CC",X"00",X"CC",X"00",X"FF",X"88",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"00",X"00",
		X"33",X"EE",X"66",X"00",X"CC",X"00",X"CC",X"EE",X"CC",X"66",X"66",X"66",X"33",X"EE",X"00",X"00",
		X"CC",X"66",X"CC",X"66",X"CC",X"66",X"FF",X"EE",X"CC",X"66",X"CC",X"66",X"CC",X"66",X"00",X"00",
		X"77",X"EE",X"11",X"88",X"11",X"88",X"11",X"88",X"11",X"88",X"11",X"88",X"77",X"EE",X"00",X"00",
		X"00",X"66",X"00",X"66",X"00",X"66",X"00",X"66",X"CC",X"66",X"CC",X"66",X"77",X"CC",X"00",X"00",
		X"CC",X"66",X"CC",X"CC",X"DD",X"88",X"FF",X"00",X"FF",X"88",X"CC",X"CC",X"CC",X"66",X"00",X"00",
		X"66",X"00",X"66",X"00",X"66",X"00",X"66",X"00",X"66",X"00",X"66",X"00",X"77",X"EE",X"00",X"00",
		X"CC",X"66",X"EE",X"EE",X"FF",X"EE",X"FF",X"EE",X"DD",X"66",X"CC",X"66",X"CC",X"66",X"00",X"00",
		X"CC",X"66",X"EE",X"66",X"FF",X"66",X"FF",X"EE",X"DD",X"EE",X"CC",X"EE",X"CC",X"66",X"00",X"00",
		X"77",X"CC",X"CC",X"66",X"CC",X"66",X"CC",X"66",X"CC",X"66",X"CC",X"66",X"77",X"CC",X"00",X"00",
		X"FF",X"CC",X"CC",X"66",X"CC",X"66",X"CC",X"66",X"FF",X"CC",X"CC",X"00",X"CC",X"00",X"00",X"00",
		X"77",X"CC",X"CC",X"66",X"CC",X"66",X"CC",X"66",X"DD",X"EE",X"CC",X"CC",X"77",X"AA",X"00",X"00",
		X"FF",X"CC",X"CC",X"66",X"CC",X"66",X"CC",X"CC",X"FF",X"88",X"DD",X"CC",X"CC",X"EE",X"00",X"00",
		X"77",X"88",X"CC",X"C4",X"CC",X"00",X"77",X"CC",X"00",X"66",X"CC",X"66",X"77",X"CC",X"00",X"00",
		X"77",X"EE",X"11",X"88",X"11",X"88",X"11",X"88",X"11",X"88",X"11",X"88",X"11",X"88",X"00",X"00",
		X"CC",X"66",X"CC",X"66",X"CC",X"66",X"CC",X"66",X"CC",X"66",X"CC",X"66",X"77",X"CC",X"00",X"00",
		X"CC",X"66",X"CC",X"66",X"CC",X"66",X"EE",X"EE",X"77",X"CC",X"33",X"88",X"11",X"00",X"00",X"00",
		X"CC",X"66",X"CC",X"66",X"DD",X"66",X"FF",X"EE",X"FF",X"EE",X"EE",X"EE",X"CC",X"66",X"00",X"00",
		X"CC",X"66",X"EE",X"EE",X"77",X"CC",X"33",X"88",X"77",X"CC",X"EE",X"EE",X"CC",X"66",X"00",X"00",
		X"66",X"66",X"66",X"66",X"66",X"66",X"33",X"CC",X"11",X"88",X"11",X"88",X"11",X"88",X"00",X"00",
		X"FF",X"EE",X"00",X"EE",X"11",X"CC",X"33",X"88",X"77",X"00",X"EE",X"00",X"FF",X"EE",X"00",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",
		X"44",X"00",X"44",X"44",X"44",X"88",X"55",X"66",X"22",X"99",X"44",X"22",X"00",X"44",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"33",X"EE",X"66",X"66",X"66",X"66",X"66",X"EE",X"33",X"66",X"00",X"00",
		X"66",X"00",X"66",X"00",X"77",X"CC",X"66",X"66",X"66",X"66",X"66",X"66",X"77",X"CC",X"00",X"00",
		X"00",X"00",X"00",X"00",X"33",X"CC",X"66",X"66",X"66",X"00",X"66",X"66",X"33",X"CC",X"00",X"00",
		X"00",X"66",X"00",X"66",X"33",X"EE",X"66",X"66",X"66",X"66",X"66",X"66",X"33",X"EE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"33",X"CC",X"66",X"66",X"77",X"EE",X"66",X"00",X"33",X"CC",X"00",X"00",
		X"11",X"CC",X"33",X"66",X"33",X"00",X"77",X"CC",X"33",X"00",X"33",X"00",X"33",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"33",X"EE",X"66",X"66",X"66",X"66",X"33",X"EE",X"00",X"66",X"33",X"CC",
		X"66",X"00",X"66",X"00",X"77",X"CC",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"00",X"00",
		X"11",X"88",X"00",X"00",X"33",X"88",X"11",X"88",X"11",X"88",X"11",X"88",X"33",X"CC",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"11",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"44",X"CC",X"33",X"88",
		X"66",X"00",X"66",X"66",X"66",X"CC",X"77",X"88",X"77",X"88",X"66",X"CC",X"66",X"66",X"00",X"00",
		X"33",X"88",X"11",X"88",X"11",X"88",X"11",X"88",X"11",X"88",X"11",X"88",X"33",X"CC",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"CC",X"DD",X"66",X"DD",X"66",X"DD",X"66",X"DD",X"66",X"00",X"00",
		X"00",X"00",X"00",X"00",X"77",X"CC",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"00",X"00",
		X"00",X"00",X"00",X"00",X"33",X"CC",X"66",X"66",X"66",X"66",X"66",X"66",X"33",X"CC",X"00",X"00",
		X"00",X"00",X"00",X"00",X"77",X"CC",X"66",X"66",X"66",X"66",X"77",X"CC",X"66",X"00",X"66",X"00",
		X"00",X"00",X"00",X"00",X"77",X"CC",X"CC",X"CC",X"CC",X"CC",X"77",X"CC",X"00",X"CC",X"00",X"EE",
		X"00",X"00",X"00",X"00",X"77",X"CC",X"76",X"62",X"66",X"00",X"66",X"00",X"66",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"73",X"CC",X"66",X"00",X"73",X"EC",X"00",X"66",X"77",X"EC",X"00",X"00",
		X"11",X"88",X"11",X"88",X"77",X"EE",X"11",X"88",X"11",X"88",X"11",X"88",X"00",X"EE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"EE",X"33",X"66",X"00",X"00",
		X"00",X"00",X"00",X"00",X"66",X"66",X"66",X"66",X"66",X"66",X"33",X"CC",X"11",X"88",X"00",X"00",
		X"00",X"00",X"00",X"00",X"DD",X"66",X"DD",X"66",X"DD",X"66",X"DD",X"66",X"76",X"CC",X"00",X"00",
		X"00",X"00",X"00",X"00",X"CC",X"CC",X"77",X"88",X"33",X"00",X"77",X"88",X"CC",X"CC",X"00",X"00",
		X"00",X"00",X"00",X"00",X"66",X"66",X"66",X"66",X"66",X"66",X"33",X"EE",X"00",X"66",X"33",X"CC",
		X"00",X"00",X"00",X"00",X"77",X"EE",X"00",X"CC",X"11",X"88",X"33",X"00",X"77",X"EE",X"00",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"72",X"00",X"F6",X"10",X"BA",X"77",X"FE",X"72",X"32",X"E4",X"32",X"C8",X"32",X"00",X"00",
		X"F7",X"88",X"C4",X"88",X"F7",X"EC",X"C4",X"62",X"C4",X"62",X"C4",X"E4",X"F7",X"C8",X"00",X"00",
		X"31",X"EE",X"72",X"00",X"E4",X"00",X"C4",X"00",X"E4",X"00",X"72",X"00",X"31",X"EE",X"00",X"00",
		X"F7",X"C8",X"C4",X"E4",X"C4",X"72",X"C4",X"32",X"C4",X"72",X"C4",X"E4",X"F7",X"C8",X"00",X"00",
		X"F7",X"88",X"C4",X"00",X"F7",X"00",X"C4",X"00",X"C4",X"00",X"C4",X"00",X"F7",X"EE",X"00",X"00",
		X"F7",X"EE",X"C4",X"00",X"F7",X"88",X"C4",X"00",X"C4",X"00",X"C4",X"00",X"C4",X"00",X"00",X"00",
		X"31",X"EE",X"72",X"00",X"E4",X"00",X"C4",X"00",X"E4",X"66",X"72",X"62",X"31",X"EC",X"00",X"00",
		X"C4",X"62",X"C4",X"62",X"F7",X"EE",X"C4",X"62",X"C4",X"62",X"C4",X"62",X"C4",X"62",X"00",X"00",
		X"73",X"EE",X"10",X"88",X"10",X"88",X"10",X"88",X"10",X"88",X"10",X"88",X"73",X"EE",X"00",X"00",
		X"00",X"62",X"00",X"62",X"00",X"62",X"00",X"62",X"00",X"62",X"C4",X"62",X"73",X"EC",X"00",X"00",
		X"D4",X"88",X"F5",X"80",X"F6",X"00",X"F5",X"80",X"D4",X"C8",X"C4",X"E4",X"C4",X"62",X"00",X"00",
		X"C4",X"00",X"C4",X"00",X"C4",X"00",X"C4",X"00",X"C4",X"00",X"C4",X"00",X"F7",X"EE",X"00",X"00",
		X"E4",X"62",X"F6",X"E6",X"D5",X"EA",X"C4",X"62",X"C4",X"62",X"C4",X"62",X"C4",X"62",X"00",X"00",
		X"C4",X"62",X"E6",X"62",X"F7",X"62",X"D5",X"EA",X"C4",X"EE",X"C4",X"66",X"C4",X"22",X"00",X"00",
		X"31",X"CC",X"62",X"62",X"C4",X"31",X"C4",X"31",X"C4",X"31",X"62",X"62",X"31",X"CC",X"00",X"00",
		X"F7",X"88",X"C4",X"C4",X"C4",X"62",X"C4",X"62",X"C4",X"C4",X"F7",X"88",X"C4",X"00",X"00",X"00",
		X"31",X"CC",X"62",X"62",X"C4",X"31",X"C4",X"31",X"C4",X"F5",X"62",X"62",X"31",X"F9",X"00",X"00",
		X"F7",X"88",X"C4",X"C4",X"C4",X"62",X"C4",X"62",X"C4",X"C4",X"F7",X"88",X"C4",X"E6",X"00",X"00",
		X"73",X"88",X"C4",X"00",X"73",X"C8",X"00",X"64",X"00",X"62",X"00",X"64",X"F7",X"C8",X"00",X"00",
		X"F7",X"FF",X"10",X"88",X"10",X"88",X"10",X"88",X"10",X"88",X"10",X"88",X"10",X"88",X"00",X"00",
		X"C4",X"62",X"C4",X"62",X"C4",X"62",X"C4",X"62",X"C4",X"62",X"C4",X"62",X"73",X"CC",X"00",X"00",
		X"C4",X"31",X"C4",X"72",X"C4",X"E4",X"D4",X"C8",X"F5",X"80",X"F6",X"00",X"E4",X"00",X"00",X"00",
		X"C4",X"62",X"C4",X"62",X"C4",X"62",X"C4",X"62",X"D5",X"EA",X"F6",X"E6",X"E4",X"62",X"00",X"00",
		X"E4",X"31",X"72",X"72",X"31",X"E4",X"10",X"C8",X"31",X"E4",X"72",X"72",X"E4",X"31",X"00",X"00",
		X"E4",X"31",X"72",X"72",X"31",X"E4",X"10",X"C8",X"31",X"80",X"72",X"00",X"E4",X"00",X"00",X"00",
		X"FF",X"EE",X"00",X"E4",X"10",X"C8",X"31",X"80",X"72",X"00",X"E4",X"00",X"FF",X"EE",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"00",X"31",X"00",X"72",X"00",X"31",X"80",X"10",X"C8",X"11",X"80",X"00",X"C8",X"00",X"44",
		X"11",X"00",X"33",X"88",X"77",X"CC",X"FF",X"EE",X"77",X"CC",X"33",X"88",X"11",X"00",X"00",X"00",
		X"FF",X"EE",X"88",X"22",X"BB",X"AA",X"BB",X"AA",X"BB",X"AA",X"88",X"22",X"FF",X"EE",X"00",X"00",
		X"FA",X"FA",X"F5",X"F5",X"FA",X"FA",X"F5",X"F5",X"FA",X"FA",X"F5",X"F5",X"FA",X"FA",X"F5",X"F5",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"03",X"0C",X"02",X"04",X"03",X"0C",X"01",X"08",X"01",X"08",X"01",X"0E",X"01",X"08",X"01",X"0E",
		X"00",X"11",X"00",X"32",X"00",X"64",X"04",X"C8",X"13",X"80",X"21",X"00",X"42",X"08",X"84",X"00",
		X"11",X"84",X"11",X"84",X"11",X"84",X"32",X"C2",X"74",X"E1",X"74",X"E1",X"32",X"C3",X"03",X"0E",
		X"00",X"00",X"99",X"77",X"99",X"44",X"FF",X"77",X"99",X"44",X"99",X"44",X"99",X"77",X"00",X"00",
		X"00",X"00",X"9B",X"99",X"22",X"55",X"22",X"55",X"33",X"DD",X"22",X"55",X"AA",X"55",X"00",X"00",
		X"00",X"00",X"11",X"FF",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"EE",X"44",X"00",X"00",
		X"00",X"00",X"44",X"88",X"44",X"88",X"77",X"88",X"44",X"88",X"44",X"88",X"44",X"88",X"00",X"00",
		X"00",X"00",X"F7",X"33",X"88",X"44",X"F6",X"44",X"11",X"44",X"11",X"44",X"EE",X"33",X"00",X"00",
		X"00",X"00",X"9B",X"9D",X"22",X"55",X"22",X"55",X"22",X"55",X"22",X"55",X"9B",X"9D",X"00",X"00",
		X"00",X"00",X"EC",X"FF",X"22",X"88",X"E4",X"EE",X"88",X"88",X"44",X"88",X"22",X"FF",X"00",X"00",
		X"00",X"00",X"88",X"9B",X"88",X"AA",X"88",X"AA",X"AA",X"BB",X"AA",X"AA",X"55",X"22",X"00",X"00",
		X"00",X"00",X"99",X"EC",X"55",X"22",X"55",X"E4",X"DD",X"88",X"55",X"44",X"55",X"22",X"00",X"00",
		X"00",X"00",X"FE",X"45",X"99",X"55",X"FA",X"55",X"CC",X"55",X"AA",X"55",X"99",X"45",X"00",X"00",
		X"00",X"00",X"CE",X"FE",X"22",X"99",X"22",X"FA",X"22",X"CC",X"22",X"AA",X"CE",X"99",X"00",X"00",
		X"00",X"00",X"88",X"99",X"88",X"AA",X"88",X"AA",X"88",X"BB",X"55",X"22",X"22",X"22",X"00",X"00",
		X"00",X"00",X"99",X"00",X"55",X"00",X"55",X"00",X"DD",X"00",X"55",X"00",X"55",X"EE",X"00",X"00",
		X"00",X"00",X"88",X"44",X"99",X"44",X"AA",X"22",X"CC",X"11",X"AA",X"11",X"99",X"11",X"00",X"00",
		X"00",X"00",X"55",X"EC",X"55",X"22",X"99",X"E4",X"11",X"88",X"11",X"44",X"11",X"22",X"00",X"00",
		X"00",X"00",X"BB",X"CC",X"AA",X"00",X"BB",X"88",X"AA",X"00",X"AA",X"00",X"BB",X"CC",X"00",X"00",
		X"00",X"00",X"88",X"AA",X"88",X"AA",X"88",X"AA",X"AA",X"AA",X"AA",X"AA",X"55",X"22",X"00",X"00",
		X"00",X"00",X"FF",X"33",X"11",X"44",X"22",X"44",X"44",X"77",X"88",X"44",X"FF",X"44",X"00",X"00",
		X"00",X"00",X"33",X"D9",X"AA",X"55",X"BA",X"D9",X"BB",X"11",X"AA",X"99",X"AA",X"55",X"00",X"00",
		X"00",X"00",X"CC",X"00",X"26",X"00",X"22",X"00",X"22",X"00",X"26",X"00",X"CC",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"44",X"88",X"44",X"EE",X"44",X"88",X"44",X"88",X"44",X"FF",X"77",X"00",X"00",
		X"00",X"00",X"33",X"CC",X"22",X"00",X"33",X"88",X"22",X"00",X"22",X"00",X"AA",X"00",X"00",X"00",
		X"00",X"00",X"00",X"70",X"10",X"F7",X"31",X"FC",X"73",X"C8",X"73",X"90",X"73",X"80",X"73",X"F0",
		X"00",X"00",X"F0",X"00",X"FF",X"F0",X"F7",X"F7",X"F6",X"71",X"EC",X"31",X"C0",X"73",X"F0",X"73",
		X"00",X"00",X"00",X"00",X"F0",X"F0",X"FF",X"FF",X"FF",X"B9",X"F9",X"FB",X"B1",X"FB",X"F1",X"FB",
		X"00",X"00",X"00",X"00",X"B0",X"E0",X"FB",X"FC",X"B8",X"EC",X"90",X"EC",X"90",X"EC",X"90",X"EC",
		X"00",X"00",X"00",X"00",X"F0",X"C0",X"FF",X"FC",X"F6",X"F7",X"F6",X"73",X"F6",X"31",X"F6",X"31",
		X"00",X"00",X"00",X"00",X"F0",X"F0",X"FF",X"FF",X"E6",X"F6",X"EA",X"F6",X"F9",X"F6",X"D8",X"F6",
		X"00",X"00",X"00",X"00",X"F0",X"70",X"FF",X"FF",X"76",X"F6",X"64",X"F6",X"C8",X"F6",X"80",X"F6",
		X"00",X"00",X"00",X"00",X"B0",X"F0",X"FB",X"FF",X"B0",X"FC",X"10",X"EC",X"10",X"EC",X"10",X"FC",
		X"00",X"00",X"00",X"00",X"F0",X"F0",X"FF",X"FF",X"F0",X"F3",X"20",X"73",X"72",X"73",X"F6",X"73",
		X"00",X"00",X"00",X"00",X"F0",X"E0",X"FF",X"EC",X"F0",X"EC",X"90",X"C8",X"B1",X"80",X"B0",X"00",
		X"73",X"FF",X"73",X"F0",X"73",X"80",X"73",X"F8",X"31",X"FF",X"10",X"FF",X"00",X"F0",X"00",X"00",
		X"FF",X"F7",X"F3",X"F6",X"73",X"F6",X"F3",X"F6",X"FF",X"F6",X"FF",X"F6",X"F3",X"F6",X"73",X"F6",
		X"FF",X"FB",X"F1",X"FB",X"31",X"FB",X"31",X"FB",X"31",X"FB",X"31",X"F9",X"31",X"D8",X"73",X"80",
		X"90",X"EC",X"90",X"EC",X"90",X"EC",X"90",X"EC",X"F9",X"FC",X"FE",X"FF",X"EC",X"F6",X"C0",X"60",
		X"F6",X"31",X"F6",X"31",X"F6",X"31",X"F6",X"B1",X"FE",X"F9",X"F7",X"F9",X"F7",X"B0",X"F6",X"00",
		X"C8",X"F6",X"C8",X"F6",X"C8",X"F6",X"C8",X"F6",X"C8",X"F6",X"C8",X"F6",X"C0",X"F0",X"00",X"00",
		X"00",X"F6",X"00",X"F6",X"00",X"F6",X"00",X"F6",X"30",X"F6",X"31",X"FF",X"30",X"F0",X"00",X"00",
		X"10",X"FF",X"30",X"FD",X"72",X"FD",X"F6",X"FC",X"FC",X"FC",X"FC",X"FF",X"D0",X"F0",X"00",X"00",
		X"EC",X"73",X"C8",X"73",X"90",X"F7",X"31",X"FB",X"F3",X"F3",X"FF",X"F3",X"F0",X"73",X"00",X"73",
		X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"B0",X"00",X"F2",X"00",X"F6",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"31",X"00",X"31",X"00",X"30",
		X"73",X"E4",X"73",X"C0",X"73",X"80",X"F6",X"00",X"EC",X"00",X"C8",X"00",X"80",X"00",X"00",X"00",
		X"72",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"00",X"10",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EC",X"00",X"C8",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"73",X"00",X"73",X"00",X"73",X"00",X"F6",X"10",X"EC",X"31",X"C8",X"31",X"80",X"30",X"00",
		X"EC",X"00",X"C8",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"33",X"77",X"77",X"33",X"EE",X"11",X"CC",X"33",X"EE",X"77",X"77",X"66",X"33",X"00",X"00",
		X"00",X"00",X"00",X"77",X"00",X"FF",X"77",X"88",X"77",X"88",X"00",X"FF",X"00",X"77",X"00",X"00",
		X"66",X"11",X"77",X"11",X"77",X"99",X"55",X"DD",X"44",X"FF",X"44",X"77",X"44",X"33",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",
		X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",
		X"00",X"00",X"22",X"FF",X"11",X"00",X"00",X"88",X"99",X"44",X"CC",X"AA",X"AA",X"88",X"99",X"00",
		X"00",X"00",X"33",X"88",X"77",X"CC",X"44",X"44",X"22",X"44",X"77",X"CC",X"77",X"CC",X"00",X"00",
		X"00",X"00",X"77",X"FF",X"77",X"FF",X"44",X"44",X"44",X"44",X"77",X"CC",X"33",X"88",X"00",X"00",
		X"00",X"00",X"33",X"88",X"77",X"CC",X"44",X"44",X"44",X"44",X"66",X"CC",X"22",X"88",X"00",X"00",
		X"00",X"00",X"33",X"88",X"77",X"CC",X"44",X"44",X"44",X"44",X"77",X"FF",X"77",X"FF",X"00",X"00",
		X"00",X"00",X"33",X"88",X"77",X"CC",X"55",X"44",X"55",X"44",X"55",X"CC",X"11",X"88",X"00",X"00",
		X"00",X"00",X"00",X"88",X"77",X"EE",X"77",X"FF",X"00",X"99",X"00",X"BB",X"00",X"22",X"00",X"00",
		X"00",X"00",X"11",X"88",X"BB",X"CC",X"AA",X"44",X"AA",X"44",X"FF",X"CC",X"77",X"CC",X"00",X"00",
		X"00",X"00",X"77",X"FF",X"77",X"FF",X"00",X"44",X"00",X"44",X"77",X"CC",X"77",X"88",X"00",X"00",
		X"00",X"00",X"00",X"00",X"44",X"44",X"77",X"DD",X"77",X"DD",X"44",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"44",X"00",X"88",X"00",X"88",X"44",X"FF",X"DD",X"77",X"DD",X"00",X"00",X"00",X"00",
		X"00",X"00",X"77",X"FF",X"77",X"FF",X"11",X"88",X"33",X"CC",X"66",X"66",X"44",X"22",X"00",X"00",
		X"00",X"00",X"00",X"00",X"44",X"11",X"77",X"FF",X"77",X"FF",X"44",X"00",X"00",X"00",X"00",X"00",
		X"77",X"CC",X"77",X"CC",X"00",X"44",X"77",X"CC",X"00",X"44",X"77",X"CC",X"77",X"88",X"00",X"00",
		X"00",X"00",X"77",X"CC",X"77",X"CC",X"00",X"44",X"00",X"44",X"77",X"CC",X"77",X"88",X"00",X"00",
		X"00",X"00",X"33",X"88",X"77",X"CC",X"44",X"44",X"44",X"44",X"77",X"CC",X"33",X"88",X"00",X"00",
		X"00",X"00",X"FF",X"CC",X"FF",X"CC",X"22",X"44",X"22",X"44",X"33",X"CC",X"11",X"88",X"00",X"00",
		X"11",X"88",X"33",X"CC",X"22",X"44",X"22",X"44",X"FF",X"CC",X"FF",X"CC",X"88",X"00",X"00",X"00",
		X"00",X"00",X"77",X"CC",X"77",X"CC",X"00",X"C4",X"00",X"44",X"00",X"44",X"00",X"C8",X"00",X"00",
		X"00",X"00",X"54",X"C8",X"55",X"CC",X"55",X"44",X"55",X"44",X"77",X"44",X"72",X"00",X"00",X"00",
		X"00",X"00",X"00",X"44",X"00",X"44",X"33",X"FF",X"77",X"FF",X"44",X"44",X"44",X"44",X"00",X"00",
		X"00",X"00",X"33",X"CC",X"77",X"CC",X"44",X"00",X"22",X"00",X"77",X"CC",X"77",X"CC",X"00",X"00",
		X"00",X"00",X"11",X"CC",X"33",X"CC",X"66",X"00",X"66",X"00",X"33",X"CC",X"11",X"CC",X"00",X"00",
		X"33",X"CC",X"77",X"CC",X"44",X"00",X"73",X"CC",X"44",X"00",X"77",X"CC",X"33",X"CC",X"00",X"00",
		X"44",X"44",X"66",X"CC",X"33",X"88",X"33",X"88",X"66",X"CC",X"44",X"44",X"00",X"00",X"00",X"00",
		X"00",X"00",X"11",X"CC",X"BB",X"CC",X"AA",X"00",X"AA",X"00",X"FF",X"CC",X"77",X"CC",X"00",X"00",
		X"00",X"00",X"44",X"44",X"66",X"44",X"77",X"44",X"55",X"CC",X"44",X"CC",X"44",X"44",X"00",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",
		X"00",X"07",X"00",X"7B",X"01",X"F6",X"12",X"ED",X"13",X"CE",X"13",X"CA",X"13",X"8C",X"13",X"8C",
		X"0F",X"08",X"FF",X"84",X"3D",X"CA",X"12",X"ED",X"01",X"EF",X"01",X"E7",X"00",X"6F",X"00",X"6F",
		X"13",X"8C",X"13",X"8C",X"13",X"CA",X"13",X"CE",X"12",X"ED",X"01",X"F6",X"00",X"7B",X"00",X"07",
		X"00",X"6F",X"00",X"6F",X"01",X"E7",X"01",X"EF",X"12",X"ED",X"3D",X"CA",X"FF",X"84",X"0F",X"08",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"13",X"00",X"37",X"00",X"07",X"00",X"01",X"00",X"01",
		X"06",X"00",X"4E",X"00",X"CE",X"00",X"CE",X"00",X"CE",X"00",X"CE",X"00",X"CE",X"00",X"CE",X"00",
		X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"16",X"00",X"7F",X"00",X"0F",
		X"CE",X"00",X"CE",X"00",X"CE",X"00",X"CE",X"00",X"CE",X"00",X"ED",X"08",X"FF",X"8C",X"0F",X"0C",
		X"00",X"07",X"00",X"7F",X"01",X"ED",X"13",X"CA",X"13",X"8C",X"01",X"08",X"00",X"00",X"00",X"01",
		X"0F",X"00",X"FE",X"08",X"3F",X"8C",X"13",X"CE",X"12",X"CE",X"13",X"CE",X"37",X"8C",X"7F",X"08",
		X"00",X"16",X"00",X"7B",X"01",X"F6",X"12",X"CF",X"13",X"8C",X"13",X"CB",X"13",X"FF",X"03",X"0F",
		X"ED",X"00",X"CA",X"00",X"0C",X"06",X"00",X"4E",X"00",X"4E",X"0F",X"C6",X"FF",X"CE",X"0F",X"0E",
		X"00",X"07",X"00",X"7F",X"01",X"ED",X"13",X"CA",X"13",X"8C",X"01",X"08",X"00",X"01",X"00",X"13",
		X"0F",X"00",X"FF",X"08",X"3D",X"8C",X"12",X"CE",X"01",X"CE",X"01",X"CE",X"1F",X"8C",X"FF",X"08",
		X"00",X"01",X"00",X"00",X"01",X"08",X"13",X"8C",X"13",X"8C",X"01",X"CF",X"00",X"7F",X"00",X"07",
		X"1F",X"8C",X"01",X"CE",X"00",X"6F",X"00",X"6F",X"01",X"E7",X"1E",X"CE",X"FF",X"8C",X"0F",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"13",X"00",X"37",X"00",X"6F",X"01",X"CE",
		X"03",X"08",X"37",X"08",X"7F",X"08",X"FF",X"08",X"BF",X"08",X"3F",X"08",X"37",X"08",X"37",X"08",
		X"13",X"8C",X"37",X"0F",X"37",X"FF",X"07",X"0F",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",
		X"37",X"08",X"3F",X"0C",X"FF",X"8C",X"3F",X"0C",X"37",X"08",X"7B",X"84",X"FF",X"CE",X"0F",X"0E",
		X"03",X"0F",X"13",X"FF",X"13",X"8F",X"13",X"8C",X"13",X"8C",X"13",X"8F",X"13",X"FB",X"13",X"ED",
		X"0F",X"0C",X"FF",X"8C",X"1E",X"8C",X"01",X"8C",X"00",X"0C",X"0E",X"00",X"FE",X"08",X"3F",X"8C",
		X"01",X"0C",X"00",X"00",X"03",X"08",X"13",X"8C",X"13",X"CA",X"01",X"ED",X"00",X"7F",X"00",X"07",
		X"13",X"CA",X"10",X"CE",X"01",X"CE",X"01",X"CE",X"13",X"CA",X"3F",X"84",X"EF",X"08",X"0E",X"00",
		X"00",X"07",X"00",X"7F",X"01",X"CF",X"12",X"8C",X"13",X"8C",X"13",X"8C",X"13",X"8F",X"13",X"FB",
		X"0F",X"00",X"FF",X"08",X"1F",X"8C",X"01",X"CA",X"01",X"CE",X"00",X"0C",X"0F",X"00",X"FF",X"08",
		X"13",X"ED",X"13",X"8E",X"13",X"8C",X"13",X"8C",X"12",X"CA",X"01",X"ED",X"00",X"7F",X"00",X"07",
		X"1F",X"8C",X"10",X"CE",X"01",X"CE",X"01",X"CE",X"03",X"CA",X"1F",X"8C",X"FF",X"08",X"0F",X"00",
		X"03",X"0F",X"13",X"FF",X"13",X"87",X"13",X"08",X"13",X"08",X"03",X"00",X"00",X"00",X"00",X"01",
		X"0F",X"0F",X"FF",X"EF",X"0F",X"6F",X"01",X"E7",X"12",X"CE",X"35",X"8C",X"7B",X"08",X"E7",X"00",
		X"00",X"01",X"00",X"12",X"00",X"13",X"00",X"13",X"00",X"13",X"00",X"13",X"00",X"13",X"00",X"03",
		X"CE",X"00",X"CA",X"00",X"8C",X"00",X"8C",X"00",X"8C",X"00",X"8C",X"00",X"8C",X"00",X"0C",X"00",
		X"00",X"07",X"00",X"7B",X"01",X"E7",X"01",X"CF",X"01",X"CE",X"01",X"ED",X"00",X"7F",X"00",X"37",
		X"0F",X"08",X"FF",X"84",X"3D",X"CA",X"12",X"CE",X"01",X"CE",X"01",X"CE",X"1E",X"CA",X"FF",X"84",
		X"00",X"7A",X"01",X"C7",X"12",X"8C",X"13",X"8C",X"13",X"CA",X"12",X"ED",X"01",X"F7",X"00",X"0F",
		X"F7",X"8C",X"3D",X"CE",X"03",X"E7",X"00",X"6F",X"00",X"6F",X"1E",X"ED",X"FF",X"CA",X"0F",X"0C",
		X"00",X"07",X"00",X"7F",X"01",X"CF",X"12",X"8E",X"13",X"8C",X"13",X"8C",X"13",X"C8",X"01",X"CF",
		X"0F",X"00",X"FF",X"08",X"3D",X"8C",X"12",X"CA",X"01",X"CE",X"01",X"CE",X"03",X"CE",X"3D",X"CE",
		X"00",X"7F",X"00",X"07",X"01",X"08",X"13",X"8C",X"12",X"8C",X"01",X"CF",X"00",X"7F",X"00",X"07",
		X"FE",X"CE",X"0F",X"CE",X"01",X"CE",X"01",X"CE",X"01",X"CA",X"1F",X"8C",X"FF",X"08",X"0F",X"00",
		X"00",X"0F",X"00",X"7F",X"00",X"35",X"00",X"36",X"00",X"6B",X"00",X"6D",X"00",X"4E",X"01",X"C6",
		X"0E",X"00",X"CE",X"00",X"ED",X"00",X"EF",X"00",X"E7",X"00",X"7E",X"08",X"7F",X"08",X"73",X"08",
		X"01",X"CB",X"01",X"FF",X"12",X"8F",X"13",X"84",X"13",X"08",X"35",X"84",X"37",X"CE",X"07",X"0E",
		X"3F",X"84",X"FF",X"8C",X"3D",X"8C",X"13",X"CA",X"13",X"CE",X"12",X"ED",X"37",X"EF",X"07",X"0F",
		X"07",X"0F",X"37",X"FF",X"12",X"ED",X"01",X"CE",X"01",X"CE",X"01",X"CE",X"01",X"CF",X"01",X"FF",
		X"01",X"CF",X"01",X"CE",X"01",X"CE",X"01",X"CE",X"01",X"CE",X"12",X"ED",X"37",X"FF",X"07",X"0F",
		X"3D",X"CA",X"03",X"ED",X"00",X"6F",X"00",X"6F",X"00",X"6F",X"0F",X"ED",X"FF",X"CA",X"0F",X"0C",
		X"0F",X"0E",X"FF",X"C6",X"3D",X"CE",X"12",X"CE",X"01",X"C6",X"00",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"27",X"00",X"6F",X"1E",X"CF",X"FF",X"8E",X"0F",X"0C",
		X"07",X"0F",X"37",X"FF",X"12",X"ED",X"01",X"CE",X"01",X"CE",X"01",X"CE",X"01",X"CE",X"01",X"CE",
		X"01",X"CE",X"01",X"CE",X"01",X"CE",X"01",X"CE",X"01",X"CE",X"12",X"ED",X"37",X"FF",X"07",X"0F",
		X"0F",X"0F",X"FF",X"EF",X"0F",X"6B",X"00",X"27",X"03",X"03",X"27",X"00",X"6B",X"00",X"EF",X"00",
		X"6B",X"00",X"27",X"00",X"03",X"00",X"00",X"03",X"00",X"27",X"0F",X"6B",X"FF",X"EF",X"0F",X"0F",
		X"6B",X"00",X"27",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"08",X"00",
		X"07",X"0F",X"37",X"EF",X"12",X"ED",X"01",X"CE",X"01",X"CE",X"1E",X"ED",X"FF",X"EF",X"0F",X"0F",
		X"0F",X"0F",X"7F",X"EF",X"35",X"CA",X"13",X"8C",X"13",X"8C",X"13",X"8C",X"1F",X"8C",X"FF",X"8C",
		X"1F",X"8C",X"13",X"8C",X"13",X"8C",X"13",X"8C",X"13",X"8C",X"35",X"CA",X"7F",X"EF",X"0F",X"0F",
		X"00",X"0F",X"00",X"7F",X"00",X"16",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",
		X"0F",X"0C",X"FF",X"8C",X"ED",X"08",X"CE",X"00",X"CE",X"00",X"CE",X"00",X"CE",X"00",X"CE",X"00",
		X"CE",X"00",X"CE",X"00",X"CE",X"00",X"CE",X"00",X"CE",X"00",X"ED",X"00",X"FF",X"8C",X"0F",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"7F",X"EF",X"35",X"CA",X"13",X"8C",X"13",X"8C",X"13",X"8C",X"13",X"8C",X"13",X"8C",
		X"00",X"00",X"00",X"00",X"03",X"08",X"13",X"8C",X"13",X"CA",X"01",X"ED",X"00",X"7F",X"00",X"07",
		X"13",X"8C",X"13",X"8C",X"13",X"8C",X"13",X"8C",X"35",X"8C",X"7B",X"84",X"FE",X"08",X"0F",X"00",
		X"0F",X"0F",X"3F",X"EF",X"12",X"CA",X"13",X"84",X"36",X"08",X"6D",X"00",X"CA",X"00",X"CE",X"00",
		X"ED",X"00",X"E7",X"00",X"7E",X"08",X"7B",X"08",X"37",X"84",X"35",X"CA",X"7F",X"EF",X"0F",X"0F",
		X"08",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"4E",X"00",X"4E",X"0F",X"C6",X"FF",X"CE",X"0F",X"0E",
		X"0F",X"08",X"7F",X"8C",X"37",X"CA",X"37",X"CE",X"36",X"ED",X"27",X"EF",X"27",X"F6",X"27",X"7F",
		X"00",X"0F",X"01",X"EF",X"12",X"CE",X"13",X"CE",X"35",X"CE",X"36",X"CE",X"6B",X"CE",X"6D",X"CE",
		X"27",X"7B",X"27",X"37",X"27",X"35",X"27",X"13",X"27",X"12",X"7A",X"09",X"7F",X"08",X"0F",X"08",
		X"C7",X"CE",X"C9",X"CE",X"8D",X"CE",X"81",X"CE",X"09",X"CE",X"12",X"ED",X"13",X"EF",X"03",X"0F",
		X"07",X"0E",X"37",X"ED",X"12",X"EF",X"01",X"FE",X"01",X"FB",X"01",X"BF",X"01",X"BD",X"01",X"9F",
		X"07",X"0F",X"37",X"EF",X"03",X"CA",X"09",X"8C",X"09",X"8C",X"85",X"8C",X"8D",X"8C",X"CB",X"8C",
		X"01",X"9E",X"01",X"8D",X"01",X"8D",X"01",X"8C",X"01",X"8C",X"12",X"CA",X"37",X"EF",X"07",X"0F",
		X"CF",X"8C",X"ED",X"8C",X"E7",X"8C",X"7E",X"8C",X"7B",X"8C",X"37",X"8C",X"35",X"8C",X"03",X"0C",
		X"0F",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"08",X"00",
		X"06",X"6F",X"6F",X"6F",X"37",X"E7",X"35",X"ED",X"12",X"CF",X"3D",X"ED",X"FF",X"E7",X"0F",X"0F",
		X"00",X"07",X"01",X"7B",X"12",X"ED",X"13",X"CA",X"13",X"CA",X"13",X"ED",X"01",X"FF",X"00",X"7B",
		X"0F",X"0E",X"FF",X"C6",X"3D",X"CE",X"12",X"CE",X"01",X"C6",X"08",X"0E",X"86",X"00",X"ED",X"08",
		X"00",X"16",X"00",X"01",X"03",X"08",X"13",X"84",X"13",X"CA",X"13",X"ED",X"13",X"F7",X"03",X"0F",
		X"FF",X"84",X"7B",X"CE",X"16",X"EF",X"01",X"E7",X"01",X"E7",X"1E",X"ED",X"FF",X"86",X"0F",X"08",
		X"03",X"0F",X"13",X"FF",X"13",X"96",X"13",X"09",X"03",X"01",X"00",X"01",X"00",X"01",X"00",X"01",
		X"0F",X"0F",X"FF",X"EF",X"ED",X"6B",X"CE",X"27",X"CE",X"03",X"CE",X"00",X"CE",X"00",X"CE",X"00",
		X"0F",X"0F",X"3F",X"EF",X"12",X"CA",X"01",X"8C",X"01",X"8C",X"01",X"8C",X"01",X"8C",X"01",X"8C",
		X"01",X"CE",X"01",X"CE",X"01",X"CE",X"01",X"CE",X"01",X"ED",X"01",X"F6",X"00",X"7B",X"00",X"07",
		X"01",X"8C",X"01",X"8C",X"01",X"8C",X"01",X"8C",X"12",X"8C",X"3D",X"84",X"FE",X"08",X"0F",X"00",
		X"0F",X"0F",X"7F",X"EF",X"35",X"CA",X"13",X"CA",X"12",X"CE",X"01",X"CE",X"01",X"ED",X"01",X"E7",
		X"07",X"0F",X"37",X"EF",X"12",X"CA",X"13",X"8C",X"13",X"84",X"13",X"08",X"35",X"08",X"36",X"08",
		X"00",X"6F",X"00",X"7E",X"00",X"7B",X"00",X"37",X"00",X"37",X"00",X"35",X"00",X"13",X"00",X"03",
		X"27",X"00",X"6B",X"00",X"6D",X"00",X"4E",X"00",X"C6",X"00",X"CA",X"00",X"8C",X"00",X"0C",X"00",
		X"0F",X"0B",X"7F",X"BF",X"7B",X"B5",X"37",X"1B",X"37",X"1B",X"37",X"1B",X"37",X"97",X"35",X"BD",
		X"0C",X"0F",X"CF",X"EF",X"CB",X"E5",X"8C",X"4E",X"8D",X"C6",X"8D",X"CE",X"CB",X"CA",X"DA",X"8C",
		X"13",X"BF",X"13",X"AF",X"13",X"EB",X"12",X"EF",X"01",X"ED",X"01",X"CE",X"01",X"CE",X"01",X"0E",
		X"DF",X"8C",X"DF",X"84",X"FD",X"08",X"F7",X"08",X"7E",X"08",X"6F",X"00",X"6F",X"00",X"0F",X"00",
		X"07",X"0F",X"37",X"EF",X"12",X"CE",X"01",X"ED",X"00",X"6F",X"00",X"7B",X"00",X"37",X"00",X"35",
		X"03",X"0F",X"13",X"EF",X"01",X"C6",X"12",X"8C",X"35",X"08",X"6B",X"00",X"C6",X"00",X"CA",X"00",
		X"00",X"13",X"00",X"35",X"00",X"6B",X"01",X"C6",X"12",X"8C",X"35",X"86",X"7F",X"EF",X"0F",X"0F",
		X"CE",X"00",X"ED",X"00",X"6F",X"00",X"7B",X"08",X"37",X"84",X"35",X"CA",X"7F",X"EF",X"0F",X"0F",
		X"03",X"0F",X"13",X"EF",X"01",X"C6",X"01",X"CA",X"12",X"8C",X"1B",X"84",X"B5",X"08",X"FA",X"08",
		X"00",X"13",X"00",X"12",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"12",X"00",X"37",X"00",X"07",
		X"EF",X"00",X"ED",X"00",X"CE",X"00",X"CE",X"00",X"CE",X"00",X"ED",X"00",X"FF",X"08",X"0F",X"08",
		X"0F",X"0E",X"FF",X"CE",X"0F",X"CE",X"01",X"CE",X"13",X"CA",X"37",X"84",X"7E",X"08",X"ED",X"00",
		X"00",X"13",X"00",X"37",X"00",X"7E",X"01",X"ED",X"12",X"CA",X"13",X"8F",X"13",X"FF",X"03",X"0F",
		X"CA",X"00",X"84",X"00",X"08",X"06",X"00",X"4E",X"00",X"4E",X"0F",X"C6",X"FF",X"CE",X"0F",X"0E",
		X"00",X"07",X"00",X"7F",X"01",X"ED",X"13",X"CA",X"13",X"8C",X"01",X"08",X"00",X"00",X"00",X"00",
		X"0F",X"00",X"FF",X"08",X"3D",X"8C",X"12",X"CE",X"12",X"CE",X"13",X"CA",X"37",X"84",X"7E",X"08",
		X"00",X"01",X"00",X"13",X"00",X"13",X"00",X"01",X"00",X"01",X"00",X"13",X"00",X"13",X"00",X"01",
		X"ED",X"00",X"CA",X"00",X"8C",X"00",X"08",X"00",X"08",X"00",X"8C",X"00",X"8C",X"00",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"0C",X"12",X"CA",X"13",X"CE",X"12",X"CA",X"01",X"0C",
		X"00",X"00",X"01",X"08",X"13",X"8C",X"13",X"8C",X"01",X"8C",X"01",X"8C",X"13",X"84",X"13",X"08",
		X"01",X"08",X"13",X"8C",X"13",X"8C",X"13",X"8C",X"13",X"8C",X"13",X"8C",X"13",X"8C",X"13",X"8C",
		X"13",X"8C",X"13",X"8C",X"12",X"8C",X"01",X"84",X"01",X"08",X"13",X"8C",X"13",X"8C",X"01",X"08",
		X"00",X"0E",X"07",X"4E",X"27",X"4F",X"27",X"F7",X"7B",X"ED",X"FE",X"4E",X"2F",X"4E",X"27",X"4E",
		X"27",X"4E",X"27",X"4F",X"27",X"F7",X"7B",X"ED",X"FE",X"4E",X"2F",X"4E",X"27",X"0E",X"07",X"00",
		X"01",X"0C",X"01",X"8C",X"74",X"F1",X"10",X"C0",X"01",X"0C",X"03",X"0E",X"02",X"02",X"66",X"33",
		X"01",X"0C",X"03",X"8E",X"74",X"F1",X"10",X"C0",X"01",X"84",X"12",X"C2",X"30",X"E0",X"01",X"04",
		X"0E",X"0E",X"0E",X"0E",X"0F",X"0E",X"27",X"8C",X"52",X"48",X"E1",X"E0",X"B4",X"A4",X"43",X"48",
		X"07",X"0C",X"0F",X"0E",X"3E",X"8E",X"5A",X"4A",X"79",X"C2",X"C3",X"68",X"D3",X"68",X"61",X"C0",
		X"07",X"0C",X"0F",X"86",X"78",X"C2",X"5E",X"8F",X"7E",X"CF",X"78",X"C3",X"69",X"C3",X"38",X"83",
		X"30",X"80",X"73",X"C8",X"97",X"2C",X"B5",X"A4",X"F6",X"EC",X"37",X"8C",X"43",X"48",X"33",X"88",
		X"C0",X"30",X"F4",X"F2",X"F7",X"FE",X"D7",X"BE",X"F7",X"FE",X"73",X"EC",X"63",X"6C",X"30",X"C0",
		X"09",X"02",X"1E",X"0E",X"28",X"C6",X"5A",X"CA",X"39",X"82",X"7A",X"42",X"24",X"84",X"03",X"08",
		X"30",X"80",X"73",X"C8",X"F7",X"EC",X"F7",X"EC",X"F7",X"EC",X"73",X"C8",X"30",X"80",X"00",X"00",
		X"60",X"C0",X"E4",X"E4",X"FE",X"EE",X"FF",X"EE",X"F7",X"EC",X"73",X"C8",X"31",X"80",X"10",X"00",
		X"E8",X"00",X"FB",X"C0",X"FB",X"FE",X"FB",X"E8",X"FB",X"80",X"F8",X"00",X"C8",X"00",X"C8",X"00",
		X"31",X"80",X"62",X"C8",X"62",X"C8",X"31",X"80",X"77",X"CC",X"31",X"00",X"31",X"00",X"31",X"00",
		X"24",X"48",X"24",X"48",X"F7",X"FE",X"E5",X"7F",X"F7",X"FE",X"24",X"48",X"24",X"48",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"08",X"FF",X"84",X"FF",X"CA",X"3D",X"ED",X"03",X"E7",X"00",X"6B",
		X"00",X"27",X"00",X"27",X"00",X"6B",X"03",X"E7",X"3D",X"ED",X"FF",X"CA",X"FF",X"84",X"0F",X"08",
		X"00",X"00",X"00",X"00",X"01",X"0F",X"12",X"FF",X"35",X"FF",X"7B",X"CB",X"7E",X"0C",X"6D",X"00",
		X"4E",X"00",X"4E",X"00",X"6D",X"00",X"7E",X"0C",X"7B",X"CB",X"35",X"FF",X"12",X"FF",X"01",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"13",X"08",X"1F",X"8C",
		X"FF",X"CE",X"FF",X"EF",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"4E",X"00",X"4E",X"00",X"6D",X"0F",
		X"7F",X"FF",X"7F",X"FF",X"6D",X"0F",X"4E",X"00",X"4E",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"08",X"13",X"8C",X"13",X"CE",X"01",X"E7",X"00",X"6B",X"08",X"27",
		X"08",X"27",X"8C",X"27",X"CF",X"6F",X"FE",X"ED",X"7F",X"CE",X"37",X"8C",X"03",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"08",X"7F",X"84",X"7F",X"CA",X"6D",X"ED",X"4E",X"6F",X"4E",X"7A",
		X"4E",X"37",X"4E",X"35",X"4E",X"12",X"4E",X"01",X"6D",X"08",X"7F",X"8C",X"0F",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"08",X"13",X"8C",X"13",X"CE",X"01",X"E7",X"08",X"6B",X"8C",X"27",
		X"8C",X"27",X"8C",X"27",X"8C",X"6B",X"CF",X"E7",X"7F",X"CE",X"37",X"8C",X"03",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"08",X"13",X"8C",X"37",X"8C",X"6F",X"08",X"4E",X"00",X"4E",X"01",
		X"4E",X"01",X"4E",X"01",X"4E",X"01",X"6D",X"13",X"7E",X"3F",X"37",X"EF",X"13",X"CE",X"01",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"8C",X"00",X"CE",X"00",X"6F",X"00",X"37",X"08",
		X"13",X"8C",X"0F",X"CE",X"FF",X"EF",X"FF",X"EF",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0E",X"00",X"6F",X"00",X"7F",X"00",X"5F",X"00",X"4F",X"00",X"4E",X"0C",X"4E",
		X"4E",X"4E",X"6D",X"4F",X"7F",X"FF",X"7F",X"FF",X"6D",X"4F",X"4E",X"0E",X"0C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"0F",X"FF",X"EF",X"FF",X"EF",X"CB",X"2F",X"C6",X"27",X"4E",X"27",
		X"4E",X"27",X"4E",X"27",X"CE",X"27",X"C8",X"6B",X"8D",X"EF",X"09",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"0C",X"13",X"8D",X"37",X"8D",X"7E",X"09",X"6D",X"00",X"4E",X"00",
		X"4E",X"00",X"4E",X"00",X"6F",X"01",X"37",X"3D",X"35",X"FF",X"12",X"FE",X"01",X"0F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"08",X"FF",X"84",X"FF",X"CE",X"87",X"6F",X"8C",X"27",X"8C",X"27",
		X"8C",X"27",X"8C",X"27",X"8C",X"27",X"8D",X"6F",X"1B",X"CE",X"13",X"84",X"01",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"0F",X"12",X"FF",X"37",X"FF",X"7E",X"1F",X"6D",X"12",X"4E",X"01",
		X"4E",X"01",X"4E",X"01",X"4F",X"01",X"6F",X"3D",X"37",X"FF",X"12",X"EF",X"01",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"0F",X"13",X"EF",X"01",X"6B",X"00",X"27",X"00",X"27",X"08",X"27",
		X"84",X"27",X"CA",X"27",X"ED",X"27",X"7E",X"2F",X"37",X"A7",X"13",X"EF",X"01",X"EF",X"00",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0E",X"7F",X"ED",
		X"7F",X"FF",X"0F",X"3D",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0C",X"37",X"CA",X"7F",X"ED",X"ED",X"6F",X"CE",X"2F",
		X"8C",X"27",X"8C",X"27",X"8C",X"6B",X"CB",X"E7",X"F7",X"ED",X"7B",X"CA",X"07",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"0C",X"35",X"CA",X"7B",X"ED",X"7E",X"3E",X"6D",X"13",X"4E",X"12",
		X"4E",X"12",X"4E",X"13",X"4E",X"35",X"6C",X"37",X"6F",X"7B",X"7B",X"EF",X"35",X"CE",X"03",X"0C",
		X"00",X"00",X"00",X"00",X"07",X"08",X"7F",X"84",X"FF",X"CE",X"CB",X"6F",X"08",X"2F",X"08",X"27",
		X"08",X"27",X"08",X"27",X"84",X"6B",X"8F",X"E7",X"FF",X"CE",X"FF",X"84",X"0F",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"08",X"12",X"8C",X"37",X"8D",X"6F",X"1B",X"4E",X"13",X"4E",X"13",
		X"4E",X"13",X"4E",X"13",X"4E",X"13",X"6F",X"1E",X"37",X"FF",X"12",X"FF",X"01",X"0F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"87",X"03",X"FE",X"2F",X"3D",X"EB",X"03",X"E7",
		X"16",X"EF",X"F7",X"EF",X"FF",X"CB",X"ED",X"0C",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0E",X"00",X"6D",X"0C",X"7F",X"CB",X"6D",X"F7",X"4E",X"3E",X"0C",X"27",X"00",X"27",
		X"00",X"27",X"0C",X"27",X"4F",X"7B",X"7D",X"FF",X"7F",X"FE",X"7F",X"87",X"6D",X"08",X"0E",X"00",
		X"00",X"00",X"00",X"03",X"00",X"27",X"0F",X"6B",X"FF",X"EF",X"FF",X"EF",X"8F",X"6B",X"8C",X"27",
		X"00",X"00",X"0C",X"00",X"4E",X"00",X"6D",X"0F",X"7F",X"FF",X"7F",X"FF",X"6D",X"0F",X"4E",X"01",
		X"4E",X"01",X"4E",X"01",X"4E",X"12",X"4E",X"13",X"6F",X"3F",X"7B",X"FE",X"35",X"ED",X"03",X"0E",
		X"00",X"27",X"00",X"27",X"00",X"6B",X"01",X"E7",X"12",X"ED",X"13",X"EF",X"03",X"0F",X"00",X"00",
		X"4E",X"00",X"4E",X"00",X"4E",X"00",X"6C",X"00",X"6F",X"00",X"3F",X"08",X"17",X"8C",X"03",X"08",
		X"00",X"00",X"00",X"03",X"00",X"27",X"0F",X"6B",X"FF",X"EF",X"FF",X"EF",X"0F",X"6B",X"00",X"27",
		X"00",X"00",X"0C",X"00",X"4E",X"00",X"6D",X"0F",X"7F",X"FF",X"7F",X"FF",X"6D",X"0F",X"4E",X"00",
		X"8C",X"27",X"CA",X"27",X"EF",X"27",X"0F",X"27",X"00",X"27",X"00",X"6B",X"01",X"EF",X"01",X"0F",
		X"4E",X"01",X"4E",X"12",X"4E",X"37",X"4E",X"07",X"4E",X"00",X"6D",X"00",X"7F",X"08",X"0F",X"08",
		X"0C",X"01",X"00",X"12",X"00",X"37",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"4E",X"00",X"4E",X"03",X"4E",X"27",X"6D",X"6B",X"7F",X"EF",X"7F",X"EF",X"6D",X"6B",X"0E",X"07",
		X"8C",X"03",X"8C",X"27",X"8F",X"6B",X"FF",X"EF",X"FF",X"EF",X"0F",X"6B",X"00",X"27",X"00",X"03",
		X"0C",X"01",X"4E",X"01",X"6D",X"0F",X"7F",X"FF",X"7F",X"FF",X"6D",X"0F",X"4E",X"00",X"0C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"27",X"00",X"27",X"0F",X"6B",
		X"FF",X"EF",X"FF",X"EF",X"0F",X"6B",X"00",X"27",X"00",X"27",X"00",X"03",X"00",X"00",X"00",X"00",
		X"7F",X"FF",X"7F",X"FF",X"6D",X"0F",X"4E",X"00",X"4C",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"00",X"27",X"0F",X"6B",X"FF",X"EF",X"FF",X"EF",X"0F",X"6B",X"00",X"27",X"00",X"03",
		X"00",X"00",X"00",X"00",X"01",X"0C",X"13",X"8C",X"37",X"8C",X"7E",X"08",X"6D",X"00",X"4E",X"00",
		X"4E",X"00",X"6D",X"00",X"7E",X"0F",X"7B",X"FF",X"35",X"FF",X"03",X"0F",X"00",X"00",X"00",X"00",
		X"CE",X"03",X"EB",X"03",X"3D",X"2F",X"12",X"EB",X"01",X"E7",X"00",X"6B",X"00",X"27",X"00",X"03",
		X"0C",X"3D",X"4F",X"F7",X"7D",X"FE",X"7F",X"CB",X"7E",X"0C",X"6D",X"00",X"4E",X"00",X"0C",X"00",
		X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"4E",X"00",X"4E",X"00",X"4E",X"00",X"4E",X"00",X"6D",X"08",X"7F",X"8C",X"0F",X"0C",X"00",X"00",
		X"00",X"03",X"0F",X"2F",X"FF",X"EF",X"1E",X"EF",X"7B",X"EF",X"FF",X"CA",X"FE",X"0C",X"CB",X"00",
		X"0C",X"00",X"CB",X"00",X"F6",X"0C",X"3D",X"CA",X"FF",X"EF",X"FF",X"EF",X"0F",X"2F",X"00",X"03",
		X"0E",X"00",X"6D",X"0F",X"7F",X"FF",X"6D",X"0F",X"0E",X"01",X"00",X"16",X"01",X"7B",X"12",X"FF",
		X"01",X"F6",X"00",X"35",X"0E",X"01",X"6D",X"0F",X"7F",X"FF",X"7F",X"FF",X"6D",X"0F",X"0E",X"00",
		X"00",X"00",X"00",X"03",X"00",X"27",X"0F",X"6B",X"FF",X"EF",X"1E",X"EF",X"7B",X"ED",X"FF",X"86",
		X"ED",X"08",X"86",X"03",X"08",X"27",X"0F",X"2F",X"FF",X"EF",X"0F",X"6B",X"00",X"27",X"00",X"03",
		X"00",X"00",X"0C",X"00",X"4E",X"00",X"6D",X"0F",X"7F",X"FF",X"6D",X"0F",X"4E",X"01",X"0C",X"16",
		X"01",X"7B",X"16",X"FF",X"7B",X"ED",X"7F",X"87",X"7F",X"FF",X"0F",X"0F",X"00",X"00",X"00",X"00",
		X"0C",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"4E",X"02",X"4E",X"2F",X"6D",X"E7",X"7E",X"CE",X"7B",X"CB",X"7F",X"FF",X"6D",X"F7",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"03",X"0C",X"37",X"CA",X"7F",X"CE",X"F6",X"E5",X"ED",X"6B",X"CE",X"27",
		X"CA",X"27",X"8C",X"27",X"84",X"6B",X"09",X"E7",X"1A",X"ED",X"13",X"EF",X"03",X"0F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"0C",X"7F",X"8C",X"7B",X"84",X"7E",X"09",X"6D",X"01",X"4E",X"12",
		X"4E",X"13",X"4E",X"35",X"4E",X"37",X"6D",X"7B",X"7A",X"F6",X"37",X"EF",X"35",X"CE",X"03",X"0C",
		X"00",X"00",X"00",X"00",X"01",X"0F",X"01",X"EF",X"00",X"6B",X"00",X"27",X"00",X"27",X"0F",X"6B",
		X"FF",X"EF",X"FF",X"EF",X"0F",X"6B",X"00",X"27",X"00",X"27",X"00",X"6B",X"01",X"EF",X"01",X"0F",
		X"00",X"03",X"00",X"03",X"00",X"27",X"0F",X"6B",X"FF",X"EF",X"0F",X"6B",X"00",X"27",X"00",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0F",X"35",X"FF",X"7B",X"FF",X"7E",X"0F",X"6D",X"00",
		X"4E",X"00",X"4E",X"00",X"6D",X"00",X"7A",X"0F",X"35",X"FF",X"03",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"03",X"00",X"27",X"01",X"6B",X"1E",X"EF",X"F7",X"EF",X"FF",X"E3",X"CB",X"2F",X"0C",X"03",
		X"00",X"00",X"0C",X"03",X"CB",X"2F",X"F7",X"EB",X"1E",X"EF",X"01",X"6B",X"00",X"27",X"00",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"03",X"7B",X"3D",X"FF",X"7F",X"ED",
		X"7E",X"0E",X"3D",X"ED",X"03",X"7B",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"0F",X"6B",X"F7",X"EF",X"FF",X"EF",X"CB",X"6B",X"0C",X"06",X"87",X"6B",X"FF",X"EF",
		X"FF",X"EF",X"C3",X"6B",X"0C",X"06",X"87",X"06",X"FE",X"6B",X"7B",X"EF",X"07",X"6B",X"00",X"07",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"F7",X"7F",X"FF",X"7F",X"CB",X"1E",X"FF",X"01",X"1F",
		X"0F",X"F7",X"7F",X"FF",X"7F",X"CB",X"1E",X"FF",X"01",X"3D",X"00",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"00",X"27",X"00",X"6B",X"03",X"EF",X"3D",X"EF",X"F7",X"A7",X"EF",X"0B",
		X"CA",X"00",X"E5",X"00",X"3E",X"0B",X"13",X"A7",X"01",X"EB",X"00",X"6F",X"00",X"27",X"00",X"03",
		X"0C",X"00",X"4E",X"00",X"6D",X"00",X"7E",X"08",X"7D",X"84",X"4F",X"CA",X"4E",X"6D",X"0C",X"37",
		X"0C",X"3F",X"4F",X"F7",X"7D",X"ED",X"7F",X"8E",X"7E",X"08",X"6D",X"00",X"4E",X"00",X"0C",X"00",
		X"CA",X"00",X"84",X"00",X"CB",X"03",X"F6",X"2F",X"3D",X"EB",X"03",X"E7",X"00",X"2F",X"00",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"4E",X"03",X"6D",X"3D",
		X"7F",X"FF",X"7F",X"FF",X"6D",X"3D",X"4E",X"03",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"8C",X"27",X"CE",X"27",X"E7",X"27",X"7B",X"2F",X"35",X"EF",X"12",X"EF",X"01",X"0F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"00",X"7E",X"08",X"7F",X"8C",X"5E",X"CE",X"4F",X"E7",X"4E",X"7B",
		X"4E",X"35",X"4E",X"12",X"4E",X"01",X"4E",X"00",X"6D",X"08",X"7F",X"8C",X"0F",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"08",X"13",X"8C",X"13",X"CE",X"01",X"E7",X"00",X"6B",X"00",X"27",
		X"08",X"27",X"8C",X"27",X"CF",X"6B",X"F6",X"E7",X"7B",X"CE",X"35",X"8C",X"03",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"6F",X"6F",
		X"6F",X"7F",X"06",X"35",X"00",X"12",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"00",X"7A",X"08",X"7F",X"08",X"7A",X"08",X"07",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"0C",X"CF",X"CE",X"7B",X"CE",X"07",X"0C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"0E",X"FF",X"EF",X"FF",X"EF",X"0F",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"07",X"6F",X"7B",X"6F",X"F7",X"06",X"0F",X"00",X"00",X"00",X"00",
		X"27",X"00",X"3E",X"0E",X"FF",X"CE",X"3D",X"0E",X"1F",X"87",X"FF",X"EF",X"1E",X"8F",X"01",X"8C",
		X"13",X"08",X"1F",X"87",X"7F",X"FF",X"1E",X"8F",X"07",X"CB",X"37",X"FF",X"07",X"C7",X"00",X"4E",
		X"00",X"00",X"88",X"44",X"8E",X"40",X"03",X"C3",X"03",X"E3",X"03",X"C3",X"8E",X"40",X"88",X"44",
		X"00",X"00",X"00",X"44",X"42",X"42",X"69",X"C3",X"70",X"E3",X"69",X"C3",X"42",X"42",X"00",X"44",
		X"60",X"07",X"B4",X"0F",X"69",X"8F",X"5A",X"0C",X"69",X"8F",X"B4",X"0F",X"60",X"07",X"00",X"00",
		X"61",X"0E",X"F0",X"87",X"96",X"4F",X"5F",X"C3",X"96",X"4F",X"F0",X"87",X"61",X"0E",X"00",X"00",
		X"0F",X"0E",X"71",X"CB",X"F1",X"4B",X"B4",X"C3",X"F1",X"E9",X"71",X"4B",X"0F",X"0E",X"0F",X"08",
		X"10",X"C0",X"53",X"2C",X"BF",X"B6",X"BE",X"FE",X"BF",X"B6",X"53",X"2C",X"10",X"C0",X"00",X"00",
		X"10",X"F0",X"71",X"FE",X"F7",X"6C",X"B7",X"EC",X"B7",X"EC",X"F7",X"6C",X"71",X"FE",X"10",X"F0",
		X"03",X"0F",X"24",X"82",X"7A",X"4A",X"39",X"A1",X"58",X"CA",X"24",X"C6",X"03",X"0F",X"00",X"00",
		X"31",X"80",X"33",X"88",X"33",X"88",X"33",X"88",X"73",X"C8",X"77",X"CC",X"55",X"44",X"00",X"00",
		X"10",X"EC",X"31",X"FE",X"73",X"FC",X"F7",X"C8",X"73",X"FC",X"31",X"FE",X"10",X"EC",X"00",X"00",
		X"FF",X"FF",X"F0",X"F0",X"31",X"FE",X"31",X"EE",X"10",X"EC",X"00",X"E4",X"00",X"C4",X"00",X"40",
		X"00",X"00",X"11",X"60",X"F1",X"F6",X"FF",X"99",X"11",X"F6",X"11",X"60",X"00",X"00",X"00",X"00",
		X"00",X"31",X"00",X"72",X"00",X"E4",X"34",X"C8",X"13",X"00",X"43",X"80",X"84",X"08",X"08",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		if addr(13) = '1' then
			data <= (others=>'0');
		else
			data <= rom_data(to_integer(unsigned(addr)));
		end if;
	end if;
end process;
end architecture;
