library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity kick_sp_bits_2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of kick_sp_bits_2 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"0E",X"0E",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"22",X"00",
		X"E0",X"00",X"22",X"00",X"E0",X"00",X"22",X"00",X"EE",X"00",X"22",X"0E",X"EE",X"00",X"00",X"EE",
		X"0E",X"00",X"00",X"EE",X"0E",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",
		X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"E0",X"0E",X"00",X"00",X"EE",X"EE",X"00",
		X"00",X"EE",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",
		X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"D0",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"E0",X"00",
		X"00",X"EE",X"EE",X"00",X"00",X"E0",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"0E",X"00",X"00",X"EE",X"0E",X"00",X"00",X"EE",
		X"EE",X"00",X"00",X"EE",X"EE",X"22",X"00",X"0E",X"E0",X"22",X"00",X"00",X"E0",X"22",X"00",X"00",
		X"E0",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"0E",X"0E",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"00",X"00",X"EE",X"EE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"E0",X"00",
		X"00",X"EE",X"EE",X"00",X"00",X"E0",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"0E",X"00",X"00",X"EE",X"0E",X"00",X"00",X"EE",
		X"EE",X"00",X"00",X"EE",X"EE",X"00",X"00",X"0E",X"E0",X"00",X"00",X"00",X"E0",X"00",X"88",X"00",
		X"70",X"00",X"88",X"00",X"75",X"00",X"88",X"00",X"05",X"E0",X"88",X"00",X"00",X"0E",X"8E",X"00",
		X"50",X"00",X"E0",X"00",X"50",X"00",X"22",X"00",X"55",X"EE",X"22",X"00",X"E5",X"EE",X"EE",X"EE",
		X"FF",X"34",X"77",X"77",X"FF",X"34",X"77",X"77",X"55",X"34",X"77",X"77",X"55",X"44",X"77",X"77",
		X"55",X"44",X"77",X"77",X"04",X"44",X"77",X"77",X"04",X"44",X"77",X"77",X"04",X"44",X"77",X"77",
		X"00",X"44",X"77",X"77",X"00",X"44",X"07",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"33",X"77",X"22",X"55",X"33",X"77",X"22",X"55",X"33",X"77",X"23",X"FF",X"33",X"77",X"23",
		X"55",X"33",X"77",X"23",X"54",X"33",X"77",X"23",X"54",X"03",X"77",X"23",X"04",X"03",X"77",X"20",
		X"04",X"00",X"BB",X"00",X"04",X"00",X"B7",X"00",X"00",X"44",X"B0",X"00",X"00",X"44",X"BB",X"00",
		X"00",X"44",X"5B",X"00",X"00",X"44",X"5B",X"00",X"00",X"44",X"BB",X"00",X"00",X"00",X"B0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"33",X"77",X"77",X"55",X"33",X"77",X"77",X"FF",X"33",X"77",X"77",X"55",X"33",X"77",X"77",
		X"55",X"33",X"B7",X"77",X"54",X"33",X"B7",X"20",X"54",X"33",X"77",X"20",X"04",X"35",X"77",X"20",
		X"04",X"04",X"77",X"00",X"00",X"44",X"07",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"44",X"BB",X"00",X"00",X"44",X"BB",X"00",X"00",X"44",X"BB",
		X"00",X"00",X"44",X"AB",X"00",X"00",X"04",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"AA",
		X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"04",X"6B",X"00",X"00",X"44",X"BB",X"00",X"00",X"44",X"B7",X"00",X"00",X"44",X"7B",
		X"00",X"00",X"44",X"BB",X"00",X"00",X"04",X"BB",X"00",X"00",X"00",X"BA",X"00",X"00",X"00",X"AA",
		X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BA",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"6B",X"00",X"00",X"00",X"BB",X"00",X"00",X"04",X"BB",
		X"00",X"00",X"44",X"BB",X"00",X"00",X"44",X"AB",X"00",X"00",X"44",X"BB",X"00",X"00",X"44",X"AB",
		X"00",X"00",X"04",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"01",X"11",
		X"00",X"00",X"01",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"01",X"00",X"00",X"77",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"70",X"40",X"53",X"77",X"77",X"44",X"55",X"77",X"77",
		X"44",X"33",X"77",X"77",X"44",X"33",X"77",X"77",X"44",X"33",X"77",X"77",X"55",X"33",X"77",X"77",
		X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",
		X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"77",X"00",X"00",X"DD",X"77",X"00",X"00",X"D0",X"77",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",
		X"00",X"0B",X"00",X"77",X"00",X"0B",X"00",X"77",X"00",X"0B",X"00",X"77",X"00",X"B0",X"00",X"77",
		X"00",X"B0",X"00",X"77",X"00",X"BB",X"00",X"77",X"00",X"BB",X"00",X"77",X"00",X"BB",X"00",X"77",
		X"0B",X"BB",X"00",X"77",X"0B",X"55",X"00",X"77",X"00",X"55",X"00",X"77",X"00",X"55",X"00",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"0E",X"0E",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",
		X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"0E",X"EE",X"00",X"00",X"EE",
		X"0E",X"00",X"00",X"EE",X"0E",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"0E",X"00",X"00",X"EE",X"EE",X"00",
		X"00",X"EE",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F5",X"EE",X"0D",X"00",X"EE",X"EE",X"DD",X"00",X"77",X"77",X"DD",X"00",X"77",X"75",X"0E",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",
		X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"EE",X"EE",X"00",X"00",X"0E",
		X"0E",X"00",X"00",X"EE",X"0E",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"0E",X"00",X"00",X"EE",X"EE",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"EE",X"EE",X"EE",X"77",X"EE",X"00",X"00",X"77",X"0E",X"E0",X"00",X"77",X"E0",X"E0",X"00",
		X"00",X"08",X"0E",X"00",X"00",X"08",X"0E",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",
		X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"0E",X"EE",X"00",X"00",X"0E",
		X"0E",X"0E",X"00",X"EE",X"0E",X"0E",X"00",X"EE",X"00",X"0E",X"00",X"E0",X"00",X"0E",X"00",X"00",
		X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"0E",X"00",X"00",X"EE",X"EE",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",
		X"00",X"B0",X"00",X"77",X"00",X"BB",X"00",X"77",X"00",X"BB",X"00",X"77",X"00",X"BB",X"00",X"77",
		X"00",X"FF",X"07",X"77",X"00",X"5F",X"07",X"77",X"00",X"5F",X"07",X"07",X"00",X"F5",X"07",X"00",
		X"00",X"44",X"77",X"00",X"50",X"44",X"77",X"00",X"50",X"44",X"77",X"21",X"55",X"44",X"77",X"21",
		X"FF",X"34",X"77",X"71",X"55",X"34",X"77",X"71",X"55",X"44",X"77",X"72",X"FF",X"44",X"77",X"72",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"B0",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"5B",X"00",X"00",X"B0",X"5B",X"00",X"00",X"B0",X"F0",X"00",
		X"00",X"B0",X"F0",X"01",X"00",X"B0",X"00",X"01",X"00",X"BB",X"07",X"11",X"00",X"BB",X"77",X"11",
		X"00",X"BB",X"77",X"11",X"50",X"BB",X"77",X"11",X"50",X"BB",X"77",X"11",X"55",X"3B",X"77",X"11",
		X"FF",X"35",X"77",X"77",X"55",X"35",X"77",X"77",X"55",X"35",X"77",X"77",X"FF",X"33",X"77",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"B0",X"00",X"00",
		X"0B",X"B0",X"00",X"10",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",
		X"00",X"50",X"00",X"11",X"00",X"F5",X"00",X"11",X"00",X"44",X"01",X"11",X"00",X"44",X"01",X"11",
		X"00",X"44",X"11",X"11",X"00",X"44",X"11",X"11",X"00",X"44",X"77",X"10",X"00",X"45",X"77",X"10",
		X"00",X"55",X"77",X"70",X"50",X"33",X"77",X"77",X"50",X"33",X"77",X"77",X"55",X"33",X"77",X"77",
		X"FF",X"33",X"77",X"77",X"55",X"33",X"77",X"77",X"55",X"33",X"77",X"77",X"FF",X"33",X"77",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"F5",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"07",X"00",X"44",X"00",X"77",X"00",X"44",X"00",X"77",
		X"00",X"44",X"00",X"77",X"00",X"45",X"00",X"77",X"00",X"55",X"77",X"77",X"00",X"33",X"77",X"77",
		X"00",X"33",X"77",X"77",X"50",X"33",X"77",X"77",X"50",X"33",X"77",X"77",X"55",X"33",X"77",X"77",
		X"FF",X"33",X"77",X"77",X"FF",X"33",X"77",X"77",X"55",X"33",X"77",X"77",X"55",X"33",X"77",X"77",
		X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",
		X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"D0",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0B",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"5B",X"00",
		X"00",X"00",X"5B",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"50",X"07",X"00",X"00",X"00",X"07",
		X"00",X"44",X"00",X"77",X"00",X"44",X"00",X"77",X"00",X"44",X"00",X"77",X"04",X"44",X"00",X"77",
		X"44",X"44",X"00",X"77",X"44",X"44",X"00",X"77",X"54",X"40",X"07",X"77",X"F4",X"00",X"77",X"77",
		X"54",X"00",X"77",X"77",X"55",X"33",X"77",X"77",X"F3",X"35",X"77",X"77",X"53",X"55",X"77",X"77",
		X"53",X"55",X"77",X"77",X"F3",X"35",X"77",X"72",X"55",X"33",X"77",X"22",X"54",X"00",X"77",X"22",
		X"F4",X"00",X"77",X"22",X"54",X"40",X"07",X"22",X"44",X"44",X"07",X"11",X"44",X"44",X"00",X"11",
		X"04",X"44",X"00",X"11",X"00",X"44",X"00",X"11",X"00",X"44",X"00",X"11",X"00",X"44",X"00",X"01",
		X"00",X"04",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"04",X"00",X"00",X"00",X"54",X"00",X"00",
		X"BB",X"FF",X"00",X"11",X"0B",X"55",X"00",X"11",X"0B",X"FF",X"00",X"11",X"00",X"54",X"00",X"11",
		X"00",X"50",X"00",X"11",X"00",X"00",X"00",X"10",X"00",X"00",X"F1",X"00",X"00",X"00",X"51",X"00",
		X"00",X"00",X"5F",X"0D",X"00",X"00",X"FF",X"DD",X"00",X"00",X"F5",X"DD",X"00",X"00",X"BD",X"DD",
		X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",
		X"77",X"77",X"BD",X"00",X"77",X"77",X"BD",X"00",X"77",X"EE",X"DD",X"00",X"77",X"00",X"DD",X"E0",
		X"00",X"00",X"0D",X"EE",X"00",X"0E",X"00",X"00",X"0E",X"0E",X"E0",X"00",X"E0",X"E0",X"E0",X"00",
		X"E0",X"E0",X"0E",X"00",X"E0",X"00",X"0E",X"00",X"EE",X"00",X"00",X"0E",X"EE",X"00",X"00",X"0E",
		X"0E",X"00",X"00",X"EE",X"0E",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"0E",X"00",X"00",X"EE",X"EE",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"BB",X"00",X"00",X"EE",X"BD",X"00",X"00",X"33",X"BD",X"E0",X"00",X"33",X"DD",X"0E",X"00",
		X"33",X"DD",X"00",X"00",X"30",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",
		X"E0",X"00",X"00",X"E0",X"E0",X"00",X"00",X"0E",X"EE",X"00",X"00",X"0E",X"EE",X"00",X"00",X"0E",
		X"0E",X"00",X"00",X"EE",X"0E",X"00",X"E0",X"EE",X"00",X"00",X"E0",X"E0",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"E0",X"0E",X"00",X"00",X"EE",X"EE",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"EE",X"EE",X"00",X"00",X"E0",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",
		X"00",X"00",X"E0",X"00",X"70",X"00",X"E0",X"E0",X"7E",X"08",X"E0",X"EE",X"7E",X"08",X"00",X"EE",
		X"77",X"08",X"80",X"0E",X"77",X"00",X"82",X"0E",X"77",X"00",X"82",X"0E",X"77",X"00",X"82",X"E0",
		X"77",X"00",X"82",X"00",X"77",X"00",X"88",X"00",X"77",X"E0",X"88",X"00",X"77",X"5E",X"58",X"00",
		X"77",X"5E",X"3E",X"00",X"77",X"F5",X"D0",X"00",X"77",X"F5",X"D0",X"00",X"37",X"BB",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"EE",X"EE",X"00",X"00",X"E0",X"0E",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"E0",X"0E",X"0E",X"00",X"EE",X"3E",X"0D",X"00",X"EE",
		X"EE",X"0D",X"00",X"0E",X"EE",X"0D",X"00",X"0E",X"E7",X"0D",X"22",X"00",X"E7",X"0D",X"22",X"00",
		X"E7",X"00",X"22",X"00",X"77",X"00",X"22",X"00",X"77",X"00",X"DD",X"00",X"77",X"00",X"DD",X"00",
		X"77",X"E0",X"DD",X"00",X"77",X"77",X"E0",X"00",X"77",X"77",X"88",X"00",X"77",X"77",X"88",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"EE",X"EE",X"00",X"00",X"E0",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"0E",X"00",X"00",X"EE",X"0E",X"00",X"00",X"EE",
		X"EE",X"00",X"00",X"0E",X"EE",X"00",X"00",X"0E",X"E0",X"80",X"0D",X"00",X"E0",X"E8",X"DD",X"00",
		X"E0",X"E8",X"DD",X"00",X"7E",X"8E",X"DD",X"00",X"70",X"8E",X"DD",X"00",X"77",X"88",X"DD",X"EE",
		X"77",X"80",X"DD",X"E0",X"77",X"EE",X"DD",X"00",X"77",X"77",X"BD",X"00",X"77",X"77",X"BD",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",
		X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",
		X"00",X"00",X"B0",X"44",X"00",X"00",X"BB",X"44",X"00",X"00",X"BB",X"44",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"44",X"AA",X"00",X"00",X"44",X"BB",X"00",X"00",X"04",X"BB",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"0B",X"B0",
		X"00",X"00",X"0B",X"B0",X"00",X"00",X"4B",X"B0",X"00",X"04",X"4B",X"B0",X"00",X"04",X"4A",X"A5",
		X"53",X"57",X"77",X"7F",X"F3",X"37",X"77",X"75",X"53",X"37",X"77",X"75",X"53",X"37",X"77",X"7F",
		X"F3",X"37",X"77",X"75",X"50",X"07",X"72",X"05",X"40",X"07",X"72",X"00",X"40",X"07",X"72",X"00",
		X"40",X"07",X"70",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"40",X"00",X"00",X"04",X"40",X"00",X"00",
		X"04",X"40",X"00",X"00",X"04",X"40",X"00",X"00",X"04",X"40",X"00",X"00",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"0B",X"B0",X"00",X"00",X"0B",
		X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"0B",X"B0",X"00",X"00",X"0B",
		X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",
		X"BB",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",
		X"BB",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",
		X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"77",X"00",
		X"04",X"00",X"77",X"20",X"54",X"00",X"77",X"20",X"55",X"00",X"77",X"20",X"FF",X"33",X"77",X"77",
		X"55",X"33",X"77",X"77",X"55",X"33",X"77",X"77",X"FF",X"33",X"77",X"77",X"55",X"35",X"77",X"77",
		X"55",X"44",X"77",X"22",X"55",X"44",X"77",X"22",X"FF",X"44",X"77",X"21",X"55",X"44",X"77",X"21",
		X"55",X"43",X"77",X"21",X"54",X"33",X"77",X"21",X"54",X"33",X"77",X"20",X"04",X"33",X"77",X"20",
		X"00",X"04",X"77",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"04",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"40",X"00",X"44",X"44",X"40",X"00",X"44",X"44",X"40",X"00",X"44",X"44",X"40",
		X"00",X"44",X"44",X"40",X"00",X"44",X"44",X"40",X"00",X"44",X"44",X"40",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"04",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"00",X"77",X"00",X"44",X"00",X"77",X"00",X"44",X"03",X"77",X"00",X"44",X"33",X"77",
		X"00",X"44",X"33",X"77",X"00",X"44",X"33",X"77",X"00",X"44",X"33",X"77",X"00",X"44",X"33",X"77",
		X"00",X"44",X"33",X"70",X"00",X"44",X"33",X"00",X"00",X"44",X"53",X"00",X"00",X"44",X"33",X"00",
		X"00",X"43",X"53",X"00",X"00",X"33",X"33",X"00",X"00",X"33",X"33",X"00",X"00",X"33",X"33",X"00",
		X"00",X"33",X"33",X"00",X"00",X"33",X"33",X"00",X"00",X"33",X"30",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"AB",X"00",X"00",X"00",X"AB",X"44",X"44",X"BB",X"BB",X"44",X"44",X"BB",X"BB",X"44",X"44",
		X"BB",X"BB",X"44",X"44",X"4B",X"BB",X"44",X"40",X"44",X"BB",X"44",X"00",X"44",X"BB",X"44",X"00",
		X"44",X"AA",X"00",X"00",X"44",X"AA",X"00",X"00",X"44",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",
		X"77",X"70",X"DD",X"0E",X"77",X"00",X"DD",X"EE",X"77",X"00",X"DD",X"EE",X"77",X"00",X"DD",X"E0",
		X"77",X"00",X"DD",X"E0",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",
		X"77",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"0E",X"EE",X"00",
		X"0E",X"E0",X"EE",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",
		X"55",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"55",X"BB",X"00",X"00",X"55",X"00",X"00",X"00",
		X"FF",X"BB",X"00",X"00",X"5B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"E0",X"00",X"EE",X"00",X"EE",X"00",X"E0",X"00",X"EE",
		X"00",X"E0",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",
		X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",
		X"E0",X"E0",X"00",X"00",X"E0",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"0E",X"00",
		X"00",X"DD",X"0E",X"00",X"00",X"FD",X"E0",X"00",X"77",X"FD",X"D0",X"00",X"77",X"F5",X"DD",X"EE",
		X"33",X"33",X"00",X"BB",X"33",X"44",X"00",X"BB",X"33",X"44",X"44",X"BB",X"33",X"44",X"44",X"BB",
		X"33",X"44",X"44",X"BB",X"33",X"44",X"44",X"5B",X"03",X"44",X"40",X"0B",X"03",X"54",X"E0",X"00",
		X"00",X"F5",X"0E",X"00",X"00",X"5F",X"00",X"00",X"00",X"F5",X"00",X"0E",X"AA",X"55",X"00",X"0E",
		X"AA",X"BB",X"00",X"EE",X"AA",X"AB",X"00",X"EE",X"AA",X"AA",X"00",X"E0",X"AA",X"BA",X"00",X"E0",
		X"0B",X"BB",X"00",X"00",X"0B",X"AB",X"4E",X"00",X"0B",X"AB",X"44",X"00",X"0B",X"6B",X"44",X"00",
		X"0B",X"60",X"44",X"BB",X"0B",X"BA",X"44",X"BB",X"0B",X"AA",X"44",X"B0",X"00",X"0A",X"44",X"BB",
		X"00",X"00",X"04",X"BB",X"00",X"04",X"00",X"B0",X"00",X"44",X"00",X"BB",X"00",X"44",X"00",X"0B",
		X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",
		X"00",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"50",X"00",X"00",
		X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"77",X"00",
		X"00",X"EE",X"77",X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"7E",X"70",
		X"00",X"00",X"7E",X"70",X"00",X"77",X"E7",X"70",X"00",X"77",X"E7",X"00",X"00",X"77",X"77",X"00",
		X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"77",X"77",X"77",X"00",X"77",X"77",X"00",X"00",
		X"77",X"77",X"00",X"E0",X"77",X"77",X"00",X"E0",X"77",X"77",X"00",X"E0",X"77",X"77",X"00",X"EE",
		X"33",X"77",X"00",X"EE",X"33",X"37",X"00",X"EE",X"33",X"33",X"EE",X"EB",X"33",X"33",X"00",X"BE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"04",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"04",X"44",X"40",X"00",X"00",X"44",X"40",X"00",X"00",X"04",X"40",X"00",X"00",X"00",X"40",
		X"00",X"00",X"04",X"40",X"00",X"00",X"44",X"40",X"00",X"04",X"44",X"40",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"04",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",
		X"00",X"44",X"40",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"4F",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"EE",X"00",X"44",X"44",X"0E",X"00",X"44",X"45",X"0E",X"00",X"44",X"55",X"00",
		X"00",X"44",X"55",X"00",X"00",X"44",X"55",X"00",X"00",X"44",X"55",X"00",X"00",X"45",X"54",X"00",
		X"00",X"55",X"40",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",
		X"00",X"66",X"60",X"00",X"00",X"66",X"66",X"00",X"00",X"F6",X"66",X"00",X"00",X"FF",X"66",X"00",
		X"00",X"FF",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"00",
		X"00",X"66",X"66",X"EE",X"00",X"66",X"66",X"0E",X"00",X"66",X"66",X"0E",X"00",X"66",X"6D",X"00",
		X"00",X"66",X"DD",X"00",X"00",X"66",X"DD",X"00",X"00",X"66",X"DD",X"00",X"00",X"6D",X"D6",X"00",
		X"00",X"DD",X"60",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CA",X"AA",X"00",X"00",X"AA",X"AA",X"00",
		X"00",X"AC",X"AA",X"00",X"00",X"CC",X"AA",X"00",X"00",X"CF",X"AA",X"00",X"00",X"CF",X"AA",X"00",
		X"00",X"CF",X"AA",X"00",X"00",X"CC",X"AA",X"00",X"00",X"AC",X"AA",X"00",X"00",X"AC",X"AA",X"00",
		X"00",X"CC",X"AA",X"00",X"00",X"CF",X"AA",X"00",X"00",X"CF",X"AA",X"00",X"00",X"CF",X"AA",X"00",
		X"00",X"CC",X"AA",X"00",X"00",X"AC",X"AA",X"00",X"00",X"AC",X"AA",X"00",X"00",X"AA",X"AA",X"00",
		X"00",X"AA",X"AA",X"00",X"00",X"CA",X"AA",X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"C6",X"66",X"00",X"00",X"66",X"66",X"00",
		X"00",X"6C",X"66",X"00",X"00",X"CC",X"66",X"00",X"00",X"CF",X"66",X"00",X"00",X"CF",X"66",X"00",
		X"00",X"CF",X"66",X"00",X"00",X"CC",X"66",X"00",X"00",X"6C",X"66",X"00",X"00",X"6C",X"66",X"00",
		X"00",X"CC",X"66",X"00",X"00",X"CF",X"66",X"00",X"00",X"CF",X"66",X"00",X"00",X"CF",X"66",X"00",
		X"00",X"CC",X"66",X"00",X"00",X"6C",X"66",X"00",X"00",X"6C",X"66",X"00",X"00",X"66",X"66",X"00",
		X"00",X"66",X"66",X"00",X"00",X"C6",X"66",X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CB",X"BB",X"00",X"00",X"BB",X"BB",X"00",
		X"00",X"BC",X"BB",X"00",X"00",X"CC",X"BB",X"00",X"00",X"CF",X"BB",X"00",X"00",X"CF",X"BB",X"00",
		X"00",X"CF",X"BB",X"00",X"00",X"CC",X"BB",X"00",X"00",X"BC",X"BB",X"00",X"00",X"BC",X"BB",X"00",
		X"00",X"CC",X"BB",X"00",X"00",X"CF",X"BB",X"00",X"00",X"CF",X"BB",X"00",X"00",X"CF",X"BB",X"00",
		X"00",X"CC",X"BB",X"00",X"00",X"BC",X"BB",X"00",X"00",X"BC",X"BB",X"00",X"00",X"BB",X"BB",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"CB",X"BB",X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",
		X"00",X"AA",X"A0",X"00",X"00",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"00",X"00",X"AF",X"AA",X"00",
		X"00",X"AF",X"AA",X"00",X"00",X"AA",X"AA",X"00",X"00",X"FA",X"AA",X"00",X"00",X"AA",X"AA",X"00",
		X"00",X"AA",X"AA",X"EE",X"00",X"AA",X"AA",X"0E",X"00",X"AA",X"A9",X"0E",X"00",X"AA",X"99",X"00",
		X"00",X"AA",X"99",X"00",X"00",X"AA",X"99",X"00",X"00",X"9A",X"99",X"00",X"00",X"A9",X"9A",X"00",
		X"00",X"99",X"A0",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"04",X"00",X"00",
		X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",
		X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"A4",X"00",X"00",X"AA",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"0A",X"00",X"00",X"00",X"F0",X"50",X"00",X"00",X"05",X"40",X"00",
		X"00",X"50",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"54",X"00",X"00",
		X"00",X"00",X"0A",X"00",X"00",X"00",X"5A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",
		X"04",X"00",X"50",X"00",X"00",X"00",X"05",X"00",X"00",X"A5",X"00",X"00",X"00",X"A5",X"00",X"00",
		X"00",X"0A",X"A0",X"40",X"00",X"0F",X"00",X"04",X"00",X"4A",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"40",X"00",X"00",X"44",X"40",X"00",X"00",X"44",X"40",X"00",X"00",X"04",X"40",
		X"00",X"00",X"44",X"40",X"00",X"00",X"44",X"40",X"00",X"00",X"44",X"40",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"04",X"00",X"00",X"44",X"04",X"00",X"00",X"44",X"04",X"00",X"00",X"44",X"04",X"00",
		X"00",X"44",X"04",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"04",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"9A",X"00",X"00",X"99",X"A9",X"00",
		X"A0",X"99",X"A9",X"90",X"AA",X"99",X"9A",X"90",X"AA",X"99",X"99",X"90",X"A6",X"99",X"99",X"90",
		X"00",X"99",X"99",X"90",X"00",X"99",X"9A",X"90",X"00",X"99",X"A9",X"90",X"00",X"99",X"A9",X"00",
		X"00",X"99",X"9A",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"04",X"00",X"00",X"44",X"04",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"04",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",
		X"00",X"A6",X"AA",X"00",X"00",X"AA",X"AA",X"00",X"00",X"AA",X"66",X"00",X"00",X"AA",X"00",X"00",
		X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"6A",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"6A",X"00",X"00",X"00",X"AA",X"60",X"00",
		X"00",X"A6",X"60",X"00",X"00",X"A6",X"A6",X"00",X"00",X"A6",X"AA",X"00",X"00",X"A6",X"AA",X"00",
		X"00",X"AA",X"6A",X"00",X"00",X"6A",X"66",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",
		X"00",X"A6",X"AA",X"00",X"00",X"AA",X"AA",X"00",X"00",X"AA",X"66",X"00",X"00",X"AA",X"00",X"00",
		X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"6A",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"6A",X"AA",X"00",
		X"00",X"AA",X"AA",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",
		X"00",X"AA",X"00",X"00",X"00",X"AA",X"AA",X"00",X"00",X"6A",X"AA",X"00",X"00",X"66",X"66",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"AA",X"AA",X"00",
		X"00",X"AA",X"AA",X"00",X"00",X"6A",X"66",X"00",X"00",X"66",X"00",X"00",X"00",X"06",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"A6",X"AA",X"00",
		X"00",X"AA",X"AA",X"00",X"00",X"AA",X"66",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",
		X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"AA",X"AA",X"00",
		X"00",X"AA",X"AA",X"00",X"00",X"6A",X"66",X"00",X"00",X"66",X"00",X"00",X"00",X"06",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"6A",X"60",X"00",X"00",X"AA",X"66",X"00",X"00",X"AA",X"A6",X"00",X"00",X"AA",X"AA",X"00",
		X"00",X"AA",X"AA",X"00",X"00",X"AA",X"6A",X"00",X"00",X"AA",X"66",X"00",X"00",X"6A",X"06",X"00",
		X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"6A",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"A6",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"6A",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",
		X"00",X"6A",X"AA",X"00",X"00",X"AA",X"AA",X"00",X"00",X"AA",X"66",X"00",X"00",X"AA",X"60",X"00",
		X"00",X"AA",X"60",X"00",X"00",X"AA",X"60",X"00",X"00",X"AA",X"60",X"00",X"00",X"6A",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"6A",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"A6",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"6A",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"A6",X"00",
		X"00",X"00",X"A6",X"00",X"00",X"66",X"A6",X"00",X"00",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"00",
		X"00",X"AA",X"A6",X"00",X"00",X"6A",X"A6",X"00",X"00",X"66",X"A6",X"00",X"00",X"06",X"A6",X"00",
		X"00",X"00",X"A6",X"00",X"00",X"00",X"A6",X"00",X"00",X"00",X"A6",X"00",X"00",X"00",X"A6",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"6A",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"A6",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"6A",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",
		X"00",X"A6",X"AA",X"00",X"00",X"AA",X"AA",X"00",X"00",X"AA",X"66",X"00",X"00",X"AA",X"00",X"00",
		X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"6A",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"6A",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"A6",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"6A",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"C5",X"55",X"00",X"00",X"55",X"55",X"00",
		X"00",X"5C",X"55",X"00",X"00",X"CC",X"55",X"00",X"00",X"CF",X"55",X"00",X"00",X"CF",X"55",X"00",
		X"00",X"CF",X"55",X"00",X"00",X"CC",X"55",X"00",X"00",X"5C",X"55",X"00",X"00",X"5C",X"55",X"00",
		X"00",X"CC",X"55",X"00",X"00",X"CF",X"55",X"00",X"00",X"CF",X"55",X"00",X"00",X"CF",X"55",X"00",
		X"00",X"CC",X"55",X"00",X"00",X"5C",X"55",X"00",X"00",X"5C",X"55",X"00",X"00",X"55",X"55",X"00",
		X"00",X"55",X"55",X"00",X"00",X"C5",X"55",X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
