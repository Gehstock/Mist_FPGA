library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity satans_hollow_bg_bits_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of satans_hollow_bg_bits_1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"AA",X"95",X"AA",X"95",X"AA",X"95",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",
		X"FF",X"AA",X"FF",X"AA",X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",X"FF",X"FA",X"FF",X"FB",
		X"6A",X"56",X"D6",X"95",X"F9",X"6A",X"FA",X"D5",X"FE",X"BE",X"FF",X"BA",X"FF",X"EA",X"FF",X"EA",
		X"BF",X"FF",X"AF",X"FF",X"AB",X"C0",X"EB",X"2A",X"E0",X"A5",X"FA",X"95",X"0A",X"55",X"A9",X"56",
		X"A9",X"55",X"59",X"54",X"68",X"00",X"68",X"00",X"A9",X"40",X"9A",X"96",X"A5",X"A5",X"AF",X"55",
		X"FE",X"AF",X"FA",X"AA",X"FA",X"FA",X"2A",X"0A",X"6A",X"55",X"59",X"55",X"59",X"A9",X"A9",X"A9",
		X"54",X"28",X"52",X"80",X"01",X"69",X"00",X"06",X"02",X"A1",X"80",X"00",X"6A",X"AA",X"55",X"55",
		X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"6A",X"50",X"6A",X"55",X"55",X"54",X"55",X"56",
		X"00",X"05",X"40",X"01",X"40",X"01",X"00",X"00",X"00",X"00",X"55",X"55",X"00",X"00",X"55",X"55",
		X"00",X"00",X"54",X"00",X"EA",X"FF",X"CA",X"00",X"28",X"A0",X"A8",X"05",X"5A",X"80",X"F5",X"55",
		X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",
		X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"AA",X"55",X"55",X"55",X"00",X"15",X"00",X"15",
		X"00",X"00",X"05",X"55",X"96",X"55",X"65",X"55",X"1A",X"AA",X"05",X"55",X"00",X"00",X"55",X"50",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"FF",X"F9",X"FC",X"06",X"00",X"01",X"00",X"00",
		X"00",X"00",X"00",X"04",X"55",X"54",X"55",X"51",X"55",X"00",X"00",X"04",X"AA",X"A8",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"54",X"00",X"50",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FC",X"00",X"01",X"00",X"55",X"00",X"55",X"01",X"55",X"05",X"55",X"15",X"55",
		X"EA",X"AA",X"FA",X"AA",X"FE",X"AA",X"FF",X"AA",X"FF",X"EA",X"FF",X"FA",X"FF",X"FA",X"FF",X"FE",
		X"FF",X"C0",X"FF",X"00",X"FC",X"00",X"F0",X"00",X"F0",X"00",X"C0",X"00",X"00",X"00",X"C0",X"00",
		X"FF",X"00",X"FF",X"F0",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FF",X"F0",
		X"FF",X"F0",X"FF",X"FC",X"FF",X"FF",X"FF",X"FC",X"FF",X"F0",X"FC",X"00",X"FF",X"00",X"F0",X"00",
		X"FF",X"C0",X"FC",X"00",X"F0",X"00",X"F0",X"00",X"C0",X"00",X"00",X"00",X"FC",X"00",X"FF",X"C0",
		X"00",X"00",X"00",X"01",X"00",X"05",X"00",X"15",X"00",X"54",X"01",X"50",X"00",X"00",X"00",X"00",
		X"15",X"55",X"55",X"55",X"00",X"55",X"C1",X"55",X"F0",X"55",X"00",X"2A",X"02",X"AA",X"00",X"00",
		X"01",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"05",X"00",X"55",X"05",X"55",
		X"15",X"6A",X"05",X"6A",X"00",X"0A",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"55",
		X"FF",X"F0",X"FF",X"00",X"FC",X"00",X"C0",X"00",X"01",X"40",X"05",X"50",X"15",X"54",X"55",X"50",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F5",X"FF",X"FC",X"FF",X"00",X"FF",X"F0",
		X"00",X"00",X"AA",X"50",X"00",X"04",X"00",X"05",X"00",X"10",X"00",X"00",X"00",X"54",X"00",X"00",
		X"55",X"00",X"54",X"00",X"50",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",
		X"55",X"00",X"AA",X"80",X"AA",X"A0",X"15",X"58",X"55",X"A8",X"55",X"2A",X"55",X"4A",X"55",X"50",
		X"00",X"28",X"00",X"80",X"2A",X"00",X"AA",X"A0",X"55",X"54",X"AA",X"A8",X"AA",X"A0",X"55",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",
		X"FF",X"C0",X"FF",X"00",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"40",X"FF",X"12",X"FF",X"06",X"FF",X"CA",X"FF",X"CA",X"FF",X"EA",X"FF",X"AA",X"FF",X"2A",
		X"FF",X"FC",X"FF",X"F0",X"FF",X"C0",X"FF",X"00",X"FF",X"01",X"FF",X"C5",X"C0",X"15",X"F0",X"55",
		X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"02",X"AA",X"0A",X"AA",X"0A",X"AA",X"2A",X"AA",
		X"00",X"2A",X"00",X"2A",X"00",X"2A",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",
		X"02",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"A2",X"AA",X"80",X"AA",X"80",X"AA",X"00",X"AA",
		X"02",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",
		X"CA",X"AA",X"CA",X"AA",X"CA",X"AA",X"CA",X"AA",X"0A",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",
		X"C2",X"A5",X"C2",X"A5",X"C2",X"A5",X"C2",X"A5",X"C2",X"A5",X"C2",X"A9",X"C2",X"A9",X"C2",X"A9",
		X"AA",X"A5",X"AA",X"A5",X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"55",X"AA",X"55",X"AA",X"95",X"AA",X"95",X"AA",X"95",X"AA",X"95",X"AA",X"A5",X"AA",X"A5",
		X"A9",X"55",X"A9",X"55",X"A9",X"55",X"A9",X"55",X"A9",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",
		X"95",X"55",X"95",X"55",X"95",X"55",X"A5",X"55",X"A5",X"55",X"A5",X"55",X"A5",X"55",X"A5",X"55",
		X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",
		X"96",X"A5",X"96",X"A5",X"96",X"A5",X"96",X"A5",X"96",X"A5",X"96",X"AA",X"96",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"A0",X"00",X"A0",X"00",X"A2",X"A8",X"A2",X"A8",X"A0",X"00",X"A0",X"00",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"A8",X"AA",X"A8",X"A0",X"00",X"A0",X"00",X"A2",X"A8",X"A2",X"A8",X"AA",X"AA",
		X"AA",X"AA",X"A0",X"28",X"A0",X"28",X"A2",X"28",X"A2",X"28",X"A2",X"00",X"A2",X"00",X"AA",X"AA",
		X"AA",X"AA",X"A0",X"00",X"A0",X"00",X"A2",X"28",X"A2",X"28",X"A2",X"28",X"A2",X"28",X"AA",X"AA",
		X"AA",X"AA",X"A0",X"00",X"A0",X"00",X"AA",X"8A",X"AA",X"8A",X"A8",X"0A",X"A8",X"0A",X"AA",X"AA",
		X"AA",X"AA",X"A2",X"00",X"A2",X"00",X"A2",X"28",X"A2",X"28",X"A2",X"28",X"A0",X"28",X"AA",X"AA",
		X"AA",X"AA",X"A2",X"80",X"A2",X"80",X"A2",X"88",X"A2",X"88",X"A0",X"00",X"A0",X"00",X"AA",X"AA",
		X"AA",X"AA",X"A0",X"00",X"A0",X"00",X"A2",X"AA",X"A2",X"AA",X"A0",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"A0",X"00",X"A0",X"00",X"A2",X"28",X"A2",X"28",X"A0",X"00",X"A0",X"00",X"AA",X"AA",
		X"AA",X"AA",X"A0",X"00",X"A0",X"00",X"A2",X"88",X"A2",X"88",X"A0",X"08",X"A0",X"08",X"AA",X"AA",
		X"5F",X"97",X"5F",X"97",X"5E",X"97",X"5E",X"A5",X"5E",X"A5",X"5E",X"A5",X"5E",X"A5",X"5E",X"A5",
		X"A9",X"7E",X"A9",X"7E",X"A9",X"7E",X"A9",X"7A",X"A9",X"7A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",
		X"97",X"FF",X"97",X"FF",X"A5",X"FF",X"A5",X"FF",X"A5",X"FF",X"A9",X"7F",X"A9",X"7F",X"A9",X"7F",
		X"A9",X"7E",X"AA",X"5E",X"AA",X"5E",X"AA",X"5E",X"AA",X"5E",X"AA",X"96",X"AA",X"9A",X"AA",X"AA",
		X"AA",X"5A",X"AA",X"5A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"A9",X"7F",X"A9",X"7F",X"A9",X"7F",X"A9",X"7F",X"A9",X"7F",X"A9",X"7F",X"A9",X"7F",X"A9",X"7F",
		X"A5",X"FF",X"A5",X"FF",X"A9",X"7F",X"A9",X"7F",X"A9",X"7F",X"AA",X"5F",X"AA",X"5F",X"AA",X"5F",
		X"AA",X"AA",X"A0",X"00",X"A0",X"00",X"A2",X"8A",X"A2",X"8A",X"A0",X"00",X"A0",X"00",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"80",X"A0",X"00",X"A0",X"88",X"A0",X"88",X"A0",X"00",X"A0",X"00",X"AA",X"AA",
		X"AA",X"AA",X"A2",X"A8",X"A2",X"A8",X"A2",X"A8",X"A2",X"A8",X"A0",X"00",X"A0",X"00",X"AA",X"AA",
		X"AA",X"AA",X"A8",X"02",X"A0",X"00",X"A0",X"A0",X"A2",X"A8",X"A0",X"00",X"A0",X"00",X"AA",X"AA",
		X"AA",X"AA",X"A2",X"A8",X"A2",X"28",X"A2",X"28",X"A2",X"28",X"A0",X"00",X"A0",X"00",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"A2",X"AA",X"A2",X"8A",X"A2",X"8A",X"A0",X"00",X"A0",X"00",X"AA",X"AA",
		X"AA",X"AA",X"A2",X"80",X"A2",X"80",X"A2",X"A8",X"A2",X"A8",X"A0",X"00",X"A0",X"00",X"AA",X"AA",
		X"AA",X"AA",X"A0",X"00",X"A0",X"00",X"AA",X"8A",X"AA",X"8A",X"A0",X"00",X"A0",X"00",X"AA",X"AA",
		X"AA",X"AA",X"A2",X"A8",X"A2",X"A8",X"A0",X"00",X"A0",X"00",X"A2",X"A8",X"A2",X"A8",X"AA",X"AA",
		X"A2",X"AA",X"A0",X"00",X"A0",X"00",X"A2",X"A8",X"A2",X"A8",X"AA",X"80",X"AA",X"80",X"AA",X"AA",
		X"AA",X"AA",X"A2",X"A8",X"A2",X"A0",X"A0",X"82",X"A8",X"0A",X"A0",X"00",X"A0",X"00",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"A0",X"AA",X"A0",X"AA",X"A8",X"AA",X"A8",X"A0",X"00",X"A0",X"00",X"AA",X"AA",
		X"AA",X"AA",X"A0",X"00",X"A2",X"AA",X"A0",X"00",X"A2",X"AA",X"A0",X"00",X"A0",X"00",X"AA",X"AA",
		X"AA",X"AA",X"A0",X"00",X"A0",X"00",X"AA",X"02",X"A8",X"2A",X"A0",X"00",X"A0",X"00",X"AA",X"AA",
		X"AA",X"AA",X"A0",X"00",X"A0",X"00",X"A2",X"A8",X"A2",X"A8",X"A0",X"00",X"A0",X"00",X"AA",X"AA",
		X"AA",X"AA",X"A0",X"0A",X"A0",X"0A",X"A2",X"8A",X"A2",X"8A",X"A0",X"00",X"A0",X"00",X"AA",X"AA",
		X"AA",X"AA",X"A0",X"00",X"A0",X"00",X"A2",X"A0",X"A2",X"A8",X"A0",X"00",X"A0",X"00",X"AA",X"AA",
		X"AA",X"AA",X"A0",X"20",X"A0",X"00",X"A2",X"0A",X"A2",X"2A",X"A0",X"00",X"A0",X"00",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"A2",X"00",X"A2",X"00",X"A2",X"28",X"A2",X"28",X"A0",X"28",X"AA",X"AA",
		X"AA",X"AA",X"A0",X"AA",X"A2",X"A8",X"A0",X"00",X"A0",X"00",X"A2",X"A8",X"A0",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"A0",X"00",X"A0",X"00",X"AA",X"A8",X"AA",X"A8",X"A0",X"00",X"A0",X"00",X"AA",X"AA",
		X"AA",X"AA",X"A2",X"AA",X"A0",X"0A",X"AA",X"80",X"A0",X"00",X"A0",X"0A",X"A2",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"A0",X"00",X"AA",X"A8",X"A0",X"00",X"AA",X"A8",X"A0",X"00",X"A0",X"00",X"AA",X"AA",
		X"AA",X"AA",X"A2",X"A8",X"A0",X"80",X"AA",X"0A",X"A0",X"2A",X"A0",X"8A",X"A2",X"A0",X"AA",X"AA",
		X"AA",X"AA",X"A2",X"AA",X"A0",X"AA",X"AA",X"00",X"A8",X"00",X"A0",X"2A",X"A2",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"A2",X"A8",X"A0",X"A8",X"A0",X"28",X"A2",X"08",X"A2",X"80",X"A2",X"A0",X"AA",X"AA",
		X"AA",X"A5",X"AA",X"A5",X"AA",X"A5",X"AA",X"A5",X"AA",X"A5",X"AA",X"A5",X"AA",X"A5",X"AA",X"A5",
		X"AA",X"AA",X"AA",X"AA",X"FE",X"AA",X"FE",X"AA",X"FE",X"AA",X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",
		X"7F",X"FA",X"7F",X"FA",X"7F",X"FA",X"7F",X"FA",X"7F",X"FE",X"7F",X"FE",X"7F",X"FE",X"7F",X"FE",
		X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"FE",X"AA",X"FE",X"AA",
		X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",
		X"FF",X"EF",X"FF",X"EF",X"FF",X"EF",X"FF",X"EF",X"FF",X"EB",X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",
		X"C1",X"55",X"01",X"55",X"02",X"55",X"02",X"55",X"0A",X"95",X"0A",X"95",X"0A",X"95",X"0A",X"A5",
		X"CA",X"A5",X"CA",X"A5",X"CA",X"A5",X"CA",X"A5",X"C2",X"95",X"C2",X"95",X"C2",X"95",X"C2",X"55",
		X"EA",X"AA",X"EA",X"AA",X"EA",X"A9",X"EA",X"A9",X"CA",X"A5",X"CA",X"A5",X"CA",X"A5",X"CA",X"A5",
		X"FF",X"EA",X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",X"FF",X"FE",
		X"55",X"55",X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",
		X"A5",X"55",X"A5",X"55",X"A5",X"55",X"A5",X"55",X"A5",X"55",X"95",X"55",X"95",X"55",X"95",X"55",
		X"A5",X"55",X"A5",X"55",X"A5",X"55",X"A5",X"55",X"A5",X"55",X"A5",X"55",X"A5",X"55",X"A5",X"55",
		X"A9",X"55",X"A9",X"55",X"A9",X"55",X"A9",X"55",X"A9",X"55",X"A9",X"55",X"A9",X"55",X"A9",X"55",
		X"AA",X"A5",X"AA",X"A5",X"AA",X"A5",X"AA",X"95",X"AA",X"95",X"AA",X"95",X"AA",X"95",X"AA",X"95",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"FF",X"FD",X"FF",X"FD",X"FF",X"D5",X"FF",X"D5",
		X"FF",X"FF",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"D5",X"FF",X"55",X"FF",X"55",X"FD",X"55",
		X"BF",X"FA",X"AF",X"EA",X"AB",X"AB",X"EA",X"AB",X"EA",X"AB",X"EA",X"AF",X"FA",X"AF",X"FA",X"BF",
		X"F7",X"77",X"5D",X"DD",X"57",X"77",X"55",X"DD",X"55",X"77",X"55",X"DD",X"55",X"77",X"55",X"55",
		X"55",X"00",X"55",X"00",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"54",X"55",X"55",
		X"50",X"00",X"50",X"01",X"40",X"05",X"50",X"0A",X"54",X"00",X"54",X"00",X"54",X"00",X"54",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"55",X"40",X"55",X"50",X"55",X"54",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"CF",X"69",X"F3",X"AB",X"F3",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"A5",X"55",X"A5",X"55",X"AA",X"55",X"AA",X"55",
		X"E5",X"FF",X"D7",X"FF",X"D5",X"7F",X"F5",X"7F",X"FD",X"BF",X"FF",X"AF",X"FF",X"5F",X"FD",X"6F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F5",X"FF",X"57",X"FF",X"5F",X"FF",X"5F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"D5",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"AA",X"55",X"AA",X"A9",X"AA",X"A9",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"7F",X"55",X"7F",X"55",X"7F",X"55",X"7F",X"55",X"7F",X"55",X"7F",X"55",X"5F",X"55",X"5F",
		X"66",X"BE",X"55",X"7E",X"EA",X"67",X"7E",X"A5",X"57",X"57",X"F7",X"F7",X"DD",X"AB",X"D5",X"FB",
		X"FF",X"FD",X"BF",X"FF",X"AF",X"FF",X"AB",X"FF",X"AA",X"C0",X"AA",X"8D",X"AA",X"87",X"AA",X"8D",
		X"7F",X"FF",X"5F",X"FF",X"D7",X"FF",X"D5",X"FF",X"F5",X"7F",X"FD",X"5F",X"FF",X"5F",X"FF",X"DF",
		X"C1",X"56",X"F0",X"5A",X"7C",X"6A",X"5C",X"6A",X"5C",X"2A",X"5F",X"0A",X"DF",X"CA",X"F7",X"CA",
		X"FF",X"06",X"F7",X"CA",X"F7",X"CA",X"D7",X"C2",X"D7",X"C2",X"F7",X"F2",X"F5",X"F2",X"FD",X"F2",
		X"FF",X"FF",X"FF",X"DF",X"FF",X"DF",X"FF",X"DF",X"FF",X"5F",X"FF",X"57",X"FD",X"57",X"55",X"55",
		X"2F",X"15",X"2F",X"15",X"2F",X"15",X"2F",X"15",X"2F",X"15",X"2F",X"15",X"3C",X"15",X"F0",X"55",
		X"AB",X"C5",X"AB",X"C5",X"AB",X"C5",X"AB",X"C5",X"AB",X"C5",X"AB",X"C5",X"AB",X"C5",X"AF",X"15",
		X"AB",X"30",X"AB",X"0C",X"AB",X"0F",X"AB",X"CF",X"AB",X"C3",X"AB",X"C7",X"AB",X"C7",X"AB",X"C7",
		X"FC",X"FF",X"5F",X"0F",X"5F",X"CF",X"5F",X"CF",X"5F",X"CF",X"9F",X"C3",X"97",X"F0",X"97",X"FC",
		X"55",X"7C",X"55",X"7F",X"AA",X"AF",X"AA",X"AF",X"AA",X"AF",X"A5",X"57",X"AA",X"AB",X"AA",X"AB",
		X"7C",X"FC",X"7C",X"FC",X"7C",X"FC",X"0F",X"3C",X"57",X"F1",X"57",X"F1",X"57",X"F1",X"57",X"05",
		X"CF",X"FF",X"CF",X"FF",X"F3",X"FF",X"F3",X"FF",X"F3",X"FF",X"F3",X"FC",X"F3",X"F1",X"F3",X"F1",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"1A",X"FF",X"16",X"FF",X"15",X"FC",X"15",X"F0",X"55",X"F1",X"55",X"F1",X"55",X"F1",X"55",
		X"FF",X"F1",X"FF",X"C1",X"FF",X"C5",X"FF",X"C5",X"FF",X"05",X"FF",X"15",X"FF",X"15",X"FF",X"16",
		X"D5",X"F3",X"F5",X"F3",X"FF",X"F0",X"FF",X"CC",X"FF",X"CC",X"FF",X"CF",X"FF",X"CF",X"FF",X"C3",
		X"F3",X"FF",X"FC",X"FF",X"FC",X"3F",X"BF",X"3F",X"AF",X"0F",X"AF",X"CF",X"AF",X"C3",X"AB",X"F3",
		X"AB",X"F3",X"AA",X"FC",X"6A",X"FC",X"6A",X"BF",X"6A",X"BF",X"6A",X"BF",X"5A",X"AF",X"5A",X"AF",
		X"F3",X"FE",X"F3",X"FB",X"F3",X"FB",X"F3",X"EE",X"F0",X"FB",X"FC",X"EE",X"FC",X"BB",X"FC",X"EE",
		X"FC",X"FB",X"FC",X"3E",X"FF",X"3B",X"FF",X"0E",X"FF",X"CF",X"FF",X"CE",X"FF",X"C1",X"7F",X"F1",
		X"7F",X"0D",X"5F",X"CD",X"5F",X"CF",X"5F",X"CF",X"5F",X"C3",X"57",X"F3",X"57",X"F3",X"57",X"F3",
		X"53",X"F3",X"43",X"F3",X"43",X"F3",X"03",X"FC",X"03",X"FC",X"43",X"F0",X"50",X"F2",X"54",X"CA",
		X"57",X"FC",X"5F",X"FC",X"5F",X"F0",X"5F",X"F1",X"5F",X"C1",X"5F",X"C6",X"7F",X"0A",X"FF",X"15",
		X"99",X"99",X"66",X"66",X"99",X"99",X"66",X"66",X"99",X"99",X"66",X"66",X"99",X"99",X"66",X"66",
		X"91",X"FC",X"64",X"FC",X"91",X"FC",X"67",X"FC",X"13",X"FC",X"47",X"FC",X"53",X"FC",X"57",X"FC",
		X"FF",X"15",X"FF",X"15",X"FF",X"15",X"FF",X"15",X"FF",X"15",X"FF",X"15",X"FF",X"15",X"FF",X"15",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"F0",X"FF",X"F1",
		X"3F",X"FF",X"1F",X"FF",X"17",X"FF",X"15",X"FF",X"15",X"7F",X"15",X"5F",X"15",X"57",X"15",X"57",
		X"BF",X"FF",X"B7",X"FF",X"FE",X"FF",X"5E",X"FF",X"E9",X"BF",X"E9",X"BF",X"76",X"BF",X"EA",X"DF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"D5",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"D7",
		X"55",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"F5",X"FF",X"F5",X"FF",X"D5",X"FF",X"D5",X"F5",X"55",X"F5",X"55",X"F5",X"55",X"FF",X"55",
		X"FF",X"FF",X"7F",X"FF",X"7F",X"FF",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"55",X"7F",X"55",X"55",
		X"55",X"5F",X"55",X"5F",X"55",X"FF",X"55",X"FF",X"5F",X"FF",X"5F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"6A",X"5A",X"AA",X"5A",X"AA",X"6A",X"AA",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"55",X"6F",X"56",X"AF",X"57",X"FF",X"5B",X"FF",X"5B",X"FF",X"AF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"59",X"55",X"59",X"55",X"65",X"55",X"65",X"55",X"95",X"6A",X"55",X"95",X"55",X"55",X"55",
		X"56",X"A5",X"55",X"A9",X"55",X"6A",X"55",X"5A",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"D5",X"55",X"F5",X"55",X"FD",X"55",X"FF",X"55",X"FF",X"D5",X"FF",X"F5",X"FF",X"FD",
		X"AA",X"AB",X"AA",X"AF",X"AA",X"BF",X"AA",X"FF",X"AB",X"FF",X"AF",X"FF",X"BF",X"FF",X"FF",X"FF",
		X"55",X"57",X"55",X"5F",X"55",X"7F",X"55",X"FF",X"57",X"FF",X"5F",X"FF",X"7F",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"77",X"77",X"DD",X"DD",X"77",X"77",X"DD",X"DD",X"77",X"77",X"DD",X"DD",X"77",X"77",X"DD",X"DD",
		X"FF",X"FC",X"FF",X"F1",X"FF",X"C7",X"FF",X"0D",X"FC",X"37",X"FC",X"DD",X"F3",X"77",X"C1",X"DD",
		X"AB",X"FF",X"AB",X"FF",X"AB",X"FF",X"AB",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"BF",X"AA",X"BF",
		X"FF",X"C0",X"FC",X"00",X"C0",X"00",X"28",X"00",X"80",X"00",X"C0",X"80",X"FE",X"00",X"FF",X"00",
		X"FF",X"C4",X"03",X"C0",X"13",X"C0",X"13",X"C0",X"10",X"01",X"15",X"55",X"15",X"55",X"15",X"55",
		X"FF",X"FD",X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"5F",X"FF",X"5F",X"7F",X"FF",
		X"FF",X"37",X"FC",X"1D",X"FC",X"77",X"FC",X"DD",X"FC",X"77",X"FC",X"DD",X"FC",X"77",X"FC",X"DD",
		X"FF",X"C7",X"FF",X"CD",X"FF",X"07",X"FF",X"1D",X"FF",X"37",X"FF",X"1D",X"FF",X"37",X"FF",X"1D",
		X"70",X"00",X"00",X"01",X"00",X"07",X"00",X"DD",X"07",X"74",X"DD",X"D1",X"77",X"07",X"DC",X"DD",
		X"77",X"00",X"00",X"01",X"00",X"55",X"05",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"55",X"40",
		X"FC",X"00",X"3C",X"1D",X"30",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"C1",X"DD",
		X"FF",X"C7",X"FF",X"CD",X"FF",X"C7",X"FF",X"CD",X"FF",X"C7",X"FF",X"CD",X"FF",X"C7",X"FF",X"0D",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"C0",X"FF",X"CD",X"FF",X"C7",X"FF",X"CD",X"FF",X"C7",X"FF",X"CD",
		X"00",X"00",X"00",X"0D",X"03",X"77",X"01",X"DD",X"77",X"77",X"DD",X"DD",X"77",X"77",X"DD",X"DD",
		X"00",X"00",X"00",X"00",X"00",X"37",X"0D",X"DD",X"77",X"77",X"DD",X"DD",X"77",X"77",X"DD",X"DD",
		X"F3",X"77",X"F1",X"DD",X"C7",X"77",X"CD",X"DD",X"C7",X"77",X"CD",X"DD",X"C7",X"77",X"DD",X"DD",
		X"FF",X"C0",X"FF",X"C1",X"FF",X"37",X"FF",X"1D",X"FC",X"77",X"FC",X"DD",X"FC",X"77",X"FC",X"00",
		X"00",X"00",X"DD",X"DD",X"77",X"77",X"DD",X"DD",X"77",X"77",X"DD",X"DD",X"77",X"77",X"DD",X"DD",
		X"00",X"77",X"1D",X"DD",X"77",X"77",X"DD",X"DD",X"77",X"77",X"DD",X"C0",X"00",X"37",X"DD",X"DD",
		X"37",X"70",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"1D",
		X"FC",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"1D",X"FC",X"37",X"FC",X"1D",X"FC",X"37",X"F0",X"DD",
		X"FF",X"F3",X"FF",X"F1",X"FF",X"C7",X"FF",X"CD",X"FF",X"37",X"FF",X"1D",X"FF",X"37",X"FF",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"FE",X"BF",X"FA",X"BF",X"EA",X"BF",X"AA",X"BF",X"AA",X"AA",
		X"FF",X"F3",X"FF",X"C3",X"FF",X"03",X"FC",X"03",X"F0",X"0F",X"C0",X"0F",X"00",X"3F",X"AA",X"AA",
		X"AA",X"AA",X"FA",X"AA",X"FA",X"AA",X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",X"FF",X"FA",X"FF",X"FE",
		X"55",X"56",X"55",X"5A",X"55",X"5A",X"55",X"6A",X"55",X"AA",X"56",X"AA",X"5A",X"AA",X"6A",X"AA",
		X"AB",X"FF",X"AB",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"BF",
		X"DD",X"DD",X"77",X"77",X"5D",X"DD",X"57",X"77",X"55",X"DD",X"55",X"77",X"55",X"5D",X"55",X"57",
		X"FF",X"FF",X"FF",X"FF",X"F3",X"00",X"F3",X"00",X"F3",X"3C",X"F3",X"3C",X"F0",X"3C",X"FF",X"FF",
		X"FF",X"FF",X"F0",X"00",X"F0",X"00",X"FF",X"CF",X"FF",X"CF",X"F0",X"00",X"F0",X"00",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"F0",X"FF",X"F0",X"FF",X"FC",X"FF",X"FC",X"F0",X"00",X"F0",X"00",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"DD",X"DF",X"77",X"7F",X"DD",X"FF",X"77",X"FF",X"DF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"77",X"7F",X"DD",X"DF",X"77",X"FF",X"DD",X"FF",X"7F",X"FF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"82",X"C0",X"00",X"C0",X"00",X"F0",X"28",X"C2",X"80",X"CA",X"00",X"20",X"00",X"00",X"08",
		X"AB",X"FF",X"AB",X"FF",X"AB",X"FF",X"AB",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"BF",X"AA",X"BF",
		X"55",X"5A",X"55",X"AA",X"56",X"AA",X"5A",X"AA",X"56",X"AA",X"55",X"AA",X"55",X"6A",X"55",X"5A",
		X"57",X"FF",X"57",X"FF",X"57",X"FF",X"55",X"FF",X"55",X"5F",X"55",X"5F",X"55",X"5F",X"55",X"5F",
		X"57",X"75",X"DF",X"FD",X"75",X"57",X"FD",X"DD",X"5D",X"FF",X"DF",X"D5",X"FD",X"5D",X"DD",X"7F",
		X"FF",X"FF",X"FF",X"FC",X"3F",X"F0",X"FF",X"02",X"C0",X"00",X"20",X"00",X"80",X"A8",X"02",X"00",
		X"14",X"51",X"14",X"51",X"14",X"54",X"15",X"14",X"45",X"44",X"51",X"44",X"51",X"45",X"11",X"45",
		X"FF",X"FF",X"FE",X"FF",X"FE",X"FF",X"FF",X"BF",X"FF",X"EF",X"FF",X"EF",X"FF",X"FB",X"FF",X"FE",
		X"55",X"51",X"15",X"51",X"15",X"51",X"15",X"11",X"15",X"11",X"15",X"15",X"55",X"15",X"55",X"15",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",X"DD",X"FF",X"F7",X"DF",X"FF",X"77",X"FF",X"DF",X"FF",
		X"FF",X"5F",X"FD",X"DF",X"FD",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"D7",X"5F",X"DD",X"DF",X"F5",
		X"FF",X"FF",X"FD",X"FF",X"DD",X"DF",X"F7",X"7F",X"5D",X"D7",X"F7",X"7F",X"DD",X"DF",X"FD",X"FF",
		X"FF",X"0A",X"FF",X"A0",X"F0",X"00",X"CA",X"00",X"20",X"02",X"80",X"0A",X"00",X"28",X"00",X"0A",
		X"15",X"5A",X"15",X"AA",X"16",X"AA",X"5A",X"AA",X"56",X"AA",X"55",X"AA",X"45",X"6A",X"45",X"5A",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EA",X"FA",X"BF",X"AB",X"FF",X"FF",X"FF",
		X"A8",X"2A",X"A8",X"A2",X"A2",X"82",X"A2",X"02",X"A2",X"82",X"A0",X"A2",X"A0",X"2A",X"A0",X"0A",
		X"77",X"7F",X"DD",X"DF",X"77",X"FF",X"DD",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"A0",X"0A",X"A0",X"2A",X"A0",X"A2",X"A0",X"82",X"A2",X"02",X"A2",X"82",X"A8",X"22",X"A8",X"2A",
		X"55",X"51",X"51",X"51",X"51",X"51",X"51",X"55",X"51",X"55",X"51",X"55",X"51",X"55",X"55",X"55",
		X"FF",X"FF",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"FF",X"FF",
		X"FF",X"FF",X"F0",X"00",X"F0",X"00",X"F3",X"FC",X"F3",X"FC",X"F0",X"00",X"F0",X"00",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FC",X"F0",X"00",X"F0",X"00",X"F3",X"FC",X"F3",X"FC",X"FF",X"FF",
		X"FF",X"FF",X"F0",X"3C",X"F0",X"3C",X"F3",X"3C",X"F3",X"3C",X"F3",X"00",X"F3",X"00",X"FF",X"FF",
		X"FF",X"FF",X"F0",X"00",X"F0",X"00",X"F3",X"3C",X"F3",X"3C",X"F3",X"3C",X"F3",X"3C",X"FF",X"FF",
		X"FF",X"FF",X"F0",X"00",X"F0",X"00",X"FF",X"CF",X"FF",X"CF",X"FC",X"0F",X"FC",X"0F",X"FF",X"FF",
		X"FF",X"FF",X"F3",X"00",X"F3",X"00",X"F3",X"3C",X"F3",X"3C",X"F3",X"3C",X"F0",X"3C",X"FF",X"FF",
		X"FF",X"FF",X"F3",X"C0",X"F3",X"C0",X"F3",X"CC",X"F3",X"CC",X"F0",X"00",X"F0",X"00",X"FF",X"FF",
		X"FF",X"FF",X"F0",X"00",X"F0",X"00",X"F3",X"FF",X"F3",X"FF",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"F0",X"00",X"F0",X"00",X"F3",X"3C",X"F3",X"3C",X"F0",X"00",X"F0",X"00",X"FF",X"FF",
		X"FF",X"FF",X"F0",X"00",X"F0",X"00",X"F3",X"CC",X"F3",X"CC",X"F0",X"0C",X"F0",X"0C",X"FF",X"FF",
		X"FF",X"0F",X"FC",X"0F",X"F0",X"8F",X"C2",X"8F",X"0A",X"8F",X"2A",X"8F",X"AA",X"80",X"AA",X"AA",
		X"FF",X"FF",X"F3",X"FC",X"F3",X"3C",X"F3",X"3C",X"F3",X"3C",X"F0",X"00",X"F0",X"00",X"FF",X"FF",
		X"80",X"02",X"2A",X"A8",X"22",X"88",X"22",X"88",X"22",X"88",X"28",X"28",X"2A",X"A8",X"80",X"02",
		X"FF",X"FF",X"FF",X"FC",X"F3",X"FC",X"F3",X"FC",X"F3",X"FC",X"F0",X"00",X"F0",X"00",X"FF",X"FF",
		X"FF",X"FF",X"F0",X"30",X"F0",X"00",X"F3",X"0F",X"F3",X"3F",X"F0",X"00",X"F0",X"00",X"FF",X"FF",
		X"FF",X"FF",X"FC",X"03",X"F0",X"00",X"F0",X"F0",X"F3",X"FC",X"F0",X"00",X"F0",X"00",X"FF",X"FF",
		X"FF",X"FF",X"F3",X"FC",X"F3",X"FC",X"F0",X"00",X"F0",X"00",X"F3",X"FC",X"F3",X"FC",X"FF",X"FF",
		X"FF",X"FF",X"F0",X"FF",X"F3",X"FC",X"F0",X"00",X"F0",X"00",X"F3",X"FC",X"F0",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
