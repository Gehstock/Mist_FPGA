library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ps02 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ps02 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"08",X"FE",X"03",X"CA",X"45",X"08",X"FE",X"02",X"CA",X"39",X"08",X"CD",X"42",X"0B",X"23",X"70",
		X"2E",X"04",X"70",X"2E",X"07",X"70",X"2E",X"14",X"70",X"2E",X"17",X"70",X"2E",X"1A",X"70",X"2E",
		X"3A",X"70",X"21",X"BE",X"20",X"70",X"CD",X"ED",X"0E",X"FE",X"03",X"D0",X"FE",X"02",X"2E",X"4D",
		X"CA",X"36",X"08",X"36",X"04",X"C9",X"36",X"02",X"C9",X"CD",X"42",X"0B",X"2E",X"0A",X"70",X"2E",
		X"1D",X"70",X"C3",X"0B",X"08",X"CD",X"42",X"0B",X"2E",X"0D",X"70",X"2E",X"20",X"70",X"2E",X"3D",
		X"70",X"21",X"C5",X"20",X"70",X"C3",X"39",X"08",X"CD",X"42",X"0B",X"2E",X"40",X"70",X"21",X"CC",
		X"20",X"70",X"C3",X"45",X"08",X"FE",X"18",X"D4",X"7F",X"08",X"CD",X"42",X"0B",X"2E",X"43",X"70",
		X"C3",X"58",X"08",X"CD",X"ED",X"0E",X"FE",X"12",X"D8",X"21",X"FA",X"20",X"36",X"01",X"C9",X"CD",
		X"42",X"0B",X"2E",X"46",X"70",X"C9",X"06",X"0A",X"C5",X"E7",X"0F",X"21",X"02",X"25",X"DA",X"93",
		X"08",X"2E",X"01",X"06",X"40",X"CD",X"CB",X"03",X"CD",X"8A",X"03",X"E7",X"0F",X"11",X"2F",X"05",
		X"21",X"02",X"25",X"DA",X"AB",X"08",X"11",X"37",X"05",X"2E",X"01",X"0E",X"08",X"CD",X"E6",X"02",
		X"CD",X"8A",X"03",X"C1",X"05",X"C2",X"88",X"08",X"E7",X"0F",X"21",X"02",X"CE",X"DA",X"C2",X"08",
		X"2E",X"01",X"11",X"01",X"0A",X"3E",X"06",X"C3",X"6E",X"0A",X"21",X"D3",X"20",X"AF",X"BE",X"C8",
		X"35",X"C9",X"21",X"D3",X"20",X"AF",X"BE",X"C9",X"E7",X"2E",X"39",X"C9",X"CD",X"09",X"0B",X"01",
		X"04",X"04",X"09",X"C9",X"E7",X"2E",X"4F",X"7E",X"C9",X"E1",X"11",X"10",X"43",X"06",X"03",X"F7",
		X"C5",X"E5",X"1A",X"D3",X"03",X"DB",X"03",X"2F",X"A6",X"77",X"23",X"13",X"AF",X"D3",X"03",X"DB",
		X"03",X"2F",X"A6",X"77",X"E1",X"01",X"20",X"00",X"09",X"C1",X"05",X"C2",X"F0",X"08",X"C9",X"F7",
		X"C5",X"E5",X"AF",X"D3",X"03",X"DB",X"03",X"77",X"23",X"0D",X"C2",X"12",X"09",X"AF",X"D3",X"03",
		X"DB",X"03",X"77",X"E1",X"01",X"20",X"00",X"09",X"C1",X"05",X"C2",X"10",X"09",X"C9",X"3A",X"0D",
		X"23",X"A7",X"C8",X"3A",X"06",X"23",X"B0",X"32",X"06",X"23",X"D3",X"04",X"C9",X"3A",X"06",X"23",
		X"A0",X"32",X"06",X"23",X"D3",X"04",X"C9",X"3A",X"07",X"23",X"A0",X"32",X"07",X"23",X"D3",X"06",
		X"C9",X"3A",X"0D",X"23",X"A7",X"C8",X"3A",X"07",X"23",X"B0",X"32",X"07",X"23",X"D3",X"06",X"C9",
		X"35",X"C3",X"87",X"00",X"21",X"F0",X"20",X"AF",X"BE",X"C2",X"60",X"09",X"21",X"4D",X"20",X"34",
		X"7E",X"E6",X"03",X"77",X"23",X"34",X"7E",X"E6",X"07",X"77",X"CD",X"FF",X"18",X"CD",X"F2",X"0E",
		X"CD",X"2C",X"0F",X"CD",X"B7",X"09",X"CD",X"04",X"0A",X"CD",X"04",X"13",X"CD",X"BD",X"05",X"CD",
		X"6B",X"16",X"2A",X"3C",X"20",X"23",X"22",X"3C",X"20",X"CD",X"F3",X"16",X"CD",X"D7",X"16",X"CD",
		X"7A",X"16",X"00",X"00",X"00",X"CD",X"38",X"16",X"CD",X"C9",X"16",X"CD",X"5B",X"16",X"00",X"00",
		X"00",X"CD",X"45",X"0A",X"C3",X"87",X"00",X"3A",X"4D",X"20",X"A7",X"CA",X"CE",X"09",X"FE",X"01",
		X"CA",X"DA",X"09",X"FE",X"02",X"CA",X"E9",X"09",X"FE",X"03",X"CA",X"F5",X"09",X"C9",X"CD",X"AD",
		X"0B",X"CD",X"CA",X"08",X"CD",X"DE",X"4A",X"C3",X"46",X"11",X"CD",X"F5",X"0C",X"CD",X"E4",X"0F",
		X"CD",X"84",X"49",X"CD",X"A9",X"17",X"C3",X"73",X"1C",X"CD",X"69",X"0D",X"CD",X"78",X"10",X"CD",
		X"FB",X"1D",X"C3",X"8E",X"18",X"CD",X"C2",X"0D",X"CD",X"DF",X"10",X"CD",X"60",X"4A",X"CD",X"39",
		X"18",X"C3",X"D5",X"18",X"3A",X"4E",X"20",X"A7",X"CA",X"1B",X"0A",X"FE",X"01",X"CA",X"27",X"0A",
		X"FE",X"02",X"CA",X"2D",X"0A",X"FE",X"03",X"CA",X"39",X"0A",X"C9",X"CD",X"AD",X"11",X"CD",X"EB",
		X"17",X"CD",X"69",X"17",X"C3",X"82",X"1D",X"CD",X"86",X"0E",X"C3",X"DA",X"13",X"CD",X"24",X"12",
		X"CD",X"2B",X"13",X"CD",X"5C",X"4B",X"C3",X"C7",X"1C",X"CD",X"94",X"12",X"CD",X"99",X"13",X"CD",
		X"27",X"1D",X"C3",X"04",X"1F",X"21",X"E5",X"20",X"AF",X"BE",X"C8",X"CD",X"ED",X"0E",X"FE",X"04",
		X"21",X"94",X"20",X"06",X"01",X"70",X"D8",X"FE",X"07",X"2E",X"9F",X"70",X"D8",X"2E",X"D4",X"70",
		X"C9",X"01",X"EB",X"43",X"0A",X"FE",X"FF",X"C8",X"CD",X"81",X"0A",X"C3",X"64",X"0A",X"D5",X"E5",
		X"77",X"23",X"1D",X"C2",X"70",X"0A",X"E1",X"01",X"80",X"00",X"09",X"D1",X"15",X"C2",X"6E",X"0A",
		X"C9",X"6F",X"03",X"0A",X"67",X"03",X"0A",X"5F",X"03",X"0A",X"57",X"03",X"0A",X"03",X"C5",X"DF",
		X"C1",X"C9",X"21",X"04",X"24",X"01",X"03",X"10",X"11",X"33",X"43",X"CD",X"A8",X"05",X"D5",X"21",
		X"04",X"26",X"CD",X"DD",X"0A",X"21",X"04",X"29",X"CD",X"E3",X"0A",X"D1",X"D5",X"21",X"04",X"2C",
		X"CD",X"DD",X"0A",X"21",X"04",X"2F",X"CD",X"E3",X"0A",X"D1",X"D5",X"21",X"04",X"32",X"CD",X"DD",
		X"0A",X"21",X"04",X"35",X"CD",X"E3",X"0A",X"D1",X"21",X"04",X"38",X"CD",X"DD",X"0A",X"21",X"04",
		X"3B",X"CD",X"E3",X"0A",X"21",X"04",X"3E",X"01",X"04",X"10",X"C3",X"A8",X"05",X"01",X"01",X"18",
		X"C3",X"A8",X"05",X"01",X"02",X"18",X"C3",X"A8",X"05",X"21",X"02",X"35",X"11",X"32",X"44",X"0E",
		X"05",X"CD",X"E6",X"02",X"CD",X"ED",X"0E",X"FE",X"0A",X"21",X"02",X"3B",X"D2",X"05",X"0B",X"24",
		X"C6",X"1C",X"C3",X"F2",X"02",X"27",X"C3",X"30",X"03",X"23",X"5E",X"23",X"56",X"EB",X"C9",X"CD",
		X"C4",X"04",X"C3",X"DA",X"03",X"73",X"23",X"72",X"23",X"C9",X"06",X"18",X"C3",X"CA",X"03",X"79",
		X"A7",X"CA",X"2C",X"0B",X"11",X"03",X"00",X"19",X"0D",X"C2",X"27",X"0B",X"7E",X"A7",X"C9",X"7D",
		X"E6",X"07",X"CD",X"DB",X"04",X"01",X"00",X"A0",X"09",X"C9",X"CD",X"09",X"0B",X"01",X"F8",X"0A",
		X"09",X"C9",X"E7",X"2E",X"00",X"C9",X"E7",X"2E",X"13",X"C9",X"F5",X"CD",X"ED",X"0E",X"FE",X"23",
		X"D2",X"94",X"0B",X"FE",X"18",X"D2",X"99",X"0B",X"FE",X"14",X"D2",X"A3",X"0B",X"FE",X"10",X"D2",
		X"76",X"0B",X"FE",X"06",X"D2",X"80",X"0B",X"FE",X"03",X"D2",X"8A",X"0B",X"F1",X"FE",X"88",X"21",
		X"FC",X"00",X"D0",X"2E",X"FE",X"C9",X"F1",X"21",X"FA",X"00",X"FE",X"88",X"D0",X"2E",X"FB",X"C9",
		X"F1",X"21",X"FB",X"00",X"FE",X"88",X"D0",X"2E",X"FC",X"C9",X"F1",X"21",X"FC",X"00",X"FE",X"88",
		X"D0",X"2E",X"FD",X"C9",X"F1",X"21",X"F8",X"00",X"C9",X"F1",X"21",X"F8",X"00",X"FE",X"88",X"D0",
		X"2E",X"F9",X"C9",X"F1",X"21",X"F9",X"00",X"FE",X"88",X"D0",X"2E",X"F8",X"C9",X"21",X"00",X"20",
		X"AF",X"BE",X"C8",X"23",X"BE",X"C2",X"BC",X"0B",X"34",X"CD",X"80",X"05",X"3A",X"0D",X"23",X"A7",
		X"C2",X"E4",X"0B",X"3A",X"20",X"23",X"3C",X"32",X"20",X"23",X"E6",X"07",X"2A",X"21",X"23",X"C2",
		X"D9",X"0B",X"7D",X"FE",X"AD",X"CC",X"E0",X"0B",X"23",X"22",X"21",X"23",X"7E",X"C3",X"E7",X"0B",
		X"21",X"91",X"44",X"C9",X"C3",X"00",X"4F",X"07",X"DA",X"52",X"0C",X"07",X"DA",X"78",X"0C",X"07",
		X"DA",X"9C",X"0C",X"07",X"DA",X"B6",X"0C",X"21",X"00",X"00",X"22",X"02",X"20",X"CD",X"80",X"05",
		X"21",X"02",X"20",X"EF",X"2A",X"04",X"20",X"7D",X"FE",X"74",X"D2",X"14",X"0C",X"FF",X"3E",X"07",
		X"11",X"02",X"07",X"DF",X"21",X"04",X"20",X"CD",X"C4",X"04",X"F7",X"C5",X"E5",X"1A",X"D3",X"03",
		X"DB",X"03",X"A6",X"CA",X"2B",X"0C",X"3E",X"01",X"32",X"37",X"20",X"DB",X"03",X"AE",X"77",X"23",
		X"13",X"0D",X"C2",X"1D",X"0C",X"AF",X"D3",X"03",X"DB",X"03",X"A6",X"CA",X"43",X"0C",X"3E",X"01",
		X"32",X"37",X"20",X"DB",X"03",X"AE",X"77",X"E1",X"01",X"20",X"00",X"09",X"C1",X"05",X"C2",X"1B",
		X"0C",X"C9",X"21",X"3E",X"20",X"3A",X"04",X"20",X"BE",X"D2",X"F7",X"0B",X"CD",X"6E",X"0C",X"C3",
		X"FA",X"0B",X"3A",X"3D",X"20",X"FE",X"18",X"C9",X"3A",X"3D",X"20",X"FE",X"20",X"C9",X"CD",X"62",
		X"0C",X"21",X"01",X"00",X"D0",X"2E",X"02",X"C9",X"21",X"40",X"20",X"3A",X"05",X"20",X"BE",X"DA",
		X"F7",X"0B",X"CD",X"8B",X"0C",X"CD",X"95",X"0C",X"C3",X"FA",X"0B",X"CD",X"62",X"0C",X"21",X"00",
		X"FE",X"D0",X"26",X"FD",X"C9",X"CD",X"68",X"0C",X"D8",X"26",X"FF",X"C9",X"21",X"3F",X"20",X"3A",
		X"04",X"20",X"BE",X"DA",X"F7",X"0B",X"CD",X"AC",X"0C",X"C3",X"FA",X"0B",X"CD",X"62",X"0C",X"21",
		X"FF",X"00",X"D0",X"2E",X"FE",X"C9",X"21",X"41",X"20",X"3A",X"05",X"20",X"BE",X"D2",X"F7",X"0B",
		X"CD",X"C9",X"0C",X"CD",X"D3",X"0C",X"C3",X"FA",X"0B",X"CD",X"62",X"0C",X"21",X"00",X"02",X"D0",
		X"26",X"03",X"C9",X"CD",X"68",X"0C",X"D8",X"26",X"01",X"C9",X"E7",X"2E",X"4B",X"7E",X"A7",X"21",
		X"00",X"03",X"C8",X"FE",X"01",X"26",X"04",X"C8",X"FE",X"02",X"26",X"05",X"C8",X"FE",X"03",X"26",
		X"06",X"C8",X"26",X"07",X"C9",X"CD",X"DA",X"0C",X"22",X"58",X"20",X"CD",X"42",X"0B",X"AF",X"BE",
		X"C8",X"0E",X"05",X"23",X"C5",X"E5",X"AF",X"BE",X"CA",X"48",X"0D",X"CD",X"09",X"0B",X"22",X"5A",
		X"20",X"21",X"5A",X"20",X"CD",X"0F",X"0B",X"21",X"5B",X"20",X"7E",X"FE",X"D8",X"D4",X"3D",X"0D",
		X"2A",X"5A",X"20",X"FF",X"3E",X"05",X"11",X"01",X"07",X"DF",X"21",X"58",X"20",X"EF",X"2A",X"5A",
		X"20",X"EB",X"E1",X"23",X"CD",X"15",X"0B",X"C1",X"0D",X"C2",X"04",X"0D",X"C9",X"E5",X"2A",X"5A",
		X"20",X"CD",X"1A",X"0B",X"E1",X"36",X"28",X"C9",X"CD",X"0D",X"1D",X"C3",X"32",X"0D",X"E7",X"2E",
		X"4C",X"7E",X"A7",X"21",X"00",X"FD",X"C8",X"FE",X"01",X"26",X"FC",X"C8",X"FE",X"02",X"26",X"FB",
		X"C8",X"FE",X"03",X"26",X"FA",X"C8",X"26",X"F9",X"C9",X"CD",X"4E",X"0D",X"22",X"60",X"20",X"CD",
		X"46",X"0B",X"AF",X"BE",X"C8",X"0E",X"05",X"23",X"C5",X"E5",X"AF",X"BE",X"CA",X"BC",X"0D",X"CD",
		X"09",X"0B",X"22",X"62",X"20",X"21",X"62",X"20",X"CD",X"0F",X"0B",X"21",X"63",X"20",X"7E",X"FE",
		X"30",X"DC",X"B1",X"0D",X"2A",X"62",X"20",X"FF",X"3E",X"04",X"11",X"01",X"07",X"DF",X"21",X"60",
		X"20",X"EF",X"2A",X"62",X"20",X"EB",X"E1",X"23",X"CD",X"15",X"0B",X"C1",X"0D",X"C2",X"78",X"0D",
		X"C9",X"E5",X"2A",X"62",X"20",X"CD",X"1A",X"0B",X"E1",X"36",X"D8",X"C9",X"CD",X"0D",X"1D",X"C3",
		X"A6",X"0D",X"21",X"4F",X"20",X"AF",X"BE",X"C8",X"23",X"BE",X"C2",X"20",X"10",X"23",X"BE",X"C2",
		X"E4",X"0D",X"34",X"23",X"BE",X"21",X"00",X"07",X"22",X"54",X"20",X"21",X"80",X"28",X"C4",X"12",
		X"0E",X"22",X"56",X"20",X"3A",X"52",X"20",X"A7",X"21",X"57",X"20",X"7E",X"C2",X"1C",X"0E",X"FE",
		X"D8",X"D2",X"24",X"0E",X"11",X"37",X"44",X"D5",X"2A",X"56",X"20",X"FF",X"3E",X"02",X"11",X"01",
		X"07",X"DF",X"01",X"01",X"18",X"D1",X"2A",X"56",X"20",X"CD",X"DA",X"03",X"21",X"54",X"20",X"C3",
		X"D8",X"02",X"21",X"00",X"F9",X"22",X"54",X"20",X"21",X"80",X"E0",X"C9",X"FE",X"28",X"DA",X"24",
		X"0E",X"C3",X"4C",X"0E",X"2A",X"56",X"20",X"CD",X"1A",X"0B",X"21",X"51",X"20",X"11",X"51",X"40",
		X"06",X"07",X"CD",X"BB",X"04",X"CD",X"52",X"0E",X"21",X"10",X"23",X"34",X"7E",X"E6",X"01",X"21",
		X"52",X"20",X"06",X"01",X"CC",X"49",X"0E",X"70",X"C9",X"06",X"00",X"C9",X"11",X"4F",X"44",X"C3",
		X"F7",X"0D",X"CD",X"ED",X"0E",X"21",X"50",X"20",X"36",X"08",X"FE",X"16",X"D0",X"FE",X"14",X"36",
		X"10",X"D0",X"FE",X"12",X"36",X"20",X"D0",X"FE",X"09",X"36",X"30",X"D0",X"FE",X"06",X"36",X"40",
		X"D0",X"FE",X"04",X"36",X"50",X"D0",X"36",X"60",X"C9",X"CD",X"ED",X"0E",X"FE",X"10",X"21",X"00",
		X"02",X"D0",X"21",X"00",X"01",X"C9",X"CD",X"79",X"0E",X"22",X"68",X"20",X"E7",X"2E",X"39",X"AF",
		X"BE",X"C8",X"0E",X"05",X"23",X"C5",X"E5",X"AF",X"BE",X"CA",X"E7",X"0E",X"CD",X"09",X"0B",X"22",
		X"6A",X"20",X"2A",X"6A",X"20",X"7C",X"D6",X"04",X"67",X"FF",X"3E",X"07",X"11",X"01",X"06",X"DF",
		X"21",X"6A",X"20",X"CD",X"0F",X"0B",X"21",X"6B",X"20",X"7E",X"FE",X"D8",X"D4",X"DC",X"0E",X"2A",
		X"6A",X"20",X"FF",X"3E",X"03",X"11",X"01",X"06",X"DF",X"21",X"68",X"20",X"EF",X"2A",X"6A",X"20",
		X"EB",X"E1",X"23",X"CD",X"15",X"0B",X"C1",X"0D",X"C2",X"95",X"0E",X"C9",X"E5",X"2A",X"6A",X"20",
		X"CD",X"1A",X"0B",X"E1",X"36",X"30",X"C9",X"CD",X"0D",X"1D",X"C3",X"D1",X"0E",X"E7",X"2E",X"4E",
		X"7E",X"C9",X"21",X"0A",X"20",X"AF",X"BE",X"C0",X"CD",X"05",X"04",X"E6",X"08",X"C2",X"0D",X"0F",
		X"21",X"0B",X"20",X"AF",X"BE",X"C2",X"0A",X"0F",X"34",X"C9",X"23",X"34",X"C9",X"21",X"0C",X"20",
		X"AF",X"BE",X"C8",X"36",X"00",X"2B",X"36",X"00",X"2E",X"0D",X"34",X"2E",X"39",X"34",X"2E",X"0F",
		X"AF",X"BE",X"C0",X"2E",X"F1",X"36",X"0A",X"21",X"0F",X"23",X"34",X"C9",X"21",X"0D",X"20",X"AF",
		X"BE",X"C8",X"23",X"BE",X"C2",X"20",X"10",X"23",X"BE",X"C2",X"47",X"0F",X"34",X"2A",X"04",X"20",
		X"01",X"0F",X"04",X"09",X"22",X"12",X"20",X"2A",X"12",X"20",X"CD",X"BC",X"0F",X"11",X"B4",X"42",
		X"CD",X"ED",X"08",X"3A",X"12",X"20",X"FE",X"F0",X"D2",X"B1",X"0F",X"21",X"10",X"20",X"06",X"02",
		X"FE",X"70",X"DA",X"67",X"0F",X"06",X"03",X"70",X"21",X"10",X"20",X"EF",X"2A",X"12",X"20",X"E5",
		X"FF",X"3E",X"06",X"11",X"02",X"02",X"DF",X"E1",X"06",X"03",X"11",X"B4",X"42",X"F7",X"C5",X"E5",
		X"1A",X"D3",X"03",X"DB",X"03",X"A6",X"CA",X"8E",X"0F",X"3E",X"01",X"32",X"38",X"20",X"DB",X"03",
		X"AE",X"77",X"23",X"13",X"AF",X"D3",X"03",X"DB",X"03",X"A6",X"CA",X"A2",X"0F",X"3E",X"01",X"32",
		X"38",X"20",X"DB",X"03",X"AE",X"77",X"E1",X"01",X"20",X"00",X"09",X"C1",X"05",X"C2",X"7E",X"0F",
		X"C9",X"21",X"0B",X"20",X"11",X"0B",X"40",X"06",X"09",X"C3",X"BB",X"04",X"7D",X"FE",X"7A",X"D2",
		X"CF",X"0F",X"C3",X"C5",X"0F",X"E5",X"FF",X"3E",X"07",X"11",X"02",X"02",X"DF",X"E1",X"C9",X"E5",
		X"FF",X"3E",X"02",X"C3",X"C9",X"0F",X"E5",X"FF",X"3E",X"06",X"C3",X"C9",X"0F",X"E5",X"FF",X"3E",
		X"04",X"C3",X"C9",X"0F",X"CD",X"D2",X"08",X"C0",X"2E",X"72",X"BE",X"C8",X"23",X"BE",X"C2",X"20",
		X"10",X"23",X"BE",X"C2",X"35",X"10",X"34",X"2A",X"70",X"20",X"4E",X"7D",X"FE",X"22",X"CC",X"22");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
