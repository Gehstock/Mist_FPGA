library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity prom_ic39 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of prom_ic39 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"42",X"42",X"7E",X"00",X"00",
		X"00",X"3C",X"42",X"42",X"42",X"42",X"3C",X"00",X"00",X"00",X"7E",X"42",X"42",X"00",X"00",X"00",
		X"00",X"08",X"04",X"7E",X"04",X"08",X"00",X"00",X"00",X"40",X"40",X"40",X"40",X"40",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"A0",X"B0",X"B8",X"BC",X"BC",X"BE",X"FE",X"00",X"C0",X"F8",X"F4",X"EC",X"DC",X"BE",X"FE",
		X"FE",X"80",X"FE",X"FC",X"F8",X"F0",X"C0",X"00",X"FE",X"BE",X"DC",X"EC",X"F4",X"F8",X"C0",X"00",
		X"FE",X"BE",X"BC",X"BC",X"B8",X"B0",X"A0",X"00",X"7F",X"7D",X"3B",X"37",X"2F",X"1F",X"03",X"00",
		X"7F",X"01",X"7F",X"3F",X"1F",X"0F",X"03",X"00",X"00",X"03",X"1F",X"2F",X"37",X"3B",X"7D",X"7F",
		X"FE",X"FE",X"FC",X"FC",X"F8",X"F0",X"C0",X"00",X"7F",X"7F",X"3F",X"3F",X"1F",X"0F",X"03",X"00",
		X"00",X"C0",X"F0",X"F8",X"FC",X"FC",X"FE",X"FE",X"00",X"03",X"0F",X"1F",X"3F",X"3F",X"7F",X"7F",
		X"3C",X"6E",X"FF",X"BB",X"FF",X"EF",X"7E",X"3C",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"A0",X"B0",X"B8",X"BC",X"BC",X"AE",X"FE",X"00",X"C0",X"F8",X"F4",X"AC",X"DC",X"AE",X"FE",
		X"FE",X"80",X"FE",X"BC",X"F8",X"F0",X"C0",X"00",X"FE",X"AE",X"DC",X"AC",X"F4",X"F8",X"C0",X"00",
		X"FE",X"AE",X"BC",X"BC",X"B8",X"B0",X"A0",X"00",X"7F",X"75",X"3B",X"35",X"2F",X"1F",X"03",X"00",
		X"7F",X"01",X"7F",X"3D",X"1F",X"0F",X"03",X"00",X"00",X"03",X"1F",X"2F",X"35",X"3B",X"75",X"7F",
		X"FE",X"EE",X"FC",X"BC",X"F8",X"F0",X"C0",X"00",X"7F",X"77",X"3F",X"3D",X"1F",X"0F",X"03",X"00",
		X"00",X"C0",X"F0",X"F8",X"BC",X"FC",X"EE",X"FE",X"00",X"03",X"0F",X"1F",X"3D",X"3F",X"77",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"7E",X"FF",X"FF",X"FF",X"FF",X"7E",X"3C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"7E",X"FF",X"FF",X"FF",X"FF",X"7E",X"3C",
		X"00",X"00",X"00",X"C0",X"00",X"00",X"08",X"04",X"00",X"02",X"00",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"20",X"10",X"00",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"10",X"01",X"08",X"00",X"0A",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"00",X"0A",
		X"80",X"10",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"08",X"00",X"00",
		X"00",X"00",X"01",X"07",X"00",X"10",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"00",X"80",X"10",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"0C",
		X"00",X"00",X"00",X"00",X"03",X"06",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"30",X"00",X"00",X"00",X"00",
		X"04",X"04",X"08",X"60",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"02",X"00",X"02",X"00",X"02",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0C",X"08",X"08",X"00",X"00",X"00",X"00",
		X"01",X"0F",X"00",X"88",X"10",X"80",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"00",X"40",X"70",X"00",X"00",X"08",X"01",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"F0",X"10",X"00",X"01",X"08",X"00",
		X"20",X"20",X"30",X"10",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"70",X"00",X"01",X"0A",X"00",X"08",X"01",
		X"10",X"F8",X"F0",X"F8",X"10",X"F0",X"40",X"00",X"09",X"19",X"09",X"19",X"0D",X"0F",X"19",X"30",
		X"00",X"00",X"00",X"00",X"04",X"4C",X"E8",X"F8",X"00",X"00",X"00",X"00",X"00",X"07",X"0D",X"19",
		X"40",X"E0",X"C0",X"60",X"40",X"C0",X"00",X"00",X"27",X"67",X"27",X"66",X"37",X"3F",X"65",X"C0",
		X"00",X"00",X"00",X"00",X"10",X"30",X"A0",X"60",X"00",X"00",X"00",X"00",X"00",X"1D",X"37",X"66",
		X"7E",X"74",X"66",X"7A",X"D3",X"01",X"00",X"00",X"06",X"02",X"06",X"03",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"50",X"FC",X"74",X"66",X"7C",X"00",X"00",X"0C",X"06",X"03",X"03",X"06",X"02",
		X"4E",X"7C",X"7E",X"5C",X"4E",X"7C",X"D6",X"03",X"06",X"02",X"06",X"02",X"06",X"03",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"50",X"FC",X"5C",X"00",X"00",X"00",X"00",X"08",X"08",X"0D",X"07",
		X"10",X"F0",X"48",X"04",X"00",X"00",X"00",X"00",X"0D",X"07",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"E0",X"F0",X"10",X"F8",X"F0",X"F8",X"20",X"17",X"0D",X"19",X"09",X"19",X"09",X"19",
		X"5C",X"FC",X"57",X"01",X"00",X"00",X"00",X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"D0",X"78",X"4C",X"5C",X"7E",X"7C",X"4E",X"0C",X"05",X"07",X"06",X"02",X"06",X"02",X"02",
		X"E0",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"67",X"25",X"24",X"77",X"5D",X"C0",X"00",X"00",
		X"00",X"00",X"10",X"30",X"E0",X"C0",X"E0",X"C0",X"00",X"00",X"00",X"05",X"1F",X"35",X"64",X"27",
		X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"26",X"77",X"DD",X"80",X"00",X"00",X"00",X"00",
		X"30",X"20",X"E0",X"40",X"60",X"C0",X"E0",X"40",X"00",X"05",X"1F",X"37",X"66",X"27",X"67",X"27",
		X"10",X"F8",X"F0",X"F8",X"10",X"F0",X"40",X"00",X"09",X"19",X"09",X"19",X"0D",X"0F",X"19",X"30",
		X"00",X"00",X"00",X"00",X"04",X"4C",X"E8",X"F8",X"00",X"00",X"00",X"00",X"00",X"07",X"0D",X"19",
		X"40",X"E0",X"C0",X"60",X"40",X"C0",X"00",X"00",X"27",X"67",X"27",X"66",X"37",X"3F",X"65",X"C0",
		X"00",X"00",X"00",X"00",X"10",X"30",X"A0",X"60",X"00",X"00",X"00",X"00",X"00",X"1D",X"37",X"66",
		X"7E",X"74",X"66",X"7A",X"D3",X"01",X"00",X"00",X"06",X"02",X"06",X"03",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"50",X"FC",X"74",X"66",X"7C",X"00",X"00",X"0C",X"06",X"03",X"03",X"06",X"02",
		X"4E",X"7C",X"7E",X"5C",X"4E",X"7C",X"D6",X"03",X"06",X"02",X"06",X"02",X"06",X"03",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"50",X"FC",X"5C",X"00",X"00",X"00",X"00",X"08",X"08",X"0D",X"07",
		X"10",X"F0",X"48",X"04",X"00",X"00",X"00",X"00",X"0D",X"07",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"E0",X"F0",X"10",X"F8",X"F0",X"F8",X"20",X"17",X"0D",X"19",X"09",X"19",X"09",X"19",
		X"5C",X"FC",X"57",X"01",X"00",X"00",X"00",X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"D0",X"78",X"4C",X"5C",X"7E",X"7C",X"4E",X"0C",X"05",X"07",X"06",X"02",X"06",X"02",X"02",
		X"E0",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"67",X"25",X"24",X"77",X"5D",X"C0",X"00",X"00",
		X"00",X"00",X"10",X"30",X"E0",X"C0",X"E0",X"C0",X"00",X"00",X"00",X"05",X"1F",X"35",X"64",X"27",
		X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"26",X"77",X"DD",X"80",X"00",X"00",X"00",X"00",
		X"30",X"20",X"E0",X"40",X"60",X"C0",X"E0",X"40",X"00",X"05",X"1F",X"37",X"66",X"27",X"67",X"27",
		X"00",X"00",X"00",X"C0",X"00",X"00",X"08",X"04",X"00",X"02",X"00",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"20",X"10",X"00",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"10",X"01",X"08",X"00",X"0A",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"00",X"0A",
		X"80",X"10",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"08",X"00",X"00",
		X"00",X"00",X"01",X"07",X"00",X"10",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"00",X"80",X"10",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"0C",
		X"00",X"00",X"00",X"00",X"03",X"06",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"30",X"00",X"00",X"00",X"00",
		X"04",X"04",X"08",X"60",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"02",X"00",X"02",X"00",X"02",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0C",X"08",X"08",X"00",X"00",X"00",X"00",
		X"01",X"0F",X"00",X"88",X"10",X"80",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"00",X"40",X"70",X"00",X"00",X"08",X"01",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"F0",X"10",X"00",X"01",X"08",X"00",
		X"20",X"20",X"30",X"10",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"70",X"00",X"01",X"0A",X"00",X"08",X"01",
		X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"FF",X"FF",X"00",X"FF",X"FF",X"00",X"FF",X"FF",
		X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"FF",X"FF",X"00",X"FF",X"FF",X"00",X"FF",X"FF",
		X"DB",X"DB",X"1B",X"FB",X"F3",X"07",X"FE",X"FC",X"FC",X"FE",X"07",X"F3",X"FB",X"1B",X"DB",X"DB",
		X"DB",X"DB",X"D8",X"DF",X"CF",X"E0",X"7F",X"3F",X"3F",X"7F",X"E0",X"CF",X"DF",X"D8",X"DB",X"DB",
		X"DB",X"DB",X"1B",X"FB",X"F3",X"07",X"FE",X"FC",X"FC",X"FE",X"07",X"F3",X"FB",X"1B",X"DB",X"DB",
		X"DB",X"DB",X"D8",X"DF",X"CF",X"E0",X"7F",X"3F",X"3F",X"7F",X"E0",X"CF",X"DF",X"D8",X"DB",X"DB",
		X"7E",X"C3",X"81",X"A5",X"A5",X"99",X"C3",X"7E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"7E",X"04",X"08",X"08",X"04",X"7E",X"00",X"00",X"42",X"42",X"7E",X"42",X"42",X"00",X"00",
		X"00",X"24",X"42",X"42",X"42",X"42",X"3C",X"00",X"00",X"44",X"2A",X"1A",X"0A",X"0A",X"7E",X"00",
		X"00",X"3C",X"42",X"42",X"42",X"42",X"3C",X"00",X"00",X"02",X"02",X"7E",X"02",X"02",X"00",X"00",
		X"00",X"44",X"2A",X"1A",X"0A",X"0A",X"7E",X"00",X"00",X"7C",X"12",X"12",X"12",X"12",X"7C",X"00",
		X"00",X"42",X"42",X"7E",X"42",X"42",X"00",X"00",X"00",X"7E",X"20",X"10",X"08",X"04",X"7E",X"00",
		X"00",X"3C",X"42",X"66",X"66",X"5A",X"3C",X"00",X"00",X"8E",X"91",X"E6",X"00",X"76",X"89",X"76",
		X"00",X"7E",X"42",X"5A",X"5A",X"42",X"7E",X"00",X"FF",X"81",X"BD",X"A5",X"A5",X"BD",X"81",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"88",X"14",X"2A",X"49",X"BE",X"49",X"2A",X"14");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
