library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_SND_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_SND_1 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"80",X"32",X"0B",X"80",X"C9",X"AF",X"32",X"00",X"80",X"32",X"01",X"80",X"C9",X"AF",X"32",X"02",
		X"80",X"32",X"03",X"80",X"C9",X"AF",X"32",X"04",X"80",X"32",X"05",X"80",X"C9",X"AF",X"32",X"06",
		X"80",X"32",X"07",X"80",X"C9",X"AF",X"32",X"08",X"80",X"32",X"09",X"80",X"C9",X"00",X"00",X"06",
		X"09",X"06",X"09",X"06",X"09",X"06",X"09",X"06",X"09",X"DA",X"0C",X"3E",X"10",X"BD",X"11",X"A6",
		X"0F",X"AD",X"0F",X"B4",X"0F",X"D5",X"0F",X"DC",X"0F",X"E3",X"0F",X"FF",X"0F",X"06",X"10",X"50",
		X"12",X"00",X"00",X"33",X"0B",X"D0",X"0B",X"5F",X"0C",X"67",X"13",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"0D",X"B7",
		X"14",X"A5",X"16",X"CD",X"10",X"4A",X"11",X"22",X"13",X"E9",X"13",X"E9",X"13",X"A5",X"16",X"A5",
		X"16",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CD",X"ED",X"0A",
		X"3E",X"03",X"32",X"1B",X"80",X"3E",X"0F",X"32",X"1C",X"80",X"3E",X"1F",X"32",X"1D",X"80",X"21",
		X"80",X"00",X"22",X"1E",X"80",X"22",X"20",X"80",X"3E",X"04",X"32",X"22",X"80",X"3E",X"40",X"32",
		X"23",X"80",X"32",X"24",X"80",X"3E",X"03",X"32",X"26",X"80",X"3E",X"0A",X"32",X"27",X"80",X"21",
		X"00",X"08",X"22",X"28",X"80",X"3E",X"08",X"32",X"2A",X"80",X"32",X"2B",X"80",X"21",X"40",X"00",
		X"22",X"2C",X"80",X"22",X"2E",X"80",X"3E",X"0C",X"32",X"30",X"80",X"3E",X"03",X"32",X"32",X"80",
		X"3E",X"0A",X"32",X"33",X"80",X"21",X"00",X"02",X"22",X"34",X"80",X"21",X"00",X"08",X"22",X"36",
		X"80",X"21",X"00",X"02",X"22",X"38",X"80",X"3E",X"08",X"32",X"3A",X"80",X"32",X"3B",X"80",X"21",
		X"20",X"00",X"22",X"3D",X"80",X"C9",X"3E",X"FF",X"C9",X"CD",X"ED",X"0A",X"3E",X"03",X"32",X"1B",
		X"80",X"3E",X"0F",X"32",X"1C",X"80",X"3E",X"1F",X"32",X"1D",X"80",X"21",X"80",X"00",X"22",X"1E",
		X"80",X"22",X"20",X"80",X"3E",X"01",X"32",X"22",X"80",X"3E",X"20",X"32",X"23",X"80",X"32",X"24",
		X"80",X"3E",X"03",X"32",X"26",X"80",X"3E",X"0D",X"32",X"27",X"80",X"21",X"00",X"08",X"22",X"28",
		X"80",X"3E",X"08",X"32",X"2A",X"80",X"32",X"2B",X"80",X"21",X"40",X"00",X"22",X"2C",X"80",X"22",
		X"2E",X"80",X"3E",X"02",X"32",X"30",X"80",X"3E",X"03",X"32",X"32",X"80",X"3E",X"0E",X"32",X"33",
		X"80",X"21",X"00",X"02",X"22",X"34",X"80",X"21",X"00",X"08",X"22",X"36",X"80",X"21",X"01",X"00",
		X"22",X"38",X"80",X"3E",X"18",X"32",X"3A",X"80",X"32",X"3B",X"80",X"21",X"00",X"01",X"22",X"3D",
		X"80",X"C9",X"CD",X"ED",X"0A",X"3E",X"02",X"32",X"1B",X"80",X"3E",X"0F",X"32",X"1C",X"80",X"3E",
		X"08",X"32",X"1D",X"80",X"21",X"80",X"00",X"22",X"1E",X"80",X"22",X"20",X"80",X"3E",X"01",X"32",
		X"22",X"80",X"3E",X"20",X"32",X"23",X"80",X"32",X"24",X"80",X"3E",X"03",X"32",X"26",X"80",X"3E",
		X"0A",X"32",X"27",X"80",X"21",X"00",X"08",X"22",X"28",X"80",X"3E",X"08",X"32",X"2A",X"80",X"32",
		X"2B",X"80",X"21",X"40",X"00",X"22",X"2C",X"80",X"22",X"2E",X"80",X"3E",X"03",X"32",X"30",X"80",
		X"3E",X"03",X"32",X"32",X"80",X"3E",X"08",X"32",X"33",X"80",X"21",X"00",X"02",X"22",X"34",X"80",
		X"21",X"00",X"08",X"22",X"36",X"80",X"21",X"01",X"00",X"22",X"38",X"80",X"3E",X"20",X"32",X"3A",
		X"80",X"32",X"3B",X"80",X"21",X"20",X"00",X"22",X"3D",X"80",X"C9",X"CD",X"ED",X"0A",X"3E",X"03",
		X"32",X"1B",X"80",X"3E",X"0E",X"32",X"1C",X"80",X"3E",X"1F",X"32",X"1D",X"80",X"21",X"80",X"00",
		X"22",X"1E",X"80",X"22",X"20",X"80",X"3E",X"01",X"32",X"22",X"80",X"3E",X"20",X"32",X"23",X"80",
		X"32",X"24",X"80",X"3E",X"03",X"32",X"26",X"80",X"3E",X"0C",X"32",X"27",X"80",X"21",X"00",X"08",
		X"22",X"28",X"80",X"3E",X"08",X"32",X"2A",X"80",X"32",X"2B",X"80",X"21",X"40",X"00",X"22",X"2C",
		X"80",X"22",X"2E",X"80",X"3E",X"03",X"32",X"30",X"80",X"3E",X"03",X"32",X"32",X"80",X"3E",X"0F",
		X"32",X"33",X"80",X"21",X"00",X"02",X"22",X"34",X"80",X"21",X"00",X"08",X"22",X"36",X"80",X"21",
		X"01",X"00",X"22",X"38",X"80",X"3E",X"20",X"32",X"3A",X"80",X"32",X"3B",X"80",X"21",X"20",X"00",
		X"22",X"3D",X"80",X"C9",X"CD",X"ED",X"0A",X"3E",X"03",X"32",X"1B",X"80",X"3E",X"0F",X"32",X"1C",
		X"80",X"3E",X"1F",X"32",X"1D",X"80",X"21",X"80",X"00",X"22",X"1E",X"80",X"22",X"20",X"80",X"3E",
		X"04",X"32",X"22",X"80",X"3E",X"40",X"32",X"23",X"80",X"32",X"24",X"80",X"3E",X"03",X"32",X"26",
		X"80",X"3E",X"0C",X"32",X"27",X"80",X"21",X"00",X"08",X"22",X"28",X"80",X"3E",X"08",X"32",X"2A",
		X"80",X"32",X"2B",X"80",X"21",X"30",X"00",X"22",X"2C",X"80",X"22",X"2E",X"80",X"3E",X"08",X"32",
		X"30",X"80",X"3E",X"03",X"32",X"32",X"80",X"3E",X"09",X"32",X"33",X"80",X"21",X"00",X"02",X"22",
		X"34",X"80",X"21",X"00",X"08",X"22",X"36",X"80",X"21",X"00",X"01",X"22",X"38",X"80",X"3E",X"01",
		X"32",X"3A",X"80",X"32",X"3B",X"80",X"21",X"20",X"00",X"22",X"3D",X"80",X"C9",X"3E",X"13",X"CD",
		X"6A",X"00",X"3E",X"14",X"CD",X"6A",X"00",X"3E",X"15",X"CD",X"6A",X"00",X"C9",X"3A",X"1B",X"80",
		X"B7",X"28",X"21",X"FE",X"01",X"28",X"22",X"FE",X"02",X"28",X"23",X"CD",X"96",X"07",X"AF",X"32",
		X"25",X"80",X"16",X"06",X"21",X"1D",X"80",X"5E",X"CD",X"34",X"05",X"CD",X"68",X"05",X"06",X"00",
		X"CD",X"D8",X"05",X"C9",X"CD",X"A1",X"06",X"18",X"E5",X"CD",X"22",X"07",X"18",X"E0",X"CD",X"5C",
		X"07",X"18",X"DB",X"16",X"06",X"21",X"1D",X"80",X"5E",X"CD",X"34",X"05",X"3A",X"25",X"80",X"B7",
		X"28",X"1E",X"FE",X"01",X"28",X"27",X"FE",X"02",X"28",X"3C",X"21",X"24",X"80",X"35",X"20",X"0E",
		X"3A",X"23",X"80",X"77",X"CD",X"25",X"06",X"3D",X"28",X"3E",X"47",X"CD",X"D8",X"05",X"AF",X"C9",
		X"3A",X"1C",X"80",X"47",X"CD",X"D8",X"05",X"21",X"25",X"80",X"34",X"18",X"DD",X"2A",X"20",X"80",
		X"2B",X"7C",X"B5",X"20",X"0C",X"2A",X"1E",X"80",X"22",X"20",X"80",X"21",X"25",X"80",X"34",X"18",
		X"C9",X"22",X"20",X"80",X"18",X"C4",X"21",X"22",X"80",X"35",X"20",X"06",X"21",X"25",X"80",X"34",
		X"18",X"B8",X"AF",X"32",X"25",X"80",X"18",X"B2",X"16",X"06",X"1E",X"04",X"CD",X"34",X"05",X"3E",
		X"FF",X"C9",X"3A",X"26",X"80",X"B7",X"28",X"19",X"FE",X"01",X"28",X"1A",X"FE",X"02",X"28",X"1B",
		X"CD",X"96",X"07",X"AF",X"32",X"31",X"80",X"2A",X"28",X"80",X"CD",X"B3",X"04",X"CD",X"FA",X"04",
		X"C9",X"CD",X"A1",X"06",X"18",X"ED",X"CD",X"22",X"07",X"18",X"E8",X"CD",X"5C",X"07",X"18",X"E3",
		X"3A",X"31",X"80",X"B7",X"28",X"1F",X"FE",X"01",X"28",X"2E",X"2A",X"2E",X"80",X"2B",X"7C",X"B5",
		X"20",X"40",X"2A",X"2C",X"80",X"22",X"2E",X"80",X"21",X"30",X"80",X"35",X"28",X"39",X"21",X"31",
		X"80",X"36",X"00",X"AF",X"C9",X"3A",X"27",X"80",X"47",X"CD",X"D8",X"05",X"3A",X"2A",X"80",X"32",
		X"2B",X"80",X"21",X"31",X"80",X"34",X"18",X"EB",X"21",X"2B",X"80",X"35",X"20",X"CC",X"3A",X"2A",
		X"80",X"77",X"CD",X"25",X"06",X"3D",X"20",X"04",X"21",X"31",X"80",X"34",X"47",X"CD",X"D8",X"05",
		X"18",X"B8",X"22",X"2E",X"80",X"18",X"CC",X"3E",X"FF",X"C9",X"3A",X"32",X"80",X"B7",X"28",X"20",
		X"FE",X"01",X"28",X"21",X"FE",X"02",X"28",X"22",X"CD",X"96",X"07",X"AF",X"32",X"3C",X"80",X"2A",
		X"36",X"80",X"CD",X"B3",X"04",X"CD",X"FA",X"04",X"3A",X"33",X"80",X"47",X"CD",X"D8",X"05",X"C9",
		X"CD",X"A1",X"06",X"18",X"E6",X"CD",X"22",X"07",X"18",X"E1",X"CD",X"5C",X"07",X"18",X"DC",X"3A",
		X"3C",X"80",X"B7",X"28",X"22",X"FE",X"01",X"28",X"32",X"CD",X"5A",X"06",X"B7",X"ED",X"5B",X"3D",
		X"80",X"ED",X"52",X"ED",X"5B",X"34",X"80",X"7C",X"BA",X"20",X"07",X"7D",X"BB",X"20",X"03",X"2A",
		X"36",X"80",X"CD",X"B3",X"04",X"AF",X"C9",X"2A",X"38",X"80",X"2B",X"7C",X"B5",X"20",X"07",X"3E",
		X"01",X"32",X"3C",X"80",X"18",X"D3",X"22",X"38",X"80",X"18",X"CE",X"21",X"3A",X"80",X"35",X"20",
		X"C8",X"3A",X"3B",X"80",X"77",X"CD",X"25",X"06",X"3D",X"28",X"06",X"47",X"CD",X"D8",X"05",X"18",
		X"B8",X"3E",X"FF",X"C9",X"CD",X"22",X"07",X"AF",X"32",X"43",X"80",X"3E",X"02",X"32",X"42",X"80",
		X"CD",X"FA",X"04",X"3E",X"08",X"32",X"3F",X"80",X"21",X"20",X"00",X"22",X"40",X"80",X"21",X"40",
		X"00",X"CD",X"B3",X"04",X"06",X"08",X"CD",X"D8",X"05",X"C9",X"3A",X"43",X"80",X"B7",X"20",X"0B",
		X"2A",X"40",X"80",X"2B",X"7C",X"B5",X"28",X"35",X"22",X"40",X"80",X"21",X"3F",X"80",X"35",X"28",
		X"1A",X"CD",X"5A",X"06",X"11",X"10",X"00",X"19",X"11",X"00",X"02",X"7C",X"BA",X"20",X"07",X"7D",
		X"BB",X"20",X"03",X"21",X"40",X"00",X"CD",X"B3",X"04",X"AF",X"C9",X"3E",X"08",X"32",X"3F",X"80",
		X"CD",X"25",X"06",X"47",X"3E",X"FF",X"05",X"C8",X"CD",X"D8",X"05",X"18",X"D4",X"21",X"20",X"00",
		X"22",X"40",X"80",X"21",X"42",X"80",X"35",X"20",X"05",X"3E",X"01",X"32",X"43",X"80",X"CD",X"C3",
		X"0C",X"18",X"A7",X"CD",X"5C",X"07",X"3E",X"08",X"32",X"44",X"80",X"21",X"00",X"0A",X"22",X"45",
		X"80",X"21",X"40",X"00",X"CD",X"B3",X"04",X"CD",X"FA",X"04",X"06",X"0B",X"CD",X"D8",X"05",X"C9",
		X"2A",X"45",X"80",X"2B",X"22",X"45",X"80",X"7C",X"B5",X"3E",X"FF",X"C8",X"3C",X"21",X"44",X"80",
		X"35",X"C0",X"36",X"08",X"CD",X"5A",X"06",X"11",X"02",X"00",X"19",X"CD",X"B3",X"04",X"AF",X"C9",
		X"DD",X"7E",X"00",X"FE",X"FF",X"C8",X"CD",X"7B",X"0D",X"AF",X"C9",X"DD",X"35",X"01",X"C0",X"3A",
		X"72",X"80",X"DD",X"77",X"01",X"DD",X"CB",X"00",X"46",X"C2",X"9B",X"0D",X"DD",X"7E",X"07",X"D6",
		X"01",X"FA",X"9B",X"0D",X"DD",X"77",X"07",X"47",X"CD",X"D8",X"05",X"DD",X"35",X"00",X"C0",X"DD",
		X"6E",X"02",X"DD",X"66",X"03",X"7E",X"47",X"E6",X"1F",X"CA",X"36",X"0E",X"FE",X"1F",X"C2",X"52",
		X"0E",X"23",X"DD",X"75",X"02",X"DD",X"74",X"03",X"78",X"E6",X"E0",X"0F",X"0F",X"0F",X"0F",X"4F",
		X"06",X"00",X"21",X"CB",X"0D",X"09",X"5E",X"23",X"56",X"EB",X"E9",X"DB",X"0D",X"F9",X"0D",X"0F",
		X"0E",X"2C",X"0E",X"2C",X"0E",X"2C",X"0E",X"2C",X"0E",X"2C",X"0E",X"DD",X"6E",X"02",X"DD",X"66",
		X"03",X"4E",X"CB",X"21",X"06",X"00",X"21",X"85",X"0E",X"09",X"5E",X"23",X"56",X"ED",X"53",X"70",
		X"80",X"DD",X"73",X"04",X"DD",X"72",X"05",X"18",X"23",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"4E",
		X"06",X"00",X"21",X"1D",X"0F",X"09",X"7E",X"32",X"72",X"80",X"DD",X"77",X"01",X"18",X"0D",X"DD",
		X"6E",X"02",X"DD",X"66",X"03",X"7E",X"DD",X"77",X"06",X"DD",X"77",X"07",X"DD",X"6E",X"02",X"DD",
		X"66",X"03",X"23",X"DD",X"75",X"02",X"DD",X"74",X"03",X"C3",X"9F",X"0D",X"06",X"00",X"CD",X"D8",
		X"05",X"DD",X"36",X"00",X"FF",X"C9",X"CD",X"40",X"0E",X"06",X"00",X"CD",X"D8",X"05",X"18",X"37",
		X"78",X"E6",X"E0",X"07",X"07",X"07",X"47",X"3E",X"01",X"18",X"01",X"07",X"10",X"FD",X"DD",X"77",
		X"00",X"C9",X"C5",X"CD",X"40",X"0E",X"C1",X"78",X"E6",X"1F",X"3D",X"07",X"4F",X"06",X"00",X"DD",
		X"6E",X"04",X"DD",X"66",X"05",X"09",X"5E",X"23",X"56",X"EB",X"CD",X"B3",X"04",X"DD",X"46",X"06",
		X"78",X"DD",X"77",X"07",X"CD",X"D8",X"05",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"23",X"DD",X"75",
		X"02",X"DD",X"74",X"03",X"C9",X"A5",X"0E",X"A9",X"0E",X"AD",X"0E",X"B1",X"0E",X"B5",X"0E",X"B9",
		X"0E",X"BD",X"0E",X"C1",X"0E",X"C5",X"0E",X"C9",X"0E",X"CD",X"0E",X"D1",X"0E",X"D5",X"0E",X"D9",
		X"0E",X"DD",X"0E",X"E1",X"0E",X"6B",X"08",X"F2",X"07",X"80",X"07",X"14",X"07",X"AE",X"06",X"4E",
		X"06",X"F3",X"05",X"9E",X"05",X"4E",X"05",X"01",X"05",X"B9",X"04",X"76",X"04",X"36",X"04",X"F9",
		X"03",X"C0",X"03",X"8A",X"03",X"57",X"03",X"27",X"03",X"FA",X"02",X"CF",X"02",X"A7",X"02",X"81",
		X"02",X"5D",X"02",X"3B",X"02",X"1B",X"02",X"FD",X"01",X"E0",X"01",X"C5",X"01",X"AC",X"01",X"94",
		X"01",X"7D",X"01",X"68",X"01",X"53",X"01",X"40",X"01",X"2E",X"01",X"1D",X"01",X"0D",X"01",X"FE",
		X"00",X"F0",X"00",X"E3",X"00",X"D6",X"00",X"CA",X"00",X"BE",X"00",X"B4",X"00",X"AA",X"00",X"A0",
		X"00",X"97",X"00",X"8F",X"00",X"87",X"00",X"7F",X"00",X"78",X"00",X"71",X"00",X"6B",X"00",X"65",
		X"00",X"5F",X"00",X"5A",X"00",X"55",X"00",X"50",X"00",X"4C",X"00",X"47",X"00",X"57",X"42",X"34",
		X"2C",X"25",X"21",X"1D",X"1A",X"0C",X"0B",X"0A",X"09",X"08",X"07",X"06",X"05",X"21",X"60",X"0F",
		X"11",X"50",X"80",X"01",X"18",X"00",X"ED",X"B0",X"3A",X"73",X"80",X"07",X"4F",X"07",X"07",X"91",
		X"4F",X"06",X"00",X"21",X"78",X"0F",X"09",X"11",X"52",X"80",X"CD",X"56",X"0F",X"11",X"5A",X"80",
		X"CD",X"56",X"0F",X"11",X"62",X"80",X"7E",X"12",X"CD",X"5D",X"0F",X"7E",X"12",X"23",X"13",X"C9",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"75",X"15",X"9C",X"15",X"C3",X"15",X"C4",X"15",
		X"E0",X"15",X"FB",X"15",X"17",X"16",X"4B",X"16",X"64",X"16",X"CD",X"A1",X"06",X"AF",X"32",X"73",
		X"80",X"CD",X"FA",X"04",X"CD",X"2D",X"0F",X"C9",X"CD",X"A1",X"06",X"CD",X"FA",X"04",X"C9",X"CD",
		X"A1",X"06",X"CD",X"FA",X"04",X"C9",X"DD",X"21",X"50",X"80",X"C3",X"70",X"0D",X"DD",X"21",X"58",
		X"80",X"C3",X"70",X"0D",X"DD",X"21",X"60",X"80",X"C3",X"70",X"0D",X"CD",X"A1",X"06",X"3E",X"01",
		X"32",X"73",X"80",X"CD",X"FA",X"04",X"C3",X"2D",X"0F",X"CD",X"A1",X"06",X"C3",X"FA",X"04",X"CD",
		X"A1",X"06",X"C3",X"FA",X"04",X"DD",X"21",X"50",X"80",X"C3",X"70",X"0D",X"DD",X"21",X"58",X"80",
		X"C3",X"70",X"0D",X"DD",X"21",X"60",X"80",X"C3",X"70",X"0D",X"CD",X"A1",X"06",X"3E",X"02",X"32",
		X"73",X"80",X"CD",X"FA",X"04",X"C3",X"2D",X"0F",X"CD",X"A1",X"06",X"CD",X"FA",X"04",X"C9",X"DD");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
