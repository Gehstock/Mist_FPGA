library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity SL31254 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(9 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of SL31254 is
	type rom is array(0 to  1023) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"04",X"9C",X"64",X"6A",X"41",X"50",X"25",X"5C",X"81",X"07",X"28",X"04",X"3F",X"20",X"5C",X"51",
		X"41",X"50",X"25",X"14",X"91",X"07",X"28",X"04",X"3F",X"20",X"14",X"51",X"6B",X"42",X"50",X"25",
		X"08",X"91",X"07",X"28",X"04",X"3F",X"20",X"09",X"52",X"42",X"50",X"25",X"2E",X"81",X"07",X"28",
		X"04",X"3F",X"20",X"2E",X"52",X"20",X"55",X"50",X"28",X"06",X"79",X"28",X"01",X"1E",X"0C",X"4C",
		X"18",X"1F",X"5C",X"20",X"40",X"B5",X"1C",X"08",X"28",X"01",X"07",X"20",X"36",X"51",X"7A",X"52",
		X"75",X"54",X"20",X"81",X"50",X"28",X"06",X"79",X"41",X"24",X"FA",X"51",X"42",X"24",X"08",X"52",
		X"34",X"94",X"F0",X"28",X"01",X"1E",X"0C",X"08",X"28",X"01",X"07",X"67",X"68",X"4C",X"22",X"00",
		X"84",X"27",X"70",X"5C",X"6A",X"71",X"50",X"18",X"DC",X"24",X"66",X"D0",X"5C",X"25",X"99",X"94",
		X"15",X"20",X"59",X"5E",X"71",X"50",X"18",X"DC",X"24",X"66",X"D0",X"25",X"99",X"94",X"06",X"28",
		X"02",X"24",X"90",X"05",X"5C",X"28",X"02",X"71",X"28",X"01",X"1E",X"0C",X"08",X"28",X"01",X"07",
		X"64",X"6F",X"71",X"FC",X"84",X"13",X"62",X"6C",X"28",X"05",X"FC",X"30",X"84",X"3B",X"62",X"69",
		X"28",X"05",X"FC",X"30",X"84",X"30",X"90",X"11",X"62",X"69",X"28",X"05",X"FC",X"30",X"84",X"26",
		X"62",X"6C",X"28",X"05",X"FC",X"30",X"84",X"21",X"64",X"6D",X"4C",X"21",X"04",X"94",X"04",X"29",
		X"05",X"9D",X"63",X"68",X"28",X"05",X"FC",X"30",X"84",X"7C",X"63",X"6A",X"28",X"05",X"FC",X"30",
		X"84",X"78",X"29",X"05",X"88",X"68",X"90",X"02",X"6B",X"62",X"4D",X"54",X"4D",X"4C",X"57",X"64",
		X"6D",X"4C",X"13",X"44",X"81",X"21",X"2A",X"05",X"0E",X"77",X"54",X"37",X"37",X"44",X"C7",X"53",
		X"42",X"18",X"1F",X"C3",X"84",X"04",X"34",X"81",X"F5",X"44",X"8E",X"16",X"90",X"0B",X"04",X"04",
		X"05",X"06",X"00",X"01",X"02",X"03",X"24",X"E9",X"2A",X"05",X"47",X"13",X"8E",X"16",X"55",X"16",
		X"56",X"64",X"6A",X"4C",X"22",X"00",X"91",X"13",X"45",X"18",X"1F",X"55",X"6D",X"4C",X"13",X"6A",
		X"91",X"05",X"46",X"18",X"1F",X"56",X"41",X"24",X"02",X"51",X"45",X"5D",X"46",X"5D",X"72",X"5C",
		X"20",X"80",X"B5",X"28",X"01",X"1E",X"0C",X"02",X"00",X"02",X"01",X"02",X"02",X"01",X"02",X"01",
		X"FE",X"02",X"FE",X"02",X"FF",X"71",X"53",X"90",X"03",X"72",X"53",X"64",X"6A",X"4C",X"33",X"84",
		X"07",X"22",X"00",X"81",X"07",X"90",X"08",X"22",X"00",X"81",X"04",X"18",X"1F",X"5C",X"20",X"80",
		X"B5",X"6B",X"4C",X"22",X"00",X"94",X"10",X"62",X"69",X"4C",X"21",X"01",X"84",X"04",X"72",X"90",
		X"03",X"20",X"FE",X"64",X"6B",X"5C",X"90",X"6C",X"42",X"25",X"14",X"81",X"0E",X"25",X"24",X"91",
		X"0A",X"41",X"25",X"14",X"81",X"14",X"25",X"5C",X"91",X"10",X"29",X"05",X"43",X"41",X"25",X"14",
		X"81",X"08",X"25",X"5C",X"91",X"04",X"29",X"05",X"43",X"64",X"6A",X"4D",X"13",X"91",X"05",X"24",
		X"02",X"90",X"03",X"24",X"FE",X"C1",X"51",X"6B",X"4C",X"C2",X"52",X"20",X"55",X"50",X"28",X"06",
		X"79",X"64",X"6B",X"70",X"5C",X"64",X"68",X"4C",X"25",X"30",X"91",X"06",X"28",X"02",X"B5",X"90",
		X"04",X"28",X"02",X"AC",X"20",X"FF",X"55",X"28",X"00",X"8F",X"63",X"6F",X"4C",X"25",X"02",X"94",
		X"10",X"62",X"6E",X"4D",X"25",X"15",X"84",X"06",X"4C",X"25",X"15",X"94",X"04",X"28",X"02",X"24",
		X"28",X"01",X"A0",X"28",X"01",X"1E",X"28",X"01",X"1E",X"29",X"00",X"37",X"08",X"28",X"01",X"07",
		X"4C",X"18",X"1F",X"C1",X"91",X"0B",X"4C",X"24",X"05",X"56",X"41",X"18",X"1F",X"CC",X"81",X"17",
		X"4C",X"18",X"1F",X"56",X"41",X"24",X"02",X"C6",X"91",X"36",X"41",X"24",X"02",X"18",X"1F",X"56",
		X"4C",X"24",X"05",X"C6",X"91",X"2A",X"4D",X"4C",X"18",X"1F",X"56",X"42",X"C6",X"91",X"0B",X"42",
		X"18",X"1F",X"56",X"4C",X"24",X"05",X"C6",X"81",X"1D",X"4C",X"18",X"1F",X"56",X"42",X"24",X"02",
		X"C6",X"91",X"0D",X"42",X"24",X"02",X"18",X"1F",X"56",X"4C",X"24",X"05",X"C6",X"81",X"07",X"70",
		X"50",X"28",X"01",X"1E",X"0C",X"71",X"90",X"F9",X"2A",X"06",X"74",X"64",X"6D",X"4C",X"21",X"20",
		X"84",X"12",X"66",X"6F",X"3C",X"94",X"0D",X"63",X"6C",X"4C",X"12",X"8E",X"16",X"66",X"6F",X"5D",
		X"67",X"71",X"5C",X"1C",X"09",X"0D",X"15",X"1C",X"1C",X"2A",X"07",X"67",X"08",X"28",X"01",X"07",
		X"0A",X"66",X"6C",X"5D",X"43",X"5D",X"44",X"5C",X"75",X"54",X"20",X"C0",X"F0",X"53",X"20",X"3F",
		X"F0",X"50",X"25",X"15",X"94",X"1F",X"64",X"68",X"72",X"54",X"28",X"06",X"EC",X"20",X"15",X"50",
		X"28",X"07",X"18",X"41",X"24",X"06",X"51",X"66",X"6D",X"4D",X"53",X"4C",X"54",X"6C",X"4C",X"0B",
		X"28",X"01",X"1E",X"0C",X"25",X"30",X"94",X"0B",X"62",X"69",X"28",X"06",X"EC",X"68",X"4D",X"50",
		X"90",X"DF",X"25",X"31",X"94",X"0B",X"62",X"6C",X"28",X"06",X"EC",X"6B",X"4D",X"50",X"90",X"D1",
		X"25",X"32",X"94",X"0B",X"63",X"68",X"28",X"06",X"EC",X"20",X"14",X"50",X"90",X"C3",X"25",X"33",
		X"94",X"BF",X"63",X"6A",X"28",X"06",X"EC",X"20",X"14",X"50",X"90",X"B5",X"08",X"28",X"01",X"07",
		X"4C",X"E1",X"94",X"06",X"4D",X"4E",X"E2",X"84",X"1C",X"41",X"55",X"42",X"56",X"4C",X"51",X"45",
		X"5D",X"4C",X"52",X"46",X"5E",X"7D",X"50",X"2A",X"07",X"67",X"28",X"07",X"18",X"2A",X"07",X"67",
		X"4D",X"51",X"4E",X"52",X"28",X"01",X"1E",X"0C",X"40",X"13",X"8E",X"C0",X"8E",X"20",X"40",X"B0",
		X"44",X"56",X"55",X"16",X"57",X"42",X"24",X"00",X"18",X"21",X"3F",X"58",X"A5",X"21",X"C0",X"C8",
		X"B5",X"41",X"24",X"FC",X"18",X"B4",X"47",X"22",X"00",X"43",X"91",X"02",X"70",X"18",X"B1",X"47",
		X"13",X"57",X"20",X"60",X"B0",X"20",X"50",X"B0",X"41",X"1F",X"51",X"74",X"58",X"38",X"94",X"FE",
		X"35",X"94",X"DF",X"42",X"1F",X"52",X"44",X"18",X"1F",X"C1",X"51",X"44",X"36",X"94",X"C4",X"44",
		X"18",X"1F",X"C2",X"52",X"70",X"B0",X"1C",X"F8",X"88",X"88",X"88",X"F8",X"20",X"20",X"20",X"20",
		X"20",X"F8",X"08",X"F8",X"80",X"F8",X"F8",X"08",X"F8",X"08",X"F8",X"88",X"88",X"F8",X"08",X"08",
		X"F8",X"80",X"F8",X"08",X"F8",X"F8",X"80",X"F8",X"88",X"F8",X"F8",X"08",X"10",X"10",X"10",X"F8",
		X"88",X"F8",X"88",X"F8",X"F8",X"88",X"F8",X"08",X"F8",X"F8",X"80",X"98",X"88",X"F8",X"F8",X"08",
		X"38",X"00",X"20",X"F8",X"20",X"20",X"20",X"20",X"00",X"00",X"00",X"00",X"00",X"F8",X"A8",X"A8",
		X"A8",X"A8",X"88",X"50",X"20",X"50",X"88",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"20",X"00",X"20",
		X"00",X"00",X"00",X"F8",X"00",X"00",X"50",X"50",X"50",X"50",X"50",X"A0",X"A0",X"A0",X"A0",X"A0",
		X"C0",X"C0",X"00",X"00",X"00",X"08",X"08",X"08",X"08",X"08",X"20",X"20",X"20",X"20",X"20",X"10",
		X"10",X"20",X"40",X"40",X"08",X"10",X"20",X"40",X"80",X"00",X"18",X"20",X"C0",X"00",X"00",X"C0",
		X"20",X"18",X"00",X"80",X"40",X"20",X"10",X"08",X"40",X"40",X"20",X"10",X"10",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
