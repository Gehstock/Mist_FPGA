library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity bwidow_pgm_rom1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of bwidow_pgm_rom1 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"28",X"43",X"29",X"20",X"41",X"54",
		X"41",X"52",X"49",X"20",X"31",X"39",X"38",X"32",X"A9",X"55",X"85",X"00",X"A9",X"00",X"8D",X"0F",
		X"60",X"8D",X"0F",X"68",X"A9",X"07",X"8D",X"0F",X"60",X"8D",X"0F",X"68",X"D8",X"8D",X"80",X"88",
		X"A9",X"38",X"8D",X"00",X"88",X"A9",X"00",X"85",X"01",X"85",X"02",X"A0",X"03",X"A9",X"00",X"91",
		X"01",X"C8",X"D0",X"F9",X"E6",X"02",X"A5",X"02",X"49",X"08",X"D0",X"F1",X"20",X"4E",X"E7",X"A9",
		X"01",X"85",X"FE",X"85",X"FF",X"A9",X"80",X"85",X"EF",X"A2",X"1F",X"8A",X"BD",X"B5",X"A5",X"9D",
		X"00",X"01",X"CA",X"10",X"F6",X"A9",X"C8",X"8D",X"00",X"88",X"85",X"99",X"A9",X"0A",X"85",X"4E",
		X"A2",X"00",X"A9",X"01",X"85",X"1B",X"85",X"1D",X"A9",X"50",X"85",X"1C",X"85",X"1E",X"A9",X"00",
		X"9D",X"D7",X"03",X"A5",X"1D",X"9D",X"D5",X"03",X"A5",X"1E",X"9D",X"D6",X"03",X"18",X"F8",X"65",
		X"1C",X"85",X"1E",X"A5",X"1D",X"65",X"1B",X"85",X"1D",X"D8",X"E8",X"E8",X"E8",X"E0",X"4B",X"90",
		X"DD",X"8D",X"0B",X"68",X"AD",X"08",X"68",X"29",X"03",X"AA",X"BD",X"25",X"9C",X"29",X"FC",X"8D",
		X"2B",X"06",X"A9",X"01",X"8D",X"01",X"02",X"20",X"95",X"9F",X"8D",X"80",X"89",X"20",X"0E",X"BE",
		X"20",X"9C",X"9D",X"20",X"54",X"99",X"A9",X"F6",X"8D",X"D0",X"03",X"58",X"A9",X"00",X"8D",X"2D",
		X"01",X"20",X"A9",X"D6",X"AD",X"2E",X"01",X"D0",X"FB",X"A9",X"00",X"8D",X"2A",X"01",X"A9",X"AA",
		X"85",X"00",X"8D",X"80",X"89",X"24",X"EF",X"10",X"2A",X"AD",X"20",X"04",X"C9",X"05",X"F0",X"23",
		X"AD",X"22",X"04",X"D0",X"1E",X"20",X"DC",X"B7",X"AE",X"23",X"04",X"BD",X"80",X"91",X"D0",X"05",
		X"A2",X"00",X"4C",X"FB",X"90",X"8D",X"22",X"04",X"BD",X"81",X"91",X"8D",X"21",X"04",X"E8",X"E8",
		X"8E",X"23",X"04",X"AD",X"21",X"04",X"F0",X"4C",X"CD",X"20",X"04",X"D0",X"08",X"A9",X"00",X"8D",
		X"21",X"04",X"4C",X"64",X"91",X"20",X"29",X"9C",X"AD",X"21",X"04",X"8D",X"20",X"04",X"0A",X"AA",
		X"20",X"3B",X"91",X"A9",X"00",X"8D",X"21",X"04",X"4C",X"64",X"91",X"BD",X"43",X"91",X"48",X"BD",
		X"42",X"91",X"48",X"60",X"51",X"91",X"E0",X"91",X"95",X"92",X"AE",X"92",X"22",X"94",X"86",X"91",
		X"D6",X"9C",X"24",X"EF",X"10",X"0B",X"A9",X"00",X"85",X"79",X"8D",X"D3",X"03",X"85",X"F7",X"85",
		X"73",X"4C",X"9C",X"9D",X"AD",X"20",X"04",X"0A",X"AA",X"BD",X"71",X"91",X"48",X"BD",X"70",X"91",
		X"48",X"60",X"52",X"98",X"8F",X"92",X"EA",X"92",X"F0",X"92",X"25",X"96",X"D8",X"91",X"F2",X"9C",
		X"24",X"01",X"0A",X"02",X"0A",X"03",X"00",X"24",X"EF",X"30",X"41",X"AD",X"C8",X"04",X"F0",X"3C",
		X"20",X"AA",X"9C",X"A2",X"02",X"20",X"B7",X"DC",X"AD",X"C9",X"04",X"18",X"69",X"01",X"20",X"AF",
		X"D7",X"20",X"C9",X"D8",X"A9",X"00",X"A0",X"00",X"20",X"EF",X"D7",X"A9",X"B0",X"A2",X"50",X"20",
		X"1D",X"D8",X"A9",X"50",X"A2",X"B0",X"20",X"1D",X"D8",X"20",X"A2",X"D7",X"A9",X"03",X"8D",X"22",
		X"04",X"A9",X"00",X"8D",X"20",X"01",X"8D",X"40",X"88",X"85",X"81",X"60",X"68",X"68",X"A9",X"01",
		X"8D",X"21",X"04",X"8D",X"D4",X"03",X"4C",X"13",X"91",X"AD",X"22",X"04",X"F0",X"F0",X"4C",X"2C",
		X"96",X"A9",X"00",X"85",X"11",X"A9",X"20",X"85",X"12",X"20",X"C9",X"D8",X"A0",X"00",X"A9",X"01",
		X"20",X"12",X"D8",X"A9",X"B0",X"A2",X"18",X"20",X"1D",X"D8",X"A0",X"00",X"A9",X"00",X"20",X"12",
		X"D8",X"A9",X"00",X"A0",X"E4",X"20",X"EF",X"D7",X"A9",X"A2",X"AA",X"A9",X"2F",X"20",X"E3",X"D7",
		X"20",X"C9",X"D8",X"A0",X"00",X"A9",X"01",X"20",X"12",X"D8",X"A9",X"A4",X"A2",X"E0",X"20",X"1D",
		X"D8",X"A0",X"20",X"A9",X"00",X"20",X"12",X"D8",X"A9",X"00",X"A0",X"E4",X"20",X"EF",X"D7",X"A9",
		X"44",X"AA",X"A9",X"30",X"20",X"E3",X"D7",X"A0",X"00",X"A9",X"01",X"20",X"12",X"D8",X"20",X"C9",
		X"D8",X"A2",X"2A",X"20",X"B7",X"DC",X"AD",X"2E",X"06",X"29",X"03",X"AA",X"BD",X"88",X"92",X"AA",
		X"20",X"B7",X"DC",X"AD",X"45",X"04",X"F0",X"22",X"A2",X"30",X"20",X"B7",X"DC",X"AD",X"2F",X"06",
		X"4A",X"4A",X"4A",X"4A",X"4A",X"4A",X"18",X"69",X"02",X"20",X"AF",X"D7",X"A9",X"04",X"85",X"1E",
		X"A9",X"00",X"18",X"20",X"AF",X"D7",X"C6",X"1E",X"D0",X"F6",X"20",X"A6",X"D7",X"A9",X"00",X"85",
		X"81",X"8D",X"20",X"01",X"8D",X"40",X"88",X"60",X"26",X"28",X"22",X"24",X"02",X"03",X"00",X"01",
		X"20",X"9C",X"96",X"4C",X"2C",X"96",X"A9",X"00",X"85",X"11",X"A9",X"20",X"85",X"12",X"20",X"7F",
		X"CB",X"20",X"A6",X"D7",X"A9",X"00",X"8D",X"20",X"01",X"8D",X"40",X"88",X"85",X"81",X"60",X"A9",
		X"00",X"85",X"11",X"85",X"A5",X"A9",X"0F",X"85",X"A8",X"A9",X"20",X"85",X"12",X"20",X"7F",X"CB",
		X"A2",X"0A",X"20",X"B7",X"DC",X"A2",X"0C",X"20",X"B7",X"DC",X"A2",X"0E",X"20",X"B7",X"DC",X"20",
		X"A6",X"D7",X"A9",X"FF",X"85",X"72",X"A9",X"00",X"85",X"71",X"8D",X"20",X"01",X"8D",X"40",X"88",
		X"85",X"81",X"8D",X"01",X"03",X"A9",X"3C",X"8D",X"22",X"04",X"60",X"20",X"9C",X"96",X"4C",X"2C",
		X"96",X"AD",X"22",X"04",X"D0",X"03",X"4C",X"D1",X"93",X"A9",X"1E",X"8D",X"24",X"04",X"E6",X"6F",
		X"A5",X"72",X"10",X"12",X"AD",X"00",X"88",X"29",X"0F",X"49",X"0F",X"F0",X"03",X"4C",X"2C",X"96",
		X"85",X"A8",X"A9",X"01",X"85",X"72",X"A5",X"6F",X"29",X"03",X"D0",X"11",X"A0",X"00",X"AD",X"0A",
		X"60",X"29",X"03",X"AA",X"BD",X"F2",X"CD",X"91",X"A3",X"A0",X"14",X"91",X"A3",X"AD",X"00",X"80",
		X"29",X"0F",X"C9",X"0F",X"F0",X"36",X"A8",X"C6",X"71",X"10",X"31",X"A9",X"05",X"85",X"71",X"98",
		X"29",X"0C",X"C9",X"0C",X"F0",X"15",X"EE",X"01",X"03",X"29",X"08",X"D0",X"06",X"CE",X"01",X"03",
		X"CE",X"01",X"03",X"AD",X"01",X"03",X"29",X"03",X"8D",X"01",X"03",X"98",X"29",X"03",X"C9",X"03",
		X"F0",X"0A",X"E6",X"72",X"29",X"01",X"F0",X"04",X"C6",X"72",X"C6",X"72",X"A5",X"72",X"29",X"1F",
		X"85",X"72",X"F0",X"03",X"0A",X"69",X"14",X"AA",X"AC",X"01",X"03",X"B9",X"F2",X"CD",X"48",X"A5",
		X"A5",X"0A",X"0A",X"18",X"69",X"08",X"A8",X"68",X"91",X"A3",X"C8",X"C8",X"BD",X"C4",X"5D",X"91",
		X"A3",X"20",X"0C",X"94",X"B0",X"03",X"4C",X"2C",X"96",X"A5",X"72",X"C9",X"1F",X"D0",X"13",X"A5",
		X"A5",X"F0",X"F3",X"0A",X"0A",X"69",X"08",X"A8",X"AD",X"C4",X"5D",X"91",X"A3",X"C6",X"A5",X"4C",
		X"2C",X"96",X"A5",X"A5",X"18",X"65",X"A9",X"AA",X"AD",X"01",X"03",X"0A",X"0A",X"0A",X"0A",X"0A",
		X"0A",X"05",X"72",X"9D",X"10",X"03",X"E6",X"A5",X"A5",X"A5",X"C9",X"03",X"F0",X"03",X"4C",X"2C",
		X"96",X"A5",X"F6",X"C9",X"03",X"F0",X"03",X"20",X"8F",X"D6",X"A9",X"1E",X"8D",X"24",X"04",X"AD",
		X"C8",X"04",X"F0",X"0B",X"AD",X"C9",X"04",X"D0",X"06",X"8D",X"20",X"04",X"4C",X"EB",X"9B",X"A9",
		X"00",X"8D",X"22",X"04",X"8D",X"23",X"04",X"8D",X"2C",X"06",X"A9",X"80",X"8D",X"20",X"04",X"85",
		X"EF",X"A9",X"01",X"8D",X"21",X"04",X"20",X"DC",X"B7",X"4C",X"13",X"91",X"AD",X"00",X"88",X"29",
		X"0F",X"49",X"0F",X"F0",X"04",X"85",X"A8",X"18",X"60",X"A5",X"A8",X"F0",X"FA",X"A9",X"00",X"85",
		X"A8",X"38",X"60",X"A9",X"02",X"85",X"11",X"A9",X"20",X"85",X"12",X"E6",X"6F",X"A5",X"6F",X"4A",
		X"90",X"04",X"A9",X"24",X"85",X"12",X"20",X"C9",X"D8",X"A0",X"00",X"A9",X"01",X"20",X"12",X"D8",
		X"20",X"C9",X"D8",X"AD",X"2E",X"01",X"0D",X"2B",X"01",X"D0",X"44",X"A2",X"46",X"20",X"B7",X"DC",
		X"A2",X"00",X"AD",X"2C",X"06",X"8E",X"2C",X"06",X"29",X"20",X"F0",X"21",X"AD",X"00",X"88",X"49",
		X"0F",X"29",X"0F",X"F0",X"0D",X"AD",X"01",X"03",X"29",X"03",X"0A",X"AA",X"20",X"EE",X"95",X"4C",
		X"99",X"94",X"EE",X"01",X"03",X"AD",X"01",X"03",X"29",X"03",X"8D",X"01",X"03",X"AD",X"01",X"03",
		X"AA",X"BD",X"8B",X"94",X"AA",X"20",X"B7",X"DC",X"4C",X"99",X"94",X"48",X"4A",X"4C",X"4E",X"A2",
		X"50",X"20",X"B7",X"DC",X"A9",X"00",X"8D",X"2C",X"06",X"A2",X"44",X"20",X"B7",X"DC",X"A5",X"7A",
		X"85",X"65",X"A5",X"7B",X"85",X"66",X"A9",X"00",X"85",X"63",X"20",X"4B",X"96",X"20",X"82",X"96",
		X"AD",X"2E",X"06",X"29",X"03",X"AA",X"BD",X"88",X"92",X"AA",X"20",X"B7",X"DC",X"AD",X"45",X"04",
		X"F0",X"22",X"A2",X"30",X"20",X"B7",X"DC",X"AD",X"2F",X"06",X"4A",X"4A",X"4A",X"4A",X"4A",X"4A",
		X"18",X"69",X"02",X"20",X"AF",X"D7",X"A9",X"04",X"85",X"1E",X"A9",X"00",X"18",X"20",X"AF",X"D7",
		X"C6",X"1E",X"D0",X"F6",X"A2",X"36",X"20",X"B7",X"DC",X"AD",X"2F",X"06",X"29",X"0C",X"4A",X"4A",
		X"69",X"03",X"20",X"AF",X"D7",X"A2",X"3A",X"20",X"B7",X"DC",X"AD",X"2F",X"06",X"29",X"03",X"AA",
		X"BD",X"25",X"9C",X"20",X"A1",X"DC",X"48",X"4A",X"4A",X"4A",X"4A",X"20",X"AF",X"D7",X"68",X"29",
		X"0F",X"20",X"AF",X"D7",X"A2",X"52",X"20",X"B7",X"DC",X"AD",X"2E",X"06",X"29",X"E0",X"4A",X"4A",
		X"4A",X"4A",X"4A",X"20",X"AF",X"D7",X"A2",X"54",X"20",X"B7",X"DC",X"AD",X"2E",X"06",X"29",X"10",
		X"4A",X"4A",X"4A",X"4A",X"18",X"69",X"01",X"20",X"AF",X"D7",X"A2",X"56",X"20",X"B7",X"DC",X"AD",
		X"2E",X"06",X"4A",X"4A",X"29",X"03",X"18",X"69",X"01",X"C9",X"01",X"F0",X"03",X"18",X"69",X"02",
		X"20",X"AF",X"D7",X"A5",X"7A",X"05",X"7B",X"D0",X"03",X"4C",X"A5",X"95",X"A2",X"38",X"20",X"B7",
		X"DC",X"A5",X"7C",X"85",X"1B",X"A5",X"7D",X"85",X"1C",X"A5",X"7E",X"85",X"1D",X"A9",X"00",X"85",
		X"65",X"85",X"66",X"E6",X"65",X"D0",X"02",X"E6",X"66",X"A5",X"1B",X"38",X"E5",X"7A",X"85",X"1B",
		X"A5",X"1C",X"E5",X"7B",X"85",X"1C",X"A5",X"1D",X"E9",X"00",X"85",X"1D",X"10",X"E5",X"A9",X"00",
		X"85",X"63",X"20",X"4B",X"96",X"A0",X"00",X"A5",X"1C",X"20",X"3F",X"CC",X"A5",X"1B",X"20",X"43",
		X"CC",X"88",X"20",X"05",X"D8",X"AD",X"2F",X"06",X"29",X"30",X"4A",X"4A",X"4A",X"4A",X"AA",X"BD",
		X"22",X"96",X"AA",X"20",X"B7",X"DC",X"AD",X"00",X"78",X"29",X"40",X"F0",X"F9",X"20",X"29",X"9C",
		X"A9",X"02",X"85",X"1B",X"A9",X"20",X"85",X"1C",X"A5",X"6F",X"4A",X"90",X"04",X"A9",X"24",X"85",
		X"1C",X"20",X"A6",X"D7",X"A9",X"00",X"85",X"11",X"A9",X"20",X"85",X"12",X"A6",X"1B",X"A5",X"1C",
		X"20",X"CF",X"D7",X"A9",X"00",X"8D",X"40",X"88",X"8D",X"20",X"01",X"85",X"81",X"60",X"BD",X"F8",
		X"95",X"48",X"BD",X"F7",X"95",X"48",X"60",X"75",X"E7",X"FE",X"95",X"08",X"96",X"1A",X"96",X"20",
		X"F6",X"CD",X"20",X"88",X"9F",X"20",X"8F",X"D6",X"60",X"78",X"A9",X"00",X"85",X"7C",X"85",X"7D",
		X"85",X"7E",X"85",X"7A",X"85",X"7B",X"58",X"20",X"93",X"D6",X"60",X"20",X"FF",X"95",X"20",X"09",
		X"96",X"60",X"3E",X"40",X"42",X"3C",X"20",X"9C",X"96",X"20",X"23",X"94",X"AD",X"20",X"01",X"D0",
		X"11",X"AD",X"00",X"78",X"29",X"40",X"D0",X"0D",X"A9",X"00",X"85",X"00",X"A9",X"AA",X"C5",X"00",
		X"D0",X"FA",X"4C",X"E2",X"90",X"8D",X"40",X"88",X"4C",X"E2",X"90",X"A9",X"00",X"85",X"1B",X"85",
		X"1C",X"85",X"1D",X"85",X"1E",X"A0",X"18",X"18",X"F8",X"A5",X"1B",X"65",X"1B",X"85",X"1B",X"A5",
		X"1C",X"65",X"1C",X"85",X"1C",X"A5",X"1D",X"65",X"1D",X"85",X"1D",X"A5",X"1E",X"65",X"1E",X"85",
		X"1E",X"D8",X"06",X"65",X"26",X"66",X"26",X"63",X"A5",X"1B",X"69",X"00",X"85",X"1B",X"88",X"D0",
		X"D6",X"60",X"A0",X"00",X"A5",X"1E",X"20",X"3F",X"CC",X"A5",X"1D",X"20",X"43",X"CC",X"A5",X"1C",
		X"20",X"43",X"CC",X"A5",X"1B",X"20",X"43",X"CC",X"88",X"4C",X"05",X"D8",X"24",X"EF",X"10",X"3F",
		X"AD",X"00",X"78",X"29",X"10",X"F0",X"20",X"AD",X"20",X"04",X"C9",X"05",X"D0",X"31",X"A9",X"00",
		X"8D",X"23",X"04",X"8D",X"22",X"04",X"8D",X"80",X"88",X"8D",X"20",X"01",X"85",X"8D",X"85",X"95",
		X"A9",X"01",X"8D",X"21",X"04",X"18",X"60",X"A9",X"05",X"8D",X"21",X"04",X"8D",X"0B",X"68",X"AD",
		X"08",X"68",X"29",X"03",X"AA",X"BD",X"25",X"9C",X"29",X"FC",X"8D",X"2B",X"06",X"18",X"60",X"AD",
		X"2F",X"06",X"29",X"C0",X"4A",X"4A",X"4A",X"4A",X"4A",X"4A",X"18",X"69",X"02",X"C9",X"05",X"D0",
		X"02",X"A9",X"00",X"8D",X"45",X"04",X"AD",X"2E",X"06",X"29",X"03",X"AA",X"4D",X"2E",X"06",X"1D",
		X"8C",X"92",X"85",X"8C",X"29",X"03",X"D0",X"0E",X"78",X"A5",X"99",X"29",X"F7",X"85",X"99",X"8D",
		X"00",X"88",X"58",X"4C",X"21",X"97",X"78",X"A5",X"99",X"09",X"08",X"85",X"99",X"8D",X"00",X"88",
		X"58",X"A5",X"8C",X"29",X"03",X"D0",X"05",X"A9",X"02",X"4C",X"3B",X"97",X"A5",X"8D",X"D0",X"0B",
		X"A5",X"99",X"09",X"F0",X"85",X"99",X"8D",X"00",X"88",X"18",X"60",X"24",X"EF",X"30",X"02",X"18",
		X"60",X"A2",X"EF",X"C9",X"02",X"90",X"02",X"A2",X"CF",X"78",X"A5",X"99",X"09",X"30",X"85",X"99",
		X"AD",X"D0",X"03",X"29",X"20",X"F0",X"05",X"8A",X"25",X"99",X"85",X"99",X"A5",X"99",X"8D",X"00",
		X"88",X"58",X"A5",X"8C",X"29",X"03",X"F0",X"06",X"A5",X"8D",X"C9",X"02",X"90",X"30",X"AD",X"2C",
		X"06",X"D0",X"07",X"18",X"A9",X"00",X"8D",X"2C",X"06",X"60",X"78",X"A2",X"00",X"8E",X"2C",X"06",
		X"58",X"29",X"20",X"D0",X"20",X"A9",X"01",X"8D",X"CA",X"04",X"8D",X"C8",X"04",X"A5",X"8C",X"29",
		X"03",X"F0",X"02",X"C6",X"8D",X"E6",X"7A",X"D0",X"02",X"E6",X"7B",X"4C",X"AF",X"97",X"AD",X"2C",
		X"06",X"29",X"20",X"F0",X"CE",X"78",X"A9",X"00",X"8D",X"2C",X"06",X"58",X"8D",X"C8",X"04",X"A9",
		X"00",X"8D",X"C9",X"04",X"A5",X"8C",X"29",X"03",X"F0",X"02",X"C6",X"8D",X"E6",X"7A",X"D0",X"02",
		X"E6",X"7B",X"68",X"68",X"A9",X"00",X"85",X"F5",X"85",X"F4",X"AD",X"2F",X"06",X"29",X"30",X"4A",
		X"4A",X"4A",X"4A",X"85",X"F6",X"C9",X"03",X"D0",X"0A",X"A5",X"8C",X"29",X"E3",X"F0",X"04",X"A9",
		X"02",X"85",X"F6",X"A9",X"00",X"8D",X"41",X"04",X"8D",X"42",X"04",X"8D",X"43",X"04",X"A9",X"07",
		X"8D",X"21",X"04",X"AD",X"2F",X"06",X"29",X"0C",X"4A",X"4A",X"69",X"02",X"8D",X"40",X"04",X"20",
		X"DC",X"B7",X"A9",X"04",X"8D",X"58",X"04",X"A9",X"FF",X"85",X"9A",X"A9",X"00",X"8D",X"47",X"04",
		X"85",X"EF",X"8D",X"2C",X"06",X"A9",X"03",X"8D",X"5C",X"04",X"20",X"0E",X"BE",X"A2",X"0F",X"A9",
		X"00",X"9D",X"48",X"04",X"CA",X"10",X"FA",X"A2",X"10",X"A9",X"03",X"9D",X"00",X"02",X"E0",X"50",
		X"90",X"06",X"9D",X"7B",X"04",X"9D",X"2B",X"05",X"8A",X"18",X"69",X"10",X"AA",X"D0",X"EA",X"A0",
		X"35",X"A2",X"00",X"BD",X"29",X"04",X"9D",X"93",X"04",X"9D",X"5E",X"04",X"E8",X"88",X"D0",X"F3",
		X"4C",X"13",X"91",X"AD",X"D4",X"03",X"D0",X"22",X"A5",X"EF",X"10",X"1B",X"20",X"9C",X"96",X"AD",
		X"00",X"02",X"C9",X"03",X"D0",X"11",X"A9",X"FF",X"85",X"9A",X"A9",X"00",X"8D",X"5D",X"04",X"A9",
		X"04",X"8D",X"58",X"04",X"4C",X"7F",X"98",X"4C",X"A2",X"98",X"A9",X"00",X"8D",X"D4",X"03",X"A9",
		X"00",X"8D",X"00",X"21",X"8D",X"06",X"21",X"A9",X"02",X"8D",X"00",X"02",X"A9",X"00",X"8D",X"28",
		X"04",X"A9",X"08",X"05",X"5E",X"85",X"5E",X"20",X"C7",X"A0",X"A9",X"00",X"8D",X"00",X"02",X"4C",
		X"63",X"99",X"A9",X"00",X"85",X"00",X"A5",X"00",X"C9",X"AA",X"D0",X"FA",X"20",X"F1",X"B1",X"C6",
		X"FF",X"D0",X"EF",X"A5",X"FE",X"85",X"FF",X"A5",X"FC",X"F0",X"0F",X"AD",X"00",X"88",X"29",X"40",
		X"A8",X"45",X"FD",X"84",X"FD",X"F0",X"DB",X"98",X"F0",X"D8",X"E6",X"6F",X"A5",X"6F",X"29",X"01",
		X"D0",X"03",X"20",X"72",X"D9",X"20",X"D2",X"A3",X"20",X"C7",X"A0",X"8D",X"80",X"89",X"20",X"F5",
		X"A5",X"8D",X"80",X"89",X"A9",X"00",X"85",X"21",X"85",X"40",X"A0",X"40",X"20",X"CF",X"CE",X"20",
		X"30",X"CF",X"A5",X"6C",X"F0",X"26",X"A2",X"10",X"A9",X"03",X"9D",X"00",X"02",X"8A",X"18",X"69",
		X"10",X"AA",X"C9",X"50",X"90",X"F2",X"A9",X"00",X"85",X"79",X"AD",X"00",X"02",X"C9",X"03",X"D0",
		X"03",X"4C",X"A6",X"99",X"A9",X"02",X"8D",X"00",X"02",X"8D",X"01",X"03",X"A9",X"00",X"85",X"40",
		X"A5",X"40",X"18",X"69",X"10",X"C9",X"50",X"D0",X"03",X"4C",X"39",X"99",X"85",X"40",X"A0",X"50",
		X"20",X"B3",X"CE",X"20",X"30",X"CF",X"4C",X"20",X"99",X"A9",X"50",X"85",X"40",X"18",X"69",X"10",
		X"90",X"03",X"4C",X"E2",X"90",X"A8",X"20",X"B3",X"CE",X"20",X"30",X"CF",X"A5",X"6E",X"18",X"69",
		X"10",X"4C",X"3B",X"99",X"A0",X"10",X"A9",X"03",X"99",X"00",X"02",X"98",X"18",X"69",X"10",X"A8",
		X"D0",X"F4",X"60",X"A9",X"00",X"85",X"73",X"24",X"EF",X"30",X"02",X"E6",X"73",X"A9",X"A2",X"8D",
		X"02",X"01",X"8D",X"03",X"01",X"A9",X"00",X"8D",X"06",X"02",X"85",X"6C",X"8D",X"0B",X"02",X"8D",
		X"09",X"02",X"A9",X"64",X"8D",X"0C",X"02",X"AD",X"C8",X"04",X"F0",X"0D",X"AD",X"C9",X"04",X"F0",
		X"08",X"A9",X"64",X"8D",X"0A",X"02",X"4C",X"9E",X"99",X"A9",X"CC",X"8D",X"0A",X"02",X"20",X"3B",
		X"9C",X"4C",X"2C",X"96",X"BF",X"00",X"A9",X"00",X"8D",X"00",X"02",X"8D",X"03",X"03",X"8D",X"D3",
		X"03",X"8D",X"06",X"02",X"8D",X"3A",X"04",X"8D",X"3B",X"04",X"8D",X"04",X"03",X"AD",X"28",X"04",
		X"F0",X"0F",X"A2",X"0F",X"A9",X"00",X"9D",X"48",X"04",X"CA",X"10",X"F8",X"A9",X"00",X"8D",X"28",
		X"04",X"AD",X"01",X"02",X"29",X"EF",X"8D",X"01",X"02",X"24",X"EF",X"10",X"03",X"4C",X"63",X"99",
		X"CE",X"40",X"04",X"10",X"6E",X"A9",X"01",X"8D",X"20",X"01",X"8D",X"80",X"88",X"20",X"AA",X"9C",
		X"A9",X"FE",X"18",X"65",X"11",X"85",X"11",X"A5",X"12",X"69",X"FF",X"85",X"12",X"A2",X"00",X"20",
		X"B7",X"DC",X"AD",X"C8",X"04",X"F0",X"0E",X"A2",X"02",X"20",X"B7",X"DC",X"AD",X"C9",X"04",X"18",
		X"69",X"01",X"20",X"AF",X"D7",X"A2",X"1A",X"20",X"B7",X"DC",X"AD",X"5D",X"04",X"18",X"69",X"01",
		X"20",X"A1",X"DC",X"48",X"4A",X"4A",X"4A",X"4A",X"38",X"20",X"AF",X"D7",X"68",X"29",X"0F",X"20",
		X"AF",X"D7",X"20",X"A2",X"D7",X"A9",X"03",X"8D",X"22",X"04",X"20",X"C1",X"91",X"AD",X"00",X"78",
		X"29",X"40",X"D0",X"0A",X"A9",X"00",X"85",X"00",X"A9",X"AA",X"C5",X"00",X"D0",X"FA",X"AD",X"22",
		X"04",X"D0",X"E7",X"A9",X"29",X"85",X"4C",X"A9",X"04",X"85",X"4D",X"AD",X"C8",X"04",X"F0",X"05",
		X"AD",X"C9",X"04",X"D0",X"18",X"A9",X"5E",X"85",X"49",X"A9",X"04",X"85",X"4A",X"A2",X"00",X"BD",
		X"50",X"02",X"9D",X"CB",X"04",X"E8",X"E0",X"B0",X"D0",X"F5",X"4C",X"92",X"9A",X"A9",X"93",X"85",
		X"49",X"A9",X"04",X"85",X"4A",X"A2",X"00",X"BD",X"50",X"02",X"9D",X"7B",X"05",X"E8",X"E0",X"B0",
		X"D0",X"F5",X"A2",X"35",X"20",X"5C",X"A0",X"AD",X"C8",X"04",X"D0",X"03",X"4C",X"22",X"9B",X"AD",
		X"C9",X"04",X"D0",X"10",X"AD",X"AA",X"04",X"30",X"79",X"A9",X"93",X"85",X"4C",X"A9",X"04",X"85",
		X"4D",X"4C",X"C1",X"9A",X"AD",X"75",X"04",X"30",X"69",X"A9",X"5E",X"85",X"4C",X"A9",X"04",X"85",
		X"4D",X"A2",X"35",X"A9",X"29",X"85",X"49",X"A9",X"04",X"85",X"4A",X"20",X"5C",X"A0",X"A9",X"FF",
		X"4D",X"C9",X"04",X"29",X"01",X"8D",X"C9",X"04",X"A2",X"00",X"AD",X"C8",X"04",X"F0",X"05",X"AD",
		X"C9",X"04",X"D0",X"0E",X"BD",X"CB",X"04",X"9D",X"50",X"02",X"E8",X"E0",X"B0",X"D0",X"F5",X"4C",
		X"FD",X"9A",X"BD",X"7B",X"05",X"9D",X"50",X"02",X"E8",X"E0",X"B0",X"D0",X"F5",X"AD",X"C9",X"04",
		X"F0",X"20",X"AD",X"CA",X"04",X"F0",X"1B",X"AD",X"C3",X"04",X"8D",X"59",X"04",X"8D",X"3E",X"04",
		X"A9",X"00",X"8D",X"CA",X"04",X"A9",X"07",X"8D",X"21",X"04",X"A9",X"1E",X"8D",X"22",X"04",X"4C",
		X"13",X"91",X"AD",X"C8",X"04",X"D0",X"08",X"AD",X"75",X"04",X"10",X"10",X"4C",X"62",X"9B",X"AD",
		X"75",X"04",X"10",X"08",X"AD",X"AA",X"04",X"10",X"03",X"4C",X"62",X"9B",X"A2",X"10",X"BD",X"01",
		X"02",X"29",X"07",X"C9",X"03",X"D0",X"07",X"BD",X"00",X"02",X"29",X"02",X"F0",X"05",X"A9",X"03",
		X"9D",X"00",X"02",X"8A",X"18",X"69",X"10",X"AA",X"D0",X"E4",X"A9",X"06",X"8D",X"21",X"04",X"4C",
		X"13",X"91",X"A5",X"F6",X"C9",X"03",X"F0",X"03",X"20",X"93",X"D6",X"A9",X"00",X"8D",X"C9",X"04",
		X"AD",X"76",X"04",X"8D",X"41",X"04",X"AD",X"77",X"04",X"8D",X"42",X"04",X"AD",X"78",X"04",X"8D",
		X"43",X"04",X"AD",X"92",X"04",X"8D",X"5D",X"04",X"AD",X"92",X"04",X"8D",X"59",X"04",X"AE",X"C8",
		X"04",X"F0",X"0B",X"AD",X"59",X"04",X"CD",X"C7",X"04",X"B0",X"03",X"AD",X"C7",X"04",X"CD",X"2B",
		X"06",X"90",X"05",X"F0",X"03",X"4C",X"BD",X"9B",X"A9",X"0D",X"85",X"19",X"AD",X"2F",X"06",X"29",
		X"03",X"AA",X"AD",X"2B",X"06",X"DD",X"25",X"9C",X"90",X"08",X"38",X"E9",X"04",X"29",X"FC",X"8D",
		X"2B",X"06",X"8D",X"59",X"04",X"8D",X"8E",X"04",X"8D",X"C3",X"04",X"20",X"90",X"CC",X"A9",X"00",
		X"8D",X"2C",X"06",X"A9",X"80",X"85",X"EF",X"AD",X"21",X"04",X"C9",X"04",X"D0",X"03",X"4C",X"13",
		X"91",X"AD",X"C8",X"04",X"F0",X"25",X"AD",X"C9",X"04",X"D0",X"20",X"A9",X"01",X"8D",X"C9",X"04",
		X"AD",X"AB",X"04",X"8D",X"41",X"04",X"AD",X"AC",X"04",X"8D",X"42",X"04",X"AD",X"AD",X"04",X"8D",
		X"43",X"04",X"AD",X"C7",X"04",X"8D",X"5D",X"04",X"4C",X"CB",X"9B",X"A9",X"1E",X"8D",X"24",X"04",
		X"A9",X"00",X"8D",X"20",X"04",X"8D",X"22",X"04",X"8D",X"23",X"04",X"8D",X"2C",X"06",X"A9",X"80",
		X"85",X"EF",X"4C",X"E2",X"90",X"0D",X"15",X"25",X"35",X"78",X"A9",X"01",X"8D",X"20",X"01",X"8D",
		X"80",X"88",X"AD",X"00",X"78",X"29",X"40",X"F0",X"F9",X"58",X"60",X"24",X"EF",X"30",X"6A",X"AD",
		X"C8",X"04",X"F0",X"30",X"A9",X"E4",X"A0",X"00",X"91",X"61",X"A9",X"00",X"A0",X"06",X"AE",X"AA",
		X"04",X"30",X"02",X"A9",X"E7",X"91",X"61",X"AD",X"C9",X"04",X"D0",X"09",X"AD",X"AA",X"04",X"18",
		X"69",X"02",X"4C",X"6B",X"9C",X"AD",X"AA",X"04",X"18",X"69",X"01",X"0A",X"AA",X"BD",X"C4",X"5D",
		X"A0",X"08",X"91",X"61",X"A9",X"E4",X"A0",X"00",X"91",X"5F",X"A0",X"06",X"A9",X"00",X"AE",X"75",
		X"04",X"30",X"02",X"A9",X"E7",X"91",X"5F",X"AD",X"C8",X"04",X"F0",X"0E",X"AD",X"C9",X"04",X"F0",
		X"09",X"AD",X"75",X"04",X"18",X"69",X"02",X"4C",X"A0",X"9C",X"AD",X"75",X"04",X"18",X"69",X"01",
		X"0A",X"AA",X"BD",X"C4",X"5D",X"A0",X"08",X"91",X"5F",X"60",X"A9",X"00",X"85",X"11",X"A9",X"20",
		X"85",X"12",X"20",X"C9",X"D8",X"A9",X"01",X"20",X"10",X"D8",X"A9",X"20",X"18",X"69",X"04",X"A2",
		X"00",X"20",X"E3",X"D7",X"20",X"A6",X"D7",X"A9",X"00",X"85",X"AA",X"85",X"11",X"A9",X"20",X"18",
		X"69",X"04",X"85",X"AB",X"85",X"12",X"60",X"AD",X"2B",X"06",X"8D",X"59",X"04",X"A9",X"0F",X"8D",
		X"22",X"04",X"20",X"AA",X"9C",X"A9",X"00",X"8D",X"5D",X"04",X"8D",X"2C",X"06",X"20",X"70",X"DA",
		X"4C",X"C1",X"91",X"A5",X"F6",X"C9",X"03",X"D0",X"15",X"A9",X"45",X"8D",X"22",X"04",X"AD",X"5D",
		X"04",X"C9",X"5D",X"B0",X"03",X"18",X"69",X"04",X"8D",X"2B",X"06",X"8D",X"59",X"04",X"E6",X"6F",
		X"A5",X"6F",X"29",X"07",X"F0",X"03",X"4C",X"69",X"9D",X"AD",X"00",X"88",X"49",X"0F",X"29",X"0F",
		X"F0",X"0A",X"A8",X"29",X"08",X"D0",X"50",X"98",X"29",X"04",X"D0",X"5C",X"AD",X"00",X"80",X"49",
		X"0F",X"29",X"0F",X"F0",X"34",X"A9",X"00",X"8D",X"2C",X"06",X"8D",X"2D",X"06",X"AD",X"00",X"88",
		X"49",X"FF",X"29",X"60",X"F0",X"23",X"A9",X"00",X"8D",X"2C",X"06",X"8D",X"5A",X"04",X"CE",X"5D",
		X"04",X"30",X"05",X"A9",X"02",X"8D",X"5A",X"04",X"AD",X"5D",X"04",X"8D",X"59",X"04",X"A9",X"01",
		X"8D",X"21",X"04",X"8D",X"D4",X"03",X"4C",X"13",X"91",X"20",X"AA",X"9C",X"20",X"70",X"DA",X"AD",
		X"22",X"04",X"F0",X"D2",X"4C",X"2C",X"96",X"AD",X"5D",X"04",X"F0",X"B0",X"38",X"E9",X"04",X"8D",
		X"5D",X"04",X"20",X"32",X"BD",X"4C",X"2C",X"9D",X"AD",X"5D",X"04",X"CD",X"59",X"04",X"B0",X"9C",
		X"18",X"69",X"04",X"8D",X"5D",X"04",X"20",X"32",X"BD",X"4C",X"2C",X"9D",X"A9",X"00",X"85",X"11",
		X"A9",X"20",X"85",X"12",X"20",X"C9",X"D8",X"A9",X"01",X"20",X"10",X"D8",X"A5",X"11",X"85",X"53",
		X"A5",X"12",X"85",X"54",X"A9",X"E4",X"A2",X"00",X"20",X"5B",X"D8",X"A9",X"80",X"85",X"08",X"A9",
		X"FE",X"85",X"09",X"A9",X"80",X"85",X"0A",X"A9",X"01",X"85",X"0B",X"20",X"E2",X"D8",X"20",X"A2",
		X"D8",X"A9",X"08",X"A2",X"04",X"20",X"1D",X"D8",X"A5",X"11",X"85",X"5F",X"A5",X"12",X"85",X"60",
		X"20",X"2F",X"A0",X"A5",X"11",X"85",X"55",X"A5",X"12",X"85",X"56",X"A9",X"E4",X"A2",X"00",X"20",
		X"5B",X"D8",X"A9",X"E0",X"85",X"08",X"A9",X"00",X"85",X"09",X"A9",X"80",X"85",X"0A",X"A9",X"01",
		X"85",X"0B",X"20",X"E2",X"D8",X"20",X"A2",X"D8",X"A9",X"08",X"A2",X"04",X"20",X"1D",X"D8",X"A5",
		X"11",X"85",X"61",X"A5",X"12",X"85",X"62",X"20",X"2F",X"A0",X"8D",X"80",X"89",X"20",X"68",X"9E",
		X"8D",X"80",X"89",X"20",X"A2",X"9E",X"A9",X"20",X"18",X"69",X"04",X"A2",X"00",X"20",X"E3",X"D7",
		X"20",X"A6",X"D7",X"A9",X"00",X"85",X"11",X"85",X"AA",X"A9",X"20",X"18",X"69",X"04",X"85",X"12",
		X"85",X"AB",X"20",X"A2",X"D7",X"A2",X"40",X"A0",X"0C",X"A5",X"F6",X"C9",X"03",X"F0",X"06",X"A9",
		X"0D",X"38",X"E5",X"F6",X"A8",X"98",X"9D",X"05",X"02",X"A9",X"04",X"9D",X"01",X"02",X"8A",X"38",
		X"E9",X"10",X"AA",X"D0",X"F0",X"4C",X"C1",X"91",X"20",X"C9",X"D8",X"A9",X"01",X"20",X"10",X"D8",
		X"A9",X"00",X"AA",X"A9",X"25",X"20",X"E3",X"D7",X"A5",X"11",X"85",X"13",X"A5",X"12",X"85",X"14",
		X"A9",X"25",X"85",X"12",X"A9",X"00",X"85",X"11",X"A9",X"40",X"85",X"0C",X"A9",X"A1",X"A2",X"00",
		X"20",X"5B",X"D8",X"20",X"76",X"BE",X"20",X"A2",X"D7",X"A5",X"13",X"85",X"11",X"A5",X"14",X"85",
		X"12",X"60",X"A2",X"00",X"A9",X"22",X"20",X"CF",X"D7",X"A5",X"11",X"48",X"A5",X"12",X"48",X"20",
		X"C9",X"D8",X"A2",X"00",X"A9",X"20",X"18",X"69",X"04",X"20",X"E3",X"D7",X"20",X"A6",X"D7",X"A2",
		X"00",X"A9",X"00",X"9D",X"00",X"22",X"9D",X"01",X"22",X"9D",X"02",X"22",X"9D",X"03",X"22",X"8A",
		X"09",X"80",X"9D",X"04",X"22",X"A9",X"A0",X"9D",X"05",X"22",X"A9",X"40",X"9D",X"06",X"22",X"A9",
		X"80",X"9D",X"07",X"22",X"8A",X"18",X"69",X"08",X"AA",X"C9",X"80",X"D0",X"D4",X"68",X"85",X"4D",
		X"68",X"85",X"4C",X"46",X"4D",X"66",X"4C",X"A5",X"4C",X"8D",X"7E",X"22",X"A5",X"4D",X"29",X"0F",
		X"09",X"E0",X"8D",X"7F",X"22",X"A2",X"00",X"A9",X"00",X"9D",X"00",X"21",X"A9",X"60",X"9D",X"01",
		X"21",X"A9",X"00",X"9D",X"02",X"21",X"A9",X"71",X"9D",X"03",X"21",X"A9",X"00",X"9D",X"04",X"21",
		X"A9",X"B4",X"9D",X"05",X"21",X"A9",X"00",X"9D",X"06",X"21",X"A9",X"60",X"9D",X"07",X"21",X"A9",
		X"00",X"9D",X"08",X"21",X"A9",X"AF",X"9D",X"09",X"21",X"A9",X"00",X"9D",X"0A",X"21",X"A9",X"71",
		X"9D",X"0B",X"21",X"A9",X"00",X"9D",X"0C",X"21",X"A9",X"60",X"9D",X"0D",X"21",X"A9",X"00",X"9D",
		X"0E",X"21",X"A9",X"C0",X"9D",X"0F",X"21",X"8A",X"18",X"69",X"10",X"AA",X"90",X"A9",X"A9",X"00",
		X"85",X"11",X"A9",X"20",X"18",X"69",X"03",X"85",X"12",X"A0",X"00",X"B9",X"69",X"D8",X"91",X"11",
		X"C8",X"C0",X"10",X"D0",X"F6",X"A5",X"11",X"18",X"69",X"10",X"85",X"11",X"90",X"EB",X"A9",X"00",
		X"85",X"73",X"A9",X"03",X"8D",X"00",X"02",X"60",X"A2",X"00",X"BD",X"A3",X"9F",X"9D",X"10",X"03",
		X"E8",X"E0",X"15",X"D0",X"F5",X"A2",X"00",X"BD",X"B8",X"9F",X"9D",X"25",X"03",X"E8",X"E0",X"77",
		X"D0",X"F5",X"60",X"C2",X"D7",X"CD",X"05",X"43",X"21",X"14",X"12",X"47",X"82",X"04",X"32",X"10",
		X"11",X"10",X"04",X"11",X"03",X"21",X"00",X"09",X"DB",X"1B",X"5B",X"01",X"08",X"01",X"11",X"C2",
		X"04",X"4D",X"01",X"01",X"01",X"11",X"D2",X"05",X"4F",X"01",X"01",X"01",X"11",X"D5",X"0E",X"52",
		X"01",X"01",X"01",X"11",X"C3",X"0E",X"47",X"01",X"01",X"01",X"11",X"C5",X"09",X"41",X"01",X"01",
		X"01",X"11",X"DB",X"13",X"4E",X"01",X"01",X"01",X"11",X"C2",X"9B",X"17",X"01",X"01",X"01",X"11",
		X"CC",X"9B",X"09",X"01",X"01",X"01",X"11",X"C1",X"9B",X"04",X"01",X"01",X"01",X"11",X"C3",X"9B");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
