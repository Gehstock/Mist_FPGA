library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity UNIWARS_1H is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of UNIWARS_1H is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",X"00",X"02",X"02",X"FE",X"FE",X"42",X"02",X"00",X"00",
		X"62",X"F2",X"BA",X"9A",X"9E",X"CE",X"46",X"00",X"8C",X"DE",X"F2",X"B2",X"92",X"86",X"04",X"00",
		X"08",X"FE",X"FE",X"C8",X"68",X"38",X"18",X"00",X"1C",X"BE",X"A2",X"A2",X"A2",X"E6",X"E4",X"00",
		X"0C",X"9E",X"92",X"92",X"D2",X"7E",X"3C",X"00",X"C0",X"E0",X"B0",X"9E",X"8E",X"C0",X"C0",X"00",
		X"0C",X"6E",X"9A",X"9A",X"B2",X"F2",X"6C",X"00",X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",X"00",
		X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",
		X"44",X"C6",X"82",X"82",X"C6",X"7C",X"38",X"00",X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",
		X"82",X"92",X"92",X"92",X"FE",X"FE",X"00",X"00",X"80",X"90",X"90",X"90",X"90",X"FE",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",
		X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",X"44",X"C6",X"82",X"82",X"C6",X"7C",X"38",X"00",
		X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",X"82",X"92",X"92",X"92",X"FE",X"FE",X"00",X"00",
		X"80",X"90",X"90",X"90",X"90",X"FE",X"FE",X"00",X"9E",X"9E",X"92",X"82",X"C6",X"7C",X"38",X"00",
		X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",X"82",X"82",X"FE",X"FE",X"82",X"82",X"00",X"00",
		X"FC",X"FE",X"02",X"02",X"02",X"06",X"04",X"00",X"82",X"C6",X"6E",X"3C",X"18",X"FE",X"FE",X"00",
		X"02",X"02",X"02",X"02",X"FE",X"FE",X"00",X"00",X"FE",X"FE",X"70",X"38",X"70",X"FE",X"FE",X"00",
		X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",X"00",
		X"70",X"F8",X"88",X"88",X"88",X"FE",X"FE",X"00",X"7A",X"FC",X"8E",X"8A",X"82",X"FE",X"7C",X"00",
		X"72",X"F6",X"9E",X"8C",X"88",X"FE",X"FE",X"00",X"0C",X"5E",X"D2",X"92",X"92",X"F6",X"64",X"00",
		X"80",X"80",X"FE",X"FE",X"80",X"80",X"00",X"00",X"FC",X"FE",X"02",X"02",X"02",X"FE",X"FC",X"00",
		X"F0",X"F8",X"1C",X"0E",X"1C",X"F8",X"F0",X"00",X"F8",X"FE",X"1C",X"38",X"1C",X"FE",X"F8",X"00",
		X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",X"C0",X"F0",X"1E",X"1E",X"F0",X"C0",X"00",X"00",
		X"C2",X"E2",X"F2",X"BA",X"9E",X"8E",X"86",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"10",X"18",X"1A",X"1E",X"1C",X"1C",X"18",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"F0",X"18",X"1C",X"1C",X"1E",X"1A",X"18",X"10",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",X"00",X"00",X"00",X"0E",X"1F",X"1C",X"0F",X"18",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",X"F0",X"18",X"0F",X"18",X"1F",X"0E",X"00",X"00",
		X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"80",X"A0",X"E0",X"C0",X"C0",X"80",
		X"0F",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"80",X"C0",X"C0",X"E0",X"A0",X"80",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"01",X"00",X"00",X"00",X"E0",X"F0",X"C0",X"F0",X"80",
		X"0F",X"01",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"80",X"F0",X"80",X"F0",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0E",X"0C",X"1E",X"1C",X"18",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"1E",X"1C",X"1E",X"0C",X"0E",X"04",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"40",X"E0",X"C0",X"E0",X"C0",X"80",
		X"0F",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"C0",X"E0",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"19",X"07",X"00",X"00",X"00",X"00",X"C0",X"E0",X"D0",X"C0",
		X"02",X"03",X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"C0",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"07",X"00",X"00",X"00",X"00",X"00",X"60",X"E0",X"F0",
		X"02",X"07",X"07",X"07",X"06",X"03",X"01",X"00",X"50",X"00",X"00",X"80",X"00",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"60",X"78",X"FC",
		X"01",X"07",X"07",X"07",X"03",X"03",X"01",X"00",X"34",X"00",X"80",X"00",X"00",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"F8",
		X"01",X"03",X"03",X"03",X"07",X"06",X"02",X"00",X"7C",X"34",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"1E",X"3C",X"38",X"28",X"00",X"00",X"00",X"F0",X"F8",X"30",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"FF",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FC",X"00",X"00",X"03",X"06",X"70",X"1E",X"00",X"60",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1E",X"70",X"06",X"03",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"0E",X"00",X"F8",X"00",X"0E",X"07",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"70",X"50",X"70",X"00",X"70",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"C3",X"A5",X"99",X"99",X"A5",X"C3",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"F0",X"7C",X"1F",
		X"00",X"00",X"01",X"04",X"06",X"02",X"05",X"0A",X"00",X"00",X"00",X"20",X"40",X"A8",X"50",X"20",
		X"04",X"06",X"06",X"05",X"01",X"00",X"00",X"00",X"E0",X"70",X"60",X"40",X"00",X"80",X"00",X"00",
		X"00",X"20",X"22",X"33",X"0B",X"0E",X"0F",X"0E",X"00",X"00",X"84",X"08",X"10",X"F6",X"E8",X"50",
		X"0A",X"07",X"02",X"04",X"08",X"10",X"10",X"20",X"60",X"E0",X"A0",X"90",X"48",X"44",X"20",X"00",
		X"00",X"00",X"3C",X"23",X"24",X"28",X"20",X"10",X"00",X"00",X"00",X"00",X"D0",X"60",X"30",X"10",
		X"08",X"0C",X"06",X"0B",X"00",X"00",X"00",X"00",X"10",X"30",X"60",X"D8",X"38",X"38",X"00",X"00",
		X"01",X"00",X"21",X"00",X"44",X"00",X"10",X"41",X"00",X"A0",X"04",X"40",X"00",X"10",X"00",X"85",
		X"A1",X"00",X"48",X"00",X"02",X"21",X"00",X"01",X"82",X"08",X"02",X"20",X"00",X"04",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"C0",
		X"00",X"01",X"0F",X"01",X"00",X"01",X"01",X"00",X"F0",X"E0",X"F0",X"E0",X"F0",X"C0",X"F0",X"E0",
		X"00",X"00",X"00",X"00",X"02",X"03",X"06",X"06",X"00",X"00",X"80",X"80",X"C0",X"E0",X"E0",X"E0",
		X"06",X"06",X"06",X"06",X"03",X"02",X"00",X"00",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"30",X"78",X"D8",X"B0",
		X"00",X"08",X"08",X"00",X"00",X"04",X"00",X"00",X"40",X"08",X"08",X"40",X"B0",X"D8",X"78",X"30",
		X"00",X"00",X"06",X"00",X"00",X"20",X"28",X"1C",X"30",X"08",X"C4",X"02",X"01",X"01",X"21",X"68",
		X"1C",X"88",X"80",X"80",X"40",X"26",X"10",X"0C",X"68",X"20",X"08",X"08",X"00",X"C0",X"00",X"00",
		X"00",X"00",X"03",X"04",X"01",X"12",X"22",X"00",X"00",X"00",X"00",X"30",X"08",X"00",X"00",X"C0",
		X"02",X"21",X"20",X"10",X"00",X"06",X"00",X"00",X"44",X"04",X"04",X"00",X"10",X"60",X"00",X"00",
		X"02",X"00",X"00",X"10",X"10",X"20",X"00",X"01",X"C0",X"00",X"10",X"08",X"00",X"00",X"84",X"40",
		X"20",X"22",X"00",X"00",X"10",X"00",X"00",X"06",X"80",X"04",X"04",X"00",X"00",X"10",X"00",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"13",X"33",X"FB",X"33",X"13",X"01",X"00",X"F8",X"81",X"BF",X"10",X"BF",X"81",X"F8",X"00",
		X"00",X"00",X"00",X"00",X"10",X"38",X"7C",X"F8",X"00",X"04",X"0E",X"07",X"0E",X"04",X"00",X"00",
		X"F3",X"F8",X"7C",X"38",X"10",X"00",X"00",X"00",X"C0",X"00",X"00",X"04",X"0E",X"07",X"0E",X"04",
		X"20",X"20",X"00",X"10",X"28",X"28",X"28",X"3E",X"2A",X"2A",X"2A",X"12",X"00",X"20",X"20",X"3E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"71",X"F3",X"E3",X"E3",X"E3",X"E3",X"E3",X"FC",X"FE",X"FF",X"FF",X"FF",X"9F",X"0F",X"07",
		X"E3",X"E3",X"E3",X"F7",X"FF",X"FF",X"7E",X"3C",X"07",X"07",X"07",X"07",X"0F",X"0F",X"0E",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"0E",X"0F",X"1F",X"5F",X"EF",X"F7",
		X"03",X"07",X"0B",X"0D",X"0E",X"07",X"03",X"01",X"FB",X"FD",X"FF",X"FF",X"FE",X"7E",X"BC",X"F8",
		X"00",X"00",X"34",X"7E",X"FD",X"DB",X"F7",X"EF",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",
		X"DF",X"BF",X"FF",X"FF",X"FF",X"FE",X"7D",X"1F",X"E0",X"E0",X"C0",X"B0",X"78",X"F8",X"F0",X"F0",
		X"03",X"07",X"07",X"06",X"01",X"03",X"01",X"00",X"F0",X"B1",X"7C",X"FE",X"FF",X"FF",X"FD",X"BB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"17",X"0F",X"07",X"03",X"00",X"00",X"00",X"00",
		X"7F",X"7D",X"FE",X"FF",X"FF",X"FF",X"BF",X"DF",X"E0",X"F0",X"F0",X"60",X"A0",X"C0",X"80",X"00",
		X"EF",X"F6",X"F8",X"E8",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"03",X"00",X"00",X"66",X"FF",X"E7",X"DB",X"BD",X"BD",
		X"03",X"07",X"07",X"0F",X"07",X"0F",X"1F",X"1F",X"BE",X"BE",X"DF",X"DB",X"EE",X"EE",X"F4",X"DC",
		X"04",X"08",X"08",X"90",X"F0",X"EC",X"DC",X"DE",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",
		X"BE",X"BE",X"FD",X"FD",X"FB",X"9B",X"37",X"37",X"40",X"80",X"C0",X"E0",X"F0",X"F0",X"E0",X"F0",
		X"5F",X"1F",X"0F",X"07",X"0F",X"0F",X"0F",X"07",X"E1",X"F3",X"E9",X"E8",X"D5",X"DF",X"BE",X"BE",
		X"07",X"07",X"03",X"03",X"00",X"00",X"00",X"00",X"BD",X"BD",X"DB",X"E7",X"FF",X"3B",X"03",X"00",
		X"8F",X"97",X"3B",X"3B",X"9D",X"ED",X"B6",X"BE",X"FC",X"F0",X"F0",X"E0",X"C0",X"C0",X"E0",X"E0",
		X"DE",X"DE",X"ED",X"F3",X"FF",X"9E",X"4A",X"00",X"E0",X"F0",X"C0",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"12",X"3F",X"9F",X"DF",X"FF",X"EF",
		X"01",X"01",X"05",X"3F",X"7F",X"3F",X"3F",X"3F",X"F7",X"FF",X"FF",X"7E",X"BC",X"F8",X"F8",X"FC",
		X"00",X"00",X"01",X"07",X"08",X"BE",X"FD",X"7D",X"00",X"00",X"80",X"C0",X"C0",X"C0",X"80",X"00",
		X"FE",X"FF",X"FF",X"FF",X"7F",X"FF",X"7F",X"7F",X"00",X"00",X"00",X"C0",X"C0",X"80",X"C0",X"C0",
		X"17",X"00",X"01",X"01",X"03",X"03",X"07",X"07",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"07",X"07",X"02",X"00",X"00",X"00",X"00",X"00",X"BF",X"1F",X"0F",X"0F",X"07",X"07",X"02",X"00",
		X"FF",X"FF",X"FE",X"FF",X"FF",X"FE",X"FE",X"FE",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"B7",X"9B",X"0D",X"0F",X"07",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"07",X"0F",X"1D",X"1E",X"00",X"0C",X"1E",X"1F",X"AE",X"EF",X"E5",X"FE",
		X"1F",X"0F",X"36",X"3B",X"1F",X"7F",X"7F",X"3F",X"7F",X"BF",X"FF",X"7F",X"FE",X"FE",X"FC",X"F8",
		X"00",X"20",X"F0",X"F6",X"EC",X"6D",X"5F",X"7B",X"00",X"00",X"00",X"00",X"C0",X"E0",X"A0",X"60",
		X"FE",X"6C",X"5F",X"3E",X"FF",X"3F",X"3F",X"7F",X"C0",X"EC",X"7A",X"F6",X"EE",X"DC",X"FC",X"F8",
		X"3F",X"7F",X"7B",X"36",X"6E",X"1D",X"2F",X"27",X"FC",X"FE",X"FF",X"7F",X"FB",X"FB",X"B7",X"6F",
		X"07",X"0D",X"1F",X"1E",X"07",X"06",X"00",X"00",X"FB",X"F7",X"77",X"EF",X"8B",X"03",X"01",X"00",
		X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FD",X"F6",X"A0",X"E0",X"F0",X"E0",X"70",X"B8",X"F0",X"F0",
		X"5F",X"5F",X"76",X"FB",X"7B",X"CD",X"87",X"00",X"60",X"F0",X"D8",X"E0",X"E0",X"80",X"00",X"00",
		X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",X"00",X"02",X"02",X"FE",X"FE",X"42",X"02",X"00",X"00",
		X"62",X"F2",X"BA",X"9A",X"9E",X"CE",X"46",X"00",X"8C",X"DE",X"F2",X"B2",X"92",X"86",X"04",X"00",
		X"08",X"FE",X"FE",X"C8",X"68",X"38",X"18",X"00",X"1C",X"BE",X"A2",X"A2",X"A2",X"E6",X"E4",X"00",
		X"0C",X"9E",X"92",X"92",X"D2",X"7E",X"3C",X"00",X"C0",X"E0",X"B0",X"9E",X"8E",X"C0",X"C0",X"00",
		X"0C",X"6E",X"9A",X"9A",X"B2",X"F2",X"6C",X"00",X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",X"00",
		X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",
		X"44",X"C6",X"82",X"82",X"C6",X"7C",X"38",X"00",X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",
		X"82",X"92",X"92",X"92",X"FE",X"FE",X"00",X"00",X"80",X"90",X"90",X"90",X"90",X"FE",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",
		X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",X"44",X"C6",X"82",X"82",X"C6",X"7C",X"38",X"00",
		X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",X"82",X"92",X"92",X"92",X"FE",X"FE",X"00",X"00",
		X"80",X"90",X"90",X"90",X"90",X"FE",X"FE",X"00",X"9E",X"9E",X"92",X"82",X"C6",X"7C",X"38",X"00",
		X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",X"82",X"82",X"FE",X"FE",X"82",X"82",X"00",X"00",
		X"FC",X"FE",X"02",X"02",X"02",X"06",X"04",X"00",X"82",X"C6",X"6E",X"3C",X"18",X"FE",X"FE",X"00",
		X"02",X"02",X"02",X"02",X"FE",X"FE",X"00",X"00",X"FE",X"FE",X"70",X"38",X"70",X"FE",X"FE",X"00",
		X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",X"00",
		X"70",X"F8",X"88",X"88",X"88",X"FE",X"FE",X"00",X"7A",X"FC",X"8E",X"8A",X"82",X"FE",X"7C",X"00",
		X"72",X"F6",X"9E",X"8C",X"88",X"FE",X"FE",X"00",X"0C",X"5E",X"D2",X"92",X"92",X"F6",X"64",X"00",
		X"80",X"80",X"FE",X"FE",X"80",X"80",X"00",X"00",X"FC",X"FE",X"02",X"02",X"02",X"FE",X"FC",X"00",
		X"F0",X"F8",X"1C",X"0E",X"1C",X"F8",X"F0",X"00",X"F8",X"FE",X"1C",X"38",X"1C",X"FE",X"F8",X"00",
		X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",X"C0",X"F0",X"1E",X"1E",X"F0",X"C0",X"00",X"00",
		X"C2",X"E2",X"F2",X"BA",X"9E",X"8E",X"86",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"10",X"10",X"18",X"7C",X"7C",X"6C",X"6E",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"6E",X"6E",X"3E",X"36",X"14",X"04",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",X"00",X"00",X"04",X"14",X"36",X"3E",X"6E",X"6E",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",X"6E",X"6C",X"7C",X"5C",X"18",X"10",X"10",X"00",
		X"00",X"00",X"00",X"08",X"04",X"00",X"00",X"08",X"30",X"78",X"C8",X"98",X"B0",X"E0",X"40",X"08",
		X"08",X"00",X"00",X"04",X"08",X"00",X"00",X"00",X"08",X"40",X"E0",X"B0",X"98",X"C8",X"78",X"30",
		X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"08",X"00",X"00",X"30",X"78",X"D8",X"B0",X"40",X"08",
		X"08",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"08",X"40",X"B0",X"D8",X"78",X"30",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"2C",X"3E",X"6E",X"6E",X"6E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"6E",X"6E",X"6E",X"3E",X"2C",X"08",X"08",X"00",
		X"00",X"08",X"08",X"2C",X"3E",X"6E",X"6E",X"6E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"6E",X"6E",X"6E",X"3E",X"2C",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"10",X"18",X"7C",X"7C",X"6C",X"6E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"6E",X"6E",X"3E",X"36",X"14",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"08",X"2C",X"3E",X"6E",X"6E",X"6E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"6E",X"6E",X"6E",X"3E",X"2C",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"04",X"14",X"36",X"3E",X"6E",X"6E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"6E",X"6C",X"7C",X"5C",X"18",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"38",X"7C",X"F8",X"00",X"04",X"0E",X"07",X"0E",X"04",X"00",X"00",
		X"F3",X"F8",X"7C",X"38",X"10",X"00",X"00",X"00",X"C0",X"00",X"00",X"04",X"0E",X"07",X"0E",X"04",
		X"00",X"00",X"00",X"00",X"00",X"07",X"0F",X"1F",X"00",X"00",X"00",X"00",X"E0",X"F0",X"DC",X"38",
		X"1C",X"27",X"3F",X"02",X"00",X"00",X"00",X"00",X"F0",X"F0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"07",X"1F",X"05",X"00",X"00",X"00",X"00",X"00",X"E0",X"F8",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"FF",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FC",X"00",X"00",X"03",X"06",X"70",X"1E",X"00",X"60",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1E",X"70",X"06",X"03",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"0E",X"00",X"F8",X"00",X"0E",X"07",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"70",X"50",X"70",X"00",X"70",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"7C",X"F0",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"F0",X"7C",X"1F",
		X"00",X"00",X"01",X"04",X"06",X"02",X"05",X"0A",X"00",X"00",X"00",X"20",X"40",X"A8",X"50",X"20",
		X"04",X"06",X"06",X"05",X"01",X"00",X"00",X"00",X"E0",X"70",X"60",X"40",X"00",X"80",X"00",X"00",
		X"00",X"20",X"22",X"33",X"0B",X"0E",X"0F",X"0E",X"00",X"00",X"84",X"08",X"10",X"F6",X"E8",X"50",
		X"0A",X"07",X"02",X"04",X"08",X"10",X"10",X"20",X"60",X"E0",X"A0",X"90",X"48",X"44",X"20",X"00",
		X"00",X"00",X"3C",X"23",X"24",X"28",X"20",X"10",X"00",X"00",X"00",X"00",X"D0",X"60",X"30",X"10",
		X"08",X"0C",X"06",X"0B",X"00",X"00",X"00",X"00",X"10",X"30",X"60",X"D8",X"38",X"38",X"00",X"00",
		X"01",X"00",X"21",X"00",X"44",X"00",X"10",X"41",X"00",X"A0",X"04",X"40",X"00",X"10",X"00",X"85",
		X"A1",X"00",X"48",X"00",X"02",X"21",X"00",X"01",X"82",X"08",X"02",X"20",X"00",X"04",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"13",X"33",X"FB",X"33",X"13",X"07",X"00",X"C0",X"01",X"BF",X"10",X"B0",X"1C",X"C4",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"13",X"33",X"FB",X"33",X"13",X"01",X"00",X"F8",X"81",X"BF",X"10",X"BF",X"81",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"13",X"33",X"FB",X"33",X"13",X"07",X"00",X"C4",X"1C",X"B0",X"10",X"BF",X"01",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"B1",X"E2",X"24",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"24",X"E2",X"B1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"04",X"01",X"12",X"22",X"00",X"00",X"00",X"00",X"30",X"08",X"00",X"00",X"C0",
		X"02",X"21",X"20",X"10",X"00",X"06",X"00",X"00",X"44",X"04",X"04",X"00",X"10",X"60",X"00",X"00",
		X"02",X"00",X"00",X"10",X"10",X"20",X"00",X"01",X"C0",X"00",X"10",X"08",X"00",X"00",X"84",X"40",
		X"20",X"22",X"00",X"00",X"10",X"00",X"00",X"06",X"80",X"04",X"04",X"00",X"00",X"10",X"00",X"40",
		X"06",X"37",X"4D",X"4D",X"59",X"79",X"36",X"00",X"3C",X"7E",X"4B",X"49",X"49",X"79",X"30",X"00",
		X"FF",X"FF",X"FF",X"C3",X"C3",X"C3",X"00",X"00",X"00",X"00",X"C3",X"C3",X"C3",X"FF",X"FF",X"FF",
		X"8E",X"DE",X"DF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"71",X"71",X"FB",X"DB",X"DB",X"8F",
		X"DB",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"C3",X"C3",X"DB",X"DB",X"DB",X"DB",
		X"0F",X"00",X"02",X"01",X"83",X"87",X"87",X"83",X"F0",X"00",X"80",X"00",X"81",X"C1",X"E1",X"E1",
		X"83",X"87",X"87",X"83",X"01",X"02",X"00",X"0F",X"E1",X"E1",X"C1",X"81",X"00",X"80",X"00",X"F0",
		X"01",X"10",X"22",X"41",X"83",X"87",X"87",X"83",X"F0",X"08",X"84",X"02",X"80",X"C0",X"E0",X"E1",
		X"83",X"07",X"07",X"03",X"41",X"22",X"10",X"0F",X"E1",X"E1",X"C1",X"81",X"02",X"84",X"08",X"80",
		X"0C",X"10",X"21",X"41",X"83",X"87",X"07",X"03",X"30",X"08",X"04",X"02",X"81",X"C1",X"E1",X"E0",
		X"03",X"87",X"87",X"83",X"41",X"21",X"10",X"0C",X"E0",X"E0",X"C1",X"81",X"02",X"04",X"08",X"70",
		X"0F",X"10",X"21",X"41",X"03",X"07",X"07",X"13",X"80",X"08",X"04",X"02",X"81",X"C1",X"E1",X"E1",
		X"83",X"87",X"87",X"83",X"41",X"21",X"10",X"01",X"E1",X"E0",X"C0",X"80",X"02",X"04",X"08",X"F0",
		X"0F",X"00",X"02",X"01",X"83",X"87",X"87",X"83",X"F0",X"00",X"80",X"00",X"81",X"C1",X"E1",X"E1",
		X"83",X"87",X"87",X"83",X"01",X"02",X"00",X"0F",X"E1",X"E1",X"C1",X"81",X"00",X"80",X"00",X"F0",
		X"01",X"10",X"22",X"41",X"83",X"87",X"87",X"83",X"F0",X"08",X"84",X"02",X"80",X"C0",X"E0",X"E1",
		X"83",X"07",X"07",X"03",X"41",X"22",X"10",X"0F",X"E1",X"E1",X"C1",X"81",X"02",X"84",X"08",X"80",
		X"0C",X"10",X"26",X"41",X"83",X"87",X"0F",X"03",X"30",X"08",X"C4",X"02",X"81",X"C1",X"E1",X"E0",
		X"03",X"87",X"87",X"83",X"41",X"26",X"10",X"0C",X"E0",X"E0",X"C1",X"81",X"02",X"C4",X"08",X"70",
		X"0F",X"10",X"21",X"41",X"03",X"07",X"07",X"83",X"80",X"08",X"04",X"02",X"81",X"C1",X"E1",X"E1",
		X"83",X"87",X"87",X"83",X"41",X"21",X"10",X"01",X"E1",X"E0",X"C0",X"80",X"02",X"04",X"08",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"0E",X"0F",X"1F",X"5F",X"EF",X"F7",
		X"03",X"07",X"0B",X"0D",X"0E",X"07",X"03",X"01",X"FB",X"FD",X"FF",X"FF",X"FE",X"7E",X"BC",X"F8",
		X"00",X"00",X"34",X"7E",X"FD",X"DB",X"F7",X"EF",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"C0",
		X"DF",X"BF",X"FF",X"FF",X"FF",X"FE",X"7D",X"1F",X"E0",X"E0",X"C0",X"B0",X"78",X"F8",X"F0",X"F0",
		X"03",X"07",X"07",X"06",X"01",X"03",X"01",X"00",X"F0",X"B1",X"7C",X"FE",X"FF",X"FF",X"FD",X"BB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"17",X"0F",X"07",X"03",X"00",X"00",X"00",X"00",
		X"7F",X"7D",X"FE",X"FF",X"FF",X"FF",X"BF",X"DF",X"E0",X"F0",X"F0",X"60",X"A0",X"C0",X"80",X"00",
		X"EF",X"F6",X"F8",X"E8",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"03",X"00",X"00",X"66",X"FF",X"E7",X"DB",X"BD",X"BD",
		X"03",X"07",X"07",X"0F",X"07",X"0F",X"1F",X"1F",X"BE",X"BE",X"DF",X"DB",X"EE",X"EE",X"F4",X"DC",
		X"04",X"08",X"08",X"90",X"F0",X"EC",X"DC",X"DE",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",
		X"BE",X"BE",X"FD",X"FD",X"FB",X"9B",X"37",X"37",X"40",X"80",X"C0",X"E0",X"F0",X"F0",X"E0",X"F0",
		X"5F",X"1F",X"0F",X"07",X"0F",X"0F",X"0F",X"07",X"E1",X"F3",X"E9",X"E8",X"D5",X"DF",X"BE",X"BE",
		X"07",X"07",X"03",X"03",X"00",X"00",X"00",X"00",X"BD",X"BD",X"DB",X"E7",X"FF",X"3B",X"03",X"00",
		X"8F",X"97",X"3B",X"3B",X"9D",X"ED",X"B6",X"BE",X"FC",X"F0",X"F0",X"E0",X"C0",X"C0",X"E0",X"E0",
		X"DE",X"DE",X"ED",X"F3",X"FF",X"9E",X"4A",X"00",X"E0",X"F0",X"C0",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"12",X"3F",X"9F",X"DF",X"FF",X"EF",
		X"01",X"01",X"05",X"3F",X"7F",X"3F",X"3F",X"3F",X"F7",X"FF",X"FF",X"7E",X"BC",X"F8",X"F8",X"FC",
		X"00",X"00",X"01",X"07",X"08",X"BE",X"FD",X"7D",X"00",X"00",X"80",X"C0",X"C0",X"C0",X"80",X"00",
		X"FE",X"FF",X"FF",X"FF",X"7F",X"FF",X"7F",X"7F",X"00",X"00",X"00",X"C0",X"C0",X"80",X"C0",X"C0",
		X"17",X"00",X"01",X"01",X"03",X"03",X"07",X"07",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"07",X"07",X"02",X"00",X"00",X"00",X"00",X"00",X"BF",X"1F",X"0F",X"0F",X"07",X"07",X"02",X"00",
		X"FF",X"FF",X"FE",X"FF",X"FF",X"FE",X"FE",X"FE",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"B7",X"9B",X"0D",X"0F",X"07",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"07",X"0F",X"1D",X"1E",X"00",X"0C",X"1E",X"1F",X"AE",X"EF",X"E5",X"FE",
		X"1F",X"0F",X"36",X"3B",X"1F",X"7F",X"7F",X"3F",X"7F",X"BF",X"FF",X"7F",X"FE",X"FE",X"FC",X"F8",
		X"00",X"20",X"F0",X"F6",X"EC",X"6D",X"5F",X"7B",X"00",X"00",X"00",X"00",X"C0",X"E0",X"A0",X"60",
		X"FE",X"6C",X"5F",X"3E",X"FF",X"3F",X"3F",X"7F",X"C0",X"EC",X"7A",X"F6",X"EE",X"DC",X"FC",X"F8",
		X"3F",X"7F",X"7B",X"36",X"6E",X"1D",X"2F",X"27",X"FC",X"FE",X"FF",X"7F",X"FB",X"FB",X"B7",X"6F",
		X"07",X"0D",X"1F",X"1E",X"07",X"06",X"00",X"00",X"FB",X"F7",X"77",X"EF",X"8B",X"03",X"01",X"00",
		X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FD",X"F6",X"A6",X"E0",X"F0",X"E0",X"70",X"B8",X"F0",X"F0",
		X"5F",X"5F",X"76",X"FB",X"7B",X"CD",X"87",X"00",X"60",X"F0",X"D8",X"E0",X"E0",X"80",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
