library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity n53xx is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(9 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of n53xx is
	type rom is array(0 to  1023) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"C7",X"C7",X"52",X"3F",X"04",X"3D",X"0B",X"80",X"90",X"58",X"1B",X"0A",X"CB",X"1B",X"71",X"B8",
		X"CA",X"12",X"23",X"1C",X"58",X"82",X"1D",X"3D",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"68",X"82",X"00",X"00",X"68",X"F9",X"00",X"00",X"69",X"1F",X"00",X"00",X"69",X"4C",X"00",X"00",
		X"6A",X"04",X"00",X"00",X"6A",X"1D",X"00",X"00",X"6A",X"37",X"00",X"00",X"6A",X"2A",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"68",X"07",X"3E",X"04",X"60",X"A2",X"5A",X"82",X"9E",X"02",X"13",X"88",X"1A",X"13",X"89",X"0A",
		X"9D",X"02",X"13",X"0A",X"13",X"1A",X"9B",X"02",X"13",X"8D",X"0A",X"97",X"02",X"13",X"0A",X"13",
		X"1D",X"C4",X"59",X"80",X"13",X"0B",X"2F",X"0F",X"08",X"1D",X"13",X"38",X"FD",X"4C",X"F7",X"5A",
		X"80",X"09",X"FD",X"08",X"09",X"FD",X"FD",X"5A",X"80",X"19",X"FD",X"08",X"19",X"59",X"81",X"39",
		X"D1",X"4D",X"CB",X"5A",X"82",X"09",X"D1",X"08",X"09",X"D1",X"D1",X"5A",X"82",X"19",X"D1",X"08",
		X"19",X"59",X"81",X"3A",X"68",X"E6",X"5A",X"84",X"4E",X"E2",X"09",X"68",X"E6",X"08",X"09",X"68",
		X"E6",X"E6",X"19",X"E6",X"08",X"19",X"59",X"81",X"3B",X"F8",X"5A",X"86",X"4F",X"F4",X"09",X"F8",
		X"08",X"09",X"F8",X"F8",X"19",X"F8",X"08",X"19",X"2C",X"3E",X"04",X"5A",X"80",X"13",X"0A",X"13",
		X"0A",X"9E",X"02",X"13",X"0A",X"13",X"1A",X"9D",X"02",X"13",X"84",X"1A",X"13",X"85",X"0A",X"9B",
		X"02",X"13",X"0A",X"13",X"1A",X"97",X"02",X"13",X"88",X"1A",X"13",X"89",X"1D",X"68",X"FC",X"3E",
		X"04",X"5A",X"80",X"9E",X"02",X"13",X"0A",X"13",X"0A",X"13",X"0A",X"13",X"0A",X"9D",X"02",X"13",
		X"0A",X"13",X"0A",X"13",X"0A",X"13",X"0A",X"9B",X"02",X"13",X"0A",X"13",X"0A",X"13",X"0A",X"13",
		X"0A",X"97",X"02",X"13",X"0A",X"13",X"0A",X"13",X"0A",X"13",X"69",X"22",X"3E",X"04",X"61",X"51",
		X"CE",X"59",X"80",X"9E",X"02",X"13",X"0A",X"13",X"0A",X"13",X"0A",X"13",X"0A",X"9D",X"02",X"13",
		X"0A",X"13",X"0A",X"13",X"0A",X"13",X"0A",X"9B",X"02",X"13",X"0A",X"13",X"0A",X"13",X"0A",X"13",
		X"0A",X"97",X"02",X"13",X"0A",X"13",X"0A",X"13",X"0A",X"13",X"0A",X"90",X"38",X"69",X"90",X"91",
		X"39",X"D0",X"92",X"3A",X"D0",X"93",X"3B",X"D0",X"08",X"69",X"7B",X"5A",X"9F",X"0A",X"1D",X"2C",
		X"1D",X"14",X"23",X"0C",X"23",X"0C",X"1F",X"1D",X"14",X"23",X"1C",X"23",X"1C",X"72",X"5B",X"1D",
		X"B2",X"FC",X"59",X"0D",X"5B",X"7F",X"69",X"F1",X"71",X"B8",X"EF",X"90",X"1D",X"69",X"FA",X"B9",
		X"F5",X"90",X"1D",X"69",X"FA",X"BA",X"69",X"E8",X"90",X"1D",X"69",X"FA",X"B5",X"69",X"D9",X"59",
		X"0D",X"5B",X"7F",X"69",X"E8",X"71",X"BB",X"CC",X"91",X"1D",X"69",X"FA",X"BD",X"D2",X"90",X"1D",
		X"69",X"FA",X"BF",X"69",X"F1",X"97",X"1D",X"69",X"FA",X"B4",X"E1",X"59",X"0D",X"5B",X"75",X"F1",
		X"E8",X"B3",X"E8",X"59",X"0D",X"5B",X"7F",X"F1",X"9E",X"02",X"12",X"4C",X"EE",X"F1",X"91",X"2F",
		X"1D",X"9D",X"02",X"12",X"4C",X"F7",X"FA",X"94",X"2F",X"1D",X"0D",X"53",X"59",X"0D",X"5A",X"80",
		X"0A",X"53",X"1D",X"2C",X"3F",X"FF",X"90",X"07",X"3E",X"20",X"61",X"51",X"5A",X"80",X"0D",X"23",
		X"01",X"08",X"0D",X"21",X"01",X"9F",X"3B",X"D9",X"90",X"07",X"3E",X"20",X"CA",X"3E",X"04",X"60",
		X"A2",X"5A",X"82",X"13",X"88",X"1A",X"13",X"89",X"1D",X"DF",X"3E",X"04",X"5A",X"80",X"13",X"0A",
		X"13",X"0A",X"13",X"0A",X"13",X"1D",X"EC",X"3E",X"04",X"59",X"80",X"9E",X"02",X"13",X"0A",X"13",
		X"1A",X"9D",X"02",X"13",X"82",X"1A",X"13",X"83",X"0A",X"9B",X"02",X"13",X"0A",X"13",X"1A",X"97",
		X"02",X"13",X"86",X"1A",X"13",X"87",X"1D",X"80",X"90",X"38",X"EF",X"71",X"39",X"EF",X"71",X"3A",
		X"EF",X"71",X"3B",X"EF",X"71",X"08",X"08",X"A8",X"D9",X"9F",X"5A",X"80",X"0A",X"1D",X"F4",X"5A",
		X"80",X"0A",X"90",X"1D",X"59",X"81",X"90",X"38",X"6A",X"91",X"71",X"39",X"6A",X"91",X"71",X"3A",
		X"6A",X"91",X"71",X"3B",X"D1",X"71",X"08",X"08",X"A9",X"6A",X"77",X"9F",X"5A",X"82",X"0A",X"1A",
		X"D6",X"5A",X"82",X"0A",X"90",X"1A",X"13",X"84",X"1A",X"13",X"85",X"1D",X"6A",X"39",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"6B",X"4A",X"00",X"00",X"6B",X"37",X"00",X"00",X"6B",X"4A",X"00",X"00",X"6B",X"02",X"00",X"00",
		X"E0",X"00",X"00",X"00",X"6B",X"37",X"00",X"00",X"6B",X"24",X"00",X"00",X"6B",X"11",X"00",X"00",
		X"52",X"3E",X"04",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"6A",X"E0",X"52",X"50",X"1B",X"51",X"54",X"5A",X"0D",X"23",X"01",X"08",X"0D",X"21",X"01",X"6B",
		X"59",X"52",X"50",X"1B",X"51",X"54",X"5A",X"0D",X"23",X"01",X"08",X"0D",X"21",X"01",X"08",X"A4",
		X"6B",X"64",X"6B",X"59",X"52",X"50",X"1B",X"51",X"54",X"5A",X"0D",X"23",X"01",X"08",X"0D",X"21",
		X"01",X"08",X"A6",X"6B",X"64",X"6B",X"59",X"52",X"50",X"1B",X"51",X"54",X"5A",X"0D",X"23",X"01",
		X"08",X"0D",X"21",X"01",X"08",X"AA",X"6B",X"64",X"6B",X"59",X"52",X"50",X"1B",X"51",X"54",X"5A",
		X"0D",X"23",X"01",X"08",X"0D",X"21",X"01",X"08",X"E4",X"25",X"DC",X"D9",X"25",X"DC",X"9F",X"23",
		X"01",X"21",X"01",X"80",X"54",X"51",X"1B",X"50",X"3E",X"04",X"3C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
