library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity gfx3 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of gfx3 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"01",X"00",X"13",X"00",X"33",X"01",X"33",X"01",X"33",X"13",X"33",X"13",X"33",X"13",X"33",
		X"11",X"11",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"11",X"33",X"00",
		X"13",X"33",X"13",X"33",X"13",X"33",X"13",X"33",X"13",X"33",X"13",X"33",X"13",X"33",X"13",X"33",
		X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"11",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"CC",X"0C",X"CC",X"CC",X"AC",X"CC",X"A5",X"C0",X"CA",X"05",X"56",X"5C",X"AA",X"5C",X"FF",
		X"A0",X"CC",X"5C",X"5C",X"FC",X"C5",X"5A",X"A5",X"FC",X"5A",X"5F",X"C5",X"5F",X"CA",X"F5",X"6F",
		X"5F",X"AF",X"C5",X"F5",X"CC",X"5A",X"C5",X"CF",X"05",X"C5",X"CC",X"5C",X"00",X"FA",X"00",X"05",
		X"AF",X"5F",X"F5",X"FF",X"54",X"65",X"AA",X"AC",X"F6",X"AA",X"AF",X"5C",X"55",X"C5",X"FC",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CF",X"00",X"55",X"00",X"FC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"CC",X"00",X"0F",X"00",X"55",X"00",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"5A",X"00",X"CC",X"C0",X"AC",X"00",X"FA",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"FF",X"0E",X"FF",X"00",X"EE",X"00",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"E0",X"FF",X"E0",X"FF",X"E0",X"FF",X"00",X"EE",X"00",X"00",X"00",
		X"00",X"0C",X"00",X"CB",X"00",X"CB",X"00",X"CB",X"0C",X"CB",X"00",X"BC",X"00",X"BB",X"00",X"BB",
		X"FF",X"C0",X"CF",X"BC",X"FF",X"FF",X"BB",X"FF",X"CF",X"FF",X"CF",X"FF",X"CC",X"FF",X"FF",X"FB",
		X"C0",X"FF",X"BC",X"FF",X"BC",X"FF",X"BB",X"FF",X"CB",X"FF",X"0C",X"BB",X"CB",X"C4",X"BB",X"04",
		X"FF",X"F4",X"FF",X"BC",X"FB",X"BC",X"F4",X"44",X"4C",X"CC",X"C0",X"00",X"00",X"00",X"4C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"05",X"00",X"0A",X"00",X"0A",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",
		X"6A",X"00",X"5F",X"00",X"F5",X"00",X"F6",X"00",X"5A",X"00",X"F6",X"00",X"50",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"56",X"00",
		X"00",X"00",X"00",X"0A",X"00",X"06",X"00",X"06",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A6",X"00",X"5F",X"00",X"56",X"00",X"5A",X"00",X"A6",X"00",X"55",X"00",X"5A",X"00",X"50",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5A",X"00",
		X"00",X"06",X"00",X"65",X"00",X"65",X"00",X"A6",X"00",X"AA",X"00",X"0A",X"00",X"00",X"00",X"00",
		X"A6",X"00",X"66",X"00",X"F6",X"00",X"AF",X"00",X"AF",X"00",X"A5",X"00",X"A0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"5A",X"00",X"A1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"56",X"00",X"FF",X"00",
		X"00",X"A5",X"00",X"65",X"00",X"65",X"00",X"AF",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"00",X"F5",X"00",X"65",X"00",X"56",X"00",X"5A",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"65",X"00",X"5F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"F6",X"00",X"66",X"00",
		X"00",X"5F",X"00",X"5F",X"00",X"65",X"00",X"66",X"00",X"6F",X"00",X"AA",X"00",X"00",X"00",X"00",
		X"FF",X"A0",X"AA",X"A0",X"FA",X"F0",X"FA",X"F0",X"5A",X"00",X"5A",X"00",X"AA",X"00",X"A0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"AF",X"00",X"F5",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"55",X"00",X"6A",X"00",X"A6",X"00",
		X"00",X"AA",X"00",X"AF",X"00",X"15",X"00",X"5F",X"00",X"55",X"00",X"66",X"00",X"5A",X"00",X"05",
		X"FF",X"00",X"55",X"A0",X"A5",X"A0",X"F5",X"A0",X"AF",X"50",X"AF",X"00",X"F5",X"00",X"56",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"6A",X"00",X"6A",X"00",X"F5",
		X"00",X"00",X"00",X"00",X"60",X"00",X"A0",X"00",X"AA",X"00",X"66",X"00",X"FF",X"50",X"55",X"F0",
		X"00",X"F5",X"00",X"F5",X"00",X"F6",X"00",X"5F",X"00",X"66",X"00",X"56",X"00",X"A5",X"00",X"00",
		X"AA",X"F5",X"A5",X"A5",X"AF",X"AA",X"66",X"AA",X"6F",X"A0",X"F5",X"50",X"5A",X"00",X"55",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"5A",X"00",X"F1",X"00",X"A1",X"00",X"A6",
		X"00",X"00",X"00",X"00",X"A0",X"00",X"65",X"00",X"65",X"00",X"FF",X"00",X"F5",X"50",X"5A",X"A0",
		X"05",X"AF",X"0F",X"6F",X"0A",X"5A",X"0A",X"FA",X"00",X"A6",X"00",X"66",X"00",X"5F",X"00",X"05",
		X"FF",X"FA",X"56",X"AF",X"55",X"AF",X"FF",X"5A",X"5F",X"50",X"55",X"A0",X"65",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"5A",X"00",X"FF",X"00",X"F1",X"00",X"F1",
		X"00",X"00",X"A0",X"00",X"55",X"00",X"5A",X"00",X"FA",X"00",X"A5",X"60",X"A5",X"56",X"AF",X"A5",
		X"0A",X"5A",X"0A",X"65",X"0A",X"6F",X"00",X"5A",X"00",X"AA",X"00",X"66",X"00",X"AA",X"00",X"00",
		X"5A",X"55",X"F5",X"A5",X"F5",X"AA",X"F6",X"5A",X"A5",X"AA",X"55",X"A0",X"F6",X"00",X"AA",X"00",
		X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"FF",X"00",X"F5",X"05",X"15",X"05",X"16",X"56",X"66",
		X"00",X"00",X"A0",X"00",X"AA",X"00",X"FF",X"00",X"55",X"A0",X"A6",X"5A",X"65",X"55",X"AA",X"A5",
		X"5F",X"A6",X"6F",X"5A",X"A6",X"5F",X"0A",X"FF",X"0A",X"AA",X"00",X"55",X"00",X"AA",X"00",X"0A",
		X"AA",X"AA",X"5A",X"5A",X"65",X"FA",X"65",X"FA",X"5A",X"FA",X"5A",X"F0",X"AA",X"00",X"A5",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"50",X"00",X"01",X"00",X"01",X"00",X"11",
		X"50",X"00",X"00",X"00",X"00",X"11",X"11",X"FE",X"1F",X"EE",X"FE",X"EE",X"EF",X"EE",X"EE",X"E0",
		X"00",X"11",X"00",X"1F",X"00",X"11",X"00",X"1F",X"00",X"11",X"00",X"01",X"55",X"01",X"00",X"00",
		X"FE",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"FE",X"00",X"1E",X"00",
		X"00",X"00",X"00",X"11",X"00",X"1F",X"00",X"F1",X"01",X"FE",X"01",X"1F",X"11",X"EE",X"1E",X"EE",
		X"1F",X"10",X"EF",X"EF",X"1E",X"EE",X"EE",X"EE",X"EE",X"0E",X"EE",X"00",X"E0",X"00",X"00",X"00",
		X"1F",X"FE",X"1E",X"FE",X"1F",X"EE",X"1E",X"FE",X"1F",X"EE",X"01",X"EE",X"01",X"EE",X"00",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"05",X"00",X"05",X"00",X"00",X"00",X"00",X"50",X"00",X"05",X"00",X"00",X"01",
		X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"00",X"00",X"00",X"01",X"10",X"11",X"11",X"1E",X"EF",
		X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"1F",X"00",X"EF",X"00",X"1E",X"00",X"FE",X"00",X"0E",
		X"FF",X"EE",X"EE",X"EE",X"EE",X"00",X"EE",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"00",X"11",X"00",X"1F",X"01",X"E1",X"01",X"EE",X"11",X"FE",X"11",X"EE",
		X"11",X"10",X"11",X"11",X"F1",X"EF",X"EE",X"EE",X"EE",X"EF",X"FE",X"EE",X"EE",X"0E",X"EE",X"00",
		X"11",X"EE",X"11",X"EE",X"1E",X"EE",X"1E",X"EE",X"01",X"E0",X"01",X"00",X"0E",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"0E",X"EE",
		X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",
		X"11",X"FE",X"11",X"EE",X"1E",X"E0",X"E1",X"00",X"1E",X"00",X"FE",X"00",X"EE",X"00",X"1E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"50",X"00",X"01",
		X"50",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"11",X"1F",X"E1",X"EE",X"FE",X"EE",X"FE",X"00",
		X"00",X"01",X"00",X"1E",X"00",X"11",X"00",X"1E",X"00",X"11",X"00",X"01",X"55",X"01",X"00",X"00",
		X"EE",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"E0",X"00",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"50",X"00",X"50",X"00",X"05",X"00",X"05",X"00",X"00",X"11",X"00",X"11",
		X"00",X"50",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"1E",X"11",X"EF",X"11",X"FE",X"1E",X"E0",X"EF",X"00",X"FE",X"00",X"FE",X"00",X"1E",X"00",
		X"00",X"50",X"00",X"50",X"00",X"05",X"00",X"05",X"00",X"00",X"00",X"00",X"50",X"01",X"05",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"01",X"11",X"11",X"1E",X"EF",X"FF",X"EE",
		X"00",X"11",X"00",X"11",X"00",X"EF",X"00",X"EF",X"00",X"1E",X"00",X"FE",X"00",X"EE",X"00",X"FE",
		X"EE",X"EE",X"EE",X"00",X"EE",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"FF",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FA",X"00",X"FF",X"C0",X"FF",X"AC",
		X"0F",X"FF",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CF",X"FF",X"0C",X"FF",X"00",X"CC",
		X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"AA",X"CC",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"AC",X"00",X"AA",X"00",X"FA",X"00",X"FA",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"CF",X"00",X"0C",
		X"FF",X"00",X"FF",X"00",X"FF",X"C0",X"FF",X"AA",X"FF",X"FF",X"FF",X"FA",X"FF",X"AC",X"CC",X"C0",
		X"00",X"FF",X"00",X"FF",X"0F",X"FF",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CF",X"AA",
		X"FC",X"00",X"FF",X"00",X"FF",X"C0",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"AA",X"FF",X"CC",X"AF",
		X"0C",X"AC",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"CA",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"FF",X"00",X"FF",X"0F",X"FF",X"0F",X"FF",X"FF",X"FF",
		X"00",X"00",X"FF",X"C0",X"FF",X"C0",X"FA",X"00",X"FA",X"00",X"AA",X"00",X"AC",X"00",X"AC",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CA",X"FA",X"0C",X"AA",X"00",X"CC",X"00",X"00",
		X"AC",X"00",X"AC",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"FF",X"00",X"F3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"32",X"00",X"33",X"C0",X"33",X"2C",
		X"03",X"33",X"03",X"33",X"33",X"33",X"33",X"33",X"33",X"32",X"33",X"22",X"03",X"2C",X"0C",X"C0",
		X"33",X"22",X"33",X"22",X"33",X"32",X"33",X"32",X"33",X"32",X"C3",X"32",X"00",X"22",X"00",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"9F",X"00",X"9F",X"00",X"99",X"00",X"99",
		X"00",X"00",X"99",X"C0",X"F9",X"8C",X"99",X"8C",X"99",X"88",X"99",X"88",X"99",X"88",X"99",X"8C",
		X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"CC",
		X"99",X"8C",X"98",X"C0",X"98",X"00",X"88",X"00",X"98",X"00",X"98",X"00",X"88",X"00",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"0F",X"00",X"6F",X"00",X"6F",X"00",X"6F",X"00",X"66",
		X"00",X"00",X"55",X"00",X"65",X"00",X"66",X"C0",X"66",X"C0",X"66",X"5C",X"66",X"5C",X"66",X"5C",
		X"00",X"66",X"00",X"66",X"00",X"66",X"00",X"66",X"00",X"66",X"00",X"66",X"00",X"C6",X"00",X"0C",
		X"66",X"5C",X"66",X"5C",X"66",X"5C",X"66",X"5C",X"66",X"5C",X"66",X"5C",X"66",X"C0",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"FA",X"00",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"AC",X"00",X"AB",X"00",X"AA",X"C0",X"AA",X"BC",X"AA",X"BC",
		X"00",X"AA",X"00",X"AA",X"00",X"0B",X"00",X"00",X"00",X"0A",X"00",X"0A",X"00",X"0C",X"00",X"00",
		X"AA",X"BB",X"AA",X"BB",X"AA",X"BB",X"AA",X"BB",X"AA",X"BB",X"AA",X"BB",X"AA",X"BC",X"CC",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"00",
		X"00",X"00",X"00",X"00",X"77",X"00",X"77",X"00",X"77",X"00",X"73",X"00",X"33",X"00",X"33",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"7F",X"00",X"71",X"00",X"77",X"00",X"07",X"00",X"00",
		X"00",X"00",X"70",X"00",X"73",X"00",X"73",X"00",X"73",X"00",X"33",X"00",X"33",X"00",X"3C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"07",X"00",X"7F",X"00",X"71",X"00",X"77",X"00",X"77",X"00",X"07",X"00",X"00",
		X"73",X"00",X"77",X"00",X"77",X"C0",X"77",X"C0",X"77",X"C0",X"73",X"C0",X"33",X"00",X"33",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",
		X"00",X"7F",X"00",X"F1",X"00",X"11",X"00",X"77",X"00",X"77",X"00",X"77",X"00",X"77",X"00",X"03",
		X"73",X"00",X"77",X"C0",X"77",X"C0",X"77",X"C0",X"73",X"C0",X"73",X"C0",X"33",X"00",X"33",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"77",X"C0",
		X"00",X"7F",X"00",X"7F",X"00",X"77",X"00",X"77",X"00",X"77",X"00",X"77",X"00",X"33",X"00",X"00",
		X"77",X"C0",X"77",X"3C",X"77",X"3C",X"77",X"3C",X"73",X"3C",X"33",X"C0",X"33",X"C0",X"33",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"F1",X"00",X"F1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"77",X"C0",X"77",X"C0",
		X"00",X"F1",X"00",X"17",X"00",X"77",X"00",X"77",X"00",X"77",X"00",X"77",X"00",X"33",X"00",X"03",
		X"77",X"3C",X"77",X"3C",X"77",X"3C",X"73",X"3C",X"33",X"3C",X"33",X"C0",X"33",X"C0",X"33",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"00",X"FF",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"77",X"C0",X"77",X"3C",X"77",X"3C",
		X"00",X"11",X"00",X"77",X"00",X"77",X"00",X"77",X"00",X"77",X"00",X"77",X"00",X"33",X"00",X"00",
		X"77",X"33",X"77",X"33",X"77",X"33",X"77",X"33",X"77",X"3C",X"33",X"3C",X"33",X"C0",X"33",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"77",X"00",X"F1",X"00",X"F1",X"07",X"17",
		X"00",X"00",X"00",X"00",X"00",X"00",X"73",X"00",X"77",X"C0",X"77",X"3C",X"77",X"3C",X"77",X"33",
		X"07",X"17",X"07",X"77",X"07",X"77",X"07",X"77",X"00",X"77",X"00",X"77",X"00",X"33",X"00",X"03",
		X"77",X"33",X"77",X"33",X"77",X"33",X"73",X"33",X"33",X"3C",X"33",X"3C",X"33",X"C0",X"33",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"00",X"FF",X"00",X"F1",X"00",X"F7",X"07",X"17",
		X"00",X"00",X"00",X"00",X"77",X"00",X"77",X"C0",X"77",X"3C",X"77",X"33",X"77",X"33",X"77",X"33",
		X"07",X"77",X"07",X"77",X"07",X"77",X"00",X"77",X"00",X"77",X"00",X"77",X"00",X"33",X"00",X"00",
		X"77",X"33",X"77",X"33",X"77",X"33",X"77",X"33",X"73",X"33",X"33",X"3C",X"33",X"C0",X"33",X"00",
		X"00",X"00",X"00",X"07",X"00",X"F1",X"00",X"F1",X"07",X"17",X"07",X"77",X"7F",X"77",X"71",X"77",
		X"00",X"00",X"73",X"00",X"77",X"C0",X"77",X"3C",X"77",X"33",X"77",X"33",X"77",X"33",X"77",X"33",
		X"77",X"77",X"77",X"77",X"77",X"77",X"07",X"77",X"03",X"77",X"00",X"33",X"00",X"33",X"00",X"03",
		X"77",X"33",X"77",X"33",X"73",X"33",X"33",X"33",X"33",X"33",X"33",X"3C",X"33",X"C0",X"33",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"30",X"00",X"30",X"00",X"30",X"33",X"30",X"33",X"30",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"33",X"00",X"33",X"00",X"BC",X"0B",X"BB",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"FF",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"03",X"3C",X"FF",X"33",X"FF",X"F3",X"FF",X"F3",X"FF",X"F3",X"FF",X"F3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"00",X"33",X"00",X"33",X"00",X"33",X"C0",
		X"FF",X"33",X"33",X"33",X"BB",X"B3",X"CC",X"CB",X"CC",X"CB",X"BB",X"CB",X"BB",X"CB",X"BB",X"CB",
		X"3F",X"FF",X"FF",X"CF",X"FF",X"CF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"FF",X"32",X"2C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"77",X"00",X"77",X"00",X"73",X"00",X"33",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"77",X"00",X"77",X"00",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BC",X"CB",X"CF",X"0C",X"FF",X"00",X"2F",X"00",X"2F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"22",X"00",X"22",X"00",X"2C",X"00",X"C2",X"00",X"22",X"00",X"CC",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"22",X"BB",X"22",X"BB",X"CC",X"BB",X"00",X"BB",X"00",X"CC",
		X"FB",X"B3",X"FF",X"F3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"FF",X"F3",X"FF",X"32",
		X"33",X"2C",X"32",X"2C",X"22",X"C0",X"22",X"00",X"22",X"22",X"22",X"22",X"22",X"CC",X"CC",X"00",
		X"FF",X"22",X"FF",X"22",X"B2",X"2C",X"BB",X"C0",X"BB",X"00",X"BC",X"00",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"99",
		X"00",X"00",X"09",X"00",X"9C",X"C0",X"99",X"99",X"99",X"98",X"98",X"88",X"88",X"44",X"84",X"41",
		X"00",X"98",X"00",X"98",X"00",X"98",X"00",X"98",X"00",X"88",X"00",X"84",X"00",X"84",X"00",X"84",
		X"44",X"11",X"41",X"1B",X"11",X"B4",X"11",X"41",X"1B",X"11",X"14",X"11",X"B4",X"1B",X"B4",X"B4",
		X"00",X"00",X"00",X"C0",X"09",X"8C",X"99",X"98",X"99",X"99",X"88",X"99",X"48",X"89",X"14",X"88",
		X"00",X"00",X"00",X"00",X"99",X"00",X"FF",X"C0",X"CF",X"C0",X"89",X"C0",X"88",X"C0",X"88",X"C0",
		X"11",X"48",X"B1",X"14",X"44",X"11",X"11",X"41",X"11",X"41",X"44",X"14",X"CC",X"14",X"CC",X"14",
		X"88",X"C0",X"88",X"C0",X"88",X"8C",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"99",
		X"00",X"00",X"09",X"00",X"9C",X"C0",X"99",X"99",X"99",X"98",X"98",X"88",X"88",X"44",X"84",X"41",
		X"00",X"98",X"00",X"98",X"00",X"98",X"00",X"98",X"00",X"88",X"00",X"84",X"00",X"84",X"00",X"84",
		X"44",X"11",X"41",X"1B",X"11",X"B4",X"11",X"41",X"1B",X"11",X"14",X"11",X"B4",X"1B",X"B4",X"B4",
		X"00",X"00",X"00",X"C0",X"09",X"8C",X"99",X"98",X"99",X"99",X"88",X"99",X"48",X"89",X"14",X"88",
		X"00",X"00",X"00",X"00",X"99",X"00",X"FF",X"C0",X"CF",X"C0",X"89",X"C0",X"88",X"C0",X"88",X"C0",
		X"11",X"48",X"B1",X"14",X"44",X"11",X"11",X"41",X"11",X"41",X"44",X"14",X"CC",X"14",X"CC",X"14",
		X"88",X"C0",X"88",X"C0",X"88",X"8C",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"00",X"84",X"00",X"84",X"00",X"84",X"00",X"88",X"00",X"88",X"00",X"F8",X"00",X"FF",X"00",X"8F",
		X"41",X"B4",X"41",X"B4",X"BC",X"55",X"C5",X"55",X"55",X"5C",X"55",X"5C",X"55",X"5C",X"55",X"C5",
		X"09",X"99",X"99",X"8C",X"88",X"8C",X"C8",X"8C",X"0C",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"41",X"CC",X"41",X"55",X"44",X"55",X"C1",X"55",X"88",X"55",X"88",X"55",X"FF",X"55",X"FF",
		X"48",X"88",X"48",X"88",X"88",X"88",X"88",X"89",X"FF",X"C9",X"CC",X"98",X"99",X"88",X"99",X"88",
		X"5C",X"FC",X"5C",X"C9",X"5C",X"09",X"C0",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"88",X"98",X"88",X"88",X"8C",X"88",X"8C",X"CC",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"84",X"00",X"84",X"00",X"84",X"00",X"88",X"00",X"88",X"00",X"88",X"00",X"88",X"00",X"88",
		X"41",X"B4",X"41",X"B4",X"BC",X"B4",X"55",X"54",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"09",X"99",X"99",X"88",X"88",X"88",X"C8",X"88",X"0C",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"CC",X"CF",X"FF",X"0C",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"41",X"CC",X"41",X"CC",X"44",X"55",X"C1",X"55",X"88",X"55",X"88",X"C5",X"FF",X"5C",X"FF",
		X"48",X"88",X"48",X"88",X"88",X"88",X"88",X"89",X"88",X"C9",X"CC",X"98",X"99",X"88",X"99",X"88",
		X"CF",X"FC",X"FF",X"C9",X"CC",X"09",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"88",X"98",X"88",X"88",X"8C",X"88",X"8C",X"CC",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"99",
		X"00",X"00",X"09",X"00",X"9C",X"C0",X"99",X"99",X"99",X"98",X"98",X"88",X"88",X"88",X"88",X"44",
		X"00",X"98",X"00",X"98",X"00",X"98",X"00",X"98",X"00",X"88",X"00",X"88",X"00",X"DD",X"00",X"FF",
		X"84",X"BB",X"4B",X"11",X"B1",X"44",X"B1",X"BB",X"55",X"55",X"55",X"55",X"55",X"CC",X"CC",X"FF",
		X"00",X"00",X"00",X"C0",X"09",X"8C",X"99",X"98",X"99",X"99",X"88",X"99",X"88",X"89",X"88",X"88",
		X"00",X"00",X"00",X"00",X"99",X"00",X"FF",X"C0",X"CF",X"C0",X"89",X"C0",X"88",X"C0",X"88",X"C0",
		X"44",X"88",X"BB",X"88",X"44",X"48",X"BB",X"B4",X"11",X"4B",X"11",X"4B",X"D1",X"B4",X"FD",X"11",
		X"88",X"C0",X"88",X"C0",X"88",X"8C",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"99",X"00",X"99",
		X"00",X"00",X"09",X"00",X"9C",X"C0",X"99",X"99",X"99",X"98",X"98",X"88",X"88",X"88",X"88",X"FF",
		X"00",X"98",X"00",X"98",X"00",X"98",X"00",X"98",X"00",X"88",X"00",X"88",X"00",X"8F",X"00",X"8F",
		X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"C0",X"09",X"8C",X"99",X"98",X"99",X"99",X"88",X"99",X"88",X"89",X"88",X"88",
		X"00",X"00",X"00",X"00",X"99",X"00",X"FF",X"C0",X"CF",X"C0",X"89",X"C0",X"88",X"C0",X"88",X"C0",
		X"FF",X"88",X"FF",X"88",X"FF",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"88",X"C0",X"88",X"C0",X"88",X"8C",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"8F",X"00",X"88",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"09",X"99",X"99",X"88",X"88",X"88",X"C8",X"8C",X"0C",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"CF",X"FF",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"DD",X"FF",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"EE",
		X"48",X"88",X"B4",X"88",X"D4",X"88",X"ED",X"89",X"E8",X"C9",X"CC",X"98",X"99",X"88",X"99",X"88",
		X"FF",X"EC",X"EE",X"C9",X"CC",X"09",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"88",X"98",X"88",X"88",X"8C",X"88",X"8C",X"CC",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"8F",X"00",X"8F",X"00",X"8F",X"00",X"88",X"00",X"88",X"00",X"88",X"00",X"88",X"00",X"88",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"09",X"99",X"99",X"88",X"88",X"88",X"C8",X"8C",X"0C",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"CC",X"FF",X"C0",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"EE",
		X"E8",X"88",X"EE",X"88",X"EE",X"88",X"EE",X"89",X"E8",X"C9",X"CC",X"98",X"99",X"88",X"99",X"88",
		X"FF",X"EC",X"EE",X"C9",X"CC",X"09",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"88",X"98",X"88",X"88",X"8C",X"88",X"8C",X"CC",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"99",X"00",X"44",X"09",X"CC",X"94",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"C9",X"44",X"44",X"CB",X"BB",X"5C",X"11",
		X"9B",X"55",X"41",X"CC",X"4C",X"FF",X"CF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"11",X"CC",X"41",X"EE",X"CC",X"FF",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"8C",X"FF",X"89",X"CF",X"48",X"FF",X"B4",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"9C",X"00",
		X"1B",X"88",X"11",X"88",X"11",X"48",X"CC",X"48",X"EE",X"B4",X"FE",X"C4",X"FF",X"EC",X"FF",X"EE",
		X"89",X"00",X"89",X"00",X"88",X"00",X"88",X"00",X"88",X"00",X"88",X"C0",X"88",X"C0",X"88",X"8C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"89",X"00",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"88",X"88",X"99",X"88",X"99",X"99",X"99",X"99",
		X"00",X"FF",X"00",X"CF",X"00",X"99",X"00",X"99",X"09",X"99",X"09",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"00",X"00",X"00",X"00",X"CC",X"C0",X"88",X"8C",X"88",X"88",X"98",X"88",X"99",X"98",X"99",X"98",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"88",X"00",X"88",X"00",X"88",X"C0",
		X"99",X"9F",X"99",X"FF",X"99",X"CC",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"98",X"99",X"88",
		X"88",X"8C",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"8C",X"88",
		X"0F",X"FF",X"0F",X"FF",X"0C",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"CC",X"00",X"00",X"00",X"09",X"00",X"99",X"00",X"99",X"00",X"98",X"00",X"88",X"00",X"C8",
		X"FF",X"FF",X"FF",X"FF",X"88",X"EE",X"8C",X"CC",X"8C",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",
		X"FF",X"EE",X"FF",X"EE",X"FF",X"EE",X"FF",X"EE",X"FF",X"EE",X"FF",X"EE",X"FF",X"EE",X"FF",X"EE",
		X"98",X"88",X"98",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"FF",X"EE",X"EE",X"EE",X"EE",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"99",
		X"98",X"8C",X"98",X"8C",X"98",X"8C",X"88",X"C0",X"88",X"C0",X"99",X"00",X"98",X"00",X"98",X"C0",
		X"99",X"89",X"99",X"89",X"18",X"99",X"41",X"98",X"C4",X"11",X"04",X"15",X"0C",X"45",X"00",X"CC",
		X"99",X"88",X"99",X"C8",X"99",X"98",X"88",X"85",X"55",X"5C",X"55",X"C1",X"55",X"44",X"55",X"CC",
		X"00",X"FF",X"09",X"9F",X"99",X"99",X"99",X"98",X"98",X"88",X"88",X"88",X"CC",X"88",X"00",X"CC",
		X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",X"CF",X"FF",X"CC",X"CC",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"99",X"88",X"88",X"18",X"11",X"1C",X"11",X"CF",X"11",X"FF",X"1C",X"FF",X"CF",X"FF",X"FF",X"FF",
		X"C9",X"88",X"98",X"88",X"88",X"88",X"88",X"88",X"88",X"8C",X"88",X"8C",X"88",X"8C",X"88",X"88",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"CC",X"FC",X"00",X"C0",X"00",X"00",X"00",X"00",X"08",X"00",X"0C",
		X"88",X"88",X"C8",X"88",X"08",X"88",X"88",X"88",X"88",X"88",X"88",X"8C",X"88",X"8C",X"88",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"33",X"03",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"33",X"00",X"33",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"BC",X"0B",X"BB",X"BB",X"BB",X"BF",X"BB",X"FF",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CB",X"00",X"FB",X"C0",
		X"33",X"F3",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"3C",X"33",X"3F",X"33",X"FF",X"33",X"FF",
		X"3B",X"BC",X"CF",X"BC",X"FF",X"C0",X"FB",X"00",X"BB",X"BC",X"BB",X"C0",X"FB",X"BB",X"F3",X"FC",
		X"00",X"00",X"0F",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",X"FF",X"03",X"33",
		X"00",X"00",X"00",X"FF",X"00",X"FF",X"80",X"FF",X"80",X"FF",X"80",X"FF",X"80",X"FF",X"80",X"33",
		X"03",X"33",X"03",X"33",X"03",X"33",X"03",X"33",X"03",X"33",X"03",X"33",X"03",X"33",X"03",X"33",
		X"80",X"33",X"80",X"33",X"80",X"33",X"80",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"33",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"33",X"33",
		X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"38",X"33",X"38",X"33",X"38",X"33",X"38",
		X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"C3",X"00",X"03",X"00",X"0C",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"C3",X"33",X"0C",X"33",X"00",X"33",X"00",X"CC",X"00",X"00",X"00",X"00",
		X"33",X"FF",X"33",X"FF",X"33",X"FF",X"33",X"3F",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"F3",X"F0",X"F3",X"FF",X"F3",X"FF",X"33",X"F3",X"33",X"33",X"33",X"30",X"33",X"30",X"33",X"30",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"30",X"00",X"00",X"00",X"00",
		X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"33",X"33",
		X"00",X"00",X"F0",X"00",X"F0",X"00",X"F8",X"00",X"F8",X"00",X"F8",X"00",X"F8",X"00",X"38",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"00",
		X"38",X"00",X"38",X"00",X"38",X"00",X"38",X"00",X"88",X"00",X"88",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"88",X"FF",X"88",X"FF",X"88",X"FF",X"88",X"33",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"88",X"33",X"88",X"33",X"88",X"33",X"88",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"03",X"33",X"03",X"33",X"00",X"88",X"00",X"88",X"00",X"00",X"00",X"FF",X"00",X"88",X"00",X"80",
		X"33",X"33",X"33",X"33",X"88",X"88",X"88",X"88",X"00",X"00",X"FF",X"FF",X"8F",X"8F",X"8F",X"8F",
		X"00",X"80",X"00",X"FF",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"8F",X"8F",X"FF",X"8F",X"88",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"00",X"33",X"00",X"88",X"00",X"88",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"8F",X"8F",X"8F",
		X"33",X"38",X"33",X"38",X"08",X"88",X"08",X"88",X"00",X"00",X"0F",X"0F",X"8F",X"0F",X"8F",X"8F",
		X"8F",X"8F",X"8F",X"0F",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"8F",X"80",X"8F",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"80",X"F8",X"80",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"FF",X"F8",X"F8",X"F8",X"F8",
		X"80",X"F8",X"00",X"FF",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"F8",X"F8",X"F8",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"88",X"88",X"88",X"88",X"00",X"00",X"F0",X"F0",X"F8",X"88",X"F8",X"80",
		X"33",X"33",X"33",X"33",X"88",X"88",X"88",X"88",X"00",X"00",X"F0",X"00",X"88",X"F0",X"F0",X"F8",
		X"F8",X"80",X"F8",X"80",X"08",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"F8",X"F0",X"08",X"88",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F7",X"00",X"AF",X"FA",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"01",X"10",X"FF",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"10",X"00",X"00",X"00",
		X"00",X"F0",X"AF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"55",X"01",X"5F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"10",X"55",X"51",X"55",X"55",
		X"88",X"88",X"88",X"A8",X"88",X"AC",X"88",X"AC",X"88",X"CC",X"8F",X"8F",X"8F",X"CF",X"8F",X"8F",
		X"A8",X"88",X"AC",X"88",X"AC",X"88",X"AC",X"88",X"8C",X"88",X"8F",X"8F",X"C8",X"CF",X"CF",X"CF",
		X"8F",X"8F",X"88",X"88",X"FF",X"8F",X"FC",X"F8",X"8F",X"FF",X"FF",X"FC",X"8C",X"8C",X"88",X"88",
		X"CF",X"8F",X"C8",X"C8",X"F8",X"88",X"FF",X"CF",X"FF",X"CF",X"8F",X"CF",X"88",X"88",X"88",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"55",X"55",X"55",X"AA",X"55",X"A0",X"55",X"00",X"0A",
		X"00",X"00",X"00",X"00",X"06",X"00",X"69",X"66",X"96",X"99",X"69",X"00",X"55",X"30",X"AA",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"A3",X"0A",X"AA",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"55",X"55",X"55",X"AA",X"55",X"A0",X"55",X"00",X"0A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"55",X"00",X"99",X"00",X"69",X"30",X"69",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"96",X"A3",X"96",X"AA",X"69",X"00",X"69",X"00",X"06",X"00",X"06",X"00",X"00",X"00",X"00",X"00",
		X"15",X"F5",X"15",X"55",X"15",X"55",X"15",X"55",X"01",X"55",X"00",X"11",X"00",X"00",X"00",X"11",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"55",X"01",X"55",X"10",X"55",X"51",X"55",X"55",
		X"01",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"01",X"55",X"00",X"55",X"00",X"15",X"00",X"01",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"11",X"11",
		X"10",X"00",X"10",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"00",X"51",X"00",X"51",X"00",X"51",X"00",X"51",X"00",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"00",X"10",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"19",X"00",X"19",X"00",X"99",X"00",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"99",X"00",X"19",X"00",X"19",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"00",X"3F",X"00",X"FF",X"01",X"FF",X"01",X"F3",X"13",X"F3",X"13",X"33",
		X"11",X"11",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"11",X"33",X"00",
		X"13",X"33",X"13",X"33",X"13",X"33",X"13",X"33",X"13",X"33",X"13",X"33",X"13",X"33",X"13",X"33",
		X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"11",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"11",X"00",X"33",X"10",X"33",X"31",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"10",X"00",X"10",X"00",
		X"13",X"33",X"13",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"11",
		X"10",X"00",X"10",X"00",X"10",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"19",X"00",X"FF",X"01",X"99",X"01",X"99",X"19",X"99",X"19",X"99",X"19",X"99",
		X"11",X"00",X"99",X"11",X"99",X"99",X"11",X"99",X"00",X"99",X"00",X"99",X"11",X"99",X"99",X"99",
		X"19",X"99",X"19",X"99",X"19",X"99",X"01",X"99",X"01",X"99",X"00",X"99",X"00",X"19",X"00",X"01",
		X"99",X"11",X"11",X"00",X"00",X"00",X"11",X"11",X"99",X"99",X"99",X"99",X"99",X"91",X"11",X"10",
		X"00",X"10",X"01",X"61",X"16",X"66",X"16",X"66",X"16",X"66",X"16",X"66",X"16",X"66",X"16",X"66",
		X"00",X"00",X"11",X"10",X"F6",X"61",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"16",X"66",
		X"16",X"66",X"16",X"66",X"16",X"66",X"16",X"66",X"16",X"66",X"16",X"66",X"01",X"61",X"00",X"10",
		X"01",X"66",X"01",X"66",X"01",X"66",X"01",X"66",X"01",X"66",X"01",X"66",X"00",X"66",X"00",X"11",
		X"13",X"33",X"13",X"33",X"13",X"33",X"13",X"33",X"13",X"33",X"13",X"33",X"13",X"33",X"13",X"33",
		X"33",X"33",X"33",X"11",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",
		X"13",X"33",X"13",X"33",X"01",X"33",X"01",X"33",X"00",X"33",X"00",X"33",X"00",X"11",X"00",X"00",
		X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"31",X"00",X"10",X"00",X"00",X"00",
		X"33",X"10",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"13",X"00",X"FF",X"01",X"F3",X"01",X"F3",X"13",X"33",X"13",X"33",X"13",X"33",
		X"11",X"00",X"33",X"10",X"33",X"31",X"33",X"33",X"33",X"33",X"13",X"33",X"01",X"33",X"01",X"33",
		X"13",X"33",X"13",X"33",X"01",X"33",X"01",X"33",X"00",X"33",X"00",X"13",X"00",X"13",X"01",X"F3",
		X"13",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"31",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"10",X"01",X"A1",X"1A",X"AA",X"1A",X"AA",X"1A",X"AA",X"1A",X"AA",X"1A",X"AA",X"1A",X"AA",
		X"00",X"11",X"00",X"AA",X"01",X"FA",X"01",X"AA",X"01",X"AA",X"01",X"AA",X"01",X"AA",X"01",X"AA",
		X"1A",X"AA",X"1A",X"AA",X"1A",X"AA",X"1A",X"AA",X"01",X"AA",X"01",X"AA",X"00",X"AA",X"00",X"11",
		X"01",X"AA",X"1A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"11",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",
		X"00",X"01",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"01",X"00",X"00",X"00",X"00",
		X"55",X"00",X"55",X"10",X"55",X"10",X"55",X"10",X"55",X"10",X"55",X"00",X"11",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"13",X"33",X"3F",X"31",X"3F",X"10",X"33",X"10",X"33",X"31",X"33",X"33",X"33",X"33",X"33",X"33",
		X"33",X"33",X"33",X"31",X"13",X"33",X"13",X"33",X"33",X"33",X"33",X"33",X"33",X"31",X"33",X"31",
		X"13",X"33",X"01",X"33",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"10",X"31",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"99",X"19",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"91",
		X"00",X"00",X"10",X"00",X"10",X"00",X"10",X"00",X"10",X"00",X"91",X"10",X"99",X"91",X"99",X"99",
		X"00",X"00",X"00",X"01",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",
		X"11",X"00",X"55",X"00",X"55",X"10",X"55",X"10",X"55",X"10",X"55",X"10",X"55",X"10",X"55",X"10",
		X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"01",X"00",X"00",X"00",X"00",
		X"55",X"10",X"55",X"10",X"55",X"10",X"55",X"10",X"55",X"10",X"55",X"00",X"11",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"01",X"77",X"17",X"77",X"1F",X"77",X"1F",X"77",X"1F",X"77",X"1F",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"17",X"77",X"17",X"77",X"17",X"77",X"17",X"77",X"17",X"77",X"17",X"77",X"17",X"77",X"17",X"77",
		X"00",X"00",X"00",X"01",X"00",X"17",X"00",X"7F",X"00",X"F7",X"01",X"77",X"17",X"77",X"77",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"00",X"77",X"00",X"77",X"00",X"77",X"00",X"77",X"00",X"77",X"00",X"77",X"00",X"71",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"AA",X"01",X"FF",X"01",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"10",X"AA",X"A1",X"AA",X"AA",X"AA",X"AA",
		X"01",X"AA",X"00",X"AA",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"A1",X"11",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"00",X"66",X"00",X"66",X"01",X"66",X"01",X"66",X"01",X"66",X"16",X"66",X"16",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"16",X"66",X"16",X"66",X"01",X"66",X"01",X"66",X"00",X"66",X"00",X"66",X"00",X"16",X"00",X"01",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"61",X"66",X"10",X"66",X"00",X"66",X"00",X"11",X"00",
		X"17",X"77",X"17",X"77",X"17",X"77",X"17",X"77",X"17",X"77",X"17",X"77",X"17",X"77",X"17",X"77",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"17",X"77",X"17",X"77",X"17",X"77",X"17",X"77",X"17",X"77",X"17",X"77",X"01",X"77",X"00",X"11",
		X"77",X"77",X"77",X"77",X"11",X"77",X"00",X"77",X"00",X"77",X"00",X"17",X"00",X"01",X"00",X"00",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"71",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"00",X"77",X"00",X"77",X"00",X"77",X"00",X"77",X"00",X"77",X"00",X"77",X"00",X"11",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"19",X"00",X"01",X"10",X"00",X"91",X"00",X"99",X"00",X"99",X"11",X"99",X"99",
		X"99",X"00",X"91",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"11",X"11",
		X"10",X"00",X"91",X"00",X"91",X"00",X"91",X"00",X"10",X"00",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"11",X"A1",X"AA",X"AA",X"AF",X"AA",X"FA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"17",
		X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"77",X"00",X"77",X"10",X"77",X"10",X"77",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"66",X"00",X"F6",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"11",X"61",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"66",X"10",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"61",X"00",
		X"00",X"01",X"00",X"01",X"00",X"1A",X"00",X"1A",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"A1",X"AA",X"A1",X"AA",X"10",X"AA",X"00",X"AA",X"00",X"AA",X"10",
		X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"1A",X"00",X"01",X"00",X"00",X"00",X"00",
		X"AA",X"A1",X"AA",X"A1",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A1",X"AA",X"11",X"11",X"00",
		X"00",X"17",X"00",X"77",X"00",X"7F",X"00",X"7F",X"00",X"77",X"01",X"77",X"01",X"77",X"17",X"77",
		X"77",X"10",X"77",X"00",X"77",X"00",X"77",X"00",X"71",X"10",X"17",X"71",X"77",X"77",X"77",X"77",
		X"17",X"77",X"17",X"77",X"17",X"77",X"17",X"77",X"17",X"77",X"01",X"77",X"00",X"11",X"00",X"00",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"17",X"77",X"01",X"77",X"00",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"01",X"99",X"19",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"91",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"01",X"77",X"17",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"01",X"77",X"17",X"77",
		X"00",X"F6",X"01",X"66",X"01",X"66",X"01",X"66",X"01",X"66",X"00",X"66",X"00",X"66",X"00",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"00",X"66",X"00",X"16",X"00",X"16",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"11",X"66",X"00",X"11",X"00",X"00",X"00",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"61",X"00",X"61",X"00",X"61",X"00",X"10",X"00",X"10",X"00",X"10",X"00",X"00",X"00",X"00",X"00",
		X"66",X"66",X"66",X"66",X"66",X"61",X"66",X"61",X"66",X"10",X"66",X"00",X"11",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"9F",X"99",X"F9",X"99",X"99",X"99",X"99",X"99",X"91",X"99",X"10",X"99",X"10",X"99",X"91",X"99",
		X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"10",X"99",X"10",X"99",X"10",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"91",X"99",X"10",X"11",X"00",X"00",X"00",
		X"99",X"91",X"99",X"91",X"99",X"99",X"99",X"99",X"99",X"99",X"19",X"91",X"01",X"10",X"00",X"00",
		X"17",X"77",X"17",X"77",X"17",X"77",X"17",X"77",X"17",X"77",X"17",X"77",X"17",X"77",X"17",X"77",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"11",X"77",X"00",X"77",X"00",
		X"17",X"77",X"17",X"77",X"17",X"77",X"17",X"77",X"01",X"77",X"00",X"77",X"00",X"11",X"00",X"00",
		X"71",X"00",X"71",X"00",X"71",X"00",X"10",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"01",X"33",X"13",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"11",X"11",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"11",X"31",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"31",X"00",X"31",X"00",X"31",X"00",X"33",X"11",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"C0",X"CC",X"5C",X"CF",X"CA",X"5C",X"55",X"CF",X"AF",X"A5",X"CF",X"AC",X"FC",X"56",X"C5",
		X"00",X"00",X"F5",X"C0",X"CA",X"CC",X"5A",X"6C",X"A5",X"C6",X"5A",X"C6",X"F5",X"CC",X"AF",X"6C",
		X"FF",X"5F",X"CF",X"C5",X"5C",X"5C",X"AA",X"FF",X"FC",X"CF",X"C5",X"5C",X"CC",X"6C",X"CC",X"CC",
		X"5A",X"FF",X"AF",X"6C",X"4F",X"5C",X"AC",X"65",X"CC",X"A0",X"54",X"5C",X"CA",X"C0",X"55",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CA",X"00",X"CC",X"00",X"5C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"06",X"00",X"55",X"0C",X"A5",X"CC",X"5A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"6C",X"00",X"A0",X"00",X"F5",X"00",X"5C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"FF",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"00",X"FE",X"00",X"FE",X"00",X"EE",X"00",
		X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"FF",X"0E",X"EE",X"00",X"00",
		X"EE",X"00",X"EE",X"00",X"FE",X"00",X"FE",X"00",X"FE",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",
		X"00",X"CF",X"00",X"BF",X"00",X"BF",X"CC",X"FC",X"BB",X"FC",X"CB",X"BF",X"0C",X"FF",X"0C",X"FF",
		X"BB",X"00",X"BB",X"C0",X"BB",X"FC",X"BF",X"FF",X"BF",X"CF",X"FF",X"FF",X"CB",X"FC",X"CC",X"4C",
		X"CB",X"FF",X"CB",X"FF",X"BF",X"FF",X"BF",X"FF",X"BB",X"FF",X"CB",X"B4",X"BB",X"BC",X"CC",X"44",
		X"FF",X"4C",X"BB",X"C0",X"44",X"00",X"CC",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"F5",X"00",X"AA",X"00",X"5A",X"00",X"F5",X"00",X"5A",X"00",X"FA",X"00",X"05",X"00",X"0F",
		X"00",X"00",X"60",X"00",X"60",X"00",X"A0",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"AF",X"00",X"6A",X"00",X"A5",X"00",X"FA",X"00",X"65",X"00",X"A6",X"00",X"0A",X"00",X"00",
		X"A0",X"00",X"A5",X"00",X"5F",X"00",X"5A",X"00",X"5F",X"00",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"65",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"55",X"00",X"5A",X"00",X"FA",X"00",X"FA",X"00",X"65",X"00",X"A6",X"00",X"AA",X"00",X"0A",
		X"A0",X"00",X"6A",X"00",X"55",X"00",X"55",X"00",X"56",X"00",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5F",X"00",X"16",X"0A",X"5F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"55",X"00",
		X"05",X"F5",X"05",X"F5",X"0A",X"5F",X"00",X"AF",X"00",X"65",X"00",X"5A",X"00",X"0A",X"00",X"00",
		X"F6",X"00",X"AF",X"00",X"6A",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"FA",X"00",X"A6",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FA",X"00",X"6A",X"00",
		X"06",X"A5",X"06",X"AA",X"0F",X"AA",X"0F",X"55",X"00",X"FF",X"00",X"55",X"00",X"AA",X"00",X"0A",
		X"65",X"00",X"F5",X"00",X"F5",X"00",X"A5",X"00",X"A5",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"66",X"00",X"6A",X"00",X"5F",X"0A",X"F6",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"AA",X"00",
		X"0A",X"FF",X"55",X"6A",X"65",X"F5",X"A6",X"55",X"A6",X"FF",X"0A",X"65",X"05",X"5F",X"00",X"FA",
		X"6A",X"00",X"55",X"00",X"F5",X"00",X"F5",X"00",X"A5",X"00",X"5A",X"00",X"6A",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"6A",X"00",X"66",X"06",X"1F",X"05",X"AF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A5",X"00",X"F6",X"00",X"5F",X"00",
		X"A5",X"AA",X"A5",X"5A",X"A5",X"AA",X"6A",X"55",X"06",X"6A",X"06",X"A6",X"00",X"A5",X"00",X"55",
		X"A6",X"00",X"AA",X"00",X"55",X"00",X"F5",X"00",X"F5",X"00",X"5A",X"00",X"A5",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0A",X"00",X"AA",X"00",X"5A",X"00",X"16",X"05",X"65",X"55",X"6F",X"6A",X"FA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"FF",X"00",X"AA",X"00",X"FF",X"00",
		X"5F",X"A6",X"F1",X"6F",X"5F",X"FA",X"A6",X"5F",X"56",X"AF",X"AA",X"F5",X"05",X"A5",X"00",X"55",
		X"6A",X"00",X"F5",X"00",X"5F",X"00",X"5F",X"00",X"F6",X"00",X"FA",X"00",X"FA",X"00",X"00",X"00",
		X"00",X"0A",X"00",X"0A",X"00",X"66",X"00",X"F6",X"00",X"15",X"0A",X"1F",X"A5",X"5F",X"A5",X"5A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"6A",X"00",X"56",X"00",X"56",X"00",X"5A",X"00",
		X"66",X"55",X"56",X"5A",X"A5",X"AA",X"AA",X"A6",X"6A",X"6F",X"06",X"65",X"00",X"A5",X"00",X"66",
		X"F6",X"60",X"AA",X"50",X"F5",X"50",X"F6",X"00",X"56",X"00",X"FA",X"00",X"AA",X"00",X"00",X"00",
		X"00",X"0A",X"00",X"A5",X"00",X"FF",X"0A",X"55",X"AF",X"55",X"AF",X"66",X"AF",X"AA",X"AA",X"6A",
		X"00",X"00",X"00",X"00",X"A0",X"00",X"FA",X"00",X"65",X"00",X"A5",X"00",X"6A",X"00",X"55",X"A0",
		X"5A",X"AA",X"55",X"AA",X"F5",X"6A",X"6F",X"AA",X"66",X"AA",X"A5",X"55",X"0A",X"5A",X"00",X"AA",
		X"A5",X"A0",X"A5",X"50",X"A5",X"50",X"A6",X"00",X"A6",X"00",X"56",X"00",X"66",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"05",X"01",X"00",X"11",X"00",X"1F",X"00",X"FE",
		X"00",X"00",X"00",X"00",X"11",X"00",X"1F",X"11",X"EE",X"E1",X"EF",X"EE",X"EE",X"0E",X"EE",X"00",
		X"00",X"11",X"00",X"1E",X"00",X"EF",X"00",X"1E",X"00",X"EF",X"00",X"1E",X"50",X"F1",X"00",X"1F",
		X"EE",X"00",X"EE",X"00",X"E0",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"E0",X"00",X"EE",X"00",
		X"00",X"11",X"00",X"1F",X"01",X"FE",X"11",X"EF",X"1F",X"EE",X"1F",X"EE",X"FE",X"EE",X"E1",X"EE",
		X"1F",X"00",X"EE",X"10",X"EE",X"EF",X"EE",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"EE",X"1F",X"E0",X"EF",X"E0",X"FE",X"00",X"EF",X"E0",X"FF",X"E0",X"1E",X"E0",X"11",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"50",X"00",X"00",X"00",X"01",X"50",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"11",X"10",X"FF",X"EF",
		X"00",X"1E",X"00",X"FF",X"01",X"EE",X"01",X"FE",X"01",X"EE",X"01",X"EE",X"00",X"EE",X"00",X"0E",
		X"EE",X"EE",X"E0",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"11",X"01",X"F1",X"11",X"E1",X"11",X"EF",X"11",X"EE",X"1E",X"EE",X"EE",X"EE",
		X"11",X"00",X"1E",X"10",X"EE",X"11",X"EF",X"F1",X"EE",X"EF",X"EE",X"EE",X"EE",X"EE",X"00",X"0E",
		X"1F",X"EE",X"EE",X"E0",X"FE",X"00",X"EE",X"00",X"FE",X"00",X"EE",X"00",X"EE",X"00",X"0E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",
		X"00",X"00",X"00",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"11",X"E0",
		X"00",X"50",X"00",X"0E",X"00",X"01",X"00",X"E1",X"00",X"11",X"00",X"01",X"55",X"01",X"00",X"00",
		X"1E",X"EE",X"EE",X"E0",X"FE",X"00",X"EE",X"00",X"EE",X"00",X"E0",X"00",X"E0",X"00",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"50",X"11",X"05",X"11",X"00",X"1E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"E1",X"00",X"FF",X"00",X"FE",X"00",X"EE",X"00",
		X"00",X"1F",X"00",X"EF",X"00",X"FE",X"00",X"FE",X"00",X"EE",X"00",X"FE",X"50",X"EE",X"00",X"FE",
		X"E0",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"10",X"11",X"11",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"11",X"00",X"11",X"00",X"0E",X"00",X"00",
		X"1E",X"EE",X"E1",X"FE",X"EF",X"EE",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"E0",X"00",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"11",X"00",X"1E",
		X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"00",X"11",X"00",X"11",X"11",X"FF",X"EF",X"EE",X"EE",
		X"50",X"FF",X"01",X"EE",X"01",X"FE",X"01",X"EE",X"01",X"EE",X"00",X"EE",X"01",X"E0",X"00",X"E0",
		X"EE",X"E0",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"0F",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"AA",X"00",X"FA",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CF",X"FF",X"00",X"CC",
		X"FA",X"C0",X"FF",X"C0",X"FF",X"AC",X"FF",X"AC",X"FA",X"AC",X"AA",X"C0",X"AA",X"00",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"AC",X"FF",X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"AC",X"00",X"AC",X"00",
		X"FF",X"FF",X"0F",X"FF",X"0F",X"FF",X"00",X"FF",X"00",X"FF",X"0F",X"FF",X"00",X"FF",X"00",X"CC",
		X"AC",X"00",X"AC",X"00",X"FA",X"00",X"FF",X"C0",X"FF",X"AC",X"FF",X"AC",X"AA",X"C0",X"CC",X"00",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"FF",X"AC",
		X"00",X"00",X"FC",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"C0",X"FF",X"C0",X"AF",X"FC",X"AA",X"FC",
		X"AA",X"C0",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"AC",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"00",X"FF",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"FF",X"00",X"FA",X"00",X"AC",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FA",X"FF",X"FA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AC",X"AA",X"C0",X"CC",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"03",X"33",X"3F",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"22",X"00",X"32",X"00",
		X"FF",X"33",X"F3",X"33",X"33",X"33",X"33",X"33",X"33",X"22",X"33",X"CC",X"32",X"00",X"CC",X"00",
		X"33",X"C0",X"33",X"C0",X"33",X"2C",X"33",X"2C",X"33",X"2C",X"33",X"2C",X"33",X"C0",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"9F",X"00",X"FF",X"00",X"F9",X"00",X"99",X"09",X"99",X"09",X"99",
		X"00",X"00",X"88",X"00",X"98",X"00",X"99",X"00",X"99",X"C0",X"99",X"C0",X"99",X"C0",X"98",X"00",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"C9",X"99",X"0C",X"CC",
		X"88",X"00",X"88",X"00",X"8C",X"00",X"C0",X"00",X"8C",X"00",X"8C",X"00",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"66",X"00",X"FF",X"00",X"F6",X"00",X"F6",X"00",X"66",X"00",X"66",X"00",X"66",
		X"00",X"00",X"C0",X"00",X"5C",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"65",X"00",X"65",X"00",
		X"00",X"66",X"00",X"66",X"00",X"66",X"00",X"66",X"00",X"66",X"00",X"66",X"00",X"66",X"00",X"CC",
		X"65",X"00",X"65",X"00",X"65",X"00",X"65",X"00",X"65",X"00",X"65",X"00",X"55",X"00",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"0A",X"AC",X"AF",X"AA",X"FF",X"AA",X"FF",X"AA",X"FA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BC",X"00",X"BB",X"00",X"AB",X"00",X"AB",X"00",
		X"AA",X"AA",X"0A",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"CC",
		X"AA",X"C0",X"AA",X"C0",X"AA",X"C0",X"AA",X"C0",X"AA",X"C0",X"AA",X"C0",X"AB",X"00",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"FF",X"00",X"F7",X"00",X"77",X"00",X"77",X"00",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"3C",X"00",X"3C",X"00",X"3C",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"77",X"00",X"F7",X"00",X"17",X"00",X"77",X"00",X"77",X"00",X"73",X"00",X"33",
		X"00",X"00",X"00",X"00",X"C0",X"00",X"3C",X"00",X"3C",X"00",X"3C",X"00",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"77",X"00",X"F1",X"00",X"17",X"00",X"17",X"00",X"77",X"00",X"77",X"00",X"77",X"00",X"33",
		X"C0",X"00",X"3C",X"00",X"73",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"3C",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",
		X"00",X"17",X"07",X"77",X"07",X"77",X"07",X"77",X"07",X"77",X"07",X"77",X"00",X"73",X"00",X"33",
		X"3C",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"3C",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"F1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"73",X"00",
		X"00",X"11",X"07",X"17",X"07",X"77",X"07",X"77",X"07",X"77",X"00",X"77",X"00",X"33",X"00",X"33",
		X"73",X"00",X"73",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"07",X"77",X"0F",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"73",X"00",X"73",X"00",
		X"7F",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"07",X"73",X"03",X"33",X"00",X"33",
		X"73",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"F7",X"07",X"17",X"07",X"17",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"73",X"00",X"77",X"00",X"77",X"00",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"07",X"77",X"07",X"77",X"00",X"33",X"00",X"33",
		X"77",X"C0",X"77",X"C0",X"73",X"C0",X"73",X"C0",X"33",X"00",X"33",X"00",X"33",X"00",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"07",X"77",X"77",X"77",X"7F",X"77",X"FF",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"33",X"00",X"73",X"00",X"73",X"00",X"73",X"C0",
		X"F1",X"77",X"71",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"73",X"07",X"33",X"00",X"33",
		X"73",X"C0",X"33",X"C0",X"33",X"C0",X"33",X"C0",X"33",X"00",X"33",X"00",X"33",X"00",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"17",X"07",X"77",X"7F",X"77",X"7F",X"77",X"71",X"77",
		X"00",X"00",X"00",X"00",X"C0",X"00",X"73",X"00",X"77",X"00",X"77",X"C0",X"77",X"C0",X"77",X"3C",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"07",X"73",X"00",X"33",X"00",X"33",
		X"77",X"3C",X"73",X"3C",X"73",X"3C",X"33",X"C0",X"33",X"C0",X"33",X"00",X"33",X"00",X"CC",X"00",
		X"00",X"00",X"00",X"77",X"07",X"77",X"7F",X"77",X"FF",X"77",X"FF",X"77",X"F1",X"77",X"17",X"77",
		X"00",X"00",X"C0",X"00",X"33",X"00",X"73",X"00",X"73",X"C0",X"73",X"C0",X"73",X"3C",X"73",X"3C",
		X"17",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"33",X"33",X"33",X"03",X"33",X"00",X"33",
		X"33",X"3C",X"33",X"3C",X"33",X"3C",X"33",X"C0",X"33",X"C0",X"33",X"00",X"33",X"00",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"3F",X"03",X"3F",X"33",X"3F",X"33",X"3F",
		X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"BB",X"3F",X"BB",X"CF",
		X"33",X"33",X"33",X"33",X"33",X"3B",X"3F",X"FB",X"FF",X"FB",X"FF",X"FB",X"FF",X"FB",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"33",X"00",X"FF",X"3C",X"CF",X"33",X"FF",X"33",X"FF",X"33",X"FF",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"3C",X"00",X"32",X"00",
		X"FF",X"33",X"33",X"33",X"BB",X"33",X"CC",X"33",X"CC",X"33",X"CC",X"33",X"BC",X"33",X"BC",X"33",
		X"FF",X"C0",X"FC",X"FC",X"FC",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"C0",X"22",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"FF",X"00",X"F7",X"00",X"77",X"00",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"3C",X"00",X"3C",X"00",X"3C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"FF",X"00",X"F7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"3C",X"00",
		X"BB",X"BC",X"BB",X"BC",X"BB",X"CF",X"BB",X"FF",X"BB",X"FF",X"C2",X"FF",X"02",X"FF",X"02",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"02",X"FF",X"02",X"2F",X"02",X"22",X"02",X"22",X"0C",X"22",X"00",X"CC",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"BC",X"FF",X"BB",X"FF",X"BB",X"2B",X"BB",X"CB",X"BB",X"0C",X"BB",X"00",X"CC",
		X"BB",X"33",X"FF",X"33",X"FF",X"33",X"FF",X"33",X"FF",X"32",X"FF",X"32",X"FF",X"22",X"FF",X"22",
		X"22",X"00",X"22",X"00",X"22",X"00",X"2C",X"00",X"22",X"2C",X"22",X"C0",X"2C",X"00",X"C0",X"00",
		X"F3",X"2C",X"32",X"C0",X"22",X"00",X"22",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"09",X"00",X"99",X"00",X"98",X"00",X"89",
		X"00",X"00",X"9C",X"00",X"C9",X"00",X"99",X"99",X"98",X"88",X"88",X"88",X"88",X"44",X"44",X"11",
		X"09",X"88",X"09",X"84",X"09",X"44",X"99",X"41",X"99",X"41",X"99",X"41",X"99",X"11",X"98",X"11",
		X"11",X"11",X"11",X"BB",X"1B",X"44",X"B4",X"11",X"41",X"1B",X"41",X"B4",X"11",X"4C",X"11",X"CC",
		X"00",X"00",X"98",X"00",X"CC",X"00",X"99",X"89",X"99",X"88",X"88",X"98",X"88",X"98",X"48",X"99",
		X"00",X"00",X"00",X"00",X"9C",X"00",X"F9",X"00",X"F8",X"00",X"88",X"00",X"98",X"00",X"88",X"00",
		X"14",X"89",X"11",X"88",X"44",X"48",X"11",X"48",X"11",X"14",X"41",X"14",X"C4",X"14",X"C4",X"14",
		X"88",X"00",X"88",X"00",X"88",X"00",X"88",X"C0",X"88",X"C0",X"88",X"C0",X"88",X"C0",X"88",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"09",X"00",X"99",X"00",X"98",X"00",X"89",
		X"00",X"00",X"9C",X"00",X"C9",X"00",X"99",X"99",X"98",X"88",X"88",X"88",X"88",X"44",X"44",X"11",
		X"09",X"88",X"09",X"84",X"09",X"44",X"99",X"41",X"99",X"41",X"99",X"41",X"99",X"11",X"98",X"11",
		X"11",X"11",X"11",X"BB",X"1B",X"44",X"B4",X"11",X"41",X"1B",X"41",X"B4",X"11",X"4C",X"11",X"CC",
		X"00",X"00",X"98",X"00",X"CC",X"00",X"99",X"89",X"99",X"88",X"88",X"98",X"88",X"98",X"48",X"99",
		X"00",X"00",X"00",X"00",X"9C",X"00",X"F9",X"00",X"F8",X"00",X"88",X"00",X"98",X"00",X"88",X"00",
		X"14",X"89",X"11",X"88",X"44",X"48",X"11",X"48",X"11",X"14",X"41",X"14",X"C4",X"14",X"C4",X"14",
		X"88",X"00",X"88",X"00",X"88",X"00",X"88",X"C0",X"88",X"C0",X"88",X"C0",X"88",X"C0",X"88",X"C0",
		X"98",X"1B",X"98",X"1B",X"98",X"11",X"98",X"44",X"88",X"8C",X"C8",X"8C",X"08",X"C5",X"09",X"C5",
		X"11",X"CC",X"11",X"CC",X"55",X"CC",X"55",X"C5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"99",X"C5",X"99",X"55",X"99",X"55",X"88",X"C5",X"CC",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"41",X"CC",X"41",X"5C",X"14",X"55",X"88",X"5C",X"88",X"5C",X"FF",X"CF",X"FF",X"CF",X"CC",
		X"88",X"8C",X"88",X"8C",X"88",X"88",X"88",X"88",X"CC",X"88",X"99",X"88",X"98",X"88",X"88",X"88",
		X"FF",X"98",X"CC",X"89",X"00",X"89",X"00",X"89",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"8C",X"89",X"8C",X"98",X"C0",X"98",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"98",X"1B",X"98",X"1B",X"98",X"11",X"98",X"44",X"88",X"85",X"C8",X"55",X"08",X"55",X"09",X"C5",
		X"11",X"CC",X"11",X"CC",X"CC",X"CC",X"55",X"CC",X"55",X"CC",X"55",X"5C",X"55",X"55",X"55",X"55",
		X"99",X"8C",X"99",X"8C",X"99",X"8C",X"88",X"C0",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"CC",X"FF",X"FF",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"41",X"CC",X"41",X"CC",X"14",X"55",X"88",X"5C",X"88",X"CF",X"FF",X"CF",X"FF",X"FF",X"CC",
		X"88",X"8C",X"88",X"8C",X"88",X"88",X"88",X"88",X"CC",X"88",X"99",X"88",X"98",X"88",X"88",X"88",
		X"FF",X"98",X"FC",X"89",X"C0",X"89",X"00",X"89",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"8C",X"89",X"8C",X"98",X"C0",X"98",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"09",X"00",X"99",X"00",X"98",X"00",X"89",
		X"00",X"00",X"8C",X"00",X"C8",X"00",X"99",X"99",X"98",X"88",X"88",X"88",X"88",X"88",X"88",X"44",
		X"09",X"88",X"09",X"88",X"09",X"84",X"99",X"84",X"99",X"45",X"99",X"55",X"99",X"C5",X"9D",X"FC",
		X"44",X"BB",X"BB",X"11",X"14",X"44",X"4B",X"BB",X"55",X"C1",X"55",X"5C",X"5C",X"CD",X"CF",X"FF",
		X"00",X"00",X"98",X"00",X"CC",X"00",X"99",X"89",X"99",X"88",X"88",X"98",X"88",X"98",X"88",X"99",
		X"00",X"00",X"00",X"00",X"9C",X"00",X"F9",X"00",X"F8",X"00",X"88",X"00",X"98",X"00",X"88",X"00",
		X"88",X"89",X"44",X"88",X"BB",X"88",X"44",X"88",X"BB",X"48",X"1B",X"48",X"11",X"B4",X"D1",X"B4",
		X"88",X"00",X"88",X"00",X"88",X"00",X"88",X"C0",X"88",X"C0",X"88",X"C0",X"88",X"C0",X"88",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"99",X"00",X"99",X"00",X"98",X"00",X"89",
		X"00",X"00",X"9C",X"00",X"C9",X"00",X"99",X"99",X"98",X"88",X"88",X"88",X"88",X"88",X"88",X"FF",
		X"09",X"88",X"09",X"88",X"09",X"8F",X"99",X"8F",X"99",X"FF",X"99",X"FF",X"99",X"FF",X"98",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"98",X"00",X"CC",X"00",X"99",X"89",X"99",X"88",X"88",X"98",X"88",X"98",X"88",X"99",
		X"00",X"00",X"00",X"00",X"9C",X"00",X"F9",X"00",X"F8",X"00",X"88",X"00",X"98",X"00",X"88",X"00",
		X"88",X"89",X"FF",X"88",X"FF",X"88",X"FF",X"88",X"FF",X"E8",X"FF",X"F8",X"FF",X"FE",X"FF",X"FF",
		X"88",X"00",X"88",X"00",X"88",X"00",X"88",X"C0",X"88",X"C0",X"88",X"C0",X"88",X"C0",X"88",X"C0",
		X"9D",X"FF",X"9F",X"FF",X"9F",X"FF",X"9F",X"FF",X"88",X"FF",X"C8",X"FF",X"08",X"FF",X"09",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"99",X"8F",X"99",X"88",X"99",X"88",X"88",X"8C",X"CC",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"ED",X"1B",X"FF",X"D1",X"FF",X"ED",X"FF",X"FE",X"FF",X"FE",X"FF",X"EE",X"FF",X"EE",X"FF",X"CC",
		X"88",X"8C",X"88",X"8C",X"88",X"88",X"88",X"88",X"CC",X"88",X"99",X"88",X"98",X"88",X"88",X"88",
		X"FE",X"98",X"EE",X"89",X"CC",X"89",X"00",X"89",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"8C",X"89",X"8C",X"98",X"C0",X"98",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"98",X"FF",X"98",X"FF",X"98",X"FF",X"98",X"FF",X"88",X"FF",X"C8",X"FF",X"08",X"8F",X"09",X"8F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"99",X"88",X"99",X"88",X"99",X"88",X"88",X"8C",X"CC",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FE",X"FF",X"EE",X"FF",X"EE",X"FF",X"CC",
		X"88",X"8C",X"88",X"8C",X"88",X"88",X"88",X"88",X"CC",X"88",X"99",X"88",X"98",X"88",X"88",X"88",
		X"FE",X"98",X"EE",X"89",X"CC",X"89",X"00",X"89",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"8C",X"89",X"8C",X"98",X"C0",X"98",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"9C",X"99",X"99",X"44",X"4B",X"CC",X"BC",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"80",X"99",X"98",X"44",X"89",X"BB",X"BB",X"41",X"1B",
		X"1C",X"55",X"1C",X"CC",X"CF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C4",X"11",X"CC",X"11",X"EE",X"C1",X"FF",X"EC",X"FF",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"8C",X"C0",X"9C",X"F8",X"88",X"88",X"88",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"48",X"88",X"B4",X"88",X"1B",X"88",X"11",X"88",X"CC",X"88",X"EE",X"88",X"EE",X"48",X"FE",X"C8",
		X"C0",X"00",X"C0",X"00",X"9C",X"00",X"9C",X"00",X"9C",X"00",X"89",X"00",X"89",X"00",X"88",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"98",X"00",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"98",X"88",X"99",X"98",X"99",X"99",
		X"0F",X"99",X"0F",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"00",X"00",X"00",X"00",X"CC",X"00",X"88",X"CC",X"88",X"88",X"89",X"88",X"89",X"88",X"99",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"8C",X"00",X"88",X"00",
		X"99",X"F8",X"99",X"FF",X"99",X"FF",X"99",X"98",X"99",X"98",X"99",X"88",X"99",X"88",X"99",X"88",
		X"88",X"00",X"88",X"C0",X"88",X"C0",X"88",X"8C",X"88",X"8C",X"88",X"8C",X"88",X"8C",X"C8",X"8C",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CF",X"FF",X"0F",X"FF",X"0C",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"FF",X"00",X"99",X"00",X"98",X"00",X"88",X"00",X"88",X"09",X"88",X"99",X"88",X"98",X"8C",
		X"FF",X"FF",X"FF",X"FF",X"CE",X"EE",X"0C",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"E9",X"FE",X"E9",X"FE",X"99",X"FE",X"98",X"FE",X"88",X"FF",X"E8",X"FF",X"EE",X"FF",X"EE",
		X"88",X"C0",X"88",X"8C",X"88",X"8C",X"88",X"8C",X"88",X"8C",X"88",X"8C",X"88",X"C0",X"88",X"C0",
		X"EE",X"EC",X"EE",X"C0",X"EC",X"09",X"C0",X"09",X"00",X"99",X"00",X"98",X"00",X"98",X"00",X"8C",
		X"88",X"00",X"88",X"00",X"88",X"00",X"88",X"00",X"88",X"00",X"8C",X"00",X"8C",X"00",X"88",X"00",
		X"98",X"99",X"9C",X"99",X"99",X"99",X"89",X"88",X"11",X"55",X"11",X"55",X"44",X"55",X"FC",X"55",
		X"99",X"99",X"99",X"99",X"99",X"88",X"88",X"C1",X"55",X"11",X"55",X"14",X"5C",X"4C",X"CC",X"CF",
		X"CF",X"CC",X"99",X"FF",X"99",X"FF",X"99",X"88",X"98",X"88",X"98",X"88",X"88",X"8C",X"CC",X"C0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"8C",X"81",X"C9",X"11",X"C9",X"11",X"C9",X"1C",X"C9",X"CF",X"C9",X"FF",X"C8",X"FF",X"FC",
		X"88",X"8C",X"88",X"8C",X"88",X"C0",X"88",X"C0",X"88",X"00",X"88",X"00",X"88",X"C0",X"88",X"8C",
		X"FF",X"FC",X"FF",X"C0",X"FF",X"00",X"CC",X"00",X"00",X"08",X"00",X"88",X"00",X"88",X"00",X"88",
		X"88",X"8C",X"88",X"8C",X"88",X"8C",X"88",X"C0",X"88",X"C0",X"88",X"00",X"88",X"00",X"88",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"FB",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"BB",X"00",X"BB",X"C0",X"BB",X"C0",X"FB",X"C0",X"FF",X"C0",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BC",X"00",X"BB",X"00",
		X"FF",X"33",X"F3",X"33",X"33",X"3C",X"33",X"CF",X"33",X"33",X"33",X"FF",X"33",X"FF",X"33",X"FC",
		X"BB",X"00",X"BB",X"00",X"FB",X"00",X"BC",X"00",X"BB",X"00",X"CC",X"00",X"BB",X"C0",X"BB",X"00",
		X"00",X"00",X"FF",X"F0",X"FF",X"F0",X"FF",X"F8",X"FF",X"F8",X"FF",X"F8",X"FF",X"F8",X"33",X"38",
		X"00",X"00",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"33",
		X"33",X"38",X"33",X"38",X"33",X"38",X"33",X"38",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"0F",X"00",X"0F",X"88",X"0F",X"88",X"0F",X"88",X"0F",X"88",X"0F",X"88",X"03",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"33",X"33",
		X"88",X"03",X"88",X"03",X"88",X"03",X"88",X"03",X"88",X"03",X"88",X"03",X"88",X"03",X"88",X"03",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"88",X"33",X"88",X"33",X"80",X"33",X"80",
		X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"C3",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"CC",X"33",X"00",X"C3",X"00",X"0C",X"00",X"00",
		X"33",X"FF",X"33",X"FF",X"33",X"FF",X"33",X"FF",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"3F",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"00",X"00",X"00",X"00",X"00",
		X"33",X"00",X"33",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"33",X"33",
		X"00",X"00",X"00",X"FF",X"00",X"FF",X"80",X"FF",X"80",X"FF",X"80",X"FF",X"80",X"FF",X"80",X"33",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"00",
		X"80",X"33",X"80",X"33",X"80",X"33",X"80",X"33",X"80",X"33",X"80",X"33",X"00",X"33",X"00",X"33",
		X"00",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"33",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"33",X"00",X"33",X"88",X"33",X"88",
		X"33",X"33",X"33",X"33",X"08",X"88",X"08",X"88",X"00",X"00",X"0F",X"0F",X"0F",X"8F",X"0F",X"0F",
		X"33",X"33",X"33",X"33",X"88",X"88",X"88",X"88",X"00",X"00",X"0F",X"F0",X"8F",X"8F",X"8F",X"8F",
		X"0F",X"0F",X"0F",X"0F",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"8F",X"8F",X"8F",X"8F",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"03",X"88",X"03",X"88",X"00",X"88",X"00",X"00",X"00",X"FF",X"FF",X"8F",X"8F",X"FF",X"FF",
		X"33",X"80",X"33",X"80",X"88",X"80",X"88",X"80",X"00",X"00",X"F0",X"0F",X"8F",X"8F",X"8F",X"FF",
		X"88",X"8F",X"80",X"8F",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"8F",X"F8",X"8F",X"F8",X"80",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"33",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"F0",X"F8",X"F8",X"F8",X"F8",
		X"00",X"00",X"00",X"F0",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"F8",X"F8",X"F8",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"88",X"88",X"88",X"88",X"00",X"00",X"FF",X"FF",X"0F",X"F8",X"0F",X"FF",
		X"33",X"88",X"33",X"88",X"88",X"88",X"88",X"88",X"00",X"00",X"FF",X"00",X"F8",X"00",X"F8",X"00",
		X"0F",X"F8",X"0F",X"FF",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"00",X"FF",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"FA",X"7F",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"01",X"00",X"11",X"11",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"01",X"00",X"10",X"00",X"00",X"00",
		X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"55",X"10",X"55",X"51",
		X"A8",X"A8",X"AA",X"AC",X"AC",X"AA",X"AA",X"8C",X"8C",X"88",X"FF",X"8F",X"CC",X"CF",X"F8",X"CF",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"FF",X"88",X"CF",X"C8",X"F8",X"C8",
		X"CC",X"FF",X"C8",X"CC",X"F8",X"88",X"CC",X"F8",X"F8",X"FC",X"FC",X"FC",X"CC",X"8C",X"88",X"88",
		X"FF",X"C8",X"CC",X"C8",X"8F",X"F8",X"FF",X"8F",X"FF",X"FF",X"FC",X"CF",X"CC",X"C8",X"88",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"56",X"F5",X"56",X"55",X"99",X"00",X"65",X"00",X"AA",
		X"00",X"00",X"00",X"00",X"66",X"00",X"66",X"00",X"69",X"66",X"99",X"00",X"23",X"00",X"A5",X"00",
		X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"30",X"AA",X"30",X"B0",X"33",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"F5",X"55",X"55",X"55",X"00",X"99",X"00",X"69",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"93",X"00",X"23",X"00",X"95",X"00",
		X"00",X"A6",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"9A",X"30",X"69",X"30",X"69",X"33",X"69",X"03",X"99",X"03",X"66",X"03",X"66",X"03",X"00",X"03",
		X"5F",X"55",X"5F",X"55",X"55",X"55",X"55",X"55",X"15",X"55",X"01",X"55",X"00",X"15",X"11",X"01",
		X"55",X"55",X"55",X"55",X"55",X"55",X"51",X"51",X"51",X"10",X"55",X"00",X"55",X"10",X"55",X"51",
		X"55",X"11",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"55",X"01",X"55",X"00",X"11",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"11",X"11",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"19",X"00",X"99",X"00",X"9F",X"00",X"99",X"00",X"99",X"01",X"99",X"01",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"99",X"01",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"11",X"00",X"00",X"00",X"00",
		X"00",X"11",X"00",X"33",X"01",X"F3",X"13",X"F3",X"3F",X"33",X"3F",X"33",X"3F",X"33",X"33",X"33",
		X"11",X"11",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"13",X"31",X"01",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"10",X"00",X"10",X"00",X"31",X"01",X"33",X"13",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"10",X"00",X"31",X"00",X"33",X"10",X"33",X"31",X"33",X"31",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"31",X"33",X"31",X"33",X"10",X"33",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"01",X"99",X"19",X"99",X"9F",X"91",X"FF",X"10",X"FF",X"10",X"9F",X"91",X"99",X"99",
		X"11",X"00",X"99",X"00",X"99",X"10",X"99",X"10",X"19",X"91",X"19",X"91",X"99",X"91",X"99",X"10",
		X"99",X"99",X"99",X"91",X"99",X"10",X"99",X"91",X"99",X"99",X"19",X"99",X"01",X"99",X"00",X"11",
		X"99",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"99",X"10",X"99",X"10",X"99",X"00",X"11",X"00",
		X"11",X"00",X"66",X"01",X"FF",X"16",X"F6",X"6F",X"F6",X"66",X"F6",X"66",X"66",X"66",X"66",X"61",
		X"00",X"00",X"11",X"00",X"66",X"00",X"66",X"10",X"66",X"61",X"66",X"61",X"66",X"61",X"66",X"61",
		X"66",X"10",X"66",X"10",X"66",X"10",X"66",X"10",X"66",X"10",X"66",X"10",X"66",X"00",X"11",X"00",
		X"66",X"61",X"66",X"61",X"66",X"61",X"66",X"61",X"66",X"61",X"66",X"61",X"16",X"10",X"01",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"33",X"33",X"33",X"11",X"31",X"00",X"10",X"00",X"10",X"00",X"10",X"00",X"31",X"00",X"31",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"13",X"33",X"01",X"33",X"00",X"11",X"00",X"00",
		X"31",X"00",X"31",X"00",X"31",X"00",X"31",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"01",X"FF",X"13",X"33",X"3F",X"33",X"3F",X"33",X"33",X"31",X"33",X"10",X"33",X"10",
		X"10",X"00",X"31",X"00",X"33",X"00",X"33",X"10",X"33",X"10",X"33",X"31",X"33",X"31",X"33",X"31",
		X"33",X"31",X"33",X"33",X"33",X"33",X"33",X"33",X"13",X"33",X"01",X"33",X"01",X"33",X"13",X"33",
		X"33",X"31",X"33",X"31",X"33",X"31",X"33",X"10",X"33",X"10",X"33",X"31",X"33",X"31",X"33",X"31",
		X"11",X"00",X"AA",X"00",X"FF",X"10",X"FA",X"10",X"FA",X"10",X"AA",X"10",X"AA",X"10",X"AA",X"10",
		X"01",X"00",X"1A",X"10",X"AF",X"A1",X"AF",X"A1",X"AF",X"A1",X"AA",X"A1",X"AA",X"A1",X"AA",X"A1",
		X"AA",X"10",X"AA",X"A1",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"11",X"AA",X"00",X"11",
		X"AA",X"A1",X"AA",X"A1",X"AA",X"A1",X"AA",X"A1",X"AA",X"A1",X"AA",X"A1",X"1A",X"A1",X"01",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",
		X"00",X"55",X"00",X"FF",X"00",X"F5",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"11",X"00",X"00",
		X"51",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"51",X"00",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"13",X"00",X"13",X"00",X"13",X"00",X"13",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"33",X"F3",X"11",X"33",X"00",X"33",X"00",X"33",X"11",X"33",X"33",X"33",X"33",X"33",X"33",
		X"33",X"10",X"33",X"00",X"33",X"10",X"33",X"10",X"33",X"10",X"33",X"10",X"33",X"00",X"33",X"00",
		X"33",X"33",X"13",X"33",X"01",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"19",X"91",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"91",X"99",X"19",X"99",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"99",X"00",X"99",X"10",
		X"00",X"11",X"00",X"55",X"00",X"FF",X"00",X"F5",X"00",X"F5",X"00",X"55",X"00",X"55",X"00",X"55",
		X"10",X"00",X"51",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",
		X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"11",X"00",X"00",
		X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"51",X"00",X"10",X"00",X"00",X"00",
		X"00",X"00",X"11",X"00",X"77",X"10",X"FF",X"71",X"F7",X"71",X"77",X"71",X"77",X"71",X"77",X"71",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"71",X"77",X"71",X"77",X"71",X"77",X"71",X"77",X"71",X"77",X"71",X"77",X"77",X"77",X"77",
		X"00",X"01",X"00",X"17",X"00",X"FF",X"01",X"77",X"17",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"00",X"71",X"00",X"71",X"00",X"71",X"00",X"71",X"00",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"11",X"1A",X"AA",X"AA",X"FA",X"AF",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"AA",X"00",X"AA",X"10",X"AA",X"10",
		X"AA",X"AA",X"1A",X"AA",X"01",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"10",X"AA",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"16",X"66",X"16",X"66",X"16",X"66",X"16",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"16",X"66",X"16",X"66",X"01",X"66",X"00",X"11",
		X"66",X"66",X"66",X"61",X"66",X"10",X"66",X"00",X"66",X"00",X"61",X"00",X"10",X"00",X"00",X"00",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"77",X"77",X"77",X"71",X"77",X"10",X"77",X"10",X"77",X"10",X"77",X"71",X"77",X"77",X"77",X"77",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"71",X"77",X"71",X"77",X"71",X"77",X"10",X"11",X"00",
		X"77",X"77",X"77",X"77",X"77",X"77",X"17",X"77",X"01",X"77",X"00",X"77",X"00",X"17",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"00",X"10",X"00",X"71",X"00",X"71",X"00",X"71",X"00",X"71",X"00",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"99",X"00",X"99",X"00",X"11",X"00",X"00",X"10",X"00",X"91",X"00",X"99",X"00",X"99",X"11",
		X"91",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"11",X"11",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"1A",X"00",X"1A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"AA",X"10",X"AA",X"10",X"AA",X"A1",X"AA",X"A1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"17",X"00",X"77",X"00",X"7F",X"00",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"71",X"00",X"77",X"00",X"77",X"00",X"77",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"01",X"66",X"16",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"01",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"01",X"66",X"16",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"AF",X"00",X"AF",X"00",X"FA",X"00",X"AA",X"01",X"AA",X"01",X"AA",X"1A",X"AA",X"1A",X"AA",
		X"AA",X"10",X"AA",X"10",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"A1",X"00",X"A1",X"00",X"AA",X"00",
		X"1A",X"AA",X"1A",X"AA",X"01",X"AA",X"01",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"11",X"00",X"00",
		X"AA",X"00",X"AA",X"00",X"AA",X"10",X"AA",X"10",X"AA",X"10",X"AA",X"00",X"AA",X"00",X"11",X"00",
		X"00",X"F7",X"01",X"F7",X"01",X"77",X"17",X"77",X"17",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"77",X"00",X"71",X"00",X"71",X"00",X"10",X"00",X"11",X"00",X"77",X"00",X"77",X"10",X"77",X"10",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"11",X"11",X"00",X"00",X"00",
		X"77",X"71",X"77",X"71",X"77",X"71",X"77",X"71",X"77",X"71",X"17",X"10",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"10",X"19",X"91",X"99",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"77",X"11",X"7F",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"17",X"10",X"77",X"71",
		X"16",X"66",X"6F",X"66",X"6F",X"66",X"66",X"66",X"66",X"66",X"16",X"66",X"16",X"66",X"01",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"01",X"66",X"00",X"66",X"00",X"66",X"00",X"66",X"00",X"66",X"00",X"16",X"00",X"01",X"00",X"00",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"11",X"11",X"00",X"00",X"00",X"00",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"61",X"66",X"61",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"10",X"66",X"10",X"66",X"00",X"66",X"00",X"66",X"00",X"61",X"00",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F9",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"19",X"99",X"01",X"99",X"01",X"99",X"19",X"99",
		X"10",X"00",X"10",X"00",X"91",X"00",X"91",X"00",X"91",X"00",X"99",X"00",X"99",X"00",X"99",X"00",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"19",X"99",X"19",X"91",X"01",X"10",X"00",X"00",X"00",
		X"99",X"00",X"99",X"00",X"99",X"10",X"99",X"10",X"99",X"10",X"99",X"00",X"11",X"00",X"00",X"00",
		X"FF",X"77",X"F7",X"77",X"F7",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"77",X"71",X"77",X"71",X"77",X"71",X"77",X"71",X"77",X"10",X"77",X"00",X"71",X"00",X"10",X"00",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"17",X"71",X"01",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
