library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity GFX1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of GFX1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"9C",X"63",X"41",X"9C",X"BE",X"BE",X"41",X"00",X"41",X"14",X"36",X"41",X"63",X"63",X"14",X"00",
		X"41",X"41",X"FF",X"00",X"41",X"41",X"FF",X"00",X"00",X"22",X"77",X"00",X"00",X"00",X"77",X"00",
		X"41",X"FF",X"DD",X"63",X"C9",X"77",X"DD",X"00",X"63",X"14",X"55",X"22",X"77",X"36",X"14",X"00",
		X"36",X"C9",X"C9",X"22",X"FF",X"63",X"C9",X"00",X"14",X"14",X"77",X"00",X"36",X"14",X"55",X"00",
		X"14",X"14",X"FF",X"9C",X"FF",X"9C",X"14",X"00",X"00",X"63",X"77",X"00",X"77",X"41",X"36",X"00",
		X"BE",X"41",X"41",X"22",X"FF",X"63",X"41",X"00",X"00",X"55",X"55",X"77",X"55",X"77",X"55",X"00",
		X"36",X"C9",X"C9",X"BE",X"FF",X"FF",X"C9",X"00",X"00",X"36",X"14",X"41",X"14",X"63",X"14",X"00",
		X"00",X"77",X"88",X"00",X"00",X"00",X"FF",X"00",X"36",X"14",X"55",X"36",X"77",X"36",X"14",X"00",
		X"36",X"C9",X"DD",X"36",X"77",X"C9",X"DD",X"00",X"00",X"55",X"14",X"63",X"63",X"77",X"14",X"00",
		X"9C",X"C9",X"EB",X"00",X"BE",X"C9",X"C9",X"00",X"63",X"14",X"14",X"63",X"77",X"77",X"14",X"00",
		X"AA",X"00",X"88",X"00",X"EB",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"EB",X"00",X"88",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"41",X"00",X"DD",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"DD",X"00",X"41",X"00",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",
		X"08",X"01",X"02",X"0C",X"0C",X"02",X"01",X"08",X"01",X"08",X"04",X"03",X"03",X"04",X"08",X"01",
		X"08",X"81",X"02",X"0C",X"0C",X"02",X"81",X"08",X"01",X"48",X"04",X"03",X"03",X"04",X"48",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"9F",X"F8",X"70",X"FE",X"FE",X"70",X"F8",X"9F",X"63",X"FF",X"BE",X"77",X"77",X"BE",X"FF",X"63",
		X"BE",X"8F",X"FF",X"6B",X"FF",X"CD",X"9F",X"BE",X"41",X"FF",X"FF",X"37",X"77",X"FF",X"FF",X"41",
		X"BE",X"8F",X"FF",X"6B",X"FF",X"CD",X"9F",X"BE",X"41",X"FF",X"FF",X"37",X"77",X"FF",X"FF",X"41",
		X"BE",X"8F",X"FF",X"6B",X"FF",X"CD",X"9F",X"BE",X"41",X"FF",X"FF",X"37",X"77",X"FF",X"FF",X"41",
		X"00",X"84",X"08",X"00",X"00",X"08",X"84",X"00",X"00",X"42",X"01",X"00",X"00",X"01",X"42",X"00",
		X"00",X"86",X"08",X"08",X"08",X"08",X"86",X"00",X"00",X"46",X"01",X"01",X"01",X"01",X"46",X"00",
		X"08",X"87",X"08",X"08",X"08",X"08",X"87",X"08",X"01",X"4E",X"01",X"01",X"01",X"01",X"4E",X"01",
		X"02",X"C8",X"04",X"22",X"02",X"14",X"78",X"22",X"14",X"B1",X"22",X"04",X"14",X"02",X"C1",X"04",
		X"20",X"49",X"10",X"02",X"20",X"04",X"F7",X"02",X"04",X"FE",X"02",X"10",X"04",X"20",X"89",X"10",
		X"22",X"81",X"14",X"20",X"22",X"10",X"8F",X"20",X"10",X"4F",X"20",X"14",X"10",X"22",X"48",X"14",
		X"08",X"B1",X"92",X"84",X"84",X"92",X"B1",X"08",X"01",X"78",X"64",X"42",X"42",X"64",X"78",X"01",
		X"00",X"92",X"84",X"08",X"08",X"84",X"92",X"00",X"00",X"64",X"42",X"01",X"01",X"42",X"64",X"00",
		X"00",X"84",X"08",X"00",X"00",X"08",X"84",X"00",X"00",X"42",X"01",X"00",X"00",X"01",X"42",X"00",
		X"00",X"04",X"08",X"00",X"00",X"08",X"04",X"00",X"00",X"02",X"01",X"00",X"00",X"01",X"02",X"00",
		X"00",X"02",X"04",X"08",X"08",X"04",X"02",X"00",X"00",X"04",X"02",X"01",X"01",X"02",X"04",X"00",
		X"08",X"01",X"02",X"04",X"04",X"02",X"01",X"08",X"01",X"08",X"04",X"02",X"02",X"04",X"08",X"01",
		X"08",X"B1",X"92",X"84",X"84",X"92",X"B1",X"08",X"01",X"78",X"64",X"42",X"42",X"64",X"78",X"01",
		X"08",X"B1",X"9E",X"8C",X"8C",X"9E",X"B1",X"08",X"01",X"78",X"67",X"43",X"43",X"67",X"78",X"01",
		X"08",X"BF",X"92",X"84",X"84",X"92",X"BF",X"08",X"01",X"7F",X"64",X"42",X"42",X"64",X"7F",X"01",
		X"0C",X"B9",X"B1",X"92",X"92",X"B1",X"B9",X"0C",X"03",X"79",X"78",X"64",X"64",X"78",X"79",X"03",
		X"0C",X"B5",X"BD",X"92",X"92",X"BD",X"B5",X"0C",X"03",X"7A",X"7B",X"64",X"64",X"7B",X"7A",X"03",
		X"0C",X"B3",X"B3",X"9E",X"9E",X"B3",X"B3",X"0C",X"03",X"7C",X"7C",X"67",X"67",X"7C",X"7C",X"03",
		X"00",X"00",X"36",X"36",X"36",X"36",X"00",X"00",X"00",X"00",X"36",X"36",X"36",X"36",X"00",X"00",
		X"88",X"55",X"22",X"14",X"14",X"AA",X"55",X"88",X"41",X"AA",X"14",X"22",X"22",X"55",X"AA",X"41",
		X"88",X"36",X"22",X"88",X"9C",X"9C",X"22",X"00",X"63",X"88",X"9C",X"63",X"77",X"77",X"88",X"00",
		X"22",X"22",X"BE",X"00",X"22",X"22",X"BE",X"00",X"00",X"14",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"22",X"BE",X"AA",X"36",X"22",X"BE",X"AA",X"00",X"36",X"C9",X"EB",X"14",X"FF",X"9C",X"C9",X"00",
		X"9C",X"22",X"22",X"14",X"BE",X"36",X"22",X"00",X"88",X"C9",X"FF",X"00",X"DD",X"88",X"EB",X"00",
		X"88",X"88",X"BE",X"88",X"BE",X"88",X"88",X"00",X"00",X"36",X"FF",X"41",X"FF",X"63",X"9C",X"00",
		X"9C",X"22",X"22",X"14",X"BE",X"36",X"22",X"00",X"41",X"AA",X"AA",X"BE",X"EB",X"BE",X"AA",X"00",
		X"9C",X"22",X"22",X"9C",X"BE",X"BE",X"22",X"00",X"00",X"DD",X"C9",X"63",X"C9",X"77",X"C9",X"00",
		X"00",X"BE",X"00",X"00",X"00",X"00",X"BE",X"00",X"9C",X"88",X"EB",X"9C",X"BE",X"9C",X"C9",X"00",
		X"9C",X"22",X"AA",X"9C",X"BE",X"22",X"AA",X"00",X"00",X"EB",X"C9",X"36",X"36",X"FF",X"C9",X"00",
		X"88",X"22",X"36",X"00",X"9C",X"22",X"22",X"00",X"77",X"C9",X"C9",X"36",X"FF",X"FF",X"C9",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BE",X"88",X"88",X"BE",X"BE",X"BE",X"88",X"00",X"63",X"9C",X"9C",X"63",X"77",X"77",X"88",X"00",
		X"9C",X"22",X"22",X"BE",X"BE",X"BE",X"22",X"00",X"36",X"C9",X"C9",X"FF",X"FF",X"FF",X"C9",X"00",
		X"14",X"36",X"22",X"88",X"36",X"9C",X"22",X"00",X"14",X"9C",X"88",X"63",X"9C",X"77",X"88",X"00",
		X"88",X"22",X"36",X"BE",X"9C",X"BE",X"22",X"00",X"63",X"88",X"9C",X"FF",X"77",X"FF",X"88",X"00",
		X"22",X"BE",X"22",X"00",X"22",X"BE",X"22",X"00",X"88",X"FF",X"C9",X"00",X"C9",X"FF",X"C9",X"00",
		X"00",X"00",X"00",X"BE",X"00",X"BE",X"00",X"00",X"88",X"C9",X"C9",X"FF",X"C9",X"FF",X"C9",X"00",
		X"BE",X"36",X"22",X"88",X"BE",X"9C",X"22",X"00",X"C9",X"9C",X"C9",X"63",X"C9",X"77",X"88",X"00",
		X"BE",X"00",X"00",X"BE",X"BE",X"BE",X"00",X"00",X"FF",X"41",X"41",X"FF",X"FF",X"FF",X"41",X"00",
		X"22",X"22",X"BE",X"00",X"22",X"22",X"BE",X"00",X"88",X"88",X"FF",X"00",X"88",X"88",X"FF",X"00",
		X"9C",X"22",X"22",X"14",X"BE",X"36",X"22",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"22",X"88",X"BE",X"BE",X"36",X"BE",X"9C",X"00",X"88",X"41",X"36",X"FF",X"9C",X"FF",X"63",X"00",
		X"22",X"BE",X"22",X"00",X"22",X"BE",X"22",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"BE",X"00",X"00",X"BE",X"BE",X"BE",X"88",X"00",X"FF",X"77",X"77",X"FF",X"FF",X"FF",X"63",X"00",
		X"BE",X"00",X"9C",X"BE",X"BE",X"BE",X"88",X"00",X"FF",X"77",X"41",X"FF",X"FF",X"FF",X"63",X"00",
		X"9C",X"22",X"22",X"9C",X"BE",X"BE",X"22",X"00",X"77",X"88",X"88",X"77",X"FF",X"FF",X"88",X"00",
		X"00",X"88",X"88",X"BE",X"88",X"BE",X"88",X"00",X"77",X"88",X"88",X"FF",X"FF",X"FF",X"88",X"00",
		X"AA",X"22",X"BE",X"9C",X"9C",X"BE",X"AA",X"00",X"77",X"88",X"88",X"77",X"FF",X"FF",X"88",X"00",
		X"22",X"88",X"BE",X"BE",X"36",X"BE",X"9C",X"00",X"77",X"88",X"C9",X"FF",X"FF",X"FF",X"88",X"00",
		X"9C",X"22",X"22",X"14",X"BE",X"36",X"22",X"00",X"00",X"C9",X"DD",X"36",X"55",X"FF",X"C9",X"00",
		X"00",X"00",X"BE",X"00",X"00",X"00",X"BE",X"00",X"88",X"88",X"FF",X"00",X"88",X"88",X"FF",X"00",
		X"9C",X"22",X"22",X"9C",X"BE",X"BE",X"22",X"00",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"9C",X"9C",X"00",X"88",X"88",X"BE",X"00",X"FF",X"41",X"41",X"FF",X"FF",X"FF",X"00",X"00",
		X"BE",X"9C",X"9C",X"BE",X"BE",X"BE",X"88",X"00",X"FF",X"41",X"41",X"FF",X"FF",X"FF",X"63",X"00",
		X"36",X"9C",X"9C",X"36",X"BE",X"BE",X"88",X"00",X"9C",X"77",X"77",X"9C",X"BE",X"BE",X"63",X"00",
		X"00",X"00",X"BE",X"00",X"00",X"00",X"BE",X"00",X"BE",X"FF",X"41",X"00",X"FF",X"BE",X"41",X"00",
		X"22",X"BE",X"22",X"36",X"22",X"BE",X"AA",X"00",X"9C",X"C9",X"FF",X"88",X"BE",X"88",X"EB",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"88",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"41",X"00",X"00",X"00",X"00",X"41",X"00",
		X"00",X"88",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"41",X"00",X"00",X"00",X"00",X"41",X"00",
		X"DF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"DF",X"FF",X"DF",X"FF",X"00",X"00",X"00",X"00",
		X"DF",X"FF",X"DF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"77",X"22",X"00",X"00",X"22",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"41",X"00",X"00",X"00",X"00",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"88",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"FF",X"FF",X"36",X"36",X"FF",X"FF",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"22",X"00",X"00",X"22",X"77",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"80",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"40",X"00",X"FF",X"FF",X"FF",X"FF",X"40",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"40",X"00",
		X"00",X"00",X"00",X"9C",X"00",X"88",X"00",X"88",X"00",X"00",X"00",X"63",X"00",X"41",X"00",X"41",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"40",X"00",X"40",X"00",X"FF",X"FF",X"FF",X"FF",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"41",
		X"9C",X"88",X"BE",X"00",X"BE",X"00",X"9C",X"00",X"63",X"41",X"77",X"00",X"77",X"00",X"63",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"88",X"9C",X"00",X"88",X"00",X"9C",X"00",X"00",X"41",X"63",X"00",X"41",X"00",X"63",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"F7",X"FF",X"00",X"00",X"00",X"00",X"F7",X"FF",X"F7",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"F7",X"FF",X"F7",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"DF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"DF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"DF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"DF",X"FF",X"DF",X"FF",X"00",X"00",X"00",X"00",
		X"DF",X"FF",X"DF",X"FF",X"00",X"00",X"00",X"00",X"DF",X"FF",X"DF",X"FF",X"00",X"00",X"00",X"00",
		X"DF",X"FF",X"DF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"DF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"40",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"40",X"00",X"40",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"40",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"40",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"40",X"00",X"FF",X"FF",X"FF",X"FF",X"40",X"00",X"40",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"02",X"00",X"00",X"00",
		X"00",X"AA",X"22",X"55",X"BE",X"55",X"AA",X"55",X"BE",X"00",X"BE",X"00",X"41",X"00",X"41",X"00",
		X"55",X"AA",X"55",X"BE",X"55",X"22",X"AA",X"00",X"00",X"41",X"00",X"41",X"00",X"BE",X"00",X"BE",
		X"77",X"00",X"77",X"00",X"88",X"00",X"88",X"00",X"00",X"55",X"14",X"AA",X"77",X"AA",X"55",X"AA",
		X"00",X"88",X"00",X"88",X"00",X"77",X"00",X"77",X"AA",X"55",X"AA",X"77",X"AA",X"14",X"55",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"63",X"FF",X"77",X"FF",X"41",X"FF",X"00",X"63",X"00",X"77",X"00",X"41",X"00",
		X"41",X"FF",X"77",X"FF",X"63",X"FF",X"FF",X"FF",X"00",X"41",X"00",X"77",X"00",X"63",X"00",X"FF",
		X"00",X"88",X"00",X"BE",X"00",X"9C",X"00",X"FF",X"88",X"FF",X"BE",X"FF",X"9C",X"FF",X"FF",X"FF",
		X"FF",X"00",X"9C",X"00",X"BE",X"00",X"88",X"00",X"FF",X"FF",X"FF",X"9C",X"FF",X"BE",X"FF",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0B",X"0F",X"0F",X"0F",X"0F",X"0F",X"03",X"0F",X"0F",X"0F",X"03",X"0E",X"0F",X"0B",
		X"00",X"08",X"00",X"68",X"00",X"08",X"00",X"68",X"0C",X"0F",X"0F",X"0F",X"0C",X"0F",X"03",X"0D",
		X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"00",X"FF",X"63",X"FF",X"00",X"FF",X"63",X"FF",
		X"9F",X"F0",X"FF",X"F0",X"9F",X"F0",X"FF",X"F0",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",
		X"0F",X"07",X"0F",X"0F",X"0C",X"0F",X"0F",X"0F",X"0F",X"92",X"93",X"93",X"0F",X"93",X"93",X"93",
		X"F0",X"60",X"F0",X"08",X"F0",X"60",X"F0",X"08",X"4E",X"0E",X"4E",X"0F",X"4E",X"02",X"4E",X"0F",
		X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"63",X"FF",X"00",X"FF",X"63",X"FF",X"00",
		X"F0",X"FF",X"F0",X"9F",X"F0",X"FF",X"F0",X"9F",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",
		X"0F",X"0F",X"0F",X"0E",X"07",X"0F",X"0D",X"0F",X"93",X"93",X"93",X"0F",X"93",X"92",X"93",X"0F",
		X"08",X"F0",X"60",X"F0",X"08",X"F0",X"60",X"F0",X"0F",X"4E",X"0A",X"4E",X"0F",X"4E",X"0E",X"4E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"00",X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"09",X"0F",X"0F",X"03",X"0F",X"0F",X"0F",X"0F",X"0B",X"03",X"0F",X"0E",X"0F",X"03",
		X"68",X"00",X"08",X"00",X"68",X"00",X"08",X"00",X"0F",X"07",X"0F",X"0C",X"0D",X"0F",X"0F",X"0C",
		X"15",X"52",X"17",X"13",X"17",X"2C",X"1F",X"1F",X"50",X"17",X"52",X"54",X"59",X"18",X"19",X"20",
		X"61",X"54",X"68",X"1C",X"69",X"15",X"63",X"1B",X"1F",X"13",X"19",X"FF",X"20",X"00",X"1E",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"DF",X"FF",X"DF",X"FF",X"02",X"00",X"00",X"00",
		X"DF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"DF",X"FF",X"DF",X"FF",X"02",X"00",X"00",X"00",
		X"DF",X"FF",X"DF",X"FF",X"00",X"00",X"00",X"00",X"DF",X"FF",X"DF",X"FF",X"00",X"00",X"00",X"00",
		X"DF",X"FF",X"DF",X"FF",X"00",X"00",X"00",X"00",X"DF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"02",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"02",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"40",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"02",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"02",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"40",X"00",X"40",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"40",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"40",X"00",X"FF",X"FF",X"FF",X"FF",X"40",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"02",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"02",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"DB",X"AF",X"06",X"20",X"09",X"00",X"50",X"5F",X"0B",X"10",X"FC",X"ED",X"56",X"19",X"D9",X"67",
		X"C3",X"C7",X"02",X"3A",X"EC",X"64",X"FE",X"00",X"E0",X"47",X"3E",X"30",X"09",X"35",X"40",X"5F",
		X"2B",X"10",X"FC",X"E1",X"3A",X"ED",X"64",X"FE",X"00",X"E0",X"47",X"3E",X"30",X"09",X"02",X"40",
		X"5F",X"0B",X"10",X"FC",X"E1",X"E1",X"25",X"66",X"20",X"F1",X"F5",X"CD",X"FD",X"CD",X"AF",X"1A",
		X"00",X"30",X"80",X"F0",X"00",X"A0",X"90",X"F0",X"00",X"40",X"20",X"FF",X"40",X"C8",X"60",X"FF",
		X"70",X"E0",X"D0",X"FC",X"E0",X"F0",X"30",X"FE",X"00",X"70",X"D0",X"B0",X"B0",X"F0",X"B0",X"F0",
		X"E0",X"B0",X"F0",X"00",X"F0",X"10",X"B0",X"00",X"88",X"00",X"88",X"00",X"88",X"00",X"00",X"41",
		X"01",X"01",X"07",X"FF",X"03",X"36",X"07",X"BE",X"60",X"03",X"0E",X"08",X"90",X"0E",X"03",X"00",
		X"00",X"30",X"80",X"F0",X"00",X"A0",X"90",X"F0",X"00",X"FE",X"20",X"C9",X"40",X"FF",X"60",X"00",
		X"70",X"E0",X"D0",X"FC",X"E0",X"F0",X"30",X"FE",X"00",X"70",X"D0",X"B0",X"B0",X"F0",X"B0",X"F0",
		X"E0",X"B0",X"F0",X"00",X"F0",X"10",X"B0",X"00",X"41",X"88",X"BE",X"00",X"77",X"00",X"88",X"41",
		X"89",X"01",X"07",X"FF",X"03",X"36",X"07",X"BE",X"60",X"03",X"0E",X"08",X"0C",X"0E",X"03",X"00",
		X"00",X"90",X"00",X"70",X"00",X"B0",X"80",X"F0",X"00",X"BF",X"E8",X"03",X"40",X"89",X"FE",X"07",
		X"F0",X"6C",X"F0",X"0F",X"E0",X"0F",X"F0",X"0F",X"90",X"F0",X"B0",X"78",X"B0",X"F0",X"70",X"6C",
		X"F0",X"80",X"B0",X"00",X"E0",X"00",X"90",X"00",X"07",X"62",X"01",X"40",X"03",X"60",X"23",X"00",
		X"0F",X"F0",X"0F",X"F0",X"0F",X"D0",X"6C",X"F0",X"6C",X"F0",X"D0",X"B0",X"78",X"A0",X"F0",X"90",
		X"00",X"90",X"00",X"E0",X"00",X"B0",X"80",X"F0",X"00",X"FE",X"C8",X"60",X"00",X"C8",X"FE",X"61",
		X"70",X"B1",X"E0",X"FF",X"F0",X"97",X"F0",X"FF",X"90",X"4C",X"B0",X"03",X"30",X"0E",X"F0",X"0F",
		X"D0",X"80",X"B0",X"00",X"F0",X"00",X"10",X"00",X"61",X"62",X"40",X"00",X"60",X"40",X"62",X"00",
		X"FF",X"70",X"97",X"F0",X"FF",X"D0",X"B1",X"70",X"0F",X"F0",X"0E",X"B0",X"03",X"B0",X"4C",X"90",
		X"00",X"00",X"00",X"BE",X"00",X"9C",X"00",X"FF",X"00",X"02",X"01",X"83",X"00",X"02",X"03",X"F0",
		X"07",X"0D",X"0B",X"0F",X"43",X"0F",X"07",X"86",X"0C",X"00",X"0F",X"77",X"07",X"63",X"08",X"FF",
		X"FF",X"00",X"63",X"00",X"FF",X"00",X"EB",X"00",X"F0",X"03",X"82",X"00",X"83",X"01",X"03",X"00",
		X"83",X"07",X"0E",X"4E",X"0F",X"4E",X"0F",X"44",X"61",X"30",X"38",X"80",X"6D",X"90",X"30",X"00",
		X"00",X"00",X"00",X"BE",X"00",X"9C",X"00",X"FF",X"00",X"B1",X"01",X"C0",X"00",X"F0",X"03",X"00",
		X"07",X"0B",X"0D",X"87",X"0B",X"0F",X"30",X"92",X"0C",X"00",X"0F",X"77",X"07",X"63",X"08",X"FF",
		X"FF",X"00",X"63",X"00",X"FF",X"00",X"EB",X"00",X"40",X"83",X"B1",X"00",X"70",X"01",X"82",X"00",
		X"85",X"0F",X"0E",X"4E",X"0F",X"46",X"0F",X"44",X"61",X"30",X"38",X"80",X"6D",X"90",X"30",X"00",
		X"00",X"9C",X"00",X"FF",X"00",X"BE",X"00",X"6F",X"00",X"F1",X"01",X"C1",X"01",X"F1",X"81",X"63",
		X"0F",X"8F",X"03",X"FF",X"0F",X"BF",X"0E",X"FF",X"00",X"30",X"08",X"0F",X"08",X"4F",X"0C",X"9F",
		X"6F",X"00",X"BE",X"00",X"FF",X"00",X"9C",X"00",X"63",X"01",X"61",X"01",X"41",X"01",X"61",X"00",
		X"FF",X"0E",X"BF",X"0F",X"FF",X"0B",X"8F",X"0F",X"9F",X"0C",X"4F",X"08",X"0F",X"08",X"0A",X"00",
		X"00",X"9C",X"00",X"63",X"00",X"BE",X"00",X"FF",X"00",X"B1",X"02",X"81",X"01",X"B1",X"83",X"03",
		X"0F",X"0F",X"0F",X"0F",X"09",X"0B",X"0E",X"0F",X"00",X"6F",X"08",X"30",X"08",X"F7",X"0C",X"F1",
		X"FF",X"00",X"BE",X"00",X"63",X"00",X"9C",X"00",X"03",X"03",X"21",X"01",X"01",X"02",X"21",X"00",
		X"0F",X"0E",X"0F",X"03",X"07",X"0F",X"0F",X"0F",X"F1",X"0C",X"F7",X"08",X"30",X"08",X"6F",X"00",
		X"00",X"9C",X"00",X"63",X"00",X"BE",X"00",X"FF",X"00",X"B1",X"02",X"81",X"01",X"B1",X"83",X"03",
		X"0F",X"0F",X"0F",X"0F",X"09",X"0B",X"0E",X"0F",X"00",X"6F",X"08",X"B0",X"08",X"F7",X"0C",X"F1",
		X"FF",X"00",X"BE",X"00",X"63",X"00",X"9C",X"00",X"03",X"83",X"B1",X"01",X"81",X"02",X"B1",X"00",
		X"0F",X"0E",X"0F",X"03",X"07",X"0F",X"0F",X"0F",X"F1",X"0C",X"F7",X"08",X"30",X"08",X"6F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"63",X"00",X"FF",X"00",X"77",X"00",X"FF",X"00",X"88",X"00",X"BE",X"00",X"9C",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"77",X"00",X"FF",X"00",X"63",X"00",X"FF",X"00",X"9C",X"00",X"BE",X"00",X"88",X"00",
		X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"63",X"00",X"FF",X"00",X"77",X"00",X"FC",X"00",X"FF",X"00",X"F8",X"00",X"FF",X"9C",X"B0",
		X"90",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"00",X"77",X"00",X"FF",X"00",X"63",X"00",X"F0",X"9C",X"FF",X"00",X"F8",X"00",X"FF",X"00",
		X"00",X"B0",X"00",X"E0",X"00",X"F0",X"10",X"F0",X"00",X"00",X"00",X"41",X"00",X"00",X"00",X"41",
		X"00",X"77",X"00",X"FF",X"00",X"77",X"41",X"FC",X"00",X"9C",X"00",X"F0",X"00",X"FF",X"9C",X"F0",
		X"F0",X"10",X"F0",X"00",X"D0",X"00",X"B0",X"00",X"41",X"00",X"00",X"00",X"41",X"00",X"00",X"00",
		X"FC",X"41",X"77",X"00",X"FF",X"00",X"77",X"00",X"D0",X"9C",X"FF",X"00",X"F0",X"00",X"9C",X"00",
		X"00",X"90",X"00",X"B0",X"00",X"B0",X"80",X"B0",X"00",X"00",X"00",X"63",X"00",X"41",X"00",X"63",
		X"00",X"FF",X"00",X"BD",X"00",X"FF",X"77",X"B2",X"00",X"FC",X"00",X"68",X"00",X"B0",X"FE",X"6C",
		X"A0",X"80",X"B0",X"00",X"B0",X"00",X"90",X"00",X"63",X"00",X"41",X"00",X"63",X"00",X"00",X"00",
		X"B2",X"77",X"FF",X"00",X"BD",X"00",X"FF",X"00",X"6C",X"FE",X"B0",X"00",X"68",X"00",X"FC",X"00",
		X"00",X"B0",X"80",X"F0",X"00",X"E0",X"90",X"F0",X"00",X"63",X"41",X"63",X"00",X"63",X"41",X"41",
		X"63",X"FE",X"FF",X"F9",X"FF",X"FD",X"FF",X"F3",X"88",X"F0",X"F8",X"03",X"BC",X"0E",X"E0",X"0F",
		X"F0",X"90",X"F0",X"00",X"D0",X"80",X"B0",X"00",X"41",X"41",X"63",X"00",X"63",X"41",X"63",X"00",
		X"F3",X"FF",X"FD",X"FF",X"F9",X"FF",X"FE",X"63",X"0F",X"F0",X"0E",X"BC",X"03",X"D8",X"F0",X"88",
		X"00",X"90",X"00",X"E0",X"00",X"B0",X"80",X"F0",X"00",X"77",X"63",X"77",X"41",X"77",X"63",X"62",
		X"74",X"BD",X"FE",X"F7",X"FE",X"9B",X"FC",X"FF",X"90",X"4C",X"B0",X"03",X"30",X"0E",X"F0",X"0F",
		X"D0",X"80",X"B0",X"00",X"F0",X"00",X"90",X"00",X"62",X"63",X"77",X"41",X"77",X"63",X"77",X"00",
		X"FF",X"FC",X"9B",X"FE",X"F7",X"FE",X"BD",X"74",X"0F",X"F0",X"0E",X"B0",X"03",X"B0",X"4C",X"90",
		X"00",X"80",X"00",X"F0",X"00",X"B0",X"80",X"F0",X"77",X"FE",X"FE",X"FC",X"77",X"FC",X"FE",X"F9",
		X"70",X"B1",X"F0",X"FF",X"F0",X"97",X"F0",X"FF",X"90",X"4C",X"B0",X"03",X"B0",X"0E",X"F0",X"0F",
		X"F0",X"80",X"B0",X"00",X"F0",X"00",X"80",X"00",X"F9",X"FE",X"FC",X"77",X"FC",X"FE",X"FE",X"77",
		X"FF",X"F0",X"97",X"F0",X"FF",X"F0",X"B1",X"70",X"0F",X"F0",X"0E",X"B0",X"03",X"B0",X"4C",X"90",
		X"00",X"90",X"00",X"E0",X"00",X"B0",X"80",X"F0",X"00",X"FE",X"C8",X"60",X"00",X"C8",X"FE",X"61",
		X"70",X"B1",X"E0",X"FF",X"F0",X"97",X"F0",X"FF",X"90",X"4C",X"B0",X"03",X"30",X"0E",X"F0",X"0F",
		X"D0",X"80",X"B0",X"00",X"F0",X"00",X"10",X"00",X"61",X"FE",X"C8",X"00",X"60",X"C8",X"FE",X"00",
		X"FF",X"70",X"97",X"F0",X"FF",X"D0",X"B1",X"70",X"0F",X"F0",X"0E",X"B0",X"03",X"B0",X"4C",X"90",
		X"15",X"52",X"17",X"13",X"17",X"2C",X"1F",X"1F",X"50",X"17",X"52",X"54",X"59",X"18",X"19",X"20",
		X"61",X"54",X"68",X"1C",X"69",X"15",X"63",X"1B",X"1F",X"13",X"19",X"EC",X"20",X"09",X"1E",X"09",
		X"3E",X"01",X"06",X"04",X"E5",X"85",X"15",X"3A",X"32",X"66",X"E3",X"67",X"28",X"25",X"11",X"ED",
		X"40",X"09",X"B4",X"09",X"3E",X"01",X"06",X"04",X"E5",X"85",X"15",X"3A",X"32",X"66",X"E3",X"57",
		X"28",X"25",X"11",X"EE",X"40",X"09",X"B4",X"09",X"3E",X"01",X"06",X"04",X"E5",X"85",X"15",X"3A",
		X"32",X"66",X"E3",X"77",X"28",X"25",X"11",X"EF",X"40",X"09",X"B4",X"09",X"3E",X"01",X"06",X"04",
		X"E5",X"85",X"15",X"3A",X"32",X"66",X"FE",X"00",X"08",X"26",X"FB",X"3E",X"01",X"1A",X"00",X"50",
		X"3E",X"02",X"E5",X"FF",X"14",X"C3",X"F1",X"02",X"1A",X"C0",X"50",X"30",X"FB",X"01",X"00",X"10",
		X"AF",X"1A",X"C0",X"50",X"86",X"0B",X"57",X"23",X"79",X"98",X"7A",X"08",X"DF",X"FE",X"FF",X"28",
		X"02",X"1F",X"E1",X"1F",X"3F",X"E1",X"20",X"CE",X"FC",X"20",X"CD",X"3E",X"11",X"E5",X"1D",X"05",
		X"C9",X"CD",X"3E",X"0A",X"E5",X"1D",X"05",X"C9",X"CD",X"3E",X"44",X"E5",X"1D",X"05",X"C9",X"3E",
		X"A0",X"E5",X"1D",X"05",X"E1",X"1A",X"C0",X"50",X"CD",X"CD",X"D1",X"13",X"01",X"FF",X"03",X"5F",
		X"ED",X"98",X"C9",X"01",X"00",X"04",X"BE",X"C4",X"53",X"05",X"0B",X"77",X"23",X"79",X"98",X"7B",
		X"08",X"DC",X"E1",X"77",X"7E",X"CE",X"27",X"57",X"7B",X"CE",X"27",X"BA",X"28",X"04",X"20",X"E3",
		X"E7",X"20",X"7E",X"CE",X"D8",X"57",X"7B",X"CE",X"D8",X"BA",X"E0",X"20",X"E3",X"C7",X"20",X"7B",
		X"E1",X"45",X"47",X"47",X"67",X"52",X"2C",X"43",X"67",X"50",X"71",X"52",X"61",X"47",X"60",X"54",
		X"08",X"19",X"39",X"38",X"1B",X"54",X"45",X"64",X"63",X"67",X"08",X"61",X"66",X"43",X"1A",X"C0",
		X"50",X"09",X"00",X"40",X"11",X"01",X"40",X"01",X"FE",X"07",X"1E",X"40",X"ED",X"98",X"1A",X"C0",
		X"50",X"09",X"00",X"64",X"11",X"01",X"64",X"01",X"FE",X"03",X"1E",X"00",X"ED",X"98",X"1A",X"C0",
		X"50",X"09",X"48",X"50",X"11",X"49",X"50",X"01",X"27",X"00",X"1E",X"00",X"ED",X"98",X"1A",X"C0",
		X"50",X"09",X"D8",X"67",X"11",X"D9",X"67",X"01",X"27",X"00",X"1E",X"00",X"ED",X"98",X"1A",X"C0",
		X"50",X"09",X"40",X"50",X"11",X"41",X"50",X"01",X"37",X"00",X"1E",X"00",X"ED",X"98",X"09",X"52",
		X"64",X"11",X"53",X"64",X"01",X"67",X"00",X"1E",X"FF",X"ED",X"98",X"09",X"D6",X"0A",X"0A",X"F1",
		X"00",X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"00",
		X"00",X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"00",
		X"15",X"7E",X"1A",X"E8",X"64",X"78",X"CE",X"18",X"09",X"B8",X"09",X"E5",X"48",X"15",X"0A",X"E9",
		X"64",X"78",X"CE",X"18",X"E3",X"3F",X"E3",X"3F",X"E3",X"3F",X"E3",X"3F",X"1A",X"EB",X"64",X"78",
		X"00",X"00",X"22",X"77",X"77",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C2",X"47",X"11",X"C3",X"47",X"01",X"34",X"00",X"1E",X"05",X"ED",X"98",X"1A",X"C0",X"50",X"09",
		X"CA",X"47",X"11",X"CB",X"47",X"01",X"34",X"00",X"1E",X"21",X"ED",X"98",X"1A",X"C0",X"50",X"09",
		X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"00",X"66",X"FF",X"FF",X"FF",X"FF",X"66",X"00",
		X"FC",X"64",X"11",X"DA",X"43",X"E5",X"D7",X"27",X"09",X"02",X"40",X"11",X"03",X"40",X"01",X"3C",
		X"00",X"1E",X"40",X"ED",X"98",X"1A",X"C0",X"50",X"09",X"02",X"44",X"11",X"03",X"44",X"01",X"34",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"77",X"77",X"22",X"00",X"00",
		X"AF",X"1A",X"24",X"40",X"3A",X"C9",X"64",X"FE",X"00",X"08",X"23",X"09",X"8C",X"35",X"11",X"24",
		X"40",X"01",X"21",X"00",X"ED",X"98",X"1A",X"C0",X"50",X"09",X"42",X"65",X"11",X"43",X"65",X"01",
		X"FF",X"00",X"1E",X"00",X"ED",X"98",X"09",X"3E",X"30",X"0A",X"73",X"65",X"0A",X"43",X"65",X"09",
		X"72",X"65",X"0A",X"62",X"65",X"09",X"58",X"30",X"0A",X"5E",X"65",X"0A",X"76",X"65",X"09",X"5D",
		X"65",X"0A",X"4D",X"65",X"09",X"8A",X"30",X"0A",X"91",X"65",X"0A",X"79",X"65",X"09",X"90",X"65",
		X"0A",X"80",X"65",X"09",X"D4",X"30",X"0A",X"AC",X"65",X"0A",X"94",X"65",X"09",X"AB",X"65",X"0A",
		X"00",X"00",X"00",X"00",X"00",X"88",X"CC",X"88",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"6A",X"31",X"0A",X"FD",X"65",X"0A",X"CD",X"65",X"09",X"FC",X"65",X"0A",X"EC",X"65",X"09",
		X"B4",X"31",X"0A",X"30",X"66",X"0A",X"00",X"66",X"09",X"17",X"66",X"0A",X"07",X"66",X"06",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",
		X"CC",X"EE",X"EE",X"CC",X"88",X"00",X"00",X"00",X"33",X"77",X"77",X"33",X"11",X"00",X"00",X"00",
		X"C0",X"21",X"09",X"F3",X"64",X"E3",X"8E",X"AF",X"1A",X"01",X"50",X"09",X"F4",X"64",X"E3",X"86",
		X"E5",X"BA",X"15",X"1A",X"C0",X"50",X"3E",X"40",X"E5",X"AD",X"14",X"3E",X"21",X"E5",X"BD",X"14",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"88",X"CC",X"CC",X"88",X"00",X"00",X"00",X"00",X"11",X"33",X"33",X"11",X"00",X"00",X"00",
		X"23",X"E5",X"B3",X"15",X"11",X"A5",X"44",X"09",X"B8",X"07",X"3E",X"20",X"06",X"30",X"E5",X"B3",
		X"15",X"11",X"4A",X"46",X"09",X"B9",X"07",X"3E",X"04",X"06",X"04",X"E5",X"B3",X"15",X"11",X"1F",
		X"45",X"09",X"B9",X"07",X"3E",X"04",X"06",X"04",X"E5",X"B3",X"15",X"11",X"20",X"41",X"09",X"A6",
		X"36",X"3E",X"01",X"06",X"10",X"E5",X"85",X"15",X"11",X"B6",X"40",X"09",X"B6",X"36",X"3E",X"01",
		X"06",X"23",X"E5",X"85",X"15",X"11",X"A5",X"40",X"09",X"A9",X"36",X"3E",X"20",X"06",X"30",X"E5",
		X"85",X"15",X"11",X"81",X"40",X"09",X"69",X"37",X"3E",X"05",X"06",X"21",X"E5",X"85",X"15",X"11",
		X"5F",X"42",X"09",X"69",X"37",X"3E",X"05",X"06",X"21",X"E5",X"85",X"15",X"11",X"4A",X"42",X"09",
		X"96",X"37",X"3E",X"04",X"06",X"04",X"E5",X"85",X"15",X"11",X"1F",X"41",X"09",X"96",X"37",X"3E",
		X"04",X"06",X"04",X"E5",X"85",X"15",X"3E",X"04",X"E5",X"FF",X"14",X"09",X"F3",X"64",X"E3",X"6E",
		X"C2",X"C0",X"21",X"E5",X"2D",X"10",X"3E",X"07",X"E5",X"FF",X"14",X"09",X"F3",X"64",X"E3",X"6E",
		X"C2",X"C0",X"21",X"3E",X"40",X"E5",X"AD",X"14",X"11",X"40",X"44",X"09",X"9B",X"07",X"3E",X"15",
		X"06",X"34",X"E5",X"B3",X"15",X"11",X"87",X"46",X"09",X"9D",X"07",X"3E",X"26",X"06",X"05",X"E5",
		X"B3",X"15",X"11",X"70",X"44",X"09",X"9D",X"07",X"3E",X"03",X"06",X"34",X"E5",X"B3",X"15",X"11",
		X"73",X"44",X"09",X"9E",X"07",X"3E",X"03",X"06",X"34",X"E5",X"B3",X"15",X"11",X"C2",X"40",X"09",
		X"8E",X"37",X"3E",X"01",X"06",X"13",X"E5",X"85",X"15",X"11",X"61",X"41",X"09",X"B9",X"37",X"3E",
		X"24",X"06",X"25",X"E5",X"85",X"15",X"3A",X"C9",X"64",X"FE",X"01",X"08",X"27",X"11",X"31",X"41",
		X"09",X"55",X"08",X"3E",X"01",X"06",X"27",X"E5",X"85",X"15",X"30",X"08",X"FE",X"02",X"08",X"27",
		X"11",X"31",X"41",X"09",X"4C",X"08",X"3E",X"01",X"06",X"27",X"E5",X"85",X"15",X"30",X"25",X"11",
		X"31",X"41",X"09",X"5B",X"08",X"3E",X"01",X"06",X"27",X"E5",X"85",X"15",X"11",X"B4",X"40",X"09",
		X"82",X"08",X"3E",X"01",X"06",X"31",X"E5",X"85",X"15",X"3A",X"EB",X"64",X"FE",X"00",X"08",X"27",
		X"11",X"7C",X"41",X"09",X"B3",X"08",X"3E",X"01",X"06",X"06",X"E5",X"85",X"15",X"30",X"1B",X"FE",
		X"01",X"08",X"27",X"11",X"7C",X"41",X"09",X"89",X"08",X"3E",X"01",X"06",X"06",X"E5",X"85",X"15",
		X"30",X"08",X"FE",X"02",X"08",X"27",X"11",X"7C",X"41",X"09",X"8F",X"08",X"3E",X"01",X"06",X"05",
		X"E5",X"85",X"15",X"30",X"25",X"11",X"7C",X"41",X"09",X"AC",X"08",X"3E",X"01",X"06",X"05",X"E5",
		X"85",X"15",X"3E",X"31",X"1A",X"4E",X"41",X"3E",X"07",X"1A",X"4E",X"45",X"3E",X"7C",X"1A",X"AA",
		X"64",X"3E",X"3B",X"1A",X"AB",X"64",X"3E",X"44",X"1A",X"AC",X"64",X"3E",X"07",X"1A",X"AD",X"64",
		X"3E",X"04",X"E5",X"FF",X"14",X"AF",X"1A",X"AA",X"64",X"09",X"F3",X"64",X"E3",X"6E",X"08",X"40",
		X"E5",X"8A",X"0A",X"E5",X"96",X"0A",X"E5",X"AA",X"0A",X"E5",X"B2",X"0A",X"E5",X"AE",X"0A",X"AF",
		X"1A",X"75",X"65",X"1A",X"78",X"65",X"1A",X"93",X"65",X"1A",X"AE",X"65",X"1A",X"E1",X"65",X"1A",
		X"CC",X"65",X"1A",X"FF",X"65",X"E5",X"C5",X"15",X"1A",X"C0",X"50",X"09",X"F3",X"64",X"E3",X"6E",
		X"08",X"26",X"09",X"F4",X"64",X"E3",X"66",X"08",X"02",X"30",X"E6",X"E3",X"A6",X"C3",X"88",X"07",
		X"E5",X"BA",X"15",X"09",X"F3",X"64",X"E3",X"CE",X"E3",X"AE",X"09",X"F4",X"64",X"E3",X"A6",X"E3",
		X"96",X"E3",X"B6",X"09",X"F5",X"64",X"E3",X"96",X"09",X"F4",X"64",X"E3",X"C6",X"09",X"52",X"64",
		X"11",X"53",X"64",X"01",X"67",X"00",X"1E",X"FF",X"ED",X"98",X"3E",X"FF",X"1A",X"01",X"50",X"09",
		X"F5",X"64",X"E3",X"56",X"08",X"27",X"3A",X"41",X"65",X"3C",X"1A",X"41",X"65",X"FE",X"14",X"08",
		X"04",X"E3",X"D6",X"E3",X"F6",X"00",X"1A",X"C0",X"50",X"3E",X"40",X"E5",X"AD",X"14",X"3E",X"03",
		X"E5",X"BD",X"14",X"3A",X"C9",X"64",X"FE",X"00",X"E2",X"B3",X"22",X"3A",X"C8",X"64",X"FE",X"02",
		X"18",X"64",X"11",X"58",X"41",X"09",X"AD",X"35",X"3E",X"01",X"06",X"23",X"E5",X"85",X"15",X"3A",
		X"40",X"50",X"E3",X"6F",X"08",X"5C",X"3A",X"C9",X"64",X"FE",X"00",X"28",X"15",X"3A",X"C8",X"64",
		X"FE",X"02",X"38",X"4E",X"D6",X"02",X"1A",X"C8",X"64",X"3A",X"CB",X"64",X"D6",X"01",X"0F",X"1A",
		X"CB",X"64",X"09",X"F4",X"64",X"E3",X"CE",X"3A",X"E8",X"64",X"1A",X"EC",X"64",X"E5",X"13",X"00",
		X"3A",X"C9",X"64",X"FE",X"00",X"E2",X"DE",X"22",X"E5",X"E5",X"14",X"C3",X"DE",X"22",X"FE",X"04",
		X"18",X"29",X"11",X"26",X"41",X"09",X"B8",X"35",X"3E",X"01",X"06",X"11",X"E5",X"85",X"15",X"11",
		X"10",X"42",X"09",X"E1",X"35",X"3E",X"01",X"06",X"02",X"E5",X"85",X"15",X"11",X"5A",X"41",X"09",
		X"AD",X"35",X"3E",X"01",X"06",X"23",X"E5",X"85",X"15",X"30",X"94",X"11",X"90",X"40",X"09",X"E3",
		X"35",X"3E",X"01",X"06",X"31",X"E5",X"85",X"15",X"30",X"85",X"3A",X"40",X"50",X"E3",X"5F",X"08",
		X"1B",X"3A",X"C9",X"64",X"FE",X"00",X"28",X"15",X"3A",X"C8",X"64",X"FE",X"04",X"38",X"0D",X"D6",
		X"04",X"1A",X"C8",X"64",X"3A",X"CB",X"64",X"D6",X"02",X"0F",X"1A",X"CB",X"64",X"09",X"F4",X"64",
		X"E3",X"8E",X"3A",X"E8",X"64",X"1A",X"EC",X"64",X"1A",X"ED",X"64",X"E5",X"13",X"00",X"E5",X"0C",
		X"00",X"C3",X"48",X"22",X"1A",X"C0",X"50",X"09",X"F3",X"64",X"E3",X"5E",X"08",X"03",X"C3",X"2F",
		X"22",X"E3",X"9E",X"C3",X"06",X"22",X"AF",X"09",X"EE",X"64",X"11",X"EF",X"64",X"01",X"05",X"00",
		X"5F",X"ED",X"98",X"1A",X"DD",X"64",X"1A",X"DE",X"64",X"3E",X"40",X"09",X"CC",X"43",X"11",X"CD",
		X"43",X"01",X"05",X"00",X"5F",X"ED",X"98",X"09",X"DE",X"43",X"11",X"DF",X"43",X"01",X"05",X"00",
		X"5F",X"ED",X"98",X"AF",X"1A",X"CC",X"43",X"1A",X"DE",X"43",X"E5",X"8E",X"0A",X"E5",X"C6",X"0A",
		X"09",X"F5",X"64",X"E3",X"E6",X"09",X"F4",X"64",X"E3",X"4E",X"28",X"02",X"30",X"32",X"3E",X"00",
		X"1A",X"03",X"50",X"E5",X"DC",X"14",X"11",X"50",X"41",X"09",X"CC",X"35",X"3E",X"01",X"06",X"25",
		X"E5",X"85",X"15",X"3E",X"03",X"E5",X"FF",X"14",X"09",X"F4",X"64",X"E3",X"EE",X"3A",X"EC",X"64",
		X"3D",X"1A",X"EC",X"64",X"3E",X"40",X"09",X"16",X"40",X"11",X"17",X"40",X"01",X"20",X"00",X"5F",
		X"ED",X"98",X"E5",X"13",X"00",X"E5",X"BA",X"0A",X"C3",X"DE",X"23",X"09",X"F4",X"64",X"E3",X"4E",
		X"08",X"D6",X"E3",X"6E",X"28",X"B8",X"3A",X"F4",X"64",X"E3",X"7F",X"08",X"1F",X"E5",X"DC",X"14",
		X"11",X"50",X"41",X"09",X"D9",X"35",X"3E",X"01",X"06",X"25",X"E5",X"85",X"15",X"3E",X"03",X"E5",
		X"FF",X"14",X"09",X"F4",X"64",X"E3",X"AE",X"3A",X"ED",X"64",X"3D",X"1A",X"ED",X"64",X"3E",X"40",
		X"09",X"02",X"40",X"11",X"03",X"40",X"01",X"20",X"00",X"5F",X"ED",X"98",X"E5",X"0C",X"00",X"E5",
		X"C2",X"0A",X"30",X"1A",X"3E",X"01",X"1A",X"03",X"50",X"30",X"C2",X"E5",X"DC",X"14",X"09",X"F4",
		X"64",X"E3",X"4E",X"08",X"A0",X"11",X"10",X"41",X"09",X"FE",X"35",X"3E",X"01",X"06",X"11",X"E5",
		X"85",X"15",X"09",X"75",X"65",X"E3",X"C6",X"3E",X"01",X"E5",X"FF",X"14",X"09",X"F4",X"64",X"E3",
		X"6E",X"28",X"9C",X"C3",X"75",X"23",X"E5",X"AA",X"0A",X"09",X"F5",X"64",X"E3",X"66",X"28",X"13",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DE",X"30",X"05",X"3E",X"02",X"E5",X"FF",X"14",X"09",X"CC",X"65",X"E3",X"C6",X"E5",X"AE",X"0A",
		X"00",X"EE",X"22",X"AA",X"AA",X"55",X"55",X"55",X"EE",X"11",X"EE",X"11",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"AA",X"AA",X"22",X"EE",X"00",X"00",X"00",X"00",X"00",X"11",X"EE",X"11",X"EE",
		X"77",X"88",X"77",X"88",X"00",X"00",X"00",X"00",X"00",X"77",X"44",X"55",X"55",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"88",X"77",X"88",X"77",X"AA",X"AA",X"AA",X"55",X"55",X"44",X"77",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"33",X"11",X"FF",X"77",X"33",X"11",X"00",X"00",X"00",X"00",
		X"11",X"33",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"11",X"33",X"77",X"FF",
		X"00",X"00",X"00",X"00",X"88",X"CC",X"EE",X"FF",X"88",X"CC",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"EE",X"CC",X"88",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"CC",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0B",X"0F",X"0F",X"0F",X"0F",X"0F",X"03",X"03",X"0F",X"0F",X"0F",X"0E",X"0F",X"0B",
		X"00",X"00",X"00",X"00",X"08",X"08",X"38",X"38",X"0C",X"0C",X"0F",X"03",X"0F",X"0F",X"0F",X"0D",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"33",X"33",X"FF",X"FF",X"FF",X"FF",
		X"CF",X"CF",X"FF",X"FF",X"F0",X"F0",X"F0",X"F0",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"0F",X"0C",X"0F",X"0F",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"C3",X"C3",X"C2",X"C3",X"C3",X"C3",
		X"F0",X"F0",X"F0",X"F0",X"30",X"30",X"08",X"08",X"1E",X"1E",X"1E",X"1E",X"0E",X"02",X"0F",X"0F",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"33",X"33",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"FF",X"FF",X"CF",X"CF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"07",X"0F",X"0D",X"0F",X"0F",X"0E",X"0F",X"C3",X"C3",X"C3",X"C3",X"C3",X"C2",X"0F",X"0F",
		X"08",X"08",X"30",X"30",X"F0",X"F0",X"F0",X"F0",X"0F",X"0F",X"0A",X"0E",X"1E",X"1E",X"1E",X"1E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"09",X"0F",X"0F",X"03",X"0F",X"0F",X"0F",X"0F",X"0B",X"0F",X"0F",X"0E",X"03",X"03",
		X"38",X"38",X"08",X"08",X"00",X"00",X"00",X"00",X"0F",X"0D",X"0F",X"0F",X"07",X"0F",X"0C",X"0C",
		X"45",X"47",X"47",X"4F",X"52",X"2C",X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",
		X"31",X"39",X"38",X"33",X"54",X"45",X"4C",X"4B",X"4F",X"20",X"49",X"4E",X"43",X"64",X"FD",X"21",
		X"FD",X"5B",X"00",X"FD",X"5A",X"01",X"FD",X"5F",X"02",X"3C",X"13",X"FD",X"5B",X"03",X"FD",X"5A",
		X"04",X"FD",X"5F",X"05",X"3A",X"8A",X"64",X"F5",X"5F",X"03",X"3A",X"8B",X"64",X"F5",X"5F",X"04",
		X"E1",X"3A",X"51",X"64",X"FE",X"00",X"E2",X"73",X"26",X"3A",X"51",X"64",X"E3",X"0F",X"C6",X"27",
		X"F5",X"46",X"05",X"80",X"C1",X"FD",X"09",X"52",X"64",X"FD",X"21",X"FD",X"5B",X"00",X"FD",X"5A",
		X"01",X"FD",X"5F",X"02",X"3C",X"09",X"08",X"00",X"31",X"EB",X"FD",X"5B",X"03",X"FD",X"5A",X"04",
		X"FD",X"5F",X"05",X"C3",X"CC",X"25",X"F5",X"7E",X"03",X"1A",X"8A",X"64",X"F5",X"7E",X"04",X"1A",
		X"8B",X"64",X"C3",X"9D",X"25",X"E5",X"CC",X"26",X"F5",X"7E",X"03",X"80",X"C3",X"AC",X"25",X"E5",
		X"CC",X"26",X"F5",X"7E",X"04",X"90",X"1A",X"8B",X"64",X"F5",X"7E",X"03",X"1A",X"8A",X"64",X"C3",
		X"9D",X"25",X"E5",X"CC",X"26",X"F5",X"7E",X"04",X"80",X"30",X"EB",X"F5",X"7E",X"05",X"C1",X"FD",
		X"09",X"52",X"64",X"FD",X"21",X"FD",X"5B",X"00",X"FD",X"5A",X"01",X"FD",X"5F",X"02",X"3A",X"8A",
		X"64",X"F5",X"5F",X"03",X"3A",X"8B",X"64",X"F5",X"5F",X"04",X"F5",X"7E",X"00",X"09",X"A7",X"26",
		X"E3",X"0F",X"E5",X"48",X"15",X"D5",X"76",X"0B",X"56",X"EB",X"D1",X"F5",X"7E",X"06",X"E9",X"B3",
		X"26",X"B3",X"26",X"B4",X"26",X"8F",X"26",X"AA",X"26",X"99",X"26",X"E1",X"13",X"FD",X"5B",X"03",
		X"FD",X"5A",X"04",X"FD",X"5F",X"05",X"E1",X"33",X"30",X"DB",X"09",X"08",X"00",X"31",X"EB",X"30",
		X"EC",X"EB",X"11",X"08",X"00",X"1F",X"3F",X"ED",X"52",X"EB",X"30",X"C9",X"3A",X"8A",X"64",X"CE",
		X"07",X"1A",X"50",X"64",X"3A",X"8B",X"64",X"CE",X"07",X"1A",X"51",X"64",X"3A",X"8A",X"64",X"E3",
		X"3F",X"E3",X"3F",X"E3",X"3F",X"57",X"3A",X"8B",X"64",X"E3",X"3F",X"E3",X"3F",X"E3",X"3F",X"77",
		X"E5",X"A7",X"14",X"E1",X"F5",X"7E",X"01",X"F5",X"86",X"02",X"47",X"CE",X"27",X"F5",X"5F",X"02",
		X"E3",X"38",X"E3",X"38",X"E3",X"38",X"E3",X"38",X"E1",X"D5",X"1F",X"3F",X"09",X"26",X"01",X"16",
		X"00",X"ED",X"52",X"7D",X"1F",X"3F",X"09",X"10",X"01",X"D1",X"72",X"16",X"00",X"ED",X"52",X"55",
		X"77",X"E1",X"7D",X"EE",X"03",X"6F",X"E1",X"09",X"F4",X"64",X"E3",X"46",X"E0",X"E3",X"6E",X"28",
		X"43",X"09",X"EE",X"64",X"7B",X"86",X"0F",X"5F",X"0B",X"7A",X"A6",X"0F",X"5F",X"0B",X"3E",X"00",
		X"A6",X"0F",X"5F",X"38",X"02",X"30",X"1A",X"09",X"F4",X"64",X"E3",X"6E",X"28",X"13",X"09",X"DE",
		X"43",X"11",X"DF",X"43",X"01",X"05",X"00",X"1E",X"40",X"ED",X"98",X"AF",X"1A",X"DE",X"43",X"30",
		X"30",X"09",X"CC",X"43",X"11",X"CD",X"43",X"01",X"05",X"00",X"1E",X"40",X"ED",X"98",X"AF",X"1A",
		X"CC",X"43",X"30",X"05",X"09",X"D9",X"64",X"30",X"BB",X"09",X"F4",X"64",X"E3",X"6E",X"28",X"74",
		X"09",X"D8",X"64",X"11",X"FB",X"43",X"3A",X"DD",X"64",X"DD",X"E5",X"D7",X"27",X"0B",X"0B",X"0B",
		X"EB",X"2A",X"E9",X"64",X"D9",X"FE",X"04",X"D0",X"E3",X"0F",X"E3",X"0F",X"3C",X"3C",X"E5",X"48",
		X"15",X"E5",X"73",X"11",X"D0",X"3A",X"DC",X"64",X"3C",X"1A",X"DC",X"64",X"09",X"75",X"65",X"E3",
		X"C6",X"09",X"F4",X"64",X"E3",X"6E",X"28",X"12",X"3A",X"DD",X"64",X"3C",X"1A",X"DD",X"64",X"3A",
		X"EC",X"64",X"3C",X"1A",X"EC",X"64",X"E5",X"13",X"00",X"E1",X"3A",X"DE",X"64",X"3C",X"1A",X"DE",
		X"64",X"3A",X"ED",X"64",X"3C",X"1A",X"ED",X"64",X"E5",X"0C",X"00",X"E1",X"09",X"DB",X"64",X"11",
		X"E9",X"43",X"3A",X"DE",X"64",X"30",X"8A",X"3E",X"03",X"DD",X"7E",X"CE",X"D8",X"E3",X"3F",X"E3",
		X"3F",X"E3",X"3F",X"E3",X"3F",X"47",X"3A",X"F4",X"64",X"E3",X"5F",X"28",X"0A",X"78",X"12",X"33",
		X"7E",X"CE",X"27",X"47",X"3A",X"F4",X"64",X"E3",X"5F",X"1A",X"F4",X"64",X"28",X"08",X"78",X"12");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
