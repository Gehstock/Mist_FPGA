library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity pooyan_sprite_grphx2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of pooyan_sprite_grphx2 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"12",X"34",X"69",
		X"00",X"00",X"00",X"00",X"0C",X"C2",X"C2",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"4B",X"4B",X"0F",X"07",X"03",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0E",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"88",X"88",X"00",X"80",X"91",X"00",X"00",X"00",X"11",X"11",X"22",X"20",X"F0",
		X"88",X"00",X"88",X"CC",X"88",X"77",X"74",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"51",X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"F0",X"20",X"22",X"11",X"11",X"00",X"00",X"00",
		X"33",X"77",X"77",X"BB",X"CC",X"88",X"00",X"88",X"00",X"80",X"88",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"10",X"30",X"30",X"00",X"00",X"00",X"70",X"F2",X"F7",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"C0",X"E8",X"EC",X"F4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"70",X"30",X"10",X"10",
		X"F0",X"F4",X"F0",X"E0",X"E0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"22",X"33",X"00",X"00",X"10",X"77",X"FD",X"77",X"FF",X"FF",
		X"00",X"00",X"80",X"CC",X"EE",X"FE",X"FE",X"FF",X"00",X"00",X"00",X"00",X"D1",X"F1",X"E0",X"E0",
		X"33",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"77",X"00",X"00",X"00",
		X"FF",X"FE",X"EE",X"CC",X"88",X"00",X"00",X"00",X"F1",X"F1",X"C0",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"00",X"33",X"33",X"00",X"00",X"00",X"77",X"77",X"FF",X"BF",X"FE",
		X"00",X"40",X"20",X"98",X"CC",X"DC",X"FE",X"F6",X"00",X"00",X"00",X"22",X"F3",X"F3",X"E2",X"E0",
		X"33",X"33",X"11",X"00",X"00",X"00",X"00",X"00",X"FE",X"BF",X"FF",X"FF",X"77",X"00",X"00",X"00",
		X"F6",X"FE",X"DC",X"CC",X"98",X"20",X"40",X"00",X"E0",X"E2",X"F3",X"F3",X"22",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"11",X"33",X"33",X"76",X"00",X"00",X"FF",X"FF",X"FE",X"FC",X"F4",X"F6",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"32",X"33",X"33",X"33",X"11",X"00",X"00",X"00",X"F7",X"FF",X"FE",X"FE",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",X"33",X"00",X"11",X"33",X"11",X"44",X"EE",X"EA",
		X"11",X"00",X"88",X"CC",X"CC",X"C8",X"64",X"70",X"88",X"00",X"00",X"00",X"00",X"60",X"30",X"10",
		X"00",X"00",X"11",X"11",X"00",X"00",X"00",X"00",X"44",X"C8",X"EE",X"EE",X"CC",X"11",X"33",X"11",
		X"F0",X"F0",X"70",X"64",X"C8",X"CC",X"CC",X"88",X"A8",X"88",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"60",X"40",X"00",X"40",X"60",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"C0",X"BB",X"66",X"00",X"00",X"00",X"00",X"66",X"EE",X"11",X"11",
		X"40",X"60",X"40",X"00",X"40",X"60",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"CC",X"FF",X"F3",X"F1",X"F1",X"F1",X"22",X"00",X"00",X"00",X"11",X"88",X"AA",X"99",
		X"66",X"66",X"44",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F3",X"FF",X"F5",X"F7",X"FF",X"EE",X"88",X"00",X"99",X"B9",X"98",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"22",X"33",X"00",X"00",X"10",X"77",X"FF",X"75",X"FF",X"FF",
		X"00",X"00",X"80",X"CC",X"EE",X"FE",X"FF",X"FF",X"00",X"00",X"00",X"40",X"C0",X"F1",X"F1",X"E0",
		X"33",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"77",X"00",X"00",X"00",
		X"FE",X"FE",X"EE",X"CC",X"88",X"00",X"00",X"00",X"E0",X"F1",X"D1",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"8C",X"10",X"10",X"10",X"00",X"10",X"10",X"10",X"00",
		X"00",X"80",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"00",X"10",X"10",X"10",X"00",
		X"00",X"80",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"CC",X"CC",X"00",X"00",X"11",X"11",X"00",X"00",X"00",X"33",X"33",X"D9",X"EE",X"EE",X"CC",
		X"00",X"00",X"00",X"88",X"CC",X"44",X"62",X"F0",X"00",X"00",X"00",X"00",X"00",X"20",X"10",X"B8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"EE",X"EE",X"51",X"33",X"33",X"00",X"11",
		X"F0",X"62",X"44",X"CC",X"88",X"00",X"00",X"99",X"E8",X"00",X"00",X"00",X"00",X"00",X"00",X"88",
		X"C4",X"88",X"00",X"11",X"73",X"E2",X"00",X"11",X"10",X"11",X"11",X"88",X"BB",X"76",X"FE",X"77",
		X"00",X"80",X"00",X"00",X"EE",X"FF",X"FF",X"F2",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"CC",
		X"66",X"DD",X"DD",X"D1",X"51",X"11",X"00",X"00",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"FC",X"33",
		X"FD",X"F7",X"F3",X"F2",X"F3",X"F7",X"FB",X"EE",X"CC",X"CC",X"CC",X"CC",X"CC",X"88",X"00",X"00",
		X"19",X"3F",X"37",X"FF",X"FF",X"FF",X"FF",X"66",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"30",X"F8",X"F8",X"BC",X"DA",X"9E",X"00",X"00",X"80",X"C0",X"C0",X"E3",X"E3",X"E3",
		X"77",X"33",X"11",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"70",X"00",X"00",X"00",X"00",
		X"3C",X"B0",X"80",X"00",X"11",X"11",X"23",X"23",X"C0",X"80",X"AC",X"8E",X"0E",X"0C",X"08",X"00",
		X"40",X"E6",X"C4",X"00",X"11",X"11",X"00",X"C4",X"00",X"20",X"60",X"66",X"DD",X"AA",X"77",X"FF",
		X"00",X"C0",X"C8",X"88",X"77",X"FC",X"F0",X"F0",X"00",X"00",X"00",X"00",X"CC",X"E2",X"E2",X"F1",
		X"C4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FD",X"FE",X"FE",X"FF",X"76",X"33",X"11",X"00",
		X"F0",X"F8",X"FC",X"F7",X"FE",X"FF",X"FF",X"00",X"F1",X"F3",X"F5",X"FF",X"EE",X"CC",X"88",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"60",X"40",X"00",X"40",X"60",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"60",X"40",X"00",X"40",X"60",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"11",X"00",X"00",X"00",X"00",
		X"00",X"88",X"CC",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"11",
		X"00",X"00",X"00",X"00",X"00",X"88",X"CC",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"8C",X"10",X"10",X"10",X"00",X"10",X"10",X"10",X"00",
		X"00",X"80",X"00",X"11",X"33",X"F7",X"77",X"77",X"00",X"00",X"77",X"FF",X"FF",X"FF",X"FF",X"FD",
		X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"00",X"10",X"10",X"10",X"00",
		X"77",X"F7",X"77",X"33",X"33",X"80",X"00",X"00",X"FD",X"F2",X"F3",X"FF",X"FF",X"FE",X"30",X"00",
		X"00",X"00",X"CC",X"EE",X"FF",X"FF",X"FF",X"FF",X"00",X"88",X"CC",X"CC",X"44",X"44",X"60",X"40",
		X"40",X"60",X"40",X"00",X"40",X"60",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FD",X"FD",X"F3",X"EE",X"CC",X"C0",X"80",X"00",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"40",X"60",X"40",X"00",X"40",X"60",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"44",X"44",X"44",X"E4",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"11",X"11",X"00",X"00",
		X"00",X"00",X"00",X"22",X"CC",X"CC",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",
		X"88",X"88",X"88",X"88",X"88",X"88",X"C8",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"11",X"55",X"33",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",
		X"00",X"00",X"98",X"DD",X"CC",X"EE",X"CC",X"CC",X"00",X"00",X"80",X"11",X"11",X"11",X"00",X"00",
		X"FF",X"77",X"76",X"33",X"11",X"00",X"00",X"00",X"FB",X"FC",X"FF",X"FF",X"FF",X"F0",X"00",X"00",
		X"C8",X"D5",X"DD",X"DD",X"BB",X"71",X"20",X"00",X"00",X"00",X"99",X"99",X"99",X"00",X"00",X"00",
		X"00",X"10",X"30",X"CC",X"EE",X"FF",X"FF",X"FE",X"00",X"00",X"88",X"CC",X"CC",X"88",X"88",X"88",
		X"40",X"60",X"40",X"00",X"40",X"60",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FD",X"F3",X"77",X"33",X"33",X"11",X"00",X"00",X"88",X"88",X"88",X"88",X"88",X"00",X"44",X"44",
		X"40",X"60",X"40",X"00",X"40",X"60",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"22",X"00",X"00",X"00",X"00",X"00",X"AA",X"FF",X"BB",
		X"77",X"00",X"22",X"33",X"11",X"CC",X"EE",X"EE",X"00",X"22",X"22",X"11",X"11",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"55",X"00",X"60",X"70",X"22",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"CC",X"EE",X"64",X"64",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"00",X"00",
		X"60",X"73",X"00",X"00",X"51",X"E2",X"11",X"33",X"00",X"00",X"00",X"00",X"00",X"FF",X"F8",X"F0",
		X"22",X"DD",X"CC",X"00",X"11",X"EE",X"FF",X"F7",X"00",X"C8",X"40",X"00",X"00",X"E8",X"40",X"88",
		X"77",X"77",X"77",X"76",X"32",X"33",X"11",X"00",X"F0",X"F8",X"FC",X"FF",X"FF",X"FD",X"FD",X"77",
		X"F3",X"F2",X"F5",X"FB",X"FB",X"FF",X"FF",X"CC",X"CC",X"C4",X"CC",X"CC",X"CC",X"88",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",
		X"00",X"11",X"22",X"00",X"00",X"00",X"00",X"00",X"FF",X"88",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"98",X"44",X"00",X"00",X"00",X"00",X"05",X"A0",X"84",X"E1",X"00",
		X"00",X"00",X"C4",X"00",X"24",X"81",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0C",
		X"10",X"30",X"20",X"00",X"00",X"00",X"00",X"00",X"E1",X"84",X"A1",X"36",X"00",X"00",X"00",X"00",
		X"04",X"81",X"24",X"00",X"44",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"11",X"00",X"EE",X"E8",X"00",
		X"33",X"88",X"88",X"88",X"44",X"40",X"71",X"F1",X"00",X"00",X"11",X"11",X"11",X"00",X"10",X"10",
		X"00",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"CC",X"EC",X"EE",X"CC",X"11",X"33",X"11",X"00",
		X"F1",X"71",X"40",X"44",X"88",X"88",X"88",X"33",X"20",X"00",X"00",X"11",X"11",X"11",X"00",X"00",
		X"00",X"00",X"11",X"B9",X"77",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"88",X"CC",X"CC",X"CC",X"DD",X"DD",X"00",X"00",X"00",X"00",X"C0",X"C8",X"99",X"99",
		X"FF",X"77",X"77",X"32",X"11",X"00",X"00",X"00",X"F7",X"FB",X"FC",X"FF",X"FF",X"F0",X"00",X"00",
		X"DD",X"C8",X"C4",X"88",X"10",X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"11",X"33",X"11",X"E2",
		X"00",X"00",X"44",X"00",X"00",X"88",X"88",X"44",X"00",X"00",X"00",X"00",X"22",X"22",X"22",X"00",
		X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"EE",X"00",X"00",X"E2",X"EE",X"11",X"33",X"11",
		X"00",X"60",X"60",X"00",X"44",X"88",X"88",X"11",X"00",X"E8",X"B8",X"10",X"20",X"22",X"22",X"22",
		X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"30",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"E0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"80",X"D1",X"E6",
		X"70",X"70",X"70",X"70",X"30",X"30",X"10",X"00",X"F0",X"F0",X"F0",X"F0",X"FA",X"F7",X"F0",X"70",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"80",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"30",X"70",X"70",X"F0",X"F0",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"C0",X"E0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"DD",
		X"F0",X"F0",X"F1",X"71",X"30",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"FC",X"FE",X"F0",X"00",X"00",
		X"F0",X"F0",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"A2",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"30",X"70",X"F0",X"F0",X"F0",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"80",X"C0",X"E0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A2",
		X"F0",X"F2",X"73",X"71",X"31",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F9",X"FB",X"F0",X"00",X"00",
		X"F0",X"F0",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"DD",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"30",X"30",X"30",X"00",X"00",X"30",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"80",X"E0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"DD",
		X"30",X"30",X"10",X"10",X"00",X"00",X"00",X"00",X"F0",X"F8",X"FC",X"F2",X"70",X"00",X"00",X"00",
		X"F0",X"F0",X"F4",X"E8",X"C0",X"00",X"00",X"00",X"A2",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"70",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"E0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"80",X"A2",X"DD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F2",X"72",X"71",X"10",X"00",X"00",X"00",X"00",
		X"F0",X"F4",X"F0",X"C0",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"8C",X"10",X"10",X"10",X"00",X"10",X"10",X"10",X"00",
		X"00",X"80",X"00",X"00",X"11",X"B3",X"33",X"77",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FD",
		X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"00",X"10",X"10",X"10",X"00",
		X"77",X"F7",X"77",X"77",X"33",X"B3",X"11",X"00",X"FD",X"FE",X"F3",X"F3",X"FF",X"FF",X"FC",X"60",
		X"D1",X"C0",X"91",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"33",
		X"00",X"CC",X"66",X"EE",X"44",X"CC",X"CC",X"EE",X"00",X"00",X"00",X"00",X"CC",X"66",X"00",X"00",
		X"11",X"00",X"00",X"33",X"00",X"00",X"00",X"00",X"F3",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"77",X"00",X"00",X"00",X"00",X"22",X"88",X"88",X"00",X"00",X"00",X"80",X"D1",X"B3",
		X"60",X"60",X"40",X"00",X"00",X"00",X"00",X"00",X"88",X"11",X"88",X"11",X"88",X"33",X"11",X"33",
		X"00",X"88",X"CC",X"CC",X"88",X"88",X"88",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"11",X"00",X"11",X"00",X"00",X"00",X"00",X"F3",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"CC",X"00",X"00",X"00",X"00",X"10",X"10",X"99",X"55",X"99",X"11",X"00",X"80",X"80",X"00",
		X"30",X"30",X"20",X"00",X"00",X"00",X"00",X"00",X"44",X"11",X"44",X"00",X"55",X"11",X"11",X"33",
		X"00",X"88",X"CC",X"CC",X"88",X"AA",X"88",X"CC",X"00",X"00",X"00",X"00",X"CC",X"66",X"00",X"00",
		X"00",X"11",X"00",X"33",X"00",X"00",X"00",X"00",X"DD",X"E2",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DD",X"DD",X"00",X"00",X"00",X"00",X"10",X"30",X"88",X"CC",X"CC",X"00",X"00",X"80",X"91",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"11",X"33",X"11",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"88",X"CC",X"44",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",
		X"00",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"E8",X"00",X"00",X"E8",X"EE",X"11",X"33",X"11",
		X"00",X"60",X"60",X"00",X"44",X"CC",X"88",X"00",X"10",X"54",X"64",X"00",X"00",X"11",X"99",X"11",
		X"D1",X"C0",X"91",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"33",
		X"00",X"CC",X"66",X"EE",X"44",X"CC",X"CC",X"EE",X"00",X"00",X"00",X"00",X"CC",X"66",X"00",X"00",
		X"11",X"00",X"00",X"33",X"00",X"00",X"00",X"00",X"D1",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"77",X"00",X"00",X"00",X"00",X"22",X"88",X"88",X"00",X"00",X"00",X"80",X"D1",X"B3",
		X"60",X"60",X"40",X"00",X"00",X"00",X"00",X"00",X"88",X"11",X"88",X"11",X"88",X"33",X"11",X"33",
		X"00",X"88",X"CC",X"CC",X"88",X"88",X"88",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"11",X"00",X"11",X"00",X"00",X"00",X"00",X"F3",X"EE",X"CC",X"00",X"00",X"22",X"00",X"00",
		X"FF",X"CC",X"00",X"00",X"00",X"00",X"10",X"10",X"99",X"55",X"11",X"11",X"00",X"80",X"80",X"00",
		X"00",X"00",X"01",X"03",X"02",X"02",X"04",X"0C",X"00",X"00",X"0C",X"0F",X"01",X"CC",X"C8",X"00",
		X"00",X"00",X"00",X"00",X"30",X"0C",X"02",X"60",X"00",X"00",X"00",X"D1",X"11",X"11",X"00",X"00",
		X"0C",X"04",X"02",X"02",X"03",X"01",X"00",X"00",X"00",X"C8",X"CC",X"01",X"0F",X"0C",X"00",X"00",
		X"60",X"02",X"0C",X"60",X"30",X"00",X"00",X"00",X"40",X"51",X"91",X"91",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"F0",X"F0",X"F0",X"70",X"30",X"10",
		X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"11",X"00",X"00",X"33",X"00",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"F3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"CC",X"00",X"22",X"22",X"22",X"00",X"00",X"11",X"33",
		X"00",X"00",X"00",X"00",X"40",X"60",X"60",X"00",X"00",X"11",X"44",X"00",X"88",X"00",X"88",X"00",
		X"CC",X"EE",X"66",X"FF",X"33",X"66",X"00",X"00",X"EE",X"00",X"11",X"11",X"11",X"00",X"00",X"00",
		X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"F9",X"11",X"00",X"11",X"00",
		X"00",X"00",X"66",X"EE",X"CC",X"CC",X"CC",X"66",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"11",X"22",X"91",X"A2",X"00",X"00",X"00",X"00",
		X"EE",X"CC",X"CC",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"07",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"07",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"04",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"0A",X"04",
		X"00",X"00",X"00",X"00",X"00",X"04",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0A",X"02",X"00",X"00",X"00",X"00",X"00",
		X"04",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"07",X"0F",X"0F",X"0F",X"0F",X"07",X"16",X"78",X"F0",X"F0",X"78",X"3C",X"0F",X"0F",
		X"19",X"3F",X"37",X"FF",X"FF",X"FF",X"FF",X"66",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"30",X"F8",X"F8",X"BC",X"8F",X"CF",X"00",X"00",X"80",X"E3",X"E3",X"C4",X"C0",X"E3",
		X"77",X"33",X"11",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"70",X"00",X"00",X"00",X"00",
		X"47",X"8B",X"10",X"10",X"11",X"11",X"23",X"23",X"E3",X"01",X"AC",X"8E",X"0E",X"0C",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"44",X"44",X"33",X"00",X"47",X"44",
		X"00",X"EE",X"11",X"11",X"EE",X"00",X"6E",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"77",X"00",X"33",X"07",X"46",X"22",X"00",
		X"99",X"9F",X"00",X"01",X"0F",X"45",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"3C",X"1E",X"0F",X"0F",X"07",X"03",X"00",X"0F",X"0F",X"3C",X"A5",X"0F",X"0F",X"0F",X"07",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0E",X"08",X"0C",X"0C",X"0C",X"0C",X"08",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"88",X"88",X"77",X"00",X"77",X"88",
		X"00",X"CC",X"22",X"22",X"CC",X"00",X"CC",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"77",X"00",X"66",X"FF",X"DD",X"66",X"11",
		X"22",X"CC",X"00",X"CC",X"EE",X"AA",X"CC",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"88",X"77",X"00",X"77",X"88",X"77",X"00",
		X"CC",X"22",X"CC",X"00",X"CC",X"22",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"99",X"77",X"00",X"00",X"FF",X"44",X"00",
		X"CC",X"22",X"CC",X"00",X"22",X"EE",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"30",X"30",X"70",X"70",X"70",X"71",X"70",X"F0",X"F7",X"F3",X"F0",X"F0",X"F0",X"F0",
		X"00",X"80",X"E8",X"FC",X"FE",X"F6",X"F6",X"F0",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",
		X"71",X"70",X"30",X"10",X"00",X"00",X"00",X"00",X"F8",X"FC",X"F0",X"F0",X"70",X"30",X"10",X"10",
		X"F2",X"F0",X"E0",X"E0",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"30",X"00",X"00",X"00",X"00",X"C0",X"E0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"30",X"30",
		X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"80",X"C0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"31",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"FC",X"F0",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"70",X"70",X"F0",X"F0",X"F0",
		X"00",X"00",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"80",X"E0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F6",X"73",X"70",X"10",X"00",X"00",X"00",X"00",
		X"F0",X"FB",X"F8",X"E0",X"00",X"00",X"00",X"00",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"16",X"16",X"12",X"07",X"00",X"00",X"0B",X"F0",X"F0",X"C3",X"87",X"4B",
		X"00",X"00",X"0B",X"B4",X"87",X"0F",X"0F",X"0F",X"00",X"00",X"08",X"84",X"C2",X"68",X"2C",X"3C",
		X"0F",X"0F",X"87",X"87",X"C3",X"E1",X"78",X"1E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"87",X"87",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"1E",X"1E",X"0F",X"0F",X"0E",X"0E",X"0E",X"0E");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
