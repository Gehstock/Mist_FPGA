library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity twotiger_sp_bits_3 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of twotiger_sp_bits_3 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"EE",X"E0",X"00",X"00",X"55",X"5E",X"00",X"00",X"55",X"55",X"E0",X"0E",X"E5",X"55",X"5E",
		X"E5",X"55",X"55",X"5E",X"E5",X"55",X"55",X"5E",X"E6",X"55",X"EF",X"5E",X"0E",X"6F",X"EE",X"5E",
		X"00",X"EE",X"E0",X"5E",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"5E",
		X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"EE",X"E0",X"00",
		X"00",X"55",X"E0",X"00",X"0E",X"5F",X"00",X"00",X"E5",X"EF",X"E0",X"00",X"E5",X"55",X"5E",X"00",
		X"0E",X"55",X"55",X"00",X"00",X"55",X"55",X"00",X"00",X"FF",X"55",X"00",X"00",X"EE",X"FE",X"00",
		X"00",X"FF",X"EE",X"00",X"00",X"FF",X"0E",X"00",X"00",X"FE",X"0E",X"00",X"00",X"FE",X"00",X"00",
		X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"FE",X"00",X"00",X"EE",X"FE",X"00",X"0E",X"55",X"FE",X"00",
		X"0E",X"E5",X"FE",X"00",X"0E",X"55",X"FE",X"00",X"00",X"55",X"FE",X"00",X"00",X"55",X"EE",X"00",
		X"00",X"F5",X"55",X"00",X"00",X"F6",X"55",X"00",X"00",X"EE",X"55",X"E0",X"00",X"EF",X"55",X"E0",
		X"00",X"FF",X"FF",X"E0",X"00",X"FF",X"EE",X"E0",X"00",X"FF",X"00",X"5E",X"00",X"FF",X"00",X"5E",
		X"00",X"FF",X"00",X"E0",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"FE",X"00",X"00",X"EE",X"FE",X"00",X"0E",X"55",X"FE",X"00",
		X"E5",X"55",X"FE",X"00",X"E5",X"55",X"EE",X"00",X"0E",X"55",X"E0",X"00",X"00",X"55",X"55",X"00",
		X"00",X"55",X"55",X"00",X"00",X"FF",X"5E",X"00",X"00",X"EE",X"5E",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"FF",X"EE",X"00",X"00",X"FF",X"0E",X"00",X"00",X"FF",X"0E",X"00",X"00",X"FF",X"0E",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"FE",X"00",X"00",X"EE",X"FE",X"00",X"00",X"E5",X"FE",X"00",X"0E",X"E5",X"FE",X"00",
		X"00",X"EE",X"FE",X"00",X"00",X"55",X"E0",X"00",X"00",X"55",X"E0",X"00",X"00",X"55",X"00",X"00",
		X"00",X"F5",X"EE",X"00",X"00",X"EF",X"EF",X"00",X"00",X"FE",X"5E",X"00",X"00",X"FF",X"55",X"00",
		X"00",X"FF",X"65",X"00",X"00",X"FF",X"E5",X"00",X"00",X"FF",X"E5",X"00",X"00",X"FE",X"E5",X"00",
		X"00",X"E0",X"E5",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"FE",X"00",X"0E",X"EE",X"FE",X"00",X"0E",X"55",X"FE",X"00",X"00",X"55",X"FE",X"00",
		X"00",X"EE",X"FE",X"00",X"00",X"55",X"FE",X"00",X"00",X"55",X"EE",X"00",X"00",X"55",X"E0",X"00",
		X"00",X"F5",X"EE",X"00",X"00",X"E5",X"55",X"00",X"00",X"EE",X"5E",X"00",X"00",X"EF",X"5E",X"00",
		X"00",X"EF",X"F5",X"00",X"00",X"EF",X"E5",X"00",X"00",X"FF",X"E5",X"00",X"00",X"FF",X"E5",X"00",
		X"00",X"EE",X"55",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"0E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"E0",X"E0",X"00",
		X"00",X"E0",X"FE",X"00",X"00",X"0E",X"FF",X"00",X"00",X"E5",X"FF",X"00",X"00",X"E5",X"FF",X"00",
		X"00",X"55",X"FF",X"00",X"00",X"55",X"FE",X"00",X"00",X"55",X"FE",X"00",X"00",X"F5",X"E0",X"00",
		X"00",X"EF",X"EE",X"00",X"00",X"0E",X"55",X"00",X"00",X"0E",X"55",X"00",X"00",X"0E",X"5E",X"00",
		X"00",X"EF",X"55",X"00",X"00",X"EF",X"EF",X"00",X"00",X"EF",X"EE",X"00",X"00",X"EF",X"0E",X"00",
		X"00",X"EE",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"0E",X"FE",X"00",X"00",X"E5",X"FF",X"00",X"00",X"E5",X"FF",X"00",
		X"00",X"5E",X"FF",X"00",X"00",X"55",X"FE",X"00",X"00",X"55",X"FE",X"00",X"00",X"55",X"E0",X"00",
		X"00",X"F5",X"E0",X"00",X"00",X"EE",X"E0",X"00",X"00",X"EF",X"5E",X"00",X"00",X"FF",X"55",X"00",
		X"00",X"FF",X"EF",X"00",X"00",X"FF",X"5E",X"00",X"00",X"FF",X"55",X"00",X"00",X"FF",X"E5",X"00",
		X"00",X"EE",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"E0",X"00",X"00",X"00",X"EE",X"EE",X"00",X"00",X"5E",X"FF",X"00",X"00",X"55",X"FF",X"00",
		X"00",X"55",X"FF",X"00",X"00",X"55",X"FF",X"00",X"00",X"F5",X"FF",X"00",X"00",X"F5",X"FE",X"00",
		X"00",X"EF",X"EE",X"00",X"00",X"EE",X"5E",X"00",X"00",X"FF",X"5E",X"00",X"00",X"FF",X"5E",X"00",
		X"00",X"FF",X"EF",X"00",X"00",X"FF",X"EF",X"00",X"00",X"FF",X"EF",X"00",X"00",X"EE",X"5E",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EF",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"5E",X"0E",X"00",X"00",X"5E",X"EF",X"00",X"00",X"55",X"FF",X"00",
		X"00",X"55",X"FF",X"00",X"00",X"55",X"FF",X"00",X"00",X"65",X"FF",X"00",X"00",X"F5",X"FF",X"00",
		X"00",X"EE",X"FE",X"00",X"00",X"E6",X"E0",X"00",X"00",X"FF",X"E0",X"00",X"00",X"FF",X"5E",X"00",
		X"00",X"FF",X"5E",X"00",X"00",X"FF",X"EF",X"00",X"00",X"EE",X"5F",X"00",X"00",X"00",X"5F",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"5E",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"55",X"0E",X"00",X"00",X"55",X"EF",X"00",
		X"00",X"55",X"FF",X"00",X"00",X"F5",X"FF",X"00",X"00",X"65",X"FF",X"00",X"00",X"E5",X"FF",X"00",
		X"00",X"E5",X"FE",X"00",X"00",X"F6",X"E0",X"00",X"00",X"FE",X"00",X"00",X"00",X"F6",X"E0",X"00",
		X"00",X"FF",X"EE",X"00",X"00",X"FF",X"FF",X"00",X"00",X"EE",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"EF",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"5E",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"5E",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"55",X"EE",X"00",X"00",X"65",X"EF",X"00",
		X"00",X"F5",X"FF",X"00",X"00",X"65",X"FF",X"00",X"00",X"EF",X"FF",X"00",X"00",X"E6",X"FF",X"00",
		X"00",X"EE",X"FE",X"00",X"00",X"FE",X"E0",X"00",X"00",X"FE",X"E0",X"00",X"00",X"FF",X"E0",X"00",
		X"00",X"FF",X"5E",X"00",X"00",X"FF",X"EE",X"00",X"00",X"EE",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"EF",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"5E",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"5E",X"00",X"00",
		X"00",X"E5",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"F5",X"EE",X"00",
		X"00",X"65",X"FE",X"00",X"00",X"F5",X"FF",X"00",X"00",X"E6",X"FF",X"00",X"00",X"E5",X"FF",X"00",
		X"00",X"FE",X"FF",X"00",X"00",X"FE",X"FE",X"00",X"00",X"FE",X"EE",X"00",X"00",X"FE",X"E0",X"00",
		X"00",X"FF",X"E0",X"00",X"00",X"FE",X"EE",X"00",X"00",X"EE",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FE",X"00",X"00",X"00",X"FE",X"00",X"00",X"00",X"5E",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"E5",X"00",X"00",X"00",X"65",X"00",X"00",X"00",X"65",X"00",X"00",X"00",X"F5",X"00",X"00",
		X"00",X"EF",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"65",X"00",X"00",
		X"00",X"EF",X"00",X"00",X"00",X"E6",X"EE",X"00",X"00",X"EF",X"FF",X"00",X"00",X"E6",X"FF",X"00",
		X"00",X"FE",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FE",X"FF",X"00",X"00",X"FE",X"EE",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"FE",X"00",
		X"00",X"00",X"FE",X"00",X"00",X"00",X"FE",X"00",X"00",X"00",X"E0",X"00",X"00",X"0E",X"E0",X"00",
		X"00",X"0E",X"E0",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"E6",X"00",X"00",X"00",X"E6",X"00",X"00",X"00",X"EF",X"FE",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"FE",X"00",X"00",X"00",X"EF",X"00",X"00",X"00",X"E6",X"00",X"00",X"00",X"EF",X"00",X"00",
		X"00",X"E6",X"00",X"00",X"00",X"EF",X"EE",X"00",X"00",X"E6",X"FF",X"00",X"00",X"E5",X"FF",X"00",
		X"00",X"FE",X"FF",X"00",X"00",X"EF",X"FF",X"00",X"00",X"E1",X"FF",X"00",X"00",X"FE",X"FF",X"00",
		X"00",X"FE",X"EE",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"FE",X"00",X"00",X"EE",X"E0",X"00",
		X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",X"EF",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"0E",X"E0",X"00",X"00",X"0E",X"E0",X"00",X"00",X"0E",X"E0",X"00",
		X"00",X"0E",X"EE",X"00",X"00",X"0E",X"EE",X"00",X"00",X"0E",X"FE",X"00",X"00",X"0E",X"FE",X"00",
		X"00",X"0F",X"FE",X"00",X"00",X"0F",X"FE",X"00",X"00",X"0F",X"FE",X"00",X"00",X"0E",X"FE",X"00",
		X"00",X"0E",X"EE",X"00",X"00",X"0E",X"E0",X"00",X"00",X"0E",X"E0",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"E0",X"99",X"00",X"00",X"E0",X"99",X"00",X"00",X"E0",X"99",X"00",X"00",
		X"BE",X"9E",X"0E",X"00",X"BE",X"99",X"EE",X"00",X"BE",X"E9",X"E9",X"00",X"BB",X"FE",X"E9",X"E0",
		X"EE",X"EB",X"EE",X"BE",X"9E",X"BB",X"BE",X"B9",X"99",X"EE",X"BB",X"B9",X"99",X"99",X"BB",X"9E",
		X"9E",X"99",X"BB",X"E0",X"9E",X"99",X"EB",X"00",X"EE",X"9E",X"EE",X"00",X"00",X"99",X"00",X"00",
		X"00",X"9E",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"E9",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"E0",X"9B",X"00",X"00",X"E0",X"BB",X"00",X"00",X"E0",X"BB",X"00",X"00",
		X"AE",X"B1",X"0E",X"00",X"AE",X"BB",X"EE",X"00",X"EA",X"B1",X"AA",X"00",X"EA",X"BB",X"EE",X"E0",
		X"BE",X"BB",X"EB",X"BE",X"BE",X"EE",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BE",X"EE",X"BB",X"BE",X"BE",X"BE",X"EB",X"E0",X"E0",X"BB",X"0E",X"00",
		X"E0",X"BE",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"9B",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"E9",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"E2",X"00",X"00",X"0F",X"22",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"E0",X"FE",X"EE",X"00",X"E0",X"EE",X"3E",X"00",X"E0",X"EF",X"EE",X"00",
		X"2E",X"EE",X"EE",X"00",X"2E",X"EE",X"EE",X"00",X"2E",X"E1",X"EE",X"00",X"22",X"11",X"EE",X"E0",
		X"EE",X"11",X"EE",X"FE",X"2E",X"EF",X"1E",X"FF",X"22",X"EF",X"1E",X"FF",X"92",X"33",X"1E",X"FE",
		X"2E",X"31",X"1E",X"E0",X"2E",X"11",X"EE",X"00",X"EE",X"F1",X"EE",X"00",X"00",X"1E",X"E0",X"00",
		X"00",X"E1",X"EE",X"00",X"00",X"EF",X"3E",X"00",X"0E",X"EF",X"31",X"00",X"FE",X"EF",X"11",X"00",
		X"0E",X"EF",X"EE",X"00",X"0E",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"E2",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"13",X"00",X"00",X"0F",X"11",X"00",X"00",
		X"00",X"F1",X"00",X"00",X"E0",X"FE",X"EE",X"00",X"E0",X"EE",X"EE",X"F0",X"E0",X"1E",X"EE",X"00",
		X"2E",X"1E",X"EE",X"00",X"31",X"1E",X"EE",X"00",X"33",X"1E",X"E1",X"00",X"22",X"EE",X"E1",X"E0",
		X"11",X"EE",X"E1",X"FE",X"11",X"EE",X"E1",X"FF",X"22",X"EE",X"EE",X"FF",X"31",X"EE",X"EE",X"FE",
		X"31",X"EE",X"EE",X"E0",X"11",X"EE",X"EE",X"00",X"11",X"EE",X"EE",X"00",X"13",X"EE",X"E3",X"0F",
		X"13",X"E3",X"E3",X"00",X"31",X"1E",X"EE",X"F0",X"33",X"1E",X"EE",X"00",X"FE",X"1E",X"EE",X"F0",
		X"0E",X"EE",X"EE",X"00",X"01",X"32",X"33",X"00",X"01",X"22",X"33",X"00",X"00",X"E2",X"13",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"AA",X"EA",X"00",X"0E",X"AA",X"AE",X"00",X"0A",X"AA",X"AE",X"00",X"0A",X"AA",X"AE",X"00",
		X"00",X"AA",X"AE",X"00",X"00",X"AA",X"B3",X"00",X"00",X"A1",X"BE",X"00",X"00",X"AA",X"EE",X"00",
		X"00",X"EE",X"EE",X"E0",X"00",X"EE",X"A3",X"E0",X"00",X"AA",X"E3",X"EE",X"00",X"AA",X"EE",X"EE",
		X"00",X"AA",X"EE",X"2E",X"00",X"AA",X"EE",X"BE",X"00",X"AA",X"E9",X"9E",X"00",X"BB",X"E9",X"E0",
		X"00",X"B9",X"EE",X"00",X"00",X"B9",X"AE",X"00",X"00",X"99",X"AE",X"00",X"00",X"9E",X"AE",X"00",
		X"00",X"E0",X"EE",X"00",X"00",X"00",X"E3",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",
		X"00",X"00",X"E3",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E3",X"00",X"00",X"00",X"EE",X"AA",X"00",
		X"00",X"AE",X"0A",X"00",X"00",X"2A",X"0A",X"00",X"00",X"EE",X"A1",X"00",X"00",X"0E",X"AA",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"0A",X"A0",X"00",X"00",X"EA",X"00",X"00",
		X"00",X"AA",X"E0",X"00",X"00",X"2A",X"E0",X"00",X"00",X"E0",X"E0",X"00",X"EE",X"00",X"00",X"00",
		X"AA",X"00",X"00",X"00",X"EA",X"22",X"00",X"00",X"E0",X"22",X"00",X"00",X"E0",X"E2",X"00",X"00",
		X"0A",X"E3",X"00",X"00",X"00",X"EA",X"00",X"00",X"0A",X"EA",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"E0",X"EE",X"00",X"00",X"E0",X"AE",X"E0",X"00",X"AE",X"3A",X"E0",X"00",X"AE",X"A3",X"E0",X"00",
		X"AA",X"EA",X"E0",X"00",X"AA",X"2A",X"AE",X"00",X"EE",X"EE",X"AE",X"00",X"0E",X"EE",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",
		X"00",X"E0",X"00",X"00",X"EE",X"AE",X"00",X"00",X"AA",X"CE",X"00",X"00",X"AE",X"CE",X"00",X"00",
		X"AA",X"EE",X"EE",X"00",X"EE",X"5E",X"77",X"00",X"EE",X"5E",X"EE",X"00",X"AA",X"55",X"AA",X"E0",
		X"EE",X"55",X"EE",X"E0",X"BB",X"AA",X"77",X"E0",X"EB",X"EE",X"BB",X"EE",X"EE",X"9B",X"EE",X"BE",
		X"0E",X"BB",X"EE",X"BE",X"00",X"BB",X"99",X"BE",X"00",X"2B",X"99",X"9E",X"00",X"B2",X"B2",X"9E",
		X"00",X"EF",X"FE",X"22",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"0F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"00",X"99",X"00",X"00",X"0E",X"99",X"00",X"00",X"E9",X"A1",X"00",X"00",X"E2",X"21",X"00",
		X"00",X"1E",X"11",X"00",X"00",X"1E",X"1E",X"F0",X"00",X"EE",X"1E",X"00",X"00",X"E1",X"EE",X"00",
		X"00",X"11",X"EE",X"00",X"F0",X"11",X"E1",X"F0",X"00",X"11",X"11",X"E0",X"0E",X"1F",X"1E",X"E0",
		X"E2",X"1F",X"1E",X"2E",X"22",X"E1",X"11",X"22",X"22",X"11",X"EE",X"22",X"E2",X"33",X"EE",X"2E",
		X"0E",X"31",X"31",X"E0",X"00",X"11",X"31",X"00",X"00",X"F1",X"33",X"00",X"F0",X"11",X"11",X"00",
		X"00",X"EE",X"EE",X"00",X"00",X"0E",X"EE",X"00",X"00",X"0E",X"EF",X"00",X"00",X"0E",X"E2",X"00",
		X"00",X"0E",X"E3",X"00",X"00",X"0E",X"EE",X"00",X"00",X"0E",X"11",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"99",X"00",X"10",X"E2",X"9E",X"00",X"10",X"11",X"E9",X"01",X"13",X"11",X"E1",X"01",X"10",
		X"01",X"EE",X"11",X"10",X"01",X"1E",X"11",X"30",X"0E",X"E1",X"1E",X"00",X"3E",X"E1",X"EE",X"00",
		X"3E",X"E1",X"EE",X"00",X"E1",X"11",X"EE",X"00",X"11",X"E1",X"EE",X"00",X"E1",X"EE",X"EE",X"01",
		X"EE",X"E1",X"E1",X"00",X"EE",X"E1",X"3E",X"00",X"11",X"E1",X"EE",X"00",X"11",X"EE",X"EE",X"00",
		X"E0",X"EE",X"EE",X"11",X"E0",X"EE",X"EE",X"11",X"E0",X"EE",X"EE",X"11",X"EE",X"EE",X"EE",X"11",
		X"EE",X"EE",X"33",X"31",X"EE",X"EE",X"3E",X"11",X"12",X"EE",X"33",X"10",X"E1",X"3E",X"33",X"30",
		X"E1",X"13",X"31",X"00",X"E1",X"33",X"31",X"00",X"EE",X"33",X"11",X"00",X"EE",X"11",X"1E",X"00",
		X"EE",X"11",X"EE",X"00",X"00",X"11",X"E0",X"00",X"00",X"EE",X"E0",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"62",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"00",
		X"00",X"F6",X"22",X"00",X"00",X"22",X"00",X"00",X"06",X"FF",X"00",X"00",X"00",X"02",X"66",X"00",
		X"00",X"22",X"60",X"00",X"00",X"00",X"20",X"00",X"00",X"20",X"20",X"00",X"06",X"20",X"22",X"00",
		X"06",X"20",X"2F",X"00",X"00",X"20",X"2F",X"60",X"00",X"20",X"FF",X"00",X"00",X"F2",X"F2",X"06",
		X"F2",X"F2",X"F2",X"02",X"02",X"F2",X"22",X"02",X"00",X"26",X"22",X"00",X"0F",X"26",X"2F",X"00",
		X"00",X"26",X"2F",X"00",X"00",X"22",X"2F",X"00",X"00",X"62",X"22",X"60",X"60",X"62",X"02",X"22",
		X"00",X"62",X"02",X"02",X"00",X"22",X"F2",X"00",X"00",X"22",X"F2",X"00",X"00",X"22",X"02",X"00",
		X"00",X"00",X"60",X"00",X"00",X"00",X"20",X"00",X"00",X"20",X"00",X"00",X"00",X"60",X"00",X"00",
		X"00",X"20",X"00",X"00",X"06",X"26",X"60",X"00",X"22",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"06",X"20",X"00",X"00",X"20",X"20",X"02",X"00",
		X"00",X"60",X"02",X"00",X"00",X"20",X"06",X"00",X"00",X"26",X"20",X"66",X"00",X"02",X"60",X"06",
		X"00",X"07",X"00",X"02",X"00",X"07",X"02",X"02",X"00",X"27",X"22",X"00",X"00",X"26",X"22",X"00",
		X"60",X"26",X"26",X"00",X"00",X"27",X"66",X"00",X"00",X"27",X"62",X"00",X"00",X"27",X"27",X"00",
		X"00",X"27",X"22",X"00",X"00",X"27",X"72",X"00",X"00",X"27",X"72",X"00",X"00",X"27",X"72",X"60",
		X"00",X"27",X"72",X"00",X"00",X"22",X"72",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"86",X"00",
		X"00",X"00",X"C4",X"00",X"00",X"00",X"64",X"00",X"00",X"00",X"64",X"00",X"00",X"00",X"64",X"00",
		X"00",X"00",X"64",X"00",X"00",X"00",X"64",X"00",X"00",X"00",X"64",X"00",X"00",X"00",X"64",X"00",
		X"00",X"00",X"64",X"00",X"00",X"00",X"64",X"00",X"00",X"00",X"64",X"00",X"00",X"00",X"64",X"00",
		X"00",X"00",X"64",X"00",X"00",X"00",X"EF",X"00",X"00",X"00",X"FF",X"00",X"00",X"70",X"FF",X"00",
		X"00",X"EF",X"F0",X"00",X"0F",X"7F",X"7F",X"00",X"00",X"00",X"0F",X"00",X"FF",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"FE",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"EF",X"E0",X"00",X"00",X"6E",X"E0",X"00",
		X"00",X"66",X"00",X"00",X"EE",X"AA",X"E0",X"00",X"66",X"FF",X"FE",X"00",X"66",X"FF",X"EE",X"E0",
		X"66",X"FF",X"FF",X"EE",X"E6",X"FF",X"66",X"FF",X"EA",X"FF",X"EE",X"FF",X"EA",X"FF",X"EB",X"BB",
		X"AA",X"FF",X"BA",X"BD",X"FF",X"FE",X"AA",X"BE",X"FF",X"EE",X"AA",X"E0",X"FF",X"EE",X"EE",X"00",
		X"EE",X"1E",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"1E",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"E1",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"DD",X"00",X"00",
		X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"ED",X"00",X"00",
		X"00",X"ED",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"EE",X"00",X"00",X"EB",X"BB",X"00",X"00",X"0E",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"EE",X"F0",X"00",X"60",X"7E",X"7F",X"F0",X"7F",X"F7",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"EA",X"00",X"0F",X"00",X"EC",X"00",X"E0",X"00",X"EC",X"0F",
		X"EE",X"00",X"EC",X"F0",X"BB",X"77",X"EC",X"97",X"77",X"70",X"7E",X"00",X"F0",X"00",X"77",X"70",
		X"00",X"00",X"10",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"EE",X"00",
		X"00",X"00",X"EA",X"00",X"00",X"00",X"AA",X"00",X"EE",X"00",X"AE",X"00",X"ED",X"00",X"AF",X"EE",
		X"DB",X"00",X"AC",X"EB",X"EB",X"00",X"AA",X"BB",X"EB",X"00",X"AE",X"EE",X"EE",X"77",X"EE",X"EE",
		X"EE",X"77",X"BB",X"BB",X"7E",X"00",X"BB",X"B7",X"77",X"70",X"E7",X"70",X"F0",X"07",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"E2",X"00",X"00",
		X"00",X"E2",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",
		X"E0",X"2E",X"E0",X"00",X"20",X"22",X"E0",X"00",X"2E",X"E2",X"EE",X"00",X"22",X"FE",X"E2",X"00",
		X"EE",X"E2",X"EE",X"00",X"2E",X"22",X"2E",X"00",X"2E",X"EE",X"22",X"00",X"2E",X"22",X"22",X"00",
		X"2E",X"22",X"EE",X"00",X"E0",X"22",X"00",X"00",X"00",X"2E",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"2E",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"22",X"00",X"00",X"00",X"E2",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"E2",X"00",X"00",X"05",X"66",X"00",X"00",
		X"00",X"55",X"00",X"00",X"E0",X"5E",X"EE",X"00",X"E0",X"EE",X"7E",X"00",X"E0",X"E5",X"EE",X"00",
		X"6E",X"EE",X"EE",X"00",X"6E",X"22",X"EE",X"00",X"2E",X"62",X"EE",X"00",X"22",X"22",X"EE",X"E0",
		X"EE",X"22",X"EE",X"5E",X"2E",X"22",X"26",X"55",X"22",X"2E",X"26",X"55",X"E2",X"22",X"2E",X"5E",
		X"6E",X"2E",X"2E",X"E0",X"6E",X"22",X"2E",X"00",X"EE",X"52",X"22",X"00",X"E0",X"26",X"22",X"00",
		X"E0",X"22",X"EE",X"00",X"E0",X"E5",X"2E",X"00",X"0E",X"E5",X"27",X"00",X"5E",X"E5",X"77",X"00",
		X"0E",X"E5",X"EE",X"00",X"0E",X"66",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"E2",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"EE",X"E0",X"00",X"00",X"CC",X"CE",X"00",X"00",X"CC",X"CC",X"E0",X"0E",X"EC",X"CC",X"CE",
		X"EC",X"CC",X"CC",X"CE",X"EC",X"CC",X"CC",X"CE",X"EB",X"CC",X"EB",X"CE",X"0E",X"BB",X"EE",X"CE",
		X"00",X"EE",X"E0",X"CE",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"CE",
		X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"EE",X"E0",X"00",
		X"00",X"CC",X"E0",X"00",X"0E",X"CD",X"00",X"00",X"EC",X"ED",X"E0",X"00",X"EC",X"CC",X"CE",X"00",
		X"0E",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"BB",X"CC",X"00",X"00",X"EE",X"BE",X"00",
		X"00",X"DD",X"EE",X"00",X"00",X"DD",X"0E",X"00",X"00",X"DE",X"0E",X"00",X"00",X"DE",X"00",X"00",
		X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"DE",X"00",X"00",X"EE",X"DE",X"00",X"0E",X"CC",X"DE",X"00",
		X"0E",X"EC",X"DE",X"00",X"0E",X"CC",X"DE",X"00",X"00",X"CC",X"DE",X"00",X"00",X"CC",X"EE",X"00",
		X"00",X"BC",X"CC",X"00",X"00",X"BB",X"CC",X"00",X"00",X"EE",X"CC",X"E0",X"00",X"ED",X"CC",X"E0",
		X"00",X"DD",X"BB",X"E0",X"00",X"DD",X"EE",X"E0",X"00",X"DD",X"00",X"CE",X"00",X"DD",X"00",X"CE",
		X"00",X"DD",X"00",X"E0",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"DE",X"00",X"00",X"EE",X"DE",X"00",X"0E",X"CC",X"DE",X"00",
		X"EC",X"CC",X"DE",X"00",X"EC",X"CC",X"EE",X"00",X"0E",X"CC",X"E0",X"00",X"00",X"CC",X"CC",X"00",
		X"00",X"CC",X"CC",X"00",X"00",X"BB",X"CE",X"00",X"00",X"EE",X"CE",X"00",X"00",X"DD",X"BB",X"00",
		X"00",X"DD",X"EE",X"00",X"00",X"DD",X"0E",X"00",X"00",X"DD",X"0E",X"00",X"00",X"DD",X"0E",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"DE",X"00",X"00",X"EE",X"DE",X"00",X"00",X"EC",X"DE",X"00",X"0E",X"EC",X"DE",X"00",
		X"00",X"EE",X"DE",X"00",X"00",X"CC",X"E0",X"00",X"00",X"CC",X"E0",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"BC",X"EE",X"00",X"00",X"EB",X"ED",X"00",X"00",X"DE",X"CE",X"00",X"00",X"DD",X"CC",X"00",
		X"00",X"DD",X"BC",X"00",X"00",X"DD",X"EC",X"00",X"00",X"DD",X"EC",X"00",X"00",X"DE",X"EC",X"00",
		X"00",X"E0",X"EC",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"DE",X"00",X"0E",X"EE",X"DE",X"00",X"0E",X"CC",X"DE",X"00",X"00",X"CC",X"DE",X"00",
		X"00",X"EE",X"DE",X"00",X"00",X"CC",X"DE",X"00",X"00",X"CC",X"EE",X"00",X"00",X"CC",X"E0",X"00",
		X"00",X"BC",X"EE",X"00",X"00",X"EC",X"CC",X"00",X"00",X"EE",X"CE",X"00",X"00",X"ED",X"CE",X"00",
		X"00",X"ED",X"BC",X"00",X"00",X"ED",X"EC",X"00",X"00",X"DD",X"EC",X"00",X"00",X"DD",X"EC",X"00",
		X"00",X"EE",X"CC",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"0E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"E0",X"E0",X"00",
		X"00",X"E0",X"DE",X"00",X"00",X"0E",X"DD",X"00",X"00",X"EC",X"DD",X"00",X"00",X"EC",X"DD",X"00",
		X"00",X"CC",X"DD",X"00",X"00",X"CC",X"DE",X"00",X"00",X"CC",X"DE",X"00",X"00",X"BC",X"E0",X"00",
		X"00",X"EB",X"EE",X"00",X"00",X"0E",X"EC",X"00",X"00",X"0E",X"CC",X"00",X"00",X"0E",X"CC",X"00",
		X"00",X"ED",X"CC",X"00",X"00",X"ED",X"EB",X"00",X"00",X"ED",X"EE",X"00",X"00",X"ED",X"0E",X"00",
		X"00",X"EE",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"0E",X"DE",X"00",X"00",X"EC",X"DD",X"00",X"00",X"EC",X"DD",X"00",
		X"00",X"CE",X"DD",X"00",X"00",X"CC",X"DE",X"00",X"00",X"CC",X"DE",X"00",X"00",X"CC",X"E0",X"00",
		X"00",X"BC",X"E0",X"00",X"00",X"EE",X"E0",X"00",X"00",X"ED",X"CE",X"00",X"00",X"DD",X"CC",X"00",
		X"00",X"DD",X"CD",X"00",X"00",X"DD",X"CD",X"00",X"00",X"DD",X"CC",X"00",X"00",X"DD",X"EC",X"00",
		X"00",X"EE",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"E0",X"00",X"00",X"00",X"EE",X"EE",X"00",X"00",X"CE",X"DD",X"00",X"00",X"CC",X"DD",X"00",
		X"00",X"CC",X"DD",X"00",X"00",X"CC",X"DD",X"00",X"00",X"BC",X"DD",X"00",X"00",X"BC",X"DE",X"00",
		X"00",X"EB",X"EE",X"00",X"00",X"EE",X"CE",X"00",X"00",X"DD",X"CE",X"00",X"00",X"DD",X"CC",X"00",
		X"00",X"DD",X"ED",X"00",X"00",X"DD",X"ED",X"00",X"00",X"DD",X"ED",X"00",X"00",X"EE",X"CE",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EF",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"CE",X"0E",X"00",X"00",X"CE",X"ED",X"00",X"00",X"CC",X"DD",X"00",
		X"00",X"CC",X"DD",X"00",X"00",X"CC",X"DD",X"00",X"00",X"BC",X"DD",X"00",X"00",X"BC",X"DD",X"00",
		X"00",X"EE",X"DE",X"00",X"00",X"EB",X"E0",X"00",X"00",X"DD",X"E0",X"00",X"00",X"DD",X"CE",X"00",
		X"00",X"DD",X"CE",X"00",X"00",X"DD",X"ED",X"00",X"00",X"EE",X"CD",X"00",X"00",X"00",X"CD",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"CE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"CC",X"0E",X"00",X"00",X"CC",X"ED",X"00",
		X"00",X"CC",X"DD",X"00",X"00",X"BC",X"DD",X"00",X"00",X"BC",X"DD",X"00",X"00",X"EC",X"DD",X"00",
		X"00",X"EC",X"DE",X"00",X"00",X"DB",X"E0",X"00",X"00",X"DE",X"00",X"00",X"00",X"DD",X"E0",X"00",
		X"00",X"DD",X"EE",X"00",X"00",X"DD",X"DD",X"00",X"00",X"EE",X"DD",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"ED",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"CE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"FC",X"00",X"00",X"00",X"CC",X"EE",X"00",X"00",X"BC",X"ED",X"00",
		X"00",X"BC",X"DD",X"00",X"00",X"BC",X"DD",X"00",X"00",X"EB",X"DD",X"00",X"00",X"EB",X"DD",X"00",
		X"00",X"EE",X"DE",X"00",X"00",X"DE",X"E0",X"00",X"00",X"DE",X"E0",X"00",X"00",X"DD",X"E0",X"00",
		X"00",X"DD",X"CE",X"00",X"00",X"DD",X"EE",X"00",X"00",X"EE",X"DD",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"DD",X"00",X"00",X"00",X"ED",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"CE",X"00",X"00",
		X"00",X"EC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"BC",X"EE",X"00",
		X"00",X"BC",X"DE",X"00",X"00",X"BC",X"DD",X"00",X"00",X"EB",X"DD",X"00",X"00",X"EC",X"DD",X"00",
		X"00",X"DE",X"DD",X"00",X"00",X"DE",X"DE",X"00",X"00",X"DE",X"EE",X"00",X"00",X"DE",X"E0",X"00",
		X"00",X"DD",X"E0",X"00",X"00",X"DE",X"EE",X"00",X"00",X"EE",X"DD",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"DD",X"00",X"00",X"00",X"DE",X"00",X"00",X"00",X"DE",X"00",X"00",X"00",X"CE",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"EC",X"00",X"00",X"00",X"BC",X"00",X"00",X"00",X"BC",X"00",X"00",X"00",X"BC",X"00",X"00",
		X"00",X"EF",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"BC",X"00",X"00",X"00",X"BC",X"00",X"00",
		X"00",X"EB",X"00",X"00",X"00",X"EB",X"EE",X"00",X"00",X"EB",X"DD",X"00",X"00",X"EB",X"DD",X"00",
		X"00",X"DE",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DE",X"DD",X"00",X"00",X"DE",X"EE",X"00",
		X"00",X"DD",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"DE",X"00",
		X"00",X"00",X"DE",X"00",X"00",X"00",X"DE",X"00",X"00",X"00",X"E0",X"00",X"00",X"0E",X"E0",X"00",
		X"00",X"0E",X"E0",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"EB",X"00",X"00",X"00",X"EB",X"00",X"00",X"00",X"EB",X"FE",X"00",X"00",X"EB",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"EB",X"00",X"00",X"00",X"EB",X"00",X"00",X"00",X"EB",X"00",X"00",
		X"00",X"EB",X"00",X"00",X"00",X"EB",X"EE",X"00",X"00",X"EB",X"DD",X"00",X"00",X"EC",X"DD",X"00",
		X"00",X"DE",X"DD",X"00",X"00",X"EF",X"DD",X"00",X"00",X"E2",X"DD",X"00",X"00",X"DE",X"DD",X"00",
		X"00",X"DE",X"EE",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"DE",X"00",X"00",X"EE",X"E0",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",X"EF",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"0E",X"E0",X"00",X"00",X"0E",X"E0",X"00",X"00",X"0E",X"E0",X"00",
		X"00",X"0E",X"EE",X"00",X"00",X"0E",X"EE",X"00",X"00",X"0E",X"DE",X"00",X"00",X"0E",X"DE",X"00",
		X"00",X"0F",X"DE",X"00",X"00",X"0F",X"DE",X"00",X"00",X"0F",X"DE",X"00",X"00",X"0E",X"DE",X"00",
		X"00",X"0E",X"EE",X"00",X"00",X"0E",X"E0",X"00",X"00",X"0E",X"E0",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"EE",X"2E",X"00",X"00",X"E2",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",
		X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"EE",X"00",X"22",X"22",X"E3",
		X"00",X"22",X"22",X"EE",X"0E",X"22",X"22",X"EE",X"E3",X"22",X"22",X"2E",X"E3",X"22",X"22",X"2E",
		X"EE",X"22",X"22",X"2E",X"00",X"22",X"22",X"2E",X"00",X"22",X"22",X"33",X"00",X"22",X"22",X"2E",
		X"00",X"E3",X"E3",X"EE",X"00",X"3E",X"EE",X"E0",X"00",X"3E",X"EE",X"E0",X"00",X"E2",X"EE",X"E0",
		X"00",X"22",X"22",X"3E",X"00",X"22",X"22",X"EE",X"00",X"22",X"22",X"00",X"00",X"77",X"07",X"00",
		X"70",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"FE",X"00",
		X"00",X"0E",X"FF",X"00",X"00",X"EF",X"FF",X"00",X"00",X"FF",X"55",X"00",X"00",X"EF",X"EE",X"00",
		X"00",X"0E",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"E5",X"E0",X"00",X"00",X"E5",X"E0",
		X"00",X"00",X"E5",X"E0",X"00",X"EE",X"EE",X"E0",X"00",X"AE",X"EE",X"00",X"00",X"AA",X"00",X"00",
		X"0E",X"4A",X"00",X"00",X"0E",X"EA",X"00",X"00",X"E0",X"4A",X"00",X"00",X"5E",X"EE",X"00",X"00",
		X"55",X"EE",X"60",X"00",X"55",X"EE",X"00",X"00",X"E5",X"5E",X"00",X"00",X"0E",X"55",X"00",X"00",
		X"00",X"E5",X"00",X"00",X"EE",X"0E",X"00",X"00",X"ED",X"00",X"00",X"00",X"ED",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"FE",X"00",
		X"00",X"0E",X"FF",X"00",X"00",X"EF",X"FF",X"00",X"00",X"FF",X"CC",X"00",X"00",X"EF",X"EE",X"00",
		X"00",X"0E",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"EC",X"E0",X"00",X"00",X"EC",X"E0",
		X"00",X"00",X"EC",X"E0",X"00",X"EE",X"EE",X"E0",X"00",X"AE",X"EE",X"00",X"00",X"AA",X"00",X"00",
		X"0E",X"4A",X"00",X"00",X"0E",X"EA",X"00",X"00",X"E0",X"4A",X"00",X"00",X"BE",X"EE",X"00",X"00",
		X"CB",X"EE",X"60",X"00",X"CC",X"EE",X"00",X"00",X"EC",X"BE",X"00",X"00",X"0E",X"CB",X"00",X"00",
		X"00",X"EC",X"00",X"00",X"EE",X"0E",X"00",X"00",X"ED",X"00",X"00",X"00",X"ED",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"EE",X"00",
		X"E5",X"55",X"55",X"00",X"9E",X"55",X"55",X"00",X"9E",X"BB",X"BB",X"00",X"AE",X"BB",X"BB",X"00",
		X"AE",X"BB",X"BB",X"00",X"A9",X"EB",X"BB",X"00",X"2A",X"EB",X"BB",X"00",X"2A",X"EB",X"BB",X"00",
		X"2A",X"EB",X"BB",X"00",X"2A",X"EA",X"AB",X"00",X"2A",X"EA",X"AB",X"00",X"22",X"BA",X"7B",X"00",
		X"00",X"07",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"0F",X"00",X"00",X"30",X"30",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"30",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",
		X"F0",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"00",X"00",X"F0",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"32",X"00",X"00",
		X"01",X"02",X"00",X"00",X"01",X"22",X"00",X"00",X"30",X"2E",X"00",X"00",X"10",X"25",X"00",X"00",
		X"10",X"55",X"00",X"00",X"20",X"25",X"00",X"00",X"20",X"52",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"22",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"22",X"55",X"00",X"00",
		X"23",X"55",X"00",X"00",X"21",X"55",X"E0",X"00",X"01",X"E5",X"6E",X"00",X"00",X"6E",X"6E",X"00",
		X"0E",X"6E",X"E0",X"00",X"0E",X"66",X"00",X"00",X"0E",X"66",X"00",X"00",X"00",X"6E",X"00",X"00",
		X"00",X"E5",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"5E",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"0E",X"FE",X"00",X"00",X"0E",X"00",X"00",X"00",X"EF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"32",X"00",X"00",
		X"01",X"02",X"00",X"00",X"01",X"22",X"00",X"00",X"30",X"2E",X"00",X"00",X"10",X"2C",X"00",X"00",
		X"10",X"CC",X"00",X"00",X"00",X"2C",X"00",X"00",X"00",X"C2",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"22",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"03",X"CC",X"00",X"00",X"01",X"CC",X"E0",X"00",X"01",X"EC",X"DE",X"00",X"00",X"DE",X"DE",X"00",
		X"0E",X"DE",X"E0",X"00",X"0E",X"DD",X"00",X"00",X"0E",X"DD",X"00",X"00",X"00",X"DE",X"00",X"00",
		X"00",X"EC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"CE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"0E",X"FE",X"00",X"00",X"0E",X"00",X"00",X"00",X"EF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
