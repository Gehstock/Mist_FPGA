library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity h1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of h1 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"31",X"00",X"24",X"C3",X"A5",X"07",X"00",X"00",X"C3",X"41",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C3",X"4D",X"00",X"00",X"00",X"00",X"00",X"00",X"7E",X"B7",X"C8",X"35",X"AF",X"3C",X"C9",X"00",
		X"3A",X"43",X"20",X"F6",X"20",X"D3",X"00",X"C9",X"7E",X"B7",X"C8",X"35",X"C0",X"37",X"C9",X"00",
		X"DB",X"02",X"07",X"07",X"07",X"C3",X"83",X"07",X"7E",X"12",X"05",X"23",X"13",X"C2",X"38",X"00",
		X"C9",X"F5",X"AF",X"32",X"11",X"20",X"2F",X"32",X"10",X"20",X"F1",X"FB",X"C9",X"F5",X"3A",X"D0",
		X"21",X"B7",X"C2",X"58",X"00",X"F1",X"FB",X"C9",X"C5",X"D5",X"E5",X"AF",X"32",X"10",X"20",X"2F",
		X"32",X"11",X"20",X"00",X"00",X"00",X"00",X"CD",X"04",X"01",X"00",X"00",X"CD",X"39",X"01",X"CD",
		X"4C",X"07",X"CD",X"C9",X"00",X"E1",X"D1",X"C1",X"F1",X"FB",X"00",X"00",X"00",X"C9",X"21",X"28",
		X"20",X"AF",X"CD",X"91",X"00",X"77",X"21",X"3D",X"20",X"CD",X"97",X"00",X"00",X"00",X"C3",X"C9",
		X"01",X"77",X"23",X"77",X"23",X"77",X"23",X"77",X"23",X"77",X"23",X"77",X"23",X"77",X"23",X"77",
		X"23",X"C9",X"21",X"01",X"20",X"3E",X"FF",X"BE",X"CA",X"00",X"1C",X"23",X"BE",X"CA",X"0C",X"1C",
		X"23",X"BE",X"CA",X"03",X"1C",X"C3",X"0F",X"1C",X"DB",X"02",X"E6",X"30",X"FE",X"10",X"CA",X"06",
		X"1C",X"00",X"00",X"00",X"00",X"00",X"C3",X"A2",X"00",X"21",X"3D",X"20",X"DB",X"00",X"E6",X"80",
		X"CC",X"DC",X"00",X"DF",X"21",X"40",X"20",X"DF",X"CC",X"E8",X"00",X"C9",X"7E",X"B7",X"36",X"04",
		X"C0",X"CD",X"98",X"07",X"34",X"2B",X"2B",X"C9",X"3A",X"43",X"20",X"1F",X"D2",X"F7",X"00",X"3F",
		X"17",X"32",X"43",X"20",X"36",X"10",X"C9",X"2B",X"7E",X"B7",X"C8",X"35",X"23",X"3A",X"43",X"20",
		X"1F",X"C3",X"EF",X"00",X"21",X"43",X"20",X"7E",X"D3",X"00",X"23",X"23",X"23",X"23",X"7E",X"D3",
		X"04",X"C9",X"21",X"49",X"01",X"DB",X"00",X"2F",X"E6",X"3F",X"85",X"D2",X"1F",X"01",X"24",X"6F",
		X"7E",X"32",X"20",X"20",X"21",X"89",X"01",X"DB",X"01",X"00",X"00",X"2F",X"E6",X"3F",X"85",X"D2",
		X"33",X"01",X"24",X"6F",X"7E",X"32",X"21",X"20",X"C9",X"CD",X"AF",X"04",X"CD",X"6F",X"05",X"CD",
		X"72",X"04",X"CD",X"07",X"05",X"CD",X"5C",X"05",X"C9",X"DA",X"DA",X"DA",X"DA",X"DA",X"DA",X"DA",
		X"DA",X"C8",X"CE",X"DA",X"D4",X"DA",X"DA",X"DA",X"DA",X"68",X"6E",X"7A",X"74",X"92",X"8C",X"80",
		X"86",X"C2",X"BC",X"B0",X"B6",X"98",X"9E",X"AA",X"A4",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"62",X"5C",X"50",X"56",X"38",X"3E",X"4A",
		X"44",X"08",X"0E",X"1A",X"14",X"32",X"2C",X"20",X"26",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"93",X"98",X"A2",X"9D",X"B6",X"B1",X"A7",
		X"AC",X"C0",X"C0",X"C0",X"C0",X"BB",X"C0",X"C0",X"C0",X"60",X"60",X"60",X"60",X"60",X"60",X"60",
		X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"8E",X"89",X"7F",X"84",X"6B",X"70",X"7A",
		X"75",X"60",X"60",X"60",X"60",X"66",X"60",X"60",X"60",X"31",X"00",X"24",X"11",X"F0",X"3F",X"21",
		X"28",X"20",X"06",X"09",X"FF",X"21",X"3D",X"20",X"06",X"05",X"FF",X"AF",X"32",X"D0",X"21",X"32",
		X"A0",X"21",X"3E",X"0A",X"00",X"00",X"AF",X"21",X"00",X"20",X"01",X"E0",X"20",X"77",X"23",X"0D",
		X"C2",X"ED",X"01",X"05",X"C2",X"ED",X"01",X"11",X"28",X"20",X"06",X"09",X"21",X"F0",X"3F",X"FF",
		X"11",X"3D",X"20",X"06",X"05",X"FF",X"3E",X"FF",X"32",X"9F",X"20",X"21",X"40",X"06",X"11",X"43",
		X"20",X"06",X"02",X"FF",X"7E",X"32",X"47",X"20",X"23",X"11",X"0A",X"20",X"06",X"05",X"FF",X"21",
		X"90",X"07",X"F7",X"7C",X"32",X"39",X"20",X"CD",X"B7",X"07",X"21",X"4C",X"06",X"11",X"68",X"20",
		X"06",X"20",X"FF",X"21",X"0C",X"07",X"11",X"C0",X"22",X"06",X"40",X"FF",X"3E",X"FF",X"32",X"4F",
		X"20",X"32",X"22",X"20",X"32",X"C4",X"21",X"21",X"00",X"01",X"22",X"E0",X"21",X"21",X"2E",X"26",
		X"22",X"37",X"20",X"21",X"00",X"04",X"22",X"5C",X"23",X"AF",X"32",X"DE",X"22",X"32",X"EE",X"22",
		X"21",X"83",X"2A",X"22",X"8A",X"21",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"FF",X"32",
		X"01",X"20",X"32",X"D0",X"21",X"00",X"C3",X"69",X"03",X"21",X"02",X"24",X"3E",X"FF",X"06",X"1B",
		X"77",X"23",X"05",X"C2",X"80",X"02",X"2B",X"11",X"20",X"00",X"3E",X"80",X"06",X"18",X"19",X"77",
		X"05",X"C2",X"8E",X"02",X"21",X"02",X"24",X"3E",X"01",X"06",X"18",X"19",X"77",X"05",X"C2",X"9B",
		X"02",X"19",X"3E",X"FF",X"06",X"1B",X"77",X"23",X"05",X"C2",X"A6",X"02",X"11",X"18",X"03",X"21",
		X"84",X"24",X"0E",X"07",X"CD",X"D9",X"02",X"11",X"34",X"03",X"21",X"98",X"24",X"0E",X"07",X"CD",
		X"D9",X"02",X"11",X"50",X"03",X"21",X"8F",X"24",X"0E",X"05",X"CD",X"03",X"03",X"11",X"5A",X"03",
		X"21",X"6E",X"25",X"0E",X"05",X"CD",X"EE",X"02",X"C9",X"06",X"04",X"1A",X"77",X"13",X"23",X"05",
		X"C2",X"DB",X"02",X"D5",X"11",X"1C",X"00",X"19",X"D1",X"0D",X"C2",X"D9",X"02",X"C9",X"06",X"03",
		X"1A",X"77",X"13",X"23",X"05",X"C2",X"F0",X"02",X"D5",X"11",X"1D",X"00",X"19",X"D1",X"0D",X"C2",
		X"EE",X"02",X"C9",X"06",X"02",X"1A",X"77",X"13",X"23",X"05",X"C2",X"05",X"03",X"D5",X"11",X"1E",
		X"00",X"19",X"D1",X"0D",X"C2",X"03",X"03",X"C9",X"1C",X"C7",X"79",X"3E",X"A2",X"28",X"8A",X"02",
		X"82",X"20",X"8A",X"02",X"9C",X"20",X"7A",X"0E",X"A0",X"20",X"2A",X"02",X"A2",X"28",X"4A",X"02",
		X"1C",X"C7",X"89",X"3E",X"F0",X"7D",X"D1",X"07",X"40",X"10",X"5B",X"00",X"40",X"10",X"55",X"00",
		X"40",X"10",X"D1",X"01",X"40",X"10",X"51",X"00",X"40",X"10",X"51",X"00",X"40",X"7C",X"D1",X"07",
		X"A8",X"03",X"28",X"01",X"38",X"01",X"28",X"01",X"A8",X"03",X"E0",X"EE",X"EE",X"20",X"A2",X"2A",
		X"E0",X"A2",X"6E",X"80",X"A2",X"26",X"E0",X"EE",X"EA",X"C3",X"E0",X"07",X"B7",X"C2",X"5A",X"04",
		X"2A",X"94",X"20",X"22",X"90",X"20",X"2A",X"96",X"20",X"22",X"92",X"20",X"3A",X"0A",X"20",X"32",
		X"99",X"20",X"3A",X"0C",X"20",X"32",X"9A",X"20",X"3A",X"0B",X"20",X"32",X"9B",X"20",X"CD",X"AA",
		X"05",X"2A",X"B4",X"20",X"22",X"B0",X"20",X"2A",X"B6",X"20",X"22",X"B2",X"20",X"3A",X"0E",X"20",
		X"32",X"D1",X"20",X"3A",X"0D",X"20",X"32",X"D2",X"20",X"21",X"99",X"20",X"3E",X"DD",X"96",X"5F",
		X"21",X"9B",X"20",X"CD",X"6D",X"04",X"21",X"C0",X"20",X"0E",X"10",X"3A",X"D1",X"20",X"47",X"AF",
		X"80",X"F5",X"07",X"07",X"E6",X"03",X"77",X"23",X"82",X"57",X"DA",X"ED",X"03",X"1D",X"CA",X"ED",
		X"03",X"F1",X"E6",X"3F",X"0D",X"C2",X"C0",X"03",X"80",X"4F",X"07",X"07",X"E6",X"03",X"82",X"57",
		X"79",X"DA",X"EE",X"03",X"E6",X"3F",X"1D",X"C2",X"D8",X"03",X"C3",X"EE",X"03",X"F1",X"3E",X"DD",
		X"93",X"CD",X"5F",X"04",X"22",X"D3",X"20",X"21",X"9A",X"20",X"3E",X"DC",X"96",X"5F",X"21",X"C0",
		X"20",X"0E",X"10",X"3A",X"D2",X"20",X"47",X"AF",X"80",X"F5",X"0F",X"0F",X"0F",X"0F",X"E6",X"0C",
		X"B6",X"77",X"23",X"1D",X"CA",X"23",X"04",X"F1",X"E6",X"3F",X"0D",X"C2",X"08",X"04",X"1E",X"00",
		X"C3",X"24",X"04",X"F1",X"3E",X"DC",X"93",X"CD",X"5F",X"04",X"22",X"D5",X"20",X"00",X"21",X"C0",
		X"20",X"11",X"A0",X"20",X"06",X"10",X"FF",X"2A",X"D5",X"20",X"22",X"B6",X"20",X"2A",X"D3",X"20",
		X"22",X"B4",X"20",X"3A",X"99",X"20",X"CD",X"5F",X"04",X"22",X"94",X"20",X"3A",X"9A",X"20",X"CD",
		X"5F",X"04",X"22",X"96",X"20",X"3E",X"FF",X"32",X"9F",X"20",X"FB",X"00",X"C3",X"69",X"03",X"0F",
		X"0F",X"0F",X"67",X"F6",X"1F",X"6F",X"7C",X"E6",X"1F",X"C6",X"24",X"67",X"C9",X"7E",X"C6",X"84",
		X"57",X"C9",X"2A",X"90",X"20",X"7E",X"E6",X"BF",X"77",X"2A",X"92",X"20",X"7E",X"E6",X"EF",X"77",
		X"2A",X"94",X"20",X"7E",X"F6",X"40",X"77",X"2A",X"96",X"20",X"7E",X"F6",X"10",X"77",X"2A",X"B0",
		X"20",X"7E",X"E6",X"DF",X"77",X"2A",X"B2",X"20",X"7E",X"E6",X"F7",X"77",X"2A",X"B4",X"20",X"7E",
		X"F6",X"20",X"77",X"2A",X"B6",X"20",X"7E",X"F6",X"08",X"77",X"AF",X"32",X"9F",X"20",X"C9",X"3A",
		X"98",X"20",X"D3",X"07",X"D3",X"07",X"3A",X"43",X"20",X"E6",X"FD",X"D3",X"00",X"21",X"A0",X"20",
		X"7E",X"D3",X"03",X"23",X"7E",X"D3",X"0B",X"23",X"7E",X"D3",X"13",X"23",X"7E",X"D3",X"1B",X"23",
		X"7E",X"D3",X"43",X"23",X"7E",X"D3",X"4B",X"23",X"7E",X"D3",X"53",X"23",X"7E",X"D3",X"5B",X"23",
		X"7E",X"D3",X"83",X"23",X"7E",X"D3",X"8B",X"23",X"7E",X"D3",X"93",X"23",X"7E",X"D3",X"9B",X"23",
		X"7E",X"D3",X"C3",X"23",X"7E",X"D3",X"CB",X"23",X"7E",X"D3",X"D3",X"23",X"7E",X"D3",X"DB",X"3A",
		X"43",X"20",X"F6",X"02",X"D3",X"00",X"C9",X"21",X"1E",X"20",X"3A",X"31",X"20",X"07",X"D2",X"12",
		X"05",X"34",X"21",X"32",X"20",X"35",X"F0",X"34",X"23",X"7E",X"B7",X"CA",X"24",X"05",X"35",X"21",
		X"1E",X"20",X"34",X"C9",X"3A",X"23",X"20",X"0F",X"0F",X"0F",X"E6",X"1F",X"11",X"2E",X"06",X"83",
		X"D2",X"34",X"05",X"14",X"5F",X"1A",X"E6",X"07",X"77",X"2B",X"1A",X"0F",X"0F",X"0F",X"E6",X"0F",
		X"77",X"2B",X"1A",X"77",X"E6",X"71",X"C0",X"C3",X"1F",X"05",X"21",X"39",X"20",X"7E",X"B7",X"C8",
		X"3D",X"77",X"E6",X"0F",X"FE",X"0F",X"C0",X"7E",X"D6",X"06",X"77",X"C9",X"3A",X"22",X"20",X"B7",
		X"C8",X"3A",X"6B",X"20",X"D6",X"60",X"D2",X"6B",X"05",X"3E",X"00",X"32",X"23",X"20",X"C9",X"11",
		X"06",X"06",X"21",X"00",X"00",X"39",X"22",X"95",X"21",X"3A",X"1E",X"20",X"4F",X"06",X"14",X"26",
		X"04",X"1A",X"81",X"6F",X"29",X"F9",X"E1",X"36",X"80",X"E1",X"36",X"80",X"13",X"05",X"C2",X"7F",
		X"05",X"06",X"14",X"26",X"04",X"1A",X"81",X"6F",X"29",X"F9",X"E1",X"36",X"00",X"E1",X"36",X"00",
		X"13",X"05",X"C2",X"93",X"05",X"2A",X"95",X"21",X"F9",X"C9",X"47",X"3A",X"99",X"20",X"D6",X"80",
		X"FA",X"F2",X"05",X"4F",X"3A",X"BF",X"21",X"B7",X"CA",X"CA",X"05",X"79",X"2F",X"4F",X"21",X"47",
		X"20",X"7E",X"91",X"5F",X"F2",X"D3",X"05",X"C3",X"EB",X"05",X"21",X"47",X"20",X"7E",X"91",X"5F",
		X"FA",X"EB",X"05",X"7E",X"D6",X"08",X"57",X"7B",X"CD",X"FC",X"05",X"FE",X"08",X"D2",X"E1",X"05",
		X"51",X"72",X"7E",X"CD",X"FC",X"05",X"80",X"32",X"98",X"20",X"C9",X"7E",X"C6",X"08",X"57",X"C3",
		X"D7",X"05",X"78",X"32",X"98",X"20",X"3E",X"00",X"32",X"47",X"20",X"C9",X"C6",X"80",X"D2",X"03",
		X"06",X"2F",X"3C",X"D6",X"80",X"C9",X"04",X"10",X"30",X"3C",X"44",X"5C",X"66",X"70",X"78",X"A0",
		X"A7",X"B5",X"C4",X"E0",X"E7",X"F0",X"F7",X"04",X"04",X"04",X"01",X"07",X"20",X"34",X"40",X"54",
		X"60",X"6C",X"74",X"88",X"A4",X"B0",X"BD",X"D0",X"E3",X"EC",X"F4",X"01",X"01",X"01",X"87",X"87",
		X"87",X"87",X"8B",X"89",X"99",X"B8",X"0D",X"0B",X"13",X"09",X"19",X"21",X"79",X"79",X"79",X"79",
		X"0E",X"01",X"00",X"40",X"20",X"50",X"20",X"80",X"00",X"00",X"00",X"00",X"80",X"D0",X"80",X"D0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"80",X"11",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"B0",X"20",
		X"B0",X"20",X"00",X"10",X"F0",X"30",X"F0",X"30",X"01",X"01",X"02",X"04",X"01",X"01",X"68",X"38",
		X"00",X"10",X"20",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0B",X"00",X"C0",X"20",X"C0",X"20",X"80",X"10",X"F0",X"30",X"F0",X"30",
		X"01",X"01",X"02",X"03",X"01",X"01",X"68",X"38",X"80",X"10",X"30",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"C0",X"20",
		X"C0",X"20",X"00",X"11",X"F0",X"30",X"F0",X"30",X"01",X"01",X"04",X"02",X"01",X"01",X"70",X"38",
		X"00",X"11",X"40",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"00",X"C0",X"20",X"C0",X"20",X"80",X"13",X"F0",X"30",X"F0",X"30",
		X"01",X"01",X"06",X"01",X"01",X"01",X"78",X"38",X"80",X"13",X"50",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"01",X"01",X"FC",X"D0",X"30",X"00",X"13",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"01",X"01",X"02",X"D0",X"10",X"00",X"13",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"01",X"01",X"02",X"D0",X"10",X"00",X"13",X"00",X"00",X"00",X"08",X"0C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"4F",X"20",X"AF",
		X"BE",X"CA",X"6E",X"07",X"77",X"21",X"12",X"20",X"34",X"CD",X"B8",X"00",X"CD",X"74",X"07",X"3E",
		X"FF",X"32",X"4F",X"20",X"21",X"65",X"20",X"7E",X"23",X"77",X"2B",X"36",X"00",X"C9",X"3E",X"FF",
		X"32",X"65",X"20",X"C9",X"21",X"A0",X"21",X"7E",X"D3",X"01",X"23",X"7E",X"D3",X"09",X"23",X"7E",
		X"D3",X"11",X"C9",X"E6",X"06",X"85",X"D2",X"8A",X"07",X"24",X"6F",X"5E",X"23",X"56",X"EB",X"C9",
		X"00",X"45",X"00",X"60",X"00",X"75",X"00",X"90",X"23",X"34",X"23",X"E5",X"CD",X"A1",X"07",X"E1",
		X"C9",X"CD",X"2D",X"50",X"C9",X"DB",X"02",X"E6",X"30",X"FE",X"10",X"CA",X"09",X"1C",X"FE",X"20",
		X"CA",X"23",X"5C",X"FB",X"C3",X"7E",X"00",X"CD",X"26",X"5C",X"B7",X"CA",X"AC",X"02",X"C3",X"79",
		X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"21",X"00",X"00",X"39",X"7C",X"FE",X"24",X"C2",X"00",X"00",X"7D",X"FE",X"00",X"C2",X"00",X"00",
		X"D3",X"02",X"3A",X"9F",X"20",X"C3",X"6C",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
