library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity tn04 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of tn04 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"58",X"10",X"00",X"90",X"31",X"0C",X"06",X"D0",X"38",X"08",X"00",X"D0",X"38",X"08",X"00",X"D0",
		X"38",X"04",X"07",X"D0",X"48",X"05",X"06",X"C8",X"50",X"04",X"05",X"BE",X"4E",X"08",X"00",X"B8",
		X"38",X"0C",X"06",X"B0",X"38",X"08",X"00",X"B0",X"38",X"04",X"07",X"B0",X"48",X"05",X"06",X"A8",
		X"50",X"04",X"05",X"9E",X"4E",X"08",X"00",X"98",X"38",X"0C",X"09",X"90",X"59",X"0C",X"0E",X"A6",
		X"67",X"08",X"00",X"98",X"60",X"0B",X"06",X"A6",X"78",X"0A",X"00",X"90",X"78",X"0B",X"06",X"A6",
		X"90",X"0A",X"00",X"90",X"90",X"0C",X"06",X"A6",X"A8",X"0A",X"00",X"A6",X"A8",X"0C",X"06",X"A6",
		X"BC",X"0B",X"00",X"90",X"A8",X"0C",X"06",X"A6",X"C0",X"0A",X"00",X"A6",X"C0",X"0C",X"06",X"A6",
		X"D4",X"0B",X"00",X"90",X"C0",X"0C",X"06",X"A6",X"D8",X"0C",X"07",X"A6",X"D8",X"0C",X"06",X"A6",
		X"F0",X"00",X"00",X"00",X"00",X"92",X"18",X"01",X"04",X"E1",X"17",X"00",X"00",X"00",X"00",X"00",
		X"17",X"00",X"1E",X"1E",X"1E",X"1E",X"FF",X"FF",X"FF",X"FF",X"36",X"00",X"CD",X"DC",X"18",X"3E",
		X"04",X"CD",X"FB",X"01",X"2A",X"33",X"20",X"CD",X"76",X"03",X"0E",X"05",X"E5",X"C5",X"11",X"D0",
		X"19",X"D5",X"06",X"02",X"C5",X"E5",X"01",X"12",X"02",X"CD",X"D5",X"01",X"3E",X"05",X"CD",X"D5",
		X"14",X"E1",X"C1",X"05",X"C2",X"B4",X"18",X"D1",X"C1",X"E1",X"0D",X"C2",X"AC",X"18",X"01",X"12",
		X"02",X"CD",X"8C",X"08",X"CD",X"C1",X"00",X"3E",X"04",X"C3",X"04",X"02",X"21",X"2F",X"20",X"36",
		X"00",X"2E",X"14",X"36",X"00",X"C9",X"3A",X"17",X"20",X"A7",X"3E",X"02",X"C2",X"FB",X"01",X"C3",
		X"04",X"02",X"3A",X"1D",X"20",X"A7",X"3E",X"01",X"C3",X"EC",X"18",X"3A",X"27",X"20",X"A7",X"3E",
		X"08",X"C3",X"EC",X"18",X"3A",X"91",X"20",X"A7",X"3E",X"08",X"C3",X"EC",X"18",X"3E",X"DF",X"CD",
		X"04",X"02",X"3E",X"DF",X"C3",X"17",X"02",X"3A",X"E4",X"20",X"A7",X"C8",X"3A",X"54",X"20",X"A7",
		X"3E",X"01",X"C2",X"0E",X"02",X"C3",X"17",X"02",X"CD",X"95",X"19",X"D8",X"CD",X"5F",X"0C",X"CD",
		X"47",X"0B",X"CD",X"17",X"19",X"C3",X"92",X"15",X"CD",X"C2",X"07",X"CD",X"95",X"19",X"D8",X"CD",
		X"81",X"09",X"CD",X"F1",X"0E",X"CD",X"4B",X"19",X"C3",X"A2",X"14",X"CD",X"5A",X"19",X"21",X"34",
		X"20",X"7E",X"2E",X"7F",X"BE",X"D8",X"C6",X"08",X"77",X"C9",X"21",X"34",X"20",X"7E",X"2E",X"7D",
		X"BE",X"D0",X"D6",X"08",X"77",X"C9",X"CD",X"79",X"19",X"CD",X"95",X"19",X"D8",X"CD",X"5F",X"0C",
		X"CD",X"9C",X"09",X"CD",X"DB",X"16",X"C3",X"6C",X"0F",X"3A",X"05",X"20",X"A7",X"3E",X"04",X"C2",
		X"0E",X"02",X"C3",X"17",X"02",X"CD",X"95",X"19",X"D8",X"CD",X"BC",X"09",X"CD",X"E2",X"0F",X"CD",
		X"56",X"0D",X"C3",X"9C",X"16",X"3A",X"7B",X"20",X"0F",X"C9",X"CD",X"71",X"03",X"C5",X"E5",X"1A",
		X"D3",X"04",X"DB",X"03",X"A6",X"CA",X"AD",X"19",X"3E",X"01",X"32",X"11",X"20",X"DB",X"03",X"AE",
		X"77",X"23",X"13",X"AF",X"D3",X"04",X"DB",X"03",X"A6",X"CA",X"C1",X"19",X"3E",X"01",X"32",X"11",
		X"20",X"DB",X"03",X"AE",X"77",X"E1",X"01",X"20",X"00",X"09",X"C1",X"05",X"C2",X"9D",X"19",X"C9",
		X"00",X"00",X"07",X"00",X"00",X"00",X"42",X"00",X"00",X"00",X"15",X"02",X"11",X"49",X"8F",X"00",
		X"EF",X"05",X"2F",X"08",X"D1",X"21",X"1D",X"20",X"00",X"00",X"17",X"00",X"09",X"11",X"07",X"00",
		X"07",X"00",X"47",X"00",X"00",X"02",X"21",X"40",X"49",X"10",X"05",X"00",X"00",X"80",X"01",X"08",
		X"09",X"40",X"07",X"00",X"03",X"00",X"01",X"00",X"49",X"02",X"49",X"44",X"00",X"80",X"09",X"02",
		X"00",X"40",X"87",X"08",X"02",X"00",X"03",X"00",X"DB",X"02",X"E6",X"03",X"21",X"27",X"21",X"F5",
		X"86",X"77",X"F1",X"2E",X"27",X"26",X"22",X"86",X"77",X"C9",X"CD",X"44",X"1A",X"7E",X"3D",X"C8",
		X"4F",X"21",X"01",X"25",X"11",X"26",X"40",X"C5",X"01",X"10",X"01",X"CD",X"D5",X"01",X"C1",X"0D",
		X"C2",X"34",X"1A",X"C9",X"CD",X"52",X"1A",X"2E",X"27",X"7E",X"C9",X"CD",X"52",X"1A",X"2E",X"25",
		X"7E",X"C9",X"3A",X"DB",X"20",X"0F",X"DA",X"5C",X"1A",X"26",X"21",X"C9",X"26",X"22",X"C9",X"3E",
		X"50",X"32",X"C2",X"20",X"C3",X"8C",X"02",X"3E",X"01",X"32",X"C1",X"20",X"C3",X"8C",X"02",X"21",
		X"01",X"50",X"22",X"C1",X"20",X"C3",X"8C",X"02",X"21",X"29",X"09",X"11",X"36",X"21",X"06",X"06",
		X"C3",X"8B",X"03",X"21",X"2F",X"09",X"C3",X"7B",X"1A",X"21",X"12",X"20",X"AF",X"BE",X"3E",X"10",
		X"CA",X"04",X"02",X"35",X"C3",X"FB",X"01",X"21",X"E9",X"20",X"3A",X"DB",X"20",X"0F",X"D0",X"23",
		X"C9",X"CD",X"97",X"1A",X"AF",X"BE",X"C8",X"CD",X"52",X"1A",X"21",X"C4",X"20",X"D2",X"B2",X"1A",
		X"2E",X"C7",X"7E",X"06",X"15",X"B8",X"D8",X"CD",X"44",X"1A",X"34",X"CD",X"2A",X"1A",X"CD",X"97",
		X"1A",X"36",X"00",X"21",X"12",X"20",X"36",X"50",X"C9",X"FE",X"FF",X"CA",X"25",X"1B",X"FE",X"FE",
		X"CA",X"1A",X"1B",X"21",X"3B",X"21",X"36",X"80",X"23",X"77",X"23",X"EB",X"21",X"5D",X"1B",X"87",
		X"4F",X"06",X"00",X"09",X"7E",X"23",X"66",X"6F",X"C3",X"F9",X"1A",X"3A",X"3B",X"21",X"A7",X"C8",
		X"21",X"3D",X"21",X"35",X"C0",X"EB",X"2A",X"3E",X"21",X"7E",X"A7",X"CA",X"25",X"1B",X"FE",X"FF",
		X"CA",X"14",X"1B",X"12",X"23",X"7E",X"06",X"08",X"D3",X"01",X"07",X"05",X"C2",X"08",X"1B",X"23",
		X"22",X"3E",X"21",X"C9",X"3A",X"3C",X"21",X"F2",X"D3",X"1A",X"3E",X"01",X"32",X"3D",X"21",X"3E",
		X"80",X"32",X"3B",X"21",X"C9",X"3E",X"FF",X"06",X"08",X"D3",X"01",X"07",X"05",X"C2",X"29",X"1B",
		X"AF",X"32",X"3B",X"21",X"C9",X"21",X"39",X"21",X"7E",X"3D",X"77",X"C0",X"2B",X"7E",X"23",X"77",
		X"23",X"7E",X"A7",X"C2",X"49",X"1B",X"C3",X"EB",X"1A",X"3A",X"36",X"21",X"CD",X"C9",X"1A",X"AF",
		X"32",X"3A",X"21",X"C9",X"AF",X"32",X"37",X"21",X"3C",X"32",X"3A",X"21",X"C9",X"08",X"45",X"9C",
		X"45",X"C6",X"45",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
