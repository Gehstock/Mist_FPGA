-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

entity CATACOMB_1H is
  port (
    CLK         : in    std_logic;
    ADDR        : in    std_logic_vector(10 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of CATACOMB_1H is


  type ROM_ARRAY is array(0 to 2047) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"38",x"7C",x"C2",x"82",x"86",x"7C",x"38",x"00", -- 0x0000
    x"02",x"02",x"FE",x"FE",x"42",x"02",x"00",x"00", -- 0x0008
    x"62",x"F2",x"BA",x"9A",x"9E",x"CE",x"46",x"00", -- 0x0010
    x"8C",x"DE",x"F2",x"B2",x"92",x"86",x"04",x"00", -- 0x0018
    x"08",x"FE",x"FE",x"C8",x"68",x"38",x"18",x"00", -- 0x0020
    x"1C",x"BE",x"A2",x"A2",x"A2",x"E6",x"E4",x"00", -- 0x0028
    x"0C",x"9E",x"92",x"92",x"D2",x"7E",x"3C",x"00", -- 0x0030
    x"C0",x"E0",x"B0",x"9E",x"8E",x"C0",x"C0",x"00", -- 0x0038
    x"0C",x"6E",x"9A",x"9A",x"B2",x"F2",x"6C",x"00", -- 0x0040
    x"78",x"FC",x"96",x"92",x"92",x"F2",x"60",x"00", -- 0x0048
    x"CF",x"0F",x"0F",x"0F",x"0F",x"0E",x"0C",x"08", -- 0x0050
    x"08",x"0C",x"0E",x"0E",x"0F",x"0F",x"0F",x"8F", -- 0x0058
    x"00",x"00",x"00",x"18",x"18",x"00",x"00",x"00", -- 0x0060
    x"18",x"28",x"38",x"2C",x"38",x"28",x"18",x"00", -- 0x0068
    x"40",x"20",x"10",x"08",x"04",x"02",x"00",x"00", -- 0x0070
    x"80",x"90",x"90",x"90",x"90",x"FE",x"FE",x"00", -- 0x0078
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0080
    x"3E",x"7E",x"C8",x"88",x"C8",x"7E",x"3E",x"00", -- 0x0088
    x"6C",x"FE",x"92",x"92",x"92",x"FE",x"FE",x"00", -- 0x0090
    x"44",x"C6",x"82",x"82",x"C6",x"7C",x"38",x"00", -- 0x0098
    x"38",x"7C",x"C6",x"82",x"82",x"FE",x"FE",x"00", -- 0x00A0
    x"82",x"92",x"92",x"92",x"FE",x"FE",x"00",x"00", -- 0x00A8
    x"80",x"90",x"90",x"90",x"90",x"FE",x"FE",x"00", -- 0x00B0
    x"9E",x"9E",x"92",x"82",x"C6",x"7C",x"38",x"00", -- 0x00B8
    x"FE",x"FE",x"10",x"10",x"10",x"FE",x"FE",x"00", -- 0x00C0
    x"82",x"82",x"FE",x"FE",x"82",x"82",x"00",x"00", -- 0x00C8
    x"FC",x"FE",x"02",x"02",x"02",x"06",x"04",x"00", -- 0x00D0
    x"82",x"C6",x"6E",x"3C",x"18",x"FE",x"FE",x"00", -- 0x00D8
    x"02",x"02",x"02",x"02",x"FE",x"FE",x"00",x"00", -- 0x00E0
    x"FE",x"FE",x"70",x"38",x"70",x"FE",x"FE",x"00", -- 0x00E8
    x"FE",x"FE",x"1C",x"38",x"70",x"FE",x"FE",x"00", -- 0x00F0
    x"7C",x"FE",x"82",x"82",x"82",x"FE",x"7C",x"00", -- 0x00F8
    x"70",x"F8",x"88",x"88",x"88",x"FE",x"FE",x"00", -- 0x0100
    x"7A",x"FC",x"8E",x"8A",x"82",x"FE",x"7C",x"00", -- 0x0108
    x"72",x"F6",x"9E",x"8C",x"88",x"FE",x"FE",x"00", -- 0x0110
    x"0C",x"5E",x"D2",x"92",x"92",x"F6",x"64",x"00", -- 0x0118
    x"80",x"80",x"FE",x"FE",x"80",x"80",x"00",x"00", -- 0x0120
    x"FC",x"FE",x"02",x"02",x"02",x"FE",x"FC",x"00", -- 0x0128
    x"F0",x"F8",x"1C",x"0E",x"1C",x"F8",x"F0",x"00", -- 0x0130
    x"F8",x"FE",x"1C",x"38",x"1C",x"FE",x"F8",x"00", -- 0x0138
    x"C6",x"EE",x"7C",x"38",x"7C",x"EE",x"C6",x"00", -- 0x0140
    x"C0",x"F0",x"1E",x"1E",x"F0",x"C0",x"00",x"00", -- 0x0148
    x"C2",x"E2",x"F2",x"BA",x"9E",x"8E",x"86",x"00", -- 0x0150
    x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00", -- 0x0158
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0160
    x"0D",x"53",x"31",x"19",x"08",x"04",x"F2",x"00", -- 0x0168
    x"3C",x"42",x"A5",x"A5",x"A5",x"99",x"42",x"3C", -- 0x0170
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0178
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0180
    x"00",x"00",x"00",x"00",x"03",x"07",x"07",x"7B", -- 0x0188
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0190
    x"07",x"07",x"03",x"00",x"00",x"00",x"00",x"00", -- 0x0198
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01B8
    x"F0",x"10",x"30",x"60",x"C0",x"C0",x"60",x"E0", -- 0x01C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01C8
    x"01",x"01",x"01",x"01",x"02",x"03",x"01",x"01", -- 0x01D0
    x"18",x"3C",x"7E",x"FF",x"3C",x"3C",x"3C",x"3C", -- 0x01D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01E0
    x"40",x"60",x"40",x"60",x"40",x"60",x"40",x"60", -- 0x01E8
    x"3C",x"42",x"81",x"A5",x"A5",x"99",x"42",x"3C", -- 0x01F0
    x"FF",x"9F",x"9F",x"9F",x"FF",x"91",x"91",x"91", -- 0x01F8
    x"80",x"40",x"20",x"10",x"00",x"02",x"26",x"24", -- 0x0200
    x"00",x"00",x"00",x"00",x"01",x"41",x"63",x"2F", -- 0x0208
    x"24",x"27",x"03",x"00",x"10",x"20",x"40",x"80", -- 0x0210
    x"2F",x"E3",x"C1",x"01",x"00",x"00",x"00",x"00", -- 0x0218
    x"07",x"08",x"08",x"08",x"07",x"00",x"07",x"08", -- 0x0220
    x"C0",x"20",x"20",x"20",x"C0",x"00",x"C0",x"20", -- 0x0228
    x"08",x"08",x"07",x"00",x"00",x"0F",x"04",x"00", -- 0x0230
    x"20",x"20",x"C0",x"00",x"20",x"E0",x"20",x"00", -- 0x0238
    x"07",x"08",x"08",x"07",x"00",x"07",x"08",x"08", -- 0x0240
    x"C0",x"20",x"20",x"C0",x"00",x"C0",x"20",x"20", -- 0x0248
    x"07",x"00",x"06",x"09",x"08",x"08",x"04",x"00", -- 0x0250
    x"C0",x"00",x"20",x"20",x"A0",x"60",x"20",x"00", -- 0x0258
    x"07",x"08",x"08",x"07",x"00",x"07",x"08",x"08", -- 0x0260
    x"C0",x"20",x"20",x"C0",x"00",x"C0",x"20",x"20", -- 0x0268
    x"07",x"00",x"07",x"09",x"09",x"08",x"04",x"00", -- 0x0270
    x"C0",x"00",x"C0",x"20",x"20",x"20",x"40",x"00", -- 0x0278
    x"01",x"07",x"1F",x"3F",x"3F",x"7F",x"7F",x"FF", -- 0x0280
    x"80",x"E0",x"F0",x"F8",x"F8",x"FC",x"FC",x"FE", -- 0x0288
    x"FF",x"7F",x"7F",x"3F",x"3F",x"1F",x"07",x"01", -- 0x0290
    x"FE",x"FC",x"FC",x"F8",x"F8",x"F0",x"E0",x"80", -- 0x0298
    x"01",x"03",x"03",x"03",x"03",x"03",x"03",x"03", -- 0x02A0
    x"80",x"C0",x"C0",x"C0",x"CE",x"D0",x"E0",x"E0", -- 0x02A8
    x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"01", -- 0x02B0
    x"E0",x"E0",x"D0",x"CE",x"C0",x"C0",x"C0",x"80", -- 0x02B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"0F", -- 0x02C0
    x"00",x"07",x"0F",x"1F",x"00",x"00",x"FF",x"FF", -- 0x02C8
    x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02D0
    x"FF",x"00",x"00",x"1F",x"0F",x"07",x"00",x"00", -- 0x02D8
    x"00",x"00",x"00",x"00",x"01",x"00",x"07",x"F8", -- 0x02E0
    x"00",x"00",x"00",x"00",x"C0",x"1C",x"FA",x"03", -- 0x02E8
    x"07",x"00",x"01",x"00",x"00",x"00",x"00",x"00", -- 0x02F0
    x"FA",x"1C",x"C0",x"00",x"00",x"00",x"00",x"00", -- 0x02F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"00", -- 0x0300
    x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E4", -- 0x0308
    x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0310
    x"E4",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0", -- 0x0318
    x"0F",x"07",x"07",x"07",x"07",x"07",x"07",x"07", -- 0x0320
    x"F0",x"80",x"C0",x"E0",x"F0",x"F8",x"F8",x"F8", -- 0x0328
    x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"0F", -- 0x0330
    x"F8",x"F8",x"F8",x"F0",x"E0",x"C0",x"80",x"F0", -- 0x0338
    x"0F",x"01",x"01",x"01",x"01",x"01",x"01",x"07", -- 0x0340
    x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"8F", -- 0x0348
    x"07",x"01",x"01",x"01",x"01",x"01",x"01",x"0F", -- 0x0350
    x"8F",x"00",x"00",x"00",x"00",x"00",x"00",x"E0", -- 0x0358
    x"01",x"07",x"1F",x"3F",x"3F",x"7F",x"7F",x"FF", -- 0x0360
    x"80",x"E0",x"F0",x"F8",x"F8",x"FC",x"FC",x"FE", -- 0x0368
    x"FF",x"7F",x"7F",x"3F",x"3F",x"1F",x"07",x"01", -- 0x0370
    x"FE",x"FC",x"FC",x"F8",x"F8",x"F0",x"E0",x"80", -- 0x0378
    x"00",x"00",x"0D",x"16",x"15",x"1B",x"3E",x"35", -- 0x0380
    x"00",x"E0",x"50",x"FC",x"AE",x"57",x"AB",x"F5", -- 0x0388
    x"6B",x"5E",x"75",x"2B",x"3D",x"16",x"0C",x"00", -- 0x0390
    x"5D",x"AB",x"F6",x"6E",x"DA",x"34",x"18",x"00", -- 0x0398
    x"00",x"00",x"00",x"00",x"01",x"00",x"07",x"F8", -- 0x03A0
    x"00",x"00",x"00",x"01",x"C6",x"1E",x"FC",x"10", -- 0x03A8
    x"07",x"00",x"01",x"00",x"00",x"00",x"00",x"00", -- 0x03B0
    x"E0",x"00",x"C0",x"00",x"00",x"00",x"00",x"00", -- 0x03B8
    x"00",x"00",x"00",x"00",x"01",x"00",x"07",x"F8", -- 0x03C0
    x"00",x"00",x"00",x"00",x"C0",x"00",x"F0",x"1C", -- 0x03C8
    x"07",x"00",x"01",x"00",x"00",x"00",x"00",x"00", -- 0x03D0
    x"FE",x"03",x"C0",x"00",x"00",x"00",x"00",x"00", -- 0x03D8
    x"0A",x"1B",x"39",x"4D",x"4C",x"FA",x"FE",x"CA", -- 0x03E0
    x"01",x"E3",x"DD",x"00",x"38",x"FC",x"E1",x"E3", -- 0x03E8
    x"CA",x"FE",x"FA",x"4C",x"4D",x"39",x"1B",x"0A", -- 0x03F0
    x"E3",x"FD",x"3C",x"38",x"00",x"C1",x"E3",x"1D", -- 0x03F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0400
    x"81",x"81",x"81",x"81",x"81",x"81",x"81",x"FF", -- 0x0408
    x"81",x"81",x"81",x"81",x"81",x"81",x"81",x"81", -- 0x0410
    x"FF",x"81",x"81",x"81",x"81",x"81",x"81",x"81", -- 0x0418
    x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01", -- 0x0420
    x"00",x"00",x"00",x"00",x"80",x"80",x"C0",x"C0", -- 0x0428
    x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0430
    x"80",x"C0",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0438
    x"02",x"03",x"00",x"00",x"03",x"03",x"02",x"02", -- 0x0440
    x"E0",x"F0",x"F0",x"F0",x"B0",x"F0",x"B0",x"B0", -- 0x0448
    x"07",x"07",x"07",x"03",x"03",x"00",x"00",x"00", -- 0x0450
    x"F0",x"B0",x"B0",x"F0",x"B0",x"A0",x"E0",x"C0", -- 0x0458
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01", -- 0x0460
    x"00",x"00",x"00",x"00",x"00",x"40",x"C0",x"C0", -- 0x0468
    x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0470
    x"80",x"80",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0478
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01", -- 0x0480
    x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"C0", -- 0x0488
    x"03",x"01",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0490
    x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0498
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02", -- 0x04A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"C0", -- 0x04A8
    x"03",x"02",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04B0
    x"F0",x"C0",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04B8
    x"0A",x"1B",x"39",x"4D",x"7C",x"CA",x"CA",x"FE", -- 0x04C0
    x"00",x"F8",x"C7",x"00",x"20",x"30",x"F0",x"F8", -- 0x04C8
    x"FE",x"CA",x"CA",x"7C",x"4D",x"3D",x"1B",x"0A", -- 0x04D0
    x"F8",x"F7",x"30",x"20",x"00",x"C0",x"F8",x"07", -- 0x04D8
    x"0F",x"09",x"01",x"03",x"01",x"01",x"02",x"02", -- 0x04E0
    x"78",x"48",x"40",x"80",x"E0",x"60",x"A0",x"80", -- 0x04E8
    x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04F0
    x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00", -- 0x04F8
    x"00",x"01",x"01",x"01",x"01",x"00",x"02",x"07", -- 0x0500
    x"80",x"C0",x"E0",x"E0",x"E0",x"C0",x"E0",x"D0", -- 0x0508
    x"06",x"26",x"3F",x"06",x"01",x"01",x"01",x"01", -- 0x0510
    x"C0",x"E0",x"C0",x"D0",x"E0",x"40",x"20",x"80", -- 0x0518
    x"0F",x"09",x"01",x"01",x"03",x"01",x"07",x"03", -- 0x0520
    x"78",x"48",x"40",x"E0",x"A0",x"E0",x"40",x"C0", -- 0x0528
    x"01",x"01",x"01",x"01",x"00",x"02",x"00",x"00", -- 0x0530
    x"C0",x"80",x"40",x"00",x"00",x"00",x"00",x"00", -- 0x0538
    x"00",x"01",x"01",x"01",x"03",x"00",x"07",x"04", -- 0x0540
    x"80",x"C0",x"C0",x"C0",x"E0",x"C0",x"D0",x"F0", -- 0x0548
    x"04",x"07",x"04",x"00",x"03",x"01",x"03",x"07", -- 0x0550
    x"D0",x"D0",x"F0",x"C0",x"E0",x"C0",x"E0",x"F0", -- 0x0558
    x"0F",x"09",x"01",x"01",x"00",x"03",x"03",x"01", -- 0x0560
    x"78",x"48",x"00",x"C0",x"E0",x"A0",x"C0",x"40", -- 0x0568
    x"01",x"00",x"00",x"01",x"01",x"00",x"00",x"00", -- 0x0570
    x"C0",x"80",x"C0",x"60",x"20",x"40",x"00",x"00", -- 0x0578
    x"00",x"01",x"01",x"01",x"03",x"03",x"04",x"04", -- 0x0580
    x"80",x"C0",x"C0",x"C0",x"E0",x"E0",x"D0",x"D0", -- 0x0588
    x"07",x"04",x"04",x"03",x"02",x"01",x"03",x"07", -- 0x0590
    x"F0",x"D0",x"C0",x"E0",x"E0",x"C0",x"E0",x"F0", -- 0x0598
    x"0F",x"09",x"01",x"01",x"03",x"01",x"02",x"01", -- 0x05A0
    x"78",x"48",x"00",x"C0",x"E0",x"80",x"C0",x"00", -- 0x05A8
    x"01",x"01",x"02",x"01",x"01",x"01",x"00",x"00", -- 0x05B0
    x"C0",x"C0",x"80",x"80",x"00",x"00",x"80",x"80", -- 0x05B8
    x"00",x"01",x"01",x"01",x"03",x"00",x"04",x"07", -- 0x05C0
    x"80",x"C0",x"C0",x"C0",x"E0",x"C0",x"F0",x"D0", -- 0x05C8
    x"04",x"04",x"07",x"00",x"01",x"01",x"03",x"07", -- 0x05D0
    x"D0",x"F0",x"D0",x"C0",x"E0",x"40",x"60",x"70", -- 0x05D8
    x"0A",x"1B",x"39",x"4D",x"7C",x"CA",x"CA",x"FE", -- 0x05E0
    x"03",x"C7",x"EB",x"00",x"3F",x"3F",x"C7",x"C7", -- 0x05E8
    x"FE",x"CA",x"CA",x"7C",x"4D",x"39",x"1B",x"0A", -- 0x05F0
    x"C7",x"FF",x"3F",x"3F",x"00",x"C3",x"C7",x"3B", -- 0x05F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0600
    x"B6",x"6D",x"DB",x"B6",x"6D",x"DB",x"B6",x"6D", -- 0x0608
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0610
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0618
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF", -- 0x0620
    x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF", -- 0x0628
    x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF", -- 0x0630
    x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF", -- 0x0638
    x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0640
    x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0648
    x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0650
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0658
    x"01",x"03",x"04",x"03",x"27",x"3E",x"6C",x"F8", -- 0x0660
    x"86",x"CF",x"2F",x"C6",x"E0",x"70",x"36",x"1F", -- 0x0668
    x"FE",x"6F",x"3F",x"27",x"03",x"04",x"03",x"01", -- 0x0670
    x"7F",x"F6",x"F0",x"E0",x"C6",x"2F",x"CF",x"86", -- 0x0678
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0680
    x"E7",x"24",x"24",x"3C",x"3C",x"24",x"24",x"E7", -- 0x0688
    x"00",x"70",x"F0",x"9B",x"8B",x"C0",x"60",x"00", -- 0x0690
    x"FF",x"D3",x"81",x"C9",x"82",x"91",x"CB",x"F3", -- 0x0698
    x"00",x"00",x"00",x"01",x"01",x"03",x"04",x"06", -- 0x06A0
    x"80",x"80",x"00",x"00",x"80",x"C0",x"C0",x"A0", -- 0x06A8
    x"15",x"0B",x"0D",x"0F",x"02",x"07",x"01",x"01", -- 0x06B0
    x"88",x"78",x"F8",x"B0",x"E0",x"B0",x"E0",x"40", -- 0x06B8
    x"00",x"02",x"03",x"0E",x"16",x"23",x"17",x"0C", -- 0x06C0
    x"48",x"B0",x"20",x"44",x"98",x"20",x"A0",x"C0", -- 0x06C8
    x"0F",x"0C",x"17",x"23",x"16",x"0F",x"02",x"02", -- 0x06D0
    x"C0",x"C0",x"A0",x"20",x"98",x"44",x"B0",x"48", -- 0x06D8
    x"00",x"1D",x"0F",x"07",x"07",x"0F",x"0F",x"0F", -- 0x06E0
    x"00",x"C0",x"80",x"00",x"00",x"80",x"80",x"C0", -- 0x06E8
    x"1F",x"1F",x"1F",x"03",x"09",x"0F",x"00",x"00", -- 0x06F0
    x"C0",x"C0",x"40",x"00",x"00",x"00",x"00",x"00", -- 0x06F8
    x"20",x"10",x"08",x"04",x"04",x"41",x"03",x"01", -- 0x0700
    x"00",x"00",x"01",x"02",x"1C",x"80",x"A2",x"60", -- 0x0708
    x"06",x"13",x"20",x"40",x"00",x"02",x"10",x"00", -- 0x0710
    x"40",x"CC",x"80",x"60",x"10",x"08",x"03",x"00", -- 0x0718
    x"08",x"04",x"04",x"02",x"81",x"43",x"22",x"15", -- 0x0720
    x"01",x"06",x"08",x"10",x"30",x"20",x"C0",x"A0", -- 0x0728
    x"0F",x"09",x"06",x"33",x"40",x"81",x"01",x"02", -- 0x0730
    x"50",x"DE",x"61",x"D0",x"10",x"18",x"08",x"04", -- 0x0738
    x"04",x"02",x"02",x"01",x"06",x"8F",x"76",x"1A", -- 0x0740
    x"04",x"08",x"10",x"C0",x"B0",x"E8",x"2F",x"98", -- 0x0748
    x"1B",x"1C",x"0A",x"07",x"07",x"08",x"08",x"10", -- 0x0750
    x"EC",x"CC",x"B8",x"F0",x"90",x"08",x"86",x"41", -- 0x0758
    x"80",x"40",x"25",x"1F",x"17",x"0D",x"5B",x"B2", -- 0x0760
    x"21",x"41",x"42",x"B4",x"FC",x"B0",x"D8",x"EE", -- 0x0768
    x"1A",x"0F",x"05",x"1E",x"1D",x"23",x"40",x"80", -- 0x0770
    x"E9",x"56",x"F8",x"DC",x"E8",x"4C",x"82",x"81", -- 0x0778
    x"00",x"03",x"0F",x"3F",x"3F",x"7F",x"FF",x"FF", -- 0x0780
    x"00",x"80",x"80",x"E0",x"E0",x"F0",x"F8",x"FE", -- 0x0788
    x"FF",x"FF",x"7F",x"7F",x"1F",x"0F",x"0F",x"06", -- 0x0790
    x"FF",x"FF",x"FE",x"FC",x"F0",x"E0",x"00",x"00", -- 0x0798
    x"28",x"44",x"00",x"08",x"08",x"10",x"00",x"40", -- 0x07A0
    x"00",x"20",x"00",x"66",x"02",x"00",x"20",x"44", -- 0x07A8
    x"0A",x"08",x"20",x"A0",x"41",x"08",x"0A",x"00", -- 0x07B0
    x"46",x"00",x"00",x"C0",x"00",x"04",x"10",x"10", -- 0x07B8
    x"20",x"0E",x"CD",x"FC",x"1F",x"E5",x"CD",x"58", -- 0x07C0
    x"3E",x"CD",x"62",x"3D",x"CD",x"F4",x"3C",x"E1", -- 0x07C8
    x"C5",x"D5",x"4F",x"CD",x"39",x"23",x"47",x"C5", -- 0x07D0
    x"E5",x"2A",x"71",x"0E",x"E3",x"06",x"82",x"C5", -- 0x07D8
    x"33",x"CD",x"2D",x"33",x"C4",x"03",x"19",x"22", -- 0x07E0
    x"79",x"0E",x"ED",x"73",x"7B",x"0E",x"7E",x"FE", -- 0x07E8
    x"3A",x"28",x"29",x"B7",x"C2",x"99",x"10",x"23", -- 0x07F0
    x"7E",x"23",x"B6",x"CA",x"37",x"10",x"23",x"5E"  -- 0x07F8
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
       DATA <= ROM(to_integer(unsigned(ADDR)));
  end process;
end RTL;
