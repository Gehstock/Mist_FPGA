library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity twotiger_bg_bits_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of twotiger_bg_bits_1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"AA",X"AF",X"FF",X"AF",X"FF",X"AF",X"FF",X"AF",X"EB",X"FF",X"CB",X"FF",
		X"AF",X"FF",X"AF",X"FF",X"AF",X"FF",X"AF",X"FF",X"AF",X"FF",X"AF",X"FF",X"AF",X"FF",X"AF",X"FF",
		X"FE",X"AF",X"FB",X"EB",X"EF",X"EA",X"FF",X"EA",X"EF",X"1A",X"EF",X"EA",X"CF",X"FA",X"FF",X"FA",
		X"FE",X"BF",X"FE",X"BF",X"FE",X"BF",X"FE",X"BF",X"FE",X"BF",X"FE",X"BF",X"FE",X"BF",X"FE",X"BF",
		X"FF",X"F7",X"FF",X"FB",X"F3",X"37",X"FC",X"FB",X"FC",X"F7",X"A0",X"FB",X"E3",X"F7",X"E9",X"9B",
		X"EB",X"FF",X"EB",X"FF",X"EB",X"FF",X"EB",X"FF",X"EB",X"FF",X"EB",X"FF",X"EB",X"FF",X"EB",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"AF",X"FF",X"AF",X"FF",X"AF",X"FF",X"AF",X"FF",X"AF",X"FF",X"AF",X"FF",
		X"AF",X"FF",X"AF",X"EB",X"AC",X"BF",X"82",X"FF",X"8A",X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",X"FF",
		X"FA",X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",X"BF",X"FE",X"BF",X"EF",X"AF",X"EB",X"EB",X"FF",X"FF",
		X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"FE",X"BF",X"FA",X"FF",X"AB",X"FF",X"EB",X"FF",
		X"FF",X"FA",X"FF",X"F0",X"FF",X"AF",X"EF",X"AF",X"EF",X"AF",X"FF",X"AA",X"FF",X"FA",X"FF",X"FA",
		X"AA",X"AF",X"FF",X"AF",X"FF",X"AF",X"FF",X"AF",X"FF",X"FF",X"FF",X"EF",X"FE",X"FF",X"EF",X"FF",
		X"FF",X"AF",X"FF",X"AF",X"FF",X"AF",X"FF",X"AF",X"0F",X"FF",X"AF",X"FF",X"AF",X"FF",X"AF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"AA",X"AB",X"FF",X"AB",X"FF",X"AB",X"FF",X"AB",X"FF",X"AB",X"FF",X"AB",
		X"FA",X"FF",X"FA",X"FF",X"03",X"FF",X"FE",X"AA",X"FF",X"FA",X"D7",X"FA",X"DB",X"7A",X"FF",X"FA",
		X"FF",X"AB",X"FF",X"AB",X"FF",X"AB",X"FF",X"AB",X"FF",X"AB",X"FF",X"AB",X"FF",X"AB",X"FF",X"AB",
		X"FA",X"BF",X"FA",X"BF",X"FF",X"AF",X"FF",X"AF",X"FF",X"EB",X"F3",X"EB",X"F3",X"FA",X"FF",X"FA",
		X"F0",X"FF",X"EC",X"0B",X"FC",X"0F",X"BF",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"EA",X"FF",X"EA",X"DA",X"BF",X"FF",X"FF",X"D0",X"3F",X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FE",
		X"FF",X"FE",X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",
		X"FF",X"D5",X"FF",X"D5",X"FF",X"D5",X"FF",X"D5",X"FF",X"D5",X"FF",X"D5",X"FF",X"D5",X"FF",X"D5",
		X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",X"FF",X"CA",X"FF",X"C2",X"FF",X"C2",X"FF",X"F2",X"FF",X"F2",
		X"FF",X"FA",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FA",
		X"FF",X"FA",X"FF",X"F8",X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",X"FF",X"CA",X"FF",X"CA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AB",X"FF",X"AF",X"FF",X"BF",X"FF",X"BF",X"FF",
		X"AA",X"AA",X"AA",X"AB",X"AA",X"AB",X"AA",X"AF",X"AA",X"AF",X"AA",X"BF",X"AA",X"BF",X"AA",X"BF",
		X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AB",X"FF",X"AB",X"FF",X"AB",X"FF",X"AB",X"FF",
		X"AF",X"FF",X"8F",X"FF",X"AF",X"FF",X"AF",X"FF",X"AF",X"FF",X"AF",X"FF",X"AF",X"FF",X"AF",X"FF",
		X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"FF",X"AB",X"FF",
		X"05",X"40",X"10",X"10",X"50",X"54",X"51",X"14",X"51",X"14",X"54",X"14",X"10",X"10",X"05",X"40",
		X"01",X"00",X"05",X"00",X"15",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"55",X"50",
		X"15",X"50",X"50",X"14",X"50",X"14",X"00",X"50",X"15",X"40",X"50",X"00",X"50",X"14",X"55",X"54",
		X"55",X"54",X"50",X"14",X"00",X"50",X"01",X"54",X"00",X"14",X"50",X"14",X"10",X"10",X"05",X"40",
		X"05",X"50",X"04",X"50",X"10",X"50",X"10",X"50",X"40",X"50",X"55",X"54",X"00",X"50",X"00",X"50",
		X"55",X"54",X"50",X"00",X"50",X"00",X"55",X"50",X"00",X"54",X"00",X"54",X"50",X"50",X"05",X"40",
		X"15",X"50",X"50",X"14",X"50",X"00",X"55",X"54",X"50",X"14",X"50",X"14",X"50",X"14",X"15",X"50",
		X"55",X"54",X"50",X"14",X"00",X"50",X"00",X"40",X"01",X"00",X"05",X"00",X"05",X"00",X"05",X"00",
		X"15",X"50",X"50",X"14",X"50",X"14",X"15",X"50",X"50",X"14",X"50",X"14",X"50",X"14",X"15",X"50",
		X"15",X"50",X"50",X"14",X"50",X"14",X"50",X"14",X"15",X"54",X"00",X"14",X"50",X"14",X"15",X"50",
		X"AF",X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"88",X"88",X"A8",X"02",X"A0",X"20",X"8A",X"03",X"A8",X"AF",X"A2",X"3F",X"A8",X"FF",X"AB",X"FF",
		X"5F",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"A8",X"AA",X"22",X"AA",X"A8",X"AA",X"23",X"AA",X"8F",X"AA",X"0F",X"AA",X"3F",X"AA",X"BF",
		X"AA",X"FF",X"AB",X"FF",X"AB",X"FF",X"AF",X"FF",X"BF",X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AB",X"AA",X"AB",X"5A",X"AF",X"AA",X"AF",X"5A",X"AF",X"66",X"BF",X"5A",X"BF",X"55",X"BF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"05",X"40",X"05",X"40",X"14",X"50",X"10",X"10",X"50",X"14",X"55",X"54",X"50",X"14",X"50",X"14",
		X"55",X"50",X"50",X"14",X"50",X"14",X"55",X"50",X"50",X"14",X"50",X"14",X"50",X"14",X"55",X"50",
		X"15",X"50",X"50",X"14",X"50",X"14",X"50",X"00",X"50",X"00",X"50",X"14",X"50",X"14",X"15",X"50",
		X"55",X"40",X"50",X"50",X"50",X"14",X"50",X"14",X"50",X"14",X"50",X"14",X"50",X"50",X"55",X"40",
		X"55",X"54",X"50",X"14",X"50",X"00",X"55",X"00",X"50",X"00",X"50",X"14",X"50",X"14",X"55",X"54",
		X"55",X"54",X"50",X"14",X"50",X"00",X"55",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",
		X"15",X"50",X"50",X"14",X"50",X"00",X"50",X"00",X"50",X"54",X"50",X"14",X"50",X"14",X"15",X"50",
		X"50",X"14",X"50",X"14",X"50",X"14",X"55",X"54",X"50",X"14",X"50",X"14",X"50",X"14",X"50",X"14",
		X"55",X"50",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"55",X"50",
		X"55",X"50",X"01",X"40",X"01",X"40",X"01",X"40",X"51",X"40",X"51",X"40",X"15",X"00",X"04",X"00",
		X"50",X"14",X"50",X"40",X"51",X"00",X"55",X"00",X"51",X"40",X"51",X"50",X"50",X"54",X"50",X"54",
		X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"14",X"55",X"54",
		X"50",X"14",X"50",X"14",X"54",X"54",X"54",X"54",X"55",X"54",X"51",X"14",X"51",X"14",X"50",X"14",
		X"40",X"14",X"50",X"14",X"54",X"14",X"54",X"14",X"51",X"14",X"50",X"54",X"50",X"54",X"50",X"14",
		X"15",X"50",X"50",X"14",X"50",X"14",X"50",X"14",X"50",X"14",X"50",X"14",X"50",X"14",X"15",X"50",
		X"55",X"50",X"50",X"14",X"50",X"14",X"50",X"14",X"55",X"50",X"50",X"00",X"50",X"00",X"50",X"00",
		X"15",X"50",X"50",X"14",X"50",X"14",X"50",X"14",X"50",X"14",X"50",X"54",X"50",X"10",X"15",X"44",
		X"55",X"50",X"50",X"14",X"50",X"14",X"50",X"50",X"55",X"00",X"51",X"40",X"50",X"50",X"50",X"14",
		X"15",X"50",X"50",X"14",X"50",X"00",X"15",X"00",X"00",X"50",X"00",X"14",X"50",X"14",X"15",X"50",
		X"55",X"50",X"45",X"10",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",
		X"50",X"14",X"50",X"14",X"50",X"14",X"50",X"14",X"50",X"14",X"50",X"14",X"50",X"14",X"15",X"50",
		X"50",X"14",X"50",X"14",X"50",X"14",X"10",X"10",X"14",X"50",X"04",X"50",X"04",X"40",X"05",X"40",
		X"51",X"14",X"51",X"14",X"51",X"14",X"51",X"14",X"51",X"14",X"15",X"50",X"14",X"50",X"04",X"10",
		X"40",X"04",X"50",X"14",X"14",X"50",X"05",X"40",X"01",X"40",X"15",X"50",X"54",X"14",X"50",X"14",
		X"40",X"04",X"50",X"14",X"14",X"50",X"15",X"40",X"05",X"40",X"05",X"00",X"05",X"00",X"05",X"00",
		X"55",X"54",X"50",X"14",X"00",X"50",X"01",X"40",X"05",X"00",X"14",X"00",X"50",X"14",X"55",X"54",
		X"5F",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"A8",X"AA",X"22",X"AA",X"A8",X"AA",X"23",X"AA",X"8F",X"AA",X"0F",X"AA",X"3F",X"AA",X"BF",
		X"AA",X"FF",X"AB",X"FF",X"AB",X"FF",X"AF",X"FF",X"BF",X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AB",X"AA",X"AB",X"5A",X"AF",X"AA",X"AF",X"5A",X"AF",X"66",X"BF",X"5A",X"BF",X"55",X"BF",
		X"FF",X"FF",X"00",X"00",X"A2",X"A8",X"65",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"AA",X"A2",X"99",X"6A",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F2",X"A0",X"2A",X"AA",X"A5",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"8A",X"AA",X"A9",X"59",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"AA",X"0A",X"51",X"A9",X"55",
		X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"FC",X"FF",X"03",X"00",X"03",X"00",X"03",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"AA",X"FE",X"29",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"A9",X"6A",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"A5",X"65",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E9",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",
		X"0F",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"F0",X"FF",X"F0",X"FF",X"F0",X"FF",X"F0",X"FF",X"FF",X"C3",X"FF",X"C3",
		X"FF",X"F0",X"FF",X"F0",X"FF",X"F0",X"FF",X"F0",X"FF",X"F0",X"FF",X"F0",X"FF",X"F0",X"FF",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",X"FF",
		X"FC",X"3F",X"FC",X"3F",X"FC",X"3F",X"FC",X"3F",X"FC",X"3F",X"FC",X"3B",X"FC",X"3F",X"FC",X"3F",
		X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"FF",X"7F",X"FF",X"B0",X"FF",X"80",X"FF",X"C0",
		X"FF",X"C0",X"FF",X"C0",X"FF",X"C0",X"FF",X"C0",X"FF",X"C0",X"FF",X"C0",X"FF",X"C0",X"FF",X"C0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"E0",X"FF",X"F0",X"FE",X"F0",X"FF",X"F0",X"EF",X"F0",X"FF",X"E0",
		X"FF",X"E0",X"FF",X"F0",X"FF",X"F0",X"FF",X"F0",X"FF",X"F2",X"FE",X"0F",X"FF",X"0F",X"FF",X"0F",
		X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",X"FC",X"FF",X"FF",X"FF",X"FB",X"FF",X"EF",X"DF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"FF",X"C0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",
		X"0F",X"FF",X"0F",X"BF",X"F0",X"FF",X"F8",X"FF",X"F8",X"FF",X"00",X"FF",X"00",X"FF",X"0F",X"FF",
		X"F0",X"FF",X"F0",X"FF",X"F0",X"FF",X"F8",X"00",X"FB",X"FF",X"FF",X"EF",X"FF",X"FE",X"FF",X"FF",
		X"F0",X"FF",X"F0",X"FF",X"F0",X"FF",X"F0",X"00",X"FF",X"F0",X"FF",X"F1",X"FF",X"F1",X"FF",X"F0",
		X"AB",X"CA",X"EB",X"F3",X"EB",X"C3",X"EB",X"83",X"EB",X"C3",X"EA",X"C3",X"AB",X"C3",X"EB",X"C3",
		X"FF",X"FF",X"FF",X"FF",X"CA",X"AA",X"C0",X"FF",X"C0",X"FF",X"C0",X"FF",X"C0",X"FF",X"C0",X"FF",
		X"FF",X"0F",X"FF",X"07",X"FF",X"C4",X"0F",X"FF",X"0F",X"FF",X"0F",X"FF",X"0E",X"FF",X"0F",X"FF",
		X"C0",X"FF",X"C0",X"FF",X"C0",X"FF",X"C0",X"FF",X"C0",X"FF",X"C0",X"FF",X"C0",X"FF",X"C0",X"FF",
		X"FC",X"0F",X"FC",X"0F",X"F0",X"FF",X"F0",X"FF",X"C3",X"FF",X"C3",X"FF",X"0F",X"F7",X"0F",X"C7",
		X"FF",X"0F",X"F0",X"3F",X"F0",X"3F",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"FF",X"FF",X"FF",
		X"FA",X"AB",X"C3",X"FB",X"C3",X"FB",X"0F",X"FB",X"0F",X"3F",X"0F",X"BB",X"0F",X"AF",X"0F",X"BF",
		X"03",X"FF",X"AB",X"FF",X"FE",X"AF",X"FC",X"0F",X"FC",X"0F",X"03",X"FF",X"03",X"FB",X"03",X"FF",
		X"55",X"55",X"55",X"15",X"55",X"55",X"11",X"14",X"55",X"55",X"55",X"15",X"55",X"55",X"55",X"15",
		X"44",X"44",X"55",X"55",X"55",X"15",X"11",X"54",X"55",X"55",X"55",X"15",X"55",X"55",X"55",X"55",
		X"55",X"58",X"55",X"54",X"55",X"60",X"55",X"51",X"55",X"81",X"55",X"45",X"56",X"05",X"55",X"15",
		X"58",X"15",X"54",X"55",X"60",X"55",X"51",X"55",X"81",X"55",X"45",X"55",X"05",X"55",X"15",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"55",
		X"7F",X"F5",X"AA",X"A5",X"EF",X"C1",X"9F",X"FD",X"E7",X"F9",X"FB",X"EF",X"FE",X"BC",X"6B",X"E9",
		X"FF",X"FD",X"AA",X"AA",X"6F",X"C3",X"CF",X"B0",X"FE",X"FC",X"FB",X"FF",X"AF",X"FD",X"AA",X"A5",
		X"FF",X"FE",X"AA",X"AA",X"43",X"F9",X"FE",X"F3",X"FE",X"BF",X"FB",X"EC",X"6F",X"FA",X"9A",X"AB",
		X"5F",X"FD",X"FA",X"A9",X"C3",X"FB",X"BF",X"F6",X"2F",X"DB",X"FB",X"EF",X"FE",X"BF",X"6B",X"E9",
		X"3F",X"FD",X"AA",X"A5",X"EF",X"C1",X"5F",X"FC",X"45",X"FB",X"39",X"EF",X"FE",X"BF",X"6B",X"E9",
		X"59",X"66",X"56",X"5A",X"59",X"66",X"55",X"AA",X"56",X"66",X"56",X"AA",X"55",X"6A",X"5A",X"AA",
		X"AA",X"AA",X"9A",X"A5",X"AA",X"95",X"AA",X"99",X"9A",X"95",X"55",X"65",X"99",X"95",X"AA",X"55",
		X"55",X"56",X"55",X"55",X"56",X"95",X"5A",X"A5",X"5A",X"A5",X"56",X"95",X"55",X"56",X"9A",X"6A",
		X"55",X"AA",X"55",X"AA",X"59",X"82",X"65",X"8A",X"45",X"09",X"4A",X"26",X"50",X"28",X"54",X"01",
		X"2A",X"8A",X"AA",X"AA",X"28",X"8A",X"AA",X"AA",X"2A",X"AA",X"0A",X"8A",X"0A",X"AA",X"00",X"8A",
		X"2A",X"AA",X"AA",X"AA",X"2A",X"AA",X"AA",X"A8",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"08",X"8A",
		X"55",X"55",X"55",X"55",X"95",X"66",X"9A",X"59",X"99",X"95",X"AA",X"A6",X"A9",X"99",X"AA",X"AA",
		X"FF",X"FF",X"FC",X"CF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FB",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"57",X"FB",X"7B",X"E5",X"FE",X"FF",X"55",X"55",
		X"FF",X"FF",X"F5",X"55",X"FF",X"FF",X"55",X"5D",X"5F",X"FB",X"7B",X"F5",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"55",X"55",X"FF",X"FF",X"FB",X"FF",X"57",X"BF",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"F5",X"55",X"FF",X"FF",X"FF",X"FF",X"57",X"BF",X"7B",X"F5",X"55",X"55",X"55",X"55",
		X"BF",X"FF",X"55",X"55",X"FF",X"57",X"FB",X"FF",X"56",X"5B",X"55",X"55",X"FF",X"F5",X"55",X"55",
		X"FF",X"FF",X"EF",X"FF",X"BE",X"57",X"FF",X"AF",X"F7",X"5F",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"EF",X"FB",X"57",X"DA",X"F5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"D5",X"EB",X"5A",X"B7",X"55",X"55",X"FF",X"F5",X"55",X"55",X"57",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"BB",X"FF",X"5F",X"F7",X"7F",X"AD",X"FA",X"F5",X"55",X"55",X"55",X"55",
		X"FF",X"FD",X"7F",X"55",X"FF",X"FF",X"5F",X"F7",X"5F",X"FD",X"57",X"F5",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"77",X"57",X"FF",X"7F",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"F5",X"55",X"FD",X"D5",X"FF",X"FD",X"FF",X"FA",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5D",X"57",X"7F",X"5F",X"FF",X"5F",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"D5",X"55",X"FF",X"55",X"FD",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"F5",X"57",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"D5",X"55",X"F7",X"55",X"FF",X"FD",X"FF",X"F5",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"DD",X"5D",X"FF",X"7F",X"FF",X"7F",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"D5",X"55",X"FF",X"D5",X"FF",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"75",X"55",X"FD",X"7F",X"FF",X"7F",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"D5",X"55",X"FF",X"D5",X"FF",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5D",X"55",X"5F",X"57",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"5D",X"55",X"7D",X"55",X"FF",X"55",X"FF",X"FF",X"FF",X"FD",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"D7",X"FD",X"77",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"5D",X"55",X"DD",X"55",X"FF",X"D5",X"FF",X"FF",X"FF",X"FD",
		X"55",X"55",X"55",X"55",X"55",X"55",X"5D",X"55",X"5F",X"7D",X"5D",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"D5",X"55",X"55",X"55",X"FF",X"D5",X"FF",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"55",X"55",X"FF",X"FF",X"5F",X"FF",X"5F",X"FF",
		X"75",X"5D",X"5D",X"75",X"57",X"D5",X"F5",X"55",X"FD",X"75",X"F5",X"5F",X"D7",X"D7",X"5F",X"F5",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"FF",X"FD",X"FF",X"F5",X"FF",X"D5",
		X"55",X"55",X"55",X"55",X"55",X"57",X"55",X"5F",X"FF",X"FF",X"5F",X"FF",X"7F",X"FF",X"7F",X"FF",
		X"75",X"55",X"7D",X"55",X"7D",X"55",X"FF",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"FF",X"FF",X"FF",X"D5",X"FF",X"55",X"FD",X"55",
		X"00",X"00",X"28",X"08",X"6A",X"2A",X"1A",X"AA",X"A6",X"AA",X"A9",X"A8",X"AA",X"60",X"AA",X"9A",
		X"20",X"00",X"98",X"08",X"9A",X"26",X"99",X"96",X"95",X"56",X"55",X"58",X"55",X"60",X"AA",X"AA",
		X"59",X"66",X"56",X"5A",X"59",X"66",X"55",X"AA",X"56",X"66",X"56",X"AA",X"55",X"6A",X"5A",X"AA",
		X"00",X"00",X"00",X"00",X"0A",X"A8",X"28",X"28",X"28",X"28",X"28",X"28",X"2A",X"A0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"80",X"0A",X"80",X"02",X"80",X"02",X"80",X"0A",X"A0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0A",X"A0",X"20",X"28",X"02",X"A0",X"28",X"00",X"2A",X"A8",X"00",X"00",
		X"00",X"00",X"00",X"00",X"2A",X"A8",X"00",X"20",X"00",X"80",X"20",X"28",X"0A",X"A8",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"A0",X"02",X"20",X"08",X"20",X"2A",X"A8",X"00",X"A0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"2A",X"A8",X"20",X"00",X"2A",X"A8",X"00",X"28",X"2A",X"A0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"2A",X"A8",X"28",X"00",X"2A",X"A0",X"28",X"28",X"2A",X"A8",X"00",X"00",
		X"00",X"00",X"00",X"00",X"2A",X"A8",X"00",X"20",X"00",X"80",X"02",X"80",X"02",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"2A",X"A8",X"28",X"28",X"0A",X"A0",X"28",X"28",X"2A",X"A8",X"00",X"00",
		X"00",X"00",X"00",X"00",X"2A",X"A8",X"28",X"28",X"0A",X"A8",X"00",X"28",X"2A",X"A8",X"00",X"00",
		X"55",X"55",X"A5",X"55",X"55",X"59",X"55",X"55",X"69",X"65",X"55",X"55",X"55",X"55",X"55",X"65",
		X"95",X"65",X"55",X"55",X"59",X"59",X"56",X"56",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"59",X"55",X"56",X"65",X"96",X"65",X"56",X"59",X"55",X"59",X"65",X"55",X"65",X"55",X"55",
		X"59",X"55",X"55",X"65",X"56",X"55",X"56",X"59",X"55",X"59",X"95",X"59",X"55",X"59",X"55",X"55",
		X"55",X"59",X"65",X"59",X"65",X"59",X"66",X"65",X"95",X"65",X"95",X"65",X"55",X"55",X"55",X"55",
		X"55",X"95",X"65",X"55",X"65",X"95",X"65",X"95",X"95",X"56",X"96",X"56",X"56",X"59",X"55",X"55",
		X"56",X"56",X"55",X"59",X"95",X"65",X"55",X"55",X"56",X"55",X"59",X"59",X"65",X"A5",X"56",X"55",
		X"55",X"56",X"5A",X"95",X"A5",X"55",X"55",X"55",X"59",X"A9",X"55",X"55",X"55",X"55",X"69",X"55",
		X"56",X"95",X"59",X"55",X"55",X"65",X"55",X"95",X"56",X"55",X"55",X"55",X"65",X"55",X"95",X"59",
		X"55",X"55",X"55",X"65",X"59",X"65",X"59",X"55",X"55",X"56",X"65",X"56",X"65",X"96",X"55",X"59",
		X"65",X"55",X"95",X"59",X"95",X"59",X"55",X"59",X"56",X"59",X"56",X"55",X"55",X"65",X"59",X"55",
		X"59",X"55",X"95",X"55",X"96",X"65",X"66",X"65",X"65",X"65",X"65",X"55",X"65",X"59",X"55",X"55",
		X"55",X"55",X"56",X"59",X"96",X"56",X"95",X"56",X"65",X"95",X"65",X"95",X"65",X"55",X"55",X"65",
		X"56",X"95",X"65",X"65",X"59",X"55",X"56",X"55",X"55",X"95",X"95",X"55",X"65",X"59",X"65",X"56",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"AA",X"A6",X"BA",X"AA",X"A9",X"E7",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"9A",X"69",X"A6",X"56",X"99",X"6A",
		X"01",X"00",X"15",X"50",X"10",X"00",X"15",X"40",X"10",X"00",X"15",X"50",X"01",X"00",X"01",X"00",
		X"FF",X"FF",X"FE",X"AA",X"FF",X"AA",X"FF",X"EA",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"AA",X"FA",X"AA",
		X"FD",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"D5",X"FF",X"F5",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"EA",X"FF",X"FA",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FE",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"AA",X"EA",X"AA",X"FA",X"AA",X"FA",X"AA",
		X"FE",X"AA",X"FE",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"EA",X"FF",X"EA",X"FF",X"FA",X"FF",X"FA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"BF",X"FF",
		X"BF",X"FF",X"AF",X"FF",X"AF",X"FF",X"AF",X"FF",X"AF",X"FF",X"AF",X"FF",X"AF",X"FF",X"AF",X"FF",
		X"AB",X"FF",X"AB",X"FF",X"AB",X"FF",X"AB",X"FF",X"AB",X"FF",X"AB",X"FF",X"AB",X"FF",X"AB",X"FF",
		X"AB",X"FF",X"AB",X"FF",X"AB",X"FF",X"A3",X"FF",X"83",X"FF",X"83",X"FF",X"8F",X"FF",X"8F",X"FF",
		X"AF",X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",X"AF",X"FF",
		X"AF",X"FF",X"2F",X"FF",X"AB",X"FF",X"AB",X"FF",X"AB",X"FF",X"AB",X"FF",X"A3",X"FF",X"A3",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A2",X"A8",X"59",X"A6",X"8A",X"99",X"99",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"6A",X"AA",X"88",X"A9",X"66",X"46",X"19",X"99",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"64",X"8A",X"9A",X"9A",
		X"AA",X"55",X"AA",X"55",X"82",X"65",X"A2",X"59",X"60",X"51",X"98",X"A1",X"28",X"05",X"40",X"15",
		X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"59",X"AA",X"9A",X"AA",X"A6",X"AA",X"A9",X"AA",X"99",
		X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"95",X"55",X"65",X"55",X"99",X"55",X"95",X"55",X"65",X"95",
		X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"AA",X"BF",X"AA",X"FF",X"AB",X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AB",X"AA",X"AF",
		X"55",X"7F",X"55",X"FF",X"55",X"FF",X"57",X"FF",X"5F",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"BF",X"AA",X"FF",X"AA",X"FF",X"AB",X"FF",X"AF",X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"BF",X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AB",X"AA",X"AB",X"AA",X"AF",X"AA",X"AF",
		X"AA",X"BF",X"AA",X"BF",X"AA",X"FF",X"AA",X"FF",X"AB",X"FF",X"AB",X"FF",X"AF",X"FF",X"AF",X"FF",
		X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"65",X"AA",X"A6",X"AA",X"9A",X"AA",X"6A",X"AA",X"66",X"AA",
		X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"55",X"A6",X"55",X"99",X"99",X"66",X"66",X"56",X"66",X"9A",
		X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"55",X"56",X"55",X"59",X"55",X"66",X"55",X"56",X"56",X"59",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"8A",X"AA",X"65",X"2A",X"A2",X"9A",X"66",X"66",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A9",X"6A",X"22",X"91",X"99",X"66",X"64",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A2",X"19",X"A6",X"A6",
		X"5A",X"6A",X"69",X"AA",X"5A",X"66",X"A6",X"AA",X"99",X"AA",X"AA",X"AA",X"A2",X"19",X"66",X"66",
		X"A9",X"A6",X"AA",X"69",X"AA",X"A5",X"AA",X"AA",X"AA",X"A6",X"AA",X"AA",X"A8",X"8A",X"99",X"98",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"59",X"9A",X"A5",
		X"A9",X"65",X"A6",X"59",X"A9",X"96",X"9A",X"69",X"A6",X"A5",X"AA",X"65",X"A9",X"AA",X"AA",X"99",
		X"65",X"55",X"95",X"55",X"69",X"55",X"99",X"59",X"66",X"95",X"9A",X"65",X"69",X"9A",X"9A",X"95",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"DF",X"47",X"FF",X"C7",X"FF",X"CF",
		X"3F",X"FF",X"8F",X"EB",X"E3",X"FB",X"F8",X"FF",X"FE",X"3F",X"FF",X"CF",X"F9",X"9A",X"FF",X"57",
		X"FF",X"FF",X"CF",X"FF",X"33",X"33",X"CF",X"FF",X"FF",X"FF",X"CC",X"CF",X"FF",X"FF",X"CF",X"FF",
		X"FB",X"FF",X"F9",X"9A",X"FF",X"CF",X"FF",X"2A",X"FC",X"BF",X"F2",X"EB",X"CB",X"EF",X"2F",X"FF",
		X"FF",X"FE",X"FF",X"FF",X"33",X"23",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"EF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0A",X"A8",X"0A",X"A8",X"0A",X"A8",X"2A",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",
		X"2A",X"A8",X"2A",X"A8",X"2A",X"A8",X"2A",X"A8",X"2A",X"A8",X"2A",X"A8",X"2A",X"A8",X"2A",X"A8",
		X"2A",X"A8",X"2A",X"A8",X"2A",X"A8",X"2A",X"A8",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"AA",X"02",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",
		X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",
		X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"02",X"AA",X"00",X"AA",
		X"AA",X"A0",X"AA",X"A8",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",
		X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",
		X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"0A",X"00",X"2A",X"00",X"AA",X"02",X"AA",X"0A",X"AA",
		X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"25",X"AA",X"25",X"69",X"09",X"56",X"02",X"56",
		X"00",X"95",X"00",X"25",X"00",X"25",X"00",X"09",X"00",X"02",X"00",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"08",X"00",X"20",X"00",X"80",X"02",X"00",X"08",X"02",
		X"2A",X"02",X"AA",X"82",X"AA",X"AA",X"AA",X"96",X"AA",X"96",X"A8",X"92",X"A0",X"A0",X"A0",X"20",
		X"80",X"A8",X"80",X"80",X"80",X"22",X"80",X"2B",X"80",X"0B",X"A0",X"0B",X"AA",X"2E",X"AA",X"BF",
		X"AA",X"AA",X"AA",X"A5",X"6A",X"A9",X"5A",X"A9",X"5A",X"A9",X"56",X"A9",X"96",X"A5",X"25",X"A5",
		X"25",X"A5",X"09",X"6A",X"09",X"6A",X"02",X"5A",X"00",X"9A",X"00",X"9A",X"00",X"9A",X"00",X"2A",
		X"00",X"2A",X"00",X"2A",X"00",X"2A",X"00",X"2A",X"00",X"2A",X"00",X"2A",X"00",X"AA",X"00",X"AA",
		X"00",X"AA",X"02",X"AA",X"09",X"A9",X"25",X"65",X"25",X"65",X"95",X"5A",X"95",X"56",X"95",X"55",
		X"25",X"55",X"25",X"55",X"09",X"55",X"09",X"55",X"25",X"55",X"95",X"55",X"95",X"55",X"95",X"55",
		X"95",X"55",X"25",X"55",X"25",X"55",X"25",X"55",X"09",X"55",X"09",X"55",X"02",X"55",X"02",X"55",
		X"02",X"55",X"02",X"55",X"00",X"AA",X"02",X"6A",X"02",X"D5",X"02",X"D5",X"0B",X"95",X"0A",X"55",
		X"09",X"55",X"0A",X"55",X"02",X"55",X"02",X"56",X"02",X"56",X"02",X"96",X"00",X"96",X"00",X"96",
		X"00",X"96",X"02",X"56",X"02",X"55",X"02",X"5D",X"00",X"B5",X"02",X"D5",X"02",X"55",X"00",X"AA",
		X"2A",X"80",X"88",X"20",X"20",X"80",X"82",X"80",X"0A",X"A2",X"0A",X"AA",X"02",X"A6",X"02",X"A5",
		X"02",X"8A",X"2A",X"8B",X"BF",X"8B",X"EA",X"0A",X"80",X"20",X"2A",X"3A",X"2B",X"02",X"00",X"02",
		X"00",X"00",X"00",X"A8",X"82",X"FE",X"8B",X"FE",X"EF",X"FE",X"FF",X"FB",X"FF",X"A0",X"BE",X"0A",
		X"E8",X"3C",X"B8",X"00",X"6E",X"00",X"6F",X"AA",X"5B",X"FF",X"56",X"FF",X"55",X"AA",X"5A",X"95",
		X"AA",X"A5",X"AA",X"A5",X"AA",X"A5",X"AA",X"A9",X"AA",X"A9",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"BE",X"AA",X"BE",X"AA",X"BE",X"AA",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A9",X"55",
		X"99",X"95",X"59",X"56",X"65",X"55",X"95",X"55",X"99",X"56",X"55",X"66",X"55",X"58",X"AA",X"A8",
		X"55",X"58",X"55",X"58",X"55",X"58",X"55",X"58",X"A9",X"58",X"65",X"56",X"65",X"56",X"65",X"56",
		X"65",X"56",X"65",X"55",X"65",X"55",X"65",X"55",X"95",X"55",X"A5",X"55",X"89",X"55",X"82",X"55",
		X"82",X"55",X"80",X"95",X"80",X"95",X"80",X"AA",X"82",X"55",X"82",X"D5",X"8B",X"55",X"89",X"75",
		X"89",X"76",X"82",X"56",X"82",X"56",X"02",X"56",X"02",X"58",X"02",X"58",X"02",X"58",X"02",X"58",
		X"02",X"58",X"02",X"5E",X"82",X"5F",X"89",X"59",X"69",X"A9",X"5A",X"A9",X"5A",X"A9",X"A0",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"00",
		X"60",X"00",X"A0",X"00",X"F8",X"00",X"BE",X"00",X"2E",X"00",X"88",X"00",X"C8",X"00",X"08",X"00",
		X"82",X"00",X"82",X"00",X"82",X"00",X"E8",X"00",X"FA",X"00",X"FE",X"00",X"BE",X"00",X"2E",X"00",
		X"A8",X"00",X"80",X"00",X"A0",X"00",X"BA",X"80",X"BA",X"A0",X"BE",X"A8",X"FE",X"AA",X"BE",X"AA",
		X"BF",X"AA",X"BF",X"A8",X"BF",X"A8",X"BF",X"AA",X"BF",X"AA",X"BF",X"AA",X"BF",X"AA",X"BF",X"AA",
		X"BF",X"AA",X"BB",X"AA",X"BB",X"A8",X"BA",X"A8",X"B9",X"A8",X"6A",X"A8",X"5A",X"A0",X"55",X"80",
		X"56",X"80",X"5A",X"80",X"6A",X"80",X"9A",X"80",X"9A",X"80",X"9A",X"00",X"9A",X"00",X"9A",X"00",
		X"A8",X"A0",X"80",X"08",X"80",X"02",X"82",X"82",X"8B",X"C2",X"82",X"E2",X"22",X"88",X"22",X"E0",
		X"22",X"80",X"88",X"80",X"88",X"80",X"68",X"80",X"68",X"80",X"58",X"80",X"58",X"80",X"58",X"80",
		X"58",X"80",X"58",X"80",X"68",X"80",X"88",X"80",X"88",X"80",X"88",X"80",X"88",X"80",X"88",X"80",
		X"08",X"80",X"08",X"80",X"08",X"80",X"08",X"80",X"08",X"80",X"08",X"80",X"08",X"80",X"08",X"80",
		X"08",X"80",X"08",X"80",X"88",X"80",X"68",X"80",X"7A",X"80",X"57",X"60",X"95",X"60",X"AA",X"80",
		X"00",X"02",X"00",X"02",X"00",X"08",X"00",X"20",X"00",X"22",X"00",X"20",X"00",X"28",X"00",X"82",
		X"00",X"88",X"02",X"02",X"02",X"20",X"00",X"A0",X"00",X"0A",X"00",X"02",X"02",X"AA",X"0B",X"EF",
		X"0B",X"BE",X"0B",X"BB",X"02",X"BB",X"0B",X"BB",X"2F",X"BB",X"2E",X"FB",X"2E",X"FB",X"2E",X"FB",
		X"2E",X"FB",X"2E",X"FB",X"2E",X"FB",X"26",X"F9",X"0A",X"F9",X"0A",X"F9",X"02",X"F9",X"02",X"F9",
		X"02",X"FB",X"02",X"FA",X"02",X"F8",X"02",X"B8",X"00",X"B8",X"00",X"A0",X"00",X"00",X"00",X"02",
		X"00",X"B0",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"09",X"00",X"AD",X"00",X"95",X"00",X"AA",
		X"28",X"00",X"AA",X"2A",X"AA",X"AA",X"A8",X"AA",X"82",X"28",X"2A",X"02",X"82",X"00",X"00",X"80",
		X"80",X"20",X"E8",X"98",X"E0",X"EA",X"80",X"E8",X"00",X"00",X"A0",X"02",X"00",X"02",X"02",X"00",
		X"A8",X"00",X"00",X"0A",X"00",X"0B",X"2A",X"AE",X"BF",X"FB",X"FF",X"EF",X"FF",X"BF",X"AA",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FA",X"AB",X"FA",X"AB",X"FA",X"AB",X"FA",X"AB",X"EF",X"BF",X"EF",X"BF",
		X"EF",X"BF",X"FA",X"FF",X"FF",X"FF",X"7F",X"FF",X"7F",X"FF",X"5F",X"FF",X"57",X"FF",X"55",X"FF",
		X"55",X"FA",X"AA",X"A0",X"2F",X"80",X"2F",X"8A",X"AA",X"AF",X"BF",X"FF",X"BB",X"FF",X"FB",X"FF",
		X"FB",X"FF",X"FB",X"FF",X"AB",X"FF",X"8A",X"AA",X"80",X"00",X"8A",X"80",X"82",X"00",X"82",X"00",
		X"82",X"00",X"82",X"00",X"80",X"80",X"80",X"80",X"20",X"80",X"20",X"80",X"20",X"80",X"20",X"80",
		X"20",X"80",X"20",X"80",X"20",X"80",X"20",X"80",X"20",X"80",X"20",X"80",X"08",X"20",X"02",X"AA",
		X"09",X"65",X"09",X"65",X"09",X"65",X"09",X"65",X"09",X"65",X"09",X"65",X"09",X"65",X"09",X"65",
		X"02",X"65",X"02",X"65",X"02",X"65",X"02",X"59",X"02",X"59",X"02",X"59",X"02",X"59",X"02",X"6D",
		X"09",X"65",X"2D",X"65",X"B5",X"67",X"D5",X"65",X"55",X"65",X"56",X"A5",X"68",X"25",X"80",X"0A",
		X"00",X"00",X"00",X"00",X"28",X"00",X"BE",X"A0",X"2F",X"80",X"BE",X"00",X"BF",X"A0",X"2F",X"F8",
		X"0B",X"F8",X"02",X"A8",X"0B",X"FA",X"A5",X"FF",X"B9",X"7F",X"FE",X"5F",X"FF",X"97",X"BE",X"25",
		X"B8",X"0A",X"F8",X"25",X"E8",X"A7",X"BE",X"9F",X"FB",X"FF",X"EF",X"FD",X"FF",X"F5",X"FF",X"D5",
		X"FF",X"D5",X"FF",X"56",X"FD",X"58",X"F5",X"60",X"D5",X"60",X"D5",X"80",X"D6",X"00",X"D8",X"00",
		X"E0",X"00",X"E0",X"00",X"E0",X"00",X"E0",X"00",X"E0",X"00",X"E8",X"00",X"E2",X"00",X"82",X"00",
		X"0A",X"00",X"2F",X"80",X"BF",X"E0",X"FF",X"F8",X"FF",X"F8",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",
		X"FF",X"FE",X"FF",X"A8",X"EA",X"80",X"80",X"80",X"00",X"80",X"02",X"00",X"02",X"00",X"02",X"00",
		X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",
		X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"20",X"00",X"80",X"00",
		X"60",X"00",X"E0",X"00",X"78",X"00",X"78",X"00",X"58",X"00",X"58",X"00",X"58",X"00",X"58",X"00",
		X"58",X"00",X"58",X"00",X"58",X"00",X"60",X"00",X"60",X"00",X"60",X"00",X"60",X"00",X"60",X"00",
		X"60",X"00",X"60",X"00",X"A0",X"00",X"A0",X"00",X"E0",X"00",X"78",X"00",X"5E",X"00",X"AA",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"E0",X"00",X"FA",X"00",X"FF",X"80",X"FF",X"E0",
		X"FF",X"58",X"FD",X"60",X"F5",X"80",X"D5",X"80",X"56",X"00",X"58",X"00",X"60",X"00",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"2A",X"00",X"2A",
		X"00",X"2A",X"00",X"2A",X"00",X"2A",X"00",X"2A",X"00",X"2A",X"00",X"2A",X"00",X"2A",X"00",X"2A",
		X"00",X"2A",X"00",X"2A",X"00",X"2A",X"00",X"2A",X"00",X"2A",X"00",X"2A",X"00",X"2A",X"A0",X"2A",
		X"98",X"2A",X"98",X"2A",X"26",X"2A",X"09",X"AA",X"09",X"6A",X"02",X"8A",X"02",X"00",X"02",X"02",
		X"02",X"0B",X"02",X"0B",X"00",X"82",X"00",X"20",X"00",X"08",X"00",X"02",X"00",X"00",X"00",X"00",
		X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"0B",X"00",X"2D",X"00",X"B5",X"00",X"95",
		X"FE",X"75",X"FE",X"55",X"FE",X"55",X"FF",X"A5",X"FF",X"F9",X"FE",X"BA",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"11",X"00",X"11",X"01",X"01",X"01",X"11",
		X"01",X"11",X"01",X"11",X"00",X"10",X"00",X"11",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"2A",X"00",X"AA",X"02",X"6A",X"02",X"6A",X"02",X"95",
		X"2A",X"AA",X"AA",X"F8",X"AB",X"FE",X"AA",X"BF",X"A8",X"2B",X"AA",X"3A",X"AA",X"0A",X"AA",X"00",
		X"AA",X"0A",X"A8",X"2F",X"AE",X"BF",X"AF",X"FE",X"9B",X"FB",X"96",X"A2",X"A5",X"60",X"A5",X"60",
		X"5A",X"5A",X"5A",X"55",X"5A",X"95",X"62",X"AA",X"62",X"AA",X"62",X"AA",X"60",X"AA",X"A0",X"AA",
		X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"9A",X"A0",X"95",X"A2",X"55",X"A2",X"55",X"A2",X"55",
		X"A2",X"56",X"A9",X"55",X"A9",X"55",X"A5",X"55",X"A5",X"55",X"89",X"55",X"02",X"55",X"82",X"55",
		X"E2",X"55",X"E2",X"55",X"89",X"55",X"25",X"55",X"A5",X"55",X"25",X"55",X"09",X"55",X"09",X"55",
		X"02",X"55",X"09",X"AA",X"2F",X"56",X"2D",X"5A",X"B5",X"58",X"95",X"68",X"95",X"60",X"95",X"A0",
		X"D5",X"80",X"D6",X"80",X"D6",X"00",X"5A",X"00",X"58",X"00",X"58",X"00",X"68",X"00",X"60",X"00",
		X"AF",X"FF",X"DB",X"FF",X"7A",X"FF",X"5F",X"AF",X"55",X"6F",X"55",X"6F",X"AA",X"BF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"10",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"10",X"11",X"10",X"11",X"00",X"10",X"00",X"10",X"00",
		X"10",X"00",X"10",X"00",X"00",X"00",X"02",X"A0",X"AA",X"A8",X"9A",X"A8",X"A6",X"A8",X"A5",X"60",
		X"0A",X"AA",X"02",X"FF",X"AB",X"FE",X"2F",X"EA",X"2F",X"B0",X"0A",X"B2",X"02",X"A2",X"00",X"02",
		X"8A",X"82",X"8B",X"E0",X"EF",X"FA",X"AA",X"FF",X"F5",X"BF",X"AA",X"2A",X"00",X"09",X"00",X"09",
		X"00",X"A5",X"AA",X"55",X"59",X"55",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"6A",X"6A",X"AA",X"AA",
		X"AA",X"AA",X"9A",X"9A",X"AA",X"AA",X"AA",X"A6",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"55",X"65",X"55",X"65",X"55",X"65",X"55",X"65",X"55",X"65",X"55",X"65",X"56",X"65",X"56",
		X"65",X"56",X"65",X"56",X"65",X"55",X"65",X"55",X"65",X"55",X"65",X"55",X"65",X"55",X"65",X"55",
		X"65",X"56",X"8A",X"A9",X"09",X"57",X"0A",X"55",X"02",X"55",X"02",X"95",X"00",X"95",X"00",X"A5",
		X"00",X"25",X"00",X"29",X"00",X"09",X"00",X"0A",X"00",X"02",X"00",X"02",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"EF",X"FF",X"FB",X"FF",X"FF",X"EA",X"FF",X"95",X"FF",X"95",X"FF",X"EA",X"FF",X"FF",
		X"00",X"00",X"A0",X"00",X"A8",X"00",X"AA",X"00",X"AA",X"80",X"AA",X"80",X"AA",X"A0",X"AA",X"A0",
		X"AA",X"A0",X"AA",X"A0",X"EA",X"A0",X"EA",X"A0",X"9A",X"A0",X"5A",X"A0",X"5A",X"A0",X"5A",X"A0",
		X"96",X"A0",X"96",X"A0",X"96",X"A0",X"96",X"A0",X"A6",X"A0",X"26",X"A0",X"26",X"A0",X"2A",X"A0",
		X"2A",X"A0",X"2A",X"A0",X"2A",X"A0",X"2A",X"A0",X"2A",X"A0",X"2A",X"A0",X"AA",X"A0",X"AA",X"A0",
		X"AA",X"A0",X"6A",X"A0",X"6A",X"A0",X"6A",X"A0",X"6A",X"A0",X"8A",X"A0",X"00",X"20",X"00",X"20",
		X"08",X"20",X"A8",X"20",X"80",X"20",X"82",X"80",X"A8",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"80",X"00",X"80",X"00",X"E0",X"00",X"78",X"00",X"58",X"00",X"5E",X"00",X"56",X"00",
		X"5E",X"00",X"5E",X"00",X"57",X"80",X"55",X"80",X"55",X"E0",X"95",X"60",X"95",X"78",X"25",X"5A",
		X"E9",X"56",X"AF",X"56",X"B5",X"56",X"F5",X"AB",X"56",X"FF",X"56",X"FF",X"AB",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"F5",X"0F",X"55",X"F5",X"55",
		X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"57",X"D7",X"57",X"FF",X"57",X"03",X"57",X"03",X"57",
		X"03",X"57",X"03",X"57",X"03",X"57",X"03",X"57",X"03",X"57",X"03",X"57",X"03",X"57",X"03",X"57",
		X"03",X"57",X"03",X"57",X"03",X"57",X"03",X"57",X"03",X"57",X"03",X"57",X"03",X"57",X"03",X"FF",
		X"00",X"0F",X"00",X"F7",X"0C",X"D7",X"FC",X"D7",X"5C",X"D7",X"5C",X"D7",X"5C",X"D7",X"5C",X"D5",
		X"5C",X"35",X"5C",X"35",X"7C",X"35",X"C0",X"35",X"00",X"35",X"00",X"35",X"00",X"35",X"00",X"35",
		X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",
		X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"FC",X"0F",X"5C",X"0D",X"5C",
		X"0D",X"57",X"0D",X"57",X"0D",X"57",X"0D",X"57",X"0D",X"57",X"0D",X"57",X"0D",X"57",X"0D",X"57",
		X"CD",X"57",X"CD",X"55",X"CD",X"55",X"CD",X"55",X"CD",X"55",X"F5",X"75",X"F5",X"75",X"75",X"75",
		X"75",X"75",X"75",X"75",X"55",X"75",X"55",X"75",X"55",X"CD",X"55",X"CD",X"55",X"CD",X"55",X"CD",
		X"57",X"0D",X"57",X"0D",X"57",X"03",X"57",X"03",X"57",X"03",X"57",X"03",X"57",X"03",X"FF",X"03",
		X"00",X"0C",X"00",X"FC",X"0F",X"5C",X"0D",X"5C",X"0D",X"5C",X"0D",X"5C",X"0D",X"5C",X"0D",X"5C",
		X"0D",X"5C",X"0D",X"5C",X"0D",X"5C",X"35",X"5C",X"35",X"5C",X"35",X"5C",X"35",X"5C",X"35",X"70",
		X"35",X"70",X"F5",X"70",X"F5",X"70",X"F5",X"70",X"D5",X"70",X"D5",X"70",X"D5",X"70",X"D5",X"70",
		X"55",X"70",X"55",X"70",X"55",X"70",X"55",X"70",X"55",X"C0",X"55",X"C0",X"55",X"C0",X"55",X"C0",
		X"55",X"C0",X"55",X"C0",X"55",X"C0",X"55",X"C0",X"55",X"C0",X"55",X"C0",X"55",X"C0",X"FF",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"3D",X"03",X"D5",X"0D",X"55",X"35",X"55",
		X"35",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"5F",
		X"D5",X"70",X"D5",X"C0",X"D5",X"C0",X"D5",X"C0",X"D5",X"C0",X"D5",X"C0",X"D5",X"C0",X"D5",X"C0",
		X"D5",X"C0",X"D5",X"C0",X"D5",X"C0",X"D5",X"C0",X"D5",X"C0",X"D5",X"C0",X"D5",X"C0",X"D5",X"C0",
		X"D5",X"C0",X"D5",X"C0",X"D5",X"C0",X"D5",X"C0",X"D5",X"7F",X"D5",X"55",X"D5",X"55",X"D5",X"55",
		X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"35",X"55",X"0F",X"FF",
		X"00",X"00",X"03",X"F0",X"3D",X"5C",X"D5",X"5C",X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"57",
		X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"57",
		X"D5",X"57",X"D5",X"57",X"D5",X"57",X"D5",X"57",X"D5",X"57",X"D5",X"57",X"D5",X"57",X"D5",X"57",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"D5",X"57",X"D5",X"57",X"D5",X"57",X"D5",X"57",X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"57",
		X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"5C",X"55",X"5C",X"55",X"70",X"FF",X"C0",
		X"FC",X"00",X"D7",X"F0",X"D5",X"5F",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",
		X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"FD",X"55",X"03",X"FD",X"00",X"0D",X"00",X"0D",
		X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",
		X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0F",
		X"00",X"00",X"00",X"00",X"C0",X"00",X"7F",X"00",X"55",X"FC",X"55",X"57",X"55",X"57",X"55",X"57",
		X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"57",X"57",X"D7",
		X"57",X"3F",X"57",X"00",X"57",X"00",X"57",X"00",X"57",X"00",X"57",X"00",X"57",X"00",X"57",X"00",
		X"57",X"00",X"57",X"00",X"57",X"00",X"57",X"00",X"57",X"00",X"57",X"00",X"57",X"00",X"57",X"00",
		X"57",X"00",X"57",X"00",X"57",X"00",X"57",X"00",X"57",X"00",X"57",X"00",X"57",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"00",X"35",X"FC",
		X"35",X"5C",X"35",X"5C",X"35",X"5C",X"35",X"5C",X"35",X"5C",X"35",X"5C",X"35",X"5C",X"35",X"5C",
		X"35",X"5C",X"35",X"5C",X"35",X"5C",X"35",X"5C",X"35",X"5C",X"35",X"5C",X"35",X"5C",X"3F",X"FC",
		X"00",X"00",X"0F",X"00",X"35",X"F0",X"D5",X"5F",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",
		X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"D5",X"D7",X"35",X"D7",X"0D",X"D7",X"0D",X"D7",X"0F",
		X"D7",X"00",X"D7",X"3C",X"D7",X"37",X"D7",X"35",X"D7",X"35",X"D7",X"35",X"D7",X"35",X"D7",X"35",
		X"D7",X"35",X"D7",X"3D",X"D7",X"0D",X"D7",X"0D",X"D7",X"0D",X"D7",X"0D",X"D5",X"F5",X"D5",X"55",
		X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"5F",X"35",X"73",X"0F",X"C3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"73",X"FC",X"73",X"57",X"73",X"55",
		X"73",X"55",X"73",X"55",X"73",X"55",X"73",X"55",X"73",X"55",X"73",X"55",X"73",X"55",X"73",X"5F",
		X"F3",X"5C",X"03",X"5C",X"C3",X"5C",X"73",X"5C",X"73",X"5F",X"73",X"55",X"73",X"55",X"73",X"55",
		X"73",X"55",X"73",X"5F",X"73",X"5C",X"73",X"5C",X"73",X"5C",X"73",X"5C",X"73",X"5C",X"73",X"5C",
		X"73",X"5F",X"73",X"55",X"73",X"55",X"73",X"55",X"73",X"55",X"73",X"55",X"73",X"55",X"F3",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"5F",X"00",
		X"57",X"3F",X"57",X"35",X"57",X"35",X"57",X"35",X"57",X"35",X"57",X"35",X"57",X"35",X"F7",X"35",
		X"0F",X"35",X"00",X"35",X"00",X"35",X"00",X"35",X"FF",X"35",X"57",X"35",X"57",X"35",X"57",X"35",
		X"57",X"35",X"57",X"35",X"FF",X"35",X"00",X"35",X"00",X"35",X"00",X"35",X"00",X"35",X"00",X"35",
		X"FF",X"35",X"57",X"35",X"57",X"35",X"57",X"35",X"57",X"35",X"57",X"35",X"57",X"35",X"FF",X"3F",
		X"00",X"00",X"F0",X"00",X"5C",X"00",X"57",X"00",X"55",X"C0",X"55",X"C3",X"55",X"7D",X"55",X"7D",
		X"55",X"7D",X"F5",X"7D",X"CD",X"7D",X"CD",X"7D",X"CD",X"7D",X"F5",X"7D",X"55",X"7D",X"55",X"7D",
		X"55",X"CD",X"57",X"0D",X"55",X"CD",X"F5",X"73",X"CD",X"70",X"CD",X"70",X"CD",X"7F",X"CD",X"7D",
		X"CD",X"7D",X"CD",X"7D",X"CD",X"7D",X"CD",X"7D",X"CD",X"7D",X"CD",X"73",X"CD",X"73",X"CD",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"00",X"57",X"F0",X"55",X"5C",X"55",X"57",
		X"55",X"57",X"55",X"57",X"55",X"57",X"5F",X"57",X"70",X"D7",X"70",X"FF",X"70",X"00",X"5C",X"00",
		X"57",X"FC",X"55",X"57",X"55",X"57",X"D5",X"57",X"3F",X"57",X"00",X"D7",X"F0",X"D7",X"70",X"D7",
		X"5F",X"57",X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"5C",X"55",X"5C",X"FF",X"F0",
		X"FC",X"00",X"FF",X"C0",X"AF",X"F0",X"FE",X"FC",X"FF",X"FF",X"FF",X"FC",X"FC",X"00",X"FF",X"C0",
		X"FF",X"C0",X"FC",X"00",X"FF",X"FC",X"FF",X"FF",X"FE",X"FC",X"AF",X"F0",X"FF",X"C0",X"FC",X"00",
		X"03",X"FF",X"00",X"3F",X"3F",X"FF",X"FF",X"FF",X"3F",X"BF",X"0F",X"FA",X"03",X"FF",X"00",X"3F",
		X"00",X"3F",X"0F",X"FF",X"3F",X"FA",X"FF",X"BF",X"FF",X"FF",X"3F",X"FF",X"0F",X"FF",X"03",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"2B",X"0A",X"BF",
		X"2F",X"FF",X"2F",X"FA",X"2E",X"A0",X"28",X"02",X"20",X"0B",X"BA",X"AF",X"BF",X"BA",X"2A",X"20",
		X"2E",X"8A",X"22",X"0F",X"22",X"00",X"08",X"00",X"0A",X"80",X"08",X"00",X"22",X"AA",X"20",X"2F",
		X"88",X"2F",X"80",X"0A",X"88",X"00",X"20",X"0A",X"0A",X"A0",X"00",X"00",X"08",X"00",X"22",X"00",
		X"20",X"80",X"82",X"20",X"80",X"20",X"80",X"A2",X"82",X"FB",X"82",X"FB",X"29",X"7B",X"09",X"7F",
		X"02",X"57",X"00",X"95",X"00",X"25",X"00",X"09",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"08",X"00",X"08",X"00",X"20",X"00",X"20",
		X"00",X"0A",X"00",X"09",X"00",X"09",X"00",X"09",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",
		X"FF",X"FF",X"FF",X"FA",X"FF",X"E7",X"FF",X"E5",X"FF",X"F9",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"E2",X"A0",X"EB",X"E0",
		X"FF",X"E0",X"BF",X"F8",X"2F",X"F8",X"0B",X"F8",X"82",X"FE",X"E2",X"F8",X"82",X"F8",X"02",X"FE",
		X"8B",X"FF",X"82",X"FF",X"00",X"BF",X"00",X"BF",X"00",X"BE",X"00",X"29",X"00",X"96",X"80",X"9B",
		X"82",X"AF",X"02",X"FF",X"0B",X"FF",X"AF",X"FF",X"2F",X"FF",X"2F",X"FF",X"0B",X"FF",X"0B",X"FF",
		X"2F",X"FF",X"2F",X"FF",X"BF",X"FF",X"BF",X"F9",X"BF",X"E5",X"BF",X"A5",X"FE",X"09",X"FE",X"02",
		X"F8",X"02",X"F8",X"02",X"E0",X"02",X"80",X"02",X"00",X"09",X"00",X"09",X"00",X"22",X"00",X"80",
		X"0A",X"00",X"20",X"00",X"80",X"00",X"00",X"01",X"00",X"05",X"00",X"55",X"01",X"6A",X"05",X"80",
		X"AA",X"00",X"56",X"00",X"5E",X"00",X"5E",X"00",X"57",X"82",X"57",X"A9",X"57",X"89",X"55",X"82",
		X"97",X"80",X"97",X"80",X"95",X"80",X"95",X"80",X"95",X"E0",X"25",X"E0",X"25",X"60",X"25",X"60",
		X"A5",X"6F",X"E5",X"6F",X"65",X"6F",X"55",X"6B",X"55",X"6E",X"A5",X"6F",X"FA",X"BF",X"FF",X"FF",
		X"80",X"00",X"80",X"00",X"80",X"28",X"82",X"BE",X"2B",X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"7F",X"FF",X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",X"5F",X"FA",
		X"AA",X"A0",X"00",X"02",X"AA",X"AB",X"77",X"FF",X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",X"9F",X"FF",
		X"97",X"FF",X"6B",X"FF",X"56",X"FF",X"55",X"AA",X"56",X"55",X"A9",X"56",X"05",X"58",X"15",X"60",
		X"55",X"80",X"56",X"00",X"6A",X"00",X"A5",X"80",X"9F",X"80",X"56",X"E0",X"55",X"F8",X"55",X"B8",
		X"95",X"5E",X"25",X"5E",X"09",X"56",X"09",X"55",X"02",X"55",X"00",X"A9",X"00",X"29",X"00",X"25",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"E8",X"00",X"FE",X"80",X"FF",X"E0",
		X"5F",X"F8",X"57",X"F6",X"9A",X"D6",X"2F",X"58",X"29",X"58",X"95",X"60",X"95",X"60",X"95",X"80",
		X"96",X"00",X"96",X"00",X"E8",X"00",X"E0",X"00",X"E0",X"00",X"E0",X"00",X"A0",X"00",X"20",X"00",
		X"E0",X"00",X"B8",X"00",X"FE",X"00",X"FE",X"00",X"EF",X"80",X"EF",X"80",X"EB",X"E0",X"EB",X"E0",
		X"EB",X"E0",X"9B",X"80",X"9A",X"00",X"A0",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"E0",X"00",X"78",X"00",X"58",X"00",
		X"56",X"FF",X"76",X"EB",X"76",X"FF",X"76",X"FF",X"56",X"EF",X"56",X"FF",X"AA",X"AB",X"FF",X"FF",
		X"6E",X"4A",X"FE",X"7A",X"01",X"C5",X"61",X"45",X"31",X"25",X"EA",X"49",X"2E",X"F9",X"75",X"FB",
		X"4D",X"C9",X"3B",X"39",X"27",X"7E",X"1C",X"3F",X"CC",X"7B",X"6E",X"49",X"FB",X"E5",X"49",X"A1",
		X"26",X"25",X"3B",X"B7",X"35",X"C9",X"1E",X"D9",X"47",X"69",X"2E",X"DE",X"0E",X"F8",X"FB",X"2B",
		X"C6",X"45",X"26",X"21",X"29",X"FB",X"4E",X"1E",X"44",X"B5",X"CE",X"42",X"6E",X"F9",X"09",X"19",
		X"22",X"71",X"45",X"36",X"D8",X"A9",X"2A",X"09",X"7A",X"E1",X"E9",X"29",X"EE",X"0E",X"D2",X"FB",
		X"02",X"39",X"49",X"C8",X"2F",X"75",X"28",X"CD",X"7E",X"F8",X"E6",X"F8",X"BD",X"6A",X"CD",X"F1",
		X"7A",X"E9",X"06",X"F8",X"B9",X"B5",X"08",X"9D",X"0C",X"74",X"69",X"09",X"21",X"4F",X"09",X"34",
		X"FE",X"3A",X"E7",X"11",X"E1",X"5A",X"48",X"FD",X"E2",X"38",X"66",X"21",X"E5",X"FA",X"FB",X"DD",
		X"C9",X"07",X"0B",X"85",X"66",X"D9",X"7A",X"F9",X"C5",X"4A",X"62",X"F8",X"0E",X"31",X"E5",X"0A",
		X"35",X"03",X"26",X"E9",X"47",X"C9",X"39",X"39",X"ED",X"C2",X"01",X"F0",X"EC",X"DA",X"6C",X"41",
		X"ED",X"03",X"2A",X"A7",X"65",X"99",X"39",X"F9",X"C8",X"C9",X"06",X"B9",X"66",X"BA",X"2F",X"F8",
		X"E1",X"07",X"47",X"BB",X"C6",X"89",X"6A",X"99",X"68",X"E1",X"E3",X"F3",X"A6",X"11",X"A5",X"79",
		X"F9",X"CD",X"16",X"C5",X"3C",X"18",X"69",X"3B",X"EA",X"D9",X"F8",X"0A",X"05",X"F1",X"E6",X"15",
		X"7E",X"00",X"78",X"39",X"09",X"3B",X"4D",X"C9",X"02",X"E9",X"39",X"BB",X"C6",X"F4",X"AE",X"C9",
		X"4B",X"2B",X"B9",X"3A",X"7E",X"F9",X"86",X"F1",X"FA",X"83",X"34",X"01",X"6A",X"79",X"EC",X"FD",
		X"6D",X"E7",X"67",X"FB",X"6E",X"29",X"F9",X"2D",X"75",X"37",X"33",X"4B",X"3F",X"D1",X"22",X"39");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
