library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity obj1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of obj1 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"04",X"1C",X"3D",X"3F",X"3F",X"3F",X"3F",X"3F",X"1E",X"1E",X"1C",X"08",X"00",X"00",
		X"00",X"00",X"05",X"1D",X"3D",X"3F",X"3E",X"3E",X"3F",X"3F",X"1E",X"1E",X"1C",X"09",X"01",X"00",
		X"00",X"00",X"00",X"02",X"0E",X"1E",X"1F",X"1F",X"1F",X"1F",X"1F",X"0F",X"0F",X"0E",X"04",X"00",
		X"00",X"03",X"07",X"07",X"1F",X"3C",X"1F",X"1F",X"1F",X"1F",X"3C",X"FF",X"FF",X"1C",X"00",X"00",
		X"00",X"10",X"30",X"20",X"40",X"60",X"70",X"70",X"60",X"40",X"70",X"30",X"18",X"1C",X"0C",X"00",
		X"00",X"03",X"04",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"03",X"1B",X"3C",X"1F",X"1F",X"1F",X"1F",X"3C",X"1B",X"03",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"04",X"1C",X"3D",X"3F",X"FF",X"FF",X"FF",X"3E",X"1E",X"1E",X"1C",X"08",X"00",X"00",
		X"00",X"00",X"04",X"1C",X"3D",X"3F",X"3F",X"3E",X"3E",X"3F",X"1E",X"1E",X"1C",X"08",X"00",X"00",
		X"00",X"00",X"04",X"1C",X"3D",X"3F",X"FF",X"FF",X"FF",X"3E",X"1E",X"1E",X"1C",X"08",X"00",X"00",
		X"00",X"00",X"04",X"1C",X"3C",X"3F",X"3F",X"3E",X"3E",X"3F",X"1E",X"1E",X"1C",X"08",X"00",X"00",
		X"00",X"00",X"00",X"02",X"0E",X"1E",X"1F",X"FF",X"FF",X"FF",X"1F",X"0F",X"0F",X"0E",X"04",X"00",
		X"00",X"00",X"00",X"02",X"0E",X"1E",X"1F",X"1F",X"1F",X"1F",X"1F",X"0F",X"0F",X"0E",X"04",X"00",
		X"00",X"01",X"01",X"02",X"0E",X"1E",X"1F",X"1F",X"1F",X"1F",X"1F",X"0F",X"0F",X"0E",X"05",X"01",
		X"01",X"03",X"07",X"1F",X"3F",X"3F",X"3E",X"3F",X"3F",X"3F",X"1F",X"1F",X"1D",X"09",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"67",X"7F",X"FF",X"FF",X"FF",X"FF",X"9E",X"1C",X"0D",X"09",X"03",X"06",X"04",
		X"01",X"01",X"21",X"6C",X"FE",X"FE",X"FE",X"FF",X"FF",X"BF",X"DE",X"66",X"20",X"00",X"00",X"00",
		X"00",X"00",X"27",X"77",X"DF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"5F",X"77",X"27",X"00",X"00",
		X"00",X"00",X"06",X"0E",X"1D",X"1B",X"1B",X"1B",X"1A",X"1A",X"1B",X"0A",X"03",X"03",X"03",X"01",
		X"00",X"00",X"03",X"04",X"08",X"0A",X"11",X"10",X"10",X"16",X"0E",X"08",X"04",X"03",X"00",X"00",
		X"02",X"0F",X"04",X"04",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"04",X"04",X"0F",X"02",
		X"05",X"0F",X"0B",X"1B",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"1B",X"0B",X"0F",X"05",
		X"00",X"00",X"00",X"00",X"4F",X"7F",X"C0",X"40",X"40",X"C0",X"7F",X"4F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"03",X"00",X"00",X"00",
		X"05",X"0F",X"0B",X"1B",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"1B",X"0B",X"0F",X"05",
		X"02",X"0F",X"04",X"04",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"04",X"04",X"0F",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"00",
		X"1F",X"3F",X"7F",X"FF",X"FF",X"BF",X"9E",X"C1",X"E1",X"C6",X"8F",X"CF",X"E6",X"73",X"1F",X"00",
		X"1F",X"3F",X"7F",X"FF",X"FF",X"BF",X"9E",X"C1",X"E1",X"C6",X"8F",X"CF",X"E6",X"73",X"1F",X"00",
		X"1F",X"3F",X"7F",X"FF",X"FF",X"BF",X"9E",X"C1",X"E1",X"C6",X"8F",X"CF",X"E6",X"73",X"1F",X"00",
		X"00",X"1E",X"36",X"60",X"C0",X"CC",X"ED",X"F1",X"ED",X"CC",X"C0",X"60",X"36",X"1E",X"0E",X"00",
		X"00",X"1E",X"36",X"60",X"C0",X"CC",X"ED",X"F1",X"ED",X"CC",X"C0",X"60",X"36",X"1E",X"0E",X"00",
		X"FE",X"47",X"87",X"14",X"85",X"04",X"89",X"F0",X"F0",X"89",X"04",X"85",X"14",X"87",X"47",X"FE",
		X"00",X"01",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"03",X"87",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",
		X"01",X"0F",X"07",X"0F",X"07",X"23",X"13",X"09",X"51",X"31",X"11",X"01",X"01",X"03",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"11",X"1F",X"1F",X"1F",X"0F",X"0F",X"07",X"03",X"03",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"07",X"07",X"03",X"01",X"01",
		X"00",X"00",X"00",X"00",X"C0",X"F8",X"FE",X"FF",X"FF",X"FF",X"FF",X"EE",X"FF",X"FC",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"0F",X"1F",X"3F",X"7F",
		X"F4",X"F9",X"FD",X"FE",X"FF",X"FF",X"FF",X"FF",X"3F",X"0F",X"07",X"01",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E6",X"E2",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"07",X"0F",X"0F",X"0F",X"1F",X"1F",X"1F",X"1F",
		X"3C",X"78",X"78",X"FC",X"F7",X"E3",X"E1",X"C0",X"CC",X"4C",X"00",X"04",X"04",X"00",X"00",X"00",
		X"00",X"00",X"01",X"01",X"03",X"03",X"03",X"07",X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"0C",X"08",
		X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",X"0F",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"0F",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",
		X"00",X"20",X"5C",X"7F",X"FF",X"7F",X"7F",X"1F",X"0F",X"07",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"03",X"07",X"07",X"07",X"0F",X"0F",X"07",X"07",X"0B",X"00",X"00",X"00",X"00",
		X"FC",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"1F",X"0E",X"00",X"00",
		X"00",X"1C",X"3E",X"7F",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"08",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"40",X"61",X"63",X"66",X"6C",X"7A",X"7A",X"6C",X"66",X"63",X"61",X"40",X"00",X"00",
		X"00",X"00",X"04",X"06",X"06",X"06",X"06",X"07",X"07",X"06",X"06",X"06",X"06",X"04",X"00",X"00",
		X"00",X"10",X"08",X"00",X"00",X"00",X"00",X"01",X"00",X"21",X"00",X"00",X"04",X"00",X"00",X"00",
		X"08",X"00",X"00",X"00",X"00",X"01",X"23",X"03",X"05",X"01",X"02",X"00",X"10",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"00",X"01",X"24",X"00",X"00",X"05",X"08",X"40",X"00",X"00",X"00",X"04",X"00",X"00",X"00",
		X"02",X"08",X"40",X"20",X"04",X"40",X"01",X"04",X"08",X"00",X"02",X"00",X"00",X"00",X"00",X"00",
		X"80",X"10",X"08",X"04",X"06",X"03",X"10",X"2F",X"03",X"01",X"01",X"0A",X"05",X"00",X"00",X"20",
		X"01",X"40",X"00",X"00",X"02",X"01",X"00",X"00",X"01",X"03",X"06",X"00",X"10",X"01",X"00",X"10",
		X"08",X"08",X"09",X"0B",X"0A",X"0B",X"09",X"08",X"08",X"08",X"09",X"0B",X"0A",X"0B",X"09",X"08",
		X"F7",X"F7",X"F7",X"F7",X"FB",X"FD",X"CE",X"B6",X"B6",X"CE",X"FD",X"FB",X"F7",X"F7",X"F7",X"F7",
		X"00",X"00",X"00",X"FF",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"F7",X"F7",X"F4",X"F4",X"F7",X"F4",X"F4",X"F7",X"F4",X"F5",X"F4",X"F7",X"FF",X"F7",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"01",X"02",X"0A",X"08",X"05",X"00",X"05",X"05",X"02",X"00",X"01",X"00",
		X"0F",X"0F",X"1F",X"1E",X"1E",X"3E",X"3C",X"3C",X"7C",X"78",X"79",X"FE",X"FE",X"70",X"30",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"06",X"07",X"06",X"03",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"06",X"07",X"06",X"03",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"1F",X"1F",X"1F",X"1C",X"1C",X"1E",X"1F",X"0F",X"0F",X"07",X"03",X"00",X"00",
		X"00",X"00",X"00",X"1F",X"1F",X"1E",X"1E",X"1E",X"1E",X"1E",X"0E",X"0F",X"07",X"03",X"00",X"00",
		X"00",X"00",X"00",X"1F",X"1F",X"1F",X"1F",X"1E",X"1C",X"1C",X"0F",X"0F",X"07",X"03",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"04",X"08",X"10",X"20",X"20",X"20",X"20",X"20",X"20",X"10",X"08",X"04",X"03",X"00",
		X"00",X"00",X"00",X"01",X"02",X"05",X"0A",X"0A",X"0A",X"0A",X"05",X"02",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"05",X"05",X"02",X"01",X"00",X"00",X"00",X"00",X"00",
		X"40",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"20",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"02",X"02",X"02",X"02",X"01",X"00",X"00",X"00",X"00",
		X"07",X"0F",X"18",X"30",X"20",X"47",X"1E",X"FE",X"FE",X"1E",X"47",X"20",X"30",X"18",X"0F",X"07",
		X"0F",X"1F",X"3F",X"3F",X"3F",X"3F",X"1F",X"0F",X"1F",X"3F",X"3F",X"3F",X"3F",X"1F",X"0F",X"00",
		X"0F",X"1F",X"3F",X"3F",X"3F",X"3F",X"1D",X"08",X"02",X"17",X"3F",X"3F",X"3F",X"3F",X"1F",X"0F",
		X"03",X"07",X"0F",X"3C",X"3D",X"3E",X"3F",X"3D",X"3D",X"3F",X"3E",X"3D",X"3C",X"0F",X"07",X"03",
		X"00",X"00",X"07",X"0F",X"1F",X"5F",X"E6",X"ED",X"7D",X"08",X"02",X"30",X"38",X"3C",X"3C",X"1C",
		X"20",X"50",X"88",X"88",X"88",X"88",X"88",X"56",X"26",X"0C",X"0C",X"0C",X"0C",X"00",X"00",X"00",
		X"07",X"08",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"08",X"07",X"00",X"00",X"0F",X"04",X"00",
		X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"07",X"00",X"06",X"09",X"08",X"08",X"04",X"00",
		X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"07",X"00",X"08",X"0D",X"0B",X"09",X"08",X"00",
		X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"07",X"00",X"09",X"0A",X"0A",X"0A",X"0E",X"00",
		X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"07",X"00",X"06",X"09",X"09",X"09",X"06",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
