library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity monitor is
    generic(
        AddrWidth   : integer := 11
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(AddrWidth-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end monitor;

architecture rtl of monitor is
    type rom2048x8 is array (0 to 2**AddrWidth-1) of std_logic_vector(7 downto 0); 
    constant romData : rom2048x8 := (
         x"C3",  x"0C",  x"00",  x"4D",  x"4F",  x"4E",  x"20",  x"20", -- 0000
         x"20",  x"20",  x"20",  x"00",  x"31",  x"C0",  x"EB",  x"CD", -- 0008
         x"C7",  x"06",  x"CD",  x"D7",  x"00",  x"C3",  x"03",  x"F0", -- 0010
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0018
         x"3E",  x"02",  x"CF",  x"C9",  x"3E",  x"00",  x"CF",  x"76", -- 0020
         x"18",  x"FD",  x"C1",  x"E1",  x"31",  x"00",  x"02",  x"E9", -- 0028
         x"C9",  x"2A",  x"2A",  x"2A",  x"20",  x"4D",  x"6F",  x"6E", -- 0030
         x"69",  x"74",  x"6F",  x"72",  x"20",  x"56",  x"30",  x"2E", -- 0038
         x"30",  x"30",  x"31",  x"20",  x"2A",  x"2A",  x"2A",  x"0A", -- 0040
         x"00",  x"FD",  x"21",  x"02",  x"00",  x"FD",  x"39",  x"FD", -- 0048
         x"66",  x"00",  x"7C",  x"57",  x"D6",  x"30",  x"38",  x"0A", -- 0050
         x"3E",  x"39",  x"94",  x"38",  x"05",  x"7A",  x"C6",  x"D0", -- 0058
         x"6F",  x"C9",  x"7C",  x"D6",  x"41",  x"38",  x"0A",  x"3E", -- 0060
         x"46",  x"94",  x"38",  x"05",  x"7A",  x"C6",  x"C9",  x"6F", -- 0068
         x"C9",  x"7C",  x"D6",  x"61",  x"38",  x"0A",  x"3E",  x"66", -- 0070
         x"94",  x"38",  x"05",  x"7A",  x"C6",  x"A9",  x"6F",  x"C9", -- 0078
         x"2E",  x"FF",  x"C9",  x"3E",  x"3E",  x"F5",  x"33",  x"CD", -- 0080
         x"BE",  x"03",  x"33",  x"C1",  x"E1",  x"E5",  x"C5",  x"2E", -- 0088
         x"00",  x"E5",  x"33",  x"CD",  x"0B",  x"04",  x"33",  x"FD", -- 0090
         x"21",  x"02",  x"00",  x"FD",  x"39",  x"FD",  x"66",  x"00", -- 0098
         x"E5",  x"33",  x"CD",  x"0B",  x"04",  x"33",  x"3E",  x"0A", -- 00A0
         x"F5",  x"33",  x"CD",  x"BE",  x"03",  x"33",  x"C9",  x"DD", -- 00A8
         x"E5",  x"DD",  x"21",  x"00",  x"00",  x"DD",  x"39",  x"DD", -- 00B0
         x"6E",  x"04",  x"DD",  x"66",  x"05",  x"E5",  x"56",  x"23", -- 00B8
         x"5E",  x"E1",  x"7A",  x"E6",  x"03",  x"28",  x"04",  x"D6", -- 00C0
         x"03",  x"20",  x"02",  x"CB",  x"FB",  x"CB",  x"3B",  x"CB", -- 00C8
         x"1A",  x"72",  x"23",  x"73",  x"DD",  x"E1",  x"C9",  x"DD", -- 00D0
         x"E5",  x"DD",  x"21",  x"00",  x"00",  x"DD",  x"39",  x"21", -- 00D8
         x"EE",  x"FF",  x"39",  x"F9",  x"DD",  x"36",  x"F6",  x"D2", -- 00E0
         x"DD",  x"36",  x"F7",  x"04",  x"DD",  x"36",  x"F4",  x"D2", -- 00E8
         x"DD",  x"36",  x"F5",  x"04",  x"DD",  x"36",  x"F2",  x"00", -- 00F0
         x"DD",  x"36",  x"F3",  x"00",  x"DD",  x"36",  x"F1",  x"01", -- 00F8
         x"DD",  x"36",  x"F0",  x"00",  x"DD",  x"36",  x"EF",  x"00", -- 0100
         x"DD",  x"36",  x"EE",  x"00",  x"DD",  x"36",  x"F8",  x"00", -- 0108
         x"21",  x"31",  x"00",  x"E5",  x"CD",  x"D4",  x"03",  x"F1", -- 0110
         x"CD",  x"CB",  x"03",  x"DD",  x"75",  x"FF",  x"7D",  x"B7", -- 0118
         x"28",  x"F6",  x"DD",  x"66",  x"FF",  x"7C",  x"FE",  x"0A", -- 0120
         x"CA",  x"C6",  x"01",  x"FE",  x"0D",  x"CA",  x"C6",  x"01", -- 0128
         x"FE",  x"3A",  x"CA",  x"DE",  x"01",  x"FE",  x"67",  x"28", -- 0130
         x"72",  x"FE",  x"6B",  x"CA",  x"B8",  x"01",  x"D6",  x"6D", -- 0138
         x"CA",  x"E5",  x"01",  x"7C",  x"FE",  x"70",  x"28",  x"55", -- 0140
         x"D6",  x"72",  x"28",  x"3F",  x"DD",  x"7E",  x"F2",  x"C6", -- 0148
         x"01",  x"DD",  x"77",  x"FD",  x"DD",  x"7E",  x"F3",  x"CE", -- 0150
         x"00",  x"DD",  x"77",  x"FE",  x"7C",  x"FE",  x"73",  x"28", -- 0158
         x"0F",  x"D6",  x"74",  x"C2",  x"97",  x"02",  x"DD",  x"36", -- 0160
         x"EF",  x"01",  x"DD",  x"36",  x"F1",  x"01",  x"18",  x"A8", -- 0168
         x"DD",  x"6E",  x"F2",  x"DD",  x"66",  x"F3",  x"66",  x"DD", -- 0170
         x"7E",  x"FD",  x"DD",  x"77",  x"F2",  x"DD",  x"7E",  x"FE", -- 0178
         x"DD",  x"77",  x"F3",  x"E5",  x"33",  x"CD",  x"0B",  x"04", -- 0180
         x"33",  x"18",  x"8D",  x"3E",  x"05",  x"D3",  x"02",  x"DD", -- 0188
         x"6E",  x"F2",  x"DD",  x"66",  x"F3",  x"E5",  x"CD",  x"2A", -- 0190
         x"00",  x"F1",  x"C3",  x"18",  x"01",  x"DD",  x"6E",  x"F2", -- 0198
         x"DD",  x"66",  x"F3",  x"E5",  x"CD",  x"83",  x"00",  x"F1", -- 01A0
         x"C3",  x"18",  x"01",  x"3E",  x"05",  x"D3",  x"02",  x"31", -- 01A8
         x"00",  x"02",  x"C3",  x"89",  x"F0",  x"C3",  x"18",  x"01", -- 01B0
         x"DD",  x"6E",  x"F2",  x"DD",  x"66",  x"F3",  x"E5",  x"CD", -- 01B8
         x"14",  x"06",  x"F1",  x"C3",  x"18",  x"01",  x"DD",  x"36", -- 01C0
         x"EE",  x"00",  x"DD",  x"36",  x"EF",  x"00",  x"DD",  x"36", -- 01C8
         x"F8",  x"00",  x"DD",  x"7E",  x"FF",  x"F5",  x"33",  x"CD", -- 01D0
         x"BE",  x"03",  x"33",  x"C3",  x"18",  x"01",  x"DD",  x"36", -- 01D8
         x"EE",  x"02",  x"C3",  x"18",  x"01",  x"F3",  x"DD",  x"36", -- 01E0
         x"FB",  x"00",  x"DD",  x"36",  x"FC",  x"00",  x"11",  x"00", -- 01E8
         x"40",  x"7A",  x"D6",  x"80",  x"30",  x"12",  x"21",  x"08", -- 01F0
         x"00",  x"39",  x"D5",  x"E5",  x"CD",  x"AF",  x"00",  x"F1", -- 01F8
         x"D1",  x"DD",  x"7E",  x"F6",  x"12",  x"13",  x"18",  x"E9", -- 0200
         x"DD",  x"36",  x"F2",  x"00",  x"DD",  x"36",  x"F3",  x"40", -- 0208
         x"DD",  x"7E",  x"F3",  x"D6",  x"80",  x"30",  x"59",  x"21", -- 0210
         x"06",  x"00",  x"39",  x"E5",  x"CD",  x"AF",  x"00",  x"F1", -- 0218
         x"DD",  x"6E",  x"F2",  x"DD",  x"66",  x"F3",  x"56",  x"DD", -- 0220
         x"5E",  x"F4",  x"7A",  x"93",  x"28",  x"38",  x"DD",  x"6E", -- 0228
         x"F2",  x"DD",  x"66",  x"F3",  x"E5",  x"CD",  x"83",  x"00", -- 0230
         x"26",  x"20",  x"E3",  x"33",  x"CD",  x"BE",  x"03",  x"33", -- 0238
         x"DD",  x"6E",  x"F2",  x"DD",  x"66",  x"F3",  x"66",  x"E5", -- 0240
         x"33",  x"CD",  x"0B",  x"04",  x"33",  x"3E",  x"20",  x"F5", -- 0248
         x"33",  x"CD",  x"BE",  x"03",  x"33",  x"DD",  x"66",  x"F4", -- 0250
         x"E5",  x"33",  x"CD",  x"0B",  x"04",  x"33",  x"3E",  x"0A", -- 0258
         x"F5",  x"33",  x"CD",  x"BE",  x"03",  x"33",  x"DD",  x"34", -- 0260
         x"F2",  x"20",  x"A5",  x"DD",  x"34",  x"F3",  x"18",  x"A0", -- 0268
         x"DD",  x"66",  x"FC",  x"2E",  x"00",  x"E5",  x"33",  x"CD", -- 0270
         x"0B",  x"04",  x"33",  x"DD",  x"66",  x"FB",  x"E5",  x"33", -- 0278
         x"CD",  x"0B",  x"04",  x"33",  x"DD",  x"34",  x"FB",  x"20", -- 0280
         x"03",  x"DD",  x"34",  x"FC",  x"21",  x"B9",  x"03",  x"E5", -- 0288
         x"CD",  x"D4",  x"03",  x"F1",  x"C3",  x"EE",  x"01",  x"DD", -- 0290
         x"7E",  x"FF",  x"F5",  x"33",  x"CD",  x"49",  x"00",  x"33", -- 0298
         x"7D",  x"3C",  x"CA",  x"18",  x"01",  x"DD",  x"7E",  x"F0", -- 02A0
         x"07",  x"07",  x"07",  x"07",  x"E6",  x"F0",  x"4F",  x"09", -- 02A8
         x"DD",  x"75",  x"F0",  x"DD",  x"7E",  x"F1",  x"D6",  x"02", -- 02B0
         x"20",  x"04",  x"3E",  x"01",  x"18",  x"01",  x"AF",  x"DD", -- 02B8
         x"77",  x"FB",  x"DD",  x"7E",  x"EF",  x"3D",  x"20",  x"5F", -- 02C0
         x"DD",  x"7E",  x"FB",  x"B7",  x"28",  x"21",  x"DD",  x"7E", -- 02C8
         x"F0",  x"DD",  x"77",  x"F9",  x"DD",  x"36",  x"FA",  x"00", -- 02D0
         x"DD",  x"7E",  x"F9",  x"DD",  x"77",  x"FA",  x"DD",  x"36", -- 02D8
         x"F9",  x"00",  x"DD",  x"36",  x"F2",  x"00",  x"DD",  x"7E", -- 02E0
         x"FA",  x"DD",  x"77",  x"F3",  x"C3",  x"B3",  x"03",  x"DD", -- 02E8
         x"7E",  x"F1",  x"D6",  x"04",  x"C2",  x"B3",  x"03",  x"DD", -- 02F0
         x"36",  x"F1",  x"00",  x"DD",  x"7E",  x"F2",  x"DD",  x"86", -- 02F8
         x"F0",  x"DD",  x"77",  x"F2",  x"DD",  x"7E",  x"F3",  x"CE", -- 0300
         x"00",  x"DD",  x"77",  x"F3",  x"3E",  x"3E",  x"F5",  x"33", -- 0308
         x"CD",  x"BE",  x"03",  x"33",  x"DD",  x"36",  x"EF",  x"00", -- 0310
         x"DD",  x"7E",  x"EE",  x"D6",  x"03",  x"C2",  x"B3",  x"03", -- 0318
         x"DD",  x"36",  x"EE",  x"04",  x"C3",  x"B3",  x"03",  x"DD", -- 0320
         x"7E",  x"FB",  x"B7",  x"CA",  x"B3",  x"03",  x"DD",  x"36", -- 0328
         x"F1",  x"00",  x"DD",  x"7E",  x"EE",  x"D6",  x"02",  x"28", -- 0330
         x"17",  x"DD",  x"7E",  x"EE",  x"D6",  x"04",  x"28",  x"28", -- 0338
         x"DD",  x"7E",  x"EE",  x"D6",  x"05",  x"28",  x"3B",  x"DD", -- 0340
         x"7E",  x"EE",  x"D6",  x"06",  x"28",  x"2A",  x"18",  x"45", -- 0348
         x"3E",  x"2A",  x"F5",  x"33",  x"CD",  x"BE",  x"03",  x"33", -- 0350
         x"DD",  x"7E",  x"F0",  x"DD",  x"77",  x"F8",  x"DD",  x"36", -- 0358
         x"EF",  x"01",  x"DD",  x"36",  x"EE",  x"03",  x"18",  x"4B", -- 0360
         x"DD",  x"36",  x"EE",  x"05",  x"DD",  x"7E",  x"F0",  x"B7", -- 0368
         x"28",  x"41",  x"DD",  x"36",  x"EE",  x"06",  x"18",  x"3B", -- 0370
         x"3E",  x"3A",  x"F5",  x"33",  x"CD",  x"BE",  x"03",  x"33", -- 0378
         x"18",  x"31",  x"DD",  x"7E",  x"F8",  x"B7",  x"20",  x"0A", -- 0380
         x"3E",  x"2D",  x"F5",  x"33",  x"CD",  x"BE",  x"03",  x"33", -- 0388
         x"18",  x"21",  x"DD",  x"35",  x"F8",  x"DD",  x"6E",  x"F2", -- 0390
         x"DD",  x"66",  x"F3",  x"DD",  x"7E",  x"F0",  x"77",  x"DD", -- 0398
         x"7E",  x"FD",  x"DD",  x"77",  x"F2",  x"DD",  x"7E",  x"FE", -- 03A0
         x"DD",  x"77",  x"F3",  x"3E",  x"2E",  x"F5",  x"33",  x"CD", -- 03A8
         x"BE",  x"03",  x"33",  x"DD",  x"34",  x"F1",  x"C3",  x"18", -- 03B0
         x"01",  x"20",  x"4F",  x"6B",  x"0A",  x"00",  x"DB",  x"00", -- 03B8
         x"B7",  x"20",  x"FB",  x"21",  x"02",  x"00",  x"39",  x"7E", -- 03C0
         x"D3",  x"00",  x"C9",  x"DB",  x"01",  x"B7",  x"28",  x"02", -- 03C8
         x"D3",  x"01",  x"6F",  x"C9",  x"C1",  x"E1",  x"E5",  x"C5", -- 03D0
         x"7E",  x"B7",  x"C8",  x"23",  x"E5",  x"F5",  x"33",  x"CD", -- 03D8
         x"BE",  x"03",  x"33",  x"E1",  x"18",  x"F2",  x"C9",  x"FD", -- 03E0
         x"21",  x"02",  x"00",  x"FD",  x"39",  x"FD",  x"56",  x"00", -- 03E8
         x"FD",  x"7E",  x"00",  x"D6",  x"0A",  x"30",  x"0A",  x"7A", -- 03F0
         x"C6",  x"30",  x"F5",  x"33",  x"CD",  x"BE",  x"03",  x"33", -- 03F8
         x"C9",  x"7A",  x"C6",  x"37",  x"F5",  x"33",  x"CD",  x"BE", -- 0400
         x"03",  x"33",  x"C9",  x"21",  x"02",  x"00",  x"39",  x"7E", -- 0408
         x"07",  x"07",  x"07",  x"07",  x"E6",  x"0F",  x"F5",  x"33", -- 0410
         x"CD",  x"E7",  x"03",  x"33",  x"21",  x"02",  x"00",  x"39", -- 0418
         x"7E",  x"E6",  x"0F",  x"F5",  x"33",  x"CD",  x"E7",  x"03", -- 0420
         x"33",  x"C9",  x"FD",  x"21",  x"02",  x"00",  x"FD",  x"39", -- 0428
         x"FD",  x"66",  x"01",  x"2E",  x"00",  x"E5",  x"33",  x"CD", -- 0430
         x"0B",  x"04",  x"33",  x"FD",  x"21",  x"02",  x"00",  x"FD", -- 0438
         x"39",  x"FD",  x"66",  x"00",  x"E5",  x"33",  x"CD",  x"0B", -- 0440
         x"04",  x"33",  x"C9",  x"21",  x"25",  x"00",  x"56",  x"7A", -- 0448
         x"B7",  x"28",  x"05",  x"21",  x"25",  x"00",  x"36",  x"00", -- 0450
         x"6A",  x"C9",  x"21",  x"00",  x"B0",  x"36",  x"00",  x"21", -- 0458
         x"00",  x"EC",  x"36",  x"20",  x"5D",  x"54",  x"13",  x"01", -- 0460
         x"BF",  x"03",  x"ED",  x"B0",  x"21",  x"00",  x"E8",  x"36", -- 0468
         x"20",  x"5D",  x"54",  x"13",  x"01",  x"BF",  x"03",  x"ED", -- 0470
         x"B0",  x"C9",  x"21",  x"02",  x"00",  x"39",  x"7E",  x"32", -- 0478
         x"00",  x"B0",  x"C9",  x"DD",  x"E5",  x"DD",  x"21",  x"00", -- 0480
         x"00",  x"DD",  x"39",  x"ED",  x"4B",  x"00",  x"B0",  x"06", -- 0488
         x"00",  x"69",  x"60",  x"29",  x"29",  x"09",  x"29",  x"29", -- 0490
         x"29",  x"11",  x"00",  x"E8",  x"19",  x"DD",  x"5E",  x"04", -- 0498
         x"16",  x"00",  x"D5",  x"01",  x"02",  x"00",  x"C5",  x"E5", -- 04A0
         x"CD",  x"9B",  x"06",  x"F1",  x"F1",  x"F1",  x"DD",  x"E1", -- 04A8
         x"C9",  x"DD",  x"E5",  x"DD",  x"21",  x"00",  x"00",  x"DD", -- 04B0
         x"39",  x"ED",  x"4B",  x"00",  x"B0",  x"06",  x"00",  x"69", -- 04B8
         x"60",  x"29",  x"29",  x"09",  x"29",  x"29",  x"29",  x"11", -- 04C0
         x"00",  x"E8",  x"19",  x"DD",  x"5E",  x"04",  x"16",  x"00", -- 04C8
         x"D5",  x"01",  x"20",  x"00",  x"C5",  x"E5",  x"CD",  x"9B", -- 04D0
         x"06",  x"F1",  x"F1",  x"F1",  x"DD",  x"E1",  x"C9",  x"DD", -- 04D8
         x"E5",  x"DD",  x"21",  x"00",  x"00",  x"DD",  x"39",  x"F5", -- 04E0
         x"F5",  x"ED",  x"4B",  x"00",  x"B0",  x"06",  x"00",  x"69", -- 04E8
         x"60",  x"29",  x"29",  x"09",  x"29",  x"29",  x"29",  x"11", -- 04F0
         x"00",  x"EC",  x"19",  x"33",  x"33",  x"E5",  x"DD",  x"7E", -- 04F8
         x"04",  x"DD",  x"77",  x"FE",  x"DD",  x"7E",  x"05",  x"DD", -- 0500
         x"77",  x"FF",  x"DD",  x"6E",  x"FE",  x"DD",  x"66",  x"FF", -- 0508
         x"7E",  x"B7",  x"28",  x"55",  x"DD",  x"34",  x"FE",  x"20", -- 0510
         x"03",  x"DD",  x"34",  x"FF",  x"5F",  x"D6",  x"09",  x"28", -- 0518
         x"20",  x"7B",  x"D6",  x"0A",  x"20",  x"36",  x"11",  x"00", -- 0520
         x"EC",  x"21",  x"00",  x"B0",  x"34",  x"ED",  x"4B",  x"00", -- 0528
         x"B0",  x"06",  x"00",  x"69",  x"60",  x"29",  x"29",  x"09", -- 0530
         x"29",  x"29",  x"29",  x"19",  x"33",  x"33",  x"E5",  x"18", -- 0538
         x"C9",  x"ED",  x"4B",  x"00",  x"B0",  x"06",  x"00",  x"69", -- 0540
         x"60",  x"29",  x"29",  x"09",  x"29",  x"29",  x"29",  x"11", -- 0548
         x"00",  x"EC",  x"19",  x"01",  x"0F",  x"00",  x"09",  x"33", -- 0550
         x"33",  x"E5",  x"18",  x"AE",  x"E1",  x"E5",  x"73",  x"DD", -- 0558
         x"34",  x"FC",  x"20",  x"A6",  x"DD",  x"34",  x"FD",  x"18", -- 0560
         x"A1",  x"3E",  x"17",  x"FD",  x"21",  x"00",  x"B0",  x"FD", -- 0568
         x"96",  x"00",  x"30",  x"05",  x"21",  x"00",  x"B0",  x"36", -- 0570
         x"00",  x"DD",  x"F9",  x"DD",  x"E1",  x"C9",  x"DD",  x"E5", -- 0578
         x"DD",  x"21",  x"00",  x"00",  x"DD",  x"39",  x"3B",  x"ED", -- 0580
         x"4B",  x"00",  x"B0",  x"06",  x"00",  x"69",  x"60",  x"29", -- 0588
         x"29",  x"09",  x"29",  x"29",  x"29",  x"11",  x"00",  x"EC", -- 0590
         x"19",  x"01",  x"12",  x"00",  x"09",  x"DD",  x"36",  x"FF", -- 0598
         x"00",  x"DD",  x"7E",  x"04",  x"E6",  x"0F",  x"4F",  x"5D", -- 05A0
         x"54",  x"1B",  x"79",  x"47",  x"D6",  x"0A",  x"30",  x"07", -- 05A8
         x"78",  x"C6",  x"30",  x"77",  x"EB",  x"18",  x"05",  x"78", -- 05B0
         x"C6",  x"37",  x"77",  x"EB",  x"06",  x"04",  x"DD",  x"CB", -- 05B8
         x"05",  x"3E",  x"DD",  x"CB",  x"04",  x"1E",  x"10",  x"F6", -- 05C0
         x"DD",  x"34",  x"FF",  x"DD",  x"7E",  x"FF",  x"D6",  x"04", -- 05C8
         x"38",  x"CF",  x"33",  x"DD",  x"E1",  x"C9",  x"ED",  x"4B", -- 05D0
         x"00",  x"B0",  x"06",  x"00",  x"69",  x"60",  x"29",  x"29", -- 05D8
         x"09",  x"29",  x"29",  x"29",  x"11",  x"00",  x"EC",  x"19", -- 05E0
         x"06",  x"28",  x"36",  x"20",  x"23",  x"10",  x"FB",  x"C9", -- 05E8
         x"01",  x"07",  x"00",  x"11",  x"00",  x"EC",  x"21",  x"FE", -- 05F0
         x"05",  x"ED",  x"B0",  x"C3",  x"00",  x"EC",  x"3E",  x"05", -- 05F8
         x"D3",  x"02",  x"C3",  x"00",  x"F0",  x"C9",  x"CD",  x"4B", -- 0600
         x"04",  x"3E",  x"05",  x"D3",  x"02",  x"31",  x"00",  x"02", -- 0608
         x"C3",  x"89",  x"F0",  x"C9",  x"3E",  x"05",  x"D3",  x"02", -- 0610
         x"C1",  x"D1",  x"ED",  x"53",  x"D7",  x"03",  x"21",  x"BD", -- 0618
         x"C0",  x"11",  x"00",  x"03",  x"01",  x"67",  x"00",  x"ED", -- 0620
         x"B0",  x"EB",  x"F9",  x"AF",  x"32",  x"AB",  x"03",  x"32", -- 0628
         x"00",  x"04",  x"2A",  x"36",  x"00",  x"11",  x"00",  x"FF", -- 0630
         x"22",  x"B0",  x"03",  x"19",  x"22",  x"56",  x"03",  x"3E", -- 0638
         x"AF",  x"32",  x"FC",  x"03",  x"CD",  x"4F",  x"C6",  x"23", -- 0640
         x"EB",  x"CD",  x"93",  x"C4",  x"CD",  x"69",  x"C6",  x"C3", -- 0648
         x"54",  x"C8",  x"C9",  x"C1",  x"D1",  x"ED",  x"53",  x"D7", -- 0650
         x"03",  x"21",  x"BD",  x"C0",  x"11",  x"00",  x"03",  x"01", -- 0658
         x"67",  x"00",  x"ED",  x"B0",  x"EB",  x"F9",  x"21",  x"C0", -- 0660
         x"01",  x"22",  x"56",  x"03",  x"CD",  x"69",  x"C6",  x"32", -- 0668
         x"AB",  x"03",  x"32",  x"00",  x"04",  x"2A",  x"36",  x"00", -- 0670
         x"11",  x"00",  x"FF",  x"22",  x"B0",  x"03",  x"19",  x"22", -- 0678
         x"56",  x"03",  x"AF",  x"32",  x"5E",  x"03",  x"CD",  x"4F", -- 0680
         x"C6",  x"3E",  x"AF",  x"32",  x"FC",  x"03",  x"31",  x"67", -- 0688
         x"03",  x"CD",  x"69",  x"C6",  x"CD",  x"4F",  x"C6",  x"C3", -- 0690
         x"54",  x"C8",  x"C9",  x"DD",  x"E5",  x"DD",  x"21",  x"00", -- 0698
         x"00",  x"DD",  x"39",  x"DD",  x"6E",  x"04",  x"DD",  x"66", -- 06A0
         x"05",  x"DD",  x"4E",  x"08",  x"DD",  x"46",  x"09",  x"51", -- 06A8
         x"58",  x"0B",  x"7B",  x"B2",  x"28",  x"07",  x"DD",  x"7E", -- 06B0
         x"06",  x"77",  x"23",  x"18",  x"F2",  x"DD",  x"6E",  x"04", -- 06B8
         x"DD",  x"66",  x"05",  x"DD",  x"E1",  x"C9",  x"00",  x"01", -- 06C0
         x"01",  x"00",  x"78",  x"B1",  x"28",  x"08",  x"11",  x"00", -- 06C8
         x"B0",  x"21",  x"C6",  x"06",  x"ED",  x"B0",  x"C9",  x"00", -- 06D0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 06D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 06E0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 06E8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 06F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 06F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0700
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0708
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0710
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0718
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0720
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0728
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0730
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0738
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0740
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0748
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0750
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0758
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0760
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0768
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0770
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0778
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0780
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0788
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0790
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0798
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 07A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 07A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 07B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 07B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 07C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 07C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 07D0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 07D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 07E0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 07E8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 07F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00"  -- 07F8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
