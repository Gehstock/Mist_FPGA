library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity time_pilot_sprite_grphx is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of time_pilot_sprite_grphx is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"91",X"23",
		X"00",X"00",X"00",X"00",X"40",X"10",X"88",X"5C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"23",X"51",X"00",X"90",X"00",X"00",X"00",X"00",
		X"4C",X"E8",X"40",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"80",X"11",X"A3",
		X"00",X"00",X"00",X"00",X"80",X"10",X"88",X"4C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"23",X"51",X"80",X"10",X"00",X"00",X"00",X"00",
		X"4C",X"A8",X"00",X"20",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"10",X"00",X"00",X"40",X"00",X"20",X"00",X"11",X"23",
		X"00",X"00",X"00",X"40",X"00",X"20",X"88",X"4C",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"40",
		X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"23",X"11",X"80",X"00",X"10",X"00",X"00",X"00",
		X"4C",X"A8",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"40",X"11",X"23",
		X"00",X"00",X"00",X"80",X"00",X"20",X"88",X"5C",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"23",X"51",X"00",X"80",X"10",X"40",X"00",X"00",
		X"4C",X"A8",X"80",X"20",X"00",X"20",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"66",X"57",X"23",X"11",X"11",X"00",X"00",X"11",X"11",X"23",X"EF",X"2F",X"0F",X"8F",
		X"88",X"4C",X"4C",X"4C",X"2E",X"3F",X"0F",X"0F",X"00",X"00",X"00",X"33",X"EF",X"1F",X"2E",X"4C",
		X"00",X"10",X"70",X"10",X"00",X"00",X"11",X"11",X"CF",X"E3",X"C7",X"C7",X"8F",X"9F",X"2E",X"4C",
		X"0F",X"1F",X"1F",X"0F",X"8F",X"67",X"11",X"00",X"C8",X"E0",X"C0",X"88",X"4C",X"3F",X"9F",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"12",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"13",X"11",X"20",X"22",X"00",X"00",X"00",X"11",
		X"48",X"4C",X"00",X"80",X"80",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"84",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"12",X"10",X"11",X"00",X"20",X"22",X"00",X"22",
		X"0C",X"08",X"00",X"40",X"44",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"84",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"00",X"10",X"11",X"00",X"11",X"22",
		X"84",X"88",X"00",X"00",X"00",X"00",X"40",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"12",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"23",X"00",X"00",X"00",X"10",X"00",X"11",
		X"C0",X"80",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"30",X"40",X"40",X"30",X"00",X"00",X"30",X"00",X"E0",X"10",X"10",X"E0",X"00",X"00",X"E0",
		X"00",X"00",X"02",X"02",X"03",X"00",X"02",X"03",X"00",X"00",X"0E",X"0A",X"0A",X"00",X"00",X"0E",
		X"40",X"40",X"30",X"00",X"00",X"70",X"20",X"00",X"10",X"10",X"E0",X"00",X"10",X"F0",X"10",X"00",
		X"02",X"00",X"03",X"02",X"03",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"0E",X"00",X"00",X"00",
		X"00",X"30",X"40",X"40",X"30",X"00",X"00",X"30",X"00",X"E0",X"10",X"10",X"E0",X"00",X"00",X"E0",
		X"00",X"00",X"02",X"02",X"03",X"00",X"02",X"03",X"00",X"00",X"0E",X"0A",X"0A",X"00",X"00",X"0E",
		X"40",X"40",X"30",X"00",X"40",X"40",X"70",X"00",X"10",X"10",X"E0",X"00",X"F0",X"90",X"90",X"00",
		X"02",X"00",X"03",X"02",X"03",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"0E",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"C9",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"84",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"83",X"32",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"BA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"74",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C8",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"81",X"00",X"00",X"00",X"00",X"00",X"00",
		X"84",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"83",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C8",X"00",X"00",X"00",X"00",X"00",X"00",X"32",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"84",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"32",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"84",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"74",X"F8",X"F8",
		X"00",X"00",X"00",X"00",X"CC",X"E2",X"F1",X"F1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"F8",X"74",X"33",X"00",X"00",X"00",X"00",
		X"F1",X"F1",X"E2",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"77",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"CC",X"EE",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"77",X"33",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"EE",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"03",X"03",X"03",X"03",
		X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"07",X"07",X"07",X"07",X"07",
		X"80",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0C",X"4A",X"4B",X"69",X"E1",X"E1",X"E1",X"E1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"E1",X"E1",X"E1",X"C3",X"C3",X"C3",X"4B",X"4B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"7F",X"7F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"CF",X"CF",X"0F",X"0F",X"0F",X"08",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",
		X"0F",X"0F",X"3F",X"7F",X"7F",X"7F",X"3F",X"0F",X"0F",X"0F",X"8F",X"CF",X"CF",X"CF",X"8F",X"0F",
		X"0F",X"0F",X"3C",X"78",X"78",X"78",X"3C",X"0F",X"0E",X"0E",X"86",X"C2",X"C2",X"C2",X"86",X"0E",
		X"0F",X"0F",X"0F",X"0F",X"3C",X"3C",X"3C",X"3C",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"F0",X"F0",X"0E",X"0E",X"0E",X"0E",X"86",X"86",X"86",X"86",
		X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"86",X"86",X"86",X"86",X"86",X"86",X"86",X"86",
		X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"86",X"86",X"86",X"86",X"86",X"86",X"86",X"86",
		X"3C",X"1E",X"0F",X"0F",X"0F",X"0F",X"0F",X"03",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"86",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"08",
		X"03",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"7F",X"7F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"CF",X"CF",X"0F",X"0F",X"0F",X"08",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",
		X"0F",X"0F",X"3C",X"78",X"78",X"78",X"3C",X"0F",X"0F",X"0F",X"87",X"C3",X"C3",X"C3",X"87",X"0F",
		X"0F",X"0F",X"3F",X"7F",X"7F",X"7F",X"3F",X"0F",X"0E",X"0E",X"8E",X"CE",X"CE",X"CE",X"8E",X"0E",
		X"03",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"78",X"78",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"C3",X"C3",X"0F",X"0F",X"0F",X"08",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",
		X"0F",X"0F",X"3F",X"7F",X"7F",X"7F",X"3F",X"0F",X"0F",X"0F",X"8F",X"CF",X"CF",X"CF",X"8F",X"0F",
		X"0F",X"0F",X"3F",X"7F",X"7F",X"7F",X"3F",X"0F",X"0E",X"0E",X"8E",X"CE",X"CE",X"CE",X"8E",X"0E",
		X"00",X"00",X"00",X"00",X"03",X"16",X"BC",X"F8",X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"7F",
		X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",X"00",X"00",X"00",X"00",X"0C",X"86",X"C3",X"E1",
		X"E9",X"E9",X"E9",X"E9",X"E9",X"F8",X"F8",X"FF",X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",
		X"11",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",X"E9",X"E9",X"E9",X"E9",X"E9",X"F0",X"F0",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",
		X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",X"00",X"00",X"00",X"00",X"0F",X"E1",X"E1",X"EF",
		X"00",X"00",X"00",X"00",X"03",X"16",X"BC",X"F8",X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",
		X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",
		X"E9",X"E9",X"E9",X"E9",X"F8",X"FC",X"76",X"33",X"08",X"00",X"00",X"08",X"0F",X"F0",X"F0",X"FF",
		X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",
		X"00",X"00",X"8F",X"F8",X"F8",X"FF",X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",X"00",X"00",
		X"00",X"00",X"0F",X"F0",X"F0",X"FF",X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"8F",X"F8",X"F8",X"FF",X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",
		X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",
		X"00",X"00",X"0F",X"F0",X"F0",X"FF",X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",X"01",X"06",
		X"00",X"00",X"0F",X"F0",X"F0",X"F8",X"F1",X"F7",X"00",X"00",X"0F",X"E1",X"E1",X"F7",X"CC",X"00",
		X"01",X"11",X"00",X"00",X"0F",X"F0",X"F0",X"FF",X"78",X"F8",X"76",X"11",X"0F",X"F0",X"F0",X"FF",
		X"84",X"84",X"87",X"E1",X"78",X"F0",X"F0",X"FF",X"00",X"00",X"00",X"0C",X"87",X"E1",X"E1",X"FF",
		X"00",X"00",X"00",X"00",X"8F",X"E9",X"E9",X"E9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"23",
		X"E9",X"E9",X"E9",X"E9",X"E9",X"F8",X"F8",X"FF",X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",
		X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",X"32",X"32",X"32",X"32",X"3E",X"F0",X"F0",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"8F",X"E9",X"E9",X"E9",
		X"84",X"84",X"84",X"84",X"87",X"F0",X"F0",X"FF",X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",
		X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",X"E9",X"E9",X"E9",X"E9",X"E9",X"E1",X"E1",X"FF",
		X"00",X"00",X"00",X"00",X"03",X"16",X"3C",X"78",X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",
		X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",X"00",X"00",X"00",X"00",X"0C",X"86",X"C3",X"F1",
		X"79",X"69",X"69",X"69",X"69",X"78",X"78",X"FF",X"88",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",
		X"11",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",X"F8",X"F8",X"F9",X"E9",X"E9",X"F0",X"F0",X"FF",
		X"00",X"00",X"00",X"00",X"03",X"16",X"3C",X"79",X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",
		X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",X"00",X"00",X"00",X"00",X"0F",X"E1",X"E1",X"FF",
		X"F3",X"E6",X"CC",X"08",X"0F",X"F0",X"F0",X"FF",X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",
		X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",X"00",X"00",X"00",X"00",X"0F",X"E1",X"E1",X"FF",
		X"00",X"00",X"00",X"00",X"03",X"16",X"BC",X"F8",X"00",X"00",X"00",X"00",X"0C",X"84",X"84",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"32",
		X"E9",X"E9",X"E9",X"E9",X"F8",X"FC",X"76",X"33",X"08",X"00",X"00",X"08",X"0F",X"F0",X"F0",X"FF",
		X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",X"32",X"32",X"32",X"16",X"3C",X"F0",X"F1",X"FF",
		X"00",X"00",X"00",X"00",X"0F",X"78",X"F0",X"F3",X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",
		X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",X"00",X"00",X"00",X"00",X"0C",X"86",X"C3",X"E1",
		X"E6",X"C4",X"C4",X"C4",X"C4",X"CC",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"00",X"00",X"01",X"23",X"32",X"32",X"33",X"E9",X"E9",X"E9",X"69",X"E1",X"C3",X"86",X"CC",
		X"00",X"00",X"00",X"00",X"8F",X"F8",X"F8",X"FF",X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",
		X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",
		X"00",X"00",X"00",X"00",X"8F",X"F8",X"F8",X"FF",X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",
		X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",
		X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",
		X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",X"00",X"00",X"00",X"00",X"0C",X"86",X"C3",X"E1",
		X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",
		X"11",X"00",X"00",X"01",X"0F",X"F0",X"F0",X"FF",X"E9",X"E9",X"E9",X"E9",X"E1",X"F3",X"E6",X"CC",
		X"00",X"00",X"00",X"00",X"03",X"16",X"BC",X"F8",X"00",X"00",X"00",X"00",X"0C",X"84",X"84",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E9",X"E9",X"E9",X"E9",X"F8",X"FC",X"76",X"33",X"08",X"00",X"00",X"08",X"0F",X"F0",X"F0",X"FF",
		X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",
		X"00",X"00",X"00",X"00",X"8F",X"F8",X"F8",X"E9",X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",
		X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",X"00",X"00",X"00",X"00",X"0C",X"86",X"C3",X"E1",
		X"E9",X"FF",X"00",X"00",X"0F",X"F0",X"F0",X"FF",X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"FF",
		X"11",X"00",X"00",X"11",X"0F",X"F0",X"F0",X"FF",X"E9",X"E9",X"E9",X"E9",X"E1",X"F3",X"E6",X"CC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"90",X"90",X"B0",X"A1",X"93",X"57",X"13",
		X"88",X"CC",X"5D",X"1D",X"3F",X"1D",X"9D",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"13",X"01",X"01",X"11",X"11",X"01",X"23",X"33",
		X"5D",X"5D",X"0C",X"08",X"08",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"90",X"90",X"B0",X"A1",X"57",X"13",
		X"00",X"88",X"DD",X"DD",X"7F",X"1D",X"1D",X"BF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"01",X"01",X"11",X"11",X"23",X"33",X"00",
		X"DD",X"1D",X"08",X"08",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"90",X"90",X"B0",X"47",X"13",
		X"00",X"00",X"88",X"DD",X"DD",X"7F",X"1D",X"BF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"01",X"01",X"11",X"23",X"33",X"00",X"00",
		X"9D",X"DD",X"08",X"08",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"90",X"B0",X"B0",X"56",X"03",
		X"00",X"00",X"88",X"CC",X"DD",X"FF",X"5D",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"01",X"01",X"33",X"00",X"00",X"00",X"00",
		X"9D",X"CC",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"90",X"B0",X"74",X"30",
		X"00",X"00",X"00",X"1D",X"6E",X"4E",X"CE",X"4E",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AE",X"1D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"43",X"E1",X"70",X"70",X"21",X"43",
		X"00",X"10",X"C3",X"2D",X"7A",X"7C",X"F8",X"E1",X"00",X"80",X"C0",X"48",X"68",X"2C",X"48",X"48",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"43",X"2D",X"F0",X"F0",X"70",X"21",X"00",X"00",
		X"E9",X"6D",X"5F",X"3C",X"5A",X"69",X"68",X"40",X"C8",X"E8",X"E0",X"C0",X"C0",X"C0",X"00",X"00",
		X"00",X"10",X"10",X"30",X"03",X"61",X"70",X"70",X"40",X"E0",X"E1",X"C3",X"C3",X"3E",X"B6",X"1F",
		X"40",X"F0",X"F0",X"87",X"3F",X"F1",X"E1",X"E1",X"00",X"00",X"80",X"68",X"2C",X"4E",X"F8",X"F8",
		X"70",X"21",X"00",X"00",X"00",X"00",X"00",X"00",X"4B",X"C3",X"E1",X"F0",X"F0",X"70",X"00",X"00",
		X"E9",X"F0",X"69",X"69",X"69",X"00",X"00",X"00",X"48",X"2C",X"4A",X"E0",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"01",X"10",X"30",X"87",X"E1",
		X"00",X"30",X"07",X"F3",X"F0",X"E1",X"E9",X"E5",X"00",X"00",X"08",X"68",X"8E",X"48",X"C0",X"68",
		X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"E1",X"C3",X"D2",X"30",X"10",X"10",X"00",X"00",
		X"3F",X"87",X"C3",X"C3",X"96",X"B4",X"78",X"00",X"68",X"68",X"E8",X"E8",X"C0",X"C0",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"30",X"21",X"13",X"57",X"93",
		X"88",X"CC",X"5D",X"1D",X"3F",X"1D",X"9D",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"93",X"81",X"81",X"91",X"91",X"01",X"23",X"33",
		X"5D",X"5D",X"0C",X"08",X"08",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"30",X"21",X"57",X"93",
		X"00",X"88",X"DD",X"DD",X"7F",X"1D",X"1D",X"BF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"91",X"81",X"81",X"91",X"91",X"23",X"33",X"00",
		X"DD",X"1D",X"08",X"08",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"30",X"47",X"93",
		X"00",X"00",X"88",X"DD",X"DD",X"7F",X"1D",X"BF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"91",X"81",X"81",X"91",X"A3",X"33",X"00",X"00",
		X"9D",X"DD",X"08",X"08",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"30",X"56",X"83",
		X"00",X"00",X"88",X"CC",X"DD",X"FF",X"5D",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"91",X"81",X"81",X"B3",X"80",X"00",X"00",X"00",
		X"9D",X"CC",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"74",X"B0",
		X"00",X"00",X"00",X"1D",X"6E",X"4E",X"CE",X"4E",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"80",X"80",X"80",X"80",X"00",X"00",X"00",
		X"AE",X"1D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"88",X"FF",X"00",X"FF",X"88",X"FF",X"00",
		X"EE",X"22",X"EE",X"00",X"EE",X"22",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"88",X"FF",X"00",X"FF",X"99",X"99",X"00",
		X"EE",X"22",X"EE",X"00",X"EE",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"88",X"FF",X"00",X"FF",X"88",X"FF",X"00",
		X"EE",X"22",X"EE",X"00",X"EE",X"22",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"88",X"FF",X"00",X"00",X"FF",X"00",X"FF",
		X"EE",X"22",X"EE",X"00",X"88",X"EE",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"88",X"FF",X"00",X"FF",X"88",X"FF",X"00",
		X"EE",X"22",X"EE",X"00",X"EE",X"22",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"88",X"FF",X"00",X"99",X"99",X"FF",X"00",
		X"EE",X"22",X"EE",X"00",X"EE",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"53",X"43",X"61",X"21",X"30",X"10",X"10",X"10",
		X"DE",X"9E",X"BC",X"2C",X"68",X"48",X"48",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"30",X"21",X"61",X"43",X"53",
		X"C0",X"48",X"48",X"68",X"2C",X"BC",X"9E",X"DE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B7",X"D3",X"43",X"61",X"21",X"30",X"10",X"10",
		X"EF",X"DE",X"9E",X"BC",X"2C",X"68",X"48",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"30",X"21",X"61",X"43",X"D3",X"B7",
		X"C0",X"48",X"68",X"2C",X"BC",X"9E",X"DE",X"EF",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"30",X"E1",X"10",X"00",X"00",X"10",X"30",X"40",X"3F",X"7F",X"B7",X"97",X"C3",X"E1",X"21",X"21",
		X"EF",X"8F",X"3C",X"68",X"2C",X"3C",X"F0",X"80",X"48",X"F0",X"80",X"00",X"00",X"00",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",
		X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"00",X"00",X"90",X"61",X"30",X"10",X"10",X"F0",X"87",X"97",X"D3",X"3F",X"1F",X"D3",X"97",
		X"48",X"48",X"78",X"0F",X"DE",X"BC",X"9E",X"DE",X"10",X"20",X"C0",X"80",X"80",X"00",X"00",X"80",
		X"F0",X"21",X"10",X"00",X"00",X"10",X"30",X"30",X"7F",X"3F",X"97",X"C3",X"D3",X"87",X"0F",X"C3",
		X"8F",X"EF",X"9E",X"BC",X"BC",X"1E",X"87",X"F0",X"80",X"48",X"F0",X"00",X"00",X"80",X"80",X"C0",
		X"60",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"61",X"30",X"10",X"10",X"10",X"10",X"10",X"00",
		X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"40",X"20",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"20",X"30",X"21",X"21",X"61",
		X"00",X"00",X"00",X"00",X"00",X"80",X"F0",X"0F",X"00",X"00",X"00",X"20",X"40",X"C0",X"80",X"80",
		X"00",X"F0",X"61",X"10",X"10",X"00",X"00",X"10",X"43",X"D3",X"1F",X"7F",X"97",X"C3",X"97",X"B7",
		X"9E",X"BC",X"9E",X"CF",X"EF",X"CF",X"9E",X"3C",X"80",X"00",X"80",X"78",X"C0",X"80",X"80",X"80",
		X"00",X"00",X"00",X"20",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"33",X"B3",X"63",X"AD",
		X"00",X"00",X"00",X"22",X"44",X"7E",X"7D",X"7B",X"00",X"00",X"00",X"40",X"80",X"00",X"00",X"88",
		X"33",X"00",X"00",X"00",X"10",X"20",X"00",X"00",X"CF",X"65",X"63",X"B3",X"11",X"00",X"00",X"00",
		X"0E",X"7B",X"7D",X"7E",X"22",X"88",X"00",X"00",X"44",X"00",X"88",X"00",X"80",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"11",X"00",X"00",X"00",X"22",X"11",X"91",X"63",X"65",
		X"00",X"00",X"00",X"00",X"10",X"20",X"C8",X"C4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"CF",X"65",X"63",X"91",X"11",X"00",X"00",X"00",
		X"6E",X"95",X"C8",X"A8",X"10",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"91",X"51",X"75",
		X"00",X"00",X"00",X"00",X"00",X"20",X"C8",X"D5",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"75",X"51",X"80",X"00",X"00",X"00",X"00",
		X"EE",X"C4",X"C8",X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"11",X"51",X"75",
		X"00",X"00",X"00",X"00",X"88",X"00",X"C8",X"C4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"75",X"73",X"22",X"00",X"00",X"00",X"00",
		X"EE",X"A2",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"80",X"60",X"30",X"31",
		X"00",X"00",X"00",X"00",X"A0",X"C0",X"C8",X"E8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"50",X"40",X"80",X"10",X"00",X"00",X"00",
		X"FC",X"C4",X"C0",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"10",X"00",X"00",X"00",X"40",X"20",X"20",X"60",X"F1",X"33",
		X"00",X"00",X"00",X"20",X"C0",X"90",X"A0",X"E8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"73",X"F0",X"60",X"20",X"20",X"40",X"00",X"00",
		X"FC",X"88",X"C0",X"40",X"20",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"20",X"10",X"00",X"40",X"30",X"00",X"00",X"10",X"20",X"B0",X"F2",X"63",X"C7",
		X"00",X"00",X"00",X"10",X"20",X"60",X"48",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"80",
		X"00",X"10",X"20",X"00",X"00",X"00",X"00",X"00",X"E7",X"F1",X"50",X"D0",X"40",X"20",X"00",X"00",
		X"6C",X"F8",X"C0",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"10",X"00",X"60",X"B0",X"00",X"00",X"00",X"00",X"A0",X"E0",X"D0",X"F2",X"E7",
		X"00",X"40",X"80",X"80",X"C0",X"F4",X"EC",X"3E",X"00",X"00",X"00",X"00",X"80",X"00",X"40",X"00",
		X"10",X"30",X"40",X"10",X"00",X"00",X"00",X"00",X"C7",X"E3",X"F2",X"70",X"50",X"90",X"00",X"00",
		X"6C",X"F8",X"E8",X"A0",X"20",X"90",X"80",X"40",X"00",X"A0",X"C0",X"00",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"61",X"61",X"25",X"16",X"16",X"05",X"05",X"05",
		X"48",X"0C",X"84",X"84",X"EE",X"0C",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"12",X"12",X"10",X"00",X"00",X"00",
		X"84",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"12",X"03",X"01",X"00",X"00",X"00",X"00",X"E0",X"D2",X"5A",X"1E",X"2D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"07",X"07",X"25",X"34",X"70",X"61",
		X"08",X"0C",X"0C",X"04",X"0C",X"0C",X"48",X"48",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"61",X"61",X"25",X"16",X"77",X"05",X"05",X"05",
		X"48",X"0C",X"84",X"84",X"84",X"0C",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"12",X"12",X"10",X"00",X"00",X"00",
		X"84",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"12",X"03",X"01",X"00",X"00",X"00",X"00",X"E0",X"D2",X"5A",X"1E",X"2D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"07",X"07",X"25",X"34",X"70",X"61",
		X"08",X"0C",X"0C",X"04",X"0C",X"0C",X"48",X"48",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"71",X"71",X"25",X"16",X"16",X"05",X"05",X"05",
		X"48",X"0C",X"84",X"84",X"EE",X"0C",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"12",X"12",X"10",X"00",X"00",X"00",
		X"84",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"12",X"03",X"01",X"00",X"00",X"00",X"00",X"E0",X"D2",X"5A",X"1E",X"2D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"07",X"07",X"67",X"76",X"FB",X"77",
		X"08",X"0C",X"0C",X"04",X"8C",X"8C",X"C8",X"48",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"71",X"71",X"25",X"16",X"77",X"05",X"05",X"05",
		X"48",X"0C",X"84",X"84",X"84",X"0C",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"12",X"12",X"10",X"00",X"00",X"00",
		X"84",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"12",X"03",X"01",X"00",X"00",X"00",X"00",X"E0",X"D2",X"5A",X"1E",X"2D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"07",X"07",X"07",X"47",X"67",X"BF",X"FF",X"73",
		X"08",X"0C",X"0C",X"44",X"CC",X"8C",X"C8",X"48",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"71",X"71",X"25",X"16",X"16",X"05",X"05",X"05",
		X"48",X"0C",X"84",X"84",X"EE",X"0C",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"12",X"12",X"10",X"00",X"00",X"00",
		X"84",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"12",X"03",X"01",X"00",X"00",X"00",X"00",X"E0",X"D2",X"5A",X"1E",X"2D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"07",X"07",X"17",X"57",X"67",X"BF",X"FF",X"73",
		X"08",X"0C",X"0C",X"44",X"4C",X"8C",X"C8",X"48",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"71",X"71",X"25",X"16",X"77",X"05",X"05",X"05",
		X"48",X"0C",X"84",X"84",X"84",X"0C",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"12",X"12",X"10",X"00",X"00",X"00",
		X"84",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"12",X"03",X"01",X"00",X"00",X"00",X"00",X"E0",X"D2",X"5A",X"1E",X"2D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DF",X"AF",X"67",X"67",X"BF",X"77",X"73",X"73",
		X"88",X"AE",X"AE",X"44",X"AE",X"EE",X"C8",X"48",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"71",X"71",X"25",X"16",X"16",X"05",X"05",X"05",
		X"48",X"0C",X"84",X"84",X"EE",X"0C",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"12",X"12",X"10",X"00",X"00",X"00",
		X"84",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"12",X"03",X"01",X"00",X"00",X"00",X"00",X"E0",X"D2",X"5A",X"1E",X"2D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9F",X"AF",X"77",X"67",X"BF",X"77",X"73",X"73",
		X"CC",X"AE",X"AE",X"44",X"9D",X"EE",X"C8",X"48",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"71",X"71",X"25",X"16",X"77",X"05",X"05",X"05",
		X"48",X"0C",X"84",X"84",X"84",X"0C",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"12",X"12",X"10",X"00",X"00",X"00",
		X"84",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"12",X"03",X"01",X"11",X"00",X"00",X"00",X"E0",X"F2",X"7A",X"9F",X"7D",
		X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"47",X"EF",X"77",X"37",X"37",X"76",X"73",X"71",
		X"88",X"8C",X"8C",X"44",X"8C",X"AE",X"EE",X"C8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"12",X"12",X"12",X"12",X"12",X"02",X"02",X"77",
		X"2C",X"C2",X"C2",X"C2",X"C0",X"E0",X"A4",X"A4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"02",X"02",X"00",X"01",X"00",X"00",
		X"2C",X"2C",X"68",X"68",X"68",X"E2",X"E2",X"C4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"30",X"03",X"01",X"00",X"00",X"00",X"00",X"E0",X"B4",X"B4",X"5A",X"4B",X"07",X"07",X"07",
		X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"12",X"12",X"12",X"12",X"30",X"23",X"27",X"32",
		X"80",X"C4",X"C6",X"C4",X"C0",X"C0",X"E0",X"68",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"12",X"12",X"12",X"12",X"12",X"02",X"02",X"03",
		X"2C",X"C2",X"C2",X"C2",X"C0",X"E0",X"E0",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"02",X"02",X"00",X"01",X"00",X"00",
		X"2C",X"2C",X"68",X"68",X"68",X"E2",X"E2",X"C4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"30",X"03",X"01",X"00",X"00",X"00",X"00",X"E0",X"B4",X"B4",X"5A",X"4B",X"07",X"07",X"07",
		X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"12",X"12",X"12",X"12",X"30",X"23",X"27",X"32",
		X"80",X"C4",X"C6",X"C4",X"C0",X"C0",X"E0",X"68",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"12",X"12",X"12",X"12",X"12",X"02",X"02",X"77",
		X"AC",X"8E",X"86",X"82",X"C0",X"E0",X"A4",X"A4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"02",X"02",X"00",X"01",X"00",X"00",
		X"2C",X"2C",X"68",X"68",X"68",X"E2",X"E2",X"C4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"30",X"03",X"01",X"00",X"00",X"00",X"00",X"E0",X"B4",X"B4",X"5A",X"4B",X"07",X"07",X"8F",
		X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9A",X"9B",X"56",X"56",X"BA",X"77",X"37",X"33",
		X"80",X"C4",X"CE",X"CC",X"C8",X"C4",X"E8",X"E8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"12",X"12",X"12",X"12",X"12",X"02",X"02",X"03",
		X"AC",X"8E",X"86",X"82",X"C0",X"E0",X"A4",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"02",X"02",X"00",X"01",X"00",X"00",
		X"2C",X"2C",X"68",X"68",X"68",X"E2",X"E2",X"C4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"30",X"03",X"01",X"00",X"00",X"00",X"00",X"E0",X"B4",X"B4",X"5A",X"4B",X"07",X"07",X"07",
		X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"13",X"13",X"57",X"32",X"B9",X"77",X"77",X"33",
		X"80",X"CC",X"C6",X"CC",X"C8",X"C8",X"E0",X"E8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"13",X"12",X"12",X"12",X"02",X"02",X"77",
		X"2C",X"86",X"86",X"82",X"C0",X"E0",X"A4",X"A4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"02",X"02",X"00",X"01",X"00",X"00",
		X"2C",X"2C",X"68",X"68",X"68",X"E2",X"E2",X"C4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"30",X"03",X"01",X"00",X"22",X"22",X"33",X"E0",X"B4",X"B4",X"5E",X"4F",X"CF",X"CF",X"67",
		X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"FE",X"FE",X"76",X"BB",X"FF",X"67",X"33",X"33",
		X"80",X"C4",X"CE",X"C4",X"C0",X"C0",X"E0",X"E8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"13",X"12",X"12",X"12",X"02",X"02",X"03",
		X"2C",X"86",X"86",X"82",X"C0",X"E0",X"A4",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"02",X"02",X"00",X"01",X"00",X"00",
		X"2C",X"2C",X"68",X"68",X"68",X"E2",X"E2",X"C4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"30",X"03",X"01",X"00",X"00",X"00",X"00",X"E0",X"B4",X"B4",X"5A",X"4B",X"47",X"47",X"23",
		X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"BA",X"BB",X"76",X"76",X"67",X"33",X"33",
		X"C4",X"CC",X"C6",X"C4",X"C8",X"C8",X"E8",X"E8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"13",X"12",X"12",X"12",X"02",X"02",X"77",
		X"2C",X"86",X"86",X"82",X"C0",X"E0",X"A4",X"A4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"02",X"02",X"00",X"01",X"00",X"00",
		X"2C",X"2C",X"68",X"68",X"68",X"E2",X"E2",X"C4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"31",X"13",X"11",X"00",X"00",X"00",X"11",X"E0",X"B4",X"F4",X"5E",X"EB",X"FF",X"67",X"23",
		X"00",X"00",X"22",X"44",X"44",X"4C",X"4C",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"76",X"FF",X"77",X"57",X"33",X"BB",X"77",X"33",
		X"88",X"C4",X"C6",X"CC",X"C0",X"CC",X"E0",X"E8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"13",X"12",X"12",X"12",X"02",X"02",X"03",
		X"2C",X"86",X"86",X"82",X"C0",X"E0",X"A4",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"02",X"02",X"00",X"01",X"00",X"00",
		X"2C",X"2C",X"68",X"68",X"68",X"E2",X"E2",X"C4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"30",X"03",X"23",X"22",X"11",X"11",X"11",X"E0",X"B4",X"F4",X"5E",X"6F",X"27",X"27",X"9F",
		X"00",X"00",X"00",X"00",X"00",X"4C",X"4C",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DF",X"76",X"BB",X"BA",X"77",X"77",X"27",X"33",
		X"C4",X"C4",X"C6",X"C4",X"C8",X"C8",X"EC",X"E8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"10",X"10",X"10",X"01",X"01",X"03",X"07",X"1E",X"3C",
		X"43",X"C3",X"C3",X"43",X"C3",X"C3",X"42",X"C3",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",
		X"11",X"11",X"11",X"11",X"11",X"11",X"00",X"00",X"3C",X"37",X"33",X"11",X"10",X"00",X"00",X"00",
		X"C2",X"E0",X"A4",X"86",X"86",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"10",X"00",X"00",X"00",X"13",X"17",X"3D",X"2D",X"0F",
		X"00",X"00",X"00",X"80",X"C0",X"84",X"86",X"86",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"00",X"0F",X"16",X"12",X"10",X"10",X"10",X"10",X"10",
		X"87",X"87",X"86",X"C3",X"C3",X"43",X"C3",X"C3",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"10",X"10",X"10",X"01",X"01",X"03",X"07",X"1E",X"3C",
		X"43",X"C3",X"C3",X"43",X"C3",X"C3",X"42",X"C3",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",
		X"11",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"3C",X"37",X"33",X"11",X"10",X"00",X"00",X"00",
		X"C2",X"E0",X"A4",X"86",X"86",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"10",X"00",X"00",X"00",X"13",X"17",X"3D",X"2D",X"0F",
		X"00",X"00",X"00",X"80",X"C0",X"84",X"86",X"86",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"0F",X"16",X"12",X"10",X"10",X"10",X"10",X"10",
		X"87",X"87",X"86",X"C3",X"C3",X"43",X"C3",X"C3",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"10",X"10",X"10",X"01",X"01",X"03",X"07",X"1E",X"3C",
		X"CB",X"CB",X"C3",X"43",X"C3",X"C3",X"42",X"C3",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",
		X"11",X"11",X"11",X"11",X"11",X"11",X"00",X"00",X"3C",X"37",X"33",X"11",X"10",X"00",X"00",X"00",
		X"C2",X"E0",X"A4",X"86",X"86",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"10",X"00",X"00",X"00",X"13",X"17",X"3D",X"2D",X"0F",
		X"00",X"00",X"00",X"80",X"C0",X"84",X"86",X"86",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"00",X"5F",X"76",X"32",X"BB",X"77",X"11",X"77",X"11",
		X"C7",X"DF",X"FF",X"CF",X"E3",X"CF",X"CB",X"CF",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"10",X"11",X"10",X"01",X"01",X"03",X"07",X"1E",X"3C",
		X"CB",X"CB",X"C3",X"43",X"C3",X"C3",X"42",X"C3",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",
		X"11",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"3C",X"37",X"33",X"11",X"10",X"00",X"00",X"00",
		X"C2",X"E0",X"A4",X"86",X"86",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"10",X"00",X"00",X"00",X"13",X"57",X"7D",X"7F",X"2F",
		X"00",X"00",X"00",X"80",X"C0",X"C4",X"E6",X"CE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"AF",X"76",X"FF",X"FF",X"32",X"55",X"77",X"11",
		X"CF",X"8F",X"E6",X"C7",X"CB",X"CB",X"CF",X"CB",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"10",X"10",X"10",X"01",X"01",X"03",X"07",X"1E",X"3C",
		X"CB",X"CB",X"C3",X"43",X"C3",X"C3",X"42",X"C3",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",
		X"11",X"11",X"11",X"11",X"11",X"11",X"00",X"00",X"3C",X"37",X"33",X"11",X"10",X"00",X"00",X"00",
		X"C2",X"E0",X"A4",X"86",X"86",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"33",X"11",X"10",X"00",X"11",X"55",X"77",X"37",X"BF",X"BF",X"AF",
		X"00",X"00",X"22",X"A2",X"EA",X"DD",X"F7",X"E6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"00",X"EF",X"37",X"FF",X"77",X"33",X"77",X"77",X"11",
		X"CF",X"FF",X"CE",X"CB",X"EB",X"EF",X"CF",X"CB",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"10",X"10",X"10",X"01",X"01",X"03",X"07",X"1E",X"3C",
		X"CB",X"CB",X"C3",X"43",X"C3",X"C3",X"42",X"C3",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",
		X"11",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"3C",X"37",X"33",X"11",X"10",X"00",X"00",X"00",
		X"C2",X"E0",X"A4",X"86",X"86",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"BB",X"77",X"77",X"33",X"11",X"11",X"32",X"00",X"AA",X"66",X"BB",X"DF",X"FF",X"6F",X"AF",
		X"22",X"AA",X"FF",X"EE",X"EA",X"AE",X"BF",X"AE",X"00",X"88",X"00",X"00",X"00",X"88",X"00",X"00",
		X"11",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"AF",X"FF",X"77",X"DD",X"33",X"99",X"77",X"11",
		X"EF",X"DF",X"EE",X"CF",X"CB",X"EF",X"CF",X"CB",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"69",X"69",X"69",X"69",X"2D",X"2D",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"9E",X"9E",X"8F",X"07",X"07",X"07",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"07",X"03",X"03",X"03",
		X"02",X"86",X"86",X"86",X"86",X"A4",X"2C",X"2C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"2D",X"2D",X"69",X"69",X"69",X"69",X"69",X"69",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"6D",X"6D",X"69",X"69",X"2D",X"2D",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"9E",X"9E",X"8F",X"07",X"07",X"07",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"07",X"03",X"03",X"03",
		X"02",X"86",X"86",X"86",X"86",X"A4",X"2C",X"2C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"23",X"33",X"11",X"55",X"33",X"01",X"33",X"01",
		X"AF",X"6F",X"7F",X"EF",X"F9",X"EF",X"ED",X"EF",X"00",X"88",X"88",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"ED",X"6D",X"69",X"69",X"2D",X"2D",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"9E",X"9E",X"8F",X"07",X"07",X"07",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"27",X"AB",X"77",X"9B",
		X"02",X"86",X"86",X"86",X"86",X"AE",X"BF",X"6E",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"BB",X"77",X"77",X"11",X"23",X"33",X"01",
		X"6F",X"6D",X"FB",X"EB",X"6D",X"FD",X"EF",X"ED",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"6D",X"6D",X"69",X"69",X"2D",X"2D",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"9E",X"9E",X"8F",X"07",X"07",X"07",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"55",X"33",X"33",X"11",X"00",X"00",X"11",X"44",X"5F",X"3F",X"DF",X"EF",X"FF",X"33",X"57",
		X"13",X"D7",X"F7",X"F7",X"D7",X"FD",X"7D",X"7D",X"00",X"44",X"88",X"00",X"00",X"44",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"77",X"33",X"67",X"11",X"45",X"33",X"01",
		X"7F",X"EF",X"FF",X"EF",X"ED",X"FF",X"EF",X"ED",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EF",X"EF",X"EF",X"77",X"23",X"01",X"01",X"01",X"3F",X"BF",X"3F",X"3F",X"3F",X"BF",X"3F",X"7F",
		X"CF",X"CF",X"FF",X"FF",X"FF",X"CF",X"CF",X"CF",X"8F",X"8F",X"8F",X"8E",X"8E",X"8E",X"8C",X"8C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"33",X"11",X"11",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"CF",X"CF",X"FF",X"FF",X"47",X"77",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"30",X"FC",
		X"70",X"70",X"F0",X"F0",X"F0",X"C7",X"F7",X"FF",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"11",X"11",X"11",X"31",X"61",X"E1",X"E7",X"EF",X"FD",X"FD",X"FF",X"3F",X"3F",X"BF",X"3F",X"7F",
		X"CF",X"CF",X"CF",X"FF",X"FF",X"FF",X"CF",X"CF",X"CC",X"CC",X"AE",X"AE",X"AE",X"9F",X"9F",X"8F",
		X"EF",X"EF",X"EF",X"67",X"23",X"01",X"01",X"11",X"3F",X"BF",X"3F",X"7F",X"3F",X"BF",X"3F",X"3F",
		X"FF",X"FF",X"FF",X"CF",X"CF",X"CF",X"FF",X"FF",X"8F",X"8F",X"8F",X"8E",X"8E",X"8E",X"8C",X"8C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"33",X"11",X"11",X"00",X"00",X"00",X"00",
		X"CF",X"CF",X"FF",X"FF",X"CF",X"CF",X"77",X"47",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"30",X"FC",
		X"70",X"70",X"F0",X"F0",X"F0",X"F0",X"C7",X"C7",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"11",X"11",X"11",X"31",X"71",X"E1",X"E1",X"F7",X"FC",X"FD",X"FD",X"FF",X"3F",X"BF",X"3F",X"3F",
		X"CF",X"FF",X"FF",X"FF",X"CF",X"CF",X"CF",X"CF",X"C4",X"CC",X"EE",X"AE",X"AE",X"BF",X"9F",X"9F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"31",X"73",X"73",X"B7",X"3F",
		X"C0",X"40",X"E8",X"64",X"56",X"56",X"CF",X"47",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"37",X"37",X"33",X"11",X"11",X"00",X"00",
		X"47",X"47",X"CF",X"46",X"46",X"44",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"30",X"71",X"73",X"B7",X"3F",
		X"C0",X"C0",X"60",X"60",X"74",X"DE",X"56",X"47",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"37",X"37",X"33",X"11",X"11",X"00",X"00",
		X"47",X"CF",X"47",X"46",X"46",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"31",X"73",X"73",X"B7",X"3F",
		X"C0",X"40",X"60",X"64",X"DE",X"56",X"47",X"47",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"37",X"37",X"33",X"11",X"11",X"00",X"00",
		X"CF",X"47",X"47",X"46",X"CE",X"44",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"30",X"71",X"73",X"B7",X"B7",
		X"C0",X"C0",X"60",X"E8",X"74",X"56",X"56",X"CF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"37",X"37",X"33",X"11",X"11",X"00",X"00",
		X"47",X"47",X"47",X"CE",X"46",X"44",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"20",X"12",X"57",X"8F",X"0F",X"0F",X"00",X"17",X"2F",X"2F",X"C7",X"2F",X"2F",X"0F",
		X"06",X"CF",X"4F",X"2F",X"1E",X"2D",X"0F",X"8F",X"00",X"20",X"40",X"84",X"8C",X"6E",X"4E",X"8F",
		X"07",X"8F",X"9F",X"36",X"21",X"41",X"11",X"00",X"5F",X"2F",X"A7",X"1F",X"0F",X"0F",X"0F",X"CC",
		X"5F",X"0F",X"4F",X"4F",X"C7",X"A7",X"84",X"80",X"4E",X"AE",X"4E",X"0E",X"0C",X"48",X"20",X"00",
		X"00",X"00",X"01",X"83",X"63",X"31",X"32",X"47",X"00",X"00",X"CD",X"1F",X"4F",X"9F",X"0F",X"2F",
		X"00",X"40",X"4B",X"4B",X"CB",X"5F",X"2F",X"8F",X"00",X"00",X"00",X"1C",X"AC",X"CA",X"86",X"0C",
		X"07",X"13",X"32",X"21",X"41",X"01",X"00",X"00",X"9F",X"8F",X"4F",X"4F",X"6D",X"2D",X"21",X"20",
		X"5F",X"0F",X"CB",X"BD",X"5E",X"3F",X"4C",X"00",X"4C",X"CC",X"4C",X"88",X"00",X"80",X"40",X"00",
		X"00",X"10",X"00",X"01",X"23",X"81",X"71",X"12",X"00",X"00",X"B3",X"6B",X"3D",X"0F",X"DF",X"0F",
		X"10",X"10",X"1C",X"6D",X"7D",X"AF",X"0F",X"9E",X"00",X"00",X"00",X"88",X"5C",X"0C",X"E0",X"88",
		X"23",X"11",X"11",X"01",X"00",X"00",X"10",X"00",X"4F",X"CF",X"3F",X"6D",X"49",X"80",X"00",X"00",
		X"9F",X"2F",X"6B",X"BD",X"1C",X"00",X"00",X"00",X"4C",X"0C",X"0C",X"08",X"00",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"10",X"00",X"00",X"00",X"10",X"76",X"1E",X"8F",X"E7",
		X"00",X"00",X"00",X"00",X"8C",X"9E",X"AC",X"6B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"43",X"4F",X"1F",X"13",X"10",X"20",X"00",X"00",
		X"8F",X"6C",X"3E",X"84",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"31",
		X"00",X"00",X"00",X"00",X"00",X"40",X"88",X"64",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"11",X"62",
		X"00",X"00",X"00",X"00",X"80",X"A8",X"44",X"3A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"A8",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"22",X"00",X"C6",
		X"00",X"00",X"00",X"80",X"98",X"2A",X"00",X"13",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"2A",X"98",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"80",X"44",X"02",X"00",X"AC",
		X"00",X"00",X"80",X"88",X"19",X"82",X"00",X"21",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"C8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"44",X"80",X"00",X"00",X"00",X"00",
		X"00",X"82",X"19",X"88",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"04",
		X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"22",X"00",X"00",X"02",X"80",X"11",X"44",X"00",X"81",
		X"00",X"00",X"88",X"20",X"00",X"15",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",
		X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"10",X"80",X"02",X"00",X"00",X"00",
		X"00",X"15",X"00",X"20",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"00",X"22",X"00",X"41",X"00",X"01",X"44",X"00",X"22",X"80",X"11",X"20",
		X"00",X"00",X"40",X"11",X"80",X"02",X"00",X"91",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"44",
		X"00",X"22",X"00",X"01",X"00",X"00",X"00",X"00",X"11",X"88",X"20",X"00",X"44",X"10",X"00",X"00",
		X"00",X"20",X"08",X"11",X"44",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"11",X"00",X"00",X"07",X"1F",
		X"00",X"00",X"01",X"CF",X"16",X"96",X"3C",X"8F",X"00",X"00",X"80",X"C4",X"00",X"00",X"80",X"08",
		X"0F",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"F1",X"70",X"00",X"00",X"11",X"00",X"00",
		X"CF",X"F8",X"E1",X"87",X"43",X"ED",X"10",X"00",X"0C",X"80",X"80",X"00",X"00",X"C4",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"11",X"01",X"37",X"7F",
		X"00",X"00",X"12",X"9E",X"1E",X"2D",X"8F",X"CB",X"00",X"00",X"88",X"00",X"00",X"08",X"0C",X"C0",
		X"07",X"0F",X"70",X"00",X"00",X"00",X"00",X"00",X"1F",X"3C",X"D0",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"87",X"87",X"C3",X"30",X"FE",X"00",X"00",X"C0",X"08",X"08",X"80",X"E2",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"10",X"13",X"3F",
		X"00",X"00",X"71",X"E1",X"C3",X"87",X"CF",X"DA",X"00",X"00",X"00",X"00",X"08",X"08",X"80",X"48",
		X"03",X"07",X"1E",X"70",X"00",X"00",X"00",X"00",X"1E",X"3C",X"F0",X"80",X"00",X"00",X"00",X"00",
		X"C3",X"87",X"F0",X"10",X"66",X"00",X"00",X"00",X"48",X"2E",X"2C",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"32",X"30",X"33",
		X"00",X"00",X"70",X"E1",X"C3",X"87",X"8F",X"DA",X"00",X"00",X"88",X"00",X"08",X"08",X"80",X"0C",
		X"00",X"01",X"03",X"07",X"34",X"00",X"00",X"00",X"37",X"1E",X"0F",X"78",X"80",X"00",X"00",X"00",
		X"C3",X"87",X"C3",X"F0",X"11",X"22",X"00",X"00",X"3D",X"2C",X"68",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"30",X"30",X"65",X"73",X"77",
		X"00",X"C4",X"84",X"1E",X"3C",X"0F",X"87",X"87",X"00",X"00",X"00",X"00",X"00",X"A2",X"0C",X"48",
		X"00",X"00",X"00",X"01",X"01",X"03",X"12",X"00",X"76",X"0F",X"1E",X"2C",X"48",X"80",X"00",X"00",
		X"B4",X"D1",X"A2",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"21",X"21",X"21",X"32",X"76",
		X"00",X"08",X"0C",X"2C",X"5A",X"0F",X"0F",X"1E",X"00",X"00",X"00",X"00",X"44",X"48",X"C0",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"76",X"74",X"07",X"1E",X"1E",X"2C",X"68",X"C0",
		X"79",X"E2",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"11",X"33",X"33",
		X"00",X"0C",X"2C",X"5A",X"0F",X"0F",X"87",X"96",X"00",X"00",X"88",X"00",X"08",X"80",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"23",X"03",X"07",X"16",X"16",X"16",X"24",X"24",
		X"F0",X"E2",X"A2",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"16",X"07",X"03",X"03",X"21",X"23",X"33",
		X"00",X"08",X"79",X"96",X"0F",X"0F",X"87",X"B4",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"13",X"03",X"03",X"03",X"03",X"12",X"02",
		X"6A",X"6A",X"08",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E1",X"0F",X"16",X"12",X"03",X"23",X"33",
		X"00",X"00",X"E2",X"68",X"1E",X"1E",X"96",X"A4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"11",X"01",X"01",X"01",X"01",X"00",X"00",
		X"6A",X"6A",X"6A",X"48",X"48",X"48",X"48",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"0F",X"1E",X"07",X"07",X"23",X"33",
		X"00",X"44",X"E0",X"1E",X"1E",X"1E",X"3D",X"B5",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"11",X"01",X"01",X"00",X"00",X"00",X"00",
		X"F1",X"0C",X"2C",X"2C",X"2C",X"2C",X"2C",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"01",X"00",X"00",X"00",X"00",X"00",X"11",X"96",X"1E",X"1E",X"87",X"63",X"33",
		X"00",X"80",X"48",X"2C",X"2C",X"2C",X"3D",X"B5",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"11",X"01",X"00",X"00",X"00",X"00",X"00",
		X"C2",X"2C",X"2C",X"1E",X"1E",X"16",X"16",X"02",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"F0",X"1E",X"0F",X"87",X"F2",
		X"00",X"C8",X"68",X"2C",X"2C",X"0E",X"1F",X"3D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"73",X"33",X"11",X"00",X"00",X"00",X"00",X"00",
		X"A4",X"96",X"9E",X"0F",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"80",X"80",X"48",X"48",X"08",
		X"00",X"00",X"00",X"00",X"01",X"01",X"32",X"10",X"11",X"10",X"21",X"C3",X"0F",X"0F",X"3C",X"F3",
		X"80",X"C0",X"48",X"6A",X"59",X"48",X"2C",X"A4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F3",X"74",X"22",X"00",X"00",X"00",X"00",X"00",
		X"DA",X"8F",X"0F",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"80",X"48",X"48",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"32",X"B8",X"43",X"87",X"87",X"87",X"0F",X"1E",X"B6",
		X"00",X"80",X"80",X"80",X"C4",X"A2",X"48",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"F7",X"F3",X"44",X"22",X"00",X"00",X"00",X"00",
		X"96",X"8F",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",X"80",X"48",X"0C",X"0E",X"00",X"00",X"00",
		X"00",X"11",X"10",X"10",X"30",X"03",X"07",X"03",X"60",X"96",X"1E",X"1E",X"96",X"0F",X"0F",X"78",
		X"00",X"00",X"00",X"88",X"44",X"80",X"C0",X"68",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"74",X"30",X"10",X"00",X"00",X"00",X"00",X"00",X"F7",X"F3",X"B4",X"66",X"00",X"00",X"00",X"00",
		X"1E",X"8F",X"0F",X"01",X"00",X"00",X"00",X"00",X"00",X"80",X"48",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"22",X"10",X"10",X"10",X"03",X"07",X"03",X"C0",X"2C",X"1E",X"1E",X"87",X"0F",X"78",X"7F",
		X"00",X"00",X"88",X"E6",X"80",X"E0",X"F0",X"96",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"74",X"30",X"10",X"00",X"00",X"00",X"00",X"00",X"F7",X"F0",X"E6",X"00",X"00",X"00",X"00",X"00",
		X"8F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"2C",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"88",X"FF",X"00",X"FF",
		X"00",X"00",X"00",X"EE",X"22",X"EE",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"FF",X"00",X"99",X"99",X"FF",X"00",X"00",
		X"22",X"EE",X"00",X"EE",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"88",X"FF",X"00",X"FF",X"88",X"FF",X"00",
		X"EE",X"22",X"EE",X"00",X"EE",X"22",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"88",X"FF",X"00",X"00",X"FF",X"44",X"00",
		X"EE",X"22",X"EE",X"00",X"22",X"EE",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"FF",X"00",X"00",X"FF",X"44",X"00",
		X"EE",X"22",X"22",X"00",X"22",X"EE",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"88",X"FF",X"00",X"FF",X"88",X"FF",X"00",
		X"EE",X"22",X"EE",X"00",X"EE",X"22",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"88",X"FF",X"00",X"FF",X"88",X"FF",X"00",
		X"EE",X"22",X"EE",X"00",X"EE",X"22",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"88",X"FF",X"00",X"FF",X"99",X"99",X"00",
		X"EE",X"22",X"EE",X"00",X"22",X"22",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"88",X"FF",X"00",X"FF",X"99",X"99",X"00",
		X"EE",X"22",X"EE",X"00",X"EE",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"88",X"FF",X"00",X"FF",X"88",X"FF",X"00",
		X"EE",X"22",X"EE",X"00",X"EE",X"22",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
