library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity obj1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of obj1 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"1F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"1F",X"1F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"07",
		X"00",X"1C",X"1E",X"14",X"00",X"0F",X"07",X"03",X"07",X"07",X"79",X"FE",X"FF",X"CF",X"CF",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"01",X"00",X"01",X"01",X"07",X"0F",X"1F",X"27",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"0F",X"00",X"3F",X"3E",X"7F",X"EF",X"CF",X"CF",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"0F",X"00",X"3F",X"3F",X"7F",X"EF",X"CF",X"CF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"07",X"3F",X"7F",X"EF",X"CF",X"CF",X"CF",X"EF",X"7F",X"3F",X"3F",X"F9",X"F7",
		X"00",X"00",X"03",X"07",X"3F",X"7F",X"EF",X"CF",X"CF",X"CF",X"EF",X"7F",X"3F",X"1F",X"3C",X"3D",
		X"00",X"00",X"04",X"1C",X"65",X"E7",X"1F",X"1F",X"1F",X"55",X"4C",X"44",X"04",X"00",X"00",X"00",
		X"00",X"00",X"04",X"1C",X"64",X"E1",X"F9",X"E9",X"C1",X"55",X"4C",X"44",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"0E",X"32",X"71",X"1F",X"1F",X"1F",X"2A",X"26",X"22",X"02",X"00",X"00",
		X"00",X"00",X"00",X"02",X"0E",X"32",X"70",X"7C",X"74",X"60",X"2A",X"26",X"22",X"02",X"00",X"00",
		X"00",X"03",X"07",X"07",X"0F",X"0F",X"1F",X"1F",X"1F",X"0F",X"0F",X"1C",X"3F",X"3F",X"7F",X"7F",
		X"00",X"00",X"00",X"78",X"FC",X"FC",X"F8",X"FC",X"7E",X"7F",X"3F",X"3F",X"3F",X"7F",X"7F",X"FF",
		X"00",X"00",X"00",X"0C",X"BF",X"FF",X"FF",X"FF",X"7F",X"E7",X"C3",X"C3",X"47",X"1F",X"3F",X"7F",
		X"1F",X"0F",X"07",X"03",X"07",X"37",X"3F",X"3F",X"3F",X"37",X"07",X"03",X"07",X"0F",X"1F",X"00",
		X"00",X"00",X"00",X"00",X"05",X"06",X"07",X"09",X"0F",X"1F",X"3F",X"7F",X"7F",X"7E",X"78",X"21",
		X"00",X"00",X"00",X"00",X"0A",X"0C",X"0F",X"13",X"1F",X"0F",X"07",X"07",X"03",X"03",X"01",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"03",X"03",X"07",X"0D",X"03",X"07",X"03",
		X"04",X"1C",X"65",X"E1",X"F9",X"E8",X"C0",X"55",X"4C",X"44",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"1C",X"65",X"E1",X"F9",X"E9",X"C1",X"55",X"4C",X"44",X"04",X"00",X"00",X"00",X"00",
		X"00",X"04",X"1C",X"65",X"E1",X"F9",X"E9",X"C1",X"54",X"4C",X"45",X"05",X"01",X"00",X"00",X"00",
		X"00",X"02",X"0E",X"32",X"70",X"7C",X"74",X"60",X"2A",X"26",X"22",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"0E",X"32",X"70",X"7C",X"74",X"60",X"2A",X"26",X"22",X"02",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"03",X"03",X"01",X"01",X"00",X"00",
		X"00",X"02",X"0D",X"06",X"07",X"03",X"03",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"07",X"07",X"3F",X"07",X"07",X"07",X"03",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"03",X"07",X"0B",X"2A",X"2B",X"2B",X"16",X"0B",X"07",X"03",X"01",X"00",X"00",
		X"03",X"07",X"05",X"08",X"1B",X"19",X"05",X"3F",X"3F",X"0F",X"05",X"37",X"3F",X"3F",X"3E",X"1C",
		X"00",X"01",X"0D",X"1C",X"61",X"C9",X"ED",X"C7",X"C7",X"ED",X"C9",X"61",X"9C",X"0D",X"01",X"00",
		X"03",X"07",X"0F",X"1F",X"3F",X"7F",X"79",X"79",X"7F",X"79",X"79",X"7F",X"3F",X"1F",X"0F",X"07",
		X"03",X"07",X"0F",X"1F",X"3F",X"7F",X"79",X"79",X"7F",X"79",X"79",X"7F",X"3F",X"1F",X"0F",X"07",
		X"00",X"80",X"00",X"80",X"00",X"85",X"44",X"88",X"70",X"88",X"44",X"85",X"00",X"80",X"00",X"80",
		X"54",X"86",X"45",X"89",X"4B",X"B7",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"1F",X"0F",X"00",X"00",
		X"00",X"00",X"00",X"01",X"07",X"8F",X"DF",X"FF",X"FF",X"FF",X"B7",X"4B",X"89",X"45",X"86",X"54",
		X"00",X"18",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"B7",X"4B",X"89",X"45",X"86",X"54",
		X"00",X"00",X"09",X"00",X"00",X"08",X"08",X"08",X"08",X"04",X"04",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"3F",X"3F",X"7F",X"5F",X"EF",X"F6",X"AC",X"CD",X"68",X"23",X"07",
		X"07",X"03",X"08",X"1A",X"33",X"2B",X"3D",X"3B",X"17",X"1F",X"0F",X"07",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"03",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"06",X"04",X"04",X"01",X"06",X"0E",
		X"00",X"00",X"00",X"00",X"C0",X"78",X"00",X"00",X"00",X"00",X"00",X"17",X"E7",X"87",X"06",X"06",
		X"7F",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"41",X"42",X"44",X"48",X"10",X"00",X"0F",X"00",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"00",X"0F",X"00",X"13",X"4B",X"53",X"53",X"4B",X"47",X"43",X"43",X"43",X"43",X"40",X"40",X"7F",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"01",X"01",X"02",X"02",X"02",X"04",X"04",X"04",X"08",X"08",X"08",X"08",X"08",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"10",X"08",X"00",X"00",X"00",X"00",X"04",X"18",X"00",X"00",X"00",X"00",X"02",X"00",X"00",
		X"17",X"2F",X"1F",X"2F",X"3F",X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"0C",X"06",X"06",X"06",X"04",X"08",X"10",X"20",X"00",X"80",X"60",X"18",X"0C",X"00",X"00",
		X"00",X"18",X"20",X"40",X"80",X"00",X"00",X"21",X"11",X"09",X"04",X"04",X"06",X"06",X"06",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3C",X"1F",X"0F",X"07",X"07",X"07",X"00",X"00",X"00",X"07",X"07",X"07",X"0F",X"1F",X"3C",X"00",
		X"01",X"03",X"05",X"06",X"00",X"00",X"00",X"0F",X"1F",X"3F",X"3F",X"3F",X"3E",X"38",X"10",X"00",
		X"01",X"03",X"05",X"06",X"00",X"00",X"00",X"03",X"07",X"07",X"07",X"03",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"03",X"01",X"00",X"01",X"03",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"00",X"11",X"02",X"05",X"0D",X"0F",X"0D",X"05",X"42",X"01",X"00",X"04",X"00",X"00",
		X"00",X"00",X"00",X"00",X"09",X"02",X"05",X"05",X"05",X"02",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"02",X"05",X"0B",X"0B",X"0B",X"0B",X"05",X"02",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"02",X"05",X"04",X"04",X"05",X"02",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"05",X"08",X"00",X"00",X"00",X"03",X"01",X"00",X"00",X"05",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"E0",X"BF",X"BF",X"E0",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"01",X"00",X"00",X"00",
		X"80",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"7F",X"80",
		X"00",X"00",X"00",X"00",X"07",X"03",X"0B",X"0C",X"0C",X"0F",X"06",X"06",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"01",X"06",X"0D",X"05",X"07",X"02",X"07",X"02",X"02",X"01",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"1F",X"3B",X"33",X"33",X"39",X"18",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"29",X"2B",X"2B",X"27",X"27",X"03",X"03",X"02",X"02",X"02",X"03",
		X"00",X"00",X"00",X"00",X"00",X"11",X"2B",X"4B",X"47",X"87",X"03",X"01",X"01",X"01",X"01",X"00",
		X"07",X"0F",X"1E",X"3F",X"3F",X"7F",X"7E",X"7E",X"7F",X"7E",X"7F",X"3F",X"3F",X"1E",X"0F",X"07",
		X"C0",X"C0",X"C1",X"C2",X"CE",X"DC",X"F0",X"F9",X"F9",X"F0",X"DC",X"CE",X"C2",X"C1",X"C0",X"C0",
		X"0C",X"0C",X"0C",X"0C",X"0D",X"0D",X"0F",X"0F",X"0F",X"0F",X"0D",X"0D",X"0C",X"0C",X"0C",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E1",X"E3",X"61",X"65",X"60",X"60",X"60",
		X"60",X"60",X"60",X"60",X"68",X"88",X"68",X"68",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",
		X"60",X"E0",X"E0",X"E1",X"E3",X"E5",X"E6",X"E1",X"C0",X"80",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C8",X"C8",X"C8",X"C8",X"C8",X"C8",X"C8",X"C8",X"C8",X"C8",X"C8",X"C8",
		X"C8",X"C8",X"C8",X"90",X"30",X"60",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"80",X"80",X"C0",X"E0",X"E0",X"E0",X"E0",X"E1",X"63",X"61",X"65",X"20",X"00",X"00",
		X"40",X"60",X"60",X"60",X"68",X"68",X"88",X"68",X"60",X"60",X"60",X"40",X"00",X"00",X"20",X"60",
		X"60",X"60",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"9F",X"9F",X"8D",X"06",X"02",X"06",X"00",X"00",
		X"40",X"80",X"89",X"01",X"18",X"18",X"4E",X"01",X"00",X"07",X"3C",X"38",X"31",X"00",X"88",X"80",
		X"01",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"32",X"18",X"00",X"00",
		X"00",X"7F",X"C0",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"C0",X"7F",X"00",
		X"00",X"03",X"04",X"08",X"10",X"20",X"20",X"20",X"20",X"20",X"20",X"10",X"08",X"04",X"03",X"00",
		X"00",X"00",X"00",X"01",X"02",X"04",X"08",X"08",X"08",X"08",X"04",X"02",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"04",X"04",X"02",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"04",X"00",X"00",X"00",X"18",X"00",X"00",X"00",X"04",X"08",X"00",X"00",
		X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"CF",X"BF",X"1E",X"1E",X"0C",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"CF",X"BF",X"1F",X"1E",X"0C",X"00",X"00",X"00",X"00",
		X"1F",X"3F",X"3F",X"7F",X"7F",X"7F",X"7F",X"67",X"DF",X"0F",X"0F",X"06",X"00",X"00",X"00",X"00",
		X"3F",X"3F",X"3F",X"3F",X"18",X"0C",X"1F",X"1F",X"3E",X"7C",X"F8",X"00",X"A0",X"F0",X"E0",X"00",
		X"63",X"77",X"7F",X"7F",X"3F",X"1F",X"07",X"0F",X"1F",X"3F",X"7E",X"00",X"A0",X"F0",X"00",X"00",
		X"CF",X"EF",X"7F",X"3E",X"3F",X"00",X"0F",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CF",X"EF",X"7F",X"3F",X"3F",X"00",X"0F",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"78",X"F0",X"F0",X"D0",X"80",X"00",X"00",X"00",X"00",X"20",X"70",X"78",X"7E",X"3E",X"1C",
		X"F7",X"E7",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"39",X"39",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"30",X"38",X"38",X"7C",X"7C",X"1E",X"1F",X"0F",X"0F",X"0F",X"07",X"07",X"27",X"8B",
		X"FB",X"8B",X"2F",X"0F",X"0F",X"1F",X"3F",X"3E",X"FC",X"F8",X"70",X"F0",X"60",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"0C",X"0E",X"0F",X"0F",X"07",X"03",X"00",
		X"7F",X"67",X"7F",X"3F",X"0F",X"7F",X"FF",X"FF",X"7E",X"F0",X"20",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"EF",X"C7",X"CF",X"47",X"2F",X"7E",X"7C",X"7C",X"2E",X"3C",X"0C",X"00",X"00",X"00",
		X"CF",X"CF",X"EF",X"CF",X"CF",X"7F",X"3F",X"5F",X"C7",X"E7",X"7F",X"FF",X"FF",X"FF",X"BF",X"0E",
		X"00",X"00",X"00",X"01",X"03",X"07",X"07",X"0F",X"0F",X"0F",X"0C",X"07",X"00",X"00",X"00",X"00",
		X"01",X"03",X"03",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"0F",X"0F",X"2F",X"8B",X"FB",
		X"FB",X"03",X"27",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"0F",X"0F",X"07",X"0F",X"06",
		X"00",X"00",X"30",X"38",X"38",X"7C",X"7C",X"1E",X"1F",X"0F",X"0F",X"0F",X"07",X"07",X"27",X"8B",
		X"07",X"08",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"08",X"07",X"00",X"00",X"0F",X"04",X"00",
		X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"07",X"00",X"06",X"09",X"08",X"08",X"04",X"00",
		X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"07",X"00",X"08",X"0D",X"0B",X"09",X"08",X"00",
		X"07",X"08",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"08",X"07",X"00",X"0F",X"04",X"02",X"01",
		X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"07",X"00",X"06",X"09",X"09",X"09",X"06",X"00",
		X"07",X"08",X"07",X"00",X"07",X"08",X"07",X"00",X"06",X"09",X"08",X"04",X"00",X"0F",X"04",X"00",
		X"07",X"08",X"07",X"00",X"07",X"08",X"07",X"00",X"04",X"09",X"09",X"07",X"00",X"0F",X"04",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
