library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity cpu3_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of cpu3_rom is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"54",X"20",X"20",X"30",X"40",X"43",X"89",X"0F",X"31",X"50",X"20",X"55",X"50",X"20",X"20",X"20",
		X"20",X"20",X"30",X"20",X"20",X"20",X"32",X"50",X"20",X"55",X"50",X"20",X"20",X"20",X"20",X"20",
		X"30",X"40",X"43",X"8B",X"0F",X"31",X"50",X"20",X"44",X"4F",X"57",X"4E",X"20",X"20",X"20",X"30",
		X"20",X"20",X"20",X"32",X"50",X"20",X"44",X"4F",X"57",X"4E",X"20",X"20",X"20",X"30",X"40",X"43",
		X"8D",X"0F",X"31",X"50",X"20",X"53",X"48",X"4F",X"54",X"31",X"20",X"20",X"30",X"20",X"20",X"20",
		X"32",X"50",X"20",X"53",X"48",X"4F",X"54",X"31",X"20",X"20",X"30",X"40",X"43",X"8F",X"0F",X"31",
		X"50",X"20",X"53",X"48",X"4F",X"54",X"32",X"20",X"20",X"30",X"20",X"20",X"20",X"32",X"50",X"20",
		X"53",X"48",X"4F",X"54",X"32",X"20",X"20",X"30",X"40",X"42",X"B2",X"0F",X"43",X"4F",X"49",X"4E",
		X"31",X"20",X"20",X"20",X"20",X"20",X"30",X"40",X"42",X"B4",X"0F",X"43",X"4F",X"49",X"4E",X"32",
		X"20",X"20",X"20",X"20",X"20",X"30",X"40",X"42",X"B6",X"0F",X"53",X"45",X"52",X"56",X"49",X"43",
		X"45",X"20",X"20",X"20",X"30",X"40",X"42",X"B8",X"0F",X"31",X"50",X"20",X"53",X"54",X"41",X"52",
		X"54",X"20",X"20",X"30",X"40",X"42",X"BA",X"0F",X"32",X"50",X"20",X"53",X"54",X"41",X"52",X"54",
		X"20",X"20",X"30",X"40",X"43",X"09",X"0F",X"43",X"4F",X"49",X"4E",X"20",X"43",X"4F",X"55",X"4E",
		X"54",X"45",X"52",X"20",X"31",X"40",X"43",X"67",X"0F",X"46",X"52",X"45",X"45",X"20",X"20",X"50",
		X"4C",X"41",X"59",X"40",X"43",X"67",X"0F",X"49",X"4E",X"56",X"41",X"4C",X"49",X"44",X"49",X"54",
		X"59",X"40",X"42",X"C3",X"0F",X"44",X"49",X"50",X"53",X"57",X"20",X"20",X"20",X"53",X"45",X"4C",
		X"45",X"43",X"54",X"40",X"43",X"66",X"0F",X"43",X"4F",X"49",X"4E",X"31",X"40",X"43",X"68",X"0F",
		X"43",X"4F",X"49",X"4E",X"32",X"40",X"43",X"6B",X"0F",X"42",X"4F",X"4E",X"55",X"53",X"20",X"20",
		X"50",X"4F",X"49",X"4E",X"54",X"40",X"42",X"CE",X"0F",X"46",X"49",X"52",X"53",X"54",X"20",X"20",
		X"20",X"20",X"30",X"30",X"30",X"30",X"20",X"50",X"4F",X"49",X"4E",X"54",X"53",X"40",X"42",X"D0",
		X"0F",X"45",X"56",X"45",X"52",X"59",X"20",X"20",X"20",X"20",X"30",X"30",X"30",X"30",X"20",X"50",
		X"4F",X"49",X"4E",X"54",X"53",X"40",X"43",X"74",X"0F",X"44",X"45",X"4D",X"4F",X"20",X"20",X"53",
		X"4F",X"55",X"4E",X"44",X"20",X"20",X"4F",X"40",X"43",X"76",X"0F",X"50",X"4C",X"41",X"59",X"45",
		X"52",X"40",X"43",X"78",X"0F",X"54",X"41",X"42",X"4C",X"45",X"20",X"20",X"20",X"40",X"43",X"78",
		X"0F",X"55",X"50",X"20",X"52",X"49",X"47",X"48",X"54",X"40",X"42",X"E5",X"0F",X"53",X"4F",X"55",
		X"4E",X"44",X"20",X"20",X"20",X"54",X"45",X"53",X"54",X"40",X"43",X"09",X"0F",X"53",X"4F",X"55",
		X"4E",X"44",X"20",X"43",X"4F",X"44",X"45",X"40",X"43",X"28",X"07",X"52",X"41",X"4D",X"20",X"20",
		X"20",X"42",X"41",X"44",X"40",X"41",X"A8",X"0F",X"52",X"41",X"4D",X"20",X"20",X"20",X"20",X"4F",
		X"4B",X"40",X"41",X"AB",X"0F",X"52",X"4F",X"4D",X"20",X"20",X"20",X"20",X"4F",X"4B",X"40",X"41",
		X"A8",X"07",X"52",X"41",X"4D",X"20",X"20",X"20",X"42",X"41",X"44",X"40",X"41",X"AB",X"07",X"52",
		X"4F",X"4D",X"20",X"20",X"20",X"42",X"41",X"44",X"40",X"42",X"E6",X"0F",X"4D",X"41",X"49",X"4E",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"53",X"55",X"42",X"40",X"42",X"26",X"0F",X"43",
		X"4F",X"49",X"4E",X"40",X"41",X"06",X"0F",X"50",X"4C",X"41",X"59",X"40",X"42",X"28",X"0F",X"43",
		X"4F",X"49",X"4E",X"40",X"41",X"08",X"0F",X"50",X"4C",X"41",X"59",X"40",X"47",X"BE",X"0F",X"54",
		X"48",X"49",X"53",X"20",X"49",X"53",X"20",X"41",X"4E",X"20",X"49",X"4C",X"4C",X"45",X"47",X"41",
		X"4C",X"20",X"44",X"55",X"50",X"4C",X"49",X"43",X"41",X"54",X"45",X"40",X"47",X"BF",X"0F",X"4F",
		X"46",X"20",X"4B",X"4F",X"4E",X"41",X"4D",X"49",X"5D",X"53",X"20",X"4F",X"52",X"49",X"47",X"49",
		X"4E",X"41",X"4C",X"20",X"50",X"43",X"42",X"4F",X"41",X"52",X"44",X"40",X"42",X"BA",X"0B",X"80",
		X"81",X"95",X"96",X"B0",X"B1",X"B2",X"F0",X"F2",X"FD",X"FE",X"40",X"42",X"BB",X"0B",X"90",X"91",
		X"A0",X"A1",X"A2",X"A3",X"C0",X"F1",X"FC",X"EF",X"FF",X"40",X"00",X"01",X"02",X"03",X"05",X"10",
		X"20",X"30",X"50",X"80",X"0B",X"10",X"11",X"40",X"14",X"70",X"15",X"80",X"14",X"A0",X"10",X"B0",
		X"0F",X"B0",X"09",X"80",X"07",X"90",X"03",X"90",X"8A",X"8B",X"8C",X"8D",X"8E",X"8F",X"80",X"81",
		X"82",X"83",X"84",X"97",X"98",X"99",X"9A",X"9B",X"9C",X"9D",X"9E",X"9F",X"90",X"91",X"92",X"93",
		X"94",X"95",X"96",X"97",X"A4",X"A5",X"A6",X"A7",X"A8",X"A9",X"AA",X"AB",X"AC",X"AD",X"AE",X"AF",
		X"A0",X"A1",X"A2",X"A3",X"A4",X"A5",X"A6",X"A7",X"B3",X"B4",X"B5",X"B6",X"B7",X"B8",X"B9",X"BA",
		X"BB",X"BC",X"BD",X"BE",X"BF",X"B0",X"B1",X"B2",X"B3",X"B4",X"B5",X"B6",X"B7",X"C1",X"C2",X"C3",
		X"C4",X"C5",X"C6",X"C7",X"C8",X"C9",X"CA",X"CB",X"CC",X"CD",X"CE",X"CF",X"C0",X"C1",X"C2",X"C3",
		X"C4",X"D0",X"D1",X"D2",X"D3",X"D4",X"D5",X"D6",X"D7",X"D8",X"D9",X"DA",X"DB",X"DC",X"DD",X"DE",
		X"DF",X"E0",X"E1",X"E2",X"E3",X"E4",X"E5",X"E6",X"E7",X"E8",X"E9",X"EA",X"EB",X"EC",X"ED",X"EE",
		X"F3",X"F4",X"F5",X"F6",X"F7",X"F8",X"F9",X"FA",X"FB",X"82",X"83",X"84",X"85",X"86",X"87",X"88",
		X"92",X"93",X"94",X"09",X"09",X"09",X"08",X"08",X"08",X"35",X"35",X"35",X"38",X"38",X"09",X"0A",
		X"0A",X"00",X"00",X"09",X"05",X"05",X"05",X"36",X"36",X"36",X"36",X"38",X"38",X"38",X"38",X"0C",
		X"01",X"0A",X"0A",X"0A",X"0A",X"09",X"03",X"05",X"05",X"05",X"05",X"36",X"36",X"36",X"36",X"36",
		X"36",X"36",X"35",X"01",X"01",X"0A",X"0A",X"0A",X"02",X"0F",X"05",X"05",X"05",X"05",X"05",X"05",
		X"37",X"36",X"36",X"36",X"37",X"37",X"37",X"37",X"01",X"01",X"01",X"0A",X"0A",X"0F",X"0F",X"0F",
		X"05",X"05",X"05",X"06",X"08",X"08",X"05",X"37",X"35",X"35",X"35",X"35",X"01",X"01",X"01",X"01",
		X"01",X"0F",X"0F",X"04",X"04",X"06",X"08",X"08",X"06",X"07",X"05",X"05",X"01",X"01",X"05",X"05",
		X"05",X"04",X"04",X"06",X"06",X"06",X"07",X"06",X"07",X"07",X"05",X"05",X"05",X"05",X"05",X"06",
		X"07",X"07",X"07",X"07",X"05",X"05",X"07",X"07",X"07",X"07",X"07",X"05",X"07",X"07",X"85",X"3B",
		X"86",X"8A",X"86",X"A1",X"86",X"EB",X"87",X"31",X"87",X"7D",X"87",X"A9",X"87",X"CE",X"89",X"02",
		X"89",X"13",X"89",X"4C",X"89",X"CA",X"8A",X"CC",X"8A",X"E4",X"8A",X"F5",X"8B",X"28",X"8B",X"C4",
		X"8B",X"C8",X"05",X"00",X"01",X"06",X"00",X"02",X"07",X"00",X"03",X"08",X"00",X"04",X"20",X"41",
		X"42",X"43",X"44",X"45",X"46",X"47",X"48",X"49",X"4A",X"4B",X"4C",X"4D",X"4E",X"4F",X"50",X"51",
		X"52",X"53",X"54",X"55",X"56",X"57",X"58",X"59",X"5A",X"2E",X"00",X"00",X"00",X"00",X"00",X"01",
		X"02",X"0E",X"8D",X"0B",X"8D",X"7A",X"8E",X"03",X"8E",X"03",X"8E",X"2C",X"8E",X"37",X"A8",X"42",
		X"4F",X"B5",X"42",X"6C",X"C2",X"42",X"5B",X"CF",X"42",X"44",X"A5",X"4C",X"41",X"B5",X"4C",X"75",
		X"A8",X"56",X"58",X"B7",X"56",X"69",X"C6",X"56",X"38",X"D5",X"56",X"54",X"A4",X"60",X"5F",X"B4",
		X"60",X"4B",X"C4",X"60",X"71",X"47",X"41",X"4D",X"45",X"20",X"4F",X"56",X"45",X"52",X"25",X"23",
		X"28",X"15",X"20",X"18",X"2C",X"15",X"1A",X"00",X"2F",X"04",X"10",X"00",X"0B",X"04",X"10",X"05",
		X"01",X"01",X"08",X"05",X"01",X"04",X"18",X"01",X"0E",X"05",X"01",X"04",X"10",X"05",X"01",X"01",
		X"06",X"04",X"0D",X"01",X"19",X"04",X"0D",X"01",X"07",X"09",X"03",X"08",X"17",X"0A",X"03",X"02",
		X"09",X"0A",X"01",X"08",X"09",X"09",X"02",X"01",X"12",X"09",X"01",X"08",X"0D",X"0A",X"03",X"02",
		X"0F",X"0A",X"01",X"08",X"0A",X"0A",X"01",X"02",X"07",X"0A",X"01",X"08",X"10",X"0A",X"01",X"02",
		X"09",X"08",X"0A",X"09",X"0B",X"08",X"10",X"0A",X"06",X"08",X"13",X"02",X"0E",X"06",X"03",X"04",
		X"18",X"02",X"08",X"0A",X"02",X"08",X"26",X"09",X"01",X"01",X"07",X"09",X"01",X"08",X"09",X"0A",
		X"06",X"02",X"03",X"08",X"05",X"09",X"0E",X"08",X"12",X"0A",X"05",X"08",X"0E",X"0A",X"01",X"02",
		X"0F",X"0A",X"01",X"08",X"0C",X"09",X"02",X"01",X"18",X"08",X"0A",X"01",X"0C",X"09",X"04",X"08",
		X"14",X"0A",X"09",X"08",X"07",X"0A",X"0B",X"02",X"10",X"08",X"0D",X"02",X"0F",X"0A",X"01",X"08",
		X"0E",X"0A",X"01",X"02",X"12",X"08",X"1E",X"09",X"07",X"01",X"24",X"04",X"0D",X"06",X"0C",X"04",
		X"07",X"06",X"02",X"02",X"18",X"06",X"07",X"02",X"10",X"06",X"01",X"04",X"06",X"06",X"01",X"02",
		X"0B",X"0A",X"07",X"02",X"0A",X"06",X"09",X"02",X"17",X"06",X"0D",X"02",X"09",X"0A",X"0F",X"02",
		X"19",X"06",X"06",X"04",X"07",X"06",X"01",X"02",X"0B",X"0A",X"01",X"08",X"19",X"0A",X"01",X"02",
		X"09",X"06",X"04",X"04",X"0C",X"05",X"02",X"01",X"23",X"05",X"01",X"04",X"17",X"06",X"02",X"02",
		X"17",X"0A",X"04",X"08",X"0E",X"0A",X"03",X"02",X"12",X"0A",X"01",X"08",X"06",X"0A",X"01",X"02",
		X"13",X"0A",X"01",X"08",X"1D",X"09",X"01",X"01",X"16",X"04",X"0A",X"06",X"01",X"02",X"1A",X"0A",
		X"07",X"08",X"1B",X"01",X"0F",X"09",X"05",X"01",X"0B",X"09",X"01",X"08",X"08",X"0A",X"0B",X"08",
		X"08",X"0A",X"04",X"02",X"15",X"06",X"03",X"04",X"11",X"01",X"11",X"05",X"01",X"04",X"07",X"06",
		X"02",X"02",X"0D",X"0A",X"03",X"08",X"27",X"09",X"02",X"01",X"23",X"04",X"13",X"06",X"02",X"02",
		X"0D",X"06",X"01",X"04",X"03",X"05",X"01",X"01",X"17",X"09",X"02",X"08",X"15",X"0A",X"02",X"02",
		X"1E",X"0A",X"02",X"08",X"07",X"0A",X"01",X"02",X"05",X"06",X"01",X"04",X"0C",X"05",X"02",X"01",
		X"1E",X"09",X"0A",X"01",X"0A",X"04",X"10",X"05",X"01",X"01",X"09",X"09",X"09",X"08",X"16",X"09",
		X"01",X"01",X"1A",X"09",X"04",X"08",X"07",X"09",X"05",X"01",X"06",X"09",X"03",X"08",X"32",X"00",
		X"65",X"00",X"1D",X"02",X"23",X"00",X"24",X"02",X"14",X"0A",X"03",X"08",X"1A",X"02",X"0D",X"08",
		X"15",X"02",X"14",X"0A",X"01",X"08",X"1D",X"02",X"11",X"06",X"02",X"04",X"0F",X"05",X"01",X"01",
		X"07",X"04",X"04",X"06",X"04",X"04",X"02",X"01",X"0D",X"09",X"01",X"08",X"0F",X"0A",X"19",X"08",
		X"11",X"02",X"23",X"06",X"0C",X"02",X"0A",X"0A",X"03",X"08",X"14",X"09",X"01",X"01",X"10",X"04",
		X"0E",X"06",X"01",X"02",X"1C",X"0A",X"04",X"08",X"0F",X"09",X"12",X"01",X"0F",X"09",X"01",X"08",
		X"0B",X"0A",X"02",X"02",X"1A",X"0A",X"01",X"08",X"09",X"0A",X"01",X"02",X"05",X"0A",X"01",X"08",
		X"0A",X"02",X"14",X"0A",X"03",X"02",X"0F",X"08",X"0E",X"09",X"03",X"01",X"16",X"04",X"15",X"01",
		X"11",X"09",X"02",X"08",X"17",X"0A",X"03",X"02",X"03",X"08",X"03",X"01",X"19",X"05",X"01",X"04",
		X"1A",X"06",X"01",X"02",X"09",X"08",X"20",X"0A",X"01",X"02",X"1C",X"06",X"03",X"04",X"0C",X"01",
		X"0F",X"04",X"0C",X"01",X"19",X"04",X"18",X"01",X"10",X"09",X"02",X"08",X"15",X"0A",X"0A",X"08",
		X"08",X"09",X"01",X"01",X"19",X"04",X"0F",X"06",X"02",X"02",X"04",X"04",X"01",X"00",X"01",X"01",
		X"1A",X"05",X"01",X"04",X"0D",X"01",X"09",X"09",X"02",X"08",X"18",X"09",X"01",X"01",X"0E",X"09",
		X"01",X"08",X"08",X"01",X"08",X"05",X"01",X"04",X"0C",X"06",X"03",X"02",X"2D",X"08",X"13",X"02",
		X"1F",X"0A",X"01",X"08",X"19",X"0A",X"01",X"02",X"12",X"06",X"01",X"04",X"1D",X"02",X"13",X"04",
		X"05",X"01",X"1B",X"09",X"02",X"08",X"0D",X"0A",X"05",X"02",X"0A",X"0A",X"02",X"08",X"0C",X"09",
		X"06",X"08",X"03",X"0A",X"01",X"02",X"1B",X"06",X"01",X"04",X"0D",X"05",X"01",X"01",X"18",X"04",
		X"08",X"06",X"01",X"02",X"15",X"0A",X"02",X"08",X"28",X"02",X"0C",X"0A",X"01",X"08",X"0A",X"0A",
		X"01",X"02",X"0C",X"0A",X"01",X"08",X"0C",X"09",X"0A",X"01",X"13",X"05",X"01",X"04",X"07",X"01",
		X"06",X"09",X"02",X"08",X"15",X"01",X"1A",X"09",X"01",X"08",X"11",X"0A",X"06",X"02",X"0E",X"06",
		X"05",X"04",X"0E",X"02",X"04",X"08",X"18",X"09",X"02",X"01",X"17",X"08",X"13",X"01",X"0E",X"05",
		X"01",X"04",X"13",X"06",X"01",X"02",X"26",X"04",X"0E",X"05",X"04",X"01",X"07",X"04",X"11",X"01",
		X"12",X"04",X"17",X"05",X"03",X"01",X"12",X"04",X"0E",X"06",X"03",X"02",X"24",X"0A",X"02",X"08",
		X"0E",X"09",X"01",X"01",X"0B",X"09",X"01",X"08",X"05",X"0A",X"06",X"02",X"17",X"08",X"17",X"09",
		X"03",X"01",X"0F",X"04",X"14",X"06",X"03",X"02",X"15",X"0A",X"02",X"08",X"0F",X"09",X"05",X"01",
		X"1E",X"04",X"09",X"01",X"1D",X"09",X"02",X"08",X"27",X"0A",X"05",X"02",X"12",X"06",X"05",X"04",
		X"13",X"01",X"1D",X"09",X"04",X"08",X"0E",X"01",X"17",X"04",X"10",X"06",X"01",X"02",X"21",X"0A",
		X"01",X"08",X"09",X"0A",X"01",X"02",X"0B",X"06",X"04",X"04",X"0E",X"05",X"01",X"01",X"11",X"00",
		X"01",X"04",X"24",X"00",X"D5",X"8E",X"44",X"8E",X"B3",X"8E",X"C9",X"30",X"31",X"32",X"33",X"34",
		X"35",X"36",X"37",X"38",X"39",X"42",X"50",X"41",X"30",X"42",X"52",X"41",X"32",X"42",X"54",X"41",
		X"34",X"42",X"56",X"41",X"36",X"42",X"58",X"41",X"38",X"00",X"01",X"02",X"03",X"04",X"00",X"01",
		X"02",X"03",X"05",X"00",X"01",X"02",X"04",X"05",X"00",X"01",X"03",X"04",X"05",X"00",X"02",X"03",
		X"04",X"05",X"01",X"02",X"03",X"04",X"05",X"1D",X"1C",X"03",X"02",X"01",X"00",X"02",X"02",X"FE",
		X"FE",X"02",X"FE",X"02",X"FE",X"F0",X"BC",X"EF",X"FA",X"E0",X"10",X"EF",X"FA",X"F0",X"BC",X"F0",
		X"5B",X"EF",X"FA",X"F0",X"BC",X"F0",X"5B",X"EB",X"CF",X"F1",X"1D",X"EF",X"FA",X"EC",X"91",X"E3",
		X"79",X"D3",X"F0",X"D0",X"E8",X"D0",X"87",X"D1",X"AA",X"D2",X"6C",X"D0",X"E8",X"D0",X"87",X"D1",
		X"AA",X"D2",X"6C",X"D3",X"2E",X"D1",X"49",X"D6",X"F8",X"E0",X"71",X"F0",X"BC",X"F1",X"1D",X"F0",
		X"5B",X"F0",X"BC",X"DA",X"00",X"F1",X"1D",X"F0",X"5B",X"EE",X"D7",X"EE",X"76",X"F1",X"1D",X"F0",
		X"BC",X"E0",X"10",X"F1",X"1D",X"F0",X"5B",X"EB",X"CF",X"EF",X"FA",X"EC",X"30",X"F1",X"1D",X"E3",
		X"DA",X"D6",X"36",X"D6",X"97",X"D1",X"49",X"D3",X"8F",X"D0",X"87",X"D2",X"0B",X"D2",X"6C",X"CF",
		X"C5",X"D2",X"CD",X"D3",X"8F",X"D0",X"E8",X"D7",X"59",X"E0",X"D2",X"EF",X"FA",X"E0",X"10",X"F0",
		X"BC",X"E0",X"10",X"DA",X"00",X"EF",X"FA",X"E0",X"10",X"EF",X"FA",X"F0",X"BC",X"EF",X"FA",X"EE",
		X"15",X"ED",X"B4",X"F0",X"BC",X"F0",X"5B",X"EB",X"CF",X"F1",X"1D",X"E0",X"10",X"F1",X"7E",X"E3",
		X"18",X"F2",X"40",X"D3",X"F0",X"D2",X"CD",X"CF",X"C5",X"D2",X"6C",X"D0",X"E8",X"D1",X"AA",X"D3",
		X"8F",X"CF",X"C5",X"D2",X"6C",X"D0",X"87",X"D7",X"BA",X"E1",X"33",X"DB",X"E5",X"DB",X"84",X"DB",
		X"E5",X"F1",X"1D",X"DA",X"00",X"F0",X"BC",X"F1",X"1D",X"EE",X"15",X"ED",X"B4",X"F1",X"1D",X"E0",
		X"10",X"F1",X"1D",X"EF",X"FA",X"F0",X"BC",X"EB",X"CF",X"EF",X"FA",X"F0",X"5B",X"F1",X"1D",X"E5",
		X"BF",X"E5",X"5E",X"D6",X"36",X"D6",X"97",X"D3",X"2E",X"D1",X"49",X"D2",X"6C",X"CF",X"C5",X"CF",
		X"C5",X"D2",X"0B",X"CF",X"C5",X"D1",X"49",X"D8",X"DD",X"E2",X"56",X"EF",X"FA",X"F0",X"BC",X"D0",
		X"26",X"EF",X"FA",X"DA",X"00",X"D9",X"9F",X"D9",X"9F",X"D9",X"9F",X"D9",X"9F",X"D9",X"9F",X"D9",
		X"9F",X"D9",X"9F",X"D9",X"9F",X"DA",X"C2",X"EB",X"6E",X"D9",X"9F",X"DD",X"08",X"DD",X"69",X"DD",
		X"CA",X"E4",X"3B",X"F2",X"40",X"D5",X"13",X"D0",X"87",X"D3",X"8F",X"D0",X"E8",X"D0",X"87",X"D2",
		X"6C",X"D0",X"E8",X"D1",X"49",X"D8",X"1B",X"E1",X"94",X"F1",X"7E",X"DB",X"84",X"DC",X"46",X"D9",
		X"9F",X"D9",X"9F",X"DA",X"61",X"F1",X"DF",X"EF",X"FA",X"F1",X"7E",X"EF",X"FA",X"F0",X"BC",X"EF",
		X"38",X"F1",X"DF",X"DB",X"E5",X"DA",X"00",X"EB",X"CF",X"E0",X"10",X"DF",X"AF",X"E0",X"10",X"DE",
		X"2B",X"E3",X"18",X"F2",X"40",X"D3",X"F0",X"D0",X"E8",X"CF",X"C5",X"D1",X"AA",X"D3",X"8F",X"D0",
		X"87",X"CF",X"C5",X"D1",X"AA",X"D7",X"BA",X"E1",X"33",X"EF",X"FA",X"F0",X"5B",X"F1",X"DF",X"DB",
		X"84",X"F0",X"5B",X"D0",X"26",X"DB",X"84",X"EF",X"38",X"F1",X"DF",X"F0",X"5B",X"D0",X"26",X"F1",
		X"DF",X"F1",X"7E",X"EF",X"99",X"DA",X"00",X"EB",X"CF",X"F0",X"BC",X"DF",X"4E",X"DE",X"ED",X"DE",
		X"8C",X"E5",X"BF",X"E5",X"5E",X"D4",X"51",X"D1",X"49",X"F3",X"63",X"CF",X"C5",X"D1",X"49",X"D0",
		X"87",X"D2",X"0B",X"D0",X"87",X"D8",X"DD",X"E2",X"56",X"E0",X"10",X"F0",X"BC",X"DB",X"E5",X"D0",
		X"26",X"F1",X"DF",X"DB",X"84",X"F0",X"BC",X"F0",X"5B",X"DB",X"E5",X"F1",X"7E",X"DB",X"84",X"DB",
		X"E5",X"F0",X"5B",X"F0",X"BC",X"DA",X"00",X"EB",X"CF",X"EF",X"FA",X"F1",X"1D",X"EC",X"30",X"DA",
		X"00",X"EC",X"F2",X"E3",X"18",X"D6",X"36",X"D6",X"97",X"D1",X"49",X"D0",X"87",X"D0",X"E8",X"D2",
		X"6C",X"D0",X"E8",X"D8",X"1B",X"E1",X"94",X"F1",X"1D",X"F0",X"5B",X"F0",X"5B",X"DB",X"84",X"F1",
		X"7E",X"EF",X"38",X"F1",X"DF",X"DB",X"84",X"DB",X"E5",X"DB",X"84",X"F0",X"BC",X"DB",X"E5",X"DB",
		X"84",X"DB",X"E5",X"DB",X"84",X"DA",X"00",X"EB",X"CF",X"DB",X"84",X"F1",X"7E",X"F0",X"BC",X"DA",
		X"00",X"ED",X"53",X"E5",X"BF",X"E5",X"5E",X"D3",X"F0",X"CF",X"C5",X"D3",X"2E",X"D0",X"87",X"D1",
		X"AA",X"CF",X"C5",X"D7",X"59",X"E0",X"D2",X"E0",X"10",X"F1",X"7E",X"F0",X"5B",X"F0",X"BC",X"F1",
		X"1D",X"EF",X"FA",X"F1",X"1D",X"D9",X"9F",X"D9",X"9F",X"DA",X"C2",X"D9",X"9F",X"D9",X"9F",X"D9",
		X"9F",X"DA",X"C2",X"DC",X"A7",X"DA",X"00",X"EB",X"CF",X"F0",X"BC",X"DB",X"E5",X"DB",X"84",X"DA",
		X"00",X"E0",X"10",X"EC",X"91",X"E3",X"18",X"D6",X"36",X"D6",X"97",X"D2",X"6C",X"D0",X"E8",X"D1",
		X"49",X"D3",X"8F",X"D7",X"BA",X"E1",X"33",X"DC",X"46",X"D9",X"9F",X"D9",X"9F",X"D9",X"9F",X"D9",
		X"9F",X"DA",X"C2",X"D9",X"9F",X"D9",X"9F",X"D9",X"9F",X"DA",X"61",X"D9",X"9F",X"D9",X"9F",X"D9",
		X"9F",X"DA",X"61",X"D9",X"9F",X"DB",X"23",X"EB",X"6E",X"D9",X"9F",X"D9",X"9F",X"D9",X"9F",X"DB",
		X"23",X"D9",X"9F",X"DC",X"A7",X"E5",X"BF",X"E5",X"5E",X"D5",X"13",X"D0",X"87",X"D2",X"6C",X"D2",
		X"CD",X"D0",X"E8",X"D3",X"2E",X"D8",X"7C",X"E1",X"F5",X"DC",X"46",X"D9",X"9F",X"D9",X"9F",X"D9",
		X"9F",X"DB",X"23",X"D9",X"9F",X"DB",X"E5",X"DB",X"84",X"F0",X"BC",X"DB",X"E5",X"DB",X"84",X"DB",
		X"E5",X"DB",X"84",X"E0",X"10",X"DA",X"00",X"EB",X"CF",X"E8",X"05",X"E7",X"A4",X"F2",X"A1",X"F3",
		X"02",X"E7",X"43",X"E7",X"43",X"E7",X"43",X"E6",X"E2",X"D3",X"F0",X"D0",X"87",X"D3",X"2E",X"F3",
		X"63",X"CF",X"C5",X"CF",X"C5",X"D1",X"49",X"D8",X"7C",X"E1",X"F5",X"EF",X"FA",X"F1",X"1D",X"EF",
		X"FA",X"DA",X"00",X"DB",X"84",X"D9",X"9F",X"D9",X"9F",X"D9",X"9F",X"D9",X"9F",X"D9",X"9F",X"D9",
		X"9F",X"D9",X"9F",X"D9",X"9F",X"DA",X"61",X"EB",X"6E",X"D9",X"9F",X"DA",X"C2",X"D9",X"9F",X"DA",
		X"61",X"D9",X"9F",X"D9",X"9F",X"DC",X"A7",X"E4",X"3B",X"D6",X"36",X"D6",X"97",X"D0",X"E8",X"D1",
		X"49",X"D1",X"AA",X"D0",X"87",X"D2",X"6C",X"D9",X"3E",X"E2",X"B7",X"DC",X"46",X"D9",X"9F",X"D9",
		X"9F",X"DA",X"61",X"D9",X"9F",X"EF",X"FA",X"F1",X"1D",X"EF",X"FA",X"F1",X"1D",X"E0",X"10",X"F0",
		X"5B",X"F0",X"BC",X"F1",X"1D",X"EF",X"FA",X"EB",X"CF",X"F1",X"1D",X"DA",X"00",X"EC",X"30",X"E4",
		X"FD",X"E6",X"81",X"E6",X"81",X"E6",X"81",X"E4",X"9C",X"F2",X"40",X"D5",X"13",X"D2",X"0B",X"CF",
		X"C5",X"D0",X"E8",X"D1",X"49",X"D0",X"E8",X"D9",X"3E",X"E2",X"B7",X"E0",X"10",X"DB",X"E5",X"F1",
		X"1D",X"F0",X"BC",X"EF",X"FA",X"F0",X"BC",X"F1",X"1D",X"F0",X"5B",X"E0",X"10",X"E0",X"10",X"E0",
		X"10",X"D0",X"26",X"F0",X"5B",X"F0",X"5B",X"EB",X"CF",X"E0",X"10",X"DA",X"00",X"EF",X"FA",X"E5",
		X"BF",X"E6",X"20",X"E5",X"5E",X"F2",X"40",X"F2",X"40",X"F2",X"40",X"D3",X"F0",X"D1",X"49",X"CF",
		X"C5",X"D3",X"2E",X"D0",X"E8",X"D2",X"0B",X"D2",X"CD",X"D8",X"7C",X"E1",X"F5",X"EF",X"FA",X"EF",
		X"38",X"DB",X"84",X"F1",X"1D",X"D9",X"9F",X"D9",X"9F",X"D9",X"9F",X"DD",X"08",X"DD",X"69",X"DD",
		X"CA",X"DB",X"84",X"F0",X"BC",X"E0",X"10",X"EB",X"CF",X"F0",X"5B",X"DA",X"00",X"F1",X"1D",X"F0",
		X"5B",X"EC",X"F2",X"E3",X"18",X"F2",X"40",X"F2",X"40",X"F2",X"40",X"D4",X"51",X"D1",X"AA",X"D0",
		X"87",X"D1",X"49",X"D2",X"CD",X"D0",X"E8",X"D1",X"49",X"D8",X"1B",X"E1",X"94",X"DC",X"46",X"D9",
		X"9F",X"D9",X"9F",X"DA",X"C2",X"F0",X"5B",X"EF",X"38",X"F0",X"5B",X"DF",X"AF",X"E0",X"10",X"DE",
		X"2B",X"EF",X"FA",X"EF",X"38",X"DB",X"84",X"EB",X"CF",X"F0",X"5B",X"DA",X"00",X"D0",X"26",X"F0",
		X"BC",X"ED",X"53",X"E5",X"BF",X"E6",X"20",X"E5",X"5E",X"F2",X"40",X"D4",X"B2",X"D1",X"49",X"CF",
		X"C5",X"D0",X"87",X"D0",X"E8",X"D1",X"49",X"D0",X"E8",X"D7",X"BA",X"E1",X"33",X"DB",X"84",X"F0",
		X"BC",X"F1",X"1D",X"DA",X"00",X"F1",X"1D",X"F0",X"BC",X"EF",X"FA",X"DF",X"4E",X"DE",X"ED",X"DE",
		X"8C",X"F0",X"BC",X"DB",X"E5",X"F0",X"5B",X"EB",X"CF",X"F0",X"5B",X"DA",X"00",X"F1",X"1D",X"DB",
		X"84",X"DB",X"E5",X"EF",X"99",X"EC",X"91",X"E4",X"3B",X"D5",X"D5",X"D5",X"74",X"D0",X"E8",X"CF",
		X"C5",X"CF",X"C5",X"CF",X"C5",X"D0",X"E8",X"D0",X"87",X"D8",X"DD",X"E2",X"56",X"F0",X"BC",X"DB",
		X"84",X"DB",X"E5",X"DA",X"00",X"EF",X"FA",X"F1",X"1D",X"F1",X"1D",X"F0",X"5B",X"EF",X"FA",X"DA",
		X"00",X"EF",X"99",X"F0",X"BC",X"DB",X"E5",X"EB",X"CF",X"EF",X"38",X"DA",X"00",X"E0",X"10",X"DB",
		X"E5",X"DB",X"84",X"EC",X"F2",X"E4",X"FD",X"E4",X"9C",X"D4",X"B2",X"D2",X"CD",X"D1",X"49",X"CF",
		X"C5",X"D0",X"87",X"CF",X"C5",X"D0",X"87",X"D9",X"3E",X"E2",X"B7",X"DB",X"84",X"DB",X"E5",X"EF",
		X"99",X"DB",X"84",X"DA",X"00",X"F1",X"1D",X"DB",X"E5",X"F0",X"BC",X"EC",X"30",X"DB",X"84",X"DA",
		X"00",X"E0",X"10",X"D0",X"26",X"DB",X"84",X"EB",X"CF",X"F1",X"1D",X"DA",X"00",X"F0",X"BC",X"DB",
		X"84",X"DB",X"E5",X"ED",X"53",X"E3",X"79",X"D5",X"D5",X"D5",X"74",X"D0",X"E8",X"D0",X"87",X"D1",
		X"49",X"CF",X"C5",X"D1",X"AA",X"CF",X"C5",X"D8",X"DD",X"E2",X"56",X"EF",X"FA",X"F1",X"1D",X"DB",
		X"84",X"EF",X"99",X"DA",X"00",X"DB",X"84",X"EF",X"FA",X"EF",X"FA",X"DB",X"E5",X"F0",X"5B",X"DA",
		X"00",X"F0",X"5B",X"DB",X"84",X"DB",X"E5",X"EB",X"CF",X"DB",X"84",X"DA",X"00",X"E0",X"10",X"EF",
		X"FA",X"DB",X"84",X"EF",X"99",X"E3",X"DA",X"D4",X"B2",X"D1",X"49",X"CF",X"C5",X"D0",X"E8",X"D0",
		X"87",X"D1",X"49",X"D2",X"0B",X"D8",X"DD",X"E2",X"56",X"EF",X"FA",X"E0",X"10",X"F0",X"5B",X"EF",
		X"FA",X"E0",X"10",X"DA",X"00",X"E8",X"66",X"E8",X"66",X"E8",X"66",X"E8",X"66",X"E8",X"C7",X"E9",
		X"28",X"E8",X"66",X"E8",X"66",X"E8",X"66",X"E9",X"89",X"E8",X"C7",X"E9",X"28",X"E8",X"66",X"E8",
		X"66",X"E8",X"66",X"E8",X"66",X"EB",X"0D",X"EA",X"AC",X"EA",X"4B",X"EA",X"4B",X"EA",X"4B",X"EA",
		X"4B",X"EA",X"4B",X"EA",X"4B",X"E9",X"EA",X"E8",X"66",X"E8",X"66",X"E8",X"66",X"E8",X"66",X"E8",
		X"66",X"E8",X"C7",X"E9",X"28",X"E0",X"10",X"EF",X"FA",X"F0",X"5B",X"F0",X"BC",X"EF",X"FA",X"DA",
		X"00",X"EF",X"FA",X"EF",X"FA",X"E0",X"10",X"EB",X"CF",X"D0",X"26",X"DA",X"00",X"DB",X"E5",X"DB",
		X"84",X"DB",X"E5",X"EC",X"30",X"E4",X"3B",X"D5",X"13",X"CF",X"C5",X"D0",X"E8",X"D1",X"49",X"CF",
		X"C5",X"D0",X"87",X"D0",X"E8",X"D8",X"7C",X"E1",X"F5",X"DB",X"84",X"DB",X"E5",X"F0",X"BC",X"F1",
		X"1D",X"EF",X"FA",X"DA",X"00",X"F0",X"BC",X"EE",X"D7",X"EE",X"76",X"F1",X"1D",X"E0",X"10",X"DA",
		X"00",X"EE",X"15",X"ED",X"B4",X"F1",X"1D",X"EB",X"CF",X"E0",X"10",X"DA",X"00",X"DB",X"E5",X"F0",
		X"BC",X"DB",X"84",X"E4",X"FD",X"E4",X"9C",X"D5",X"13",X"D0",X"87",X"CF",X"C5",X"D1",X"49",X"D3",
		X"2E",X"CF",X"C5",X"D2",X"CD",X"D8",X"1B",X"E1",X"94",X"DB",X"E5",X"DB",X"84",X"DB",X"E5",X"F0",
		X"BC",X"F1",X"1D",X"DA",X"00",X"D9",X"9F",X"D9",X"9F",X"D9",X"9F",X"D9",X"9F",X"D9",X"9F",X"DB",
		X"23",X"D9",X"9F",X"D9",X"9F",X"D9",X"9F",X"EB",X"6E",X"D9",X"9F",X"DA",X"61",X"D9",X"9F",X"D9",
		X"9F",X"DC",X"A7",X"E3",X"DA",X"D5",X"D5",X"D5",X"74",X"D1",X"AA",X"D0",X"87",X"CF",X"C5",X"D0",
		X"E8",X"D0",X"87",X"D2",X"0B",X"D7",X"59",X"E0",X"D2",X"DC",X"46",X"D9",X"9F",X"D9",X"9F",X"D9",
		X"9F",X"DA",X"C2",X"DB",X"23",X"EF",X"FA",X"EE",X"15",X"EE",X"76",X"EF",X"FA",X"E0",X"10",X"DA",
		X"00",X"EE",X"D7",X"EE",X"76",X"E0",X"10",X"EB",X"CF",X"DB",X"84",X"F0",X"BC",X"DB",X"84",X"DB",
		X"E5",X"E4",X"FD",X"E4",X"9C",X"D4",X"B2",X"D0",X"87",X"CF",X"C5",X"D2",X"CD",X"D0",X"E8",X"D0",
		X"87",X"D2",X"6C",X"D1",X"49",X"D7",X"BA",X"E1",X"33",X"EF",X"FA",X"F1",X"1D",X"DB",X"84",X"DB",
		X"E5",X"DA",X"00",X"DA",X"00",X"F1",X"1D",X"F0",X"BC",X"F0",X"5B",X"F1",X"1D",X"F0",X"BC",X"DA",
		X"00",X"F1",X"1D",X"E0",X"10",X"EF",X"FA",X"EB",X"CF",X"F0",X"BC",X"DB",X"E5",X"F0",X"BC",X"EC",
		X"F2",X"E3",X"79",X"D5",X"D5",X"D5",X"74",X"D2",X"6C",X"D0",X"87",X"D1",X"49",X"D3",X"8F",X"D1",
		X"49",X"CF",X"C5",X"D0",X"E8",X"D2",X"0B",X"D8",X"7C",X"E1",X"F5",X"F0",X"BC",X"F1",X"1D",X"DB",
		X"84",X"DA",X"00",X"DA",X"00",X"D9",X"9F",X"D9",X"9F",X"D9",X"9F",X"D9",X"9F",X"D9",X"9F",X"DA",
		X"61",X"DC",X"A7",X"F1",X"1D",X"F0",X"BC",X"EB",X"CF",X"F1",X"1D",X"DB",X"84",X"DB",X"E5",X"ED",
		X"53",X"E3",X"79",X"D4",X"51",X"CF",X"C5",X"D1",X"AA",X"D0",X"E8",X"D2",X"6C",X"D0",X"87",X"D1",
		X"AA",X"F3",X"63",X"D1",X"49",X"D2",X"6C",X"D8",X"1B",X"E1",X"94",X"EF",X"FA",X"E0",X"10",X"DC",
		X"46",X"DA",X"61",X"DB",X"23",X"E0",X"10",X"E0",X"10",X"E0",X"10",X"E0",X"10",X"EF",X"FA",X"F1",
		X"1D",X"F0",X"5B",X"EF",X"FA",X"DB",X"E5",X"EB",X"CF",X"EF",X"FA",X"F0",X"BC",X"E0",X"10",X"F1",
		X"1D",X"E3",X"DA",X"D4",X"B2",X"D0",X"87",X"CF",X"C5",X"D3",X"8F",X"D1",X"49",X"D2",X"6C",X"D0",
		X"87",X"D2",X"6C",X"CF",X"C5",X"D2",X"CD",X"D7",X"BA",X"E1",X"33",X"DB",X"E5",X"EF",X"FA",X"E0",
		X"10",X"F1",X"1D",X"DA",X"00",X"E0",X"10",X"E0",X"10",X"E0",X"10",X"F0",X"BC",X"F1",X"1D",X"F0",
		X"5B",X"EE",X"D7",X"EE",X"76",X"DB",X"84",X"EB",X"CF",X"F1",X"1D",X"DB",X"E5",X"EF",X"FA",X"E4",
		X"FD",X"E4",X"9C",X"D5",X"13",X"D0",X"E8",X"D3",X"8F",X"D2",X"6C",X"D0",X"E8",X"D2",X"0B",X"CF",
		X"C5",X"D0",X"E8",X"D3",X"8F",X"D0",X"87",X"D8",X"DD",X"E2",X"56",X"DB",X"84",X"E0",X"10",X"F0",
		X"BC",X"EF",X"FA",X"DA",X"00",X"D9",X"9F",X"D9",X"9F",X"D9",X"9F",X"D9",X"9F",X"D9",X"9F",X"D9",
		X"9F",X"D9",X"9F",X"D9",X"9F",X"D9",X"9F",X"EB",X"6E",X"D9",X"9F",X"D9",X"9F",X"DC",X"A7",X"E3",
		X"79",X"D5",X"D5",X"D5",X"74",X"D2",X"6C",X"D0",X"87",X"D3",X"2E",X"D3",X"8F",X"D1",X"49",X"D2",
		X"6C",X"D1",X"AA",X"D0",X"E8",X"D1",X"49",X"D8",X"7C",X"E1",X"F5",X"DC",X"46",X"D9",X"9F",X"D9",
		X"9F",X"D9",X"9F",X"DB",X"23",X"F1",X"1D",X"E0",X"10",X"EE",X"D7",X"ED",X"B4",X"DB",X"84",X"DB",
		X"E5",X"DB",X"84",X"F0",X"BC",X"F1",X"1D",X"EB",X"CF",X"F0",X"5B",X"F0",X"BC",X"DB",X"84",X"E3",
		X"79",X"D4",X"B2",X"CF",X"C5",X"D0",X"E8",X"D1",X"AA",X"D0",X"E8",X"CF",X"C5",X"D0",X"87",X"CF",
		X"C5",X"D3",X"8F",X"D0",X"87",X"D2",X"6C",X"D9",X"3E",X"E2",X"B7",X"DB",X"E5",X"DB",X"84",X"F0",
		X"BC",X"E0",X"10",X"DA",X"00",X"0C",X"0D",X"0E",X"0F",X"1C",X"1D",X"1E",X"1F",X"1C",X"1D",X"1E",
		X"1F",X"0C",X"0D",X"0E",X"0F",X"1E",X"1F",X"0C",X"0D",X"0E",X"0F",X"1C",X"1D",X"0E",X"0F",X"1C",
		X"1D",X"1E",X"1F",X"0C",X"0D",X"0C",X"0D",X"0E",X"0F",X"1C",X"1D",X"1E",X"1F",X"1C",X"1D",X"1E",
		X"1F",X"0C",X"0D",X"0E",X"0F",X"1E",X"1E",X"0C",X"0D",X"0E",X"0F",X"1C",X"1D",X"0E",X"0F",X"1C",
		X"1D",X"1E",X"1F",X"0C",X"0D",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"10",X"21",
		X"22",X"21",X"22",X"21",X"22",X"12",X"32",X"8C",X"8D",X"8E",X"8F",X"AD",X"AE",X"30",X"60",X"65",
		X"65",X"65",X"65",X"65",X"65",X"61",X"32",X"BC",X"BD",X"BE",X"BF",X"30",X"51",X"51",X"00",X"01",
		X"01",X"01",X"02",X"00",X"01",X"02",X"30",X"49",X"49",X"49",X"32",X"30",X"49",X"32",X"10",X"21",
		X"21",X"21",X"12",X"10",X"21",X"12",X"10",X"33",X"33",X"33",X"33",X"36",X"66",X"66",X"63",X"30",
		X"00",X"00",X"03",X"44",X"44",X"44",X"44",X"30",X"00",X"03",X"33",X"33",X"33",X"33",X"33",X"3C",
		X"CC",X"33",X"C3",X"36",X"66",X"33",X"63",X"0C",X"0D",X"0E",X"0F",X"1C",X"1D",X"1E",X"1F",X"1C",
		X"1D",X"1E",X"1F",X"0C",X"43",X"0E",X"0F",X"1E",X"64",X"5A",X"0D",X"0E",X"0F",X"1C",X"1D",X"0E",
		X"74",X"6A",X"1D",X"1E",X"1F",X"0C",X"0D",X"0C",X"0D",X"0E",X"0F",X"1C",X"1D",X"1E",X"1F",X"1C",
		X"1D",X"1E",X"1F",X"0C",X"0D",X"4C",X"4D",X"1E",X"1F",X"0C",X"70",X"0E",X"0F",X"5C",X"5D",X"0E",
		X"0F",X"1C",X"1D",X"1E",X"0A",X"0C",X"0D",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"70",X"0E",X"0F",X"1C",X"1D",X"1E",X"1F",
		X"1C",X"1D",X"1E",X"1F",X"0C",X"0D",X"0E",X"0F",X"1E",X"1F",X"0C",X"0D",X"0E",X"0F",X"1C",X"EB",
		X"0E",X"0F",X"1C",X"1D",X"1E",X"1F",X"0C",X"0D",X"0C",X"0D",X"0E",X"0F",X"43",X"1D",X"1E",X"1F",
		X"1C",X"1D",X"1E",X"1F",X"0C",X"0D",X"0E",X"0F",X"1E",X"1F",X"0C",X"0D",X"0E",X"0F",X"1C",X"1D",
		X"0E",X"0F",X"1C",X"1D",X"1E",X"1F",X"0C",X"0D",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0D",X"0E",X"0F",X"1C",X"1D",X"1E",
		X"1F",X"1C",X"1D",X"6E",X"6F",X"0C",X"0D",X"0E",X"0F",X"1E",X"1F",X"7E",X"7F",X"0E",X"0F",X"1C",
		X"1D",X"0E",X"0F",X"1C",X"1D",X"1E",X"1F",X"0A",X"0D",X"0C",X"0D",X"0E",X"0F",X"1C",X"1D",X"1E",
		X"1F",X"1C",X"1D",X"1E",X"04",X"0C",X"0D",X"0E",X"0F",X"1E",X"1F",X"0C",X"69",X"2F",X"0F",X"1C",
		X"1D",X"0E",X"0F",X"1C",X"3F",X"4F",X"1F",X"0C",X"0D",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"8C",X"8D",X"8E",X"8F",X"9C",X"9D",
		X"9E",X"9A",X"9C",X"9D",X"9E",X"9F",X"8C",X"8D",X"8E",X"8F",X"9E",X"9F",X"8C",X"8D",X"8E",X"8F",
		X"9C",X"9D",X"8E",X"8F",X"C9",X"CA",X"CB",X"9F",X"8C",X"8D",X"8C",X"8D",X"DC",X"EA",X"ED",X"EE",
		X"9E",X"9F",X"9C",X"9D",X"EF",X"F6",X"F7",X"FF",X"8E",X"8F",X"9E",X"9F",X"8C",X"43",X"6F",X"7F",
		X"9C",X"9D",X"8E",X"8F",X"9C",X"9D",X"9E",X"9F",X"8C",X"8D",X"30",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"10",X"00",X"00",X"00",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0D",X"0E",X"40",X"41",
		X"42",X"1E",X"1F",X"1C",X"1D",X"1E",X"50",X"51",X"52",X"53",X"0F",X"1E",X"1F",X"0C",X"60",X"61",
		X"62",X"63",X"1D",X"0E",X"0F",X"1C",X"1D",X"71",X"72",X"73",X"0D",X"0C",X"0D",X"0E",X"0F",X"1C",
		X"1D",X"1E",X"1F",X"1C",X"1D",X"1E",X"1F",X"0C",X"0D",X"0E",X"0F",X"6C",X"6D",X"0C",X"0D",X"0E",
		X"0F",X"1C",X"1D",X"7C",X"7D",X"1C",X"1D",X"1E",X"1F",X"0C",X"0D",X"20",X"00",X"01",X"11",X"00",
		X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0D",X"0E",X"0F",
		X"1C",X"1D",X"1E",X"1F",X"1C",X"1D",X"1E",X"1F",X"0C",X"0D",X"0E",X"0F",X"1E",X"1F",X"0C",X"0D",
		X"00",X"01",X"02",X"03",X"40",X"41",X"42",X"1D",X"10",X"11",X"12",X"13",X"50",X"51",X"52",X"53",
		X"20",X"21",X"22",X"23",X"60",X"61",X"62",X"63",X"30",X"31",X"32",X"33",X"1E",X"71",X"72",X"73",
		X"0E",X"0F",X"1C",X"1D",X"A0",X"0F",X"1C",X"1D",X"1E",X"1F",X"0C",X"0D",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"10",X"11",X"10",X"10",X"00",X"10",X"00",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0D",X"0E",
		X"0F",X"1C",X"1D",X"1E",X"0A",X"1C",X"00",X"01",X"02",X"03",X"0D",X"0E",X"0F",X"1E",X"10",X"11",
		X"12",X"13",X"0F",X"1C",X"1D",X"0E",X"20",X"21",X"22",X"23",X"1F",X"0C",X"0D",X"0C",X"30",X"31",
		X"32",X"33",X"1D",X"1E",X"1F",X"1C",X"1D",X"1E",X"1F",X"0C",X"0D",X"0E",X"0F",X"1E",X"1F",X"0C",
		X"0D",X"0E",X"0F",X"6E",X"6F",X"0E",X"0F",X"1C",X"1D",X"1E",X"1F",X"7E",X"7F",X"20",X"00",X"00",
		X"00",X"00",X"01",X"11",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"8C",X"8D",
		X"8E",X"8F",X"9C",X"9D",X"9E",X"9F",X"9C",X"9D",X"99",X"9F",X"8C",X"8D",X"8E",X"8F",X"9E",X"9F",
		X"8C",X"8D",X"8E",X"8F",X"9C",X"9D",X"8E",X"8F",X"9C",X"9D",X"9E",X"9F",X"8C",X"8D",X"8C",X"8D",
		X"8E",X"85",X"86",X"87",X"88",X"9F",X"9C",X"98",X"9E",X"89",X"8A",X"A8",X"A9",X"8F",X"9E",X"9F",
		X"8C",X"AA",X"B8",X"B9",X"BA",X"9D",X"8E",X"8F",X"9C",X"C5",X"C6",X"C7",X"C8",X"8D",X"30",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"11",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",
		X"05",X"06",X"07",X"08",X"09",X"1E",X"1F",X"14",X"15",X"16",X"17",X"18",X"19",X"1A",X"0F",X"24",
		X"25",X"26",X"27",X"28",X"29",X"2A",X"2B",X"34",X"35",X"36",X"37",X"38",X"39",X"3A",X"3B",X"44",
		X"45",X"46",X"47",X"48",X"49",X"4A",X"4B",X"54",X"55",X"56",X"57",X"58",X"59",X"A8",X"5B",X"1E",
		X"65",X"66",X"67",X"68",X"A8",X"A8",X"6B",X"0E",X"75",X"76",X"77",X"78",X"79",X"7A",X"0D",X"20",
		X"00",X"11",X"00",X"00",X"01",X"11",X"10",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"03",X"30",X"00",X"00",X"00",X"00",
		X"FB",X"FB",X"FB",X"8C",X"8D",X"1D",X"1E",X"1F",X"FB",X"FB",X"FB",X"9C",X"9D",X"0D",X"0E",X"0F",
		X"FB",X"FB",X"FB",X"AC",X"AD",X"0F",X"1C",X"1D",X"FB",X"FB",X"FB",X"BC",X"BD",X"1F",X"0C",X"0D",
		X"FB",X"FB",X"FB",X"CC",X"CD",X"1D",X"1E",X"1F",X"FB",X"FB",X"FB",X"FB",X"DD",X"DE",X"DF",X"0F",
		X"FB",X"FB",X"FB",X"FB",X"FB",X"EE",X"EF",X"1D",X"FB",X"FB",X"FB",X"FB",X"FB",X"FE",X"FF",X"0D",
		X"20",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",
		X"00",X"22",X"22",X"20",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",
		X"00",X"FB",X"FB",X"FB",X"FB",X"FB",X"89",X"8A",X"1F",X"FB",X"FB",X"FB",X"FB",X"FB",X"99",X"9A",
		X"0F",X"FB",X"FB",X"FB",X"FB",X"FB",X"A9",X"AA",X"1D",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"BA",
		X"BB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"CA",X"CB",X"FB",X"FB",X"FB",X"FB",X"FB",X"D9",X"DA",
		X"DB",X"FB",X"FB",X"FB",X"FB",X"FB",X"E9",X"EA",X"1D",X"FB",X"FB",X"FB",X"FB",X"FB",X"F9",X"FA",
		X"0D",X"20",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"22",X"22",
		X"22",X"20",X"22",X"22",X"22",X"20",X"22",X"22",X"22",X"20",X"22",X"22",X"22",X"00",X"22",X"22",
		X"22",X"00",X"FB",X"FB",X"FB",X"FB",X"FB",X"84",X"85",X"1F",X"FB",X"FB",X"FB",X"FB",X"FB",X"94",
		X"95",X"0F",X"FB",X"FB",X"FB",X"FB",X"A3",X"A4",X"A5",X"1D",X"FB",X"FB",X"FB",X"FB",X"FB",X"B4",
		X"B5",X"0D",X"FB",X"FB",X"FB",X"FB",X"FB",X"C4",X"C5",X"1F",X"FB",X"FB",X"FB",X"FB",X"D3",X"D4",
		X"0E",X"0F",X"FB",X"FB",X"FB",X"E2",X"E3",X"E4",X"1C",X"1D",X"FB",X"FB",X"FB",X"F2",X"F3",X"1F",
		X"0C",X"0D",X"20",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"20",X"00",X"22",
		X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"20",X"00",X"22",X"22",X"00",X"00",X"22",
		X"22",X"00",X"00",X"FB",X"FB",X"FB",X"86",X"87",X"1D",X"1E",X"1F",X"FB",X"FB",X"FB",X"96",X"97",
		X"0D",X"0E",X"0F",X"FB",X"FB",X"FB",X"A6",X"A7",X"0F",X"1C",X"1D",X"FB",X"FB",X"FB",X"B6",X"B7",
		X"1F",X"0C",X"0D",X"FB",X"FB",X"FB",X"FB",X"C7",X"C8",X"1E",X"1F",X"FB",X"FB",X"FB",X"FB",X"D7",
		X"D8",X"0E",X"0F",X"FB",X"FB",X"FB",X"FB",X"E7",X"E8",X"1C",X"1D",X"FB",X"FB",X"FB",X"F6",X"F7",
		X"F8",X"0C",X"0D",X"20",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",
		X"22",X"22",X"00",X"00",X"22",X"22",X"20",X"00",X"22",X"22",X"20",X"00",X"22",X"22",X"20",X"00",
		X"22",X"22",X"00",X"00",X"FB",X"FB",X"FB",X"8E",X"8F",X"1D",X"1E",X"1F",X"FB",X"FB",X"FB",X"9E",
		X"9F",X"0D",X"0E",X"0F",X"FB",X"FB",X"FB",X"AE",X"AF",X"0F",X"1C",X"1D",X"FB",X"FB",X"FB",X"BE",
		X"BF",X"1F",X"0C",X"0D",X"80",X"81",X"82",X"CE",X"CF",X"1D",X"1E",X"1F",X"90",X"91",X"92",X"93",
		X"0C",X"0D",X"0E",X"0F",X"1E",X"1F",X"0C",X"0D",X"0E",X"0F",X"4C",X"4D",X"0E",X"0F",X"1C",X"1D",
		X"1E",X"1F",X"5C",X"5D",X"20",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",
		X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",
		X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",
		X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"B2",X"FB",X"FB",X"FB",
		X"FB",X"FB",X"FB",X"C1",X"C2",X"FB",X"FB",X"FB",X"FB",X"FB",X"D0",X"D1",X"D2",X"FB",X"FB",X"FB",
		X"FB",X"FB",X"E0",X"E1",X"0D",X"20",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"20",X"22",X"22",
		X"22",X"00",X"22",X"22",X"22",X"00",X"FB",X"FB",X"FB",X"FB",X"FB",X"DC",X"83",X"1F",X"FB",X"FB",
		X"FB",X"FB",X"FB",X"EC",X"ED",X"0F",X"FB",X"FB",X"FB",X"FB",X"FB",X"FC",X"FD",X"1D",X"FB",X"FB",
		X"FB",X"FB",X"FB",X"FB",X"A1",X"A2",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",
		X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",
		X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"20",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"22",
		X"22",X"22",X"00",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"0C",X"0D",X"0E",X"0A",X"1C",X"1D",X"1E",X"1F",X"1C",
		X"1D",X"1E",X"1F",X"0C",X"0D",X"0E",X"0F",X"B0",X"B1",X"0C",X"0D",X"0E",X"0F",X"1C",X"1D",X"C0",
		X"F0",X"F1",X"C6",X"8B",X"1F",X"43",X"0D",X"FB",X"FB",X"FB",X"D6",X"9B",X"1D",X"1E",X"1F",X"FB",
		X"FB",X"FB",X"E6",X"AB",X"0D",X"0E",X"0F",X"FB",X"FB",X"FB",X"D5",X"B9",X"0F",X"1C",X"04",X"FB",
		X"FB",X"FB",X"E5",X"C9",X"1F",X"0C",X"0D",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",
		X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"0C",X"0D",X"0E",X"0F",X"0B",X"B3",X"7B",X"A8",
		X"1C",X"1D",X"1E",X"1F",X"1B",X"B3",X"A8",X"A8",X"1E",X"4C",X"4D",X"0D",X"0E",X"2C",X"2D",X"B3",
		X"0E",X"5C",X"5D",X"1D",X"7B",X"1F",X"0C",X"0B",X"0C",X"0D",X"0E",X"0F",X"1C",X"1D",X"1E",X"1B",
		X"1C",X"1D",X"1E",X"1F",X"0C",X"04",X"0E",X"0B",X"1E",X"1F",X"0C",X"0D",X"0E",X"0F",X"1C",X"1B",
		X"0E",X"0F",X"1C",X"7B",X"1E",X"2C",X"2D",X"B3",X"20",X"00",X"00",X"45",X"74",X"00",X"00",X"45",
		X"44",X"00",X"00",X"04",X"45",X"00",X"00",X"70",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",
		X"04",X"00",X"00",X"00",X"04",X"00",X"07",X"04",X"45",X"0C",X"0D",X"0E",X"0F",X"0B",X"B3",X"7B",
		X"A8",X"1C",X"1D",X"70",X"1F",X"1B",X"B3",X"A8",X"3C",X"1E",X"1F",X"0C",X"0D",X"0B",X"B3",X"A8",
		X"4E",X"0E",X"7B",X"1C",X"1D",X"1B",X"B3",X"A8",X"4E",X"0C",X"0D",X"2C",X"2D",X"B3",X"A8",X"7B",
		X"4E",X"1C",X"0B",X"B3",X"A8",X"A8",X"3C",X"3D",X"3E",X"1E",X"1B",X"B3",X"A8",X"A8",X"5E",X"5F",
		X"5F",X"7B",X"0F",X"2C",X"2D",X"B3",X"A8",X"A8",X"A8",X"20",X"00",X"00",X"45",X"74",X"00",X"00",
		X"45",X"44",X"00",X"00",X"45",X"44",X"07",X"00",X"45",X"44",X"00",X"44",X"54",X"74",X"04",X"54",
		X"44",X"44",X"04",X"54",X"44",X"44",X"70",X"44",X"54",X"44",X"0C",X"0D",X"0E",X"0F",X"0B",X"B3",
		X"A8",X"A8",X"1C",X"1D",X"1E",X"1F",X"1B",X"B3",X"A8",X"3C",X"1E",X"1F",X"0C",X"0D",X"0E",X"0B",
		X"B3",X"5E",X"0E",X"0F",X"1C",X"7B",X"1E",X"1B",X"B3",X"A8",X"0C",X"04",X"0E",X"0F",X"1C",X"1D",
		X"0B",X"B3",X"1C",X"1D",X"1E",X"1F",X"43",X"0D",X"1B",X"B3",X"1E",X"1F",X"0C",X"0D",X"0E",X"0F",
		X"1C",X"0B",X"0E",X"0F",X"1C",X"1D",X"1E",X"7B",X"0C",X"1B",X"20",X"00",X"00",X"45",X"44",X"00",
		X"00",X"45",X"44",X"00",X"00",X"04",X"54",X"00",X"07",X"04",X"54",X"00",X"00",X"00",X"45",X"00",
		X"00",X"00",X"45",X"00",X"00",X"00",X"04",X"00",X"00",X"07",X"04",X"0C",X"64",X"5A",X"0F",X"1C",
		X"1D",X"1E",X"0B",X"1C",X"74",X"6A",X"1F",X"0C",X"0D",X"0E",X"1B",X"1E",X"1F",X"0C",X"0D",X"0E",
		X"2C",X"2D",X"B3",X"0E",X"7B",X"1C",X"2C",X"2D",X"B3",X"A8",X"A8",X"0C",X"0D",X"0B",X"B3",X"A8",
		X"7B",X"A8",X"3C",X"1C",X"1D",X"1B",X"B3",X"A8",X"A8",X"3C",X"3E",X"1E",X"1F",X"0C",X"0B",X"B3",
		X"A8",X"5E",X"5F",X"0E",X"7B",X"1C",X"1B",X"B3",X"A8",X"A8",X"A8",X"20",X"00",X"00",X"00",X"04",
		X"00",X"00",X"00",X"04",X"00",X"00",X"04",X"45",X"07",X"04",X"45",X"44",X"00",X"45",X"47",X"44",
		X"00",X"45",X"44",X"44",X"00",X"04",X"54",X"44",X"07",X"04",X"54",X"44",X"0B",X"B3",X"5E",X"5F",
		X"5F",X"5F",X"5F",X"2E",X"1B",X"B3",X"A8",X"A8",X"A8",X"A8",X"A8",X"5E",X"1E",X"2C",X"2D",X"2C",
		X"2D",X"B3",X"A8",X"A8",X"0E",X"0F",X"1C",X"1D",X"1E",X"2C",X"2D",X"B3",X"0C",X"0D",X"0E",X"7B",
		X"1C",X"1D",X"1E",X"0B",X"6C",X"6D",X"1E",X"1F",X"0C",X"0D",X"0E",X"1B",X"7C",X"7D",X"0C",X"0D",
		X"0E",X"0F",X"1C",X"0B",X"0E",X"0F",X"1C",X"1D",X"1E",X"7B",X"0C",X"1B",X"20",X"45",X"44",X"44",
		X"44",X"45",X"44",X"44",X"44",X"04",X"44",X"45",X"44",X"00",X"00",X"04",X"45",X"00",X"07",X"00",
		X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"07",X"04",X"0C",X"0D",X"0E",
		X"04",X"1C",X"1D",X"0B",X"7B",X"1C",X"1D",X"1E",X"1F",X"0C",X"0D",X"1B",X"B3",X"70",X"1F",X"0C",
		X"0D",X"2C",X"2D",X"B3",X"A8",X"0E",X"7B",X"1C",X"0B",X"B3",X"A8",X"A8",X"A8",X"0C",X"0D",X"0E",
		X"1B",X"B3",X"7B",X"3C",X"3D",X"1C",X"2C",X"2D",X"B3",X"A8",X"A8",X"4E",X"FB",X"0B",X"B3",X"A8",
		X"A8",X"A8",X"3C",X"3E",X"FB",X"1B",X"B3",X"3C",X"3D",X"3D",X"3E",X"FB",X"FB",X"20",X"00",X"00",
		X"00",X"47",X"00",X"00",X"00",X"45",X"00",X"00",X"44",X"54",X"07",X"04",X"54",X"44",X"00",X"04",
		X"57",X"44",X"04",X"45",X"44",X"44",X"45",X"44",X"44",X"44",X"45",X"44",X"44",X"44",X"0C",X"0D",
		X"0E",X"0F",X"1C",X"1D",X"1E",X"0B",X"1C",X"1D",X"1E",X"0A",X"0C",X"0D",X"0E",X"1B",X"1E",X"1F",
		X"0C",X"0D",X"0E",X"2C",X"2D",X"B3",X"0E",X"0F",X"7B",X"1D",X"0B",X"B3",X"A8",X"A8",X"0C",X"0D",
		X"0E",X"0F",X"1B",X"B3",X"A8",X"7B",X"1C",X"4C",X"4D",X"1F",X"0C",X"2C",X"2D",X"B3",X"1E",X"5C",
		X"5D",X"0D",X"0E",X"0F",X"1C",X"0B",X"0E",X"0F",X"1C",X"1D",X"1E",X"7B",X"0C",X"1B",X"20",X"00",
		X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"04",X"45",X"00",X"70",X"45",X"44",X"00",
		X"00",X"45",X"47",X"00",X"00",X"04",X"45",X"00",X"00",X"00",X"04",X"00",X"00",X"07",X"04",X"19",
		X"81",X"82",X"19",X"19",X"81",X"82",X"19",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",
		X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"92",X"92",X"C4",X"C5",X"92",X"92",X"C4",X"C5",X"51",
		X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"62",X"00",X"01",X"01",X"01",X"01",X"02",X"62",X"64",
		X"30",X"51",X"51",X"51",X"51",X"32",X"64",X"72",X"10",X"22",X"22",X"22",X"22",X"12",X"72",X"10",
		X"39",X"93",X"39",X"93",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"AA",X"33",X"AA",
		X"33",X"33",X"33",X"33",X"43",X"33",X"33",X"34",X"43",X"33",X"33",X"34",X"43",X"66",X"66",X"34",
		X"17",X"51",X"51",X"A1",X"51",X"00",X"01",X"02",X"A3",X"51",X"51",X"B1",X"51",X"30",X"51",X"32",
		X"B3",X"51",X"51",X"94",X"51",X"10",X"11",X"12",X"17",X"51",X"51",X"94",X"51",X"60",X"65",X"61",
		X"17",X"51",X"51",X"A1",X"51",X"00",X"01",X"02",X"A3",X"51",X"51",X"B1",X"51",X"30",X"51",X"43",
		X"B3",X"51",X"51",X"94",X"51",X"30",X"51",X"43",X"17",X"51",X"51",X"94",X"51",X"10",X"22",X"12",
		X"10",X"33",X"3A",X"33",X"33",X"93",X"3A",X"33",X"33",X"93",X"33",X"33",X"33",X"33",X"33",X"34",
		X"44",X"33",X"3A",X"33",X"33",X"93",X"3A",X"33",X"36",X"93",X"33",X"33",X"36",X"33",X"33",X"33",
		X"63",X"A0",X"51",X"51",X"A4",X"19",X"81",X"82",X"19",X"51",X"51",X"51",X"51",X"51",X"51",X"51",
		X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"92",X"92",X"C4",X"C5",X"92",X"92",X"C4",
		X"C5",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"34",X"35",X"35",X"36",X"51",
		X"51",X"51",X"51",X"44",X"51",X"51",X"46",X"51",X"51",X"51",X"51",X"54",X"55",X"55",X"56",X"51",
		X"51",X"10",X"33",X"33",X"39",X"93",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"AA",
		X"33",X"AA",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"33",X"33",X"19",X"81",X"82",X"19",X"19",X"81",X"82",X"19",X"51",X"51",X"51",X"51",X"51",X"51",
		X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"93",X"51",X"51",X"91",X"92",X"92",
		X"C4",X"C5",X"17",X"51",X"51",X"A1",X"51",X"51",X"51",X"51",X"A3",X"51",X"51",X"B1",X"34",X"35",
		X"36",X"51",X"B3",X"51",X"51",X"94",X"44",X"51",X"46",X"51",X"17",X"51",X"51",X"94",X"54",X"55",
		X"56",X"51",X"10",X"39",X"93",X"39",X"93",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"33",X"33",X"AA",X"33",X"3A",X"33",X"33",X"93",X"3A",X"33",X"33",X"93",X"33",X"33",X"33",X"33",
		X"33",X"33",X"33",X"A0",X"51",X"51",X"A4",X"19",X"81",X"82",X"19",X"51",X"51",X"51",X"51",X"51",
		X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"93",X"51",X"51",X"91",X"92",
		X"92",X"C4",X"C5",X"17",X"51",X"51",X"A1",X"51",X"51",X"51",X"51",X"A3",X"51",X"51",X"B1",X"51",
		X"34",X"35",X"36",X"B3",X"51",X"51",X"94",X"51",X"44",X"51",X"46",X"17",X"51",X"51",X"94",X"51",
		X"54",X"55",X"56",X"10",X"33",X"33",X"39",X"93",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"33",X"33",X"33",X"AA",X"33",X"3A",X"33",X"33",X"93",X"3A",X"33",X"33",X"93",X"33",X"33",X"33",
		X"33",X"33",X"33",X"33",X"51",X"51",X"51",X"51",X"51",X"51",X"EC",X"51",X"00",X"01",X"01",X"01",
		X"01",X"02",X"EC",X"51",X"10",X"22",X"22",X"22",X"22",X"12",X"EC",X"51",X"51",X"51",X"51",X"51",
		X"51",X"51",X"51",X"51",X"51",X"50",X"51",X"50",X"51",X"50",X"51",X"51",X"51",X"51",X"00",X"01",
		X"01",X"01",X"01",X"02",X"51",X"51",X"10",X"22",X"22",X"22",X"22",X"12",X"51",X"49",X"49",X"49",
		X"49",X"49",X"49",X"49",X"10",X"33",X"33",X"33",X"C3",X"33",X"33",X"33",X"C3",X"36",X"66",X"66",
		X"C3",X"33",X"33",X"33",X"33",X"39",X"39",X"39",X"33",X"33",X"33",X"33",X"33",X"33",X"36",X"66",
		X"63",X"3C",X"CC",X"CC",X"CC",X"51",X"51",X"51",X"51",X"51",X"00",X"01",X"02",X"00",X"01",X"02",
		X"51",X"50",X"30",X"51",X"43",X"30",X"50",X"43",X"51",X"51",X"30",X"51",X"43",X"30",X"51",X"43",
		X"51",X"50",X"30",X"51",X"43",X"30",X"50",X"43",X"51",X"51",X"30",X"51",X"43",X"30",X"51",X"43",
		X"51",X"50",X"30",X"51",X"43",X"30",X"50",X"43",X"51",X"51",X"10",X"11",X"12",X"10",X"11",X"12",
		X"51",X"51",X"51",X"51",X"51",X"10",X"33",X"33",X"33",X"33",X"33",X"33",X"93",X"36",X"39",X"63",
		X"33",X"36",X"33",X"63",X"93",X"36",X"39",X"63",X"33",X"36",X"33",X"63",X"93",X"36",X"39",X"63",
		X"33",X"33",X"33",X"33",X"33",X"33",X"51",X"04",X"05",X"05",X"06",X"80",X"19",X"19",X"51",X"14",
		X"15",X"15",X"16",X"17",X"A2",X"51",X"51",X"14",X"15",X"15",X"16",X"17",X"A2",X"51",X"51",X"24",
		X"25",X"25",X"26",X"C3",X"92",X"92",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"00",X"01",
		X"01",X"02",X"00",X"01",X"01",X"02",X"30",X"51",X"51",X"32",X"30",X"51",X"51",X"32",X"10",X"11",
		X"11",X"12",X"10",X"11",X"11",X"12",X"10",X"35",X"55",X"33",X"33",X"35",X"55",X"33",X"43",X"35",
		X"55",X"33",X"43",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"19",X"19",X"84",X"51",X"04",X"05",X"05",X"06",X"51",
		X"A2",X"94",X"51",X"14",X"15",X"15",X"16",X"51",X"A2",X"94",X"51",X"14",X"15",X"15",X"16",X"92",
		X"92",X"C1",X"51",X"24",X"25",X"25",X"26",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"00",
		X"01",X"01",X"02",X"00",X"01",X"01",X"02",X"30",X"51",X"51",X"32",X"30",X"51",X"51",X"32",X"10",
		X"11",X"11",X"12",X"10",X"11",X"11",X"12",X"10",X"33",X"33",X"55",X"53",X"34",X"33",X"55",X"53",
		X"34",X"33",X"55",X"53",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"19",X"81",X"82",X"19",X"19",X"81",X"82",X"19",
		X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",
		X"93",X"51",X"51",X"91",X"92",X"92",X"C4",X"C5",X"17",X"51",X"51",X"A1",X"51",X"51",X"51",X"51",
		X"A3",X"51",X"51",X"B1",X"51",X"91",X"92",X"92",X"B3",X"51",X"51",X"94",X"51",X"94",X"68",X"69",
		X"17",X"51",X"51",X"94",X"51",X"94",X"78",X"79",X"10",X"39",X"93",X"39",X"93",X"33",X"33",X"33",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"AA",X"33",X"3A",X"33",X"33",X"93",X"3A",X"33",
		X"33",X"93",X"33",X"33",X"74",X"33",X"33",X"33",X"43",X"19",X"81",X"82",X"19",X"19",X"81",X"82",
		X"19",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",
		X"51",X"92",X"92",X"C4",X"C5",X"92",X"92",X"C4",X"C5",X"51",X"51",X"51",X"51",X"51",X"51",X"51",
		X"51",X"92",X"92",X"92",X"92",X"92",X"92",X"92",X"92",X"68",X"69",X"68",X"69",X"68",X"69",X"68",
		X"69",X"78",X"79",X"78",X"79",X"78",X"79",X"78",X"79",X"10",X"39",X"93",X"39",X"93",X"33",X"33",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"AA",X"33",X"AA",X"33",X"33",X"33",X"33",X"33",X"33",
		X"33",X"33",X"74",X"74",X"74",X"74",X"43",X"43",X"43",X"43",X"19",X"81",X"82",X"19",X"19",X"81",
		X"82",X"84",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"94",X"51",X"51",X"51",X"51",X"51",X"51",
		X"51",X"94",X"92",X"92",X"C4",X"C5",X"93",X"51",X"51",X"94",X"51",X"51",X"51",X"51",X"17",X"51",
		X"51",X"A1",X"92",X"92",X"93",X"51",X"A3",X"51",X"51",X"B1",X"68",X"69",X"17",X"51",X"B3",X"51",
		X"51",X"94",X"78",X"79",X"17",X"51",X"17",X"51",X"51",X"94",X"10",X"39",X"93",X"39",X"93",X"33",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"AA",X"33",X"33",X"33",X"33",X"33",X"3A",X"33",
		X"33",X"93",X"3A",X"74",X"33",X"93",X"33",X"43",X"33",X"33",X"33",X"68",X"69",X"17",X"51",X"17",
		X"51",X"51",X"A1",X"78",X"79",X"17",X"51",X"A3",X"51",X"51",X"B1",X"68",X"69",X"17",X"51",X"B3",
		X"51",X"51",X"94",X"78",X"79",X"17",X"51",X"17",X"51",X"51",X"94",X"68",X"69",X"17",X"51",X"17",
		X"51",X"51",X"A1",X"78",X"79",X"17",X"51",X"A3",X"51",X"51",X"B1",X"68",X"69",X"17",X"51",X"B3",
		X"51",X"51",X"94",X"78",X"79",X"17",X"51",X"17",X"51",X"51",X"94",X"10",X"74",X"33",X"33",X"3A",
		X"43",X"33",X"93",X"3A",X"74",X"33",X"93",X"33",X"43",X"33",X"33",X"33",X"74",X"33",X"33",X"3A",
		X"43",X"33",X"93",X"3A",X"74",X"33",X"93",X"33",X"43",X"33",X"33",X"33",X"68",X"69",X"17",X"51",
		X"17",X"51",X"51",X"A1",X"78",X"79",X"17",X"51",X"A3",X"51",X"51",X"B1",X"19",X"19",X"A0",X"51",
		X"B3",X"51",X"51",X"94",X"51",X"51",X"51",X"51",X"17",X"51",X"51",X"94",X"19",X"81",X"82",X"19",
		X"A0",X"51",X"51",X"A1",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"B1",X"51",X"51",X"51",X"51",
		X"51",X"51",X"51",X"94",X"93",X"51",X"51",X"91",X"92",X"92",X"92",X"C1",X"10",X"74",X"33",X"33",
		X"3A",X"43",X"33",X"93",X"3A",X"33",X"33",X"93",X"33",X"33",X"33",X"33",X"33",X"39",X"93",X"33",
		X"3A",X"33",X"33",X"33",X"3A",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"68",X"69",X"68",
		X"69",X"68",X"69",X"68",X"69",X"78",X"79",X"78",X"79",X"78",X"79",X"78",X"79",X"19",X"19",X"19",
		X"19",X"19",X"19",X"19",X"19",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"19",X"81",X"82",
		X"19",X"19",X"81",X"82",X"19",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"51",
		X"51",X"51",X"51",X"51",X"51",X"92",X"92",X"C4",X"C5",X"92",X"92",X"C4",X"C5",X"10",X"74",X"74",
		X"74",X"74",X"43",X"43",X"43",X"43",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"39",X"93",
		X"39",X"93",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"AA",X"33",X"AA",X"17",X"51",
		X"51",X"A1",X"51",X"94",X"68",X"69",X"A3",X"51",X"51",X"B1",X"51",X"94",X"78",X"79",X"B3",X"51",
		X"51",X"94",X"51",X"A4",X"19",X"19",X"17",X"51",X"51",X"94",X"51",X"51",X"51",X"51",X"17",X"51",
		X"51",X"A4",X"19",X"81",X"82",X"19",X"A3",X"51",X"51",X"51",X"51",X"51",X"51",X"51",X"B3",X"51",
		X"51",X"51",X"51",X"51",X"51",X"51",X"C3",X"92",X"C4",X"C5",X"92",X"92",X"C4",X"C5",X"10",X"33",
		X"3A",X"33",X"74",X"93",X"3A",X"33",X"43",X"93",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"33",X"39",X"93",X"93",X"33",X"33",X"33",X"93",X"33",X"33",X"33",X"33",X"AA",X"33",X"AA",X"17",
		X"51",X"51",X"A1",X"51",X"94",X"68",X"69",X"A3",X"51",X"51",X"B1",X"51",X"94",X"78",X"79",X"B3",
		X"51",X"51",X"94",X"51",X"94",X"68",X"69",X"17",X"51",X"51",X"94",X"51",X"94",X"78",X"79",X"17",
		X"51",X"51",X"A1",X"51",X"94",X"68",X"69",X"A3",X"51",X"51",X"B1",X"51",X"94",X"78",X"79",X"B3",
		X"51",X"51",X"94",X"51",X"94",X"68",X"69",X"17",X"51",X"51",X"94",X"51",X"94",X"78",X"79",X"10",
		X"33",X"3A",X"33",X"74",X"93",X"3A",X"33",X"43",X"93",X"33",X"33",X"74",X"33",X"33",X"33",X"43");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
