library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity bagman_tile_bit1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of bagman_tile_bit1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",X"00",X"02",X"02",X"FE",X"FE",X"42",X"02",X"00",X"00",
		X"62",X"F2",X"BA",X"9A",X"9E",X"CE",X"46",X"00",X"8C",X"DE",X"F2",X"B2",X"92",X"86",X"04",X"00",
		X"08",X"FE",X"FE",X"C8",X"68",X"38",X"18",X"00",X"1C",X"BE",X"A2",X"A2",X"A2",X"E6",X"E4",X"00",
		X"0C",X"9E",X"92",X"92",X"D2",X"7E",X"3C",X"00",X"C0",X"E0",X"B0",X"9E",X"8E",X"C0",X"C0",X"00",
		X"0C",X"6E",X"9A",X"9A",X"B2",X"F2",X"6C",X"00",X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"18",X"24",X"62",X"51",X"85",X"46",X"24",X"18",X"18",X"24",X"46",X"89",X"91",X"62",X"24",X"18",
		X"18",X"24",X"42",X"D5",X"AB",X"42",X"24",X"18",X"00",X"00",X"80",X"80",X"80",X"80",X"FF",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",
		X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",X"44",X"C6",X"82",X"82",X"C6",X"7C",X"38",X"00",
		X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",X"82",X"92",X"92",X"92",X"FE",X"FE",X"00",X"00",
		X"80",X"90",X"90",X"90",X"90",X"FE",X"FE",X"00",X"9E",X"9E",X"92",X"82",X"C6",X"7C",X"38",X"00",
		X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",X"82",X"82",X"FE",X"FE",X"82",X"82",X"00",X"00",
		X"FC",X"FE",X"02",X"02",X"02",X"06",X"04",X"00",X"82",X"C6",X"6E",X"3C",X"18",X"FE",X"FE",X"00",
		X"02",X"02",X"02",X"02",X"FE",X"FE",X"00",X"00",X"FE",X"FE",X"70",X"38",X"70",X"FE",X"FE",X"00",
		X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",X"00",
		X"70",X"F8",X"88",X"88",X"88",X"FE",X"FE",X"00",X"7A",X"FC",X"8E",X"8A",X"82",X"FE",X"7C",X"00",
		X"72",X"F6",X"9E",X"8C",X"88",X"FE",X"FE",X"00",X"0C",X"5E",X"D2",X"92",X"92",X"F6",X"64",X"00",
		X"80",X"80",X"FE",X"FE",X"80",X"80",X"00",X"00",X"FC",X"FE",X"02",X"02",X"02",X"FE",X"FC",X"00",
		X"F0",X"F8",X"1C",X"0E",X"1C",X"F8",X"F0",X"00",X"F8",X"FE",X"1C",X"38",X"1C",X"FE",X"F8",X"00",
		X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",X"C0",X"F0",X"1E",X"1E",X"F0",X"C0",X"00",X"00",
		X"C2",X"E2",X"F2",X"BA",X"9E",X"8E",X"86",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",
		X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"00",X"40",X"40",X"40",X"40",X"40",X"40",X"00",
		X"00",X"00",X"00",X"00",X"28",X"00",X"00",X"00",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"00",X"00",X"82",X"C6",X"6C",X"38",X"00",X"00",X"00",X"00",X"38",X"6C",X"C6",X"82",X"00",X"00",
		X"00",X"00",X"82",X"FE",X"FE",X"82",X"00",X"00",X"82",X"FE",X"FE",X"82",X"82",X"FE",X"FE",X"82",
		X"00",X"28",X"28",X"28",X"28",X"28",X"28",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"00",
		X"F6",X"F6",X"00",X"00",X"F6",X"F6",X"00",X"00",X"FA",X"FA",X"00",X"00",X"FA",X"FA",X"00",X"00",
		X"00",X"00",X"00",X"F6",X"F6",X"00",X"00",X"00",X"00",X"00",X"00",X"FA",X"FA",X"00",X"00",X"00",
		X"00",X"00",X"00",X"E0",X"C0",X"00",X"00",X"00",X"00",X"E0",X"C0",X"00",X"E0",X"C0",X"00",X"00",
		X"00",X"60",X"E0",X"00",X"60",X"E0",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"1F",X"20",X"40",X"80",X"80",X"80",X"80",X"80",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"40",X"20",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"36",X"00",X"00",X"00",X"09",X"3B",X"2B",X"2B",X"A8",
		X"7F",X"6B",X"62",X"46",X"00",X"07",X"06",X"00",X"A9",X"AB",X"AB",X"AB",X"80",X"80",X"00",X"00",
		X"00",X"00",X"C8",X"EA",X"02",X"42",X"62",X"60",X"00",X"00",X"00",X"20",X"A8",X"A8",X"A8",X"A0",
		X"60",X"62",X"42",X"02",X"02",X"00",X"00",X"00",X"A1",X"AB",X"AB",X"AA",X"A0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"36",X"7F",X"6B",X"00",X"00",X"00",X"09",X"3B",X"2B",X"AB",X"A8",
		X"62",X"46",X"01",X"07",X"07",X"03",X"00",X"00",X"A9",X"AB",X"AB",X"AB",X"80",X"80",X"00",X"00",
		X"00",X"10",X"38",X"10",X"00",X"40",X"02",X"07",X"D7",X"D0",X"D7",X"80",X"0F",X"20",X"3F",X"00",
		X"02",X"20",X"70",X"21",X"00",X"04",X"0E",X"04",X"07",X"0C",X"1F",X"39",X"2C",X"18",X"1F",X"0F",
		X"00",X"00",X"00",X"10",X"38",X"10",X"00",X"40",X"D7",X"D0",X"D7",X"80",X"0F",X"10",X"1F",X"00",
		X"04",X"0E",X"04",X"00",X"20",X"70",X"21",X"00",X"07",X"0C",X"1F",X"39",X"2C",X"18",X"1F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D7",X"D0",X"D7",X"80",X"0F",X"10",X"1F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"0C",X"1F",X"39",X"2C",X"18",X"1F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D7",X"D0",X"D7",X"80",X"0F",X"00",X"3F",X"D0",
		X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"FF",X"A0",X"AE",X"12",X"0A",X"0A",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"06",X"1F",X"00",X"00",X"00",X"11",X"17",X"97",X"07",X"05",
		X"1D",X"1D",X"01",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"D5",X"54",X"54",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"36",X"FF",X"00",X"00",X"00",X"00",X"09",X"2B",X"2B",X"AB",
		X"EA",X"EA",X"46",X"00",X"00",X"00",X"00",X"00",X"A8",X"A9",X"AB",X"AB",X"2B",X"00",X"00",X"00",
		X"00",X"03",X"01",X"00",X"01",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",X"80",
		X"0C",X"36",X"7F",X"6B",X"62",X"46",X"00",X"00",X"00",X"E0",X"00",X"C0",X"00",X"00",X"00",X"00",
		X"0F",X"07",X"00",X"07",X"00",X"0F",X"80",X"EF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"E8",X"1F",X"68",X"FF",X"D4",X"C7",X"8C",X"00",X"00",X"80",X"00",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"70",X"75",X"00",X"F0",X"70",X"00",X"70",X"40",X"40",X"41",
		X"05",X"1D",X"6D",X"FF",X"D5",X"C5",X"8C",X"00",X"57",X"57",X"56",X"40",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"18",X"6C",X"FE",X"00",X"00",X"78",X"B8",X"90",X"D0",X"50",X"50",
		X"D7",X"C5",X"8D",X"01",X"00",X"00",X"01",X"00",X"50",X"50",X"50",X"50",X"50",X"90",X"B8",X"3C",
		X"00",X"00",X"00",X"00",X"06",X"1B",X"3F",X"35",X"00",X"00",X"00",X"30",X"20",X"35",X"97",X"D7",
		X"31",X"23",X"00",X"00",X"00",X"00",X"00",X"00",X"53",X"50",X"50",X"54",X"54",X"54",X"DC",X"1E",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"36",X"7F",X"00",X"00",X"3C",X"DC",X"88",X"88",X"88",X"A8",
		X"6B",X"62",X"46",X"00",X"00",X"00",X"00",X"00",X"A8",X"A8",X"A8",X"A9",X"2F",X"2F",X"66",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"36",X"7F",X"00",X"00",X"00",X"00",X"09",X"2B",X"3B",X"AB",
		X"6B",X"62",X"46",X"00",X"00",X"00",X"00",X"00",X"A8",X"A9",X"AB",X"AB",X"2B",X"00",X"00",X"00",
		X"00",X"10",X"38",X"10",X"00",X"40",X"02",X"07",X"C0",X"C0",X"C0",X"80",X"00",X"3F",X"3F",X"0F",
		X"02",X"20",X"70",X"21",X"00",X"04",X"0E",X"04",X"07",X"0F",X"1F",X"7F",X"2F",X"1F",X"00",X"00",
		X"00",X"00",X"00",X"10",X"38",X"10",X"00",X"40",X"C0",X"C0",X"C0",X"80",X"00",X"1F",X"1F",X"0F",
		X"04",X"0E",X"04",X"00",X"20",X"70",X"21",X"00",X"07",X"0F",X"1F",X"7F",X"2F",X"1F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"80",X"00",X"1F",X"1F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"0F",X"1F",X"7F",X"2F",X"1F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"80",X"00",X"10",X"38",X"5C",
		X"02",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"7C",X"FC",X"FE",X"FF",X"FF",X"3F",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"13",X"00",X"00",X"00",X"01",X"03",X"23",X"F3",X"F0",
		X"1F",X"1F",X"07",X"07",X"01",X"00",X"00",X"00",X"F0",X"F8",X"FC",X"FC",X"FC",X"5C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"0C",X"16",X"9F",X"00",X"00",X"00",X"00",X"01",X"23",X"63",X"E3",
		X"FF",X"FF",X"3F",X"3E",X"0E",X"02",X"00",X"00",X"E0",X"E1",X"E3",X"E3",X"63",X"00",X"00",X"00",
		X"00",X"00",X"DC",X"FF",X"1F",X"3D",X"1C",X"1E",X"00",X"00",X"00",X"00",X"08",X"88",X"88",X"00",
		X"1E",X"1C",X"3D",X"1B",X"03",X"01",X"00",X"00",X"01",X"83",X"83",X"82",X"C0",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"16",X"00",X"00",X"10",X"11",X"13",X"33",X"33",X"20",
		X"1F",X"1F",X"1F",X"3F",X"3E",X"0F",X"06",X"00",X"E1",X"F3",X"F3",X"E3",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"04",X"0C",X"16",X"1F",X"1F",X"00",X"00",X"10",X"11",X"13",X"73",X"F3",X"E0",
		X"10",X"3F",X"3E",X"0E",X"07",X"03",X"00",X"00",X"E1",X"F3",X"F3",X"E3",X"C0",X"80",X"00",X"00",
		X"08",X"04",X"02",X"01",X"04",X"0C",X"16",X"1F",X"00",X"00",X"00",X"80",X"C0",X"61",X"E3",X"E3",
		X"1F",X"1F",X"3F",X"3E",X"0E",X"02",X"00",X"00",X"C3",X"C0",X"E0",X"E1",X"67",X"07",X"06",X"00",
		X"00",X"00",X"00",X"1F",X"01",X"04",X"0C",X"16",X"00",X"00",X"00",X"80",X"80",X"C1",X"E3",X"E3",
		X"1F",X"1F",X"1F",X"3F",X"3E",X"0E",X"02",X"00",X"E3",X"C0",X"C0",X"E1",X"E7",X"67",X"06",X"00",
		X"08",X"04",X"02",X"01",X"00",X"04",X"0C",X"16",X"00",X"00",X"00",X"80",X"C0",X"41",X"63",X"E3",
		X"1F",X"1F",X"1F",X"3F",X"3E",X"0E",X"02",X"00",X"E3",X"C0",X"C0",X"E1",X"E7",X"67",X"06",X"00",
		X"00",X"00",X"00",X"00",X"04",X"0C",X"16",X"1F",X"20",X"20",X"20",X"60",X"60",X"41",X"E3",X"E3",
		X"1F",X"1F",X"3F",X"3E",X"0E",X"02",X"00",X"00",X"C3",X"C0",X"E0",X"E1",X"67",X"07",X"06",X"00",
		X"00",X"00",X"00",X"02",X"06",X"0B",X"0F",X"0F",X"10",X"10",X"10",X"30",X"30",X"21",X"B3",X"F3",
		X"0F",X"1F",X"1F",X"07",X"01",X"00",X"00",X"00",X"F3",X"E0",X"E0",X"60",X"60",X"40",X"DC",X"DE",
		X"00",X"00",X"00",X"00",X"04",X"0C",X"16",X"1F",X"00",X"80",X"BC",X"DC",X"C0",X"60",X"60",X"E0",
		X"1F",X"1F",X"3F",X"3E",X"0E",X"02",X"00",X"00",X"E0",X"E0",X"E0",X"60",X"40",X"DC",X"DE",X"DE",
		X"00",X"00",X"00",X"00",X"04",X"0C",X"16",X"1F",X"40",X"40",X"7C",X"DC",X"C0",X"80",X"C0",X"C0",
		X"1F",X"1F",X"3F",X"3E",X"0E",X"02",X"00",X"00",X"C0",X"C0",X"E0",X"E1",X"67",X"27",X"66",X"60",
		X"00",X"00",X"00",X"00",X"04",X"0C",X"16",X"1F",X"00",X"00",X"00",X"10",X"11",X"13",X"33",X"33",
		X"1F",X"1F",X"3F",X"3E",X"0E",X"02",X"00",X"00",X"E0",X"E1",X"F3",X"F3",X"63",X"00",X"00",X"00",
		X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"C0",X"20",X"20",X"C0",X"00",X"C0",X"20",X"20",
		X"00",X"00",X"0E",X"8C",X"CC",X"EA",X"00",X"00",X"01",X"01",X"00",X"00",X"20",X"60",X"F0",X"F0",
		X"1F",X"20",X"40",X"80",X"80",X"80",X"80",X"80",X"FF",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"80",X"80",X"80",X"80",X"80",X"40",X"20",X"1F",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5C",X"FE",X"54",X"FE",X"54",X"74",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9C",X"C8",X"E8",X"F2",X"F3",X"F2",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F2",X"F3",X"F2",X"E8",X"C8",X"9C",
		X"01",X"01",X"00",X"00",X"3F",X"7F",X"FF",X"FF",X"01",X"01",X"00",X"00",X"E0",X"E0",X"F0",X"F0",
		X"01",X"01",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"01",X"00",X"00",X"01",X"01",X"00",X"00",
		X"07",X"02",X"02",X"02",X"02",X"02",X"02",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"F0",X"F0",
		X"01",X"01",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"07",X"07",X"03",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",
		X"7F",X"7F",X"3F",X"3F",X"1F",X"0F",X"0F",X"07",X"07",X"07",X"03",X"03",X"01",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"FF",X"FF",X"01",X"01",X"01",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",X"A0",X"A0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"B0",X"B8",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E0",X"E0",X"F0",X"F0",X"F8",X"FC",X"BE",X"BF",
		X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"80",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"A0",X"80",
		X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"A0",X"A0",X"80",X"80",X"80",X"80",X"C0",X"C0",X"80",X"80",
		X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"BF",X"BF",X"F8",X"F8",X"F8",X"F8",X"FC",X"FC",X"BC",X"BC",
		X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"B0",X"B8",X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",X"A0",X"A0",
		X"80",X"80",X"80",X"C0",X"C0",X"C0",X"80",X"80",X"C0",X"C0",X"80",X"80",X"80",X"80",X"80",X"80",
		X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"A0",X"A0",
		X"FE",X"FC",X"FC",X"F8",X"F8",X"F8",X"B0",X"B0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"BE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"C0",X"E0",X"F0",X"F8",X"F8",X"BC",X"BE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"9F",X"F8",X"FC",X"FC",X"FE",X"FE",X"FF",X"BF",X"BF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E0",X"F0",X"F0",X"F0",X"F0",X"F8",X"B8",X"B8",X"F8",X"F0",X"F0",X"F0",X"F0",X"E0",X"A0",X"A0",
		X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"B8",X"B8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"BF",
		X"8F",X"9F",X"BF",X"BF",X"FF",X"FF",X"BF",X"BF",X"80",X"81",X"81",X"83",X"83",X"87",X"87",X"8F",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"83",X"81",X"81",X"80",X"80",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"07",X"06",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"04",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"20",X"20",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0E",X"1F",X"1F",X"0E",X"04",X"04",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"14",X"0C",X"0C",X"0A",X"18",X"10",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0E",X"0F",X"0F",X"0E",X"04",X"04",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"0C",X"0C",X"0A",X"09",X"08",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"D8",X"5C",X"76",X"74",X"2C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"F5",X"FA",X"F5",X"FA",X"F5",X"FA",X"75",
		X"7A",X"35",X"3A",X"15",X"1A",X"05",X"0A",X"05",X"1A",X"15",X"1A",X"15",X"0A",X"05",X"0A",X"05",
		X"FA",X"F5",X"7A",X"75",X"7A",X"35",X"3A",X"35",X"FA",X"F5",X"FA",X"75",X"7A",X"35",X"3A",X"15",
		X"EA",X"E5",X"CA",X"C5",X"CA",X"C5",X"CA",X"C5",X"CA",X"C5",X"8A",X"85",X"8A",X"85",X"8A",X"85",
		X"8A",X"85",X"8A",X"C5",X"CA",X"C5",X"CA",X"C5",X"CA",X"C5",X"EA",X"E5",X"EA",X"E5",X"EA",X"E5",
		X"7A",X"75",X"7A",X"75",X"FA",X"F5",X"FA",X"F5",X"1A",X"15",X"3A",X"35",X"3A",X"35",X"7A",X"75",
		X"7A",X"75",X"7A",X"75",X"3A",X"35",X"3A",X"35",X"3A",X"35",X"3A",X"35",X"7A",X"75",X"7A",X"75",
		X"EA",X"C5",X"CA",X"85",X"8A",X"05",X"0A",X"05",X"FA",X"F5",X"FA",X"F5",X"FA",X"F5",X"FA",X"E5",
		X"0A",X"85",X"CA",X"E5",X"FA",X"F5",X"FA",X"F5",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",
		X"FA",X"F5",X"FA",X"E5",X"EA",X"E5",X"CA",X"C5",X"CA",X"C5",X"8A",X"85",X"8A",X"85",X"8A",X"85",
		X"8A",X"85",X"8A",X"85",X"8A",X"85",X"8A",X"C5",X"CA",X"C5",X"CA",X"C5",X"CA",X"C5",X"EA",X"E5",
		X"0A",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"1A",X"15",X"1A",X"15",X"3A",X"75",X"7A",X"75",
		X"FA",X"F5",X"FA",X"F5",X"FA",X"F5",X"FA",X"F5",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"40",X"20",X"10",X"08",X"04",X"FF",X"04",X"08",X"10",X"20",X"40",X"80",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"40",X"A0",X"50",
		X"A0",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"50",
		X"A0",X"50",X"A0",X"40",X"A0",X"50",X"A0",X"50",X"AF",X"5F",X"AF",X"5F",X"AF",X"FF",X"FF",X"FF",
		X"04",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"04",X"08",X"10",X"3E",X"00",X"1A",
		X"24",X"24",X"24",X"3E",X"00",X"3E",X"02",X"02",X"02",X"3E",X"00",X"20",X"20",X"3E",X"20",X"20",
		X"00",X"22",X"2A",X"2A",X"2A",X"3E",X"00",X"1A",X"24",X"24",X"24",X"3E",X"00",X"00",X"00",X"00",
		X"00",X"02",X"02",X"02",X"02",X"3E",X"00",X"3E",X"02",X"02",X"02",X"3E",X"00",X"22",X"22",X"22",
		X"22",X"3E",X"00",X"22",X"2A",X"2A",X"2A",X"3E",X"00",X"1A",X"24",X"24",X"24",X"3E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"22",X"2A",X"2A",X"2A",X"3E",X"00",X"2E",X"2A",X"2A",X"2A",X"3A",
		X"00",X"1E",X"24",X"24",X"24",X"1E",X"00",X"1A",X"24",X"24",X"24",X"3E",X"00",X"22",X"2A",X"2A",
		X"2A",X"3E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",
		X"20",X"3E",X"20",X"20",X"00",X"3E",X"04",X"08",X"10",X"3E",X"00",X"22",X"2A",X"2A",X"2A",X"3E",
		X"00",X"3E",X"10",X"08",X"10",X"3E",X"00",X"22",X"2A",X"2A",X"2A",X"3E",X"00",X"22",X"22",X"22",
		X"22",X"3E",X"20",X"1E",X"24",X"24",X"24",X"1E",X"00",X"20",X"28",X"28",X"28",X"3E",X"00",X"20",
		X"28",X"28",X"28",X"3E",X"00",X"22",X"2A",X"2A",X"2A",X"3E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"2A",X"2A",X"2A",X"3E",X"00",X"22",X"22",X"22",X"22",
		X"3E",X"00",X"3E",X"04",X"08",X"10",X"3E",X"00",X"1E",X"24",X"24",X"24",X"1E",X"00",X"38",X"04",
		X"02",X"04",X"38",X"00",X"1C",X"22",X"22",X"22",X"3E",X"00",X"1E",X"24",X"24",X"24",X"1E",X"00",
		X"00",X"00",X"00",X"00",X"22",X"2A",X"2A",X"2A",X"3E",X"00",X"22",X"22",X"22",X"22",X"3E",X"00",
		X"3E",X"04",X"08",X"10",X"3E",X"00",X"1E",X"24",X"24",X"24",X"1E",X"00",X"38",X"04",X"02",X"04",
		X"38",X"00",X"1E",X"24",X"24",X"24",X"1A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"2A",
		X"2A",X"2A",X"3E",X"00",X"1A",X"24",X"24",X"24",X"3E",X"00",X"3E",X"02",X"02",X"02",X"3E",X"00",
		X"20",X"20",X"3E",X"20",X"20",X"00",X"3E",X"00",X"00",X"1A",X"24",X"24",X"24",X"3E",X"00",X"22",
		X"22",X"22",X"22",X"3E",X"00",X"22",X"2A",X"2A",X"2A",X"3E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"2A",X"2A",X"2A",X"3E",X"00",X"20",X"20",X"3E",
		X"20",X"20",X"00",X"3E",X"00",X"1A",X"24",X"24",X"24",X"3E",X"00",X"38",X"04",X"02",X"3C",X"02",
		X"08",X"08",X"08",X"08",X"08",X"0C",X"06",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"08",X"08",X"08",X"08",X"08",X"18",X"30",X"E0",X"E0",X"30",X"18",X"08",X"08",X"08",X"08",X"08",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"06",X"0C",X"08",X"08",X"08",X"08",X"08",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"F8",X"E4",X"E2",X"E2",X"E2",X"E3",X"E3",X"FE",X"E0",X"0E",X"31",X"61",X"E1",
		X"E1",X"E1",X"E1",X"EE",X"F0",X"E0",X"FE",X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",X"E2",X"FC",X"00",
		X"F8",X"E6",X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",X"EE",X"F0",X"E0",X"E0",X"F0",X"E8",X"E4",
		X"E2",X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",X"72",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"07",X"04",X"02",X"01",X"02",X"04",X"07",
		X"00",X"04",X"04",X"07",X"04",X"04",X"E0",X"FC",X"E2",X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",X"E2",
		X"FC",X"E0",X"80",X"00",X"FC",X"E2",X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",X"E6",X"F8",X"00",X"F8",
		X"E6",X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",X"E2",X"EC",X"F0",X"E0",X"E0",X"E0",X"F8",X"E4",
		X"E2",X"E3",X"E3",X"E3",X"E3",X"E3",X"7B",X"06",X"E0",X"FC",X"E2",X"E3",X"E3",X"E3",X"E3",X"E3",
		X"E2",X"FE",X"00",X"80",X"C0",X"E0",X"E0",X"C0",X"80",X"00",X"EC",X"E2",X"E3",X"E3",X"E3",X"E3",
		X"E3",X"E3",X"E6",X"E8",X"00",X"E0",X"E8",X"E4",X"E2",X"E2",X"E2",X"E3",X"E3",X"63",X"63",X"63",
		X"63",X"E3",X"E3",X"E3",X"E3",X"E3",X"E2",X"E2",X"E2",X"EC",X"F0",X"00",X"F8",X"E6",X"E3",X"E3",
		X"E3",X"E3",X"E3",X"E3",X"E3",X"E2",X"EC",X"F0",X"E0",X"E0",X"E0",X"E8",X"E4",X"E2",X"E2",X"E3",
		X"E3",X"E3",X"E3",X"7B",X"06",X"E0",X"E8",X"E4",X"E2",X"E3",X"E3",X"E3",X"E3",X"23",X"23",X"23",
		X"23",X"E3",X"E3",X"E3",X"E3",X"E3",X"E2",X"E2",X"FC",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",
		X"11",X"71",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"FF",X"00",X"00",
		X"07",X"19",X"71",X"F1",X"F1",X"F1",X"F1",X"F1",X"FD",X"F3",X"E1",X"F1",X"F9",X"F7",X"F1",X"F1",
		X"F1",X"F1",X"71",X"19",X"07",X"01",X"00",X"00",X"FF",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",
		X"F1",X"F1",X"F1",X"F1",X"71",X"11",X"11",X"71",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",
		X"F1",X"F1",X"F1",X"FF",X"00",X"07",X"C9",X"E9",X"E9",X"E9",X"E9",X"E9",X"E9",X"E9",X"C9",X"86",
		X"80",X"C0",X"E1",X"FF",X"F1",X"F1",X"F1",X"F1",X"F1",X"71",X"31",X"0E",X"00",X"07",X"19",X"71",
		X"F1",X"F1",X"F1",X"F1",X"F1",X"FD",X"F3",X"E1",X"F1",X"F9",X"F7",X"F1",X"F1",X"F1",X"F1",X"71",
		X"19",X"07",X"01",X"00",X"00",X"01",X"03",X"05",X"05",X"09",X"09",X"C9",X"F1",X"F1",X"F1",X"91",
		X"91",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"04",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"07",
		X"00",X"00",X"03",X"04",X"04",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"06",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"02",X"02",X"04",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"04",
		X"06",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"04",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"0C",X"04",X"04",X"03",X"00",X"00",X"00",X"00",X"03",X"04",X"04",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"0C",X"0C",X"06",X"01",X"00",X"00",X"00",X"01",X"02",X"02",X"04",X"04",X"0C",X"0C",X"0C",X"0C",
		X"0C",X"0C",X"0C",X"0C",X"04",X"04",X"02",X"01",X"00",X"01",X"02",X"02",X"04",X"0C",X"0C",X"0C",
		X"0C",X"0C",X"0C",X"0C",X"04",X"06",X"01",X"00",X"00",X"00",X"00",X"01",X"02",X"04",X"04",X"0C",
		X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"04",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"E0",X"E0",X"E0",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"0F",X"3F",X"FF",X"FF",X"FF",X"E7",X"87",X"07",X"07",X"07",X"07",X"87",X"E7",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"03",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"E0",X"E0",X"20",X"00",X"00",X"00",
		X"3F",X"0F",X"07",X"07",X"07",X"07",X"07",X"07",X"00",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"80",
		X"07",X"3F",X"3F",X"3F",X"1F",X"1F",X"1F",X"0F",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"E0",
		X"0F",X"0F",X"07",X"07",X"07",X"07",X"07",X"3F",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"80",X"00",X"00",X"00",
		X"3F",X"07",X"07",X"07",X"07",X"C7",X"F7",X"FF",X"FF",X"7F",X"1F",X"07",X"01",X"00",X"00",X"00",
		X"00",X"01",X"07",X"1F",X"7F",X"FF",X"FC",X"F8",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"07",X"07",X"07",X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"07",X"07",X"07",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"12",X"01",X"00",X"22",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"50",X"00",X"00",X"00",X"00",X"02",X"15",X"2A",X"55",
		X"00",X"00",X"00",X"00",X"80",X"40",X"A8",X"55",X"00",X"01",X"02",X"15",X"AA",X"55",X"AA",X"55",
		X"80",X"40",X"80",X"50",X"A8",X"55",X"AA",X"55",X"0A",X"15",X"2A",X"55",X"AA",X"55",X"AA",X"55",
		X"0A",X"50",X"A8",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",
		X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"FF",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"FF",
		X"0F",X"07",X"07",X"07",X"00",X"00",X"00",X"00",X"07",X"07",X"03",X"03",X"01",X"01",X"01",X"00",
		X"7F",X"7F",X"3F",X"3F",X"1F",X"1F",X"0F",X"0F",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"FC",X"FC",
		X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"0F",X"1F",X"1F",X"1F",X"3F",X"3F",X"3F",X"7F",
		X"E0",X"F0",X"F0",X"F8",X"F8",X"F8",X"FC",X"FC",X"C0",X"E0",X"E0",X"F0",X"F8",X"F8",X"FC",X"FE",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F8",X"F8",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"80",X"FC",X"FC",X"FC",X"F8",X"F8",X"F0",X"F0",X"F0",
		X"01",X"01",X"00",X"00",X"FE",X"FE",X"FE",X"FE",X"01",X"01",X"00",X"00",X"03",X"03",X"03",X"03",
		X"7F",X"3F",X"3F",X"1F",X"1F",X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",
		X"80",X"C0",X"C0",X"C0",X"E0",X"E0",X"E0",X"F0",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",
		X"FF",X"FE",X"FE",X"FE",X"00",X"00",X"10",X"10",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"07",X"07",X"07",X"07",X"00",X"00",X"10",X"10",X"E0",X"C0",X"00",X"00",X"00",X"00",X"10",X"10",
		X"01",X"01",X"00",X"00",X"E0",X"E0",X"E0",X"E0",X"01",X"01",X"00",X"00",X"1F",X"1F",X"0F",X"0F",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"E0",X"E0",X"F0",X"F0",
		X"FE",X"FE",X"FC",X"FC",X"FC",X"F8",X"F8",X"F8",X"07",X"07",X"06",X"04",X"00",X"00",X"10",X"10",
		X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"F0",X"F0",X"E0",X"E0",X"C0",X"C0",X"80",X"00",
		X"80",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"80",
		X"1F",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"07",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"E0",
		X"00",X"80",X"80",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FE",X"FE",X"FE",
		X"C0",X"C0",X"C0",X"E0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"FC",X"FC",
		X"FE",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"00",X"00",X"10",X"10",X"01",X"01",X"00",X"00",X"80",X"80",X"80",X"80",
		X"FF",X"FF",X"7F",X"7F",X"7F",X"3F",X"3F",X"3F",X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"03",
		X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"01",X"01",X"00",X"00",X"7F",X"3F",X"1F",X"1F",
		X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"3F",X"3F",X"3F",X"3F",X"7F",X"7F",X"7F",X"7F",
		X"03",X"03",X"03",X"03",X"00",X"00",X"10",X"10",X"01",X"01",X"00",X"00",X"0F",X"0F",X"0F",X"0F",
		X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",X"3F",X"1F",
		X"7F",X"7F",X"3F",X"3F",X"3F",X"1F",X"1F",X"1F",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"C0",X"E0",X"E0",X"F0",X"F0",X"F8",X"FC",X"C0",X"E0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F8",
		X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",X"FE",X"FE",
		X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",
		X"7F",X"3F",X"3F",X"1F",X"1F",X"0F",X"0F",X"07",X"07",X"03",X"03",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"1F",X"0F",X"0F",X"07",X"03",X"03",X"01",X"01",
		X"FF",X"FF",X"7F",X"7F",X"3F",X"3F",X"1F",X"1F",X"0F",X"07",X"07",X"03",X"03",X"03",X"01",X"01",
		X"7F",X"3F",X"3F",X"1F",X"1F",X"1F",X"0F",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",
		X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"01",X"1F",X"1F",X"1F",X"1F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"E0",X"E0",X"F0",X"F0",X"F8",X"FC",X"FE",X"FF",
		X"C0",X"C0",X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"F0",X"F0",X"F0",X"00",X"00",X"10",X"10",
		X"7F",X"7F",X"7F",X"7F",X"00",X"00",X"10",X"10",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"03",X"03",X"03",X"07",X"07",X"07",X"0F",X"0F",X"0F",X"1F",X"1F",X"1F",X"3F",
		X"3F",X"3F",X"7F",X"3F",X"00",X"00",X"10",X"10",X"01",X"01",X"00",X"00",X"F0",X"F0",X"F0",X"F0",
		X"01",X"01",X"00",X"00",X"F0",X"F0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"C0",
		X"FE",X"FC",X"7C",X"38",X"00",X"00",X"10",X"10",X"01",X"01",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"10",X"10",X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"7F",X"3F",X"00",X"00",X"10",X"10",X"01",X"01",X"00",X"00",X"3F",X"7F",X"FF",X"FF",
		X"FF",X"FF",X"FE",X"FC",X"00",X"00",X"10",X"10",X"01",X"01",X"00",X"00",X"FC",X"FE",X"FF",X"FF",
		X"01",X"01",X"00",X"00",X"01",X"01",X"00",X"00",X"7F",X"7F",X"7F",X"3F",X"3F",X"3F",X"1F",X"1F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"3F",X"3F",X"3F",X"00",X"00",X"10",X"10",
		X"01",X"01",X"00",X"00",X"07",X"07",X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",X"3F",X"3F",X"00",X"01",X"01",X"01",X"01",X"03",X"03",X"03",
		X"03",X"07",X"07",X"07",X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"7F",X"7F",X"1F",X"1F",X"1F",X"1F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"07",X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"03",X"01",X"01",X"00",X"00",X"10",X"10",
		X"01",X"01",X"00",X"00",X"01",X"01",X"00",X"00",X"7F",X"7F",X"3F",X"3F",X"1F",X"1F",X"1F",X"0F",
		X"0F",X"0F",X"07",X"07",X"07",X"03",X"03",X"03",X"03",X"03",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"03",X"03",X"03",X"03",X"03",X"03",X"07",X"07",X"07",X"07",X"0F",
		X"80",X"C0",X"E0",X"F0",X"F8",X"F8",X"FC",X"FE",X"00",X"80",X"C0",X"E0",X"F0",X"F8",X"FC",X"FE",
		X"00",X"80",X"C0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FE",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",X"F0",X"F0",X"E0",X"E0",X"C0",X"80",X"00",
		X"FE",X"FC",X"F8",X"F0",X"E0",X"C0",X"80",X"00",X"FF",X"FE",X"FC",X"FC",X"F8",X"F0",X"F0",X"E0",
		X"E0",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"FE",X"FC",X"FC",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",
		X"80",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"F0",
		X"F8",X"F8",X"F8",X"F8",X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"E0",X"E0",X"00",X"00",X"10",X"10",
		X"01",X"01",X"00",X"00",X"C0",X"E0",X"E0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",
		X"F8",X"F8",X"F8",X"F8",X"00",X"00",X"10",X"10",X"01",X"01",X"00",X"00",X"C0",X"C0",X"C0",X"80",
		X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"03",X"03",X"03",X"07",
		X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",X"3F",X"3F",X"7F",X"7F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"1F",X"1F",X"00",X"00",X"10",X"10",X"0F",X"0F",X"0F",X"07",X"07",X"07",X"03",X"03",
		X"03",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"03",
		X"03",X"03",X"03",X"07",X"07",X"07",X"0F",X"0F",X"0F",X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",X"3F",
		X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",
		X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"C0",X"C0",
		X"C0",X"C0",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"C0",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",X"F0",X"F0",X"00",X"00",X"10",X"10",
		X"00",X"00",X"07",X"03",X"01",X"01",X"00",X"00",X"FC",X"FC",X"FC",X"FE",X"FE",X"FE",X"FF",X"FF",
		X"01",X"01",X"00",X"00",X"20",X"60",X"F0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",X"1F",X"1F",X"0F",X"07",X"03",X"03",
		X"00",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"C0",X"C0",X"E0",X"F0",X"F0",X"F8",X"F8",
		X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"E0",
		X"F0",X"F0",X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"80",X"C0",X"E0",X"F0",X"F0",X"F8",X"F8",X"FC",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",
		X"03",X"03",X"03",X"03",X"03",X"07",X"07",X"07",X"07",X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"03",X"03",X"03",
		X"03",X"01",X"01",X"01",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"03",X"03",X"03",X"07",X"07",X"0F",X"0F",X"0F",X"1F",X"1F",X"1F",X"3F",X"3F",X"7F",X"7F",X"7F",
		X"FF",X"FF",X"FE",X"FC",X"00",X"00",X"10",X"10",X"01",X"01",X"00",X"00",X"0C",X"06",X"07",X"03",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"01",X"03",X"03",X"07",X"07",X"0F",X"0F",X"1F",X"3F",X"3F",X"7F",X"7F",X"FF",X"FF",
		X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",
		X"E0",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",
		X"1F",X"0F",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"01",X"01",X"01",X"01",X"01",X"01",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"F0",X"F0",
		X"01",X"01",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"07",X"07",X"03",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",
		X"7F",X"7F",X"3F",X"3F",X"1F",X"1F",X"0F",X"0F",X"07",X"07",X"03",X"03",X"01",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"FF",X"FF",X"01",X"01",X"01");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
