library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_OBJ_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_OBJ_1 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"7C",X"C6",X"C6",X"82",X"C6",X"C6",X"7C",X"00",X"00",X"00",X"FE",X"FE",X"8E",X"00",X"00",
		X"00",X"66",X"F2",X"BA",X"9E",X"8E",X"C6",X"62",X"00",X"FE",X"FE",X"92",X"92",X"82",X"C6",X"C6",
		X"00",X"18",X"FE",X"1E",X"1A",X"D8",X"F8",X"F8",X"00",X"9C",X"BE",X"B2",X"B2",X"B2",X"F6",X"F6",
		X"00",X"4C",X"DE",X"92",X"92",X"92",X"FE",X"7C",X"00",X"E0",X"F0",X"98",X"8E",X"86",X"C2",X"E0",
		X"00",X"6C",X"FE",X"92",X"92",X"92",X"FE",X"6C",X"00",X"7C",X"FE",X"92",X"92",X"92",X"F6",X"64",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"3C",X"42",X"81",X"A5",X"A5",X"99",X"42",X"3C",
		X"00",X"00",X"00",X"18",X"18",X"04",X"03",X"02",X"00",X"00",X"00",X"18",X"18",X"20",X"C0",X"40",
		X"02",X"03",X"04",X"18",X"18",X"00",X"00",X"00",X"40",X"C0",X"20",X"18",X"18",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7E",X"D6",X"D0",X"D0",X"D0",X"D6",X"7E",
		X"00",X"44",X"EE",X"BA",X"92",X"82",X"FE",X"FE",X"00",X"44",X"C6",X"82",X"82",X"82",X"FE",X"7C",
		X"00",X"7C",X"FE",X"82",X"82",X"BA",X"FE",X"FE",X"00",X"C6",X"C6",X"92",X"92",X"92",X"FE",X"FE",
		X"00",X"C0",X"C0",X"90",X"92",X"96",X"FE",X"FE",X"00",X"6C",X"EE",X"8A",X"8A",X"82",X"FE",X"7C",
		X"00",X"FE",X"FE",X"D0",X"10",X"16",X"FE",X"FE",X"00",X"00",X"C6",X"FE",X"FE",X"FE",X"C6",X"00",
		X"00",X"FC",X"FE",X"C2",X"06",X"0E",X"0C",X"08",X"00",X"82",X"C6",X"EE",X"38",X"92",X"FE",X"FE",
		X"00",X"1E",X"0E",X"06",X"02",X"E2",X"FE",X"FE",X"00",X"FE",X"C6",X"60",X"30",X"60",X"C6",X"FE",
		X"00",X"FE",X"CE",X"9C",X"38",X"72",X"E6",X"FE",X"00",X"7C",X"EE",X"C6",X"C6",X"C6",X"EE",X"7C",
		X"00",X"60",X"F0",X"90",X"90",X"92",X"FE",X"FE",X"00",X"06",X"7E",X"F6",X"CE",X"C6",X"DE",X"7C",
		X"00",X"62",X"F6",X"9E",X"90",X"96",X"FE",X"FE",X"00",X"C4",X"8E",X"9A",X"9A",X"B2",X"F2",X"66",
		X"00",X"F0",X"C2",X"FE",X"FE",X"FE",X"C2",X"F0",X"00",X"FC",X"FE",X"FA",X"02",X"02",X"FE",X"FC",
		X"00",X"C0",X"F8",X"FC",X"0E",X"FC",X"F8",X"C0",X"00",X"FE",X"C6",X"0C",X"18",X"0C",X"C6",X"FE",
		X"00",X"C6",X"C6",X"28",X"10",X"28",X"C6",X"C6",X"00",X"FE",X"FE",X"D2",X"12",X"16",X"F6",X"F6",
		X"00",X"CE",X"E2",X"F2",X"BA",X"9E",X"8E",X"E6",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"00",X"00",X"04",X"00",X"70",X"89",X"8F",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",
		X"00",X"00",X"00",X"08",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"1C",X"08",X"00",X"00",
		X"00",X"00",X"08",X"1C",X"34",X"08",X"00",X"00",X"00",X"00",X"0C",X"28",X"04",X"2E",X"14",X"00",
		X"00",X"08",X"A0",X"88",X"7C",X"20",X"48",X"00",X"38",X"60",X"8A",X"8A",X"22",X"58",X"38",X"00",
		X"10",X"24",X"00",X"40",X"44",X"42",X"28",X"10",X"02",X"10",X"04",X"02",X"00",X"20",X"02",X"0C",
		X"01",X"08",X"00",X"01",X"00",X"10",X"01",X"06",X"04",X"01",X"00",X"01",X"00",X"09",X"01",X"02",
		X"07",X"0F",X"1F",X"1E",X"1E",X"1F",X"0F",X"07",X"19",X"3B",X"7C",X"78",X"78",X"7C",X"3B",X"19",
		X"31",X"72",X"9C",X"F0",X"F0",X"9C",X"72",X"31",X"19",X"3B",X"4C",X"78",X"78",X"4C",X"3B",X"19",
		X"1C",X"31",X"5F",X"F8",X"F8",X"5F",X"31",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"0E",
		X"00",X"00",X"00",X"00",X"0E",X"EE",X"E0",X"EE",X"00",X"00",X"E0",X"EE",X"0E",X"EE",X"E0",X"EE",
		X"0E",X"EE",X"E0",X"EE",X"0E",X"EE",X"E0",X"EE",X"0E",X"EE",X"E0",X"EE",X"0E",X"EE",X"00",X"00",
		X"0E",X"EE",X"E0",X"EE",X"00",X"00",X"00",X"00",X"0E",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3B",X"44",X"92",X"BA",X"92",X"44",X"B8",X"81",X"F0",X"08",X"04",X"02",X"C1",X"21",X"11",X"91",
		X"89",X"88",X"84",X"83",X"40",X"20",X"10",X"0F",X"91",X"11",X"21",X"C1",X"02",X"04",X"08",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"05",X"08",X"09",X"02",X"05",X"05",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"03",X"03",X"08",X"10",X"03",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"1B",X"38",X"3F",X"00",X"00",X"3C",X"1C",X"08",X"88",X"F8",X"40",
		X"2F",X"09",X"0D",X"00",X"00",X"00",X"00",X"00",X"24",X"2C",X"1C",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"1F",X"3F",X"3F",X"00",X"00",X"3C",X"1C",X"08",X"88",X"F8",X"C0",
		X"2E",X"0B",X"0B",X"03",X"02",X"00",X"00",X"00",X"64",X"6C",X"3C",X"04",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"1F",X"3F",X"3D",X"00",X"00",X"3C",X"1C",X"08",X"88",X"F8",X"40",
		X"2E",X"0B",X"0D",X"01",X"00",X"00",X"00",X"00",X"64",X"6C",X"BC",X"84",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"25",X"20",X"12",X"03",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"05",X"48",X"88",X"10",X"03",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"A1",X"82",X"46",X"04",X"00",X"00",X"01",
		X"00",X"00",X"00",X"02",X"04",X"00",X"00",X"00",X"00",X"21",X"21",X"44",X"81",X"02",X"00",X"04",
		X"20",X"98",X"8B",X"64",X"00",X"2E",X"42",X"44",X"30",X"88",X"48",X"7E",X"19",X"34",X"44",X"43",
		X"30",X"08",X"08",X"66",X"81",X"A5",X"14",X"23",X"83",X"4C",X"69",X"1E",X"18",X"24",X"42",X"C1",
		X"02",X"12",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"18",X"20",X"20",X"00",X"00",X"00",
		X"00",X"06",X"24",X"48",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"0C",X"02",X"40",X"00",
		X"08",X"08",X"04",X"20",X"10",X"00",X"00",X"00",X"00",X"20",X"10",X"00",X"00",X"00",X"00",X"00",
		X"18",X"50",X"A0",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"40",X"20",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"00",X"09",X"14",X"02",X"00",X"40",X"C0",X"20",X"00",X"40",X"80",X"00",
		X"00",X"4C",X"11",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",
		X"3C",X"4E",X"A7",X"96",X"67",X"0E",X"1F",X"18",X"3C",X"4E",X"87",X"86",X"97",X"6E",X"1F",X"18",
		X"3D",X"4E",X"86",X"87",X"86",X"8E",X"9D",X"40",X"3D",X"4E",X"86",X"87",X"96",X"6E",X"1D",X"00",
		X"00",X"00",X"00",X"01",X"02",X"02",X"63",X"00",X"00",X"00",X"00",X"40",X"90",X"A0",X"E0",X"00",
		X"00",X"63",X"02",X"02",X"01",X"00",X"00",X"00",X"00",X"E0",X"A0",X"90",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"0D",X"00",X"00",X"00",X"40",X"00",X"00",X"E0",X"F8",
		X"0D",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"E0",X"00",X"00",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"33",X"0D",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"F8",
		X"0D",X"33",X"01",X"00",X"00",X"00",X"00",X"00",X"F8",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"20",X"10",X"16",X"09",X"61",X"93",X"96",X"80",X"40",X"40",X"C0",X"00",X"8C",X"CA",X"72",
		X"0E",X"03",X"05",X"88",X"68",X"10",X"01",X"02",X"69",X"C9",X"84",X"48",X"20",X"C0",X"00",X"00",
		X"00",X"00",X"22",X"51",X"11",X"0D",X"03",X"06",X"20",X"40",X"40",X"80",X"00",X"88",X"D6",X"71",
		X"1E",X"D3",X"31",X"02",X"01",X"00",X"01",X"01",X"60",X"C0",X"B0",X"08",X"10",X"96",X"08",X"00",
		X"7E",X"87",X"81",X"87",X"81",X"87",X"81",X"7E",X"3C",X"4E",X"42",X"4E",X"42",X"4E",X"42",X"3C",
		X"18",X"3C",X"24",X"3C",X"24",X"3C",X"24",X"18",X"3C",X"4E",X"42",X"4E",X"42",X"4E",X"42",X"3C",
		X"00",X"00",X"00",X"00",X"00",X"49",X"5B",X"ED",X"00",X"00",X"00",X"00",X"00",X"24",X"6C",X"B6",
		X"6D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B6",X"00",X"04",X"04",X"0A",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"24",X"6D",X"6D",X"00",X"00",X"00",X"00",X"00",X"92",X"B6",X"B6",
		X"6D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B6",X"00",X"04",X"0A",X"11",X"00",X"00",X"00",
		X"00",X"01",X"01",X"00",X"01",X"01",X"00",X"01",X"00",X"C0",X"E0",X"00",X"C0",X"E0",X"00",X"C0",
		X"01",X"00",X"01",X"11",X"08",X"05",X"09",X"10",X"E0",X"00",X"C0",X"E0",X"00",X"C0",X"E0",X"00",
		X"00",X"01",X"01",X"00",X"01",X"01",X"00",X"01",X"80",X"E0",X"80",X"40",X"E0",X"80",X"40",X"E0",
		X"01",X"00",X"01",X"01",X"10",X"0D",X"11",X"00",X"80",X"40",X"E0",X"80",X"40",X"E0",X"80",X"00",
		X"00",X"1F",X"20",X"40",X"9C",X"91",X"92",X"82",X"00",X"F0",X"08",X"44",X"A4",X"14",X"8C",X"2C",
		X"82",X"9E",X"91",X"90",X"40",X"20",X"1F",X"00",X"8C",X"2C",X"14",X"A4",X"44",X"08",X"F0",X"00",
		X"00",X"1F",X"20",X"40",X"90",X"99",X"9D",X"81",X"00",X"F0",X"08",X"44",X"A4",X"14",X"94",X"34",
		X"81",X"91",X"99",X"9C",X"40",X"20",X"1F",X"00",X"14",X"94",X"34",X"A4",X"44",X"08",X"F0",X"00",
		X"00",X"1F",X"20",X"40",X"84",X"8C",X"9C",X"80",X"00",X"F0",X"08",X"44",X"A4",X"A4",X"A4",X"A4",
		X"80",X"84",X"8C",X"9C",X"40",X"20",X"1F",X"00",X"A4",X"A4",X"A4",X"A4",X"44",X"08",X"F0",X"00",
		X"00",X"1F",X"20",X"40",X"9C",X"8C",X"84",X"80",X"00",X"F0",X"08",X"44",X"44",X"44",X"44",X"44",
		X"80",X"9C",X"8C",X"84",X"40",X"20",X"1F",X"00",X"44",X"44",X"44",X"44",X"44",X"08",X"F0",X"00",
		X"00",X"03",X"07",X"0F",X"1F",X"1F",X"3F",X"3F",X"00",X"C0",X"E0",X"F0",X"F8",X"F8",X"FC",X"FC",
		X"3F",X"3F",X"1F",X"1F",X"0F",X"07",X"03",X"00",X"FC",X"FC",X"F8",X"F8",X"F0",X"E0",X"C0",X"00",
		X"00",X"03",X"07",X"0F",X"1F",X"1F",X"3E",X"3E",X"00",X"C0",X"E0",X"F0",X"F8",X"F8",X"7C",X"7C",
		X"3E",X"3E",X"1F",X"1F",X"0F",X"07",X"03",X"00",X"7C",X"7C",X"F8",X"F8",X"F0",X"E0",X"C0",X"00",
		X"00",X"03",X"07",X"0F",X"1F",X"1F",X"3C",X"3C",X"00",X"C0",X"E0",X"F0",X"F8",X"F8",X"3C",X"3C",
		X"3C",X"3C",X"1F",X"1F",X"0F",X"07",X"03",X"00",X"3C",X"3C",X"F8",X"F8",X"F0",X"E0",X"C0",X"00",
		X"00",X"03",X"07",X"0F",X"1F",X"1F",X"3C",X"3C",X"00",X"C0",X"E0",X"F0",X"F8",X"F8",X"3C",X"3C",
		X"3C",X"3C",X"1F",X"1F",X"0F",X"07",X"03",X"00",X"3C",X"3C",X"F8",X"F8",X"F0",X"E0",X"C0",X"00",
		X"01",X"01",X"01",X"01",X"01",X"00",X"01",X"1B",X"80",X"80",X"80",X"80",X"80",X"00",X"80",X"D8",
		X"1B",X"01",X"00",X"01",X"01",X"01",X"01",X"01",X"D8",X"80",X"00",X"80",X"80",X"80",X"80",X"80",
		X"00",X"20",X"50",X"28",X"14",X"0A",X"05",X"03",X"00",X"00",X"00",X"00",X"20",X"70",X"A0",X"C0",
		X"03",X"05",X"0E",X"04",X"00",X"00",X"00",X"00",X"C0",X"A0",X"50",X"28",X"14",X"0A",X"04",X"00",
		X"00",X"00",X"00",X"01",X"01",X"00",X"01",X"FB",X"00",X"00",X"00",X"80",X"80",X"00",X"80",X"DF",
		X"FB",X"01",X"00",X"01",X"01",X"00",X"00",X"00",X"DF",X"80",X"00",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"04",X"03",X"0B",X"00",X"00",X"00",X"00",X"80",X"20",X"C0",X"D0",
		X"0B",X"03",X"04",X"01",X"00",X"00",X"00",X"00",X"D0",X"C0",X"20",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"06",X"0F",X"08",X"18",X"18",X"1F",X"01",X"01",X"01",X"01",X"80",X"80",X"C0",X"C0",
		X"18",X"18",X"08",X"0F",X"06",X"00",X"00",X"00",X"C0",X"80",X"80",X"01",X"01",X"01",X"01",X"01",
		X"00",X"00",X"30",X"78",X"44",X"C6",X"C7",X"FF",X"00",X"00",X"00",X"04",X"1C",X"10",X"20",X"00",
		X"C7",X"C6",X"44",X"78",X"30",X"00",X"00",X"00",X"20",X"10",X"1C",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"03",X"01",X"01",X"C1",X"E1",X"11",X"10",X"18",X"F8",
		X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"18",X"10",X"11",X"E1",X"C1",X"01",X"01",X"01",
		X"00",X"00",X"01",X"02",X"16",X"2D",X"7B",X"7F",X"00",X"C4",X"06",X"0A",X"12",X"E2",X"E0",X"C0",
		X"53",X"1B",X"1A",X"00",X"00",X"00",X"00",X"00",X"C0",X"50",X"70",X"10",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"1E",X"3F",X"7F",X"7F",X"00",X"18",X"20",X"70",X"10",X"E0",X"C0",X"C0",
		X"53",X"1B",X"1A",X"00",X"00",X"00",X"00",X"00",X"C0",X"40",X"20",X"18",X"10",X"60",X"00",X"00",
		X"00",X"00",X"00",X"00",X"1E",X"3F",X"7F",X"77",X"00",X"00",X"00",X"00",X"74",X"2C",X"DC",X"84",
		X"53",X"1B",X"1A",X"00",X"00",X"00",X"00",X"00",X"E8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"1E",X"3F",X"7B",X"7D",X"00",X"18",X"20",X"70",X"10",X"20",X"C4",X"8C",
		X"56",X"1B",X"1D",X"00",X"00",X"00",X"00",X"00",X"FC",X"04",X"88",X"80",X"00",X"00",X"00",X"00",
		X"00",X"03",X"07",X"1C",X"3E",X"3F",X"7F",X"7D",X"00",X"80",X"00",X"04",X"04",X"FC",X"CC",X"84",
		X"7E",X"7D",X"3F",X"3F",X"1C",X"07",X"03",X"00",X"20",X"F0",X"F8",X"88",X"08",X"00",X"C0",X"00",
		X"00",X"03",X"07",X"1C",X"3F",X"3F",X"7D",X"7E",X"00",X"C0",X"00",X"04",X"04",X"FC",X"CC",X"00",
		X"7D",X"7F",X"3F",X"3F",X"1C",X"07",X"03",X"00",X"80",X"CC",X"FC",X"04",X"04",X"00",X"C0",X"00",
		X"00",X"03",X"07",X"1C",X"3E",X"27",X"6F",X"7F",X"00",X"80",X"00",X"04",X"04",X"FC",X"CC",X"80",
		X"7F",X"6F",X"27",X"3F",X"1C",X"07",X"03",X"00",X"A0",X"F0",X"F0",X"98",X"08",X"00",X"C0",X"00",
		X"00",X"03",X"07",X"1C",X"3F",X"27",X"6D",X"79",X"00",X"C0",X"00",X"04",X"04",X"FC",X"CC",X"80",
		X"79",X"6D",X"27",X"3F",X"1C",X"07",X"03",X"00",X"80",X"CC",X"FC",X"04",X"04",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"0E",X"1F",X"1F",X"3E",X"3F",X"00",X"00",X"00",X"02",X"82",X"FE",X"E6",X"00",
		X"3E",X"3F",X"1F",X"1F",X"0E",X"00",X"00",X"00",X"C0",X"E6",X"FE",X"82",X"02",X"00",X"00",X"00",
		X"00",X"00",X"07",X"1C",X"3F",X"25",X"6D",X"78",X"00",X"00",X"84",X"C4",X"7C",X"3C",X"80",X"00",
		X"78",X"6D",X"25",X"3F",X"1C",X"07",X"00",X"00",X"00",X"80",X"3C",X"7C",X"C4",X"84",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
