library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity TRIPLEDRAWPOKER_ROM_PGM_0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of TRIPLEDRAWPOKER_ROM_PGM_0 is
	type rom is array(0 to  12287) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"ED",X"56",X"31",X"00",X"44",X"C3",X"7B",X"00",X"E5",X"C5",X"F5",X"04",X"0C",X"C3",X"71",X"00",
		X"85",X"6F",X"30",X"01",X"24",X"7E",X"C9",X"FF",X"E5",X"B7",X"ED",X"52",X"E1",X"C9",X"28",X"28",
		X"E5",X"77",X"23",X"10",X"FC",X"E1",X"C9",X"AD",X"E1",X"87",X"85",X"6F",X"30",X"3C",X"18",X"39",
		X"47",X"00",X"FD",X"36",X"41",X"00",X"28",X"E1",X"C3",X"29",X"0B",X"D5",X"F5",X"BE",X"30",X"05",
		X"16",X"00",X"5F",X"19",X"19",X"23",X"5E",X"23",X"56",X"EB",X"F1",X"D1",X"E9",X"A7",X"C8",X"E5",
		X"D5",X"C5",X"06",X"00",X"4F",X"09",X"EB",X"09",X"41",X"1B",X"2B",X"1A",X"BE",X"20",X"02",X"10",
		X"F8",X"79",X"C1",X"D1",X"E1",X"C9",X"C3",X"27",X"08",X"24",X"7E",X"23",X"66",X"6F",X"E9",X"77",
		X"23",X"0D",X"C2",X"6F",X"00",X"10",X"F8",X"F1",X"C1",X"E1",X"C9",X"FD",X"21",X"8E",X"40",X"21",
		X"84",X"00",X"18",X"04",X"CD",X"BC",X"00",X"E9",X"F3",X"CD",X"6C",X"0A",X"01",X"00",X"04",X"11",
		X"00",X"40",X"AF",X"CD",X"7B",X"0A",X"12",X"13",X"0D",X"20",X"FB",X"10",X"F6",X"CD",X"35",X"07",
		X"CD",X"DD",X"02",X"CD",X"8E",X"04",X"CD",X"2E",X"06",X"CD",X"FC",X"15",X"CD",X"C2",X"02",X"28",
		X"07",X"38",X"05",X"CD",X"C1",X"08",X"18",X"03",X"CD",X"BA",X"08",X"E9",X"F5",X"18",X"1C",X"D5",
		X"E5",X"FD",X"E5",X"D1",X"21",X"02",X"00",X"7D",X"21",X"00",X"00",X"19",X"36",X"00",X"21",X"48",
		X"00",X"19",X"EB",X"3D",X"20",X"F2",X"CD",X"AE",X"0E",X"E1",X"D1",X"3A",X"45",X"40",X"E6",X"08",
		X"20",X"06",X"CD",X"AE",X"02",X"28",X"D8",X"AF",X"CD",X"A9",X"01",X"CD",X"F0",X"00",X"F1",X"C9",
		X"FD",X"E5",X"E5",X"D5",X"C5",X"F5",X"01",X"02",X"00",X"41",X"4F",X"FD",X"E5",X"D1",X"AF",X"C5",
		X"21",X"02",X"00",X"19",X"01",X"07",X"04",X"48",X"06",X"00",X"CF",X"21",X"02",X"00",X"19",X"CF",
		X"21",X"48",X"00",X"19",X"EB",X"C1",X"10",X"E7",X"FD",X"E5",X"D1",X"41",X"3A",X"4A",X"40",X"21",
		X"01",X"00",X"19",X"77",X"79",X"90",X"3C",X"21",X"00",X"00",X"19",X"77",X"21",X"48",X"00",X"19",
		X"EB",X"05",X"20",X"E8",X"CD",X"DF",X"18",X"41",X"FD",X"E5",X"D1",X"FD",X"E5",X"AF",X"21",X"01",
		X"00",X"19",X"BE",X"28",X"2E",X"21",X"01",X"00",X"19",X"35",X"79",X"90",X"3C",X"21",X"00",X"00",
		X"19",X"77",X"D5",X"FD",X"E1",X"C5",X"CD",X"2A",X"03",X"CD",X"96",X"28",X"C1",X"21",X"01",X"00",
		X"19",X"7E",X"A7",X"20",X"0E",X"79",X"90",X"3C",X"D5",X"FD",X"E1",X"C5",X"CD",X"2A",X"03",X"CD",
		X"D0",X"11",X"C1",X"21",X"48",X"00",X"19",X"EB",X"10",X"C3",X"D1",X"D5",X"AF",X"41",X"21",X"01",
		X"00",X"19",X"BE",X"20",X"C0",X"21",X"48",X"00",X"19",X"EB",X"10",X"F2",X"FD",X"E1",X"41",X"11",
		X"48",X"00",X"79",X"90",X"3C",X"CD",X"15",X"06",X"FD",X"19",X"10",X"F6",X"CD",X"35",X"0B",X"CD",
		X"D3",X"10",X"F1",X"C1",X"D1",X"E1",X"FD",X"E1",X"C9",X"E5",X"C5",X"F5",X"4F",X"06",X"FF",X"18",
		X"0B",X"CD",X"15",X"08",X"CD",X"AE",X"02",X"CD",X"58",X"12",X"06",X"00",X"CD",X"81",X"0A",X"28",
		X"F0",X"0C",X"0D",X"20",X"16",X"6F",X"CD",X"AE",X"02",X"BD",X"38",X"E5",X"CD",X"15",X"08",X"45",
		X"CD",X"8F",X"02",X"10",X"FB",X"7D",X"21",X"45",X"40",X"CB",X"E6",X"6F",X"F1",X"7D",X"C1",X"E1",
		X"C9",X"E5",X"F5",X"21",X"45",X"40",X"3A",X"3D",X"40",X"E6",X"03",X"FE",X"03",X"20",X"0F",X"7E",
		X"E6",X"40",X"28",X"3C",X"D5",X"11",X"8E",X"40",X"CD",X"47",X"03",X"D1",X"18",X"32",X"FE",X"01",
		X"20",X"2E",X"7E",X"E6",X"30",X"FE",X"30",X"20",X"27",X"CB",X"A6",X"D5",X"C5",X"21",X"44",X"40",
		X"ED",X"5B",X"CA",X"12",X"01",X"02",X"01",X"CD",X"FC",X"08",X"7A",X"C6",X"10",X"57",X"3A",X"45",
		X"40",X"E6",X"02",X"3E",X"20",X"28",X"04",X"01",X"20",X"00",X"79",X"CD",X"CC",X"0B",X"C1",X"D1",
		X"CD",X"65",X"04",X"F1",X"E1",X"C9",X"F5",X"CD",X"7A",X"08",X"28",X"14",X"E5",X"21",X"45",X"40",
		X"CB",X"5E",X"20",X"0B",X"CD",X"52",X"02",X"3D",X"20",X"FA",X"CB",X"E6",X"CD",X"3F",X"1C",X"E1",
		X"F1",X"C9",X"E5",X"D5",X"C5",X"F5",X"11",X"44",X"40",X"21",X"45",X"40",X"CB",X"56",X"28",X"13",
		X"1A",X"FE",X"99",X"38",X"04",X"CB",X"CE",X"18",X"21",X"CB",X"4E",X"20",X"04",X"CB",X"CE",X"18",
		X"19",X"CB",X"8E",X"7E",X"E6",X"01",X"3C",X"47",X"1A",X"80",X"27",X"30",X"02",X"3E",X"99",X"12",
		X"4F",X"AF",X"90",X"27",X"47",X"79",X"B8",X"D4",X"C1",X"08",X"F1",X"C1",X"D1",X"E1",X"C9",X"E5",
		X"F5",X"21",X"44",X"40",X"3A",X"45",X"40",X"E6",X"01",X"28",X"05",X"7E",X"FE",X"99",X"30",X"03",
		X"CD",X"BA",X"08",X"7E",X"A7",X"28",X"03",X"D6",X"01",X"27",X"77",X"F1",X"E1",X"C9",X"3A",X"44",
		X"40",X"A7",X"C0",X"3A",X"45",X"40",X"E6",X"04",X"C8",X"3A",X"45",X"40",X"E6",X"02",X"C8",X"AF",
		X"37",X"C9",X"C5",X"4F",X"3A",X"45",X"40",X"47",X"E6",X"08",X"20",X"0E",X"78",X"E6",X"01",X"20",
		X"05",X"78",X"E6",X"04",X"20",X"03",X"37",X"18",X"01",X"AF",X"79",X"C1",X"C9",X"F5",X"AF",X"32",
		X"44",X"40",X"3E",X"01",X"CD",X"F0",X"0A",X"3E",X"02",X"20",X"0C",X"CD",X"F0",X"0A",X"20",X"03",
		X"AF",X"18",X"0F",X"3E",X"01",X"18",X"0B",X"CD",X"F0",X"0A",X"20",X"04",X"3E",X"04",X"18",X"02",
		X"3E",X"08",X"32",X"45",X"40",X"3E",X"06",X"CD",X"F0",X"0A",X"28",X"08",X"3A",X"45",X"40",X"F6",
		X"80",X"32",X"45",X"40",X"F1",X"C9",X"E5",X"21",X"45",X"40",X"CB",X"E6",X"CB",X"EE",X"E1",X"C9",
		X"E5",X"21",X"45",X"40",X"CB",X"A6",X"CB",X"AE",X"E1",X"C9",X"E5",X"F5",X"21",X"45",X"40",X"CB",
		X"7E",X"28",X"0C",X"3D",X"E6",X"01",X"28",X"07",X"06",X"02",X"CD",X"2B",X"0B",X"18",X"05",X"06",
		X"01",X"CD",X"35",X"0B",X"F1",X"E1",X"C9",X"C5",X"01",X"02",X"00",X"41",X"21",X"00",X"00",X"19",
		X"7E",X"A7",X"28",X"2F",X"3D",X"4F",X"D5",X"C5",X"21",X"02",X"00",X"19",X"EB",X"01",X"02",X"00",
		X"09",X"01",X"07",X"04",X"78",X"CD",X"DC",X"03",X"C1",X"28",X"17",X"C5",X"06",X"00",X"21",X"CE",
		X"12",X"09",X"09",X"7E",X"23",X"66",X"6F",X"01",X"07",X"04",X"EB",X"CD",X"FC",X"08",X"C1",X"CD",
		X"A8",X"1D",X"D1",X"21",X"48",X"00",X"19",X"EB",X"10",X"C2",X"C1",X"C9",X"F5",X"BE",X"30",X"2F",
		X"C5",X"D5",X"E5",X"EB",X"21",X"00",X"00",X"FD",X"E5",X"C1",X"09",X"4F",X"7E",X"A7",X"28",X"1C",
		X"EB",X"06",X"00",X"09",X"09",X"23",X"4E",X"23",X"46",X"11",X"02",X"00",X"FD",X"E5",X"E1",X"19",
		X"11",X"07",X"04",X"7A",X"54",X"5D",X"CD",X"C1",X"03",X"CD",X"D2",X"10",X"E1",X"D1",X"C1",X"F1",
		X"C9",X"A7",X"C8",X"E5",X"D5",X"C5",X"F5",X"F5",X"0A",X"8E",X"27",X"12",X"03",X"13",X"23",X"E3",
		X"25",X"E3",X"C2",X"C8",X"03",X"E1",X"E1",X"7C",X"C1",X"D1",X"E1",X"C9",X"A7",X"C8",X"E5",X"D5",
		X"C5",X"F5",X"0E",X"00",X"47",X"1A",X"BE",X"28",X"2E",X"0C",X"C5",X"4F",X"46",X"C5",X"E6",X"F0",
		X"4F",X"78",X"E6",X"F0",X"B9",X"C1",X"79",X"28",X"10",X"C6",X"10",X"27",X"4F",X"C5",X"E6",X"0F",
		X"4F",X"78",X"E6",X"0F",X"B9",X"C1",X"79",X"28",X"0C",X"E6",X"F0",X"47",X"79",X"E6",X"0F",X"C6",
		X"01",X"27",X"E6",X"0F",X"B0",X"12",X"C1",X"13",X"23",X"10",X"CA",X"79",X"C1",X"A7",X"78",X"C1",
		X"D1",X"E1",X"C9",X"E5",X"21",X"45",X"40",X"CB",X"F6",X"E1",X"C9",X"E5",X"21",X"45",X"40",X"CB",
		X"B6",X"E1",X"C9",X"F5",X"A7",X"28",X"2C",X"E5",X"D5",X"C5",X"47",X"0E",X"00",X"21",X"8E",X"40",
		X"11",X"02",X"00",X"19",X"C5",X"EB",X"06",X"00",X"21",X"CE",X"12",X"09",X"09",X"7E",X"23",X"66",
		X"6F",X"01",X"07",X"04",X"EB",X"CD",X"FC",X"08",X"11",X"48",X"00",X"19",X"C1",X"0C",X"10",X"E4",
		X"C1",X"D1",X"E1",X"F1",X"C9",X"21",X"3D",X"40",X"34",X"23",X"7E",X"3C",X"FE",X"3C",X"38",X"1C",
		X"36",X"00",X"23",X"7E",X"3C",X"FE",X"3C",X"38",X"13",X"36",X"00",X"23",X"7E",X"3C",X"FE",X"3C",
		X"38",X"0A",X"36",X"00",X"23",X"7E",X"3C",X"FE",X"18",X"38",X"01",X"AF",X"77",X"C9",X"E5",X"F5",
		X"21",X"3D",X"40",X"AF",X"77",X"23",X"77",X"23",X"77",X"23",X"77",X"23",X"77",X"F1",X"E1",X"C9",
		X"21",X"3D",X"40",X"23",X"5E",X"23",X"56",X"23",X"7E",X"23",X"66",X"6F",X"3A",X"3D",X"40",X"C9",
		X"F5",X"C5",X"4F",X"7E",X"A7",X"28",X"38",X"D5",X"E5",X"47",X"23",X"7E",X"23",X"A1",X"BE",X"23",
		X"20",X"08",X"23",X"5E",X"23",X"56",X"23",X"23",X"18",X"09",X"BE",X"20",X"1A",X"23",X"23",X"23",
		X"5E",X"23",X"56",X"23",X"C5",X"4E",X"23",X"46",X"23",X"7E",X"23",X"E5",X"66",X"6F",X"EB",X"CD",
		X"E2",X"0B",X"E1",X"23",X"C1",X"18",X"04",X"11",X"09",X"00",X"19",X"10",X"CE",X"E1",X"D1",X"C1",
		X"F1",X"C9",X"F5",X"7E",X"A7",X"28",X"23",X"C5",X"D5",X"E5",X"47",X"23",X"23",X"23",X"23",X"5E",
		X"23",X"56",X"23",X"23",X"23",X"C5",X"4E",X"23",X"46",X"23",X"7E",X"23",X"E5",X"66",X"6F",X"EB",
		X"CD",X"E2",X"0B",X"E1",X"C1",X"10",X"E4",X"E1",X"D1",X"C1",X"F1",X"C9",X"E5",X"C5",X"4F",X"B7",
		X"CD",X"2C",X"05",X"1F",X"FE",X"64",X"30",X"F8",X"B9",X"C1",X"E1",X"C9",X"E5",X"D5",X"2A",X"48",
		X"40",X"5E",X"23",X"56",X"3E",X"F1",X"CD",X"93",X"05",X"7B",X"C6",X"19",X"5F",X"7A",X"CE",X"36",
		X"77",X"2B",X"73",X"D1",X"E1",X"C9",X"E5",X"2A",X"48",X"40",X"36",X"36",X"23",X"36",X"23",X"E1",
		X"C9",X"E5",X"C5",X"F5",X"42",X"4B",X"11",X"00",X"00",X"CB",X"38",X"79",X"1F",X"4F",X"30",X"03",
		X"EB",X"19",X"EB",X"29",X"B0",X"C2",X"59",X"05",X"F1",X"C1",X"E1",X"C9",X"F5",X"C5",X"7C",X"2F",
		X"47",X"7D",X"2F",X"4F",X"03",X"21",X"00",X"00",X"3E",X"11",X"E5",X"09",X"30",X"01",X"E3",X"E1",
		X"CB",X"13",X"CB",X"12",X"CB",X"15",X"CB",X"14",X"3D",X"C2",X"7A",X"05",X"CB",X"1C",X"CB",X"1D",
		X"C1",X"F1",X"C9",X"E5",X"F5",X"EB",X"11",X"00",X"00",X"B7",X"1F",X"30",X"03",X"EB",X"19",X"EB",
		X"29",X"B7",X"C2",X"9A",X"05",X"F1",X"E1",X"C9",X"E5",X"C5",X"F5",X"FD",X"E5",X"C1",X"21",X"02",
		X"00",X"09",X"EB",X"01",X"07",X"04",X"78",X"01",X"0A",X"00",X"04",X"CD",X"4D",X"00",X"38",X"0E",
		X"D5",X"11",X"09",X"00",X"19",X"D1",X"0D",X"20",X"F2",X"10",X"F0",X"04",X"18",X"2E",X"05",X"0B",
		X"78",X"B1",X"28",X"1B",X"D5",X"E5",X"E5",X"60",X"69",X"11",X"09",X"00",X"CD",X"51",X"05",X"42",
		X"4B",X"D1",X"21",X"09",X"00",X"19",X"09",X"2B",X"EB",X"09",X"2B",X"ED",X"B8",X"E1",X"D1",X"EB",
		X"01",X"07",X"04",X"48",X"06",X"00",X"ED",X"B0",X"CD",X"0B",X"07",X"BF",X"C1",X"78",X"C1",X"E1",
		X"C9",X"E5",X"D5",X"C5",X"2A",X"CC",X"12",X"EB",X"2A",X"46",X"40",X"01",X"07",X"04",X"CD",X"FC",
		X"08",X"C1",X"D1",X"E1",X"C9",X"D5",X"C5",X"F5",X"ED",X"5B",X"46",X"40",X"CD",X"A8",X"05",X"20",
		X"09",X"CD",X"2A",X"03",X"CD",X"1B",X"19",X"CD",X"0B",X"07",X"F1",X"C1",X"D1",X"C9",X"E5",X"D5",
		X"C5",X"F5",X"21",X"04",X"48",X"01",X"FC",X"03",X"CD",X"F9",X"06",X"21",X"00",X"48",X"BE",X"20",
		X"2E",X"01",X"02",X"00",X"21",X"04",X"48",X"06",X"0A",X"11",X"66",X"00",X"79",X"4E",X"B9",X"28",
		X"11",X"0C",X"0D",X"28",X"4B",X"19",X"10",X"F5",X"01",X"00",X"04",X"21",X"00",X"48",X"AF",X"CF",
		X"18",X"28",X"23",X"22",X"46",X"40",X"21",X"02",X"48",X"22",X"48",X"40",X"C3",X"F4",X"06",X"AF",
		X"CD",X"7B",X"0A",X"C6",X"08",X"21",X"00",X"48",X"01",X"05",X"01",X"18",X"05",X"77",X"BE",X"20",
		X"32",X"23",X"10",X"F9",X"0D",X"20",X"F6",X"A7",X"20",X"E6",X"21",X"04",X"48",X"01",X"02",X"00",
		X"71",X"23",X"22",X"46",X"40",X"21",X"02",X"48",X"22",X"48",X"40",X"CD",X"46",X"05",X"18",X"4E",
		X"77",X"23",X"22",X"46",X"40",X"21",X"02",X"48",X"22",X"48",X"40",X"CD",X"36",X"16",X"CD",X"0B",
		X"07",X"18",X"41",X"21",X"84",X"58",X"01",X"66",X"00",X"CD",X"F9",X"06",X"01",X"02",X"00",X"21",
		X"80",X"58",X"BE",X"20",X"14",X"3A",X"84",X"58",X"B9",X"20",X"0E",X"21",X"85",X"58",X"22",X"46",
		X"40",X"21",X"42",X"40",X"22",X"48",X"40",X"18",X"1B",X"21",X"80",X"58",X"06",X"6A",X"AF",X"E7",
		X"21",X"84",X"58",X"71",X"23",X"22",X"46",X"40",X"21",X"42",X"40",X"22",X"48",X"40",X"CD",X"36",
		X"16",X"CD",X"0B",X"07",X"F1",X"C1",X"D1",X"E1",X"C9",X"E5",X"C5",X"3E",X"A5",X"04",X"0C",X"18",
		X"02",X"86",X"23",X"0D",X"20",X"FB",X"10",X"F9",X"C1",X"E1",X"C9",X"E5",X"C5",X"F5",X"2A",X"46",
		X"40",X"01",X"00",X"4C",X"B7",X"ED",X"42",X"21",X"04",X"48",X"01",X"FC",X"03",X"38",X"06",X"21",
		X"84",X"58",X"01",X"66",X"00",X"CD",X"F9",X"06",X"01",X"FC",X"FF",X"09",X"77",X"F1",X"C1",X"E1",
		X"C9",X"2A",X"46",X"40",X"C9",X"E5",X"C5",X"F5",X"01",X"04",X"80",X"21",X"00",X"58",X"AF",X"E7",
		X"06",X"08",X"7C",X"80",X"67",X"0D",X"20",X"F6",X"3E",X"FF",X"ED",X"47",X"77",X"3E",X"20",X"CD",
		X"BD",X"09",X"CD",X"35",X"0B",X"CD",X"73",X"0A",X"CD",X"E1",X"1A",X"CD",X"15",X"08",X"CD",X"13",
		X"0C",X"20",X"D5",X"F1",X"C1",X"E1",X"C9",X"E5",X"C5",X"F5",X"21",X"00",X"40",X"06",X"20",X"AF",
		X"E7",X"3E",X"FC",X"32",X"21",X"40",X"3E",X"1C",X"32",X"20",X"40",X"21",X"22",X"40",X"06",X"10",
		X"AF",X"E7",X"32",X"32",X"40",X"3E",X"FE",X"32",X"34",X"40",X"3E",X"0C",X"32",X"33",X"40",X"F1",
		X"C1",X"E1",X"C9",X"21",X"00",X"40",X"11",X"40",X"58",X"01",X"20",X"00",X"ED",X"B0",X"21",X"22",
		X"40",X"1C",X"ED",X"A0",X"1C",X"ED",X"A0",X"1C",X"ED",X"A0",X"1C",X"ED",X"A0",X"1C",X"ED",X"A0",
		X"1C",X"ED",X"A0",X"1C",X"ED",X"A0",X"1C",X"ED",X"A0",X"1C",X"ED",X"A0",X"1C",X"ED",X"A0",X"1C",
		X"ED",X"A0",X"1C",X"ED",X"A0",X"1C",X"ED",X"A0",X"1C",X"ED",X"A0",X"1C",X"ED",X"A0",X"1C",X"7E",
		X"12",X"C9",X"E5",X"C5",X"F5",X"21",X"20",X"40",X"06",X"00",X"4E",X"3E",X"1C",X"91",X"28",X"11",
		X"CB",X"3F",X"CB",X"3F",X"36",X"1C",X"21",X"04",X"40",X"09",X"0E",X"04",X"70",X"09",X"3D",X"20",
		X"FB",X"3A",X"32",X"40",X"A7",X"20",X"03",X"32",X"30",X"40",X"21",X"33",X"40",X"4E",X"3E",X"0C",
		X"91",X"28",X"0E",X"CB",X"3F",X"36",X"0C",X"21",X"24",X"40",X"09",X"70",X"23",X"23",X"3D",X"20",
		X"FA",X"F1",X"C1",X"E1",X"C9",X"F5",X"3A",X"00",X"78",X"ED",X"57",X"A7",X"20",X"01",X"76",X"CD",
		X"D2",X"07",X"CD",X"E1",X"01",X"F1",X"C9",X"E5",X"D5",X"C5",X"F5",X"CD",X"6C",X"0A",X"CD",X"93",
		X"07",X"CD",X"36",X"02",X"CD",X"C9",X"08",X"CD",X"EC",X"1A",X"CD",X"51",X"08",X"CD",X"73",X"0A",
		X"F1",X"C1",X"D1",X"E1",X"ED",X"45",X"C5",X"4F",X"7B",X"B2",X"A1",X"4F",X"7B",X"A2",X"B1",X"C1",
		X"C9",X"3A",X"3A",X"40",X"5F",X"3A",X"00",X"60",X"57",X"32",X"3A",X"40",X"3A",X"3C",X"40",X"CD",
		X"46",X"08",X"32",X"3C",X"40",X"3A",X"39",X"40",X"5F",X"3A",X"00",X"68",X"57",X"32",X"39",X"40",
		X"3A",X"3B",X"40",X"CD",X"46",X"08",X"32",X"3B",X"40",X"C9",X"E5",X"C5",X"21",X"35",X"40",X"01",
		X"00",X"02",X"78",X"CD",X"16",X"0B",X"28",X"0C",X"7E",X"F6",X"80",X"77",X"FE",X"A1",X"30",X"22",
		X"3C",X"77",X"18",X"1E",X"7E",X"A7",X"28",X"1A",X"CB",X"BE",X"CB",X"7F",X"20",X"14",X"FE",X"02",
		X"38",X"0E",X"FE",X"21",X"30",X"0A",X"0C",X"3A",X"37",X"40",X"3C",X"28",X"03",X"32",X"37",X"40",
		X"36",X"00",X"23",X"10",X"CD",X"79",X"A7",X"C1",X"E1",X"C9",X"F5",X"AF",X"32",X"05",X"70",X"F1",
		X"C9",X"F5",X"3E",X"FF",X"32",X"05",X"70",X"F1",X"C9",X"3A",X"38",X"40",X"A7",X"28",X"19",X"FE",
		X"10",X"38",X"10",X"D6",X"10",X"32",X"38",X"40",X"C0",X"3E",X"04",X"32",X"38",X"40",X"AF",X"32",
		X"03",X"60",X"C9",X"3D",X"32",X"38",X"40",X"C9",X"3A",X"37",X"40",X"A7",X"C8",X"3D",X"32",X"37",
		X"40",X"3E",X"40",X"32",X"38",X"40",X"3E",X"FF",X"32",X"03",X"60",X"C9",X"E5",X"D5",X"C5",X"F5",
		X"79",X"87",X"87",X"87",X"82",X"57",X"78",X"A7",X"79",X"20",X"11",X"A7",X"28",X"61",X"7A",X"C6",
		X"F8",X"57",X"3E",X"30",X"CD",X"CC",X"0B",X"0D",X"28",X"55",X"18",X"3E",X"A7",X"28",X"49",X"7A",
		X"C6",X"F8",X"57",X"7E",X"E6",X"0F",X"C6",X"30",X"CD",X"CC",X"0B",X"0D",X"28",X"3A",X"7A",X"C6",
		X"F8",X"57",X"7E",X"E6",X"F0",X"0F",X"0F",X"0F",X"0F",X"28",X"0F",X"C6",X"30",X"CD",X"CC",X"0B",
		X"0D",X"28",X"29",X"CD",X"75",X"09",X"28",X"12",X"18",X"0D",X"CD",X"75",X"09",X"28",X"0F",X"C6",
		X"30",X"CD",X"CC",X"0B",X"0D",X"28",X"15",X"23",X"10",X"C5",X"7A",X"C6",X"F8",X"57",X"3E",X"20",
		X"CD",X"CC",X"0B",X"0D",X"20",X"F4",X"18",X"07",X"AF",X"BE",X"20",X"03",X"23",X"10",X"F9",X"C1",
		X"78",X"C1",X"D1",X"E1",X"C9",X"E5",X"C5",X"4F",X"AF",X"18",X"04",X"23",X"BE",X"20",X"02",X"10",
		X"FA",X"79",X"C1",X"E1",X"C9",X"E5",X"D5",X"C5",X"4F",X"47",X"87",X"87",X"87",X"82",X"57",X"7A",
		X"D6",X"08",X"57",X"D5",X"EB",X"21",X"0A",X"00",X"CD",X"6C",X"05",X"7D",X"C6",X"30",X"EB",X"D1",
		X"CD",X"CC",X"0B",X"7D",X"B4",X"28",X"04",X"10",X"E6",X"18",X"0D",X"05",X"28",X"0A",X"7A",X"D6",
		X"08",X"57",X"3E",X"20",X"CD",X"CC",X"0B",X"BF",X"79",X"C1",X"D1",X"E1",X"C9",X"E5",X"D5",X"C5",
		X"F5",X"21",X"B2",X"12",X"4F",X"06",X"00",X"09",X"4E",X"21",X"00",X"50",X"71",X"11",X"01",X"50",
		X"01",X"FF",X"03",X"ED",X"B0",X"CD",X"67",X"07",X"F1",X"C1",X"D1",X"E1",X"C9",X"E5",X"D5",X"F5",
		X"C5",X"CB",X"38",X"CB",X"38",X"CB",X"38",X"28",X"7E",X"CB",X"39",X"CB",X"39",X"CB",X"39",X"28",
		X"76",X"D5",X"21",X"B2",X"12",X"85",X"6F",X"30",X"01",X"24",X"7E",X"F5",X"CD",X"AE",X"0B",X"F1",
		X"16",X"00",X"E5",X"59",X"77",X"23",X"1D",X"20",X"FB",X"E1",X"1E",X"20",X"19",X"10",X"F3",X"D1",
		X"3A",X"21",X"40",X"C6",X"04",X"E6",X"3C",X"28",X"4E",X"0F",X"0F",X"C1",X"C5",X"F5",X"78",X"B7",
		X"1F",X"82",X"C6",X"16",X"2F",X"57",X"79",X"B7",X"1F",X"83",X"C6",X"F8",X"5F",X"78",X"C6",X"10",
		X"47",X"79",X"C6",X"10",X"4F",X"21",X"00",X"40",X"F1",X"F5",X"7A",X"96",X"E5",X"6F",X"78",X"CB",
		X"3F",X"85",X"E1",X"23",X"23",X"23",X"B8",X"30",X"19",X"7B",X"96",X"E5",X"6F",X"79",X"CB",X"3F",
		X"85",X"E1",X"B9",X"30",X"0D",X"E5",X"D5",X"C5",X"CD",X"96",X"0E",X"C1",X"D1",X"E1",X"2B",X"2B",
		X"2B",X"2B",X"23",X"F1",X"3D",X"20",X"D2",X"C1",X"F1",X"D1",X"E1",X"C9",X"F5",X"AF",X"32",X"01",
		X"70",X"F1",X"C9",X"F5",X"3E",X"FF",X"32",X"01",X"70",X"F1",X"C9",X"F5",X"3A",X"00",X"78",X"F1",
		X"C9",X"3A",X"3B",X"40",X"E6",X"01",X"20",X"09",X"3A",X"3B",X"40",X"E6",X"02",X"C8",X"3E",X"02",
		X"C9",X"3E",X"01",X"C9",X"F5",X"E5",X"3D",X"20",X"30",X"21",X"D5",X"0A",X"3A",X"3C",X"40",X"57",
		X"A6",X"23",X"20",X"15",X"7A",X"A6",X"20",X"15",X"1E",X"00",X"23",X"7A",X"A6",X"20",X"12",X"23",
		X"7A",X"A6",X"20",X"11",X"16",X"00",X"E1",X"F1",X"C9",X"1E",X"01",X"18",X"ED",X"1E",X"FF",X"18",
		X"E9",X"16",X"01",X"18",X"F1",X"16",X"FF",X"18",X"ED",X"21",X"D9",X"0A",X"3A",X"3B",X"40",X"57",
		X"3A",X"3C",X"40",X"18",X"CB",X"80",X"20",X"08",X"04",X"40",X"20",X"08",X"04",X"3D",X"28",X"08",
		X"3A",X"3B",X"40",X"E6",X"10",X"3E",X"02",X"C9",X"3A",X"3C",X"40",X"E6",X"10",X"3E",X"01",X"C9",
		X"E5",X"C5",X"F5",X"E6",X"07",X"4F",X"FE",X"03",X"30",X"05",X"3A",X"00",X"68",X"18",X"03",X"3A",
		X"00",X"70",X"47",X"79",X"21",X"0E",X"0B",X"D7",X"A0",X"C1",X"78",X"C1",X"E1",X"C9",X"00",X"40",
		X"80",X"01",X"02",X"04",X"08",X"00",X"3D",X"28",X"08",X"3A",X"00",X"60",X"E6",X"02",X"3E",X"02",
		X"C9",X"3A",X"00",X"60",X"E6",X"01",X"3E",X"01",X"C9",X"ED",X"4D",X"F5",X"AF",X"32",X"07",X"70",
		X"32",X"06",X"70",X"F1",X"C9",X"F5",X"3E",X"FF",X"32",X"07",X"70",X"32",X"06",X"70",X"F1",X"C9",
		X"04",X"05",X"C8",X"E5",X"C5",X"67",X"79",X"E6",X"F8",X"0F",X"0F",X"6F",X"7C",X"26",X"58",X"77",
		X"2C",X"2C",X"10",X"FB",X"C1",X"E1",X"C9",X"E5",X"E6",X"F8",X"0F",X"0F",X"6F",X"26",X"58",X"7E",
		X"E1",X"C9",X"E5",X"C5",X"4C",X"21",X"00",X"58",X"06",X"20",X"71",X"23",X"23",X"10",X"FB",X"C1",
		X"E1",X"C9",X"E5",X"C5",X"F5",X"6F",X"26",X"00",X"29",X"01",X"DB",X"15",X"09",X"7E",X"23",X"66",
		X"6F",X"7E",X"CB",X"6F",X"20",X"18",X"D5",X"E6",X"1F",X"3C",X"47",X"16",X"58",X"23",X"7E",X"E6",
		X"F8",X"0F",X"0F",X"3C",X"5F",X"7E",X"E6",X"07",X"12",X"10",X"F2",X"D1",X"18",X"0C",X"E6",X"07",
		X"06",X"20",X"21",X"01",X"58",X"77",X"2C",X"2C",X"10",X"FB",X"F1",X"C1",X"E1",X"C9",X"7A",X"E6",
		X"F8",X"6F",X"26",X"00",X"54",X"29",X"29",X"CB",X"3B",X"CB",X"3B",X"CB",X"3B",X"19",X"11",X"40",
		X"50",X"19",X"C9",X"E5",X"D5",X"CD",X"AE",X"0B",X"7E",X"D1",X"E1",X"C9",X"E5",X"D5",X"F5",X"21",
		X"B2",X"12",X"85",X"6F",X"30",X"01",X"24",X"7E",X"F5",X"CD",X"AE",X"0B",X"F1",X"77",X"F1",X"D1",
		X"E1",X"C9",X"E5",X"D5",X"C5",X"F5",X"AF",X"B9",X"28",X"24",X"B8",X"28",X"21",X"E5",X"CD",X"AE",
		X"0B",X"D1",X"C5",X"E5",X"D5",X"1A",X"11",X"B2",X"12",X"83",X"5F",X"30",X"01",X"14",X"1A",X"77",
		X"11",X"20",X"00",X"19",X"D1",X"13",X"10",X"EC",X"E1",X"23",X"C1",X"0D",X"20",X"E4",X"F1",X"C1",
		X"D1",X"E1",X"C9",X"E5",X"D5",X"C5",X"4F",X"21",X"BC",X"1A",X"46",X"04",X"05",X"28",X"0E",X"23",
		X"5E",X"23",X"56",X"23",X"DD",X"1A",X"A6",X"23",X"BE",X"00",X"00",X"00",X"00",X"AF",X"ED",X"47",
		X"79",X"C1",X"D1",X"E1",X"C9",X"E5",X"D5",X"C5",X"F5",X"29",X"01",X"0D",X"13",X"09",X"4E",X"23",
		X"46",X"0A",X"E6",X"03",X"21",X"4F",X"0C",X"CD",X"3B",X"00",X"F1",X"C1",X"D1",X"E1",X"C9",X"04",
		X"3D",X"0D",X"58",X"0C",X"0F",X"0D",X"F4",X"0C",X"69",X"60",X"23",X"46",X"2B",X"CB",X"7E",X"28",
		X"19",X"78",X"E6",X"07",X"3C",X"4F",X"1F",X"2F",X"3C",X"83",X"5F",X"78",X"E6",X"F8",X"0F",X"0F",
		X"0F",X"3C",X"47",X"1F",X"2F",X"3C",X"82",X"57",X"18",X"0C",X"78",X"CB",X"38",X"CB",X"38",X"CB",
		X"38",X"04",X"E6",X"07",X"3C",X"4F",X"7E",X"23",X"E5",X"E6",X"18",X"0F",X"0F",X"0F",X"EF",X"97",
		X"0C",X"AD",X"0C",X"C4",X"0C",X"DD",X"0C",X"CD",X"AE",X"0B",X"D1",X"13",X"1A",X"16",X"00",X"59",
		X"E5",X"77",X"23",X"1D",X"20",X"FB",X"E1",X"1E",X"20",X"19",X"10",X"F3",X"C9",X"CD",X"AE",X"0B",
		X"D1",X"13",X"1A",X"11",X"20",X"00",X"E5",X"C5",X"77",X"3C",X"19",X"10",X"FB",X"C1",X"E1",X"23",
		X"0D",X"20",X"F3",X"C9",X"CD",X"AE",X"0B",X"D1",X"E5",X"C5",X"13",X"1A",X"77",X"7D",X"C6",X"20",
		X"6F",X"30",X"01",X"24",X"10",X"F4",X"C1",X"E1",X"23",X"0D",X"20",X"EC",X"C9",X"CD",X"AE",X"0B",
		X"D1",X"13",X"1A",X"11",X"E0",X"FF",X"E5",X"C5",X"77",X"3D",X"19",X"10",X"FB",X"C1",X"E1",X"23",
		X"0D",X"20",X"F3",X"C9",X"0A",X"CB",X"7F",X"20",X"02",X"1D",X"1D",X"CB",X"77",X"20",X"01",X"AF",
		X"21",X"32",X"40",X"77",X"2B",X"3E",X"FC",X"93",X"77",X"2B",X"3E",X"F0",X"92",X"77",X"C9",X"21",
		X"33",X"40",X"7E",X"23",X"BE",X"C8",X"0A",X"CB",X"7F",X"28",X"02",X"1D",X"1D",X"CB",X"77",X"28",
		X"06",X"7E",X"C6",X"02",X"77",X"18",X"04",X"2B",X"7E",X"35",X"35",X"21",X"22",X"40",X"85",X"6F",
		X"30",X"01",X"24",X"3E",X"F0",X"92",X"77",X"23",X"3E",X"FC",X"93",X"77",X"C9",X"21",X"20",X"40",
		X"7E",X"23",X"BE",X"C8",X"0A",X"CB",X"7F",X"28",X"09",X"7A",X"D6",X"08",X"57",X"7B",X"D6",X"08",
		X"5F",X"0A",X"CB",X"77",X"28",X"06",X"7E",X"C6",X"04",X"77",X"18",X"07",X"2B",X"7E",X"C6",X"FC",
		X"77",X"C6",X"04",X"21",X"00",X"40",X"85",X"6F",X"30",X"01",X"24",X"7A",X"C6",X"1E",X"2F",X"77",
		X"23",X"03",X"0A",X"77",X"23",X"0B",X"0A",X"E6",X"38",X"0F",X"0F",X"0F",X"77",X"23",X"73",X"C9",
		X"E5",X"D5",X"C5",X"F5",X"29",X"01",X"0D",X"13",X"09",X"4E",X"23",X"46",X"0A",X"E6",X"03",X"21",
		X"9A",X"0D",X"CD",X"3B",X"00",X"F1",X"C1",X"D1",X"E1",X"C9",X"04",X"4B",X"0E",X"A3",X"0D",X"0C",
		X"0E",X"F1",X"0D",X"69",X"60",X"23",X"46",X"2B",X"CB",X"7E",X"28",X"19",X"78",X"E6",X"07",X"3C",
		X"4F",X"1F",X"2F",X"3C",X"83",X"5F",X"78",X"E6",X"F8",X"0F",X"0F",X"0F",X"3C",X"47",X"1F",X"2F",
		X"3C",X"82",X"57",X"18",X"0C",X"78",X"CB",X"38",X"CB",X"38",X"CB",X"38",X"04",X"E6",X"07",X"3C",
		X"4F",X"21",X"B2",X"12",X"7D",X"C6",X"20",X"6F",X"30",X"01",X"24",X"7E",X"F5",X"CD",X"AE",X"0B",
		X"F1",X"16",X"00",X"59",X"E5",X"77",X"23",X"1D",X"20",X"FB",X"E1",X"1E",X"20",X"19",X"10",X"F3",
		X"C9",X"0A",X"E6",X"80",X"28",X"02",X"1D",X"1D",X"21",X"31",X"40",X"3E",X"FC",X"93",X"BE",X"C0",
		X"2B",X"3E",X"F0",X"92",X"96",X"C0",X"77",X"23",X"77",X"23",X"77",X"C9",X"0A",X"E6",X"80",X"28",
		X"02",X"1D",X"1D",X"3A",X"34",X"40",X"4F",X"C6",X"02",X"CB",X"3F",X"C8",X"47",X"3E",X"FC",X"93",
		X"5F",X"3E",X"F0",X"92",X"57",X"21",X"22",X"40",X"BE",X"23",X"28",X"04",X"23",X"10",X"F9",X"C9",
		X"7B",X"BE",X"7A",X"20",X"F7",X"79",X"D6",X"02",X"32",X"34",X"40",X"06",X"00",X"EB",X"21",X"22",
		X"40",X"09",X"7E",X"12",X"70",X"23",X"13",X"7E",X"12",X"70",X"C9",X"69",X"60",X"7A",X"C6",X"1E",
		X"2F",X"57",X"CB",X"7E",X"28",X"07",X"C6",X"08",X"57",X"7B",X"C6",X"F8",X"5F",X"23",X"4E",X"3A",
		X"21",X"40",X"C6",X"04",X"E6",X"FC",X"C8",X"0F",X"0F",X"47",X"2B",X"7E",X"E6",X"38",X"0F",X"0F",
		X"0F",X"F5",X"21",X"00",X"40",X"7A",X"BE",X"23",X"20",X"15",X"79",X"BE",X"20",X"11",X"23",X"7E",
		X"E3",X"BC",X"E3",X"23",X"20",X"0B",X"7B",X"BE",X"20",X"07",X"CD",X"96",X"0E",X"18",X"05",X"23",
		X"23",X"23",X"10",X"E1",X"F1",X"C9",X"EB",X"21",X"21",X"40",X"7E",X"D6",X"04",X"77",X"C6",X"07",
		X"4F",X"06",X"00",X"21",X"00",X"40",X"09",X"0E",X"04",X"ED",X"B8",X"23",X"71",X"C9",X"E5",X"C5",
		X"F5",X"21",X"00",X"00",X"22",X"5F",X"40",X"CD",X"B5",X"12",X"3E",X"01",X"CD",X"37",X"29",X"3E",
		X"00",X"CD",X"58",X"11",X"FD",X"34",X"02",X"CD",X"73",X"2C",X"CD",X"2C",X"05",X"CD",X"AE",X"02",
		X"20",X"33",X"CD",X"24",X"2E",X"CD",X"15",X"08",X"CD",X"AE",X"02",X"20",X"28",X"CD",X"BA",X"21",
		X"3E",X"01",X"CD",X"27",X"17",X"CD",X"09",X"0F",X"21",X"4E",X"10",X"CD",X"F2",X"04",X"0E",X"01",
		X"CD",X"D3",X"10",X"CD",X"AE",X"02",X"20",X"0D",X"CD",X"19",X"10",X"CD",X"AE",X"02",X"20",X"05",
		X"0E",X"01",X"CD",X"D0",X"11",X"F1",X"C1",X"E1",X"C9",X"E5",X"D5",X"C5",X"F5",X"21",X"53",X"0F",
		X"11",X"10",X"18",X"01",X"09",X"16",X"CD",X"E2",X"0B",X"21",X"15",X"58",X"11",X"43",X"0F",X"01",
		X"2C",X"01",X"CD",X"15",X"08",X"79",X"E6",X"1F",X"FE",X"1F",X"20",X"03",X"1A",X"13",X"77",X"CD",
		X"AE",X"02",X"20",X"05",X"0B",X"78",X"B1",X"20",X"E9",X"CD",X"B5",X"12",X"36",X"01",X"F1",X"C1",
		X"D1",X"E1",X"C9",X"02",X"04",X"05",X"01",X"02",X"04",X"05",X"01",X"02",X"04",X"05",X"01",X"02",
		X"04",X"05",X"01",X"44",X"45",X"53",X"49",X"47",X"4E",X"20",X"4C",X"41",X"42",X"53",X"20",X"49",
		X"4E",X"43",X"20",X"21",X"20",X"31",X"39",X"38",X"33",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"50",
		X"48",X"4F",X"4E",X"45",X"20",X"20",X"34",X"30",X"38",X"20",X"20",X"37",X"34",X"38",X"20",X"37",
		X"36",X"30",X"32",X"20",X"20",X"53",X"41",X"4E",X"54",X"41",X"20",X"43",X"4C",X"41",X"52",X"41",
		X"20",X"43",X"41",X"4C",X"49",X"46",X"20",X"20",X"20",X"20",X"20",X"54",X"48",X"4F",X"4D",X"41",
		X"53",X"20",X"41",X"55",X"54",X"4F",X"4D",X"41",X"54",X"49",X"43",X"53",X"20",X"49",X"4E",X"43",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"46",X"4F",X"52",X"20",X"41",X"4D",X"55",X"53",
		X"45",X"4D",X"45",X"4E",X"54",X"20",X"4F",X"4E",X"4C",X"59",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"54",X"52",X"49",X"50",X"4C",X"45",X"20",X"44",X"52",X"41",X"57",
		X"20",X"50",X"4F",X"4B",X"45",X"52",X"20",X"20",X"20",X"E5",X"C5",X"F5",X"06",X"78",X"3E",X"00",
		X"21",X"4E",X"10",X"CD",X"F2",X"04",X"CD",X"15",X"08",X"4F",X"CD",X"AE",X"02",X"20",X"1B",X"79",
		X"3C",X"10",X"F3",X"06",X"78",X"3E",X"00",X"21",X"4E",X"10",X"CD",X"B0",X"04",X"CD",X"15",X"08",
		X"4F",X"CD",X"AE",X"02",X"20",X"04",X"79",X"3C",X"10",X"F0",X"F1",X"C1",X"E1",X"C9",X"01",X"1F",
		X"00",X"0F",X"5A",X"10",X"96",X"10",X"03",X"14",X"40",X"20",X"20",X"20",X"42",X"45",X"20",X"41",
		X"20",X"42",X"49",X"47",X"20",X"57",X"49",X"4E",X"4E",X"45",X"52",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"54",X"52",X"49",X"50",X"4C",X"45",X"20",X"44",X"52",X"41",X"57",X"20",X"50",
		X"4F",X"4B",X"45",X"52",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"C9",X"E5",X"D5",X"C5",X"F5",X"0D",X"28",X"08",X"3E",X"01",X"CD",X"33",X"04",X"CD",
		X"58",X"11",X"3E",X"04",X"CD",X"72",X"0B",X"21",X"44",X"11",X"11",X"40",X"20",X"01",X"01",X"14",
		X"CD",X"E2",X"0B",X"06",X"05",X"11",X"30",X"00",X"CD",X"31",X"07",X"C5",X"01",X"07",X"04",X"CD",
		X"FC",X"08",X"CD",X"B9",X"11",X"01",X"09",X"00",X"09",X"7A",X"C6",X"78",X"57",X"01",X"07",X"04",
		X"CD",X"FC",X"08",X"CD",X"B9",X"11",X"7A",X"D6",X"78",X"57",X"CD",X"81",X"0A",X"20",X"22",X"3E",
		X"2D",X"CD",X"FA",X"26",X"7B",X"D6",X"08",X"5F",X"01",X"09",X"00",X"09",X"C1",X"10",X"CC",X"CD",
		X"81",X"0A",X"20",X"05",X"3E",X"78",X"CD",X"FA",X"26",X"CD",X"E8",X"1A",X"F1",X"C1",X"D1",X"E1",
		X"C9",X"C1",X"18",X"F5",X"41",X"4C",X"4C",X"20",X"54",X"49",X"4D",X"45",X"20",X"48",X"49",X"47",
		X"48",X"20",X"53",X"43",X"4F",X"52",X"45",X"53",X"E5",X"D5",X"C5",X"F5",X"3D",X"28",X"0E",X"3A",
		X"8C",X"40",X"FE",X"02",X"20",X"2C",X"FD",X"E5",X"E1",X"11",X"48",X"00",X"19",X"11",X"02",X"00",
		X"19",X"01",X"07",X"04",X"11",X"E8",X"A0",X"CD",X"FC",X"08",X"21",X"97",X"11",X"11",X"F0",X"A8",
		X"01",X"01",X"06",X"CD",X"E2",X"0B",X"21",X"9D",X"11",X"11",X"F8",X"00",X"01",X"01",X"1C",X"CD",
		X"E2",X"0B",X"F1",X"C1",X"D1",X"E1",X"C9",X"50",X"4F",X"49",X"4E",X"54",X"53",X"50",X"4C",X"41",
		X"59",X"45",X"52",X"20",X"4F",X"4E",X"45",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"50",
		X"4C",X"41",X"59",X"45",X"52",X"20",X"54",X"57",X"4F",X"E5",X"D5",X"C5",X"F5",X"01",X"04",X"00",
		X"09",X"7A",X"C6",X"40",X"57",X"01",X"01",X"05",X"CD",X"E2",X"0B",X"F1",X"C1",X"D1",X"E1",X"C9",
		X"E5",X"C5",X"F5",X"CD",X"B5",X"12",X"CD",X"EA",X"11",X"06",X"78",X"3E",X"00",X"CD",X"B0",X"04",
		X"CD",X"15",X"08",X"3C",X"10",X"F7",X"F1",X"C1",X"E1",X"C9",X"0D",X"21",X"F8",X"11",X"C8",X"3D",
		X"21",X"04",X"12",X"C8",X"21",X"38",X"12",X"C9",X"01",X"1F",X"00",X"0F",X"1B",X"12",X"24",X"12",
		X"01",X"09",X"48",X"40",X"01",X"1F",X"00",X"0F",X"10",X"12",X"24",X"12",X"01",X"14",X"48",X"20",
		X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"4F",X"4E",X"45",X"20",X"47",X"41",X"4D",X"45",X"20",
		X"4F",X"56",X"45",X"52",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"01",X"1F",X"00",X"0F",X"44",X"12",X"24",X"12",
		X"01",X"14",X"48",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"54",X"57",X"4F",X"20",X"47",
		X"41",X"4D",X"45",X"20",X"4F",X"56",X"45",X"52",X"E5",X"D5",X"C5",X"F5",X"04",X"05",X"28",X"03",
		X"CD",X"B5",X"12",X"0C",X"0D",X"20",X"15",X"FE",X"01",X"20",X"11",X"21",X"8A",X"12",X"11",X"48",
		X"28",X"01",X"01",X"12",X"CD",X"E2",X"0B",X"F1",X"C1",X"D1",X"E1",X"C9",X"21",X"9C",X"12",X"11",
		X"48",X"08",X"01",X"01",X"19",X"CD",X"E2",X"0B",X"18",X"ED",X"50",X"52",X"45",X"53",X"53",X"20",
		X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"53",X"54",X"41",X"52",X"54",X"50",X"52",X"45",X"53",
		X"53",X"20",X"31",X"20",X"4F",X"52",X"20",X"32",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",
		X"53",X"54",X"41",X"52",X"54",X"D5",X"C5",X"F5",X"01",X"50",X"E0",X"11",X"08",X"00",X"3E",X"20",
		X"CD",X"DD",X"09",X"CD",X"15",X"08",X"F1",X"C1",X"D1",X"C9",X"00",X"C8",X"E8",X"58",X"E8",X"00",
		X"E8",X"00",X"E7",X"ED",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C3",X"C4",X"C5",X"C6",X"C7",X"C8",X"C9",X"CA",X"CB",X"CC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"CD",X"CE",X"CF",X"D0",X"D1",X"D2",X"D3",X"D4",X"D5",X"D6",X"D7",X"D8",X"D9",
		X"DA",X"DB",X"DC",X"DD",X"DE",X"DF",X"E0",X"E1",X"E2",X"E3",X"E4",X"E5",X"E6",X"7B",X"13",X"A7",
		X"13",X"BB",X"13",X"CF",X"13",X"E3",X"13",X"F7",X"13",X"0B",X"14",X"1F",X"14",X"33",X"14",X"47",
		X"14",X"5B",X"14",X"6F",X"14",X"83",X"14",X"97",X"14",X"91",X"13",X"00",X"00",X"7B",X"13",X"B1",
		X"13",X"C5",X"13",X"D9",X"13",X"ED",X"13",X"01",X"14",X"15",X"14",X"29",X"14",X"3D",X"14",X"51",
		X"14",X"65",X"14",X"79",X"14",X"8D",X"14",X"A1",X"14",X"E3",X"14",X"F7",X"14",X"01",X"15",X"0F",
		X"15",X"1D",X"15",X"29",X"15",X"35",X"15",X"3F",X"15",X"53",X"15",X"5B",X"15",X"6B",X"15",X"7B",
		X"15",X"8B",X"15",X"9B",X"15",X"AB",X"15",X"B7",X"15",X"C3",X"15",X"CF",X"15",X"C7",X"14",X"D5",
		X"14",X"B9",X"14",X"AB",X"14",X"ED",X"14",X"49",X"15",X"63",X"15",X"51",X"1C",X"E7",X"E7",X"E7",
		X"E7",X"E7",X"E7",X"E7",X"E7",X"E7",X"E7",X"E7",X"E7",X"E7",X"E7",X"E7",X"E7",X"E7",X"E7",X"E7",
		X"E7",X"51",X"1C",X"80",X"82",X"82",X"81",X"82",X"82",X"82",X"82",X"83",X"84",X"85",X"86",X"82",
		X"82",X"82",X"82",X"7E",X"82",X"82",X"7F",X"51",X"19",X"05",X"6A",X"6C",X"07",X"00",X"6B",X"6D",
		X"00",X"51",X"19",X"05",X"6E",X"70",X"07",X"00",X"6F",X"71",X"00",X"51",X"19",X"05",X"0A",X"0C",
		X"07",X"00",X"0B",X"0D",X"00",X"51",X"19",X"05",X"0E",X"10",X"07",X"00",X"0F",X"11",X"00",X"51",
		X"19",X"05",X"12",X"3C",X"07",X"00",X"13",X"3D",X"00",X"51",X"19",X"05",X"16",X"40",X"07",X"00",
		X"17",X"41",X"00",X"51",X"19",X"05",X"1A",X"1C",X"07",X"00",X"1B",X"1D",X"00",X"51",X"19",X"05",
		X"1E",X"20",X"07",X"00",X"1F",X"21",X"00",X"51",X"19",X"05",X"22",X"3C",X"07",X"00",X"23",X"25",
		X"00",X"51",X"19",X"05",X"26",X"40",X"07",X"00",X"27",X"29",X"00",X"51",X"19",X"05",X"2A",X"3C",
		X"07",X"00",X"2B",X"2D",X"00",X"51",X"19",X"05",X"2E",X"40",X"07",X"00",X"2F",X"31",X"00",X"51",
		X"19",X"05",X"32",X"34",X"07",X"00",X"33",X"35",X"00",X"51",X"19",X"05",X"36",X"38",X"07",X"00",
		X"37",X"39",X"00",X"51",X"19",X"05",X"3A",X"3C",X"07",X"00",X"3B",X"3D",X"00",X"51",X"19",X"05",
		X"3E",X"40",X"07",X"00",X"3F",X"41",X"00",X"51",X"19",X"05",X"42",X"44",X"07",X"00",X"43",X"45",
		X"00",X"51",X"19",X"05",X"46",X"48",X"07",X"00",X"47",X"49",X"00",X"51",X"19",X"05",X"4A",X"4C",
		X"07",X"00",X"4B",X"4D",X"00",X"51",X"19",X"05",X"4E",X"50",X"07",X"00",X"4F",X"51",X"00",X"51",
		X"19",X"05",X"52",X"54",X"07",X"00",X"53",X"55",X"00",X"51",X"19",X"05",X"56",X"58",X"07",X"00",
		X"57",X"59",X"00",X"51",X"19",X"05",X"5A",X"5C",X"07",X"00",X"5B",X"5D",X"00",X"51",X"19",X"05",
		X"5E",X"60",X"07",X"00",X"5F",X"61",X"00",X"51",X"19",X"05",X"62",X"64",X"07",X"00",X"63",X"65",
		X"00",X"51",X"19",X"05",X"66",X"68",X"07",X"00",X"67",X"69",X"00",X"51",X"1A",X"00",X"00",X"00",
		X"00",X"00",X"72",X"74",X"00",X"06",X"73",X"75",X"08",X"51",X"1A",X"00",X"00",X"00",X"00",X"00",
		X"76",X"78",X"00",X"06",X"77",X"79",X"08",X"51",X"1A",X"00",X"00",X"00",X"00",X"00",X"01",X"02",
		X"00",X"06",X"03",X"04",X"08",X"51",X"1A",X"00",X"00",X"00",X"00",X"00",X"7A",X"7C",X"00",X"06",
		X"7B",X"7D",X"08",X"51",X"19",X"87",X"89",X"8B",X"8D",X"88",X"8A",X"8C",X"8E",X"51",X"19",X"14",
		X"18",X"24",X"30",X"15",X"19",X"28",X"2C",X"51",X"19",X"E8",X"EC",X"EC",X"EA",X"E9",X"EC",X"EC",
		X"EB",X"51",X"29",X"8F",X"91",X"93",X"95",X"97",X"99",X"90",X"92",X"94",X"96",X"98",X"9A",X"51",
		X"29",X"E8",X"EC",X"EC",X"EC",X"EC",X"EA",X"E9",X"EC",X"EC",X"EC",X"EC",X"EB",X"51",X"21",X"9B",
		X"9D",X"9F",X"A1",X"8D",X"9C",X"9E",X"A0",X"A2",X"8E",X"51",X"21",X"E8",X"EC",X"EC",X"EC",X"EA",
		X"E9",X"EC",X"EC",X"EC",X"EB",X"51",X"19",X"A3",X"97",X"91",X"99",X"A4",X"98",X"92",X"9A",X"51",
		X"19",X"E8",X"EC",X"EC",X"EA",X"E9",X"EC",X"EC",X"EB",X"51",X"19",X"F5",X"F1",X"F7",X"F9",X"F6",
		X"F2",X"F8",X"FA",X"51",X"11",X"A5",X"97",X"A7",X"A6",X"98",X"A8",X"51",X"11",X"E8",X"EC",X"EA",
		X"E9",X"EC",X"EB",X"51",X"11",X"EE",X"F1",X"F3",X"EF",X"F2",X"F4",X"51",X"31",X"AD",X"AF",X"B1",
		X"B3",X"B5",X"B7",X"B9",X"AE",X"B0",X"B2",X"B4",X"B6",X"B8",X"BA",X"51",X"31",X"E8",X"EC",X"EC",
		X"EC",X"EC",X"EC",X"EA",X"E9",X"EC",X"EC",X"EC",X"EC",X"EC",X"EB",X"51",X"31",X"8F",X"89",X"A9",
		X"A9",X"97",X"95",X"A7",X"90",X"8A",X"AA",X"AA",X"98",X"96",X"A8",X"51",X"31",X"E8",X"EC",X"EC",
		X"EC",X"EC",X"EC",X"EA",X"E9",X"EC",X"EC",X"EC",X"EC",X"EC",X"EB",X"51",X"21",X"A5",X"8B",X"9F",
		X"AB",X"BB",X"A6",X"8C",X"A0",X"AC",X"BC",X"51",X"21",X"E8",X"EC",X"EC",X"EC",X"EA",X"E9",X"EC",
		X"EC",X"EC",X"EB",X"51",X"21",X"05",X"BD",X"BF",X"C1",X"07",X"06",X"BE",X"C0",X"C2",X"08",X"51",
		X"21",X"E8",X"EC",X"EC",X"EC",X"EA",X"E9",X"EC",X"EC",X"EC",X"EB",X"E5",X"15",X"E6",X"15",X"E9",
		X"15",X"F3",X"15",X"F6",X"15",X"21",X"01",X"EA",X"F2",X"08",X"91",X"99",X"A1",X"A9",X"B1",X"B9",
		X"C1",X"C9",X"D1",X"01",X"15",X"1D",X"04",X"11",X"19",X"21",X"29",X"35",X"E5",X"D5",X"C5",X"F5",
		X"3E",X"20",X"CD",X"BD",X"09",X"CD",X"25",X"16",X"CD",X"61",X"16",X"CD",X"16",X"03",X"21",X"1F",
		X"16",X"01",X"01",X"06",X"11",X"00",X"90",X"CD",X"E2",X"0B",X"F1",X"C1",X"D1",X"E1",X"C9",X"43",
		X"52",X"45",X"44",X"49",X"54",X"F5",X"3E",X"05",X"CD",X"F0",X"0A",X"3E",X"05",X"28",X"02",X"3E",
		X"0A",X"32",X"4A",X"40",X"F1",X"C9",X"E5",X"D5",X"C5",X"F5",X"3E",X"0A",X"CD",X"31",X"07",X"EB",
		X"21",X"58",X"16",X"01",X"04",X"00",X"ED",X"B0",X"21",X"5C",X"16",X"01",X"05",X"00",X"ED",X"B0",
		X"3D",X"20",X"ED",X"F1",X"C1",X"D1",X"E1",X"C9",X"00",X"50",X"00",X"00",X"50",X"4F",X"4B",X"45",
		X"52",X"F5",X"3E",X"00",X"CD",X"72",X"0B",X"CD",X"77",X"16",X"CD",X"EB",X"16",X"3E",X"00",X"CD",
		X"27",X"17",X"CD",X"58",X"18",X"F1",X"C9",X"E5",X"D5",X"C5",X"F5",X"3E",X"01",X"CD",X"72",X"0B",
		X"11",X"F0",X"08",X"21",X"9D",X"16",X"01",X"01",X"1A",X"CD",X"E2",X"0B",X"CD",X"D1",X"16",X"FD",
		X"7E",X"37",X"CD",X"33",X"04",X"CD",X"B7",X"16",X"F1",X"C1",X"D1",X"E1",X"C9",X"50",X"4F",X"49",
		X"4E",X"54",X"53",X"20",X"20",X"20",X"42",X"45",X"53",X"54",X"20",X"47",X"41",X"4D",X"45",X"20",
		X"20",X"20",X"48",X"41",X"4E",X"44",X"53",X"E5",X"D5",X"C5",X"CD",X"01",X"06",X"CD",X"31",X"07",
		X"01",X"04",X"00",X"09",X"11",X"E0",X"60",X"01",X"01",X"05",X"CD",X"E2",X"0B",X"C1",X"D1",X"E1",
		X"C9",X"E5",X"D5",X"F5",X"FD",X"E5",X"E1",X"11",X"01",X"00",X"19",X"6E",X"26",X"00",X"23",X"11",
		X"E8",X"B8",X"3E",X"02",X"CD",X"85",X"09",X"F1",X"D1",X"E1",X"C9",X"E5",X"D5",X"C5",X"F5",X"FD",
		X"E5",X"E1",X"11",X"06",X"00",X"19",X"06",X"24",X"3E",X"00",X"77",X"23",X"10",X"FC",X"F1",X"C1",
		X"D1",X"E1",X"C9",X"01",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"07",
		X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"70",
		X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"E5",X"D5",X"C5",X"F5",X"CD",X"31",X"18",X"4F",X"3E",
		X"02",X"CD",X"72",X"0B",X"FD",X"7E",X"2A",X"FE",X"09",X"20",X"02",X"0E",X"00",X"79",X"FD",X"E5",
		X"E1",X"01",X"2A",X"00",X"09",X"4E",X"06",X"00",X"11",X"90",X"08",X"21",X"51",X"17",X"C3",X"3B",
		X"00",X"02",X"56",X"17",X"E2",X"17",X"01",X"09",X"0E",X"21",X"64",X"17",X"CD",X"E2",X"0B",X"F1",
		X"C1",X"D1",X"E1",X"C9",X"50",X"41",X"49",X"52",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"32",X"20",X"50",X"41",X"49",X"52",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"33",X"20",X"4F",X"46",X"20",X"41",X"20",X"4B",X"49",X"4E",X"44",X"20",X"20",X"20",X"53",X"54",
		X"52",X"41",X"49",X"47",X"48",X"54",X"20",X"20",X"20",X"20",X"20",X"20",X"46",X"4C",X"55",X"53",
		X"48",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"46",X"55",X"4C",X"4C",X"20",X"48",
		X"4F",X"55",X"53",X"45",X"20",X"20",X"20",X"20",X"34",X"20",X"4F",X"46",X"20",X"41",X"20",X"4B",
		X"49",X"4E",X"44",X"20",X"20",X"20",X"53",X"54",X"52",X"41",X"49",X"47",X"48",X"54",X"20",X"46",
		X"4C",X"55",X"53",X"48",X"52",X"4F",X"59",X"41",X"4C",X"20",X"46",X"4C",X"55",X"53",X"48",X"20",
		X"20",X"20",X"21",X"64",X"17",X"78",X"B9",X"C5",X"CC",X"23",X"18",X"01",X"01",X"0E",X"CD",X"E2",
		X"0B",X"01",X"0E",X"00",X"09",X"47",X"3E",X"08",X"83",X"5F",X"78",X"C1",X"3C",X"FE",X"09",X"20",
		X"E5",X"79",X"FE",X"09",X"CA",X"5F",X"17",X"21",X"10",X"18",X"CD",X"3B",X"00",X"C3",X"5F",X"17",
		X"09",X"DB",X"1D",X"0D",X"1E",X"55",X"1E",X"AA",X"1E",X"06",X"1F",X"68",X"1F",X"D2",X"1F",X"44",
		X"20",X"BD",X"20",X"E5",X"F5",X"79",X"87",X"21",X"25",X"58",X"85",X"6F",X"36",X"00",X"F1",X"E1",
		X"C9",X"E5",X"D5",X"C5",X"F5",X"3E",X"09",X"11",X"90",X"A0",X"FD",X"E5",X"E1",X"01",X"06",X"00",
		X"09",X"01",X"07",X"04",X"CD",X"FC",X"08",X"47",X"3E",X"08",X"83",X"5F",X"78",X"01",X"04",X"00",
		X"3D",X"20",X"ED",X"F1",X"C1",X"D1",X"E1",X"C9",X"E5",X"D5",X"C5",X"F5",X"FD",X"E5",X"E1",X"01",
		X"2B",X"00",X"09",X"11",X"60",X"10",X"06",X"05",X"CD",X"77",X"18",X"3E",X"28",X"82",X"57",X"23",
		X"10",X"F6",X"F1",X"C1",X"D1",X"E1",X"C9",X"E5",X"D5",X"C5",X"F5",X"7E",X"47",X"E6",X"0F",X"4F",
		X"78",X"E6",X"20",X"0F",X"B1",X"6F",X"26",X"00",X"CD",X"35",X"0C",X"3E",X"00",X"B1",X"28",X"17",
		X"FE",X"0E",X"28",X"13",X"21",X"30",X"00",X"78",X"E6",X"30",X"0F",X"0F",X"0F",X"0F",X"85",X"6F",
		X"3E",X"10",X"83",X"5F",X"CD",X"35",X"0C",X"F1",X"C1",X"D1",X"E1",X"C9",X"E5",X"D5",X"C5",X"F5",
		X"CD",X"A0",X"04",X"3E",X"05",X"85",X"5F",X"D6",X"3C",X"38",X"03",X"24",X"18",X"01",X"7B",X"6F",
		X"22",X"8A",X"40",X"F1",X"C1",X"D1",X"E1",X"C9",X"E5",X"D5",X"C5",X"F5",X"CD",X"A0",X"04",X"ED",
		X"5B",X"8A",X"40",X"97",X"ED",X"52",X"38",X"01",X"AF",X"C1",X"78",X"C1",X"D1",X"E1",X"C9",X"FD",
		X"E5",X"E5",X"D5",X"C5",X"F5",X"CD",X"FC",X"15",X"CD",X"15",X"08",X"79",X"32",X"8C",X"40",X"CD",
		X"EB",X"16",X"FD",X"E5",X"E1",X"11",X"02",X"00",X"19",X"EB",X"21",X"17",X"19",X"01",X"04",X"00",
		X"ED",X"B0",X"11",X"48",X"00",X"FD",X"19",X"3D",X"CD",X"15",X"08",X"20",X"E2",X"CD",X"23",X"04",
		X"F1",X"C1",X"D1",X"E1",X"FD",X"E1",X"C9",X"10",X"00",X"00",X"00",X"E5",X"D5",X"C5",X"F5",X"CD",
		X"39",X"21",X"CD",X"AC",X"18",X"FD",X"70",X"32",X"CD",X"B5",X"12",X"CD",X"63",X"19",X"EB",X"CD",
		X"11",X"1A",X"11",X"18",X"50",X"3E",X"05",X"01",X"75",X"1A",X"CD",X"C8",X"18",X"28",X"1C",X"CD",
		X"39",X"21",X"CD",X"20",X"1A",X"CD",X"2D",X"1A",X"CD",X"90",X"1A",X"CD",X"15",X"08",X"28",X"EA",
		X"3D",X"20",X"E4",X"3E",X"3C",X"CD",X"FA",X"26",X"CD",X"B5",X"12",X"CD",X"0B",X"07",X"F1",X"C1",
		X"D1",X"E1",X"C9",X"E5",X"D5",X"C5",X"F5",X"0D",X"28",X"12",X"21",X"FD",X"19",X"3D",X"28",X"03",
		X"21",X"07",X"1A",X"11",X"50",X"48",X"01",X"01",X"0A",X"CD",X"E2",X"0B",X"21",X"8D",X"19",X"11",
		X"28",X"00",X"01",X"04",X"1C",X"CD",X"E2",X"0B",X"F1",X"C1",X"D1",X"E1",X"C9",X"54",X"48",X"45",
		X"20",X"4A",X"4F",X"59",X"53",X"54",X"49",X"43",X"4B",X"20",X"41",X"4E",X"44",X"20",X"46",X"49",
		X"52",X"45",X"20",X"42",X"55",X"54",X"54",X"4F",X"4E",X"45",X"4E",X"54",X"45",X"52",X"20",X"59",
		X"4F",X"55",X"52",X"20",X"4E",X"41",X"4D",X"45",X"20",X"55",X"53",X"49",X"4E",X"47",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"41",X"20",X"4E",X"45",X"57",X"20",X"48",X"49",X"47",X"48",X"20",
		X"53",X"43",X"4F",X"52",X"45",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"43",X"4F",X"4E",X"47",X"52",X"41",X"54",X"55",X"4C",X"41",X"54",X"49",X"4F",X"4E",X"53",
		X"20",X"59",X"4F",X"55",X"52",X"53",X"20",X"49",X"53",X"20",X"20",X"20",X"20",X"50",X"4C",X"41",
		X"59",X"45",X"52",X"20",X"4F",X"4E",X"45",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"54",X"57",
		X"4F",X"E5",X"C5",X"06",X"04",X"0E",X"20",X"71",X"10",X"FD",X"CD",X"0B",X"07",X"C1",X"E1",X"C9",
		X"C5",X"F5",X"0A",X"77",X"01",X"01",X"01",X"CD",X"E2",X"0B",X"F1",X"C1",X"C9",X"E5",X"D5",X"F5",
		X"3E",X"00",X"FD",X"B6",X"34",X"28",X"05",X"FD",X"35",X"34",X"18",X"27",X"FD",X"7E",X"32",X"CD",
		X"94",X"0A",X"3E",X"00",X"B2",X"28",X"1C",X"CD",X"53",X"1D",X"CD",X"AC",X"18",X"CD",X"0B",X"07",
		X"FD",X"36",X"34",X"14",X"15",X"28",X"10",X"0B",X"C5",X"E1",X"11",X"75",X"1A",X"DF",X"30",X"03",
		X"01",X"8F",X"1A",X"F1",X"D1",X"E1",X"C9",X"03",X"C5",X"E1",X"11",X"8F",X"1A",X"DF",X"38",X"F3",
		X"01",X"75",X"1A",X"18",X"EE",X"41",X"42",X"43",X"44",X"45",X"46",X"47",X"48",X"49",X"4A",X"4B",
		X"4C",X"4D",X"4E",X"4F",X"50",X"51",X"52",X"53",X"54",X"55",X"56",X"57",X"58",X"59",X"5A",X"20",
		X"C5",X"F5",X"3E",X"00",X"FD",X"B6",X"35",X"28",X"06",X"FD",X"35",X"35",X"AF",X"18",X"19",X"FD",
		X"7E",X"32",X"CD",X"DD",X"0A",X"28",X"11",X"CD",X"36",X"1D",X"CD",X"AC",X"18",X"FD",X"36",X"35",
		X"14",X"23",X"F5",X"3E",X"08",X"82",X"57",X"F1",X"C1",X"78",X"C1",X"C9",X"09",X"00",X"2F",X"00",
		X"00",X"40",X"2F",X"3F",X"3F",X"C0",X"2F",X"3F",X"3E",X"80",X"2F",X"3F",X"3D",X"C0",X"2F",X"3F",
		X"3B",X"40",X"2F",X"3F",X"37",X"40",X"2F",X"3F",X"2F",X"80",X"2F",X"3F",X"1F",X"40",X"2F",X"3F",
		X"00",X"F5",X"AF",X"32",X"4B",X"40",X"F1",X"C9",X"CD",X"E1",X"1A",X"C9",X"F5",X"C5",X"01",X"FF",
		X"00",X"3A",X"4B",X"40",X"A7",X"28",X"38",X"D5",X"E5",X"11",X"1E",X"41",X"F5",X"1A",X"13",X"21",
		X"3E",X"1B",X"CD",X"3B",X"00",X"20",X"1F",X"21",X"4B",X"40",X"35",X"F1",X"FE",X"01",X"28",X"17",
		X"1B",X"C5",X"D5",X"6F",X"26",X"00",X"29",X"29",X"4D",X"44",X"6B",X"62",X"23",X"23",X"23",X"23",
		X"ED",X"B0",X"D1",X"C1",X"18",X"04",X"F1",X"13",X"13",X"13",X"3D",X"20",X"CF",X"E1",X"D1",X"79",
		X"32",X"00",X"78",X"78",X"32",X"06",X"68",X"0F",X"32",X"07",X"68",X"C1",X"F1",X"C9",X"0C",X"1F",
		X"1C",X"1F",X"1C",X"1F",X"1C",X"1F",X"1C",X"1F",X"1C",X"1F",X"1C",X"1F",X"1C",X"1F",X"1C",X"1F",
		X"1C",X"1F",X"1C",X"2F",X"1C",X"2F",X"1C",X"D5",X"C5",X"F5",X"4F",X"A7",X"28",X"0B",X"FD",X"7E",
		X"00",X"A7",X"20",X"05",X"21",X"23",X"41",X"18",X"35",X"21",X"1E",X"41",X"3A",X"4B",X"40",X"A7",
		X"28",X"0B",X"47",X"79",X"11",X"04",X"00",X"BE",X"30",X"07",X"19",X"10",X"FA",X"71",X"EB",X"18",
		X"17",X"28",X"1A",X"79",X"EB",X"68",X"26",X"00",X"29",X"29",X"4D",X"44",X"19",X"5D",X"54",X"2B",
		X"13",X"13",X"13",X"ED",X"B8",X"23",X"77",X"EB",X"21",X"4B",X"40",X"34",X"EB",X"23",X"F1",X"C1",
		X"D1",X"C9",X"E5",X"A7",X"28",X"04",X"4F",X"1A",X"18",X"0E",X"13",X"1A",X"FE",X"FF",X"28",X"19",
		X"07",X"07",X"07",X"E6",X"07",X"3C",X"4F",X"1A",X"E6",X"1F",X"21",X"00",X"1C",X"85",X"6F",X"30",
		X"01",X"24",X"0D",X"AF",X"3C",X"79",X"4E",X"06",X"03",X"E1",X"C9",X"E5",X"A7",X"28",X"07",X"3D",
		X"28",X"21",X"4F",X"1A",X"18",X"11",X"13",X"1A",X"FE",X"FF",X"28",X"1A",X"07",X"07",X"07",X"E6",
		X"07",X"21",X"F8",X"1B",X"D7",X"4F",X"1A",X"E6",X"1F",X"21",X"00",X"1C",X"85",X"6F",X"30",X"01",
		X"24",X"79",X"4E",X"06",X"02",X"04",X"E1",X"C9",X"57",X"4C",X"41",X"36",X"2B",X"20",X"15",X"0A",
		X"0C",X"1A",X"27",X"33",X"3E",X"49",X"53",X"5D",X"66",X"6F",X"77",X"7F",X"86",X"8D",X"93",X"99",
		X"9F",X"A5",X"AA",X"AF",X"B3",X"B7",X"BC",X"BF",X"C3",X"C6",X"CA",X"CD",X"D0",X"D2",X"FF",X"EB",
		X"7E",X"23",X"5E",X"23",X"56",X"CD",X"A2",X"1B",X"72",X"2B",X"73",X"2B",X"77",X"EB",X"C9",X"EB",
		X"7E",X"23",X"5E",X"23",X"56",X"CD",X"CB",X"1B",X"72",X"2B",X"73",X"2B",X"77",X"EB",X"C9",X"E5",
		X"D5",X"F5",X"3E",X"00",X"CD",X"57",X"1B",X"11",X"53",X"1C",X"36",X"00",X"23",X"73",X"23",X"72",
		X"F1",X"D1",X"E1",X"C9",X"2C",X"70",X"73",X"B5",X"FF",X"E5",X"D5",X"F5",X"3E",X"03",X"CD",X"57",
		X"1B",X"11",X"6D",X"1C",X"36",X"00",X"23",X"73",X"23",X"72",X"F1",X"D1",X"E1",X"C9",X"60",X"61",
		X"62",X"63",X"7E",X"FF",X"E5",X"D5",X"F5",X"3E",X"03",X"CD",X"57",X"1B",X"11",X"88",X"1C",X"36",
		X"00",X"23",X"73",X"23",X"72",X"F1",X"D1",X"E1",X"C9",X"62",X"63",X"64",X"65",X"7E",X"FF",X"E5",
		X"D5",X"F5",X"3E",X"03",X"CD",X"57",X"1B",X"11",X"A3",X"1C",X"36",X"00",X"23",X"73",X"23",X"72",
		X"F1",X"D1",X"E1",X"C9",X"64",X"65",X"66",X"67",X"7E",X"FF",X"E5",X"D5",X"F5",X"3E",X"03",X"CD",
		X"57",X"1B",X"11",X"BE",X"1C",X"36",X"00",X"23",X"73",X"23",X"72",X"F1",X"D1",X"E1",X"C9",X"66",
		X"67",X"68",X"69",X"7E",X"FF",X"E5",X"D5",X"F5",X"3A",X"4B",X"40",X"B7",X"20",X"0E",X"3E",X"07",
		X"CD",X"57",X"1B",X"11",X"DF",X"1C",X"36",X"00",X"23",X"73",X"23",X"72",X"F1",X"D1",X"E1",X"C9",
		X"FE",X"80",X"82",X"83",X"FF",X"E5",X"D5",X"F5",X"3E",X"02",X"CD",X"57",X"1B",X"11",X"F9",X"1C",
		X"36",X"00",X"23",X"73",X"23",X"72",X"F1",X"D1",X"E1",X"C9",X"40",X"3E",X"40",X"FF",X"E5",X"D5",
		X"F5",X"3E",X"01",X"CD",X"57",X"1B",X"11",X"12",X"1D",X"36",X"00",X"23",X"73",X"23",X"72",X"F1",
		X"D1",X"E1",X"C9",X"9E",X"85",X"86",X"87",X"BE",X"FF",X"E5",X"D5",X"F5",X"3E",X"06",X"CD",X"57",
		X"1B",X"11",X"2D",X"1D",X"36",X"00",X"23",X"73",X"23",X"72",X"F1",X"D1",X"E1",X"C9",X"9E",X"6D",
		X"6C",X"6B",X"6A",X"69",X"68",X"FF",X"E5",X"D5",X"F5",X"3E",X"04",X"CD",X"57",X"1B",X"11",X"4A",
		X"1D",X"36",X"00",X"23",X"73",X"23",X"72",X"F1",X"D1",X"E1",X"C9",X"BE",X"68",X"69",X"6A",X"6B",
		X"6C",X"5E",X"FF",X"E5",X"D5",X"F5",X"3E",X"05",X"CD",X"57",X"1B",X"11",X"67",X"1D",X"36",X"00",
		X"23",X"73",X"23",X"72",X"F1",X"D1",X"E1",X"C9",X"BE",X"8C",X"BE",X"FF",X"E5",X"D5",X"F5",X"3E",
		X"09",X"CD",X"57",X"1B",X"11",X"80",X"1D",X"36",X"00",X"23",X"73",X"23",X"72",X"F1",X"D1",X"E1",
		X"C9",X"A0",X"A1",X"A2",X"A3",X"A4",X"A5",X"A6",X"A7",X"FF",X"E5",X"D5",X"F5",X"3E",X"08",X"CD",
		X"57",X"1B",X"11",X"9E",X"1D",X"36",X"00",X"23",X"73",X"23",X"72",X"F1",X"D1",X"E1",X"C9",X"A7",
		X"A6",X"A5",X"A4",X"A3",X"A2",X"A1",X"A0",X"FF",X"C9",X"E5",X"D5",X"F5",X"CD",X"E8",X"1A",X"3E",
		X"0A",X"CD",X"57",X"1B",X"11",X"C0",X"1D",X"36",X"00",X"23",X"73",X"23",X"72",X"F1",X"D1",X"E1",
		X"C9",X"F4",X"F5",X"F1",X"EE",X"EE",X"F0",X"CC",X"E8",X"E9",X"E5",X"E2",X"E2",X"E4",X"C0",X"E8",
		X"E9",X"E5",X"E2",X"E2",X"E4",X"E2",X"E2",X"C0",X"DE",X"CC",X"FF",X"E5",X"D5",X"F5",X"3E",X"0B",
		X"CD",X"57",X"1B",X"11",X"F2",X"1D",X"36",X"00",X"23",X"73",X"23",X"72",X"01",X"1E",X"00",X"F1",
		X"D1",X"E1",X"C9",X"CC",X"E7",X"E8",X"E9",X"C5",X"E9",X"C5",X"E9",X"E5",X"85",X"E5",X"F1",X"F3",
		X"F4",X"F5",X"F1",X"F3",X"F5",X"F5",X"F0",X"D3",X"D1",X"F5",X"EC",X"D1",X"FF",X"E5",X"D5",X"F5",
		X"3E",X"0B",X"CD",X"57",X"1B",X"11",X"24",X"1E",X"36",X"00",X"23",X"73",X"23",X"72",X"01",X"3C",
		X"00",X"F1",X"D1",X"E1",X"C9",X"CC",X"E7",X"E8",X"E9",X"C5",X"E9",X"C5",X"E9",X"E5",X"85",X"E5",
		X"F1",X"F3",X"F4",X"F5",X"F1",X"F3",X"F5",X"F5",X"F0",X"D3",X"D1",X"F5",X"EC",X"D1",X"E7",X"E8",
		X"E9",X"C5",X"E9",X"C5",X"E9",X"E5",X"85",X"C5",X"EE",X"EC",X"EB",X"EE",X"F1",X"F5",X"F5",X"F3",
		X"F1",X"EE",X"93",X"D3",X"FF",X"E5",X"D5",X"F5",X"3E",X"0B",X"CD",X"57",X"1B",X"11",X"6C",X"1E",
		X"36",X"00",X"23",X"73",X"23",X"72",X"01",X"2D",X"00",X"F1",X"D1",X"E1",X"C9",X"CC",X"E7",X"E8",
		X"E9",X"C5",X"E9",X"C5",X"E9",X"E5",X"85",X"E5",X"F1",X"F3",X"F4",X"F5",X"F1",X"F3",X"F5",X"F5",
		X"F0",X"D3",X"D1",X"F5",X"EC",X"D1",X"E7",X"E8",X"E9",X"C5",X"E9",X"C5",X"E9",X"E5",X"85",X"C5",
		X"EE",X"EC",X"EB",X"EE",X"F1",X"F5",X"F5",X"F3",X"F1",X"EE",X"93",X"D3",X"E7",X"E8",X"E9",X"C5",
		X"E9",X"C5",X"E9",X"E5",X"85",X"E5",X"F1",X"F3",X"F4",X"FF",X"E5",X"D5",X"F5",X"3E",X"0B",X"CD",
		X"57",X"1B",X"11",X"C1",X"1E",X"36",X"00",X"23",X"73",X"23",X"72",X"01",X"64",X"00",X"F1",X"D1",
		X"E1",X"C9",X"CC",X"E7",X"E8",X"E9",X"C5",X"E9",X"C5",X"E9",X"E5",X"85",X"E5",X"F1",X"F3",X"F4",
		X"F5",X"F1",X"F3",X"F5",X"F5",X"F0",X"D3",X"D1",X"F5",X"EC",X"D1",X"E7",X"E8",X"E9",X"C5",X"E9",
		X"C5",X"E9",X"E5",X"85",X"C5",X"EE",X"EC",X"EB",X"EE",X"F1",X"F5",X"F5",X"F3",X"F1",X"EE",X"93",
		X"D3",X"E7",X"E8",X"E9",X"C5",X"E9",X"C5",X"E9",X"E5",X"85",X"E5",X"F1",X"F3",X"F4",X"F5",X"F1",
		X"F3",X"F5",X"F5",X"F0",X"D3",X"FF",X"E5",X"D5",X"F5",X"3E",X"0B",X"CD",X"57",X"1B",X"11",X"1D",
		X"1F",X"36",X"00",X"23",X"73",X"23",X"72",X"01",X"78",X"00",X"F1",X"D1",X"E1",X"C9",X"CC",X"E7",
		X"E8",X"E9",X"C5",X"E9",X"C5",X"E9",X"E5",X"85",X"E5",X"F1",X"F3",X"F4",X"F5",X"F1",X"F3",X"F5",
		X"F5",X"F0",X"D3",X"D1",X"F5",X"EC",X"D1",X"E7",X"E8",X"E9",X"C5",X"E9",X"C5",X"E9",X"E5",X"85",
		X"C5",X"EE",X"EC",X"EB",X"EE",X"F1",X"F5",X"F5",X"F3",X"F1",X"EE",X"93",X"D3",X"E7",X"E8",X"E9",
		X"C5",X"E9",X"C5",X"E9",X"E5",X"85",X"E5",X"F1",X"F3",X"F4",X"F5",X"F1",X"F3",X"F5",X"F5",X"F0",
		X"D3",X"D1",X"E9",X"E0",X"D1",X"F1",X"F3",X"FF",X"E5",X"D5",X"F5",X"3E",X"0B",X"CD",X"57",X"1B",
		X"11",X"7F",X"1F",X"36",X"00",X"23",X"73",X"23",X"72",X"01",X"8C",X"00",X"F1",X"D1",X"E1",X"C9",
		X"CC",X"E7",X"E8",X"E9",X"C5",X"E9",X"C5",X"E9",X"E5",X"85",X"E5",X"F1",X"F3",X"F4",X"F5",X"F1",
		X"F3",X"F5",X"F5",X"F0",X"D3",X"D1",X"F5",X"EC",X"D1",X"E7",X"E8",X"E9",X"C5",X"E9",X"C5",X"E9",
		X"E5",X"85",X"C5",X"EE",X"EC",X"EB",X"EE",X"F1",X"F5",X"F5",X"F3",X"F1",X"EE",X"93",X"D3",X"E7",
		X"E8",X"E9",X"C5",X"E9",X"C5",X"E9",X"E5",X"85",X"E5",X"F1",X"F3",X"F4",X"F5",X"F1",X"F3",X"F5",
		X"F5",X"F0",X"D3",X"D1",X"E9",X"E0",X"D1",X"F1",X"F3",X"F5",X"F1",X"F3",X"F5",X"F5",X"F1",X"F3",
		X"F1",X"FF",X"E5",X"D5",X"F5",X"3E",X"0B",X"CD",X"57",X"1B",X"11",X"E9",X"1F",X"36",X"00",X"23",
		X"73",X"23",X"72",X"01",X"A0",X"00",X"F1",X"D1",X"E1",X"C9",X"CC",X"E7",X"E8",X"E9",X"C5",X"E9",
		X"C5",X"E9",X"E5",X"85",X"E5",X"F1",X"F3",X"F4",X"F5",X"F1",X"F3",X"F5",X"F5",X"F0",X"D3",X"D1",
		X"F5",X"EC",X"D1",X"E7",X"E8",X"E9",X"C5",X"E9",X"C5",X"E9",X"E5",X"85",X"C5",X"EE",X"EC",X"EB",
		X"EE",X"F1",X"F5",X"F5",X"F3",X"F1",X"EE",X"93",X"D3",X"E7",X"E8",X"E9",X"C5",X"E9",X"C5",X"E9",
		X"E5",X"85",X"E5",X"F1",X"F3",X"F4",X"F5",X"F1",X"F3",X"F5",X"F5",X"F0",X"D3",X"D1",X"E9",X"E0",
		X"D1",X"F1",X"F3",X"F5",X"F1",X"F3",X"F5",X"F5",X"F1",X"F3",X"F1",X"F5",X"F1",X"F3",X"F5",X"F5",
		X"F1",X"F3",X"F1",X"FF",X"E5",X"D5",X"F5",X"3E",X"0B",X"CD",X"57",X"1B",X"11",X"5B",X"20",X"36",
		X"00",X"23",X"73",X"23",X"72",X"01",X"B4",X"00",X"F1",X"D1",X"E1",X"C9",X"CC",X"E7",X"E8",X"E9",
		X"C5",X"E9",X"C5",X"E9",X"E5",X"85",X"E5",X"F1",X"F3",X"F4",X"F5",X"F1",X"F3",X"F5",X"F5",X"F0",
		X"D3",X"D1",X"F5",X"EC",X"D1",X"E7",X"E8",X"E9",X"C5",X"E9",X"C5",X"E9",X"E5",X"85",X"C5",X"EE",
		X"EC",X"EB",X"EE",X"F1",X"F5",X"F5",X"F3",X"F1",X"EE",X"93",X"D3",X"E7",X"E8",X"E9",X"C5",X"E9",
		X"C5",X"E9",X"E5",X"85",X"E5",X"F1",X"F3",X"F4",X"F5",X"F1",X"F3",X"F5",X"F5",X"F0",X"D3",X"D1",
		X"E9",X"E0",X"D1",X"F1",X"F3",X"F5",X"F1",X"F3",X"F5",X"F5",X"F1",X"F3",X"F1",X"F5",X"F1",X"F3",
		X"F5",X"F5",X"F1",X"F3",X"F1",X"F5",X"F1",X"F3",X"F5",X"F5",X"F0",X"D3",X"FF",X"E5",X"D5",X"F5",
		X"3E",X"0B",X"CD",X"57",X"1B",X"11",X"D4",X"20",X"36",X"00",X"23",X"73",X"23",X"72",X"01",X"C8",
		X"00",X"F1",X"D1",X"E1",X"C9",X"CC",X"E7",X"E8",X"E9",X"C5",X"E9",X"C5",X"E9",X"E5",X"85",X"E5",
		X"F1",X"F3",X"F4",X"F5",X"F1",X"F3",X"F5",X"F5",X"F0",X"D3",X"D1",X"F5",X"EC",X"D1",X"E7",X"E8",
		X"E9",X"C5",X"E9",X"C5",X"E9",X"E5",X"85",X"C5",X"EE",X"EC",X"EB",X"EE",X"F1",X"F5",X"F5",X"F3",
		X"F1",X"EE",X"93",X"D3",X"E7",X"E8",X"E9",X"C5",X"E9",X"C5",X"E9",X"E5",X"85",X"E5",X"F1",X"F3",
		X"F4",X"F5",X"F1",X"F3",X"F5",X"F5",X"F0",X"D3",X"D1",X"E9",X"E0",X"D1",X"F1",X"F3",X"F5",X"F1",
		X"F3",X"F5",X"F5",X"F1",X"F3",X"F1",X"F5",X"F1",X"F3",X"F5",X"F5",X"F1",X"F3",X"F1",X"F5",X"F1",
		X"F3",X"F5",X"F5",X"F0",X"D3",X"91",X"D1",X"E7",X"FF",X"E5",X"D5",X"F5",X"3A",X"4B",X"40",X"B7",
		X"20",X"0E",X"3E",X"0B",X"CD",X"57",X"1B",X"11",X"53",X"21",X"36",X"00",X"23",X"73",X"23",X"72",
		X"F1",X"D1",X"E1",X"C9",X"D0",X"CC",X"EC",X"F7",X"F5",X"F4",X"F2",X"D0",X"EE",X"EE",X"EB",X"E9",
		X"E7",X"E9",X"EB",X"EE",X"EE",X"F0",X"F2",X"F4",X"D5",X"8E",X"DE",X"CE",X"8E",X"D0",X"F2",X"D0",
		X"F2",X"F0",X"F2",X"D0",X"F7",X"D5",X"F7",X"F5",X"F7",X"F5",X"F0",X"10",X"CE",X"8E",X"D0",X"F2",
		X"D0",X"F2",X"F0",X"D0",X"F0",X"F0",X"CB",X"F0",X"EF",X"F0",X"D2",X"90",X"F0",X"DE",X"EE",X"CE",
		X"8E",X"D0",X"F2",X"D0",X"F2",X"F0",X"F2",X"D0",X"F7",X"D5",X"F7",X"F5",X"F5",X"F7",X"EC",X"8C",
		X"CC",X"F4",X"EC",X"F7",X"D5",X"F7",X"F5",X"F7",X"F5",X"F0",X"F0",X"F2",X"F0",X"EE",X"EE",X"D0",
		X"F0",X"F0",X"CE",X"F0",X"EE",X"EE",X"D0",X"89",X"9E",X"FF",X"CD",X"DC",X"21",X"CD",X"1E",X"22",
		X"CD",X"43",X"22",X"CD",X"A6",X"22",X"CD",X"C0",X"22",X"CD",X"DE",X"22",X"CD",X"EB",X"22",X"CD",
		X"F8",X"22",X"CD",X"CF",X"22",X"CD",X"10",X"23",X"CD",X"23",X"23",X"C9",X"E5",X"D5",X"C5",X"F5",
		X"FD",X"36",X"39",X"00",X"FD",X"36",X"3A",X"00",X"FD",X"36",X"3B",X"00",X"FD",X"36",X"3C",X"00",
		X"FD",X"E5",X"E1",X"01",X"39",X"00",X"09",X"EB",X"FD",X"E5",X"E1",X"01",X"2B",X"00",X"09",X"06",
		X"04",X"7E",X"E6",X"0F",X"4F",X"C5",X"23",X"E5",X"7E",X"E6",X"0F",X"B9",X"20",X"03",X"1A",X"3C",
		X"12",X"23",X"10",X"F4",X"E1",X"C1",X"13",X"10",X"E8",X"F1",X"C1",X"D1",X"E1",X"C9",X"E5",X"C5",
		X"F5",X"FD",X"36",X"3D",X"00",X"FD",X"E5",X"E1",X"01",X"2B",X"00",X"09",X"7E",X"E6",X"F0",X"4F",
		X"06",X"04",X"23",X"7E",X"E6",X"F0",X"B9",X"20",X"06",X"10",X"F7",X"FD",X"36",X"3D",X"FF",X"F1",
		X"C1",X"E1",X"C9",X"E5",X"C5",X"F5",X"FD",X"36",X"3E",X"00",X"FD",X"E5",X"E1",X"01",X"2B",X"00",
		X"09",X"CD",X"79",X"22",X"FE",X"01",X"20",X"0B",X"3E",X"02",X"CD",X"8F",X"22",X"3E",X"01",X"28",
		X"02",X"3E",X"09",X"06",X"04",X"3C",X"FE",X"0E",X"30",X"0B",X"CD",X"8F",X"22",X"20",X"06",X"10",
		X"F4",X"FD",X"36",X"3E",X"FF",X"F1",X"C1",X"E1",X"C9",X"E5",X"C5",X"7E",X"E6",X"0F",X"4F",X"06",
		X"04",X"23",X"7E",X"E6",X"0F",X"B9",X"30",X"01",X"4F",X"10",X"F6",X"79",X"C1",X"E1",X"C9",X"E5",
		X"C5",X"F5",X"06",X"05",X"4F",X"7E",X"E6",X"0F",X"B9",X"28",X"06",X"23",X"10",X"F7",X"3E",X"01",
		X"B7",X"C1",X"78",X"C1",X"E1",X"C9",X"F5",X"FD",X"36",X"2A",X"09",X"3E",X"01",X"CD",X"4A",X"23",
		X"B7",X"28",X"0B",X"FE",X"02",X"3E",X"00",X"20",X"02",X"3E",X"01",X"FD",X"77",X"2A",X"F1",X"C9",
		X"F5",X"3E",X"02",X"CD",X"4A",X"23",X"B7",X"28",X"04",X"FD",X"36",X"2A",X"02",X"F1",X"C9",X"F5",
		X"3E",X"03",X"CD",X"4A",X"23",X"B7",X"28",X"04",X"FD",X"36",X"2A",X"06",X"F1",X"C9",X"F5",X"FD",
		X"7E",X"3E",X"3C",X"20",X"04",X"FD",X"36",X"2A",X"03",X"F1",X"C9",X"F5",X"FD",X"7E",X"3D",X"3C",
		X"20",X"04",X"FD",X"36",X"2A",X"04",X"F1",X"C9",X"F5",X"3E",X"02",X"CD",X"4A",X"23",X"B7",X"28",
		X"0D",X"3E",X"01",X"CD",X"4A",X"23",X"FE",X"02",X"20",X"04",X"FD",X"36",X"2A",X"05",X"F1",X"C9",
		X"F5",X"FD",X"7E",X"3E",X"3C",X"20",X"0A",X"FD",X"7E",X"3D",X"3C",X"20",X"04",X"FD",X"36",X"2A",
		X"07",X"F1",X"C9",X"E5",X"C5",X"F5",X"FD",X"7E",X"2A",X"FE",X"07",X"20",X"19",X"FD",X"E5",X"E1",
		X"01",X"2B",X"00",X"09",X"3E",X"01",X"CD",X"8F",X"22",X"20",X"0B",X"3E",X"0D",X"CD",X"8F",X"22",
		X"20",X"04",X"FD",X"36",X"2A",X"08",X"F1",X"C1",X"E1",X"C9",X"E5",X"C5",X"FD",X"E5",X"E1",X"01",
		X"39",X"00",X"09",X"01",X"00",X"04",X"BE",X"20",X"01",X"0C",X"23",X"10",X"F9",X"79",X"C1",X"E1",
		X"C9",X"E5",X"D5",X"C5",X"F5",X"CD",X"AC",X"18",X"21",X"D0",X"23",X"11",X"E4",X"23",X"01",X"14",
		X"00",X"CD",X"28",X"2A",X"CD",X"4F",X"2A",X"3E",X"08",X"32",X"8D",X"40",X"FD",X"36",X"36",X"00",
		X"FD",X"36",X"40",X"00",X"FD",X"36",X"33",X"00",X"FD",X"36",X"46",X"00",X"3E",X"00",X"CD",X"C8",
		X"18",X"28",X"23",X"CD",X"88",X"2A",X"CD",X"F0",X"2A",X"CD",X"7B",X"28",X"20",X"06",X"21",X"BB",
		X"23",X"CD",X"EF",X"2B",X"CD",X"15",X"08",X"3C",X"67",X"CD",X"2C",X"05",X"7C",X"FD",X"6E",X"36",
		X"2C",X"20",X"DB",X"CD",X"25",X"2C",X"F1",X"C1",X"D1",X"E1",X"C9",X"0A",X"4A",X"24",X"77",X"24",
		X"A4",X"24",X"D1",X"24",X"FE",X"24",X"2B",X"25",X"49",X"24",X"70",X"25",X"49",X"24",X"24",X"2E",
		X"F8",X"A8",X"1E",X"00",X"1E",X"00",X"1E",X"00",X"1E",X"00",X"1E",X"00",X"20",X"00",X"22",X"00",
		X"24",X"00",X"00",X"00",X"F9",X"23",X"03",X"24",X"0D",X"24",X"17",X"24",X"21",X"24",X"2B",X"24",
		X"F8",X"23",X"35",X"24",X"F8",X"23",X"3F",X"24",X"00",X"01",X"0F",X"00",X"09",X"1E",X"00",X"1F",
		X"00",X"40",X"10",X"01",X"0F",X"00",X"09",X"1E",X"00",X"1F",X"00",X"40",X"38",X"01",X"0F",X"00",
		X"09",X"1E",X"00",X"1F",X"00",X"40",X"60",X"01",X"0F",X"00",X"09",X"1E",X"00",X"1F",X"00",X"40",
		X"88",X"01",X"0F",X"00",X"09",X"1E",X"00",X"1F",X"00",X"40",X"B0",X"01",X"0F",X"00",X"09",X"20",
		X"00",X"21",X"00",X"28",X"10",X"01",X"0F",X"00",X"09",X"22",X"00",X"23",X"00",X"28",X"60",X"01",
		X"0F",X"00",X"09",X"24",X"00",X"25",X"00",X"28",X"B0",X"C9",X"E5",X"F5",X"3E",X"01",X"FD",X"B6",
		X"3F",X"FD",X"77",X"3F",X"FD",X"36",X"41",X"00",X"21",X"34",X"00",X"22",X"61",X"40",X"21",X"6D",
		X"24",X"22",X"75",X"40",X"CD",X"4F",X"2A",X"CD",X"36",X"1D",X"F1",X"E1",X"C9",X"01",X"0F",X"00",
		X"09",X"34",X"00",X"1F",X"00",X"40",X"10",X"E5",X"F5",X"3E",X"02",X"FD",X"B6",X"3F",X"FD",X"77",
		X"3F",X"FD",X"36",X"41",X"00",X"21",X"34",X"00",X"22",X"63",X"40",X"21",X"9A",X"24",X"22",X"77",
		X"40",X"CD",X"4F",X"2A",X"CD",X"36",X"1D",X"F1",X"E1",X"C9",X"01",X"0F",X"00",X"09",X"34",X"00",
		X"1F",X"00",X"40",X"38",X"E5",X"F5",X"3E",X"04",X"FD",X"B6",X"3F",X"FD",X"77",X"3F",X"FD",X"36",
		X"41",X"00",X"21",X"34",X"00",X"22",X"65",X"40",X"21",X"C7",X"24",X"22",X"79",X"40",X"CD",X"4F",
		X"2A",X"CD",X"36",X"1D",X"F1",X"E1",X"C9",X"01",X"0F",X"00",X"09",X"34",X"00",X"1F",X"00",X"40",
		X"60",X"E5",X"F5",X"3E",X"08",X"FD",X"B6",X"3F",X"FD",X"77",X"3F",X"FD",X"36",X"41",X"00",X"21",
		X"34",X"00",X"22",X"67",X"40",X"21",X"F4",X"24",X"22",X"7B",X"40",X"CD",X"4F",X"2A",X"CD",X"36",
		X"1D",X"F1",X"E1",X"C9",X"01",X"0F",X"00",X"09",X"34",X"00",X"1F",X"00",X"40",X"88",X"E5",X"F5",
		X"3E",X"10",X"FD",X"B6",X"3F",X"FD",X"77",X"3F",X"FD",X"36",X"41",X"00",X"21",X"34",X"00",X"22",
		X"69",X"40",X"21",X"21",X"25",X"22",X"7D",X"40",X"CD",X"4F",X"2A",X"CD",X"36",X"1D",X"F1",X"E1",
		X"C9",X"01",X"0F",X"00",X"09",X"34",X"00",X"1F",X"00",X"40",X"B0",X"E5",X"D5",X"C5",X"21",X"5C",
		X"25",X"11",X"61",X"40",X"01",X"0A",X"00",X"ED",X"B0",X"21",X"66",X"25",X"11",X"75",X"40",X"01",
		X"0A",X"00",X"ED",X"B0",X"FD",X"36",X"3F",X"00",X"FD",X"7E",X"47",X"3C",X"20",X"04",X"FD",X"36",
		X"41",X"FF",X"CD",X"4F",X"2A",X"CD",X"53",X"1D",X"C1",X"D1",X"E1",X"C9",X"1E",X"00",X"1E",X"00",
		X"1E",X"00",X"1E",X"00",X"1E",X"00",X"F9",X"23",X"03",X"24",X"0D",X"24",X"17",X"24",X"21",X"24",
		X"FD",X"36",X"3F",X"1F",X"FD",X"36",X"36",X"FF",X"FD",X"36",X"41",X"00",X"C9",X"F5",X"FD",X"7E",
		X"2A",X"FE",X"09",X"C4",X"88",X"25",X"F1",X"C9",X"E5",X"D5",X"C5",X"F5",X"CD",X"AC",X"18",X"CD",
		X"BB",X"27",X"FD",X"36",X"36",X"00",X"FD",X"36",X"33",X"01",X"FD",X"36",X"46",X"00",X"21",X"E5",
		X"25",X"11",X"ED",X"25",X"01",X"08",X"00",X"CD",X"28",X"2A",X"CD",X"4F",X"2A",X"3E",X"00",X"CD",
		X"C8",X"18",X"28",X"23",X"CD",X"88",X"2A",X"CD",X"F0",X"2A",X"CD",X"7B",X"28",X"20",X"06",X"21",
		X"DC",X"25",X"CD",X"EF",X"2B",X"CD",X"15",X"08",X"3C",X"67",X"CD",X"2C",X"05",X"7C",X"FD",X"6E",
		X"36",X"2C",X"20",X"DB",X"CD",X"25",X"2C",X"F1",X"C1",X"D1",X"E1",X"C9",X"04",X"0A",X"26",X"10",
		X"26",X"0A",X"26",X"0B",X"26",X"50",X"00",X"28",X"00",X"2A",X"00",X"00",X"00",X"F5",X"25",X"F6",
		X"25",X"F5",X"25",X"00",X"26",X"00",X"01",X"0F",X"00",X"09",X"28",X"00",X"29",X"00",X"40",X"38",
		X"01",X"0F",X"00",X"09",X"2A",X"00",X"2B",X"00",X"40",X"88",X"C9",X"FD",X"36",X"36",X"FF",X"C9",
		X"E5",X"D5",X"C5",X"F5",X"CD",X"AC",X"18",X"CD",X"9D",X"26",X"CD",X"25",X"2C",X"CD",X"CA",X"26",
		X"21",X"79",X"26",X"11",X"81",X"26",X"01",X"08",X"00",X"CD",X"28",X"2A",X"CD",X"4F",X"2A",X"FD",
		X"36",X"33",X"01",X"FD",X"36",X"36",X"00",X"FD",X"36",X"46",X"00",X"3E",X"00",X"CD",X"C8",X"18",
		X"28",X"29",X"CD",X"88",X"2A",X"CD",X"F0",X"2A",X"CD",X"7B",X"28",X"20",X"06",X"21",X"70",X"26",
		X"CD",X"EF",X"2B",X"CD",X"15",X"08",X"3C",X"67",X"CD",X"2C",X"05",X"7C",X"FD",X"6E",X"36",X"2C",
		X"20",X"DB",X"CD",X"25",X"2C",X"CD",X"B3",X"26",X"CD",X"58",X"18",X"F1",X"C1",X"D1",X"E1",X"C9",
		X"04",X"0A",X"26",X"03",X"27",X"0A",X"26",X"0B",X"27",X"50",X"00",X"2E",X"00",X"2C",X"00",X"00",
		X"00",X"F5",X"25",X"89",X"26",X"F5",X"25",X"93",X"26",X"01",X"0F",X"00",X"09",X"2E",X"00",X"2F",
		X"00",X"40",X"38",X"01",X"0F",X"00",X"09",X"2C",X"00",X"2D",X"00",X"40",X"88",X"E5",X"D5",X"C5",
		X"FD",X"E5",X"E1",X"11",X"2B",X"00",X"19",X"11",X"4D",X"40",X"01",X"05",X"00",X"ED",X"B0",X"C1",
		X"D1",X"E1",X"C9",X"E5",X"D5",X"C5",X"FD",X"E5",X"E1",X"11",X"2B",X"00",X"19",X"EB",X"21",X"4D",
		X"40",X"01",X"05",X"00",X"ED",X"B0",X"C1",X"D1",X"E1",X"C9",X"C5",X"F5",X"FD",X"7E",X"3F",X"FD",
		X"36",X"3F",X"00",X"CD",X"59",X"2E",X"FD",X"77",X"3F",X"FD",X"36",X"2D",X"0E",X"CD",X"58",X"18",
		X"CD",X"2C",X"05",X"4F",X"E6",X"0F",X"28",X"F8",X"FE",X"0E",X"30",X"F4",X"79",X"E6",X"3F",X"CD",
		X"D4",X"2E",X"28",X"EC",X"FD",X"77",X"2D",X"F1",X"C1",X"C9",X"F5",X"CD",X"15",X"08",X"3D",X"20",
		X"FA",X"F1",X"C9",X"F5",X"3E",X"00",X"CD",X"13",X"27",X"F1",X"C9",X"F5",X"3E",X"20",X"CD",X"13",
		X"27",X"F1",X"C9",X"F5",X"CD",X"58",X"18",X"CD",X"2B",X"27",X"3E",X"78",X"CD",X"88",X"2A",X"CD",
		X"15",X"08",X"3D",X"20",X"F7",X"FD",X"36",X"36",X"FF",X"F1",X"C9",X"E5",X"D5",X"C5",X"F5",X"4F",
		X"FD",X"7E",X"2D",X"E6",X"20",X"B9",X"FD",X"E5",X"E1",X"11",X"42",X"00",X"19",X"28",X"1B",X"06",
		X"04",X"36",X"00",X"23",X"10",X"FB",X"21",X"74",X"27",X"11",X"28",X"50",X"01",X"01",X"08",X"CD",
		X"E2",X"0B",X"CD",X"8A",X"1D",X"F1",X"C1",X"D1",X"E1",X"C9",X"44",X"4D",X"54",X"5D",X"3E",X"04",
		X"CD",X"C1",X"03",X"21",X"7C",X"27",X"11",X"28",X"40",X"01",X"01",X"0B",X"CD",X"E2",X"0B",X"CD",
		X"6C",X"1D",X"18",X"E1",X"57",X"49",X"4E",X"20",X"4C",X"4F",X"53",X"54",X"57",X"49",X"4E",X"20",
		X"44",X"4F",X"55",X"42",X"4C",X"45",X"44",X"E5",X"D5",X"C5",X"F5",X"FD",X"7E",X"2A",X"FE",X"09",
		X"28",X"13",X"FD",X"E5",X"E1",X"11",X"42",X"00",X"19",X"E5",X"3E",X"00",X"06",X"04",X"BE",X"23",
		X"20",X"08",X"10",X"FA",X"E1",X"F1",X"C1",X"D1",X"E1",X"C9",X"FD",X"E5",X"E1",X"01",X"02",X"00",
		X"09",X"C1",X"54",X"5D",X"3E",X"04",X"CD",X"C1",X"03",X"18",X"EA",X"E5",X"D5",X"C5",X"F5",X"FD",
		X"E5",X"E1",X"11",X"42",X"00",X"19",X"EB",X"FD",X"E5",X"E1",X"01",X"06",X"00",X"09",X"FD",X"7E",
		X"2A",X"07",X"07",X"4F",X"06",X"00",X"09",X"01",X"04",X"00",X"ED",X"B0",X"F1",X"C1",X"D1",X"E1",
		X"C9",X"E5",X"C5",X"F5",X"CD",X"A9",X"1D",X"CD",X"B5",X"12",X"CD",X"01",X"28",X"06",X"78",X"3E",
		X"00",X"CD",X"B0",X"04",X"CD",X"15",X"08",X"3C",X"10",X"F7",X"CD",X"B5",X"12",X"F1",X"C1",X"E1",
		X"C9",X"0D",X"21",X"0F",X"28",X"C8",X"3D",X"21",X"33",X"28",X"C8",X"21",X"5F",X"28",X"C9",X"01",
		X"1F",X"00",X"0F",X"1B",X"28",X"27",X"28",X"01",X"0C",X"48",X"40",X"50",X"4C",X"41",X"59",X"45",
		X"52",X"20",X"52",X"45",X"41",X"44",X"59",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"01",X"1F",X"00",X"0F",X"3F",X"28",X"4F",X"28",X"01",X"10",X"48",X"30",X"50",
		X"4C",X"41",X"59",X"45",X"52",X"20",X"4F",X"4E",X"45",X"20",X"52",X"45",X"41",X"44",X"59",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"01",
		X"1F",X"00",X"0F",X"6B",X"28",X"4F",X"28",X"01",X"10",X"48",X"30",X"50",X"4C",X"41",X"59",X"45",
		X"52",X"20",X"54",X"57",X"4F",X"20",X"52",X"45",X"41",X"44",X"59",X"C5",X"F5",X"FD",X"7E",X"46",
		X"3C",X"28",X"0F",X"06",X"FF",X"FD",X"7E",X"32",X"CD",X"DD",X"0A",X"28",X"02",X"06",X"00",X"FD",
		X"70",X"46",X"C1",X"78",X"C1",X"C9",X"D5",X"C5",X"F5",X"CD",X"F8",X"28",X"CD",X"37",X"29",X"CD",
		X"95",X"29",X"CD",X"C8",X"18",X"28",X"42",X"CD",X"BA",X"21",X"3E",X"01",X"CD",X"27",X"17",X"CD",
		X"61",X"23",X"CD",X"C8",X"18",X"28",X"32",X"CD",X"BA",X"21",X"3E",X"01",X"CD",X"27",X"17",X"7A",
		X"FD",X"46",X"41",X"04",X"FD",X"36",X"47",X"00",X"FD",X"36",X"41",X"00",X"28",X"E1",X"3E",X"01",
		X"CD",X"27",X"17",X"CD",X"7D",X"25",X"CD",X"C8",X"18",X"28",X"0E",X"CD",X"87",X"27",X"FD",X"7E",
		X"37",X"CD",X"33",X"04",X"3E",X"64",X"CD",X"FA",X"26",X"CD",X"78",X"29",X"28",X"04",X"F1",X"C1",
		X"D1",X"C9",X"FD",X"36",X"01",X"00",X"18",X"F6",X"E5",X"D5",X"C5",X"F5",X"21",X"19",X"29",X"0D",
		X"28",X"09",X"21",X"23",X"29",X"3D",X"28",X"03",X"21",X"2D",X"29",X"11",X"F8",X"48",X"01",X"01",
		X"0A",X"CD",X"E2",X"0B",X"F1",X"C1",X"D1",X"E1",X"C9",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"4F",X"4E",X"45",X"50",X"4C",X"41",
		X"59",X"45",X"52",X"20",X"54",X"57",X"4F",X"E5",X"D5",X"C5",X"FD",X"36",X"35",X"00",X"FD",X"36",
		X"34",X"00",X"FD",X"36",X"38",X"00",X"FD",X"36",X"41",X"FF",X"FD",X"36",X"47",X"FF",X"FD",X"36",
		X"3F",X"00",X"FD",X"70",X"32",X"FD",X"77",X"37",X"21",X"4D",X"40",X"22",X"5D",X"40",X"21",X"4D",
		X"40",X"11",X"4E",X"40",X"01",X"0A",X"00",X"36",X"00",X"ED",X"B0",X"CD",X"59",X"2E",X"CD",X"33",
		X"04",X"CD",X"61",X"16",X"C1",X"D1",X"E1",X"C9",X"E5",X"C5",X"F5",X"FD",X"E5",X"E1",X"01",X"02",
		X"00",X"09",X"3E",X"00",X"06",X"04",X"BE",X"20",X"07",X"23",X"10",X"FA",X"FD",X"36",X"33",X"02",
		X"C1",X"78",X"C1",X"E1",X"C9",X"E5",X"F5",X"CD",X"AC",X"18",X"CD",X"73",X"2C",X"CD",X"E1",X"27",
		X"3E",X"02",X"32",X"8D",X"40",X"21",X"FD",X"29",X"11",X"03",X"2A",X"01",X"06",X"00",X"CD",X"28",
		X"2A",X"CD",X"4F",X"2A",X"3E",X"00",X"32",X"89",X"40",X"FD",X"36",X"33",X"01",X"FD",X"36",X"36",
		X"00",X"FD",X"36",X"46",X"00",X"CD",X"C8",X"18",X"28",X"29",X"CD",X"88",X"2A",X"CD",X"F0",X"2A",
		X"CD",X"3D",X"2A",X"CD",X"7B",X"28",X"20",X"06",X"21",X"F6",X"29",X"CD",X"EF",X"2B",X"67",X"CD",
		X"2C",X"05",X"7C",X"CD",X"15",X"08",X"3C",X"CD",X"78",X"29",X"FD",X"6E",X"36",X"2C",X"20",X"D5",
		X"CD",X"25",X"2C",X"F1",X"E1",X"C9",X"03",X"F3",X"2C",X"73",X"2C",X"24",X"2E",X"60",X"00",X"26",
		X"00",X"24",X"00",X"09",X"2A",X"0A",X"2A",X"14",X"2A",X"00",X"01",X"0F",X"00",X"09",X"26",X"00",
		X"27",X"00",X"40",X"38",X"01",X"0F",X"00",X"09",X"24",X"00",X"25",X"00",X"40",X"60",X"01",X"0F",
		X"00",X"09",X"36",X"00",X"36",X"00",X"40",X"38",X"E5",X"D5",X"C5",X"D5",X"11",X"5F",X"40",X"C5",
		X"ED",X"B0",X"C1",X"E1",X"11",X"75",X"40",X"ED",X"B0",X"C1",X"D1",X"E1",X"C9",X"E5",X"F5",X"3E",
		X"00",X"FD",X"B6",X"35",X"20",X"06",X"21",X"0A",X"2A",X"22",X"77",X"40",X"F1",X"E1",X"C9",X"E5",
		X"D5",X"C5",X"F5",X"21",X"5F",X"40",X"11",X"40",X"10",X"7E",X"23",X"06",X"02",X"E5",X"23",X"0E",
		X"05",X"07",X"DC",X"7C",X"2A",X"F5",X"3E",X"28",X"82",X"57",X"F1",X"0D",X"20",X"F3",X"D1",X"1A",
		X"11",X"28",X"10",X"E5",X"10",X"E9",X"E1",X"F1",X"C1",X"D1",X"E1",X"C9",X"D5",X"5E",X"23",X"56",
		X"23",X"E3",X"EB",X"CD",X"35",X"0C",X"E1",X"C9",X"E5",X"D5",X"C5",X"F5",X"21",X"75",X"40",X"CD",
		X"C5",X"1C",X"FD",X"7E",X"33",X"87",X"5F",X"16",X"00",X"19",X"7E",X"23",X"66",X"6F",X"F1",X"CD",
		X"37",X"2C",X"F5",X"3E",X"03",X"CD",X"72",X"0B",X"21",X"C5",X"2A",X"11",X"18",X"20",X"01",X"01",
		X"13",X"CD",X"E2",X"0B",X"21",X"D8",X"2A",X"11",X"10",X"10",X"01",X"01",X"18",X"CD",X"E2",X"0B",
		X"F1",X"C1",X"D1",X"E1",X"C9",X"53",X"45",X"4C",X"45",X"43",X"54",X"20",X"43",X"48",X"4F",X"49",
		X"43",X"45",X"20",X"55",X"53",X"49",X"4E",X"47",X"4A",X"4F",X"59",X"53",X"54",X"49",X"43",X"4B",
		X"20",X"41",X"4E",X"44",X"20",X"46",X"49",X"52",X"45",X"20",X"42",X"55",X"54",X"54",X"4F",X"4E",
		X"D5",X"F5",X"3E",X"00",X"FD",X"B6",X"34",X"28",X"05",X"FD",X"35",X"34",X"18",X"1B",X"21",X"5F",
		X"40",X"FD",X"7E",X"32",X"CD",X"94",X"0A",X"3E",X"00",X"B2",X"20",X"10",X"B3",X"20",X"1F",X"18",
		X"08",X"CD",X"4F",X"2A",X"3E",X"14",X"FD",X"77",X"34",X"F1",X"D1",X"C9",X"7A",X"07",X"38",X"07",
		X"3E",X"00",X"CD",X"40",X"2B",X"18",X"EA",X"3E",X"01",X"CD",X"40",X"2B",X"18",X"E3",X"7B",X"07",
		X"38",X"07",X"3E",X"01",X"CD",X"96",X"2B",X"18",X"D8",X"3E",X"00",X"CD",X"96",X"2B",X"18",X"D1",
		X"E5",X"D5",X"C5",X"F5",X"0F",X"FD",X"7E",X"33",X"38",X"26",X"FE",X"05",X"01",X"00",X"05",X"38",
		X"03",X"01",X"05",X"0A",X"3C",X"B8",X"20",X"01",X"79",X"CD",X"D3",X"2B",X"20",X"F6",X"CD",X"E8",
		X"1A",X"CD",X"19",X"1D",X"FD",X"36",X"46",X"00",X"CD",X"AC",X"18",X"FD",X"77",X"33",X"18",X"21",
		X"FE",X"05",X"01",X"FF",X"04",X"38",X"03",X"01",X"04",X"09",X"3D",X"B9",X"20",X"01",X"78",X"CD",
		X"D3",X"2B",X"20",X"F6",X"CD",X"E8",X"1A",X"CD",X"19",X"1D",X"FD",X"36",X"46",X"00",X"FD",X"77",
		X"33",X"F1",X"C1",X"D1",X"E1",X"C9",X"C5",X"F5",X"0F",X"38",X"1D",X"FD",X"7E",X"33",X"3E",X"09",
		X"FE",X"0A",X"30",X"2C",X"CD",X"D3",X"2B",X"20",X"27",X"CD",X"E8",X"1A",X"CD",X"19",X"1D",X"FD",
		X"36",X"46",X"00",X"FD",X"77",X"33",X"18",X"18",X"FD",X"7E",X"33",X"D6",X"05",X"38",X"11",X"CD",
		X"D3",X"2B",X"20",X"0C",X"CD",X"E8",X"1A",X"CD",X"19",X"1D",X"CD",X"AC",X"18",X"FD",X"77",X"33",
		X"F1",X"C1",X"C9",X"E5",X"C5",X"F5",X"FE",X"05",X"38",X"03",X"23",X"D6",X"05",X"3C",X"47",X"7E",
		X"07",X"10",X"FD",X"3E",X"00",X"38",X"02",X"3E",X"01",X"B7",X"C1",X"78",X"C1",X"E1",X"C9",X"E5",
		X"F5",X"3E",X"00",X"FD",X"B6",X"35",X"28",X"05",X"FD",X"35",X"35",X"18",X"25",X"FD",X"7E",X"32",
		X"CD",X"DD",X"0A",X"3E",X"00",X"28",X"18",X"CD",X"E8",X"1A",X"CD",X"AC",X"18",X"3E",X"00",X"CD",
		X"88",X"2A",X"FD",X"7E",X"33",X"CD",X"3B",X"00",X"3E",X"0A",X"FD",X"77",X"35",X"3E",X"FF",X"FD",
		X"77",X"38",X"F1",X"E1",X"C9",X"D5",X"C5",X"F5",X"01",X"50",X"C0",X"11",X"10",X"10",X"3E",X"20",
		X"CD",X"DD",X"09",X"F1",X"C1",X"D1",X"C9",X"E5",X"D5",X"C5",X"F5",X"4F",X"7E",X"A7",X"28",X"2E",
		X"47",X"23",X"7E",X"23",X"A1",X"BE",X"23",X"20",X"08",X"23",X"5E",X"23",X"56",X"23",X"23",X"18",
		X"09",X"BE",X"20",X"14",X"23",X"23",X"23",X"5E",X"23",X"56",X"23",X"7E",X"23",X"E5",X"66",X"6F",
		X"EB",X"CD",X"35",X"0C",X"E1",X"23",X"18",X"04",X"11",X"07",X"00",X"19",X"10",X"D4",X"F1",X"C1",
		X"D1",X"E1",X"C9",X"E5",X"D5",X"F5",X"21",X"1E",X"2A",X"22",X"77",X"40",X"CD",X"93",X"2C",X"CD",
		X"31",X"18",X"3E",X"00",X"FD",X"BE",X"08",X"38",X"04",X"F1",X"D1",X"E1",X"C9",X"F1",X"D1",X"E1",
		X"C3",X"24",X"2E",X"F5",X"FD",X"7E",X"38",X"3C",X"CA",X"A3",X"2C",X"3E",X"00",X"32",X"89",X"40",
		X"C3",X"D6",X"2C",X"FD",X"7E",X"02",X"E6",X"0F",X"C2",X"D6",X"2C",X"3A",X"89",X"40",X"E6",X"01",
		X"CA",X"D6",X"2C",X"FD",X"7E",X"02",X"E6",X"F0",X"C2",X"F4",X"2C",X"3A",X"89",X"40",X"E6",X"02",
		X"CA",X"F4",X"2C",X"FD",X"7E",X"03",X"E6",X"0F",X"C2",X"3A",X"2D",X"3A",X"89",X"40",X"E6",X"04",
		X"CA",X"3A",X"2D",X"C3",X"80",X"2D",X"3A",X"89",X"40",X"F6",X"01",X"32",X"89",X"40",X"21",X"EF",
		X"2C",X"CD",X"E9",X"2D",X"21",X"03",X"17",X"CD",X"BE",X"2D",X"CD",X"59",X"1C",X"F1",X"C9",X"01",
		X"00",X"00",X"00",X"C9",X"3A",X"89",X"40",X"F6",X"02",X"32",X"89",X"40",X"3E",X"0A",X"CD",X"FA",
		X"26",X"21",X"12",X"2D",X"CD",X"E9",X"2D",X"21",X"16",X"2D",X"CD",X"BE",X"2D",X"CD",X"74",X"1C",
		X"F1",X"C9",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"04",
		X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"20",X"00",X"00",X"3A",X"89",X"40",X"F6",X"04",X"32",
		X"89",X"40",X"3E",X"0A",X"CD",X"FA",X"26",X"21",X"58",X"2D",X"CD",X"E9",X"2D",X"21",X"5C",X"2D",
		X"CD",X"BE",X"2D",X"CD",X"8F",X"1C",X"F1",X"C9",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",
		X"00",X"02",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"10",X"00",X"00",
		X"00",X"20",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"02",X"00",
		X"3E",X"0A",X"CD",X"FA",X"26",X"21",X"96",X"2D",X"CD",X"E9",X"2D",X"21",X"9A",X"2D",X"CD",X"BE",
		X"2D",X"CD",X"AA",X"1C",X"F1",X"C9",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"20",
		X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"02",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"20",X"00",X"E5",X"D5",
		X"C5",X"F5",X"E5",X"FD",X"E5",X"E1",X"11",X"06",X"00",X"19",X"EB",X"6B",X"62",X"C1",X"3E",X"09",
		X"F5",X"3E",X"04",X"CD",X"C1",X"03",X"03",X"03",X"03",X"03",X"23",X"23",X"23",X"23",X"5D",X"54",
		X"F1",X"3D",X"20",X"EC",X"F1",X"C1",X"D1",X"E1",X"C9",X"E5",X"D5",X"C5",X"F5",X"E5",X"FD",X"E5",
		X"E1",X"01",X"02",X"00",X"09",X"EB",X"42",X"4B",X"E1",X"3E",X"04",X"CD",X"09",X"2E",X"FD",X"7E",
		X"37",X"CD",X"33",X"04",X"F1",X"C1",X"D1",X"E1",X"C9",X"A7",X"C8",X"E5",X"D5",X"C5",X"F5",X"F5",
		X"97",X"0A",X"9E",X"27",X"12",X"03",X"13",X"23",X"E3",X"25",X"E3",X"20",X"F4",X"E1",X"E1",X"7C",
		X"C1",X"D1",X"E1",X"C9",X"E5",X"D5",X"C5",X"F5",X"21",X"5F",X"40",X"3A",X"8D",X"40",X"87",X"4F",
		X"06",X"00",X"09",X"11",X"35",X"00",X"73",X"23",X"72",X"CD",X"4F",X"2A",X"3E",X"00",X"CD",X"27",
		X"17",X"FD",X"36",X"36",X"FF",X"CD",X"59",X"2E",X"CD",X"77",X"2E",X"CD",X"A0",X"2E",X"CD",X"FE",
		X"1C",X"CD",X"58",X"18",X"F1",X"C1",X"D1",X"E1",X"C9",X"E5",X"C5",X"F5",X"FD",X"7E",X"3F",X"FD",
		X"E5",X"E1",X"01",X"2B",X"00",X"09",X"06",X"05",X"0F",X"38",X"02",X"36",X"00",X"23",X"10",X"F8",
		X"CD",X"58",X"18",X"F1",X"C1",X"E1",X"C9",X"E5",X"C5",X"F5",X"FD",X"7E",X"3F",X"FD",X"E5",X"E1",
		X"01",X"2B",X"00",X"09",X"06",X"05",X"0F",X"38",X"10",X"36",X"0E",X"CD",X"58",X"18",X"CD",X"E5",
		X"1C",X"0E",X"1E",X"CD",X"15",X"08",X"0D",X"20",X"FA",X"23",X"10",X"EA",X"F1",X"C1",X"E1",X"C9",
		X"E5",X"D5",X"C5",X"F5",X"FD",X"7E",X"3F",X"FD",X"E5",X"E1",X"01",X"2B",X"00",X"09",X"5D",X"54",
		X"06",X"05",X"0F",X"F5",X"38",X"15",X"CD",X"2C",X"05",X"4F",X"E6",X"0F",X"28",X"F8",X"FE",X"0E",
		X"30",X"F4",X"79",X"E6",X"3F",X"CD",X"D4",X"2E",X"28",X"EC",X"12",X"13",X"F1",X"10",X"E3",X"F1",
		X"C1",X"D1",X"E1",X"C9",X"E5",X"C5",X"F5",X"21",X"4D",X"40",X"06",X"0E",X"BE",X"23",X"28",X"0D",
		X"10",X"FA",X"2A",X"5D",X"40",X"77",X"23",X"22",X"5D",X"40",X"3E",X"01",X"B7",X"C1",X"78",X"C1",
		X"E1",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"FF",X"FF",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"7F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"7F",X"FF",X"FF",X"3F",X"FF",X"FF",X"FF",X"3F",X"3F",X"3F",X"FF",X"FF",X"FF",X"7F",X"3F",X"3F",
		X"FF",X"3F",X"BF",X"FF",X"BF",X"3F",X"3F",X"3F",X"3F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
