library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity bwidow_pgm_rom3 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of bwidow_pgm_rom3 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"C9",X"10",X"B0",X"03",X"9D",X"05",X"02",X"20",X"31",X"B1",X"20",X"B4",X"C9",X"20",X"DE",X"C3",
		X"4C",X"5C",X"A6",X"16",X"20",X"14",X"60",X"61",X"D0",X"99",X"14",X"EB",X"58",X"D1",X"76",X"00",
		X"80",X"6A",X"6A",X"A9",X"FF",X"85",X"47",X"4A",X"85",X"46",X"A9",X"00",X"A8",X"48",X"F0",X"18",
		X"B9",X"00",X"02",X"29",X"03",X"C9",X"02",X"B0",X"14",X"B9",X"01",X"02",X"29",X"0F",X"C9",X"0B",
		X"D0",X"0B",X"A5",X"9A",X"29",X"03",X"F0",X"05",X"A6",X"40",X"20",X"03",X"CE",X"68",X"18",X"69",
		X"10",X"90",X"D9",X"A5",X"47",X"60",X"A9",X"FF",X"85",X"47",X"4A",X"85",X"46",X"A9",X"00",X"A8",
		X"48",X"F0",X"16",X"B9",X"00",X"02",X"29",X"03",X"C9",X"02",X"B0",X"12",X"B9",X"01",X"02",X"29",
		X"0F",X"C9",X"01",X"F0",X"04",X"C9",X"0B",X"D0",X"05",X"A6",X"40",X"20",X"03",X"CE",X"68",X"18",
		X"69",X"10",X"90",X"DB",X"A5",X"47",X"60",X"A9",X"FF",X"85",X"47",X"A9",X"7F",X"85",X"46",X"A0",
		X"50",X"84",X"1C",X"B9",X"00",X"02",X"29",X"02",X"D0",X"16",X"24",X"EF",X"30",X"0D",X"B9",X"01",
		X"02",X"29",X"0F",X"AA",X"BD",X"13",X"B0",X"29",X"10",X"F0",X"05",X"A6",X"40",X"20",X"03",X"CE",
		X"A5",X"1C",X"18",X"69",X"10",X"A8",X"D0",X"D9",X"A5",X"47",X"30",X"4A",X"A6",X"40",X"9D",X"0E",
		X"02",X"20",X"31",X"B1",X"60",X"A9",X"FF",X"85",X"47",X"4A",X"85",X"46",X"A0",X"00",X"A6",X"40",
		X"20",X"03",X"CE",X"A6",X"40",X"A0",X"50",X"84",X"1C",X"20",X"49",X"AF",X"90",X"05",X"A6",X"40",
		X"20",X"03",X"CE",X"A5",X"1C",X"18",X"69",X"10",X"A8",X"D0",X"EC",X"A6",X"40",X"A5",X"47",X"10",
		X"11",X"A6",X"40",X"BD",X"06",X"02",X"18",X"69",X"10",X"29",X"3F",X"9D",X"0E",X"02",X"20",X"31",
		X"B1",X"60",X"9D",X"0E",X"02",X"60",X"A6",X"40",X"20",X"12",X"B1",X"9D",X"0E",X"02",X"20",X"31",
		X"B1",X"60",X"A9",X"00",X"38",X"FD",X"0A",X"02",X"C9",X"80",X"6A",X"85",X"42",X"A9",X"00",X"38",
		X"FD",X"0C",X"02",X"C9",X"80",X"6A",X"AA",X"A4",X"42",X"20",X"69",X"A2",X"29",X"3F",X"A6",X"40",
		X"60",X"AD",X"44",X"04",X"09",X"01",X"85",X"1B",X"BD",X"0E",X"02",X"38",X"FD",X"06",X"02",X"F0",
		X"16",X"30",X"1F",X"C9",X"21",X"B0",X"11",X"C5",X"1B",X"90",X"02",X"A5",X"1B",X"18",X"7D",X"06",
		X"02",X"29",X"3F",X"9D",X"06",X"02",X"A8",X"60",X"85",X"1C",X"A9",X"40",X"38",X"E5",X"1C",X"4C",
		X"67",X"B1",X"49",X"FF",X"18",X"69",X"01",X"C9",X"21",X"90",X"06",X"38",X"E9",X"20",X"4C",X"47",
		X"B1",X"85",X"1C",X"C5",X"1B",X"90",X"04",X"A5",X"1B",X"85",X"1C",X"BD",X"06",X"02",X"38",X"E5",
		X"1C",X"29",X"3F",X"9D",X"06",X"02",X"A8",X"60",X"E7",X"60",X"08",X"76",X"E4",X"60",X"07",X"75",
		X"E3",X"60",X"4A",X"74",X"E6",X"60",X"11",X"74",X"E2",X"60",X"59",X"73",X"E4",X"60",X"24",X"73",
		X"E5",X"60",X"71",X"72",X"E1",X"60",X"3F",X"72",X"E7",X"60",X"0F",X"72",X"03",X"00",X"74",X"04",
		X"40",X"73",X"05",X"00",X"73",X"07",X"40",X"72",X"09",X"00",X"72",X"0D",X"40",X"71",X"0F",X"20",
		X"71",X"11",X"00",X"71",X"EE",X"00",X"0A",X"00",X"05",X"02",X"05",X"00",X"05",X"FE",X"0A",X"00",
		X"05",X"02",X"05",X"00",X"FF",X"14",X"20",X"02",X"20",X"FE",X"14",X"00",X"FF",X"14",X"10",X"02",
		X"0F",X"00",X"08",X"FC",X"0F",X"00",X"FF",X"1E",X"20",X"02",X"10",X"FC",X"08",X"08",X"FF",X"14",
		X"00",X"24",X"EF",X"30",X"03",X"4C",X"26",X"B4",X"A5",X"5E",X"D0",X"2B",X"A5",X"79",X"C9",X"02",
		X"B0",X"15",X"A5",X"F7",X"29",X"01",X"D0",X"0E",X"A2",X"10",X"A9",X"03",X"9D",X"00",X"02",X"8A",
		X"18",X"69",X"10",X"AA",X"D0",X"F4",X"60",X"A9",X"00",X"85",X"73",X"A5",X"F7",X"0A",X"AA",X"BD",
		X"29",X"B2",X"48",X"BD",X"28",X"B2",X"48",X"60",X"37",X"B2",X"BA",X"B2",X"62",X"B2",X"BA",X"B2",
		X"7D",X"B2",X"BA",X"B2",X"9D",X"B2",X"BA",X"B2",X"A9",X"E6",X"85",X"4C",X"A9",X"B2",X"85",X"4D",
		X"A2",X"40",X"A9",X"00",X"8D",X"09",X"02",X"8D",X"0B",X"02",X"8D",X"0A",X"02",X"A9",X"28",X"8D",
		X"0C",X"02",X"4C",X"55",X"B2",X"A9",X"50",X"85",X"49",X"A9",X"02",X"85",X"4A",X"20",X"5C",X"A0",
		X"4C",X"CE",X"B2",X"A9",X"26",X"85",X"4C",X"A9",X"B3",X"85",X"4D",X"A2",X"60",X"A9",X"00",X"8D",
		X"09",X"02",X"8D",X"0B",X"02",X"8D",X"0A",X"02",X"8D",X"0C",X"02",X"4C",X"55",X"B2",X"A9",X"86",
		X"85",X"4C",X"A9",X"B3",X"85",X"4D",X"A2",X"60",X"A9",X"00",X"8D",X"09",X"02",X"8D",X"0B",X"02",
		X"8D",X"0A",X"02",X"8D",X"03",X"03",X"A9",X"40",X"8D",X"0C",X"02",X"4C",X"55",X"B2",X"A9",X"E6",
		X"85",X"4C",X"A9",X"B3",X"85",X"4D",X"A2",X"40",X"A9",X"00",X"8D",X"09",X"02",X"8D",X"0B",X"02",
		X"8D",X"0C",X"02",X"A9",X"18",X"8D",X"0A",X"02",X"4C",X"55",X"B2",X"A2",X"50",X"BD",X"00",X"02",
		X"29",X"03",X"C9",X"03",X"F0",X"01",X"60",X"8A",X"18",X"69",X"10",X"AA",X"D0",X"EF",X"A9",X"00",
		X"85",X"79",X"E6",X"F7",X"A5",X"F7",X"C9",X"08",X"B0",X"01",X"60",X"A9",X"02",X"8D",X"23",X"04",
		X"A9",X"00",X"8D",X"22",X"04",X"60",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"18",X"00",X"03",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"10",X"00",X"03",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"D0",X"08",X"00",X"03",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"06",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",
		X"28",X"00",X"50",X"01",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",
		X"64",X"00",X"14",X"01",X"00",X"02",X"00",X"02",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",
		X"50",X"00",X"C4",X"01",X"00",X"03",X"00",X"02",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",
		X"D8",X"00",X"B0",X"01",X"00",X"03",X"00",X"07",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",
		X"9C",X"00",X"EC",X"01",X"00",X"04",X"00",X"07",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",
		X"B0",X"00",X"3C",X"01",X"00",X"04",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"18",X"00",X"03",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"00",X"E0",X"14",X"00",X"03",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"00",X"C0",X"10",X"00",X"03",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"28",X"00",X"E0",X"0C",X"00",X"03",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"D8",X"08",X"00",X"03",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"B8",X"00",X"C8",X"04",X"00",X"03",X"00",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A0",X"00",X"18",X"04",X"00",X"03",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"98",X"00",X"30",X"04",X"00",X"03",X"00",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A8",X"00",X"E0",X"04",X"00",X"03",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"98",X"00",X"D8",X"04",X"00",X"03",X"AD",X"01",X"03",X"05",X"73",X"05",X"6C",X"F0",X"01",X"60",
		X"A5",X"5E",X"D0",X"FB",X"A2",X"0F",X"A9",X"00",X"18",X"7D",X"48",X"04",X"CA",X"10",X"F9",X"8D",
		X"36",X"04",X"AD",X"28",X"04",X"D0",X"08",X"AD",X"36",X"04",X"F0",X"36",X"4C",X"B2",X"B4",X"AD",
		X"36",X"04",X"D0",X"09",X"AD",X"3A",X"04",X"D0",X"03",X"4C",X"D2",X"B4",X"60",X"CE",X"21",X"01",
		X"30",X"01",X"60",X"AE",X"58",X"04",X"E0",X"08",X"90",X"02",X"A2",X"07",X"BD",X"D4",X"B7",X"8D",
		X"21",X"01",X"A9",X"0B",X"38",X"ED",X"51",X"04",X"0A",X"0A",X"0A",X"0A",X"69",X"50",X"AA",X"4C",
		X"EB",X"B6",X"AD",X"3A",X"04",X"0D",X"04",X"03",X"D0",X"03",X"4C",X"D2",X"B4",X"A5",X"79",X"29",
		X"0F",X"F0",X"01",X"60",X"A5",X"6F",X"29",X"1F",X"D0",X"F9",X"EE",X"44",X"04",X"AD",X"44",X"04",
		X"C9",X"08",X"90",X"03",X"CE",X"44",X"04",X"AD",X"3D",X"04",X"C9",X"0B",X"B0",X"03",X"EE",X"3D",
		X"04",X"60",X"AD",X"3A",X"04",X"18",X"6D",X"04",X"03",X"CD",X"3D",X"04",X"90",X"06",X"20",X"8D",
		X"B4",X"4C",X"9F",X"B6",X"AD",X"3A",X"04",X"F0",X"03",X"4C",X"94",X"B6",X"4C",X"9F",X"B6",X"4C",
		X"8E",X"B5",X"20",X"DC",X"B7",X"A9",X"A0",X"8D",X"00",X"25",X"A9",X"00",X"85",X"4B",X"A9",X"0D",
		X"85",X"5E",X"A9",X"00",X"8D",X"01",X"03",X"85",X"4B",X"8D",X"03",X"03",X"8D",X"D3",X"03",X"85",
		X"79",X"EE",X"5D",X"04",X"24",X"EF",X"30",X"D7",X"AD",X"5A",X"04",X"D0",X"D2",X"AD",X"5D",X"04",
		X"F0",X"CD",X"4A",X"B0",X"CA",X"4A",X"B0",X"C7",X"38",X"E9",X"01",X"85",X"19",X"0A",X"65",X"19",
		X"AA",X"A9",X"00",X"85",X"A5",X"A9",X"0E",X"85",X"5E",X"38",X"AD",X"43",X"04",X"FD",X"D7",X"03",
		X"AD",X"42",X"04",X"FD",X"D6",X"03",X"AD",X"41",X"04",X"FD",X"D5",X"03",X"90",X"52",X"AD",X"41",
		X"04",X"9D",X"D5",X"03",X"85",X"1B",X"AD",X"42",X"04",X"9D",X"D6",X"03",X"85",X"1C",X"AD",X"43",
		X"04",X"9D",X"D7",X"03",X"85",X"1D",X"A5",X"1C",X"F8",X"18",X"69",X"50",X"85",X"1C",X"A5",X"1B",
		X"69",X"01",X"85",X"1B",X"D8",X"E8",X"E8",X"E8",X"E0",X"4B",X"B0",X"24",X"BD",X"D7",X"03",X"38",
		X"E5",X"1D",X"BD",X"D6",X"03",X"E5",X"1C",X"BD",X"D5",X"03",X"E5",X"1B",X"B0",X"D8",X"A5",X"1D",
		X"9D",X"D7",X"03",X"A5",X"1C",X"9D",X"D6",X"03",X"A5",X"1B",X"9D",X"D5",X"03",X"4C",X"46",X"B5",
		X"A5",X"9A",X"8D",X"5B",X"04",X"AD",X"5D",X"04",X"8D",X"59",X"04",X"20",X"56",X"BD",X"AD",X"5D",
		X"04",X"C9",X"21",X"90",X"11",X"29",X"07",X"D0",X"0D",X"EE",X"5C",X"04",X"AD",X"5C",X"04",X"C9",
		X"08",X"90",X"03",X"CE",X"5C",X"04",X"AD",X"5D",X"04",X"29",X"03",X"49",X"03",X"D0",X"35",X"8D",
		X"34",X"01",X"A9",X"01",X"8D",X"28",X"04",X"06",X"9A",X"E6",X"9A",X"A2",X"10",X"A9",X"03",X"9D",
		X"00",X"02",X"8A",X"18",X"69",X"10",X"AA",X"D0",X"F4",X"A9",X"01",X"8D",X"21",X"01",X"AD",X"58",
		X"04",X"18",X"69",X"01",X"C9",X"0A",X"B0",X"03",X"8D",X"58",X"04",X"8D",X"44",X"04",X"A9",X"0B",
		X"8D",X"51",X"04",X"60",X"AD",X"5D",X"04",X"85",X"19",X"38",X"E9",X"3C",X"30",X"07",X"29",X"07",
		X"18",X"69",X"34",X"85",X"19",X"A5",X"19",X"0A",X"65",X"19",X"AA",X"BD",X"AF",X"B8",X"29",X"0F",
		X"0A",X"09",X"01",X"8D",X"3F",X"04",X"BD",X"AF",X"B8",X"4A",X"4A",X"4A",X"4A",X"8D",X"44",X"04",
		X"BD",X"B0",X"B8",X"8D",X"3D",X"04",X"BD",X"B1",X"B8",X"8D",X"21",X"01",X"8D",X"3C",X"04",X"A0",
		X"00",X"8C",X"28",X"04",X"A2",X"00",X"8E",X"36",X"04",X"A4",X"19",X"F0",X"13",X"BD",X"63",X"B9",
		X"F0",X"0A",X"29",X"F0",X"C9",X"E0",X"B0",X"04",X"E8",X"4C",X"2D",X"B6",X"E8",X"88",X"D0",X"ED",
		X"BD",X"63",X"B9",X"4A",X"4A",X"4A",X"4A",X"A8",X"BD",X"63",X"B9",X"29",X"0F",X"C0",X"0D",X"B0",
		X"0C",X"85",X"19",X"A5",X"F6",X"F0",X"1D",X"C9",X"02",X"F0",X"23",X"A5",X"19",X"99",X"48",X"04",
		X"18",X"6D",X"36",X"04",X"8D",X"36",X"04",X"BD",X"63",X"B9",X"29",X"F0",X"C9",X"E0",X"B0",X"14",
		X"E8",X"4C",X"40",X"B6",X"A5",X"19",X"0A",X"65",X"19",X"4A",X"4A",X"4C",X"5D",X"B6",X"A5",X"19",
		X"0A",X"4C",X"76",X"B6",X"AD",X"5A",X"04",X"F0",X"0A",X"CE",X"5A",X"04",X"D0",X"05",X"A9",X"01",
		X"8D",X"4D",X"04",X"60",X"CE",X"21",X"01",X"D0",X"24",X"AD",X"3C",X"04",X"8D",X"21",X"01",X"A2",
		X"50",X"BD",X"00",X"02",X"29",X"03",X"C9",X"03",X"F0",X"3C",X"18",X"8A",X"69",X"10",X"AA",X"C9",
		X"00",X"D0",X"EE",X"AD",X"04",X"03",X"F0",X"06",X"A5",X"79",X"8D",X"3E",X"04",X"60",X"A5",X"79",
		X"38",X"ED",X"3E",X"04",X"C9",X"0F",X"90",X"F5",X"AD",X"0A",X"60",X"29",X"F0",X"C9",X"50",X"90",
		X"F7",X"A8",X"B9",X"01",X"02",X"29",X"0F",X"C9",X"05",X"F0",X"ED",X"A9",X"03",X"99",X"00",X"02",
		X"A5",X"79",X"8D",X"3E",X"04",X"60",X"AD",X"28",X"04",X"F0",X"1C",X"AD",X"51",X"04",X"C9",X"0B",
		X"F0",X"06",X"AD",X"36",X"01",X"4C",X"2B",X"B7",X"AD",X"0A",X"60",X"29",X"0F",X"C9",X"0C",X"B0",
		X"F7",X"8D",X"36",X"01",X"4C",X"2B",X"B7",X"A9",X"00",X"85",X"1B",X"AD",X"D1",X"03",X"C9",X"0B",
		X"F0",X"04",X"85",X"1B",X"E6",X"1B",X"AD",X"0A",X"60",X"29",X"0F",X"C9",X"0C",X"90",X"03",X"38",
		X"E9",X"0C",X"CD",X"D1",X"03",X"F0",X"EF",X"C5",X"1B",X"F0",X"EB",X"A8",X"B9",X"C8",X"B7",X"9D",
		X"06",X"02",X"A9",X"01",X"9D",X"0D",X"02",X"98",X"0A",X"0A",X"A8",X"B9",X"E7",X"B7",X"9D",X"09",
		X"02",X"B9",X"E8",X"B7",X"9D",X"0A",X"02",X"B9",X"E9",X"B7",X"9D",X"0B",X"02",X"B9",X"EA",X"B7",
		X"9D",X"0C",X"02",X"8A",X"A8",X"AD",X"28",X"04",X"F0",X"17",X"AD",X"44",X"04",X"99",X"05",X"02",
		X"A9",X"C6",X"9D",X"02",X"02",X"A9",X"B1",X"9D",X"03",X"02",X"A2",X"09",X"86",X"19",X"4C",X"AC",
		X"B7",X"AD",X"44",X"04",X"99",X"05",X"02",X"AD",X"0A",X"60",X"29",X"0F",X"AA",X"85",X"19",X"C9",
		X"0E",X"90",X"24",X"AD",X"3A",X"04",X"D0",X"0D",X"AD",X"36",X"04",X"CD",X"56",X"04",X"F0",X"2F",
		X"CD",X"57",X"04",X"F0",X"2A",X"A5",X"79",X"C9",X"05",X"90",X"23",X"A9",X"00",X"99",X"02",X"02",
		X"AD",X"44",X"04",X"4A",X"99",X"05",X"02",X"BD",X"48",X"04",X"F0",X"CB",X"DE",X"48",X"04",X"B9",
		X"01",X"02",X"29",X"F0",X"05",X"19",X"99",X"01",X"02",X"A9",X"00",X"99",X"00",X"02",X"60",X"A9",
		X"00",X"8D",X"56",X"04",X"8D",X"57",X"04",X"60",X"25",X"29",X"2E",X"32",X"37",X"3B",X"05",X"09",
		X"0E",X"12",X"17",X"1B",X"10",X"09",X"08",X"07",X"06",X"05",X"04",X"03",X"A2",X"0B",X"A9",X"00",
		X"9D",X"29",X"04",X"CA",X"10",X"FA",X"60",X"00",X"28",X"00",X"50",X"00",X"50",X"00",X"3C",X"00",
		X"64",X"00",X"14",X"00",X"64",X"00",X"EC",X"00",X"50",X"00",X"C4",X"00",X"28",X"00",X"B0",X"00",
		X"D8",X"00",X"B0",X"00",X"B0",X"00",X"C4",X"00",X"9C",X"00",X"EC",X"00",X"9C",X"00",X"14",X"00",
		X"B0",X"00",X"3C",X"00",X"D8",X"00",X"50",X"5E",X"5E",X"58",X"5E",X"5E",X"5E",X"5E",X"5E",X"58",
		X"5E",X"5E",X"5E",X"6A",X"64",X"5E",X"58",X"52",X"4C",X"52",X"58",X"5E",X"64",X"6A",X"6A",X"5E",
		X"5E",X"98",X"5E",X"5E",X"98",X"5E",X"5E",X"98",X"5E",X"5E",X"98",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5E",X"9E",X"5E",X"9E",X"5E",X"9E",X"5E",X"9E",X"5E",
		X"9E",X"5E",X"9E",X"5E",X"98",X"5E",X"98",X"5E",X"98",X"5E",X"98",X"5E",X"98",X"5E",X"98",X"98",
		X"9E",X"A4",X"AA",X"AA",X"AA",X"AA",X"AA",X"92",X"92",X"92",X"92",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"98",X"98",X"98",X"9E",X"9E",X"9E",X"9E",X"9E",X"98",
		X"98",X"98",X"98",X"92",X"92",X"92",X"9E",X"9E",X"9E",X"9E",X"9E",X"92",X"92",X"92",X"92",X"9E",
		X"9E",X"52",X"9E",X"9E",X"9E",X"9E",X"9E",X"52",X"9E",X"9E",X"9E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"BB",X"AA",X"30",X"5F",X"EE",X"3D",X"A8",X"0F",
		X"04",X"19",X"1F",X"05",X"19",X"1F",X"06",X"19",X"00",X"00",X"00",X"1F",X"07",X"19",X"2F",X"08",
		X"19",X"2F",X"09",X"19",X"00",X"00",X"00",X"3F",X"0A",X"18",X"3F",X"0A",X"17",X"3F",X"0A",X"16",
		X"00",X"00",X"00",X"37",X"0A",X"15",X"37",X"0A",X"14",X"47",X"0A",X"14",X"00",X"00",X"00",X"47",
		X"0A",X"14",X"47",X"0A",X"14",X"47",X"0A",X"14",X"00",X"00",X"00",X"47",X"0A",X"14",X"47",X"0A",
		X"14",X"47",X"0A",X"14",X"00",X"00",X"00",X"47",X"0A",X"14",X"47",X"0A",X"14",X"47",X"0A",X"14",
		X"00",X"00",X"00",X"57",X"0A",X"14",X"57",X"0A",X"14",X"57",X"0A",X"14",X"00",X"00",X"00",X"57",
		X"0A",X"14",X"57",X"0A",X"14",X"57",X"0A",X"14",X"00",X"00",X"00",X"57",X"0A",X"0F",X"57",X"0A",
		X"0F",X"57",X"0A",X"0F",X"00",X"00",X"00",X"57",X"0A",X"0F",X"57",X"0A",X"0F",X"57",X"0A",X"0F",
		X"00",X"00",X"00",X"57",X"0B",X"0F",X"57",X"0B",X"0F",X"57",X"0B",X"05",X"00",X"00",X"00",X"57",
		X"0A",X"0F",X"57",X"0A",X"0F",X"57",X"0A",X"0F",X"00",X"00",X"00",X"57",X"0B",X"07",X"57",X"0B",
		X"07",X"67",X"0B",X"07",X"00",X"00",X"00",X"57",X"0B",X"07",X"67",X"0B",X"07",X"77",X"0B",X"07",
		X"00",X"00",X"00",X"25",X"75",X"05",X"E1",X"25",X"75",X"05",X"E1",X"25",X"75",X"05",X"E1",X"00",
		X"25",X"75",X"05",X"E1",X"25",X"75",X"05",X"E1",X"25",X"75",X"05",X"E1",X"00",X"25",X"75",X"05",
		X"D1",X"E1",X"25",X"75",X"05",X"D2",X"E1",X"25",X"75",X"05",X"D4",X"E1",X"00",X"DB",X"E1",X"25",
		X"75",X"05",X"D1",X"E1",X"25",X"75",X"05",X"D2",X"E1",X"00",X"0A",X"F1",X"0A",X"F2",X"0A",X"F3",
		X"00",X"25",X"75",X"05",X"D1",X"F1",X"25",X"75",X"05",X"D2",X"F1",X"25",X"75",X"05",X"D4",X"F1",
		X"00",X"25",X"75",X"05",X"D1",X"F1",X"25",X"75",X"05",X"D2",X"F1",X"25",X"75",X"05",X"D4",X"F1",
		X"00",X"25",X"75",X"05",X"D2",X"F1",X"25",X"75",X"05",X"D4",X"F1",X"25",X"75",X"05",X"D8",X"F1",
		X"00",X"25",X"75",X"05",X"D2",X"F1",X"25",X"75",X"05",X"D4",X"F1",X"25",X"75",X"05",X"D8",X"F1",
		X"00",X"25",X"75",X"05",X"D2",X"F1",X"25",X"75",X"05",X"D2",X"F2",X"25",X"75",X"05",X"D4",X"F4",
		X"00",X"25",X"75",X"05",X"D2",X"F1",X"25",X"75",X"05",X"D4",X"F2",X"25",X"75",X"05",X"D8",X"F4",
		X"00",X"25",X"75",X"05",X"D2",X"F1",X"25",X"75",X"05",X"D4",X"F2",X"25",X"75",X"05",X"D8",X"F4",
		X"00",X"25",X"75",X"05",X"D2",X"F2",X"25",X"75",X"05",X"D4",X"F2",X"25",X"75",X"05",X"D4",X"F2",
		X"00",X"02",X"7A",X"2A",X"D4",X"F3",X"04",X"7A",X"2A",X"D4",X"F3",X"06",X"7A",X"2A",X"D4",X"F3",
		X"00",X"06",X"7A",X"2A",X"D4",X"F3",X"08",X"7A",X"2A",X"D4",X"F3",X"0A",X"7A",X"2A",X"D4",X"F3",
		X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"6B",X"6E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"ED",X"F4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"29",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"5A",X"00",X"00",X"00",X"00",
		X"00",X"00",X"19",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"71",X"86",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9F",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"4C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"9C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B5",X"C6",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"8B",X"92",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B5",X"C6",X"D9",X"DC",
		X"00",X"00",X"E1",X"E6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"01",X"0F",X"00",X"00",X"2F",X"02",X"FF",X"0F",X"00",X"00",X"00",X"04",
		X"0E",X"03",X"79",X"04",X"0E",X"03",X"00",X"04",X"0E",X"03",X"51",X"04",X"0E",X"07",X"00",X"00",
		X"8F",X"04",X"00",X"03",X"AF",X"04",X"FF",X"03",X"8B",X"04",X"FF",X"03",X"A6",X"04",X"FF",X"07",
		X"00",X"00",X"06",X"30",X"00",X"03",X"00",X"00",X"AF",X"18",X"00",X"01",X"A0",X"18",X"00",X"01",
		X"AF",X"18",X"00",X"01",X"A0",X"18",X"00",X"01",X"AF",X"18",X"00",X"01",X"A0",X"18",X"00",X"01",
		X"00",X"00",X"00",X"08",X"00",X"02",X"10",X"08",X"10",X"03",X"20",X"08",X"10",X"03",X"30",X"08",
		X"10",X"03",X"40",X"08",X"10",X"03",X"50",X"08",X"10",X"03",X"60",X"08",X"10",X"03",X"00",X"00",
		X"2F",X"08",X"00",X"02",X"AF",X"08",X"00",X"04",X"AD",X"08",X"FF",X"0E",X"00",X"00",X"60",X"10",
		X"00",X"01",X"50",X"10",X"F8",X"01",X"48",X"10",X"18",X"01",X"60",X"18",X"F0",X"01",X"60",X"10",
		X"F8",X"01",X"60",X"10",X"08",X"10",X"00",X"00",X"8C",X"20",X"02",X"01",X"8E",X"10",X"00",X"04",
		X"8E",X"38",X"FF",X"04",X"00",X"18",X"00",X"01",X"00",X"00",X"00",X"04",X"10",X"0A",X"00",X"04",
		X"10",X"0A",X"00",X"00",X"05",X"04",X"05",X"02",X"CF",X"04",X"00",X"02",X"0F",X"04",X"00",X"02",
		X"00",X"04",X"00",X"04",X"C5",X"04",X"05",X"02",X"0F",X"04",X"00",X"02",X"CF",X"04",X"00",X"02",
		X"00",X"04",X"00",X"04",X"00",X"00",X"0F",X"04",X"00",X"01",X"00",X"00",X"A8",X"04",X"40",X"01",
		X"00",X"00",X"F0",X"09",X"F0",X"02",X"D0",X"09",X"10",X"02",X"F0",X"09",X"F0",X"02",X"D0",X"09",
		X"10",X"02",X"F0",X"09",X"F0",X"02",X"D0",X"09",X"10",X"02",X"F0",X"09",X"F0",X"02",X"D0",X"09",
		X"10",X"02",X"F0",X"09",X"F0",X"02",X"D0",X"09",X"10",X"02",X"00",X"00",X"AF",X"09",X"FF",X"0A",
		X"A7",X"09",X"01",X"0A",X"00",X"00",X"08",X"04",X"20",X"0A",X"08",X"04",X"01",X"09",X"10",X"0C",
		X"04",X"0C",X"00",X"00",X"0F",X"04",X"00",X"0A",X"6F",X"04",X"00",X"09",X"6F",X"10",X"FF",X"09",
		X"00",X"00",X"B0",X"02",X"00",X"11",X"00",X"00",X"C0",X"02",X"02",X"11",X"00",X"00",X"60",X"01",
		X"00",X"01",X"60",X"01",X"FF",X"40",X"48",X"01",X"FF",X"30",X"30",X"01",X"FF",X"20",X"24",X"01",
		X"FF",X"18",X"1E",X"01",X"FF",X"14",X"1B",X"01",X"FF",X"12",X"18",X"01",X"FF",X"10",X"00",X"00",
		X"A8",X"DE",X"00",X"01",X"A0",X"01",X"00",X"01",X"00",X"00",X"00",X"04",X"00",X"06",X"1B",X"04",
		X"0E",X"03",X"00",X"04",X"00",X"01",X"51",X"04",X"0E",X"03",X"00",X"04",X"00",X"01",X"87",X"04",
		X"0E",X"03",X"00",X"04",X"00",X"01",X"BD",X"04",X"0E",X"02",X"00",X"00",X"4F",X"04",X"00",X"03",
		X"8F",X"04",X"00",X"03",X"AE",X"04",X"FF",X"03",X"4B",X"04",X"00",X"01",X"AA",X"04",X"FF",X"03",
		X"47",X"04",X"00",X"01",X"A6",X"04",X"FF",X"03",X"43",X"04",X"00",X"01",X"A2",X"04",X"FE",X"02",
		X"00",X"00",X"0A",X"FF",X"00",X"10",X"00",X"00",X"40",X"20",X"01",X"0A",X"4A",X"10",X"01",X"06",
		X"00",X"00",X"20",X"01",X"00",X"03",X"70",X"01",X"10",X"06",X"00",X"00",X"AF",X"01",X"FE",X"02",
		X"A0",X"01",X"00",X"01",X"A2",X"02",X"FF",X"03",X"00",X"00",X"36",X"10",X"00",X"03",X"43",X"10",
		X"0E",X"0A",X"D0",X"10",X"00",X"07",X"00",X"00",X"A3",X"10",X"04",X"04",X"AF",X"10",X"FF",X"10",
		X"00",X"00",X"A9",X"0F",X"D0",X"36",X"A9",X"9F",X"D0",X"32",X"A9",X"3F",X"D0",X"2E",X"A9",X"4F",
		X"D0",X"2A",X"A9",X"1F",X"D0",X"26",X"A9",X"5F",X"D0",X"22",X"A9",X"6F",X"D0",X"1E",X"A9",X"7F",
		X"D0",X"1A",X"A9",X"AF",X"D0",X"16",X"A9",X"BF",X"D0",X"12",X"A9",X"CF",X"D0",X"0E",X"A9",X"2F",
		X"D0",X"0A",X"A9",X"DF",X"D0",X"06",X"A9",X"8F",X"D0",X"02",X"A9",X"EF",X"24",X"EF",X"30",X"22",
		X"86",X"ED",X"84",X"EE",X"A8",X"A2",X"0F",X"B9",X"42",X"BA",X"F0",X"0E",X"86",X"F3",X"95",X"AD",
		X"A9",X"01",X"95",X"CD",X"95",X"DD",X"A9",X"FF",X"85",X"F3",X"88",X"CA",X"10",X"E9",X"A6",X"ED",
		X"A4",X"EE",X"60",X"A2",X"0F",X"B5",X"AD",X"F0",X"7E",X"E4",X"F3",X"F0",X"7A",X"D6",X"CD",X"D0",
		X"76",X"D6",X"DD",X"D0",X"38",X"F6",X"AD",X"F6",X"AD",X"B5",X"AD",X"0A",X"A8",X"B0",X"10",X"B9",
		X"2C",X"BB",X"95",X"BD",X"B9",X"2F",X"BB",X"95",X"DD",X"B9",X"2D",X"BB",X"4C",X"BC",X"BD",X"B9",
		X"2C",X"BC",X"95",X"BD",X"B9",X"2F",X"BC",X"95",X"DD",X"B9",X"2D",X"BC",X"95",X"CD",X"D0",X"0A",
		X"95",X"AD",X"B5",X"BD",X"F0",X"04",X"95",X"AD",X"D0",X"CB",X"4C",X"F8",X"BD",X"0A",X"A8",X"B0",
		X"0B",X"B9",X"2D",X"BB",X"95",X"CD",X"B9",X"2E",X"BB",X"4C",X"E4",X"BD",X"B9",X"2D",X"BC",X"95",
		X"CD",X"B9",X"2E",X"BC",X"B4",X"BD",X"18",X"75",X"BD",X"95",X"BD",X"8A",X"4A",X"90",X"09",X"98",
		X"55",X"BD",X"29",X"F0",X"55",X"BD",X"95",X"BD",X"B5",X"BD",X"E0",X"08",X"90",X"06",X"9D",X"F8",
		X"67",X"4C",X"07",X"BE",X"9D",X"00",X"60",X"CA",X"30",X"03",X"4C",X"85",X"BD",X"60",X"A9",X"00",
		X"8D",X"0F",X"60",X"8D",X"0F",X"68",X"A9",X"07",X"8D",X"0F",X"60",X"8D",X"0F",X"68",X"A2",X"07",
		X"A9",X"00",X"9D",X"00",X"60",X"9D",X"00",X"68",X"95",X"AD",X"95",X"BD",X"CA",X"10",X"F3",X"A9",
		X"00",X"8D",X"08",X"60",X"A2",X"00",X"8E",X"08",X"68",X"60",X"02",X"04",X"04",X"FE",X"C4",X"04",
		X"03",X"02",X"FC",X"00",X"05",X"01",X"00",X"FC",X"F8",X"05",X"FF",X"FE",X"FC",X"F8",X"04",X"FD",
		X"FC",X"FE",X"F0",X"02",X"FC",X"FC",X"00",X"EC",X"FE",X"FC",X"FC",X"02",X"E4",X"FC",X"FD",X"FE",
		X"04",X"E0",X"FB",X"FF",X"00",X"04",X"D8",X"FB",X"01",X"02",X"04",X"D8",X"FC",X"03",X"04",X"02",
		X"D0",X"FE",X"04",X"04",X"00",X"CC",X"A2",X"00",X"A9",X"01",X"85",X"6D",X"20",X"C9",X"D8",X"8A",
		X"48",X"BD",X"3A",X"BE",X"85",X"15",X"E8",X"BD",X"3A",X"BE",X"85",X"16",X"A5",X"4E",X"85",X"02",
		X"A5",X"15",X"85",X"03",X"20",X"67",X"A0",X"85",X"09",X"A5",X"01",X"85",X"08",X"A5",X"16",X"85",
		X"03",X"20",X"67",X"A0",X"85",X"0B",X"A5",X"01",X"85",X"0A",X"A9",X"00",X"85",X"0C",X"20",X"E2",
		X"D8",X"A9",X"A0",X"85",X"0C",X"A9",X"58",X"85",X"02",X"A5",X"15",X"85",X"03",X"20",X"67",X"A0",
		X"85",X"09",X"A5",X"01",X"85",X"08",X"A5",X"16",X"85",X"03",X"20",X"67",X"A0",X"85",X"0B",X"A5",
		X"01",X"85",X"0A",X"20",X"E2",X"D8",X"68",X"18",X"69",X"05",X"AA",X"C9",X"3C",X"90",X"9D",X"20",
		X"C9",X"D8",X"A5",X"11",X"85",X"74",X"A5",X"12",X"85",X"75",X"A5",X"4E",X"8D",X"80",X"89",X"85",
		X"05",X"A9",X"00",X"85",X"0C",X"85",X"07",X"AA",X"BD",X"3A",X"BE",X"85",X"03",X"A5",X"05",X"85",
		X"02",X"20",X"67",X"A0",X"85",X"09",X"A5",X"01",X"85",X"08",X"E8",X"BD",X"3A",X"BE",X"85",X"03",
		X"20",X"67",X"A0",X"85",X"0B",X"A5",X"01",X"85",X"0A",X"20",X"E2",X"D8",X"A9",X"A1",X"A2",X"00",
		X"20",X"5B",X"D8",X"A9",X"A0",X"85",X"0C",X"A5",X"07",X"18",X"69",X"05",X"C9",X"3C",X"90",X"C5",
		X"AD",X"3A",X"BE",X"85",X"03",X"20",X"67",X"A0",X"85",X"09",X"A5",X"01",X"85",X"08",X"AD",X"3C",
		X"BE",X"85",X"03",X"20",X"67",X"A0",X"85",X"0B",X"A5",X"01",X"85",X"0A",X"20",X"E2",X"D8",X"A9",
		X"00",X"85",X"0C",X"20",X"C9",X"D8",X"E6",X"6D",X"A5",X"05",X"18",X"65",X"4E",X"C9",X"58",X"90",
		X"8B",X"60",X"29",X"36",X"00",X"09",X"16",X"20",X"29",X"36",X"00",X"09",X"16",X"20",X"80",X"0C",
		X"00",X"0A",X"80",X"1B",X"00",X"19",X"00",X"14",X"00",X"37",X"80",X"25",X"00",X"1E",X"80",X"52",
		X"00",X"32",X"00",X"28",X"00",X"6E",X"80",X"3E",X"00",X"32",X"80",X"89",X"00",X"4B",X"00",X"3C",
		X"00",X"A5",X"80",X"57",X"00",X"46",X"80",X"C0",X"00",X"64",X"00",X"50",X"00",X"DC",X"00",X"00",
		X"5A",X"00",X"00",X"00",X"B4",X"00",X"00",X"00",X"0E",X"01",X"00",X"00",X"68",X"01",X"00",X"00",
		X"C2",X"01",X"00",X"00",X"1C",X"02",X"00",X"00",X"76",X"02",X"00",X"00",X"D0",X"02",X"00",X"00",
		X"2A",X"03",X"00",X"00",X"84",X"03",X"00",X"00",X"DE",X"03",X"00",X"00",X"38",X"04",X"00",X"00",
		X"92",X"04",X"00",X"00",X"EC",X"04",X"00",X"00",X"46",X"05",X"00",X"00",X"A0",X"05",X"06",X"00",
		X"5A",X"00",X"0C",X"00",X"B4",X"00",X"12",X"00",X"0E",X"01",X"18",X"00",X"68",X"01",X"1E",X"00",
		X"C2",X"01",X"24",X"00",X"1C",X"02",X"2A",X"00",X"76",X"02",X"30",X"00",X"D0",X"02",X"36",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
