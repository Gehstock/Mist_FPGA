library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity mpe_43f is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of mpe_43f is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"11",X"7F",X"FF",X"9C",X"08",X"00",
		X"00",X"E0",X"F8",X"FC",X"FC",X"C8",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"0F",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"F0",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"0F",X"FF",X"F1",X"FD",X"FB",X"F7",X"F1",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"30",X"78",X"FC",X"FC",X"FC",X"78",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"FF",X"DF",X"EF",X"07",X"EF",X"DF",X"00",X"00",X"FF",X"1F",X"7F",X"3F",X"7F",X"1F",
		X"00",X"00",X"FF",X"1F",X"BF",X"BF",X"BF",X"7F",X"00",X"00",X"FF",X"1F",X"5F",X"5F",X"5F",X"1F",
		X"00",X"00",X"FF",X"1F",X"BF",X"BF",X"BF",X"BF",X"FF",X"07",X"07",X"07",X"07",X"FF",X"FF",X"FF",
		X"FF",X"07",X"07",X"07",X"07",X"FF",X"FF",X"FF",X"FF",X"07",X"07",X"07",X"07",X"FF",X"FF",X"FF",
		X"FF",X"07",X"07",X"07",X"07",X"FF",X"FF",X"FF",X"FF",X"07",X"07",X"07",X"07",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",
		X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",
		X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",
		X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",
		X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"36",X"63",X"63",X"7F",X"63",X"63",
		X"00",X"7E",X"63",X"63",X"7E",X"63",X"63",X"7E",X"00",X"1E",X"33",X"60",X"60",X"60",X"33",X"1E",
		X"00",X"7C",X"66",X"63",X"63",X"63",X"66",X"7C",X"00",X"7E",X"60",X"60",X"7C",X"60",X"60",X"7F",
		X"00",X"7F",X"60",X"60",X"7E",X"60",X"60",X"60",X"00",X"1F",X"30",X"60",X"67",X"63",X"33",X"1F",
		X"00",X"63",X"63",X"63",X"7F",X"63",X"63",X"63",X"00",X"7E",X"18",X"18",X"18",X"18",X"18",X"7E",
		X"00",X"03",X"03",X"03",X"03",X"03",X"63",X"3C",X"00",X"63",X"66",X"6C",X"78",X"7C",X"6E",X"67",
		X"00",X"60",X"60",X"60",X"60",X"60",X"60",X"7F",X"00",X"63",X"77",X"7F",X"7F",X"6B",X"63",X"63",
		X"00",X"63",X"73",X"7B",X"7F",X"6F",X"67",X"63",X"00",X"3E",X"63",X"63",X"63",X"63",X"63",X"3E",
		X"00",X"7E",X"63",X"63",X"63",X"7E",X"60",X"60",X"00",X"3E",X"63",X"63",X"63",X"6B",X"67",X"3D",
		X"00",X"7E",X"63",X"63",X"67",X"7C",X"6E",X"67",X"00",X"3C",X"66",X"60",X"3E",X"03",X"63",X"3E",
		X"00",X"7E",X"18",X"18",X"18",X"18",X"18",X"18",X"00",X"63",X"63",X"63",X"63",X"63",X"63",X"3E",
		X"00",X"63",X"63",X"63",X"77",X"3E",X"1C",X"08",X"00",X"63",X"63",X"6B",X"7F",X"7F",X"77",X"63",
		X"00",X"63",X"77",X"3E",X"1C",X"3E",X"77",X"63",X"00",X"66",X"66",X"66",X"3C",X"18",X"18",X"18",
		X"00",X"7E",X"7E",X"0C",X"18",X"30",X"7E",X"7E",X"03",X"07",X"06",X"0C",X"08",X"00",X"60",X"60",
		X"3C",X"42",X"99",X"A1",X"A5",X"99",X"42",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"50",X"50",X"50",X"50",X"50",X"50",X"40",X"40",
		X"00",X"00",X"00",X"00",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"F8",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",
		X"00",X"33",X"73",X"73",X"00",X"00",X"00",X"00",X"7E",X"7F",X"7F",X"3F",X"1F",X"0F",X"1F",X"0F",
		X"00",X"00",X"80",X"80",X"C0",X"C1",X"E1",X"E3",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"1F",X"01",X"03",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"80",X"E0",X"F8",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"0F",X"3F",X"FF",X"FF",X"FF",X"FF",X"0F",X"07",X"07",X"C7",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"F0",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"66",X"00",X"00",X"C0",X"E0",X"F0",X"F0",X"F8",
		X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"70",
		X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"67",X"03",X"01",X"03",X"03",X"00",X"01",X"03",
		X"66",X"00",X"00",X"03",X"07",X"1F",X"3F",X"3F",X"C0",X"C0",X"E1",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"C3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"C0",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"F8",X"FF",X"FF",X"FF",X"FF",
		X"00",X"03",X"0F",X"3F",X"FF",X"FF",X"FF",X"FF",X"C0",X"F1",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"01",X"C7",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C7",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"C0",X"C0",X"C0",X"80",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"7E",X"FE",
		X"FC",X"FC",X"FC",X"FC",X"F8",X"F8",X"F8",X"F8",X"FC",X"FC",X"FC",X"FC",X"F8",X"F8",X"F8",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"3F",X"3F",X"3F",X"7E",X"7E",X"7E",X"7E",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"E0",
		X"00",X"00",X"C0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"80",X"80",X"C0",X"C0",X"E0",X"F0",X"F8",X"F8",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"01",X"0F",X"1F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"03",X"03",X"07",X"0F",X"0F",X"0F",X"0F",X"1F",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"C0",X"F0",X"FC",X"FE",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"C0",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"01",X"01",X"03",X"07",X"0F",X"0F",X"0F",X"9F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"03",X"07",X"0F",X"0F",X"1F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"F0",X"F0",X"F0",X"F8",X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",
		X"80",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"80",X"81",X"81",X"C3",X"E7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"01",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"03",
		X"07",X"07",X"0F",X"1F",X"3F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"1F",X"1F",X"3F",X"3F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"F0",X"F0",X"F0",X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"98",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"03",X"03",X"07",X"07",X"0F",X"1F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"01",X"0F",X"0F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"1F",X"3F",X"3F",X"3F",X"3F",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"1F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"F8",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"0F",X"3F",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"03",X"1F",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"C0",X"FC",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"E1",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"07",X"3F",X"FF",X"FF",X"FF",X"FF",X"80",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"F8",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"7F",X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"E0",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"80",X"E0",X"F8",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"C3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"F0",X"FF",X"FF",
		X"00",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"F0",X"FF",X"FF",X"FF",X"FF",X"00",X"3E",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"03",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"0F",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"C3",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"C7",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"03",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"01",X"01",X"01",X"01",X"03",X"03",X"03",X"03",X"07",X"07",X"07",X"07",X"0F",X"0F",X"0F",X"0F",
		X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",X"3F",X"3F",X"7E",X"7E",X"7E",X"7E",X"FC",X"FC",X"FC",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"F8",X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"CF",X"CF",X"C7",X"C7",X"83",X"83",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"0F",X"0F",
		X"BF",X"BF",X"FF",X"FF",X"FD",X"FD",X"F1",X"F1",X"C3",X"C3",X"03",X"03",X"07",X"07",X"07",X"07",
		X"0F",X"0F",X"0F",X"0F",X"1F",X"1F",X"1F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"3F",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"FC",X"FC",X"F8",X"F8",X"F8",X"F8",
		X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"07",X"0F",X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",X"3F",X"3F",X"7E",X"7E",X"7E",X"7E",
		X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"3F",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E1",
		X"80",X"00",X"00",X"00",X"01",X"01",X"01",X"03",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F8",X"FC",X"FC",X"FE",X"FE",X"FE",X"FE",
		X"F0",X"F0",X"F0",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"01",X"03",X"07",X"07",X"07",X"07",
		X"3F",X"3F",X"3F",X"1F",X"1F",X"1F",X"0F",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"E0",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"80",
		X"C3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",
		X"3F",X"3F",X"3F",X"3F",X"7E",X"7E",X"7E",X"FE",X"FC",X"FC",X"FC",X"FC",X"F8",X"F0",X"E0",X"80",
		X"00",X"00",X"00",X"00",X"81",X"81",X"81",X"81",X"03",X"03",X"03",X"03",X"07",X"07",X"07",X"07",
		X"FC",X"FC",X"FD",X"FF",X"FF",X"FF",X"FC",X"F8",X"3C",X"FF",X"FF",X"FF",X"FF",X"0F",X"07",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"E0",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",
		X"E0",X"E0",X"E0",X"E0",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"01",X"03",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"C0",X"F0",X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"FC",X"FC",X"F8",X"F8",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"07",X"0F",X"0F",X"0F",X"0F",X"7F",X"7F",X"7F",X"3F",X"3F",X"3F",X"1F",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",
		X"C0",X"80",X"80",X"80",X"00",X"00",X"00",X"01",X"87",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E7",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"FC",X"FC",
		X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"07",X"07",X"07",X"07",
		X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"3F",X"3F",X"3F",X"3F",X"7E",X"7E",X"7E",X"7E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"E0",X"E0",
		X"F8",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"87",X"9F",X"BF",X"FF",X"FF",X"FF",X"C0",X"00",
		X"80",X"80",X"81",X"03",X"07",X"07",X"07",X"07",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"FC",X"FC");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
