library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity bootrom is
    generic(
        AddrWidth   : integer := 14
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(AddrWidth-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end bootrom;

architecture rtl of bootrom is
    signal romAddr : integer range 0 to 2**AddrWidth-1;
    type rom16384x8 is array (0 to 2**AddrWidth-1) of std_logic_vector(7 downto 0); 
    constant romData : rom16384x8 := (
         x"31",  x"c0",  x"eb",  x"21",  x"8c",  x"00",  x"11",  x"00", -- 0000
         x"f0",  x"cd",  x"2c",  x"00",  x"21",  x"dc",  x"0e",  x"11", -- 0008
         x"00",  x"c0",  x"cd",  x"2c",  x"00",  x"21",  x"a6",  x"31", -- 0010
         x"11",  x"00",  x"80",  x"cd",  x"2c",  x"00",  x"01",  x"07", -- 0018
         x"00",  x"11",  x"00",  x"ec",  x"21",  x"85",  x"00",  x"ed", -- 0020
         x"b0",  x"c3",  x"00",  x"ec",  x"3e",  x"80",  x"d9",  x"11", -- 0028
         x"01",  x"00",  x"d9",  x"cd",  x"7f",  x"00",  x"38",  x"04", -- 0030
         x"ed",  x"a0",  x"18",  x"f7",  x"4e",  x"23",  x"06",  x"00", -- 0038
         x"cb",  x"79",  x"28",  x"10",  x"cd",  x"7f",  x"00",  x"cd", -- 0040
         x"7d",  x"00",  x"cd",  x"7d",  x"00",  x"cd",  x"7d",  x"00", -- 0048
         x"38",  x"02",  x"cb",  x"b9",  x"03",  x"d9",  x"62",  x"6b", -- 0050
         x"43",  x"d9",  x"cd",  x"7f",  x"00",  x"d9",  x"30",  x"0a", -- 0058
         x"04",  x"18",  x"f6",  x"d9",  x"cd",  x"7f",  x"00",  x"d9", -- 0060
         x"ed",  x"6a",  x"10",  x"f7",  x"23",  x"d9",  x"d8",  x"e5", -- 0068
         x"d9",  x"e5",  x"d9",  x"62",  x"6b",  x"ed",  x"42",  x"c1", -- 0070
         x"ed",  x"b0",  x"e1",  x"18",  x"b6",  x"cb",  x"10",  x"87", -- 0078
         x"c0",  x"7e",  x"23",  x"17",  x"c9",  x"3e",  x"01",  x"d3", -- 0080
         x"02",  x"c3",  x"00",  x"80",  x"04",  x"c3",  x"64",  x"f6", -- 0088
         x"c3",  x"ae",  x"02",  x"56",  x"12",  x"f7",  x"c3",  x"7f", -- 0090
         x"02",  x"83",  x"02",  x"29",  x"9e",  x"f7",  x"0e",  x"02", -- 0098
         x"a8",  x"02",  x"20",  x"c4",  x"02",  x"de",  x"f5",  x"c3", -- 00A0
         x"0b",  x"12",  x"f8",  x"c3",  x"fc",  x"08",  x"df",  x"02", -- 00A8
         x"09",  x"34",  x"f4",  x"c3",  x"6f",  x"02",  x"a4",  x"08", -- 00B0
         x"27",  x"33",  x"02",  x"37",  x"1a",  x"09",  x"d2",  x"05", -- 00B8
         x"d9",  x"02",  x"22",  x"e5",  x"02",  x"f4",  x"f7",  x"43", -- 00C0
         x"00",  x"09",  x"f0",  x"0c",  x"f0",  x"15",  x"f0",  x"12", -- 00C8
         x"f0",  x"00",  x"0f",  x"f0",  x"18",  x"f0",  x"39",  x"f0", -- 00D0
         x"3c",  x"f0",  x"00",  x"e2",  x"f3",  x"65",  x"f3",  x"06", -- 00D8
         x"f0",  x"f3",  x"f3",  x"00",  x"f8",  x"f3",  x"2d",  x"f4", -- 00E0
         x"45",  x"f4",  x"6a",  x"f4",  x"08",  x"3c",  x"f7",  x"3b", -- 00E8
         x"f7",  x"33",  x"27",  x"f0",  x"00",  x"2a",  x"f0",  x"1e", -- 00F0
         x"f0",  x"21",  x"f0",  x"a8",  x"f4",  x"00",  x"e3",  x"fa", -- 00F8
         x"24",  x"f0",  x"3f",  x"f0",  x"42",  x"f0",  x"02",  x"3e", -- 0100
         x"f7",  x"3d",  x"f7",  x"b9",  x"f5",  x"19",  x"00",  x"d8", -- 0108
         x"f4",  x"21",  x"89",  x"f0",  x"e5",  x"21",  x"80",  x"00", -- 0110
         x"00",  x"22",  x"1b",  x"00",  x"3e",  x"3e",  x"cd",  x"05", -- 0118
         x"00",  x"f3",  x"cd",  x"5c",  x"f3",  x"38",  x"23",  x"cd", -- 0120
         x"b9",  x"80",  x"18",  x"21",  x"ea",  x"f5",  x"e5",  x"cd", -- 0128
         x"ea",  x"00",  x"f1",  x"ca",  x"e6",  x"f5",  x"c5",  x"cd", -- 0130
         x"8e",  x"f2",  x"04",  x"c1",  x"28",  x"07",  x"cd",  x"26", -- 0138
         x"14",  x"2a",  x"00",  x"71",  x"00",  x"e9",  x"08",  x"30", -- 0140
         x"2a",  x"cd",  x"fe",  x"22",  x"f2",  x"da",  x"bc",  x"00", -- 0148
         x"06",  x"04",  x"21",  x"e9",  x"ef",  x"11",  x"d5",  x"fb", -- 0150
         x"46",  x"cd",  x"74",  x"3e",  x"3a",  x"3a",  x"02",  x"d5", -- 0158
         x"5e",  x"23",  x"56",  x"23",  x"33",  x"85",  x"0d",  x"e1", -- 0160
         x"d1",  x"13",  x"00",  x"23",  x"83",  x"10",  x"e5",  x"c9", -- 0168
         x"41",  x"03",  x"28",  x"2c",  x"08",  x"da",  x"44",  x"0b", -- 0170
         x"01",  x"09",  x"2e",  x"2b",  x"00",  x"b8",  x"f2",  x"58", -- 0178
         x"c1",  x"20",  x"50",  x"02",  x"3e",  x"04",  x"93",  x"87", -- 0180
         x"32",  x"33",  x"74",  x"00",  x"40",  x"00",  x"79",  x"fe", -- 0188
         x"3a",  x"20",  x"05",  x"cd",  x"01",  x"c4",  x"f1",  x"fe", -- 0190
         x"3d",  x"c2",  x"e2",  x"f5",  x"2d",  x"a9",  x"5b",  x"6e", -- 0198
         x"b2",  x"6e",  x"80",  x"17",  x"cd",  x"ab",  x"f0",  x"d8", -- 01A0
         x"00",  x"00",  x"e5",  x"d5",  x"7c",  x"84",  x"85",  x"87", -- 01A8
         x"16",  x"00",  x"00",  x"5f",  x"21",  x"c9",  x"ef",  x"19", -- 01B0
         x"71",  x"23",  x"02",  x"70",  x"d1",  x"e1",  x"3a",  x"04", -- 01B8
         x"00",  x"80",  x"22",  x"37",  x"3a",  x"3b",  x"00",  x"47", -- 01C0
         x"4d",  x"bc",  x"28",  x"0a",  x"95",  x"3c",  x"fe",  x"00", -- 01C8
         x"06",  x"28",  x"04",  x"3d",  x"b8",  x"20",  x"25",  x"d5", -- 01D0
         x"20",  x"58",  x"21",  x"19",  x"06",  x"09",  x"3c",  x"cb", -- 01D8
         x"02",  x"1e",  x"3d",  x"20",  x"07",  x"cb",  x"39",  x"06", -- 01E0
         x"80",  x"03",  x"05",  x"10",  x"f2",  x"43",  x"cd",  x"ce", -- 01E8
         x"02",  x"f2",  x"d1",  x"30",  x"0b",  x"08",  x"32",  x"1b", -- 01F0
         x"84",  x"72",  x"37",  x"c9",  x"c3",  x"87",  x"48",  x"2a", -- 01F8
         x"72",  x"73",  x"23",  x"00",  x"72",  x"c3",  x"bd",  x"f0", -- 0200
         x"08",  x"38",  x"34",  x"06",  x"02",  x"03",  x"3e",  x"17", -- 0208
         x"32",  x"2f",  x"00",  x"70",  x"a2",  x"76",  x"93",  x"08", -- 0210
         x"e3",  x"d8",  x"5f",  x"3a",  x"0b",  x"bb",  x"3e",  x"04", -- 0218
         x"03",  x"d8",  x"4d",  x"6c",  x"63",  x"1c",  x"10",  x"04", -- 0220
         x"3e",  x"3b",  x"10",  x"e3",  x"c3",  x"92",  x"44",  x"22", -- 0228
         x"1e",  x"a2",  x"40",  x"32",  x"1d",  x"00",  x"b7",  x"c9", -- 0230
         x"51",  x"1e",  x"77",  x"cf",  x"48",  x"e4",  x"11",  x"12", -- 0238
         x"01",  x"01",  x"cd",  x"c6",  x"46",  x"e4",  x"22",  x"c3", -- 0240
         x"df",  x"00",  x"21",  x"81",  x"00",  x"23",  x"7e",  x"fe", -- 0248
         x"20",  x"28",  x"00",  x"fa",  x"cd",  x"d7",  x"f1",  x"4f", -- 0250
         x"c0",  x"fe",  x"01",  x"00",  x"d8",  x"bf",  x"c9",  x"7e", -- 0258
         x"b7",  x"c8",  x"e5",  x"c5",  x"00",  x"21",  x"ab",  x"fc", -- 0260
         x"01",  x"05",  x"00",  x"ed",  x"b1",  x"00",  x"c1",  x"e1", -- 0268
         x"36",  x"20",  x"23",  x"c9",  x"11",  x"52",  x"00",  x"01", -- 0270
         x"af",  x"06",  x"51",  x"12",  x"1b",  x"10",  x"fc",  x"46", -- 0278
         x"e5",  x"e7",  x"00",  x"38",  x"0d",  x"28",  x"0b",  x"12", -- 0280
         x"04",  x"13",  x"c0",  x"31",  x"20",  x"f8",  x"cd",  x"d0", -- 0288
         x"00",  x"f1",  x"78",  x"32",  x"00",  x"01",  x"79",  x"e1", -- 0290
         x"08",  x"41",  x"3a",  x"55",  x"fe",  x"30",  x"38",  x"16", -- 0298
         x"8b",  x"21",  x"30",  x"12",  x"3e",  x"21",  x"11",  x"12", -- 02A0
         x"cd",  x"15",  x"f8",  x"3c",  x"12",  x"38",  x"02",  x"4f", -- 02A8
         x"bf",  x"82",  x"30",  x"fe",  x"40",  x"22",  x"38",  x"f8", -- 02B0
         x"bb",  x"82",  x"17",  x"cd",  x"4d",  x"f2",  x"f5",  x"d5", -- 02B8
         x"23",  x"18",  x"06",  x"09",  x"90",  x"cd",  x"69",  x"f2", -- 02C0
         x"f1",  x"80",  x"23",  x"f5",  x"b7",  x"ed",  x"52",  x"f1", -- 02C8
         x"c9",  x"88",  x"31",  x"04",  x"af",  x"07",  x"3c",  x"30", -- 02D0
         x"01",  x"fb",  x"21",  x"c1",  x"ef",  x"d6",  x"08",  x"23", -- 02D8
         x"07",  x"02",  x"c6",  x"08",  x"2b",  x"28",  x"fb",  x"8d", -- 02E0
         x"40",  x"cb",  x"16",  x"3d",  x"c8",  x"21",  x"10",  x"fa", -- 02E8
         x"3a",  x"d5",  x"eb",  x"1a",  x"a6",  x"18",  x"04",  x"c0", -- 02F0
         x"48",  x"02",  x"e6",  x"df",  x"be",  x"00",  x"13",  x"23", -- 02F8
         x"20",  x"0c",  x"10",  x"ee",  x"d1",  x"d1",  x"00",  x"6b", -- 0300
         x"62",  x"2b",  x"7e",  x"2b",  x"6e",  x"67",  x"c9",  x"90", -- 0308
         x"d4",  x"c9",  x"21",  x"44",  x"00",  x"9c",  x"3e",  x"01", -- 0310
         x"c3",  x"ed",  x"a1",  x"20",  x"12",  x"23",  x"23",  x"a9", -- 0318
         x"32",  x"0b",  x"7f",  x"9a",  x"a6",  x"82",  x"60",  x"0c", -- 0320
         x"af",  x"2b",  x"2b",  x"04",  x"be",  x"20",  x"e8",  x"e1", -- 0328
         x"25",  x"9b",  x"80",  x"24",  x"c9",  x"c1",  x"c9",  x"01", -- 0330
         x"04",  x"06",  x"02",  x"21",  x"26",  x"fc",  x"ff",  x"60", -- 0338
         x"c5",  x"41",  x"05",  x"99",  x"b1",  x"6c",  x"20",  x"09", -- 0340
         x"c8",  x"79",  x"23",  x"eb",  x"00",  x"fc",  x"10",  x"f0", -- 0348
         x"f6",  x"01",  x"c9",  x"4c",  x"f5",  x"a2",  x"58",  x"27", -- 0350
         x"78",  x"b7",  x"9b",  x"22",  x"64",  x"cb",  x"3f",  x"e8", -- 0358
         x"20",  x"cb",  x"23",  x"e6",  x"03",  x"4e",  x"83",  x"b3", -- 0360
         x"85",  x"f1",  x"19",  x"19",  x"e5",  x"95",  x"20",  x"21", -- 0368
         x"ff",  x"ff",  x"02",  x"eb",  x"cd",  x"bc",  x"fc",  x"d1", -- 0370
         x"3f",  x"8a",  x"30",  x"c5",  x"ed",  x"05",  x"b0",  x"18", -- 0378
         x"0e",  x"3e",  x"0d",  x"af",  x"21",  x"3e",  x"0a",  x"0d", -- 0380
         x"85",  x"4f",  x"cd",  x"fc",  x"48",  x"c1",  x"81",  x"c0", -- 0388
         x"3e",  x"20",  x"18",  x"f1",  x"00",  x"ed",  x"73",  x"0b", -- 0390
         x"00",  x"31",  x"c0",  x"01",  x"37",  x"40",  x"3f",  x"17", -- 0398
         x"f5",  x"ed",  x"43",  x"0d",  x"00",  x"02",  x"32",  x"0f", -- 03A0
         x"00",  x"21",  x"45",  x"f3",  x"98",  x"21",  x"21",  x"b9", -- 03A8
         x"da",  x"a9",  x"53",  x"06",  x"0b",  x"00",  x"f0",  x"09", -- 03B0
         x"09",  x"7e",  x"23",  x"66",  x"08",  x"6f",  x"4b",  x"42", -- 03B8
         x"3a",  x"19",  x"e5",  x"2e",  x"05",  x"03",  x"c9",  x"30", -- 03C0
         x"06",  x"cd",  x"a5",  x"45",  x"f1",  x"37",  x"02",  x"97", -- 03C8
         x"49",  x"11",  x"11",  x"ed",  x"4b",  x"32",  x"ed",  x"7b", -- 03D0
         x"42",  x"48",  x"8e",  x"80",  x"98",  x"ed",  x"50",  x"12", -- 03D8
         x"c8",  x"11",  x"e1",  x"81",  x"23",  x"4d",  x"44",  x"03", -- 03E0
         x"36",  x"48",  x"29",  x"35",  x"c9",  x"24",  x"b5",  x"6a", -- 03E8
         x"7f",  x"69",  x"d8",  x"ed",  x"a0",  x"17",  x"00",  x"34", -- 03F0
         x"35",  x"00",  x"e1",  x"20",  x"2b",  x"fe",  x"03",  x"20", -- 03F8
         x"03",  x"af",  x"90",  x"d8",  x"fe",  x"1f",  x"05",  x"28", -- 0400
         x"1b",  x"fe",  x"02",  x"20",  x"df",  x"40",  x"c6",  x"f3", -- 0408
         x"20",  x"fb",  x"18",  x"26",  x"d7",  x"fe",  x"a0",  x"00", -- 0410
         x"20",  x"fe",  x"0b",  x"28",  x"cf",  x"fe",  x"0a",  x"28", -- 0418
         x"15",  x"cb",  x"fe",  x"08",  x"9b",  x"90",  x"16",  x"18", -- 0420
         x"c2",  x"fe",  x"02",  x"10",  x"28",  x"03",  x"34",  x"02", -- 0428
         x"03",  x"b4",  x"30",  x"d8",  x"1a",  x"90",  x"92",  x"b3", -- 0430
         x"3a",  x"46",  x"35",  x"9b",  x"d2",  x"81",  x"40",  x"47", -- 0438
         x"c8",  x"0b",  x"0a",  x"fe",  x"09",  x"92",  x"aa",  x"de", -- 0440
         x"40",  x"38",  x"f4",  x"3e",  x"08",  x"b5",  x"bf",  x"38", -- 0448
         x"10",  x"f3",  x"07",  x"01",  x"35",  x"c9",  x"1a",  x"b7", -- 0450
         x"20",  x"06",  x"3a",  x"6a",  x"50",  x"90",  x"af",  x"d0", -- 0458
         x"36",  x"13",  x"18",  x"ef",  x"21",  x"00",  x"03",  x"01", -- 0460
         x"18",  x"38",  x"cd",  x"93",  x"f5",  x"3c",  x"88",  x"82", -- 0468
         x"af",  x"32",  x"17",  x"6c",  x"00",  x"cd",  x"da",  x"2d", -- 0470
         x"e1",  x"f5",  x"24",  x"0c",  x"11",  x"be",  x"c2",  x"19", -- 0478
         x"11",  x"6d",  x"f4",  x"62",  x"08",  x"00",  x"9a",  x"41", -- 0480
         x"d1",  x"21",  x"5c",  x"c5",  x"52",  x"0b",  x"dd",  x"52", -- 0488
         x"a1",  x"40",  x"37",  x"c0",  x"3a",  x"73",  x"c1",  x"3d", -- 0490
         x"32",  x"c0",  x"ef",  x"9e",  x"34",  x"1d",  x"22",  x"8a", -- 0498
         x"db",  x"cc",  x"cb",  x"ad",  x"98",  x"d8",  x"31",  x"21", -- 04A0
         x"93",  x"3b",  x"34",  x"fe",  x"53",  x"67",  x"f7",  x"73", -- 04A8
         x"4c",  x"32",  x"97",  x"bd",  x"b1",  x"92",  x"22",  x"73", -- 04B0
         x"43",  x"70",  x"17",  x"5a",  x"4d",  x"6b",  x"0b",  x"02", -- 04B8
         x"5f",  x"71",  x"72",  x"5f",  x"d9",  x"23",  x"ff",  x"11", -- 04C0
         x"09",  x"01",  x"a0",  x"5c",  x"5b",  x"0c",  x"24",  x"3a", -- 04C8
         x"4c",  x"b7",  x"a2",  x"c4",  x"3e",  x"09",  x"f5",  x"49", -- 04D0
         x"2a",  x"95",  x"04",  x"d5",  x"11",  x"7f",  x"14",  x"52", -- 04D8
         x"4e",  x"d1",  x"98",  x"4c",  x"89",  x"38",  x"4c",  x"ed", -- 04E0
         x"a0",  x"3b",  x"2a",  x"f2",  x"30",  x"a1",  x"36",  x"d6", -- 04E8
         x"fe",  x"61",  x"30",  x"46",  x"7e",  x"e0",  x"18",  x"34", -- 04F0
         x"c3",  x"ae",  x"15",  x"d5",  x"01",  x"fc",  x"09",  x"16", -- 04F8
         x"03",  x"21",  x"f5",  x"80",  x"e5",  x"2b",  x"36",  x"3a", -- 0500
         x"23",  x"0a",  x"40",  x"c5",  x"3e",  x"07",  x"47",  x"af", -- 0508
         x"c6",  x"01",  x"00",  x"27",  x"10",  x"fb",  x"77",  x"3e", -- 0510
         x"33",  x"ed",  x"67",  x"10",  x"23",  x"77",  x"23",  x"48", -- 0518
         x"c1",  x"03",  x"15",  x"2e",  x"20",  x"e2",  x"f4",  x"06", -- 0520
         x"0e",  x"08",  x"c3",  x"f7",  x"f2",  x"57",  x"71",  x"56", -- 0528
         x"6d",  x"bc",  x"59",  x"36",  x"d8",  x"58",  x"71",  x"26", -- 0530
         x"30",  x"1d",  x"a5",  x"0b",  x"cd",  x"59",  x"ff",  x"cd", -- 0538
         x"51",  x"d6",  x"08",  x"c0",  x"c4",  x"3a",  x"61",  x"be", -- 0540
         x"40",  x"e1",  x"74",  x"28",  x"09",  x"fe",  x"ff",  x"28", -- 0548
         x"08",  x"05",  x"f1",  x"3e",  x"0b",  x"90",  x"a3",  x"04", -- 0550
         x"0c",  x"d8",  x"15",  x"11",  x"3c",  x"c7",  x"0c",  x"20", -- 0558
         x"01",  x"3c",  x"7c",  x"c5",  x"ba",  x"12",  x"c8",  x"21", -- 0560
         x"e6",  x"2d",  x"3a",  x"bc",  x"29",  x"e1",  x"08",  x"d0", -- 0568
         x"11",  x"e4",  x"a5",  x"d7",  x"0b",  x"88",  x"f5",  x"fc", -- 0570
         x"a0",  x"66",  x"21",  x"43",  x"4f",  x"22",  x"40",  x"64", -- 0578
         x"0e",  x"4d",  x"32",  x"66",  x"00",  x"18",  x"60",  x"16", -- 0580
         x"c0",  x"2e",  x"62",  x"e1",  x"ba",  x"66",  x"ab",  x"ae", -- 0588
         x"c8",  x"bc",  x"16",  x"b8",  x"d8",  x"11",  x"19",  x"26", -- 0590
         x"58",  x"d2",  x"d2",  x"c4",  x"ce",  x"d0",  x"85",  x"30", -- 0598
         x"09",  x"06",  x"b7",  x"37",  x"c8",  x"cd",  x"a3",  x"b9", -- 05A0
         x"48",  x"18",  x"99",  x"92",  x"6d",  x"a6",  x"b2",  x"f5", -- 05A8
         x"86",  x"30",  x"05",  x"10",  x"a2",  x"af",  x"c9",  x"be", -- 05B0
         x"c3",  x"22",  x"d9",  x"2a",  x"47",  x"7e",  x"f5",  x"5a", -- 05B8
         x"13",  x"a6",  x"0b",  x"11",  x"48",  x"fc",  x"d7",  x"cd", -- 05C0
         x"80",  x"44",  x"2a",  x"26",  x"d0",  x"92",  x"b5",  x"80", -- 05C8
         x"32",  x"41",  x"54",  x"99",  x"28",  x"c7",  x"95",  x"7f", -- 05D0
         x"93",  x"45",  x"c0",  x"0e",  x"95",  x"86",  x"31",  x"f2", -- 05D8
         x"87",  x"04",  x"13",  x"1a",  x"38",  x"1e",  x"a1",  x"d8", -- 05E0
         x"e5",  x"32",  x"00",  x"47",  x"0e",  x"00",  x"eb",  x"3e", -- 05E8
         x"1f",  x"be",  x"80",  x"4e",  x"ed",  x"a0",  x"03",  x"03", -- 05F0
         x"2b",  x"23",  x"41",  x"10",  x"74",  x"71",  x"eb",  x"79", -- 05F8
         x"b7",  x"ff",  x"12",  x"c0",  x"cc",  x"23",  x"3e",  x"07", -- 0600
         x"03",  x"18",  x"02",  x"03",  x"01",  x"91",  x"03",  x"d0", -- 0608
         x"e2",  x"45",  x"82",  x"d0",  x"19",  x"88",  x"18",  x"f5", -- 0610
         x"99",  x"9c",  x"15",  x"81",  x"14",  x"74",  x"f1",  x"01", -- 0618
         x"11",  x"5b",  x"fc",  x"d6",  x"05",  x"30",  x"0c",  x"5f", -- 0620
         x"42",  x"6f",  x"f1",  x"c6",  x"35",  x"9f",  x"90",  x"18", -- 0628
         x"4d",  x"02",  x"d6",  x"02",  x"d8",  x"f5",  x"11",  x"56", -- 0630
         x"81",  x"37",  x"cc",  x"58",  x"9d",  x"df",  x"02",  x"20", -- 0638
         x"04",  x"06",  x"08",  x"18",  x"03",  x"e3",  x"c0",  x"0f", -- 0640
         x"21",  x"cc",  x"fb",  x"00",  x"11",  x"09",  x"00",  x"cb", -- 0648
         x"38",  x"04",  x"19",  x"10",  x"00",  x"fd",  x"eb",  x"18", -- 0650
         x"1f",  x"11",  x"62",  x"fc",  x"3d",  x"50",  x"28",  x"b2", -- 0658
         x"73",  x"c1",  x"05",  x"13",  x"11",  x"81",  x"05",  x"83", -- 0660
         x"0d",  x"11",  x"92",  x"05",  x"06",  x"07",  x"11",  x"9d", -- 0668
         x"05",  x"11",  x"01",  x"1b",  x"c4",  x"b5",  x"63",  x"d9", -- 0670
         x"60",  x"f3",  x"31",  x"00",  x"45",  x"02",  x"a3",  x"91", -- 0678
         x"38",  x"5d",  x"0a",  x"54",  x"13",  x"06",  x"01",  x"dc", -- 0680
         x"22",  x"91",  x"01",  x"ed",  x"47",  x"3c",  x"d3",  x"8a", -- 0688
         x"3e",  x"cf",  x"03",  x"22",  x"af",  x"02",  x"d3",  x"88", -- 0690
         x"f5",  x"f0",  x"06",  x"40",  x"05",  x"7e",  x"2f",  x"77", -- 0698
         x"56",  x"ba",  x"03",  x"dd",  x"10",  x"28",  x"06",  x"0d", -- 06A0
         x"24",  x"2b",  x"22",  x"2b",  x"23",  x"e5",  x"60",  x"10", -- 06A8
         x"ea",  x"21",  x"08",  x"14",  x"f3",  x"22",  x"06",  x"aa", -- 06B0
         x"82",  x"e0",  x"f6",  x"11",  x"30",  x"92",  x"37",  x"49", -- 06B8
         x"70",  x"9f",  x"ca",  x"ab",  x"e3",  x"85",  x"05",  x"9c", -- 06C0
         x"1b",  x"f9",  x"0b",  x"22",  x"01",  x"00",  x"eb",  x"c2", -- 06C8
         x"e6",  x"fc",  x"f9",  x"e0",  x"cd",  x"12",  x"f7",  x"11", -- 06D0
         x"72",  x"f7",  x"81",  x"92",  x"21",  x"23",  x"dd",  x"29", -- 06D8
         x"82",  x"30",  x"84",  x"b9",  x"ac",  x"1c",  x"c2",  x"d2", -- 06E0
         x"2f",  x"e9",  x"fc",  x"00",  x"11",  x"ca",  x"ef",  x"01", -- 06E8
         x"1f",  x"00",  x"2a",  x"36",  x"ff",  x"78",  x"e0",  x"b0", -- 06F0
         x"ba",  x"08",  x"b0",  x"fc",  x"0e",  x"0c",  x"09",  x"21", -- 06F8
         x"24",  x"02",  x"fc",  x"22",  x"eb",  x"ef",  x"22",  x"ed", -- 0700
         x"02",  x"58",  x"ef",  x"8f",  x"b4",  x"09",  x"f7",  x"22", -- 0708
         x"cd",  x"ef",  x"92",  x"15",  x"27",  x"55",  x"96",  x"52", -- 0710
         x"a9",  x"6e",  x"a3",  x"62",  x"df",  x"10",  x"22",  x"e9", -- 0718
         x"17",  x"f1",  x"f8",  x"22",  x"40",  x"cb",  x"20",  x"e3", -- 0720
         x"ef",  x"ed",  x"5e",  x"11",  x"c0",  x"b8",  x"1b",  x"7b", -- 0728
         x"5d",  x"b2",  x"96",  x"b6",  x"28",  x"3d",  x"00",  x"e9", -- 0730
         x"2e",  x"07",  x"18",  x"07",  x"2e",  x"05",  x"59",  x"20", -- 0738
         x"50",  x"2c",  x"00",  x"7d",  x"cd",  x"58",  x"f7",  x"5c", -- 0740
         x"d8",  x"bf",  x"c8",  x"bb",  x"dd",  x"ff",  x"65",  x"d0", -- 0748
         x"9a",  x"a0",  x"fe",  x"04",  x"c8",  x"09",  x"ed",  x"53", -- 0750
         x"bc",  x"01",  x"ef",  x"2c",  x"bc",  x"d9",  x"ce",  x"d5", -- 0758
         x"f4",  x"bc",  x"14",  x"04",  x"c1",  x"af",  x"28",  x"c9", -- 0760
         x"ea",  x"1b",  x"6f",  x"f7",  x"e3",  x"e2",  x"80",  x"e9", -- 0768
         x"c1",  x"4f",  x"38",  x"f0",  x"dc",  x"de",  x"b9",  x"e7", -- 0770
         x"d0",  x"cd",  x"b4",  x"8a",  x"e4",  x"98",  x"e0",  x"18", -- 0778
         x"d5",  x"79",  x"b9",  x"d5",  x"20",  x"f9",  x"a4",  x"59", -- 0780
         x"ee",  x"a9",  x"7a",  x"04",  x"9b",  x"18",  x"c5",  x"53", -- 0788
         x"e1",  x"32",  x"4d",  x"d8",  x"10",  x"f4",  x"c8",  x"0d", -- 0790
         x"06",  x"06",  x"22",  x"18",  x"b6",  x"4d",  x"18",  x"f8", -- 0798
         x"28",  x"c8",  x"f6",  x"18",  x"ac",  x"c0",  x"0f",  x"04", -- 07A0
         x"18",  x"a6",  x"fe",  x"91",  x"a3",  x"f0",  x"cc",  x"30", -- 07A8
         x"20",  x"e4",  x"cd",  x"54",  x"aa",  x"7c",  x"9f",  x"03", -- 07B0
         x"18",  x"dc",  x"cd",  x"8f",  x"fe",  x"f3",  x"03",  x"13", -- 07B8
         x"00",  x"aa",  x"34",  x"c3",  x"e9",  x"4a",  x"fa",  x"91", -- 07C0
         x"62",  x"5a",  x"4f",  x"5f",  x"a9",  x"07",  x"5f",  x"13", -- 07C8
         x"1b",  x"05",  x"85",  x"69",  x"60",  x"fb",  x"68",  x"01", -- 07D0
         x"38",  x"01",  x"71",  x"3d",  x"74",  x"0e",  x"29",  x"4f", -- 07D8
         x"c2",  x"85",  x"3a",  x"d2",  x"98",  x"0f",  x"2a",  x"e0", -- 07E0
         x"d1",  x"4c",  x"45",  x"ce",  x"e6",  x"23",  x"0e",  x"68", -- 07E8
         x"61",  x"e7",  x"92",  x"18",  x"52",  x"1a",  x"a3",  x"40", -- 07F0
         x"6a",  x"cd",  x"36",  x"f8",  x"d8",  x"01",  x"01",  x"02", -- 07F8
         x"00",  x"1a",  x"13",  x"d6",  x"30",  x"d8",  x"85",  x"90", -- 0800
         x"3f",  x"d8",  x"80",  x"00",  x"0d",  x"c8",  x"87",  x"47", -- 0808
         x"87",  x"87",  x"80",  x"47",  x"28",  x"18",  x"ec",  x"f7", -- 0810
         x"11",  x"13",  x"be",  x"c8",  x"e2",  x"01",  x"4e",  x"38", -- 0818
         x"13",  x"77",  x"91",  x"09",  x"d5",  x"39",  x"cc",  x"a0", -- 0820
         x"b8",  x"c1",  x"eb",  x"14",  x"36",  x"30",  x"eb",  x"a4", -- 0828
         x"8d",  x"f0",  x"84",  x"b6",  x"bb",  x"d8",  x"e6",  x"30", -- 0830
         x"20",  x"69",  x"0a",  x"db",  x"86",  x"70",  x"1b",  x"79", -- 0838
         x"12",  x"0a",  x"f1",  x"18",  x"d1",  x"f1",  x"83",  x"01", -- 0840
         x"d6",  x"14",  x"38",  x"15",  x"28",  x"cc",  x"10",  x"f8", -- 0848
         x"7b",  x"a0",  x"01",  x"b1",  x"c9",  x"7b",  x"06",  x"8f", -- 0850
         x"cb",  x"21",  x"01",  x"cf",  x"c8",  x"40",  x"db",  x"88", -- 0858
         x"06",  x"c7",  x"cd",  x"28",  x"79",  x"f8",  x"85",  x"87", -- 0860
         x"27",  x"0e",  x"3a",  x"27",  x"e1",  x"9d",  x"b9",  x"5c", -- 0868
         x"8c",  x"cd",  x"27",  x"68",  x"f8",  x"8d",  x"02",  x"af", -- 0870
         x"77",  x"c9",  x"79",  x"9d",  x"a2",  x"28",  x"39",  x"53", -- 0878
         x"02",  x"05",  x"7b",  x"ee",  x"80",  x"18",  x"ed",  x"07", -- 0880
         x"3a",  x"1d",  x"f3",  x"b9",  x"e8",  x"ad",  x"0d",  x"ff", -- 0888
         x"11",  x"01",  x"30",  x"00",  x"c0",  x"38",  x"ff",  x"a6", -- 0890
         x"24",  x"ea",  x"b8",  x"97",  x"15",  x"03",  x"d3",  x"80", -- 0898
         x"42",  x"1e",  x"3f",  x"4c",  x"62",  x"0a",  x"e8",  x"b8", -- 08A0
         x"c9",  x"91",  x"c5",  x"77",  x"09",  x"34",  x"03",  x"a6", -- 08A8
         x"83",  x"2d",  x"02",  x"79",  x"77",  x"3d",  x"9a",  x"e0", -- 08B0
         x"cd",  x"7d",  x"f9",  x"3a",  x"4a",  x"16",  x"ca",  x"0c", -- 08B8
         x"18",  x"c3",  x"7b",  x"d4",  x"06",  x"fa",  x"18",  x"a7", -- 08C0
         x"f5",  x"a3",  x"3c",  x"8d",  x"ca",  x"a7",  x"32",  x"eb", -- 08C8
         x"01",  x"22",  x"3b",  x"00",  x"26",  x"29",  x"22",  x"3d", -- 08D0
         x"04",  x"51",  x"b1",  x"b4",  x"48",  x"25",  x"95",  x"02", -- 08D8
         x"13",  x"02",  x"29",  x"4c",  x"16",  x"e6",  x"38",  x"4c", -- 08E0
         x"f1",  x"24",  x"40",  x"04",  x"49",  x"3a",  x"14",  x"c9", -- 08E8
         x"06",  x"21",  x"06",  x"8f",  x"b7",  x"dc",  x"2d",  x"b4", -- 08F0
         x"22",  x"07",  x"32",  x"13",  x"02",  x"64",  x"14",  x"94", -- 08F8
         x"b7",  x"80",  x"57",  x"f1",  x"fe",  x"39",  x"30",  x"e6", -- 0900
         x"d6",  x"2e",  x"31",  x"38",  x"de",  x"c8",  x"ff",  x"3d", -- 0908
         x"ca",  x"2a",  x"8d",  x"f8",  x"e0",  x"90",  x"05",  x"33", -- 0910
         x"34",  x"ca",  x"f3",  x"f9",  x"99",  x"31",  x"08",  x"74", -- 0918
         x"f8",  x"83",  x"2b",  x"3c",  x"0b",  x"28",  x"18",  x"a1", -- 0920
         x"42",  x"3d",  x"c0",  x"6d",  x"32",  x"ec",  x"eb",  x"8b", -- 0928
         x"c0",  x"93",  x"28",  x"00",  x"f6",  x"9e",  x"04",  x"19", -- 0930
         x"2c",  x"67",  x"0e",  x"53",  x"96",  x"1f",  x"21",  x"2c", -- 0938
         x"af",  x"13",  x"34",  x"79",  x"ab",  x"c1",  x"d8",  x"28", -- 0940
         x"4e",  x"28",  x"24",  x"30",  x"02",  x"3b",  x"02",  x"53", -- 0948
         x"b4",  x"c7",  x"81",  x"02",  x"1e",  x"fe",  x"13",  x"d8", -- 0950
         x"71",  x"8f",  x"28",  x"12",  x"11",  x"18",  x"1a",  x"3a", -- 0958
         x"a7",  x"64",  x"88",  x"2c",  x"01",  x"00",  x"47",  x"3a", -- 0960
         x"3c",  x"00",  x"90",  x"47",  x"9d",  x"40",  x"4f",  x"fa", -- 0968
         x"c1",  x"45",  x"10",  x"d2",  x"b6",  x"13",  x"32",  x"3f", -- 0970
         x"23",  x"02",  x"11",  x"3e",  x"9e",  x"4e",  x"8a",  x"00", -- 0978
         x"c0",  x"1b",  x"1a",  x"3c",  x"77",  x"21",  x"58",  x"2c", -- 0980
         x"0a",  x"23",  x"3d",  x"06",  x"be",  x"d0",  x"77",  x"18", -- 0988
         x"77",  x"1a",  x"cc",  x"23",  x"35",  x"1a",  x"c1",  x"a8", -- 0990
         x"3d",  x"1a",  x"ac",  x"35",  x"46",  x"11",  x"be",  x"d8", -- 0998
         x"3c",  x"1a",  x"5d",  x"3a",  x"1a",  x"18",  x"4f",  x"3a", -- 09A0
         x"4f",  x"21",  x"d2",  x"92",  x"90",  x"32",  x"ca",  x"f1", -- 09A8
         x"41",  x"b4",  x"88",  x"fd",  x"2c",  x"22",  x"2d",  x"cb", -- 09B0
         x"09",  x"c8",  x"ef",  x"cb",  x"6f",  x"c3",  x"34",  x"f2", -- 09B8
         x"5a",  x"3f",  x"ad",  x"7e",  x"cb",  x"22",  x"e5",  x"ac", -- 09C0
         x"92",  x"0b",  x"34",  x"16",  x"27",  x"9a",  x"a9",  x"f4", -- 09C8
         x"81",  x"ae",  x"e6",  x"f0",  x"78",  x"cc",  x"c0",  x"21", -- 09D0
         x"77",  x"e1",  x"b2",  x"b7",  x"29",  x"72",  x"9f",  x"4d", -- 09D8
         x"28",  x"77",  x"27",  x"fc",  x"fc",  x"27",  x"3a",  x"34", -- 09E0
         x"0a",  x"eb",  x"be",  x"a1",  x"af",  x"f5",  x"56",  x"cc", -- 09E8
         x"b4",  x"6a",  x"4f",  x"8d",  x"34",  x"47",  x"f1",  x"dc", -- 09F0
         x"ab",  x"30",  x"01",  x"41",  x"66",  x"c1",  x"f5",  x"0a", -- 09F8
         x"78",  x"91",  x"28",  x"37",  x"0f",  x"2e",  x"98",  x"9d", -- 0A00
         x"19",  x"18",  x"c3",  x"83",  x"f2",  x"6d",  x"ad",  x"11", -- 0A08
         x"c5",  x"c8",  x"81",  x"3c",  x"47",  x"2b",  x"1b",  x"f8", -- 0A10
         x"98",  x"fc",  x"a2",  x"2e",  x"cb",  x"29",  x"91",  x"4f", -- 0A18
         x"b4",  x"3e",  x"f9",  x"a4",  x"53",  x"9f",  x"62",  x"42", -- 0A20
         x"02",  x"c1",  x"a9",  x"e3",  x"c1",  x"e1",  x"4d",  x"06", -- 0A28
         x"10",  x"ca",  x"f1",  x"28",  x"91",  x"4f",  x"47",  x"a8", -- 0A30
         x"94",  x"ee",  x"38",  x"2b",  x"28",  x"02",  x"0d",  x"36", -- 0A38
         x"20",  x"c5",  x"f5",  x"c4",  x"2d",  x"8c",  x"80",  x"c6", -- 0A40
         x"7e",  x"27",  x"96",  x"40",  x"bf",  x"77",  x"f1",  x"c1", -- 0A48
         x"c8",  x"ac",  x"8c",  x"88",  x"33",  x"c9",  x"0e",  x"0d", -- 0A50
         x"27",  x"cb",  x"22",  x"19",  x"07",  x"00",  x"e6",  x"7f", -- 0A58
         x"ee",  x"82",  x"f3",  x"f5",  x"53",  x"20",  x"fa",  x"f1", -- 0A60
         x"04",  x"15",  x"fb",  x"3e",  x"83",  x"30",  x"d3",  x"93", -- 0A68
         x"f1",  x"0a",  x"90",  x"f1",  x"fb",  x"c9",  x"b6",  x"53", -- 0A70
         x"d3",  x"82",  x"ff",  x"14",  x"80",  x"3e",  x"06",  x"c7", -- 0A78
         x"d3",  x"83",  x"3e",  x"40",  x"03",  x"23",  x"27",  x"10", -- 0A80
         x"3e",  x"96",  x"03",  x"3e",  x"cf",  x"cc",  x"99",  x"2b", -- 0A88
         x"92",  x"af",  x"02",  x"b8",  x"ac",  x"2e",  x"0a",  x"98", -- 0A90
         x"03",  x"ff",  x"03",  x"17",  x"d2",  x"3a",  x"93",  x"3d", -- 0A98
         x"3d",  x"00",  x"c9",  x"18",  x"1e",  x"1f",  x"5d",  x"00", -- 0AA0
         x"08",  x"09",  x"0f",  x"0a",  x"0b",  x"02",  x"0d",  x"b9", -- 0AA8
         x"92",  x"19",  x"de",  x"38",  x"5e",  x"0c",  x"62",  x"1b", -- 0AB0
         x"0c",  x"00",  x"9a",  x"90",  x"1c",  x"1d",  x"00",  x"7d", -- 0AB8
         x"ab",  x"8d",  x"82",  x"85",  x"86",  x"84",  x"cf",  x"00", -- 0AC0
         x"c3",  x"96",  x"90",  x"9b",  x"9c",  x"af",  x"c4",  x"95", -- 0AC8
         x"00",  x"92",  x"ae",  x"87",  x"ac",  x"8c",  x"91",  x"83", -- 0AD0
         x"ad",  x"09",  x"80",  x"81",  x"c2",  x"00",  x"00",  x"93", -- 0AD8
         x"02",  x"00",  x"ec",  x"ed",  x"ee",  x"ef",  x"f0",  x"ca", -- 0AE0
         x"cc",  x"00",  x"d0",  x"d1",  x"da",  x"de",  x"fc",  x"df", -- 0AE8
         x"fd",  x"db",  x"00",  x"b3",  x"a0",  x"a1",  x"9e",  x"9f", -- 0AF0
         x"c0",  x"c7",  x"b4",  x"2e",  x"b0",  x"b1",  x"c7",  x"00", -- 0AF8
         x"dc",  x"ff",  x"dd",  x"be",  x"b2",  x"a3",  x"f9",  x"aa", -- 0B00
         x"00",  x"a5",  x"a9",  x"88",  x"c8",  x"c6",  x"bc",  x"b6", -- 0B08
         x"bb",  x"00",  x"ba",  x"fb",  x"fa",  x"bd",  x"b8",  x"a8", -- 0B10
         x"c1",  x"a6",  x"00",  x"89",  x"b5",  x"f8",  x"a4",  x"a2", -- 0B18
         x"a7",  x"c5",  x"98",  x"00",  x"00",  x"d7",  x"b9",  x"d2", -- 0B20
         x"d3",  x"f2",  x"e0",  x"e2",  x"00",  x"f4",  x"e8",  x"f5", -- 0B28
         x"f6",  x"8a",  x"d4",  x"8b",  x"d8",  x"60",  x"d9",  x"e3", -- 0B30
         x"d5",  x"00",  x"d6",  x"ea",  x"e7",  x"f3",  x"e6",  x"c9", -- 0B38
         x"e1",  x"e9",  x"00",  x"e3",  x"e4",  x"cb",  x"94",  x"9d", -- 0B40
         x"97",  x"9a",  x"99",  x"cb",  x"b9",  x"97",  x"a1",  x"4e", -- 0B48
         x"53",  x"54",  x"8d",  x"16",  x"e0",  x"40",  x"52",  x"45", -- 0B50
         x"41",  x"44",  x"45",  x"32",  x"52",  x"00",  x"e6",  x"05", -- 0B58
         x"50",  x"55",  x"4e",  x"43",  x"48",  x"11",  x"ec",  x"91", -- 0B60
         x"4c",  x"49",  x"19",  x"95",  x"08",  x"9c",  x"c4",  x"4f", -- 0B68
         x"53",  x"03",  x"00",  x"c8",  x"d6",  x"c3",  x"ba",  x"05", -- 0B70
         x"f0",  x"41",  x"53",  x"47",  x"4e",  x"12",  x"14",  x"80", -- 0B78
         x"c3",  x"81",  x"f1",  x"54",  x"49",  x"39",  x"4d",  x"45", -- 0B80
         x"0b",  x"05",  x"22",  x"f5",  x"43",  x"4c",  x"4f",  x"3d", -- 0B88
         x"0b",  x"b3",  x"8e",  x"06",  x"43",  x"52",  x"54",  x"00", -- 0B90
         x"89",  x"04",  x"42",  x"41",  x"05",  x"14",  x"01",  x"01", -- 0B98
         x"0c",  x"72",  x"6f",  x"62",  x"6f",  x"74",  x"04",  x"22", -- 0BA0
         x"6e",  x"19",  x"5a",  x"20",  x"83",  x"c2",  x"30",  x"31", -- 0BA8
         x"47",  x"20",  x"14",  x"02",  x"50",  x"73",  x"74",  x"61", -- 0BB0
         x"72",  x"23",  x"74",  x"20",  x"04",  x"70",  x"65",  x"57", -- 0BB8
         x"08",  x"07",  x"42",  x"5e",  x"2d",  x"65",  x"40",  x"72", -- 0BC0
         x"24",  x"72",  x"07",  x"00",  x"6d",  x"65",  x"41",  x"6d", -- 0BC8
         x"06",  x"79",  x"20",  x"70",  x"72",  x"34",  x"17",  x"65", -- 0BD0
         x"63",  x"02",  x"96",  x"80",  x"65",  x"6e",  x"64",  x"20", -- 0BD8
         x"6f",  x"39",  x"66",  x"20",  x"17",  x"2a",  x"00",  x"72", -- 0BE0
         x"14",  x"06",  x"10",  x"20",  x"6e",  x"6f",  x"3c",  x"66", -- 0BE8
         x"6f",  x"75",  x"6e",  x"8b",  x"1e",  x"62",  x"61",  x"0d", -- 0BF0
         x"14",  x"90",  x"00",  x"66",  x"69",  x"6c",  x"79",  x"65", -- 0BF8
         x"19",  x"01",  x"20",  x"2c",  x"2e",  x"3a",  x"43",  x"ff", -- 0C00
         x"bf",  x"20",  x"fb",  x"fc",  x"c2",  x"05",  x"fc",  x"e4", -- 0C08
         x"fc",  x"bd",  x"ff",  x"f7",  x"2d",  x"f2",  x"0a",  x"fb", -- 0C10
         x"c4",  x"28",  x"f3",  x"8b",  x"a4",  x"9e",  x"40",  x"3e", -- 0C18
         x"3c",  x"2b",  x"34",  x"28",  x"be",  x"20",  x"96",  x"a0", -- 0C20
         x"ad",  x"f7",  x"3e",  x"6a",  x"18",  x"0a",  x"02",  x"0a", -- 0C28
         x"50",  x"f1",  x"be",  x"ed",  x"3e",  x"4d",  x"f5",  x"fd", -- 0C30
         x"34",  x"32",  x"23",  x"d9",  x"12",  x"7f",  x"32",  x"24", -- 0C38
         x"04",  x"a5",  x"e4",  x"79",  x"a2",  x"82",  x"16",  x"51", -- 0C40
         x"fb",  x"fe",  x"ad",  x"c8",  x"35",  x"eb",  x"bb",  x"a5", -- 0C48
         x"c3",  x"a6",  x"20",  x"82",  x"00",  x"cd",  x"30",  x"fd", -- 0C50
         x"28",  x"2e",  x"1c",  x"be",  x"ad",  x"1b",  x"2b",  x"36", -- 0C58
         x"28",  x"df",  x"17",  x"36",  x"06",  x"97",  x"42",  x"0e", -- 0C60
         x"0d",  x"23",  x"77",  x"fb",  x"f1",  x"fe",  x"cd",  x"82", -- 0C68
         x"04",  x"87",  x"c9",  x"07",  x"e1",  x"34",  x"ac",  x"7e", -- 0C70
         x"c9",  x"00",  x"e5",  x"d5",  x"c5",  x"21",  x"68",  x"fe", -- 0C78
         x"6a",  x"e5",  x"f5",  x"24",  x"7a",  x"0c",  x"7b",  x"02", -- 0C80
         x"3a",  x"62",  x"26",  x"9e",  x"00",  x"06",  x"cb",  x"c3", -- 0C88
         x"cb",  x"fa",  x"cb",  x"bd",  x"8b",  x"1b",  x"5a",  x"0e", -- 0C90
         x"fd",  x"80",  x"81",  x"fe",  x"67",  x"cd",  x"89",  x"fe", -- 0C98
         x"07",  x"6f",  x"d1",  x"c1",  x"c0",  x"c5",  x"cf",  x"40", -- 0CA0
         x"af",  x"cd",  x"83",  x"fe",  x"f5",  x"06",  x"84",  x"67", -- 0CA8
         x"f1",  x"85",  x"bf",  x"13",  x"d8",  x"12",  x"e0",  x"00", -- 0CB0
         x"5f",  x"7d",  x"fe",  x"48",  x"28",  x"6e",  x"fe",  x"44", -- 0CB8
         x"41",  x"34",  x"fe",  x"46",  x"af",  x"40",  x"3e",  x"a9", -- 0CC0
         x"d6",  x"2c",  x"6f",  x"00",  x"7c",  x"fe",  x"38",  x"c0", -- 0CC8
         x"7d",  x"c3",  x"38",  x"fe",  x"00",  x"fe",  x"40",  x"28", -- 0CD0
         x"6b",  x"d0",  x"d6",  x"39",  x"d8",  x"01",  x"84",  x"cb", -- 0CD8
         x"78",  x"28",  x"2d",  x"01",  x"90",  x"9b",  x"97",  x"d4", -- 0CE0
         x"ce",  x"61",  x"ae",  x"80",  x"60",  x"0d",  x"ed",  x"41", -- 0CE8
         x"cb",  x"7c",  x"00",  x"c8",  x"3c",  x"fe",  x"0c",  x"38", -- 0CF0
         x"64",  x"28",  x"60",  x"00",  x"fe",  x"0e",  x"38",  x"5e", -- 0CF8
         x"28",  x"5a",  x"fe",  x"0f",  x"00",  x"28",  x"58",  x"d6", -- 0D00
         x"2b",  x"38",  x"4e",  x"fe",  x"0d",  x"01",  x"d0",  x"21", -- 0D08
         x"33",  x"fb",  x"18",  x"55",  x"3d",  x"fe",  x"90",  x"d8", -- 0D10
         x"d6",  x"06",  x"04",  x"c8",  x"30",  x"0d",  x"fe",  x"fa", -- 0D18
         x"f8",  x"40",  x"d6",  x"1f",  x"cb",  x"73",  x"c8",  x"69", -- 0D20
         x"d6",  x"b3",  x"50",  x"00",  x"1b",  x"38",  x"34",  x"fe", -- 0D28
         x"1e",  x"c0",  x"18",  x"50",  x"2f",  x"60",  x"3b",  x"26", -- 0D30
         x"28",  x"26",  x"c1",  x"3b",  x"20",  x"28",  x"20",  x"37", -- 0D38
         x"82",  x"18",  x"21",  x"40",  x"34",  x"05",  x"20",  x"78", -- 0D40
         x"a9",  x"ba",  x"c0",  x"ef",  x"40",  x"a4",  x"7c",  x"20", -- 0D48
         x"c2",  x"b7",  x"00",  x"20",  x"a2",  x"3e",  x"5f",  x"18", -- 0D50
         x"08",  x"c6",  x"20",  x"0a",  x"c6",  x"2b",  x"c6",  x"10", -- 0D58
         x"05",  x"3e",  x"03",  x"28",  x"1d",  x"21",  x"53",  x"fb", -- 0D60
         x"06",  x"a9",  x"01",  x"09",  x"7e",  x"fe",  x"6d",  x"70", -- 0D68
         x"ee",  x"5d",  x"0d",  x"28",  x"ec",  x"b7",  x"e1",  x"d3", -- 0D70
         x"a5",  x"c4",  x"90",  x"0a",  x"18",  x"43",  x"e1",  x"22", -- 0D78
         x"fe",  x"7e",  x"ba",  x"d9",  x"96",  x"40",  x"aa",  x"a3", -- 0D80
         x"af",  x"11",  x"64",  x"b2",  x"14",  x"31",  x"fe",  x"7d", -- 0D88
         x"1e",  x"8a",  x"a7",  x"c5",  x"64",  x"04",  x"18",  x"15", -- 0D90
         x"ea",  x"c1",  x"d1",  x"21",  x"33",  x"e0",  x"10",  x"60", -- 0D98
         x"20",  x"03",  x"1d",  x"d6",  x"21",  x"3c",  x"e8",  x"96", -- 0DA0
         x"fa",  x"c9",  x"3e",  x"25",  x"ff",  x"2c",  x"ec",  x"34", -- 0DA8
         x"93",  x"e0",  x"af",  x"18",  x"d7",  x"00",  x"3e",  x"f7", -- 0DB0
         x"06",  x"08",  x"81",  x"cb",  x"3b",  x"d8",  x"05",  x"10", -- 0DB8
         x"fa",  x"c0",  x"81",  x"bf",  x"ab",  x"c1",  x"db",  x"91", -- 0DC0
         x"2f",  x"57",  x"9c",  x"79",  x"ef",  x"62",  x"fb",  x"2c", -- 0DC8
         x"86",  x"0b",  x"67",  x"3e",  x"fe",  x"06",  x"af",  x"6f", -- 0DD0
         x"90",  x"6f",  x"85",  x"25",  x"03",  x"cf",  x"85",  x"f0", -- 0DD8
         x"d3",  x"02",  x"91",  x"db",  x"90",  x"2f",  x"5f",  x"3e", -- 0DE0
         x"c1",  x"ed",  x"07",  x"dc",  x"92",  x"bc",  x"be",  x"e2", -- 0DE8
         x"09",  x"fe",  x"cb",  x"e4",  x"cc",  x"65",  x"a4",  x"46", -- 0DF0
         x"5f",  x"69",  x"0b",  x"0a",  x"5c",  x"fb",  x"2a",  x"ad", -- 0DF8
         x"9c",  x"aa",  x"c8",  x"e3",  x"fe",  x"cd",  x"08",  x"29", -- 0E00
         x"ff",  x"3a",  x"6b",  x"15",  x"18",  x"ff",  x"28",  x"2a", -- 0E08
         x"1b",  x"ad",  x"31",  x"80",  x"7e",  x"08",  x"3a",  x"24", -- 0E10
         x"33",  x"86",  x"28",  x"d4",  x"06",  x"f2",  x"0c",  x"28", -- 0E18
         x"7a",  x"b3",  x"31",  x"3e",  x"85",  x"8e",  x"10",  x"40", -- 0E20
         x"03",  x"fb",  x"57",  x"c9",  x"22",  x"c5",  x"4f",  x"96", -- 0E28
         x"08",  x"cb",  x"09",  x"f5",  x"dc",  x"3b",  x"f1",  x"d4", -- 0E30
         x"02",  x"2d",  x"ff",  x"10",  x"f4",  x"c1",  x"1e",  x"cd", -- 0E38
         x"41",  x"06",  x"1e",  x"20",  x"b6",  x"90",  x"1e",  x"40", -- 0E40
         x"7a",  x"23",  x"cd",  x"38",  x"2c",  x"32",  x"6a",  x"e2", -- 0E48
         x"2a",  x"02",  x"b5",  x"43",  x"fa",  x"53",  x"ef",  x"ac", -- 0E50
         x"cc",  x"5d",  x"3a",  x"ca",  x"10",  x"04",  x"79",  x"a9", -- 0E58
         x"05",  x"a8",  x"5c",  x"f3",  x"7e",  x"60",  x"e1",  x"3e", -- 0E60
         x"63",  x"05",  x"1c",  x"b0",  x"03",  x"18",  x"0f",  x"0b", -- 0E68
         x"0a",  x"c5",  x"03",  x"e7",  x"03",  x"d7",  x"20",  x"16", -- 0E70
         x"cd",  x"d1",  x"00",  x"ff",  x"38",  x"f9",  x"fe",  x"90", -- 0E78
         x"38",  x"f5",  x"10",  x"55",  x"f5",  x"b9",  x"ad",  x"1a", -- 0E80
         x"4f",  x"c0",  x"37",  x"cd",  x"e0",  x"ff",  x"fe",  x"00", -- 0E88
         x"52",  x"30",  x"f1",  x"10",  x"ef",  x"cd",  x"e8",  x"ff", -- 0E90
         x"11",  x"d8",  x"32",  x"6b",  x"a5",  x"91",  x"aa",  x"9a", -- 0E98
         x"0b",  x"77",  x"8f",  x"a9",  x"06",  x"f1",  x"0e",  x"b0", -- 0EA0
         x"47",  x"0e",  x"b8",  x"c8",  x"44",  x"37",  x"79",  x"db", -- 0EA8
         x"80",  x"7c",  x"07",  x"e5",  x"5f",  x"f1",  x"77",  x"d2", -- 0EB0
         x"af",  x"99",  x"3a",  x"e9",  x"b0",  x"4f",  x"0a",  x"e2", -- 0EB8
         x"81",  x"06",  x"c9",  x"16",  x"08",  x"af",  x"5f",  x"73", -- 0EC0
         x"08",  x"3f",  x"30",  x"04",  x"74",  x"d8",  x"37",  x"0a", -- 0EC8
         x"cb",  x"1b",  x"15",  x"20",  x"49",  x"0e",  x"3f",  x"7b", -- 0ED0
         x"c9",  x"00",  x"ff",  x"e0",  x"00",  x"18",  x"0b",  x"c3", -- 0ED8
         x"8c",  x"c0",  x"7f",  x"7f",  x"42",  x"00",  x"41",  x"53", -- 0EE0
         x"49",  x"43",  x"00",  x"21",  x"bd",  x"c0",  x"00",  x"11", -- 0EE8
         x"00",  x"03",  x"01",  x"67",  x"00",  x"ed",  x"b0",  x"00", -- 0EF0
         x"eb",  x"f9",  x"cd",  x"69",  x"c6",  x"32",  x"ab",  x"03", -- 0EF8
         x"00",  x"32",  x"00",  x"04",  x"21",  x"92",  x"c0",  x"cd", -- 0F00
         x"c9",  x"1a",  x"d1",  x"21",  x"ae",  x"05",  x"cd",  x"00", -- 0F08
         x"ae",  x"c5",  x"21",  x"62",  x"03",  x"cd",  x"86",  x"c9", -- 0F10
         x"08",  x"7a",  x"d6",  x"06",  x"21",  x"2a",  x"2b",  x"30", -- 0F18
         x"00",  x"03",  x"11",  x"ff",  x"bf",  x"23",  x"cd",  x"89", -- 0F20
         x"c6",  x"00",  x"28",  x"09",  x"7e",  x"47",  x"2f",  x"77", -- 0F28
         x"be",  x"70",  x"10",  x"28",  x"f2",  x"2b",  x"42",  x"ff", -- 0F30
         x"22",  x"b0",  x"08",  x"03",  x"19",  x"22",  x"56",  x"27", -- 0F38
         x"41",  x"c6",  x"20",  x"2a",  x"56",  x"21",  x"ef",  x"fb", -- 0F40
         x"19",  x"cd",  x"0d",  x"29",  x"d8",  x"21",  x"a0",  x"40", -- 0F48
         x"00",  x"2a",  x"04",  x"e0",  x"7e",  x"fe",  x"78",  x"20", -- 0F50
         x"01",  x"00",  x"3e",  x"af",  x"32",  x"fc",  x"03",  x"31", -- 0F58
         x"67",  x"03",  x"23",  x"18",  x"0a",  x"7c",  x"52",  x"45", -- 0F60
         x"7e",  x"9c",  x"71",  x"00",  x"c3",  x"88",  x"c3",  x"0c", -- 0F68
         x"0a",  x"0d",  x"48",  x"43",  x"71",  x"2d",  x"11",  x"09", -- 0F70
         x"00",  x"00",  x"20",  x"42",  x"59",  x"54",  x"45",  x"53", -- 0F78
         x"26",  x"20",  x"46",  x"23",  x"45",  x"0d",  x"00",  x"4d", -- 0F80
         x"45",  x"4d",  x"4f",  x"52",  x"59",  x"20",  x"00",  x"45", -- 0F88
         x"4e",  x"44",  x"20",  x"3f",  x"20",  x"3a",  x"00",  x"01", -- 0F90
         x"c3",  x"89",  x"c0",  x"c3",  x"67",  x"c9",  x"00",  x"00", -- 0F98
         x"a0",  x"d6",  x"00",  x"6f",  x"7c",  x"de",  x"10",  x"00", -- 0FA0
         x"67",  x"78",  x"03",  x"47",  x"3e",  x"00",  x"d0",  x"12", -- 0FA8
         x"35",  x"4a",  x"ca",  x"99",  x"00",  x"39",  x"1c",  x"76", -- 0FB0
         x"98",  x"22",  x"95",  x"b3",  x"98",  x"00",  x"0a",  x"dd", -- 0FB8
         x"47",  x"98",  x"53",  x"d1",  x"99",  x"99",  x"00",  x"0a", -- 0FC0
         x"1a",  x"9f",  x"98",  x"65",  x"bc",  x"cd",  x"98",  x"00", -- 0FC8
         x"d6",  x"77",  x"3e",  x"98",  x"52",  x"c7",  x"4f",  x"80", -- 0FD0
         x"06",  x"0b",  x"ff",  x"1b",  x"00",  x"0a",  x"01",  x"28", -- 0FD8
         x"00",  x"49",  x"d7",  x"9d",  x"00",  x"00",  x"83",  x"65", -- 0FE0
         x"04",  x"fe",  x"ff",  x"00",  x"43",  x"4c",  x"01",  x"04", -- 0FE8
         x"0d",  x"48",  x"c5",  x"6b",  x"c6",  x"73",  x"ce",  x"45", -- 0FF0
         x"00",  x"58",  x"54",  x"c4",  x"41",  x"54",  x"41",  x"c9", -- 0FF8
         x"4e",  x"20",  x"50",  x"55",  x"08",  x"49",  x"4d",  x"d2", -- 1000
         x"45",  x"04",  x"41",  x"44",  x"cc",  x"45",  x"54",  x"43", -- 1008
         x"54",  x"02",  x"4f",  x"d2",  x"55",  x"4e",  x"c9",  x"46", -- 1010
         x"0f",  x"51",  x"53",  x"09",  x"a3",  x"41",  x"0f",  x"53", -- 1018
         x"55",  x"42",  x"d2",  x"17",  x"08",  x"55",  x"52",  x"4e", -- 1020
         x"05",  x"4d",  x"d3",  x"88",  x"12",  x"50",  x"cf",  x"2e", -- 1028
         x"cf",  x"4e",  x"01",  x"ce",  x"55",  x"4c",  x"4c",  x"d7", -- 1030
         x"41",  x"49",  x"38",  x"00",  x"45",  x"46",  x"d0",  x"4f", -- 1038
         x"4b",  x"45",  x"c4",  x"c2",  x"03",  x"c1",  x"55",  x"1c", -- 1040
         x"10",  x"cc",  x"49",  x"4e",  x"36",  x"c3",  x"4c",  x"53", -- 1048
         x"00",  x"d7",  x"49",  x"44",  x"54",  x"48",  x"c2",  x"59", -- 1050
         x"45",  x"11",  x"a1",  x"c3",  x"41",  x"27",  x"d0",  x"52", -- 1058
         x"15",  x"0a",  x"54",  x"c3",  x"4f",  x"03",  x"1d",  x"a9", -- 1060
         x"52",  x"1c",  x"67",  x"52",  x"04",  x"20",  x"4f",  x"6c", -- 1068
         x"c3",  x"53",  x"41",  x"56",  x"44",  x"45",  x"85",  x"57", -- 1070
         x"00",  x"d4",  x"41",  x"42",  x"28",  x"d4",  x"4f",  x"c6", -- 1078
         x"4e",  x"11",  x"d3",  x"50",  x"43",  x"07",  x"48",  x"45", -- 1080
         x"5a",  x"45",  x"81",  x"66",  x"00",  x"45",  x"50",  x"ab", -- 1088
         x"ad",  x"aa",  x"af",  x"de",  x"44",  x"c1",  x"aa",  x"cf", -- 1090
         x"02",  x"52",  x"be",  x"bd",  x"bc",  x"d3",  x"47",  x"91", -- 1098
         x"28",  x"3f",  x"c1",  x"42",  x"04",  x"53",  x"d5",  x"53", -- 10A0
         x"52",  x"c6",  x"94",  x"51",  x"b3",  x"90",  x"75",  x"53", -- 10A8
         x"d3",  x"51",  x"20",  x"52",  x"d2",  x"1f",  x"cc",  x"4e", -- 10B0
         x"c5",  x"58",  x"55",  x"50",  x"5d",  x"0d",  x"64",  x"49", -- 10B8
         x"02",  x"4e",  x"c1",  x"54",  x"4e",  x"d0",  x"d7",  x"44", -- 10C0
         x"4b",  x"96",  x"50",  x"03",  x"d0",  x"49",  x"cc",  x"a1", -- 10C8
         x"4c",  x"49",  x"52",  x"24",  x"d6",  x"83",  x"10",  x"c1", -- 10D0
         x"53",  x"43",  x"28",  x"c3",  x"48",  x"09",  x"10",  x"46", -- 10D8
         x"54",  x"04",  x"24",  x"d2",  x"49",  x"47",  x"48",  x"05", -- 10E0
         x"cd",  x"8a",  x"a1",  x"0e",  x"8c",  x"85",  x"22",  x"d4", -- 10E8
         x"52",  x"98",  x"c0",  x"03",  x"46",  x"46",  x"c5",  x"44", -- 10F0
         x"89",  x"cd",  x"c5",  x"b9",  x"10",  x"45",  x"80",  x"1a", -- 10F8
         x"00",  x"c9",  x"de",  x"c7",  x"dc",  x"cc",  x"48",  x"ca", -- 1100
         x"ec",  x"00",  x"cb",  x"01",  x"cf",  x"1f",  x"cc",  x"5d", -- 1108
         x"ca",  x"07",  x"00",  x"ca",  x"eb",  x"c9",  x"cf",  x"ca", -- 1110
         x"df",  x"c8",  x"f6",  x"13",  x"c9",  x"25",  x"ca",  x"81", -- 1118
         x"00",  x"18",  x"c9",  x"ec",  x"d3",  x"b3",  x"ca",  x"c0", -- 1120
         x"01",  x"cb",  x"f7",  x"d3",  x"c4",  x"d0",  x"37",  x"d4", -- 1128
         x"3a",  x"00",  x"fa",  x"c5",  x"ea",  x"c6",  x"d0",  x"dd", -- 1130
         x"b9",  x"10",  x"cb",  x"f4",  x"df",  x"1b",  x"38",  x"db", -- 1138
         x"fa",  x"00",  x"ca",  x"48",  x"c9",  x"f2",  x"c6",  x"aa", -- 1140
         x"c9",  x"43",  x"00",  x"dc",  x"41",  x"dd",  x"40",  x"c6", -- 1148
         x"2d",  x"c6",  x"b7",  x"04",  x"c7",  x"b8",  x"c7",  x"e7", -- 1150
         x"c3",  x"19",  x"a6",  x"00",  x"d6",  x"70",  x"d7",  x"bc", -- 1158
         x"d6",  x"03",  x"03",  x"90",  x"00",  x"d0",  x"e3",  x"d3", -- 1160
         x"bd",  x"d0",  x"1f",  x"d9",  x"fd",  x"00",  x"d9",  x"59", -- 1168
         x"d5",  x"6d",  x"d9",  x"70",  x"da",  x"76",  x"01",  x"da", -- 1170
         x"d7",  x"da",  x"ec",  x"da",  x"31",  x"d4",  x"86",  x"10", -- 1178
         x"d5",  x"d6",  x"2c",  x"00",  x"d3",  x"56",  x"d1",  x"bf", -- 1180
         x"d3",  x"3b",  x"d3",  x"4b",  x"00",  x"d3",  x"5b",  x"d3", -- 1188
         x"89",  x"d3",  x"92",  x"d3",  x"79",  x"00",  x"11",  x"d8", -- 1190
         x"79",  x"6a",  x"d4",  x"7c",  x"98",  x"d5",  x"00",  x"7c", -- 1198
         x"f3",  x"d5",  x"7f",  x"28",  x"d9",  x"50",  x"5e",  x"00", -- 11A0
         x"ce",  x"46",  x"5d",  x"ce",  x"4e",  x"46",  x"53",  x"4e", -- 11A8
         x"00",  x"52",  x"47",  x"4f",  x"44",  x"46",  x"43",  x"4f", -- 11B0
         x"56",  x"26",  x"4f",  x"4d",  x"84",  x"90",  x"91",  x"44", -- 11B8
         x"44",  x"25",  x"2f",  x"30",  x"ed",  x"28",  x"c5",  x"45", -- 11C0
         x"53",  x"bc",  x"de",  x"20",  x"43",  x"4e",  x"55",  x"45", -- 11C8
         x"46",  x"0a",  x"49",  x"4f",  x"d0",  x"04",  x"52",  x"52", -- 11D0
         x"bd",  x"ca",  x"07",  x"ec",  x"24",  x"95",  x"09",  x"20", -- 11D8
         x"00",  x"46",  x"49",  x"f4",  x"28",  x"ef",  x"24",  x"4f", -- 11E0
         x"55",  x"ac",  x"4d",  x"0d",  x"a7",  x"f2",  x"41",  x"42", -- 11E8
         x"52",  x"82",  x"30",  x"4b",  x"00",  x"e5",  x"00",  x"2a", -- 11F0
         x"db",  x"03",  x"06",  x"00",  x"09",  x"09",  x"3e",  x"00", -- 11F8
         x"e5",  x"3e",  x"d0",  x"95",  x"6f",  x"3e",  x"ff",  x"9c", -- 1200
         x"00",  x"38",  x"04",  x"67",  x"39",  x"e1",  x"d8",  x"1e", -- 1208
         x"0c",  x"00",  x"18",  x"14",  x"2a",  x"ca",  x"03",  x"22", -- 1210
         x"58",  x"03",  x"04",  x"1e",  x"02",  x"01",  x"1e",  x"14", -- 1218
         x"02",  x"00",  x"92",  x"02",  x"12",  x"02",  x"22",  x"bb", -- 1220
         x"d5",  x"43",  x"fe",  x"50",  x"55",  x"cb",  x"21",  x"00", -- 1228
         x"dd",  x"c2",  x"57",  x"19",  x"44",  x"4d",  x"0b",  x"3e", -- 1230
         x"25",  x"3f",  x"1e",  x"0e",  x"d6",  x"c4",  x"85",  x"05", -- 1238
         x"c3",  x"83",  x"ac",  x"2e",  x"11",  x"a2",  x"e2",  x"b4", -- 1240
         x"d0",  x"ca",  x"0d",  x"00",  x"c0",  x"7c",  x"a5",  x"3c", -- 1248
         x"c4",  x"21",  x"d8",  x"3e",  x"3a",  x"c1",  x"af",  x"2f", -- 1250
         x"68",  x"1d",  x"20",  x"37",  x"dc",  x"fd",  x"06",  x"dd", -- 1258
         x"cd",  x"df",  x"c6",  x"2b",  x"57",  x"00",  x"21",  x"ea", -- 1260
         x"03",  x"3a",  x"4d",  x"03",  x"b7",  x"00",  x"28",  x"6b", -- 1268
         x"ed",  x"5b",  x"4e",  x"03",  x"f2",  x"f0",  x"02",  x"c3", -- 1270
         x"d5",  x"cd",  x"2a",  x"d8",  x"d1",  x"04",  x"00",  x"bb", -- 1278
         x"c4",  x"3e",  x"2a",  x"38",  x"02",  x"3e",  x"20",  x"b9", -- 1280
         x"8f",  x"c6",  x"92",  x"78",  x"d1",  x"28",  x"30",  x"06", -- 1288
         x"3f",  x"25",  x"18",  x"ba",  x"2c",  x"2a",  x"50",  x"f7", -- 1290
         x"06",  x"38",  x"f4",  x"d5",  x"11",  x"f9",  x"5d",  x"c5", -- 1298
         x"15",  x"ea",  x"22",  x"33",  x"ae",  x"78",  x"f5",  x"05", -- 12A0
         x"18",  x"47",  x"c8",  x"cd",  x"97",  x"28",  x"b5",  x"71", -- 12A8
         x"c0",  x"c1",  x"39",  x"80",  x"30",  x"58",  x"d5",  x"7e", -- 12B0
         x"23",  x"13",  x"b6",  x"23",  x"28",  x"3e",  x"7f",  x"34", -- 12B8
         x"23",  x"0a",  x"66",  x"6f",  x"26",  x"2c",  x"94",  x"00", -- 12C0
         x"de",  x"d1",  x"c2",  x"96",  x"c3",  x"38",  x"b7",  x"3f", -- 12C8
         x"0e",  x"18",  x"cd",  x"3e",  x"3e",  x"56",  x"51",  x"da", -- 12D0
         x"0f",  x"21",  x"61",  x"19",  x"02",  x"bd",  x"c8",  x"3c", -- 12D8
         x"3d",  x"ca",  x"0a",  x"64",  x"f5",  x"3f",  x"78",  x"da", -- 12E0
         x"00",  x"c4",  x"47",  x"d1",  x"f1",  x"d2",  x"8a",  x"c8", -- 12E8
         x"d5",  x"4d",  x"c5",  x"71",  x"cd",  x"1b",  x"50",  x"b7", -- 12F0
         x"17",  x"52",  x"38",  x"08",  x"f1",  x"00",  x"f5",  x"b7", -- 12F8
         x"20",  x"03",  x"c3",  x"20",  x"ca",  x"c5",  x"00",  x"30", -- 1300
         x"11",  x"eb",  x"2a",  x"d7",  x"03",  x"1a",  x"02",  x"23", -- 1308
         x"03",  x"13",  x"82",  x"02",  x"20",  x"f7",  x"ed",  x"43", -- 1310
         x"0c",  x"8c",  x"30",  x"28",  x"22",  x"13",  x"00",  x"e3", -- 1318
         x"c1",  x"09",  x"e5",  x"cd",  x"ab",  x"c4",  x"e1",  x"40", -- 1320
         x"22",  x"0a",  x"eb",  x"36",  x"ff",  x"d1",  x"23",  x"01", -- 1328
         x"23",  x"73",  x"23",  x"72",  x"23",  x"11",  x"62",  x"2b", -- 1330
         x"0b",  x"77",  x"23",  x"13",  x"3c",  x"ef",  x"0a",  x"d5", -- 1338
         x"84",  x"23",  x"eb",  x"21",  x"67",  x"e5",  x"23",  x"62", -- 1340
         x"6b",  x"9e",  x"08",  x"c8",  x"23",  x"04",  x"a6",  x"3c", -- 1348
         x"80",  x"05",  x"af",  x"be",  x"23",  x"20",  x"fc",  x"eb", -- 1350
         x"c0",  x"29",  x"18",  x"e8",  x"cd",  x"30",  x"2c",  x"c3", -- 1358
         x"c5",  x"43",  x"55",  x"00",  x"7e",  x"02",  x"c8",  x"0b", -- 1360
         x"2b",  x"18",  x"f6",  x"2a",  x"24",  x"5f",  x"03",  x"d9", -- 1368
         x"c2",  x"2a",  x"2b",  x"c8",  x"4a",  x"8d",  x"c5",  x"c3", -- 1370
         x"19",  x"60",  x"69",  x"08",  x"40",  x"3f",  x"c8",  x"3f", -- 1378
         x"d0",  x"18",  x"e4",  x"88",  x"9f",  x"af",  x"03",  x"32", -- 1380
         x"0e",  x"05",  x"5f",  x"08",  x"44",  x"fb",  x"e5",  x"fe", -- 1388
         x"88",  x"9a",  x"71",  x"c5",  x"00",  x"47",  x"fe",  x"22", -- 1390
         x"ca",  x"91",  x"c5",  x"b7",  x"ca",  x"10",  x"97",  x"c5", -- 1398
         x"3a",  x"1b",  x"b7",  x"7e",  x"20",  x"01",  x"73",  x"fe", -- 13A0
         x"3f",  x"3e",  x"9e",  x"28",  x"6d",  x"1c",  x"17",  x"30", -- 13A8
         x"38",  x"f3",  x"09",  x"3c",  x"38",  x"64",  x"b8",  x"00", -- 13B0
         x"20",  x"c1",  x"c5",  x"01",  x"6d",  x"c5",  x"10",  x"c5", -- 13B8
         x"06",  x"7f",  x"13",  x"61",  x"38",  x"07",  x"32",  x"fe", -- 13C0
         x"7b",  x"df",  x"04",  x"e6",  x"5f",  x"77",  x"4e",  x"eb", -- 13C8
         x"64",  x"f2",  x"00",  x"26",  x"c5",  x"04",  x"7e",  x"e6", -- 13D0
         x"7f",  x"20",  x"15",  x"64",  x"3a",  x"b6",  x"a7",  x"11", -- 13D8
         x"c8",  x"3a",  x"fb",  x"04",  x"c0",  x"3c",  x"57",  x"83", -- 13E0
         x"2a",  x"0c",  x"e0",  x"15",  x"00",  x"c8",  x"b9",  x"20", -- 13E8
         x"dd",  x"eb",  x"e5",  x"00",  x"13",  x"1a",  x"b7",  x"fa", -- 13F0
         x"69",  x"c5",  x"4f",  x"78",  x"09",  x"fe",  x"88",  x"20", -- 13F8
         x"04",  x"98",  x"43",  x"2b",  x"23",  x"43",  x"50",  x"02", -- 1400
         x"3f",  x"b9",  x"28",  x"e5",  x"05",  x"e1",  x"18",  x"bb", -- 1408
         x"48",  x"f1",  x"98",  x"82",  x"eb",  x"79",  x"c1",  x"f6", -- 1410
         x"20",  x"12",  x"13",  x"0c",  x"d6",  x"24",  x"3a",  x"28", -- 1418
         x"6f",  x"49",  x"af",  x"91",  x"a1",  x"80",  x"d6",  x"54", -- 1420
         x"28",  x"05",  x"d6",  x"12",  x"0e",  x"c2",  x"e3",  x"d6", -- 1428
         x"1a",  x"7e",  x"b7",  x"c3",  x"08",  x"b8",  x"28",  x"e0", -- 1430
         x"1f",  x"0c",  x"13",  x"25",  x"18",  x"f3",  x"f7",  x"2c", -- 1438
         x"27",  x"01",  x"31",  x"c9",  x"4c",  x"85",  x"0a",  x"00", -- 1440
         x"52",  x"8c",  x"8c",  x"00",  x"43",  x"92",  x"4a",  x"86", -- 1448
         x"a7",  x"cd",  x"00",  x"e3",  x"cd",  x"e4",  x"dd",  x"e3", -- 1450
         x"fe",  x"00",  x"1c",  x"11",  x"9f",  x"c5",  x"28",  x"0e", -- 1458
         x"fe",  x"1d",  x"28",  x"11",  x"a4",  x"06",  x"a7",  x"80", -- 1460
         x"1e",  x"11",  x"a8",  x"c5",  x"20",  x"14",  x"c9",  x"34", -- 1468
         x"c9",  x"24",  x"cd",  x"49",  x"a7",  x"cb",  x"a3",  x"ba", -- 1470
         x"f1",  x"00",  x"c5",  x"e1",  x"c3",  x"5e",  x"cb",  x"cd", -- 1478
         x"0f",  x"df",  x"00",  x"20",  x"02",  x"e1",  x"c9",  x"cd", -- 1480
         x"27",  x"df",  x"38",  x"90",  x"e1",  x"32",  x"df",  x"2a", -- 1488
         x"18",  x"c1",  x"66",  x"8b",  x"00",  x"d5",  x"dd",  x"23", -- 1490
         x"18",  x"f7",  x"11",  x"c8",  x"f7",  x"d5",  x"28",  x"4e", -- 1498
         x"17",  x"d4",  x"09",  x"eb",  x"e3",  x"28",  x"b3",  x"aa", -- 14A0
         x"9c",  x"51",  x"c8",  x"e1",  x"bd",  x"41",  x"28",  x"06", -- 14A8
         x"10",  x"80",  x"c2",  x"48",  x"c3",  x"eb",  x"7d",  x"34", -- 14B0
         x"b4",  x"ca",  x"d9",  x"45",  x"22",  x"10",  x"cb",  x"ff", -- 14B8
         x"a3",  x"22",  x"e1",  x"a0",  x"90",  x"c1",  x"c3",  x"54", -- 14C0
         x"96",  x"9a",  x"5f",  x"12",  x"de",  x"3a",  x"09",  x"91", -- 14C8
         x"45",  x"25",  x"f3",  x"3e",  x"89",  x"00",  x"b2",  x"dc", -- 14D0
         x"f1",  x"af",  x"18",  x"27",  x"ea",  x"c0",  x"85",  x"24", -- 14D8
         x"e0",  x"26",  x"5e",  x"03",  x"c3",  x"a7",  x"01",  x"d8", -- 14E0
         x"32",  x"0d",  x"b5",  x"a4",  x"cf",  x"06",  x"b0",  x"b1", -- 14E8
         x"93",  x"c4",  x"17",  x"30",  x"cd",  x"87",  x"9c",  x"f7", -- 14F0
         x"25",  x"22",  x"d9",  x"02",  x"db",  x"3f",  x"89",  x"c9", -- 14F8
         x"97",  x"12",  x"b4",  x"0a",  x"44",  x"b2",  x"9a",  x"1d", -- 1500
         x"02",  x"de",  x"af",  x"6f",  x"67",  x"22",  x"d5",  x"ff", -- 1508
         x"24",  x"cc",  x"0e",  x"df",  x"08",  x"03",  x"e5",  x"c5", -- 1510
         x"2a",  x"31",  x"c9",  x"7c",  x"e0",  x"e5",  x"7d",  x"93", -- 1518
         x"48",  x"c9",  x"b2",  x"41",  x"02",  x"d8",  x"fe",  x"5b", -- 1520
         x"3f",  x"c9",  x"3a",  x"51",  x"93",  x"e5",  x"8f",  x"95", -- 1528
         x"6e",  x"74",  x"4c",  x"d6",  x"3e",  x"2b",  x"08",  x"18", -- 1530
         x"eb",  x"11",  x"c3",  x"b6",  x"24",  x"f5",  x"de",  x"98", -- 1538
         x"c8",  x"38",  x"13",  x"00",  x"3a",  x"41",  x"03",  x"47", -- 1540
         x"3a",  x"ac",  x"03",  x"04",  x"90",  x"ba",  x"05",  x"b8", -- 1548
         x"13",  x"cc",  x"61",  x"cb",  x"88",  x"48",  x"0b",  x"79", -- 1550
         x"d4",  x"c1",  x"c1",  x"f1",  x"c9",  x"e7",  x"65",  x"ba", -- 1558
         x"61",  x"3e",  x"09",  x"bf",  x"5b",  x"bf",  x"66",  x"ca", -- 1560
         x"15",  x"fd",  x"5c",  x"d3",  x"22",  x"42",  x"61",  x"64", -- 1568
         x"63",  x"03",  x"65",  x"82",  x"40",  x"6c",  x"c9",  x"ed", -- 1570
         x"53",  x"56",  x"46",  x"68",  x"89",  x"a0",  x"25",  x"de", -- 1578
         x"cd",  x"c8",  x"dd",  x"23",  x"28",  x"12",  x"c5",  x"85", -- 1580
         x"2a",  x"13",  x"a6",  x"6a",  x"ff",  x"ea",  x"b4",  x"08", -- 1588
         x"5b",  x"e1",  x"a3",  x"60",  x"c5",  x"cd",  x"91",  x"c7", -- 1590
         x"e1",  x"00",  x"4e",  x"23",  x"46",  x"23",  x"78",  x"b1", -- 1598
         x"28",  x"59",  x"00",  x"cd",  x"67",  x"c7",  x"cd",  x"f9", -- 15A0
         x"c8",  x"c5",  x"5e",  x"13",  x"23",  x"56",  x"23",  x"80", -- 15A8
         x"22",  x"ea",  x"be",  x"af",  x"71",  x"84",  x"22",  x"8f", -- 15B0
         x"aa",  x"2c",  x"65",  x"ee",  x"28",  x"d2",  x"26",  x"28", -- 15B8
         x"14",  x"b9",  x"12",  x"d3",  x"f2",  x"3c",  x"23",  x"9a", -- 15C0
         x"02",  x"95",  x"11",  x"1a",  x"cb",  x"03",  x"f2",  x"4e", -- 15C8
         x"c7",  x"18",  x"e6",  x"1c",  x"89",  x"18",  x"ba",  x"1f", -- 15D0
         x"83",  x"d7",  x"18",  x"f2",  x"bf",  x"02",  x"44",  x"03", -- 15D8
         x"d2",  x"49",  x"9a",  x"13",  x"44",  x"62",  x"c0",  x"5a", -- 15E0
         x"27",  x"c2",  x"02",  x"fe",  x"03",  x"20",  x"ea",  x"84", -- 15E8
         x"35",  x"0c",  x"4e",  x"b7",  x"ee",  x"22",  x"2a",  x"82", -- 15F0
         x"cf",  x"7f",  x"8b",  x"ca",  x"29",  x"8f",  x"33",  x"26", -- 15F8
         x"01",  x"c9",  x"d6",  x"7f",  x"fe",  x"56",  x"d7",  x"61", -- 1600
         x"d6",  x"55",  x"96",  x"35",  x"e3",  x"0c",  x"18",  x"b0", -- 1608
         x"06",  x"21",  x"c1",  x"47",  x"5a",  x"85",  x"ac",  x"c7", -- 1610
         x"10",  x"f8",  x"f0",  x"11",  x"e7",  x"48",  x"f3",  x"0a", -- 1618
         x"89",  x"ca",  x"21",  x"a0",  x"d2",  x"39",  x"81",  x"30", -- 1620
         x"81",  x"c0",  x"8d",  x"a9",  x"02",  x"e5",  x"69",  x"60", -- 1628
         x"7a",  x"b3",  x"eb",  x"d8",  x"84",  x"eb",  x"b0",  x"a3", -- 1630
         x"01",  x"b7",  x"20",  x"e1",  x"c8",  x"09",  x"18",  x"12", -- 1638
         x"e3",  x"3e",  x"64",  x"e2",  x"8d",  x"cd",  x"95",  x"96", -- 1640
         x"c1",  x"f8",  x"6c",  x"a2",  x"22",  x"44",  x"c8",  x"e5", -- 1648
         x"02",  x"82",  x"30",  x"cd",  x"c1",  x"c7",  x"d1",  x"ab", -- 1650
         x"80",  x"09",  x"d5",  x"2b",  x"56",  x"2c",  x"2b",  x"5e", -- 1658
         x"b8",  x"ac",  x"6e",  x"15",  x"30",  x"00",  x"e1",  x"20", -- 1660
         x"e8",  x"d1",  x"f9",  x"eb",  x"0e",  x"08",  x"a2",  x"a7", -- 1668
         x"ff",  x"cc",  x"11",  x"4a",  x"e3",  x"04",  x"58",  x"e8", -- 1670
         x"40",  x"29",  x"cd",  x"cd",  x"cc",  x"04",  x"c8",  x"a6", -- 1678
         x"cd",  x"26",  x"cd",  x"3e",  x"eb",  x"00",  x"d6",  x"e1", -- 1680
         x"c5",  x"d5",  x"01",  x"00",  x"81",  x"51",  x"4c",  x"5a", -- 1688
         x"a2",  x"ab",  x"0a",  x"3e",  x"01",  x"20",  x"0e",  x"e1", -- 1690
         x"ce",  x"18",  x"a4",  x"d0",  x"d2",  x"1b",  x"f5",  x"33", -- 1698
         x"33",  x"40",  x"cf",  x"33",  x"06",  x"81",  x"c5",  x"33", -- 16A0
         x"cd",  x"25",  x"16",  x"de",  x"af",  x"29",  x"86",  x"2a", -- 16A8
         x"2a",  x"e8",  x"8a",  x"28",  x"b7",  x"ce",  x"45",  x"23", -- 16B0
         x"a6",  x"e4",  x"7f",  x"c9",  x"4a",  x"23",  x"c2",  x"4d", -- 16B8
         x"83",  x"59",  x"22",  x"3a",  x"bb",  x"91",  x"99",  x"0f", -- 16C0
         x"ca",  x"a2",  x"3c",  x"a7",  x"76",  x"ca",  x"53",  x"ef", -- 16C8
         x"16",  x"cd",  x"48",  x"50",  x"11",  x"54",  x"c0",  x"d7", -- 16D0
         x"c8",  x"d6",  x"22",  x"80",  x"da",  x"b0",  x"00",  x"fe", -- 16D8
         x"25",  x"38",  x"14",  x"d6",  x"50",  x"38",  x"34",  x"05", -- 16E0
         x"fe",  x"05",  x"38",  x"0a",  x"47",  x"f2",  x"a8",  x"28", -- 16E8
         x"29",  x"c3",  x"03",  x"03",  x"e0",  x"c6",  x"25",  x"07", -- 16F0
         x"4f",  x"85",  x"6c",  x"a4",  x"04",  x"40",  x"c2",  x"09", -- 16F8
         x"f1",  x"62",  x"c5",  x"96",  x"ec",  x"60",  x"50",  x"d0", -- 1700
         x"90",  x"28",  x"5c",  x"f7",  x"c0",  x"3f",  x"ca",  x"a3", -- 1708
         x"bc",  x"86",  x"e3",  x"ac",  x"15",  x"cb",  x"10",  x"ea", -- 1710
         x"c3",  x"6f",  x"3e",  x"2c",  x"be",  x"c0",  x"9f",  x"3e", -- 1718
         x"29",  x"45",  x"18",  x"d2",  x"90",  x"59",  x"a6",  x"62", -- 1720
         x"eb",  x"d6",  x"71",  x"e5",  x"d5",  x"39",  x"9e",  x"81", -- 1728
         x"d1",  x"d2",  x"87",  x"84",  x"85",  x"cc",  x"dd",  x"80", -- 1730
         x"a8",  x"86",  x"01",  x"f3",  x"dd",  x"c0",  x"fe",  x"13", -- 1738
         x"28",  x"08",  x"87",  x"32",  x"c0",  x"8d",  x"70",  x"18", -- 1740
         x"0f",  x"9d",  x"92",  x"0a",  x"1e",  x"c8",  x"fe",  x"0a", -- 1748
         x"02",  x"30",  x"02",  x"02",  x"18",  x"f1",  x"c0",  x"f6", -- 1750
         x"c0",  x"c0",  x"30",  x"21",  x"f6",  x"25",  x"ff",  x"c1", -- 1758
         x"89",  x"02",  x"f5",  x"7d",  x"a4",  x"3c",  x"9c",  x"e2", -- 1760
         x"22",  x"d3",  x"d7",  x"aa",  x"12",  x"b6",  x"b3",  x"ab", -- 1768
         x"78",  x"ab",  x"c3",  x"ae",  x"70",  x"f1",  x"21",  x"00", -- 1770
         x"21",  x"c3",  x"c2",  x"71",  x"c3",  x"c3",  x"88",  x"c3", -- 1778
         x"42",  x"2a",  x"16",  x"7c",  x"b5",  x"1e",  x"5c",  x"27", -- 1780
         x"56",  x"c3",  x"72",  x"d3",  x"90",  x"2e",  x"61",  x"4b", -- 1788
         x"a1",  x"12",  x"9d",  x"80",  x"f2",  x"6f",  x"c9",  x"1e", -- 1790
         x"08",  x"58",  x"c3",  x"19",  x"0d",  x"3a",  x"00",  x"e8", -- 1798
         x"03",  x"fe",  x"90",  x"da",  x"45",  x"d7",  x"01",  x"04", -- 17A0
         x"80",  x"90",  x"11",  x"00",  x"00",  x"93",  x"40",  x"18", -- 17A8
         x"d7",  x"e1",  x"51",  x"c8",  x"19",  x"18",  x"e1",  x"2b", -- 17B0
         x"0c",  x"2e",  x"80",  x"d0",  x"e5",  x"f5",  x"21",  x"98", -- 17B8
         x"4e",  x"19",  x"8e",  x"22",  x"da",  x"c2",  x"d0",  x"85", -- 17C0
         x"19",  x"29",  x"80",  x"01",  x"f1",  x"d6",  x"30",  x"5f", -- 17C8
         x"16",  x"00",  x"30",  x"19",  x"eb",  x"c0",  x"24",  x"e0", -- 17D0
         x"28",  x"ad",  x"44",  x"5e",  x"53",  x"be",  x"c8",  x"e6", -- 17D8
         x"88",  x"b0",  x"a1",  x"8b",  x"10",  x"e1",  x"b0",  x"ca", -- 17E0
         x"bd",  x"9b",  x"6c",  x"10",  x"df",  x"28",  x"e3",  x"58", -- 17E8
         x"eb",  x"bb",  x"5f",  x"04",  x"7c",  x"9a",  x"57",  x"da", -- 17F0
         x"3e",  x"be",  x"e5",  x"f1",  x"87",  x"01",  x"28",  x"aa", -- 17F8
         x"58",  x"45",  x"d2",  x"85",  x"0d",  x"eb",  x"22",  x"56", -- 1800
         x"bd",  x"e5",  x"30",  x"8a",  x"83",  x"53",  x"ed",  x"84", -- 1808
         x"4f",  x"ec",  x"91",  x"05",  x"01",  x"54",  x"6f",  x"09", -- 1810
         x"10",  x"0e",  x"03",  x"e8",  x"ca",  x"94",  x"27",  x"e5", -- 1818
         x"82",  x"3e",  x"8c",  x"ba",  x"6a",  x"ee",  x"97",  x"86", -- 1820
         x"49",  x"f8",  x"9b",  x"0f",  x"8c",  x"4a",  x"23",  x"09", -- 1828
         x"dc",  x"be",  x"c4",  x"d4",  x"ae",  x"57",  x"2b",  x"e1", -- 1830
         x"48",  x"0e",  x"b8",  x"c1",  x"c0",  x"16",  x"ff",  x"9d", -- 1838
         x"10",  x"c7",  x"f9",  x"fe",  x"05",  x"8c",  x"1e",  x"04", -- 1840
         x"20",  x"f0",  x"4e",  x"24",  x"22",  x"23",  x"eb",  x"1b", -- 1848
         x"20",  x"07",  x"3a",  x"ff",  x"4c",  x"db",  x"87",  x"e2", -- 1850
         x"a2",  x"50",  x"81",  x"43",  x"e1",  x"01",  x"3a",  x"0e", -- 1858
         x"00",  x"9a",  x"30",  x"79",  x"48",  x"47",  x"c4",  x"df", -- 1860
         x"2d",  x"b8",  x"c8",  x"95",  x"40",  x"f3",  x"18",  x"f4", -- 1868
         x"cd",  x"06",  x"cf",  x"a4",  x"c0",  x"09",  x"b4",  x"d5", -- 1870
         x"3a",  x"ae",  x"c2",  x"22",  x"fa",  x"c9",  x"91",  x"e3", -- 1878
         x"d2",  x"28",  x"1f",  x"04",  x"cd",  x"2b",  x"cd",  x"28", -- 1880
         x"35",  x"69",  x"e5",  x"b9",  x"f7",  x"23",  x"8f",  x"4b", -- 1888
         x"a0",  x"39",  x"72",  x"86",  x"30",  x"12",  x"9e",  x"27", -- 1890
         x"b3",  x"71",  x"e8",  x"53",  x"c0",  x"10",  x"8f",  x"ea", -- 1898
         x"02",  x"d1",  x"cd",  x"1b",  x"d3",  x"b9",  x"66",  x"66", -- 18A0
         x"06",  x"c4",  x"ed",  x"fa",  x"a2",  x"e3",  x"c2",  x"71", -- 18A8
         x"f7",  x"c2",  x"e6",  x"cb",  x"60",  x"21",  x"d4",  x"7e", -- 18B0
         x"45",  x"47",  x"8b",  x"fc",  x"76",  x"5b",  x"1f",  x"88", -- 18B8
         x"2b",  x"a2",  x"09",  x"78",  x"ca",  x"92",  x"e8",  x"01", -- 18C0
         x"87",  x"c9",  x"fe",  x"2c",  x"c0",  x"b7",  x"a6",  x"65", -- 18C8
         x"50",  x"93",  x"88",  x"e1",  x"1a",  x"a9",  x"67",  x"25", -- 18D0
         x"29",  x"fd",  x"44",  x"20",  x"08",  x"23",  x"93",  x"60", -- 18D8
         x"fe",  x"d4",  x"20",  x"4a",  x"f8",  x"e1",  x"02",  x"da", -- 18E0
         x"07",  x"ca",  x"c3",  x"91",  x"2d",  x"48",  x"be",  x"83", -- 18E8
         x"07",  x"99",  x"c5",  x"fd",  x"68",  x"60",  x"88",  x"28", -- 18F0
         x"42",  x"5e",  x"1b",  x"d5",  x"38",  x"09",  x"e3",  x"98", -- 18F8
         x"82",  x"0f",  x"06",  x"e0",  x"fe",  x"a5",  x"4e",  x"02", -- 1900
         x"cb",  x"fe",  x"a8",  x"28",  x"78",  x"e5",  x"50",  x"01", -- 1908
         x"28",  x"5d",  x"fe",  x"3b",  x"ca",  x"b2",  x"cb",  x"90", -- 1910
         x"84",  x"55",  x"e5",  x"8c",  x"c3",  x"eb",  x"a4",  x"ef", -- 1918
         x"c0",  x"34",  x"d8",  x"cd",  x"8a",  x"11",  x"d1",  x"36", -- 1920
         x"20",  x"be",  x"8c",  x"34",  x"03",  x"cd",  x"88",  x"c8", -- 1928
         x"85",  x"0a",  x"04",  x"cc",  x"8c",  x"0b",  x"86",  x"3d", -- 1930
         x"b8",  x"d4",  x"c9",  x"c2",  x"cc",  x"d1",  x"aa",  x"66", -- 1938
         x"a0",  x"0e",  x"21",  x"b7",  x"61",  x"05",  x"36",  x"00", -- 1940
         x"91",  x"b8",  x"3e",  x"66",  x"0d",  x"91",  x"b2",  x"0a", -- 1948
         x"04",  x"70",  x"40",  x"ac",  x"30",  x"40",  x"03",  x"3d", -- 1950
         x"c8",  x"f5",  x"62",  x"af",  x"0d",  x"f1",  x"a0",  x"a3", -- 1958
         x"3a",  x"42",  x"c6",  x"38",  x"d0",  x"37",  x"30",  x"29", -- 1960
         x"d6",  x"0d",  x"e0",  x"ab",  x"20",  x"fa",  x"12",  x"2f", -- 1968
         x"18",  x"15",  x"a9",  x"07",  x"1e",  x"d4",  x"cd",  x"db", -- 1970
         x"be",  x"13",  x"fa",  x"11",  x"a8",  x"e5",  x"91",  x"60", -- 1978
         x"1f",  x"2f",  x"83",  x"30",  x"2a",  x"0b",  x"3c",  x"a8", -- 1980
         x"7f",  x"47",  x"ed",  x"05",  x"10",  x"fb",  x"a8",  x"ad", -- 1988
         x"8b",  x"94",  x"69",  x"85",  x"8a",  x"32",  x"7d",  x"8c", -- 1990
         x"57",  x"88",  x"b1",  x"40",  x"08",  x"00",  x"3f",  x"52", -- 1998
         x"45",  x"44",  x"4f",  x"20",  x"46",  x"0e",  x"52",  x"4f", -- 19A0
         x"4d",  x"20",  x"b1",  x"06",  x"41",  x"52",  x"54",  x"81", -- 19A8
         x"04",  x"3a",  x"ce",  x"9f",  x"e2",  x"42",  x"e6",  x"62", -- 19B0
         x"21",  x"c9",  x"2c",  x"09",  x"c9",  x"d1",  x"c3",  x"85", -- 19B8
         x"fd",  x"8d",  x"37",  x"d1",  x"c1",  x"ca",  x"bd",  x"d4", -- 19C0
         x"7e",  x"9f",  x"c1",  x"20",  x"10",  x"cd",  x"8b",  x"0e", -- 19C8
         x"48",  x"a6",  x"3b",  x"91",  x"d5",  x"cc",  x"07",  x"04", -- 19D0
         x"d4",  x"c6",  x"18",  x"04",  x"08",  x"cf",  x"0e",  x"c6", -- 19D8
         x"c1",  x"38",  x"36",  x"bb",  x"49",  x"af",  x"1c",  x"2b", -- 19E0
         x"d5",  x"08",  x"37",  x"36",  x"2c",  x"c2",  x"a6",  x"a7", -- 19E8
         x"b1",  x"ab",  x"f6",  x"31",  x"4c",  x"49",  x"e3",  x"82", -- 19F0
         x"a9",  x"f1",  x"27",  x"d0",  x"0a",  x"e3",  x"d5",  x"3c", -- 19F8
         x"98",  x"46",  x"1e",  x"5c",  x"9a",  x"20",  x"7d",  x"ee", -- 1A00
         x"c6",  x"36",  x"03",  x"d1",  x"c1",  x"da",  x"1f",  x"c9", -- 1A08
         x"38",  x"a1",  x"ca",  x"47",  x"ca",  x"f0",  x"3b",  x"e0", -- 1A10
         x"72",  x"21",  x"a8",  x"31",  x"57",  x"f2",  x"e9",  x"e2", -- 1A18
         x"96",  x"2c",  x"ac",  x"57",  x"d5",  x"09",  x"16",  x"3a", -- 1A20
         x"06",  x"2c",  x"94",  x"8b",  x"8e",  x"d1",  x"c0",  x"88", -- 1A28
         x"88",  x"cc",  x"46",  x"c3",  x"77",  x"5a",  x"ca",  x"a1", -- 1A30
         x"89",  x"a1",  x"d7",  x"e3",  x"d6",  x"c4",  x"e1",  x"92", -- 1A38
         x"e4",  x"b5",  x"d0",  x"58",  x"c2",  x"db",  x"cb",  x"a1", -- 1A40
         x"0e",  x"0a",  x"20",  x"93",  x"d1",  x"33",  x"a2",  x"eb", -- 1A48
         x"c2",  x"f4",  x"e4",  x"a0",  x"b6",  x"21",  x"ab",  x"cc", -- 1A50
         x"27",  x"c4",  x"c9",  x"f7",  x"00",  x"3f",  x"45",  x"58", -- 1A58
         x"54",  x"52",  x"41",  x"04",  x"20",  x"49",  x"47",  x"4e", -- 1A60
         x"4f",  x"eb",  x"64",  x"df",  x"59",  x"d2",  x"91",  x"82", -- 1A68
         x"31",  x"11",  x"da",  x"4b",  x"1e",  x"06",  x"f7",  x"4c", -- 1A70
         x"dc",  x"64",  x"ca",  x"03",  x"c0",  x"54",  x"fe",  x"83", -- 1A78
         x"20",  x"e2",  x"a9",  x"b6",  x"cc",  x"d4",  x"68",  x"c4", -- 1A80
         x"8a",  x"b0",  x"f3",  x"92",  x"bc",  x"b0",  x"c2",  x"4e", -- 1A88
         x"12",  x"c3",  x"f9",  x"d5",  x"2a",  x"f5",  x"b3",  x"c3", -- 1A90
         x"dd",  x"d6",  x"dd",  x"2d",  x"f3",  x"16",  x"d4",  x"71", -- 1A98
         x"75",  x"97",  x"ee",  x"d6",  x"83",  x"c1",  x"c1",  x"90", -- 1AA0
         x"09",  x"97",  x"e1",  x"66",  x"9b",  x"e8",  x"c5",  x"c3", -- 1AA8
         x"0c",  x"50",  x"c8",  x"f9",  x"2a",  x"bc",  x"d8",  x"8d", -- 1AB0
         x"aa",  x"da",  x"8d",  x"a2",  x"29",  x"df",  x"cc",  x"80", -- 1AB8
         x"08",  x"f6",  x"37",  x"d4",  x"c0",  x"8f",  x"b7",  x"e8", -- 1AC0
         x"1e",  x"5e",  x"18",  x"c9",  x"a2",  x"cc",  x"ad",  x"3c", -- 1AC8
         x"2b",  x"16",  x"bf",  x"2d",  x"0e",  x"01",  x"c7",  x"01", -- 1AD0
         x"cd",  x"ad",  x"cd",  x"22",  x"d1",  x"9a",  x"84",  x"02", -- 1AD8
         x"c1",  x"f8",  x"fa",  x"78",  x"d4",  x"55",  x"29",  x"80", -- 1AE0
         x"18",  x"06",  x"d6",  x"b3",  x"38",  x"15",  x"c7",  x"15", -- 1AE8
         x"cb",  x"01",  x"fe",  x"01",  x"17",  x"aa",  x"ba",  x"57", -- 1AF0
         x"cd",  x"78",  x"22",  x"46",  x"c6",  x"97",  x"89",  x"18", -- 1AF8
         x"e7",  x"7a",  x"91",  x"86",  x"84",  x"ce",  x"7e",  x"0d", -- 1B00
         x"1d",  x"d6",  x"ac",  x"e7",  x"0c",  x"07",  x"d0",  x"5f", -- 1B08
         x"53",  x"00",  x"3d",  x"b3",  x"7b",  x"ca",  x"b3",  x"d2", -- 1B10
         x"07",  x"83",  x"2e",  x"5f",  x"21",  x"c9",  x"02",  x"19", -- 1B18
         x"78",  x"56",  x"ba",  x"d0",  x"23",  x"b7",  x"b0",  x"c5", -- 1B20
         x"01",  x"47",  x"49",  x"03",  x"43",  x"4a",  x"a0",  x"03", -- 1B28
         x"d6",  x"58",  x"51",  x"dc",  x"77",  x"a2",  x"c8",  x"32", -- 1B30
         x"18",  x"90",  x"99",  x"88",  x"ae",  x"46",  x"a4",  x"1e", -- 1B38
         x"24",  x"ee",  x"62",  x"da",  x"b8",  x"42",  x"cd",  x"8f", -- 1B40
         x"a6",  x"c0",  x"37",  x"fe",  x"ac",  x"28",  x"08",  x"e8", -- 1B48
         x"fe",  x"2e",  x"ca",  x"0d",  x"fe",  x"ad",  x"24",  x"28", -- 1B50
         x"19",  x"ec",  x"4c",  x"ca",  x"d4",  x"fe",  x"00",  x"aa", -- 1B58
         x"ca",  x"e3",  x"ce",  x"fe",  x"a7",  x"ca",  x"f0",  x"00", -- 1B60
         x"d0",  x"d6",  x"b6",  x"30",  x"28",  x"cd",  x"36",  x"cd", -- 1B68
         x"50",  x"c3",  x"cd",  x"16",  x"08",  x"7d",  x"cd",  x"3d", -- 1B70
         x"cd",  x"a2",  x"c8",  x"ed",  x"8c",  x"c0",  x"d6",  x"5e", -- 1B78
         x"b4",  x"c4",  x"91",  x"98",  x"e5",  x"9c",  x"85",  x"c1", -- 1B80
         x"64",  x"a9",  x"e2",  x"cc",  x"92",  x"4a",  x"10",  x"bc", -- 1B88
         x"ed",  x"db",  x"18",  x"c5",  x"5c",  x"79",  x"0b",  x"fe", -- 1B90
         x"33",  x"38",  x"07",  x"8d",  x"5d",  x"e3",  x"13",  x"e0", -- 1B98
         x"bb",  x"80",  x"1e",  x"fe",  x"2d",  x"38",  x"17",  x"c9", -- 1BA0
         x"43",  x"fc",  x"d6",  x"2a",  x"ec",  x"d5",  x"f3",  x"8a", -- 1BA8
         x"e3",  x"37",  x"f4",  x"91",  x"eb",  x"90",  x"47",  x"ac", -- 1BB0
         x"12",  x"bf",  x"16",  x"e3",  x"11",  x"f2",  x"70",  x"96", -- 1BB8
         x"94",  x"dd",  x"8f",  x"08",  x"66",  x"69",  x"e9",  x"15", -- 1BC0
         x"83",  x"90",  x"c8",  x"2f",  x"c8",  x"14",  x"fe",  x"4a", -- 1BC8
         x"2b",  x"06",  x"ac",  x"c1",  x"94",  x"c9",  x"b9",  x"2f", -- 1BD0
         x"f5",  x"83",  x"72",  x"fe",  x"08",  x"f1",  x"eb",  x"c1", -- 1BD8
         x"e3",  x"35",  x"e0",  x"d6",  x"b0",  x"0e",  x"0b",  x"c1", -- 1BE0
         x"79",  x"00",  x"21",  x"b0",  x"d0",  x"20",  x"05",  x"a3", -- 1BE8
         x"4f",  x"78",  x"10",  x"a2",  x"e9",  x"b3",  x"04",  x"b2", -- 1BF0
         x"e9",  x"21",  x"23",  x"96",  x"ce",  x"86",  x"06",  x"1f", -- 1BF8
         x"7a",  x"17",  x"ea",  x"44",  x"64",  x"78",  x"ff",  x"40", -- 1C00
         x"c3",  x"97",  x"cd",  x"98",  x"ce",  x"05",  x"79",  x"b7", -- 1C08
         x"1f",  x"c1",  x"d1",  x"2e",  x"ae",  x"40",  x"21",  x"d9", -- 1C10
         x"ce",  x"26",  x"e5",  x"ca",  x"a2",  x"8d",  x"fa",  x"98", -- 1C18
         x"bb",  x"fe",  x"d2",  x"61",  x"7e",  x"b4",  x"8f",  x"28", -- 1C20
         x"d1",  x"44",  x"c5",  x"1a",  x"02",  x"d3",  x"b3",  x"e0", -- 1C28
         x"f1",  x"57",  x"e1",  x"00",  x"7b",  x"b2",  x"c8",  x"7a", -- 1C30
         x"d6",  x"01",  x"d8",  x"af",  x"03",  x"bb",  x"3c",  x"d0", -- 1C38
         x"15",  x"1d",  x"0a",  x"81",  x"8d",  x"9c",  x"00",  x"ed", -- 1C40
         x"3f",  x"c3",  x"a2",  x"d6",  x"3c",  x"00",  x"8f",  x"c1", -- 1C48
         x"a0",  x"c6",  x"ff",  x"9f",  x"c3",  x"a9",  x"11",  x"d6", -- 1C50
         x"16",  x"5a",  x"fb",  x"91",  x"87",  x"c8",  x"7b",  x"2f", -- 1C58
         x"4f",  x"11",  x"7a",  x"2f",  x"cd",  x"7d",  x"c1",  x"c3", -- 1C60
         x"de",  x"25",  x"e6",  x"22",  x"c8",  x"d5",  x"30",  x"01", -- 1C68
         x"fa",  x"2b",  x"ce",  x"c5",  x"e1",  x"04",  x"ad",  x"03", -- 1C70
         x"46",  x"ce",  x"a4",  x"a9",  x"e1",  x"af",  x"4f",  x"e4", -- 1C78
         x"2c",  x"98",  x"38",  x"05",  x"0f",  x"38",  x"35",  x"0b", -- 1C80
         x"4f",  x"0a",  x"fb",  x"e9",  x"2a",  x"f6",  x"06",  x"d6", -- 1C88
         x"24",  x"20",  x"0a",  x"3c",  x"1c",  x"1a",  x"0f",  x"81", -- 1C90
         x"14",  x"3a",  x"f0",  x"d8",  x"3d",  x"ca",  x"01",  x"dd", -- 1C98
         x"cf",  x"f2",  x"48",  x"cf",  x"7e",  x"d6",  x"e4",  x"d2", -- 1CA0
         x"6f",  x"41",  x"81",  x"0f",  x"e5",  x"50",  x"59",  x"2a", -- 1CA8
         x"df",  x"bc",  x"9a",  x"11",  x"01",  x"e1",  x"03",  x"ca", -- 1CB0
         x"e0",  x"d5",  x"2a",  x"d9",  x"84",  x"c6",  x"8c",  x"e6", -- 1CB8
         x"0f",  x"6c",  x"ae",  x"79",  x"04",  x"96",  x"23",  x"20", -- 1CC0
         x"02",  x"78",  x"04",  x"28",  x"31",  x"38",  x"23",  x"00", -- 1CC8
         x"18",  x"cf",  x"b5",  x"ff",  x"4b",  x"11",  x"55",  x"f0", -- 1CD0
         x"37",  x"d8",  x"a9",  x"d0",  x"26",  x"ed",  x"90",  x"fd", -- 1CD8
         x"2a",  x"db",  x"9f",  x"3f",  x"09",  x"a7",  x"86",  x"ab", -- 1CE0
         x"c4",  x"e0",  x"96",  x"0a",  x"fa",  x"89",  x"22",  x"3d", -- 1CE8
         x"2b",  x"c0",  x"86",  x"21",  x"64",  x"b7",  x"d1",  x"08", -- 1CF0
         x"73",  x"23",  x"72",  x"23",  x"32",  x"c9",  x"32",  x"74", -- 1CF8
         x"e8",  x"90",  x"20",  x"a2",  x"ca",  x"82",  x"6d",  x"8a", -- 1D00
         x"42",  x"2a",  x"ad",  x"88",  x"62",  x"57",  x"d5",  x"b0", -- 1D08
         x"61",  x"5b",  x"c9",  x"c1",  x"dc",  x"24",  x"92",  x"e1", -- 1D10
         x"3c",  x"57",  x"96",  x"7a",  x"ee",  x"c4",  x"b8",  x"ac", -- 1D18
         x"8b",  x"a2",  x"41",  x"1d",  x"1e",  x"00",  x"61",  x"e2", -- 1D20
         x"ce",  x"83",  x"30",  x"3e",  x"19",  x"28",  x"ed",  x"5b", -- 1D28
         x"50",  x"85",  x"db",  x"aa",  x"11",  x"b9",  x"85",  x"85", -- 1D30
         x"7e",  x"b8",  x"a9",  x"ac",  x"08",  x"e8",  x"55",  x"3a", -- 1D38
         x"24",  x"8d",  x"00",  x"51",  x"c3",  x"f1",  x"44",  x"4d", -- 1D40
         x"ca",  x"aa",  x"02",  x"cf",  x"96",  x"28",  x"5f",  x"1e", -- 1D48
         x"10",  x"d9",  x"b0",  x"11",  x"04",  x"00",  x"00",  x"f1", -- 1D50
         x"ca",  x"67",  x"c9",  x"71",  x"23",  x"70",  x"2b",  x"23", -- 1D58
         x"4f",  x"db",  x"22",  x"ab",  x"ac",  x"ab",  x"b0",  x"0c", -- 1D60
         x"2a",  x"17",  x"79",  x"01",  x"01",  x"0b",  x"00",  x"30", -- 1D68
         x"02",  x"c1",  x"03",  x"1a",  x"a4",  x"f5",  x"e5",  x"4f", -- 1D70
         x"d7",  x"88",  x"91",  x"f1",  x"3d",  x"01",  x"20",  x"ea", -- 1D78
         x"f5",  x"42",  x"4b",  x"eb",  x"19",  x"f7",  x"c8",  x"cd", -- 1D80
         x"45",  x"30",  x"99",  x"66",  x"47",  x"b2",  x"65",  x"03", -- 1D88
         x"57",  x"b0",  x"60",  x"5e",  x"eb",  x"29",  x"08",  x"09", -- 1D90
         x"eb",  x"2b",  x"2b",  x"bd",  x"d0",  x"f1",  x"38",  x"22", -- 1D98
         x"47",  x"4c",  x"4f",  x"bb",  x"16",  x"69",  x"e1",  x"7a", -- 1DA0
         x"e3",  x"f5",  x"e0",  x"ba",  x"90",  x"d2",  x"43",  x"d1", -- 1DA8
         x"19",  x"43",  x"a2",  x"7f",  x"8b",  x"15",  x"29",  x"29", -- 1DB0
         x"c1",  x"2a",  x"9f",  x"62",  x"c9",  x"ab",  x"35",  x"21", -- 1DB8
         x"b7",  x"73",  x"39",  x"c1",  x"18",  x"4e",  x"0d",  x"f0", -- 1DC0
         x"0b",  x"cd",  x"09",  x"d2",  x"13",  x"9b",  x"81",  x"2a", -- 1DC8
         x"c4",  x"03",  x"e2",  x"d3",  x"4f",  x"e2",  x"a1",  x"41", -- 1DD0
         x"50",  x"1e",  x"d5",  x"a4",  x"1b",  x"73",  x"06",  x"06", -- 1DD8
         x"90",  x"c3",  x"ae",  x"d6",  x"9c",  x"a0",  x"47",  x"af", -- 1DE0
         x"18",  x"0c",  x"ed",  x"cd",  x"45",  x"d1",  x"da",  x"c6", -- 1DE8
         x"01",  x"8e",  x"05",  x"c5",  x"d5",  x"98",  x"ed",  x"da", -- 1DF0
         x"70",  x"2b",  x"09",  x"56",  x"2b",  x"5e",  x"e1",  x"f4", -- 1DF8
         x"d9",  x"90",  x"3b",  x"82",  x"64",  x"63",  x"e3",  x"b7", -- 1E00
         x"61",  x"c3",  x"84",  x"28",  x"55",  x"2b",  x"24",  x"18", -- 1E08
         x"19",  x"88",  x"e3",  x"8a",  x"d0",  x"7a",  x"b3",  x"ca", -- 1E10
         x"54",  x"2a",  x"c3",  x"7e",  x"bb",  x"27",  x"6f",  x"e5", -- 1E18
         x"b9",  x"3a",  x"9e",  x"84",  x"03",  x"2a",  x"e3",  x"03", -- 1E20
         x"0a",  x"e1",  x"95",  x"03",  x"21",  x"03",  x"27",  x"a1", -- 1E28
         x"8b",  x"c1",  x"f9",  x"e2",  x"ec",  x"49",  x"d3",  x"11", -- 1E30
         x"55",  x"03",  x"1d",  x"03",  x"24",  x"4a",  x"ff",  x"fb", -- 1E38
         x"84",  x"01",  x"e1",  x"c0",  x"1e",  x"16",  x"8e",  x"8c", -- 1E40
         x"8a",  x"a7",  x"3e",  x"80",  x"81",  x"40",  x"b6",  x"47", -- 1E48
         x"cd",  x"0b",  x"33",  x"cf",  x"c3",  x"75",  x"02",  x"39", -- 1E50
         x"a9",  x"88",  x"c0",  x"c0",  x"01",  x"57",  x"d3",  x"c5", -- 1E58
         x"ac",  x"b5",  x"59",  x"e5",  x"75",  x"c3",  x"56",  x"ba", -- 1E60
         x"60",  x"9e",  x"d1",  x"01",  x"e5",  x"6f",  x"cd",  x"f2", -- 1E68
         x"d2",  x"d1",  x"c9",  x"10",  x"9d",  x"eb",  x"85",  x"e5", -- 1E70
         x"77",  x"1b",  x"a1",  x"29",  x"52",  x"00",  x"2b",  x"06", -- 1E78
         x"22",  x"50",  x"e5",  x"0e",  x"ff",  x"99",  x"a4",  x"0c", -- 1E80
         x"f8",  x"10",  x"06",  x"ba",  x"28",  x"e0",  x"96",  x"20", -- 1E88
         x"f4",  x"b0",  x"ff",  x"cc",  x"bd",  x"f2",  x"dc",  x"fa", -- 1E90
         x"66",  x"79",  x"34",  x"21",  x"11",  x"2a",  x"2a",  x"b2", -- 1E98
         x"03",  x"fc",  x"38",  x"3e",  x"56",  x"01",  x"a0",  x"f9", -- 1EA0
         x"8f",  x"c3",  x"28",  x"22",  x"88",  x"10",  x"e1",  x"7e", -- 1EA8
         x"82",  x"8c",  x"1e",  x"c3",  x"fd",  x"ce",  x"6c",  x"6d", -- 1EB0
         x"92",  x"07",  x"1c",  x"1d",  x"c8",  x"ed",  x"28",  x"fe", -- 1EB8
         x"0d",  x"cc",  x"30",  x"66",  x"cb",  x"b3",  x"04",  x"f2", -- 1EC0
         x"b7",  x"0e",  x"f1",  x"f5",  x"c0",  x"b5",  x"fc",  x"50", -- 1EC8
         x"06",  x"ff",  x"09",  x"ab",  x"28",  x"37",  x"e0",  x"94", -- 1ED0
         x"22",  x"0d",  x"56",  x"f1",  x"b8",  x"8b",  x"1e",  x"1a", -- 1ED8
         x"01",  x"28",  x"c2",  x"bf",  x"f5",  x"01",  x"e3",  x"d1", -- 1EE0
         x"e0",  x"82",  x"b0",  x"5c",  x"4a",  x"c4",  x"fa",  x"c5", -- 1EE8
         x"da",  x"2c",  x"44",  x"fe",  x"b4",  x"56",  x"03",  x"34", -- 1EF0
         x"5d",  x"2b",  x"02",  x"01",  x"1a",  x"d2",  x"20",  x"3f", -- 1EF8
         x"c6",  x"b2",  x"0e",  x"53",  x"d9",  x"c4",  x"08",  x"0a", -- 1F00
         x"cb",  x"c0",  x"b7",  x"cd",  x"68",  x"d2",  x"14",  x"18", -- 1F08
         x"ee",  x"c1",  x"d7",  x"db",  x"49",  x"75",  x"15",  x"7b", -- 1F10
         x"bc",  x"05",  x"b7",  x"f2",  x"3b",  x"d2",  x"ad",  x"24", -- 1F18
         x"e4",  x"55",  x"cc",  x"2b",  x"09",  x"66",  x"1c",  x"f2", -- 1F20
         x"33",  x"1c",  x"02",  x"da",  x"01",  x"59",  x"d2",  x"e0", -- 1F28
         x"c6",  x"80",  x"35",  x"4a",  x"ef",  x"bc",  x"f0",  x"97", -- 1F30
         x"9a",  x"8a",  x"8a",  x"33",  x"19",  x"2a",  x"e2",  x"59", -- 1F38
         x"d8",  x"85",  x"07",  x"95",  x"bc",  x"4a",  x"09",  x"d0", -- 1F40
         x"c4",  x"8a",  x"f1",  x"e5",  x"cd",  x"b7",  x"e5",  x"0c", -- 1F48
         x"7d",  x"b4",  x"b7",  x"02",  x"46",  x"2b",  x"4e",  x"e5", -- 1F50
         x"b6",  x"82",  x"6e",  x"26",  x"46",  x"b1",  x"d0",  x"2b", -- 1F58
         x"2e",  x"ca",  x"ae",  x"95",  x"c9",  x"bf",  x"cd",  x"9b", -- 1F60
         x"84",  x"2b",  x"c3",  x"0c",  x"4d",  x"e5",  x"cd",  x"85", -- 1F68
         x"d4",  x"f5",  x"92",  x"03",  x"2a",  x"98",  x"68",  x"0c", -- 1F70
         x"e5",  x"86",  x"1e",  x"27",  x"1c",  x"da",  x"86",  x"09", -- 1F78
         x"7b",  x"d1",  x"83",  x"30",  x"96",  x"88",  x"16",  x"01", -- 1F80
         x"d3",  x"15",  x"c2",  x"03",  x"c0",  x"f0",  x"e9",  x"d2", -- 1F88
         x"c4",  x"02",  x"21",  x"f2",  x"91",  x"62",  x"18",  x"6f", -- 1F90
         x"6b",  x"63",  x"ba",  x"22",  x"6f",  x"2c",  x"2d",  x"9f", -- 1F98
         x"40",  x"12",  x"03",  x"13",  x"18",  x"66",  x"f8",  x"3d", -- 1FA0
         x"3b",  x"40",  x"25",  x"1b",  x"d3",  x"eb",  x"c0",  x"d5", -- 1FA8
         x"88",  x"69",  x"1b",  x"4e",  x"97",  x"e7",  x"99",  x"22", -- 1FB0
         x"47",  x"09",  x"89",  x"52",  x"90",  x"69",  x"ee",  x"48", -- 1FB8
         x"8a",  x"d8",  x"89",  x"b1",  x"14",  x"c0",  x"ea",  x"28", -- 1FC0
         x"c9",  x"16",  x"01",  x"c0",  x"d0",  x"f0",  x"04",  x"fb", -- 1FC8
         x"d2",  x"af",  x"57",  x"80",  x"e7",  x"e9",  x"5c",  x"0e", -- 1FD0
         x"84",  x"30",  x"d3",  x"28",  x"55",  x"da",  x"70",  x"1a", -- 1FD8
         x"4d",  x"c9",  x"98",  x"80",  x"18",  x"cd",  x"30",  x"24", -- 1FE0
         x"d4",  x"7a",  x"73",  x"c1",  x"c2",  x"f7",  x"0a",  x"02", -- 1FE8
         x"da",  x"d3",  x"af",  x"e3",  x"4f",  x"e5",  x"ef",  x"c5", -- 1FF0
         x"38",  x"f9",  x"c2",  x"11",  x"0e",  x"00",  x"2b",  x"78", -- 1FF8
         x"e1",  x"a6",  x"e1",  x"4a",  x"e5",  x"2c",  x"46",  x"ee", -- 2000
         x"12",  x"68",  x"a2",  x"91",  x"d8",  x"4e",  x"d5",  x"53", -- 2008
         x"89",  x"11",  x"b3",  x"86",  x"18",  x"cf",  x"2d",  x"54", -- 2010
         x"99",  x"1a",  x"34",  x"90",  x"18",  x"e3",  x"02",  x"7e", -- 2018
         x"cd",  x"de",  x"d3",  x"04",  x"05",  x"84",  x"f0",  x"c5", -- 2020
         x"1e",  x"14",  x"ff",  x"fe",  x"29",  x"8b",  x"6a",  x"fa", -- 2028
         x"e9",  x"f0",  x"c8",  x"58",  x"f1",  x"14",  x"e3",  x"01", -- 2030
         x"61",  x"cb",  x"12",  x"3d",  x"be",  x"3c",  x"d0",  x"cb", -- 2038
         x"c0",  x"91",  x"bb",  x"47",  x"d8",  x"30",  x"43",  x"c9", -- 2040
         x"7f",  x"ca",  x"cf",  x"2a",  x"d4",  x"5f",  x"54",  x"c3", -- 2048
         x"e0",  x"19",  x"46",  x"28",  x"72",  x"e3",  x"eb",  x"f4", -- 2050
         x"d2",  x"86",  x"67",  x"70",  x"c9",  x"eb",  x"31",  x"26", -- 2058
         x"c1",  x"d7",  x"c8",  x"23",  x"92",  x"82",  x"4f",  x"ed", -- 2060
         x"78",  x"c3",  x"ad",  x"21",  x"cd",  x"14",  x"d4",  x"81", -- 2068
         x"f0",  x"03",  x"4f",  x"7b",  x"29",  x"ed",  x"79",  x"13", -- 2070
         x"0a",  x"f5",  x"c8",  x"67",  x"f4",  x"af",  x"5e",  x"4d", -- 2078
         x"c1",  x"19",  x"82",  x"25",  x"ab",  x"a0",  x"28",  x"fa", -- 2080
         x"1c",  x"96",  x"0e",  x"32",  x"0d",  x"17",  x"45",  x"f9", -- 2088
         x"fd",  x"d9",  x"80",  x"68",  x"61",  x"76",  x"c9",  x"b7", -- 2090
         x"45",  x"8f",  x"2e",  x"8b",  x"7b",  x"04",  x"c5",  x"40", -- 2098
         x"1a",  x"18",  x"b2",  x"cd",  x"1c",  x"6c",  x"c9",  x"d5", -- 20A0
         x"38",  x"9a",  x"d1",  x"12",  x"12",  x"eb",  x"44",  x"46", -- 20A8
         x"81",  x"c3",  x"3b",  x"b1",  x"d0",  x"16",  x"95",  x"06", -- 20B0
         x"e3",  x"d3",  x"c0",  x"21",  x"04",  x"d9",  x"a4",  x"9b", -- 20B8
         x"31",  x"18",  x"09",  x"04",  x"21",  x"8b",  x"17",  x"fb", -- 20C0
         x"21",  x"78",  x"b7",  x"b8",  x"a2",  x"e8",  x"d9",  x"e7", -- 20C8
         x"ca",  x"8a",  x"00",  x"90",  x"30",  x"0c",  x"2f",  x"3c", -- 20D0
         x"76",  x"eb",  x"e0",  x"72",  x"97",  x"c3",  x"1b",  x"fe", -- 20D8
         x"19",  x"d0",  x"95",  x"00",  x"03",  x"d7",  x"67",  x"f1", -- 20E0
         x"98",  x"93",  x"d5",  x"b4",  x"4c",  x"21",  x"96",  x"f2", -- 20E8
         x"44",  x"ab",  x"f1",  x"0a",  x"00",  x"d5",  x"30",  x"4b", -- 20F0
         x"23",  x"34",  x"28",  x"63",  x"2e",  x"90",  x"d8",  x"3e", -- 20F8
         x"d5",  x"00",  x"18",  x"40",  x"af",  x"90",  x"47",  x"7e", -- 2100
         x"9b",  x"5f",  x"88",  x"67",  x"9a",  x"57",  x"03",  x"99", -- 2108
         x"4f",  x"01",  x"dc",  x"16",  x"d5",  x"68",  x"63",  x"af", -- 2110
         x"47",  x"a7",  x"c0",  x"20",  x"16",  x"4a",  x"00",  x"54", -- 2118
         x"65",  x"6f",  x"78",  x"d6",  x"08",  x"fe",  x"e0",  x"36", -- 2120
         x"20",  x"f0",  x"86",  x"80",  x"5d",  x"c9",  x"05",  x"29", -- 2128
         x"cb",  x"12",  x"cb",  x"01",  x"11",  x"f2",  x"d4",  x"d4", -- 2130
         x"78",  x"5c",  x"45",  x"cb",  x"61",  x"08",  x"21",  x"12", -- 2138
         x"00",  x"86",  x"77",  x"30",  x"e5",  x"c8",  x"78",  x"21", -- 2140
         x"c1",  x"79",  x"fc",  x"fd",  x"d4",  x"aa",  x"18",  x"e6", -- 2148
         x"08",  x"80",  x"a9",  x"4f",  x"c3",  x"76",  x"1c",  x"c0", -- 2150
         x"00",  x"14",  x"c0",  x"0c",  x"c0",  x"0e",  x"80",  x"34", -- 2158
         x"c0",  x"06",  x"c3",  x"53",  x"d6",  x"7e",  x"83",  x"5b", -- 2160
         x"30",  x"8a",  x"5b",  x"89",  x"4f",  x"89",  x"b7",  x"e9", -- 2168
         x"e0",  x"30",  x"2f",  x"77",  x"af",  x"49",  x"6f",  x"71", -- 2170
         x"7d",  x"71",  x"7d",  x"70",  x"2f",  x"7d",  x"6f",  x"a0", -- 2178
         x"4a",  x"62",  x"b8",  x"c1",  x"43",  x"5a",  x"51",  x"ca", -- 2180
         x"30",  x"18",  x"f5",  x"c6",  x"6c",  x"09",  x"f1",  x"2d", -- 2188
         x"f0",  x"ab",  x"1f",  x"4f",  x"02",  x"cb",  x"1a",  x"cb", -- 2190
         x"1b",  x"cb",  x"18",  x"e6",  x"c4",  x"00",  x"00",  x"81", -- 2198
         x"00",  x"03",  x"aa",  x"56",  x"19",  x"80",  x"f1",  x"22", -- 21A0
         x"76",  x"00",  x"80",  x"45",  x"aa",  x"38",  x"82",  x"cd", -- 21A8
         x"97",  x"d6",  x"24",  x"b7",  x"ea",  x"b3",  x"c0",  x"73", -- 21B0
         x"7e",  x"01",  x"35",  x"80",  x"f0",  x"a6",  x"04",  x"90", -- 21B8
         x"37",  x"f5",  x"70",  x"af",  x"08",  x"6f",  x"d4",  x"eb", -- 21C0
         x"80",  x"04",  x"cd",  x"f5",  x"d5",  x"21",  x"48",  x"90", -- 21C8
         x"a8",  x"66",  x"d4",  x"20",  x"21",  x"4c",  x"05",  x"ce", -- 21D0
         x"d9",  x"01",  x"80",  x"ac",  x"1f",  x"3e",  x"1a",  x"60", -- 21D8
         x"f1",  x"bd",  x"d8",  x"22",  x"01",  x"31",  x"0c",  x"18", -- 21E0
         x"72",  x"ad",  x"56",  x"40",  x"20",  x"c8",  x"2e",  x"15", -- 21E8
         x"58",  x"d6",  x"79",  x"32",  x"54",  x"f7",  x"a5",  x"22", -- 21F0
         x"d1",  x"d2",  x"01",  x"23",  x"01",  x"50",  x"58",  x"21", -- 21F8
         x"bc",  x"d4",  x"e5",  x"03",  x"14",  x"d5",  x"e5",  x"04", -- 2200
         x"a3",  x"93",  x"f3",  x"45",  x"dd",  x"06",  x"00",  x"2e", -- 2208
         x"08",  x"1f",  x"67",  x"79",  x"30",  x"0b",  x"aa",  x"f1", -- 2210
         x"21",  x"6c",  x"19",  x"92",  x"3a",  x"91",  x"2b",  x"89", -- 2218
         x"95",  x"d8",  x"2d",  x"7c",  x"20",  x"4d",  x"e4",  x"83", -- 2220
         x"b1",  x"19",  x"bc",  x"14",  x"e7",  x"a0",  x"01",  x"20", -- 2228
         x"84",  x"d9",  x"65",  x"ec",  x"5c",  x"5a",  x"06",  x"ca", -- 2230
         x"4b",  x"c3",  x"2e",  x"ff",  x"5c",  x"00",  x"34",  x"34", -- 2238
         x"2b",  x"7e",  x"32",  x"14",  x"03",  x"c6",  x"04",  x"10", -- 2240
         x"04",  x"87",  x"0c",  x"03",  x"41",  x"eb",  x"81",  x"80", -- 2248
         x"57",  x"5f",  x"32",  x"17",  x"03",  x"e9",  x"95",  x"7d", -- 2250
         x"8e",  x"10",  x"03",  x"de",  x"00",  x"19",  x"3f",  x"30", -- 2258
         x"07",  x"0d",  x"9f",  x"71",  x"37",  x"d2",  x"d5",  x"40", -- 2260
         x"79",  x"3c",  x"3d",  x"01",  x"1f",  x"fa",  x"ec",  x"d4", -- 2268
         x"17",  x"cb",  x"13",  x"e1",  x"2b",  x"e6",  x"21",  x"10", -- 2270
         x"3a",  x"19",  x"30",  x"17",  x"1d",  x"79",  x"b2",  x"34", -- 2278
         x"b3",  x"20",  x"f4",  x"8c",  x"eb",  x"03",  x"35",  x"e1", -- 2280
         x"20",  x"c7",  x"1e",  x"0a",  x"8f",  x"31",  x"78",  x"e3", -- 2288
         x"30",  x"7c",  x"d6",  x"7d",  x"c0",  x"11",  x"ae",  x"80", -- 2290
         x"47",  x"1f",  x"00",  x"a8",  x"78",  x"f2",  x"7b",  x"d6", -- 2298
         x"c6",  x"80",  x"77",  x"f4",  x"94",  x"9c",  x"e3",  x"11", -- 22A0
         x"77",  x"2b",  x"c9",  x"80",  x"80",  x"2f",  x"e1",  x"b7", -- 22A8
         x"e1",  x"f2",  x"a8",  x"ba",  x"18",  x"d1",  x"aa",  x"f0", -- 22B0
         x"95",  x"94",  x"c6",  x"02",  x"12",  x"38",  x"c7",  x"47", -- 22B8
         x"82",  x"99",  x"31",  x"8d",  x"31",  x"18",  x"bc",  x"a4", -- 22C0
         x"4b",  x"a9",  x"40",  x"e7",  x"03",  x"fe",  x"06",  x"2f", -- 22C8
         x"17",  x"9f",  x"c0",  x"3c",  x"2f",  x"91",  x"06",  x"88", -- 22D0
         x"bd",  x"98",  x"1d",  x"4f",  x"4c",  x"70",  x"88",  x"23", -- 22D8
         x"03",  x"36",  x"80",  x"17",  x"c3",  x"b9",  x"d4",  x"15", -- 22E0
         x"08",  x"f0",  x"21",  x"23",  x"7e",  x"ee",  x"aa",  x"59", -- 22E8
         x"80",  x"c5",  x"93",  x"92",  x"83",  x"0d",  x"f4",  x"8b", -- 22F0
         x"b8",  x"99",  x"49",  x"82",  x"05",  x"11",  x"db",  x"0f", -- 22F8
         x"18",  x"03",  x"f6",  x"21",  x"ed",  x"53",  x"17",  x"15", -- 2300
         x"ed",  x"43",  x"16",  x"df",  x"d3",  x"8a",  x"59",  x"09", -- 2308
         x"82",  x"ab",  x"4e",  x"80",  x"c2",  x"c9",  x"11",  x"0b", -- 2310
         x"01",  x"06",  x"04",  x"1a",  x"77",  x"13",  x"23",  x"10", -- 2318
         x"ee",  x"56",  x"42",  x"81",  x"07",  x"37",  x"1f",  x"77", -- 2320
         x"3f",  x"1f",  x"c6",  x"61",  x"77",  x"79",  x"09",  x"81", -- 2328
         x"4f",  x"1f",  x"ae",  x"c9",  x"bf",  x"19",  x"5d",  x"06", -- 2330
         x"21",  x"a0",  x"d6",  x"e5",  x"64",  x"18",  x"79",  x"c8", -- 2338
         x"22",  x"ae",  x"60",  x"79",  x"b0",  x"32",  x"00",  x"d7", -- 2340
         x"1f",  x"a9",  x"c9",  x"23",  x"78",  x"be",  x"c0",  x"31", -- 2348
         x"2b",  x"79",  x"03",  x"7a",  x"03",  x"81",  x"7b",  x"96", -- 2350
         x"c0",  x"e1",  x"e2",  x"22",  x"47",  x"b1",  x"52",  x"ae", -- 2358
         x"2a",  x"2a",  x"c9",  x"28",  x"de",  x"c0",  x"ae",  x"67", -- 2360
         x"fc",  x"69",  x"0a",  x"d7",  x"3e",  x"98",  x"90",  x"c8", -- 2368
         x"c1",  x"7c",  x"17",  x"dc",  x"ee",  x"44",  x"ae",  x"55", -- 2370
         x"aa",  x"90",  x"23",  x"1b",  x"7a",  x"a3",  x"14",  x"3c", -- 2378
         x"c0",  x"0b",  x"8f",  x"c0",  x"fe",  x"98",  x"3a",  x"97", -- 2380
         x"7e",  x"d0",  x"a7",  x"00",  x"45",  x"d7",  x"36",  x"98", -- 2388
         x"7b",  x"f5",  x"79",  x"22",  x"17",  x"cd",  x"ca",  x"db", -- 2390
         x"8a",  x"f9",  x"50",  x"78",  x"b1",  x"03",  x"c8",  x"3e", -- 2398
         x"10",  x"29",  x"38",  x"06",  x"b6",  x"c0",  x"eb",  x"30", -- 23A0
         x"04",  x"09",  x"1e",  x"da",  x"0b",  x"d0",  x"de",  x"40", -- 23A8
         x"17",  x"fe",  x"2d",  x"f5",  x"28",  x"05",  x"0b",  x"fe", -- 23B0
         x"2b",  x"28",  x"01",  x"8c",  x"a4",  x"ad",  x"5b",  x"47", -- 23B8
         x"67",  x"c4",  x"5e",  x"94",  x"00",  x"38",  x"3d",  x"fe", -- 23C0
         x"2e",  x"28",  x"16",  x"fe",  x"17",  x"45",  x"20",  x"15", -- 23C8
         x"a1",  x"a6",  x"4d",  x"ce",  x"12",  x"80",  x"4b",  x"14", -- 23D0
         x"20",  x"07",  x"af",  x"93",  x"5f",  x"00",  x"0c",  x"0c", -- 23D8
         x"28",  x"de",  x"e5",  x"7b",  x"90",  x"f4",  x"05",  x"ed", -- 23E0
         x"d7",  x"f2",  x"e4",  x"d7",  x"d2",  x"80",  x"e7",  x"d5", -- 23E8
         x"f1",  x"3c",  x"20",  x"0b",  x"f2",  x"d1",  x"f1",  x"cc", -- 23F0
         x"fb",  x"24",  x"97",  x"47",  x"c8",  x"0f",  x"82",  x"d6", -- 23F8
         x"f0",  x"97",  x"a3",  x"03",  x"57",  x"78",  x"89",  x"47", -- 2400
         x"c5",  x"f0",  x"4d",  x"0d",  x"29",  x"d6",  x"30",  x"f4", -- 2408
         x"14",  x"e1",  x"93",  x"14",  x"18",  x"a8",  x"a3",  x"85", -- 2410
         x"cd",  x"a9",  x"9d",  x"22",  x"c3",  x"85",  x"60",  x"7b", -- 2418
         x"07",  x"07",  x"83",  x"21",  x"07",  x"86",  x"1a",  x"5f", -- 2420
         x"18",  x"a5",  x"d5",  x"33",  x"0d",  x"d8",  x"4d",  x"98", -- 2428
         x"ca",  x"96",  x"0d",  x"06",  x"98",  x"86",  x"a4",  x"92", -- 2430
         x"22",  x"c8",  x"d1",  x"11",  x"ea",  x"03",  x"96",  x"55", -- 2438
         x"36",  x"57",  x"04",  x"42",  x"d8",  x"36",  x"2d",  x"8c", -- 2440
         x"c0",  x"30",  x"ca",  x"ef",  x"d8",  x"e5",  x"49",  x"fc", -- 2448
         x"60",  x"af",  x"5e",  x"f5",  x"bf",  x"50",  x"43",  x"91", -- 2450
         x"11",  x"44",  x"f8",  x"a3",  x"18",  x"02",  x"d7",  x"b7", -- 2458
         x"e2",  x"6e",  x"d8",  x"f1",  x"81",  x"68",  x"83",  x"88", -- 2460
         x"18",  x"ec",  x"85",  x"e3",  x"1c",  x"42",  x"cd",  x"5e", -- 2468
         x"d4",  x"3c",  x"f6",  x"32",  x"84",  x"b0",  x"01",  x"06", -- 2470
         x"a0",  x"d2",  x"81",  x"3c",  x"04",  x"fa",  x"89",  x"d8", -- 2478
         x"fe",  x"08",  x"eb",  x"40",  x"3c",  x"47",  x"3e",  x"02", -- 2480
         x"3d",  x"00",  x"3d",  x"e1",  x"f5",  x"11",  x"08",  x"d9", -- 2488
         x"05",  x"20",  x"18",  x"06",  x"36",  x"2e",  x"52",  x"23", -- 2490
         x"42",  x"05",  x"06",  x"cc",  x"f5",  x"d6",  x"a4",  x"35", -- 2498
         x"eb",  x"85",  x"f0",  x"06",  x"2f",  x"04",  x"91",  x"e9", -- 24A0
         x"5f",  x"ad",  x"f2",  x"9e",  x"9e",  x"e1",  x"79",  x"9e", -- 24A8
         x"4f",  x"91",  x"b1",  x"30",  x"f0",  x"9c",  x"88",  x"23", -- 24B0
         x"c6",  x"46",  x"eb",  x"e8",  x"40",  x"23",  x"c1",  x"0d", -- 24B8
         x"20",  x"d2",  x"09",  x"05",  x"28",  x"0b",  x"2b",  x"d7", -- 24C0
         x"19",  x"30",  x"bc",  x"48",  x"97",  x"c4",  x"81",  x"35", -- 24C8
         x"f1",  x"28",  x"1a",  x"36",  x"45",  x"44",  x"24",  x"2b", -- 24D0
         x"81",  x"8c",  x"9f",  x"c3",  x"e5",  x"3d",  x"00",  x"d6", -- 24D8
         x"0a",  x"30",  x"fb",  x"c6",  x"3a",  x"5e",  x"23",  x"2c", -- 24E0
         x"ed",  x"14",  x"71",  x"e1",  x"9f",  x"02",  x"74",  x"94", -- 24E8
         x"11",  x"f7",  x"23",  x"a3",  x"34",  x"e1",  x"e2",  x"17", -- 24F0
         x"65",  x"d8",  x"e9",  x"bb",  x"80",  x"80",  x"a0",  x"86", -- 24F8
         x"01",  x"10",  x"26",  x"27",  x"00",  x"9c",  x"25",  x"00", -- 2500
         x"64",  x"0c",  x"0a",  x"02",  x"eb",  x"68",  x"21",  x"88", -- 2508
         x"d0",  x"e3",  x"e9",  x"94",  x"93",  x"cd",  x"c3",  x"5b", -- 2510
         x"dd",  x"b4",  x"20",  x"78",  x"ca",  x"6d",  x"d9",  x"f2", -- 2518
         x"28",  x"38",  x"d9",  x"9a",  x"b2",  x"bc",  x"03",  x"2e", -- 2520
         x"d0",  x"d4",  x"ce",  x"11",  x"79",  x"f6",  x"7f",  x"9e", -- 2528
         x"82",  x"f2",  x"55",  x"d9",  x"d9",  x"f0",  x"70",  x"d7", -- 2530
         x"98",  x"23",  x"f5",  x"53",  x"e1",  x"0a",  x"7c",  x"1f", -- 2538
         x"e1",  x"22",  x"af",  x"29",  x"03",  x"e3",  x"84",  x"dc", -- 2540
         x"1a",  x"d9",  x"f7",  x"a6",  x"1b",  x"18",  x"59",  x"d5", -- 2548
         x"3f",  x"9a",  x"5e",  x"d5",  x"85",  x"83",  x"38",  x"81", -- 2550
         x"11",  x"3b",  x"aa",  x"0b",  x"2b",  x"e1",  x"01",  x"fe", -- 2558
         x"88",  x"d2",  x"76",  x"d6",  x"37",  x"96",  x"99",  x"54", -- 2560
         x"fd",  x"da",  x"98",  x"09",  x"f5",  x"93",  x"aa",  x"61", -- 2568
         x"d5",  x"92",  x"91",  x"ac",  x"6a",  x"49",  x"6c",  x"09", -- 2570
         x"8c",  x"3b",  x"21",  x"ad",  x"7c",  x"56",  x"d9",  x"f9", -- 2578
         x"08",  x"c1",  x"4a",  x"c3",  x"33",  x"08",  x"40",  x"00", -- 2580
         x"2e",  x"94",  x"74",  x"70",  x"4f",  x"2e",  x"77",  x"6e", -- 2588
         x"00",  x"02",  x"88",  x"7a",  x"e6",  x"a0",  x"2a",  x"7c", -- 2590
         x"50",  x"01",  x"aa",  x"aa",  x"7e",  x"ff",  x"ff",  x"7f", -- 2598
         x"7f",  x"c0",  x"18",  x"81",  x"cd",  x"81",  x"c0",  x"60", -- 25A0
         x"11",  x"98",  x"d5",  x"d5",  x"ae",  x"89",  x"26",  x"2e", -- 25A8
         x"e1",  x"0e",  x"61",  x"a3",  x"bc",  x"18",  x"06",  x"c2", -- 25B0
         x"50",  x"3d",  x"c8",  x"87",  x"25",  x"f5",  x"18",  x"15", -- 25B8
         x"b6",  x"95",  x"53",  x"07",  x"e3",  x"11",  x"e1",  x"18", -- 25C0
         x"dd",  x"56",  x"e2",  x"00",  x"1b",  x"03",  x"fa",  x"5d", -- 25C8
         x"da",  x"21",  x"3c",  x"66",  x"03",  x"26",  x"0b",  x"05", -- 25D0
         x"c8",  x"86",  x"e6",  x"07",  x"b0",  x"52",  x"a4",  x"0d", -- 25D8
         x"87",  x"87",  x"4f",  x"b4",  x"d8",  x"a7",  x"d0",  x"1a", -- 25E0
         x"03",  x"3c",  x"e6",  x"41",  x"03",  x"13",  x"fe",  x"01", -- 25E8
         x"88",  x"32",  x"0a",  x"0e",  x"21",  x"60",  x"da",  x"1a", -- 25F0
         x"23",  x"a6",  x"20",  x"62",  x"7b",  x"59",  x"ee",  x"4f", -- 25F8
         x"5d",  x"4f",  x"8a",  x"a4",  x"e4",  x"03",  x"21",  x"5c", -- 2600
         x"19",  x"b6",  x"7e",  x"00",  x"d6",  x"ab",  x"20",  x"04", -- 2608
         x"77",  x"0c",  x"15",  x"1c",  x"65",  x"cd",  x"a3",  x"50", -- 2610
         x"82",  x"c3",  x"f7",  x"d6",  x"e9",  x"ec",  x"01",  x"6c", -- 2618
         x"18",  x"a7",  x"b1",  x"00",  x"46",  x"68",  x"99",  x"e9", -- 2620
         x"92",  x"69",  x"10",  x"d1",  x"06",  x"75",  x"68",  x"21", -- 2628
         x"ba",  x"da",  x"3c",  x"ca",  x"88",  x"17",  x"49",  x"83", -- 2630
         x"a3",  x"99",  x"8e",  x"ce",  x"8e",  x"94",  x"fb",  x"b2", -- 2638
         x"c0",  x"b1",  x"f5",  x"84",  x"21",  x"be",  x"21",  x"66", -- 2640
         x"bd",  x"db",  x"15",  x"37",  x"f2",  x"a6",  x"09",  x"b0", -- 2648
         x"1a",  x"c8",  x"a4",  x"f5",  x"f4",  x"8a",  x"a3",  x"be", -- 2650
         x"39",  x"4c",  x"f1",  x"d4",  x"09",  x"1a",  x"c2",  x"da", -- 2658
         x"c3",  x"b5",  x"48",  x"3c",  x"49",  x"f3",  x"d0",  x"7f", -- 2660
         x"05",  x"ba",  x"d7",  x"00",  x"1e",  x"86",  x"64",  x"26", -- 2668
         x"99",  x"87",  x"58",  x"34",  x"88",  x"b6",  x"e0",  x"5d", -- 2670
         x"13",  x"a5",  x"86",  x"da",  x"18",  x"83",  x"4f",  x"4c", -- 2678
         x"76",  x"da",  x"b0",  x"b9",  x"df",  x"aa",  x"5b",  x"31", -- 2680
         x"52",  x"f3",  x"64",  x"49",  x"fc",  x"91",  x"6a",  x"a8", -- 2688
         x"c9",  x"fb",  x"50",  x"81",  x"da",  x"09",  x"db",  x"48", -- 2690
         x"01",  x"b1",  x"51",  x"6e",  x"59",  x"8c",  x"d5",  x"6f", -- 2698
         x"d4",  x"1b",  x"13",  x"db",  x"8a",  x"91",  x"9e",  x"80", -- 26A0
         x"c9",  x"09",  x"4a",  x"d7",  x"3b",  x"00",  x"78",  x"02", -- 26A8
         x"6e",  x"84",  x"7b",  x"fe",  x"c1",  x"2f",  x"00",  x"7c", -- 26B0
         x"74",  x"31",  x"9a",  x"7d",  x"84",  x"3d",  x"5a",  x"00", -- 26B8
         x"7d",  x"c8",  x"7f",  x"91",  x"7e",  x"e4",  x"bb",  x"4c", -- 26C0
         x"24",  x"7e",  x"6c",  x"f1",  x"4b",  x"7f",  x"e9",  x"01", -- 26C8
         x"49",  x"db",  x"28",  x"03",  x"e7",  x"d9",  x"37",  x"18", -- 26D0
         x"47",  x"db",  x"f1",  x"17",  x"e9",  x"e1",  x"a7",  x"1a", -- 26D8
         x"ae",  x"c0",  x"de",  x"b7",  x"88",  x"5c",  x"89",  x"0b", -- 26E0
         x"2f",  x"fe",  x"94",  x"9c",  x"00",  x"47",  x"d2",  x"48", -- 26E8
         x"c3",  x"d6",  x"07",  x"b1",  x"c3",  x"da",  x"06",  x"5d", -- 26F0
         x"d0",  x"00",  x"80",  x"b5",  x"6f",  x"eb",  x"18",  x"e0", -- 26F8
         x"30",  x"7b",  x"87",  x"00",  x"f6",  x"0d",  x"04",  x"57", -- 2700
         x"1e",  x"ef",  x"18",  x"d4",  x"a6",  x"c4",  x"36",  x"00", -- 2708
         x"9d",  x"c1",  x"89",  x"c6",  x"20",  x"f8",  x"b3",  x"90", -- 2710
         x"cd",  x"fe",  x"d2",  x"06",  x"cd",  x"09",  x"d2",  x"2a", -- 2718
         x"c4",  x"ab",  x"40",  x"5b",  x"56",  x"03",  x"af",  x"ed", -- 2720
         x"14",  x"52",  x"d1",  x"e3",  x"03",  x"14",  x"28",  x"58", -- 2728
         x"dd",  x"c8",  x"e4",  x"18",  x"dd",  x"47",  x"e1",  x"04", -- 2730
         x"12",  x"03",  x"13",  x"2b",  x"7d",  x"b4",  x"20",  x"f6", -- 2738
         x"0a",  x"58",  x"5f",  x"03",  x"57",  x"c1",  x"23",  x"38", -- 2740
         x"44",  x"2a",  x"2b",  x"54",  x"40",  x"0c",  x"ae",  x"c2", -- 2748
         x"1b",  x"7b",  x"b2",  x"1b",  x"a8",  x"33",  x"e8",  x"21", -- 2750
         x"f8",  x"dc",  x"38",  x"42",  x"20",  x"2d",  x"26",  x"02", -- 2758
         x"77",  x"dd",  x"e3",  x"2b",  x"d5",  x"4c",  x"c6",  x"50", -- 2760
         x"b8",  x"82",  x"90",  x"05",  x"e1",  x"42",  x"4b",  x"00", -- 2768
         x"03",  x"d1",  x"2b",  x"70",  x"2b",  x"71",  x"2b",  x"35", -- 2770
         x"16",  x"03",  x"20",  x"fc",  x"ab",  x"6a",  x"76",  x"f0", -- 2778
         x"25",  x"2f",  x"fd",  x"dd",  x"d9",  x"23",  x"85",  x"b0", -- 2780
         x"18",  x"29",  x"cd",  x"87",  x"03",  x"dc",  x"e5",  x"e2", -- 2788
         x"7b",  x"db",  x"eb",  x"7b",  x"e6",  x"d4",  x"5e",  x"e1", -- 2790
         x"5e",  x"e1",  x"00",  x"28",  x"c7",  x"cd",  x"1d",  x"de", -- 2798
         x"21",  x"3f",  x"dc",  x"01",  x"c3",  x"71",  x"c3",  x"42", -- 27A0
         x"41",  x"44",  x"00",  x"f9",  x"10",  x"28",  x"c6",  x"cd", -- 27A8
         x"20",  x"b0",  x"dc",  x"6c",  x"d7",  x"03",  x"1b",  x"1b", -- 27B0
         x"cc",  x"c6",  x"08",  x"39",  x"01",  x"d1",  x"ff",  x"41", -- 27B8
         x"09",  x"44",  x"63",  x"4d",  x"43",  x"6f",  x"3e",  x"0c", -- 27C0
         x"67",  x"e5",  x"33",  x"1e",  x"d2",  x"3e",  x"c3",  x"49", -- 27C8
         x"31",  x"91",  x"46",  x"2a",  x"21",  x"12",  x"d6",  x"28", -- 27D0
         x"c3",  x"8a",  x"c4",  x"39",  x"1e",  x"26",  x"ae",  x"04", -- 27D8
         x"cd",  x"ac",  x"dc",  x"69",  x"cc",  x"02",  x"c8",  x"3b", -- 27E0
         x"3e",  x"01",  x"32",  x"cc",  x"d6",  x"43",  x"06",  x"cf", -- 27E8
         x"05",  x"24",  x"94",  x"1d",  x"60",  x"69",  x"eb",  x"d1", -- 27F0
         x"28",  x"4e",  x"fa",  x"07",  x"09",  x"09",  x"23",  x"3a", -- 27F8
         x"ae",  x"8f",  x"00",  x"c9",  x"3e",  x"d4",  x"23",  x"01", -- 2800
         x"00",  x"3e",  x"d3",  x"f5",  x"3a",  x"5d",  x"03",  x"a7", -- 2808
         x"3e",  x"20",  x"00",  x"32",  x"05",  x"28",  x"04",  x"f1", -- 2810
         x"c6",  x"58",  x"04",  x"a8",  x"be",  x"d0",  x"81",  x"3a", -- 2818
         x"cd",  x"50",  x"f1",  x"2e",  x"09",  x"3f",  x"d3",  x"21", -- 2820
         x"54",  x"f7",  x"aa",  x"0d",  x"64",  x"2b",  x"99",  x"10", -- 2828
         x"00",  x"fb",  x"d5",  x"11",  x"82",  x"dc",  x"73",  x"23", -- 2830
         x"72",  x"12",  x"d1",  x"23",  x"f1",  x"9e",  x"6a",  x"01", -- 2838
         x"eb",  x"47",  x"00",  x"79",  x"fe",  x"09",  x"38",  x"04", -- 2840
         x"0d",  x"23",  x"18",  x"13",  x"f7",  x"ed",  x"b0",  x"b7", -- 2848
         x"0d",  x"af",  x"47",  x"86",  x"ac",  x"84",  x"dd",  x"20", -- 2850
         x"fa",  x"b9",  x"c1",  x"4f",  x"30",  x"01",  x"04",  x"81", -- 2858
         x"2a",  x"79",  x"43",  x"c9",  x"5a",  x"07",  x"03",  x"cb", -- 2860
         x"bc",  x"ca",  x"7d",  x"06",  x"00",  x"3e",  x"13",  x"20", -- 2868
         x"02",  x"c6",  x"08",  x"32",  x"08",  x"66",  x"03",  x"ec", -- 2870
         x"06",  x"f1",  x"c3",  x"d5",  x"dd",  x"19",  x"8d",  x"47", -- 2878
         x"cb",  x"c7",  x"19",  x"70",  x"12",  x"19",  x"09",  x"d4", -- 2880
         x"19",  x"c3",  x"d2",  x"51",  x"fd",  x"8a",  x"24",  x"d8", -- 2888
         x"25",  x"80",  x"51",  x"2a",  x"d4",  x"04",  x"11",  x"ff", -- 2890
         x"fb",  x"19",  x"f7",  x"48",  x"11",  x"4f",  x"cd",  x"b5", -- 2898
         x"28",  x"dd",  x"e1",  x"9a",  x"c1",  x"33",  x"8e",  x"11", -- 28A0
         x"43",  x"cf",  x"11",  x"f6",  x"df",  x"65",  x"4a",  x"db", -- 28A8
         x"09",  x"e2",  x"89",  x"dd",  x"c1",  x"49",  x"dd",  x"4a", -- 28B0
         x"87",  x"18",  x"e5",  x"e0",  x"88",  x"7e",  x"95",  x"8e", -- 28B8
         x"34",  x"81",  x"f2",  x"23",  x"85",  x"59",  x"f4",  x"1f", -- 28C0
         x"b1",  x"33",  x"c5",  x"1d",  x"9c",  x"3b",  x"11",  x"c1", -- 28C8
         x"79",  x"cd",  x"72",  x"78",  x"eb",  x"04",  x"99",  x"eb", -- 28D0
         x"70",  x"95",  x"28",  x"09",  x"b4",  x"56",  x"2b",  x"5e", -- 28D8
         x"b8",  x"86",  x"28",  x"f3",  x"1a",  x"10",  x"01",  x"13", -- 28E0
         x"0b",  x"18",  x"f5",  x"23",  x"e5",  x"1f",  x"26",  x"0d", -- 28E8
         x"1f",  x"e1",  x"1f",  x"c8",  x"cf",  x"1a",  x"48",  x"13", -- 28F0
         x"d1",  x"c9",  x"45",  x"3a",  x"a9",  x"b9",  x"75",  x"d4", -- 28F8
         x"94",  x"46",  x"99",  x"c3",  x"3e",  x"0c",  x"f5",  x"e0", -- 2900
         x"6c",  x"0f",  x"31",  x"5f",  x"7a",  x"78",  x"7b",  x"d8", -- 2908
         x"b2",  x"3c",  x"c3",  x"e5",  x"09",  x"0c",  x"0b",  x"b1", -- 2910
         x"b4",  x"80",  x"7a",  x"18",  x"06",  x"d5",  x"1e",  x"62", -- 2918
         x"80",  x"0c",  x"cb",  x"19",  x"89",  x"ef",  x"e5",  x"93", -- 2920
         x"81",  x"11",  x"42",  x"b1",  x"21",  x"06",  x"7a",  x"aa", -- 2928
         x"1a",  x"3e",  x"41",  x"dc",  x"15",  x"1c",  x"10",  x"f8", -- 2930
         x"c1",  x"91",  x"41",  x"3e",  x"f5",  x"df",  x"29",  x"2b", -- 2938
         x"64",  x"06",  x"8e",  x"d7",  x"47",  x"83",  x"5a",  x"d9", -- 2940
         x"0a",  x"23",  x"20",  x"31",  x"da",  x"c2",  x"30",  x"38", -- 2948
         x"79",  x"48",  x"e6",  x"f6",  x"12",  x"c1",  x"2d",  x"87", -- 2950
         x"fe",  x"04",  x"07",  x"01",  x"30",  x"16",  x"cb",  x"4e", -- 2958
         x"cb",  x"ce",  x"8e",  x"2a",  x"3c",  x"c2",  x"27",  x"e1", -- 2960
         x"c3",  x"89",  x"60",  x"cb",  x"5e",  x"cb",  x"de",  x"00", -- 2968
         x"18",  x"ee",  x"cb",  x"6e",  x"cb",  x"ee",  x"18",  x"e8", -- 2970
         x"92",  x"e2",  x"03",  x"d6",  x"39",  x"30",  x"39",  x"5a", -- 2978
         x"8b",  x"7a",  x"3a",  x"00",  x"10",  x"38",  x"14",  x"cb", -- 2980
         x"66",  x"cb",  x"e6",  x"96",  x"c9",  x"b2",  x"8a",  x"00", -- 2988
         x"c4",  x"cb",  x"56",  x"cb",  x"d6",  x"18",  x"f0",  x"cb", -- 2990
         x"06",  x"46",  x"cb",  x"c6",  x"18",  x"ea",  x"38",  x"24", -- 2998
         x"ea",  x"8b",  x"74",  x"2a",  x"95",  x"23",  x"c0",  x"00", -- 29A0
         x"01",  x"61",  x"03",  x"c5",  x"fc",  x"c9",  x"24",  x"d7", -- 29A8
         x"de",  x"ae",  x"2c",  x"fe",  x"22",  x"d6",  x"02",  x"b7", -- 29B0
         x"28",  x"1f",  x"f2",  x"a7",  x"de",  x"1d",  x"19",  x"9a", -- 29B8
         x"c7",  x"c1",  x"13",  x"fa",  x"10",  x"b7",  x"f2",  x"bb", -- 29C0
         x"9d",  x"70",  x"e4",  x"1e",  x"92",  x"d8",  x"b7",  x"ca", -- 29C8
         x"00",  x"3e",  x"20",  x"03",  x"18",  x"0c",  x"03",  x"02", -- 29D0
         x"90",  x"fd",  x"56",  x"fc",  x"11",  x"09",  x"e1",  x"d0", -- 29D8
         x"cb",  x"25",  x"2a",  x"a5",  x"05",  x"af",  x"02",  x"e1", -- 29E0
         x"81",  x"0a",  x"e5",  x"a4",  x"14",  x"c5",  x"8e",  x"55", -- 29E8
         x"ed",  x"9e",  x"48",  x"cd",  x"9c",  x"b7",  x"01",  x"0a", -- 29F0
         x"20",  x"05",  x"cd",  x"12",  x"df",  x"3c",  x"b1",  x"21", -- 29F8
         x"0f",  x"df",  x"c0",  x"40",  x"27",  x"df",  x"d8",  x"f8", -- 2A00
         x"dd",  x"df",  x"18",  x"03",  x"e7",  x"fe",  x"0d",  x"c0", -- 2A08
         x"3e",  x"09",  x"30",  x"09",  x"23",  x"7e",  x"49",  x"f6", -- 2A10
         x"d1",  x"c8",  x"20",  x"8a",  x"a1",  x"30",  x"44",  x"c3", -- 2A18
         x"d4",  x"fe",  x"88",  x"ba",  x"02",  x"a7",  x"a3",  x"2a", -- 2A20
         x"2f",  x"37",  x"c9",  x"b0",  x"a2",  x"28",  x"44",  x"c8", -- 2A28
         x"80",  x"28",  x"2a",  x"fe",  x"1f",  x"00",  x"28",  x"47", -- 2A30
         x"fe",  x"19",  x"ca",  x"c5",  x"df",  x"fe",  x"10",  x"18", -- 2A38
         x"ca",  x"cf",  x"04",  x"02",  x"ca",  x"db",  x"80",  x"04", -- 2A40
         x"1a",  x"28",  x"48",  x"fe",  x"0b",  x"c8",  x"a5",  x"5a", -- 2A48
         x"02",  x"01",  x"02",  x"f8",  x"11",  x"05",  x"3f",  x"4a", -- 2A50
         x"87",  x"c9",  x"77",  x"4f",  x"38",  x"9e",  x"14",  x"ab", -- 2A58
         x"03",  x"e5",  x"85",  x"28",  x"07",  x"7e",  x"84",  x"19", -- 2A60
         x"d2",  x"18",  x"a2",  x"54",  x"c6",  x"60",  x"15",  x"6e", -- 2A68
         x"18",  x"11",  x"df",  x"e5",  x"23",  x"9a",  x"9e",  x"fb", -- 2A70
         x"0d",  x"c6",  x"d1",  x"af",  x"cb",  x"28",  x"2d",  x"17", -- 2A78
         x"78",  x"20",  x"54",  x"f7",  x"6b",  x"0e",  x"b0",  x"6f", -- 2A80
         x"34",  x"26",  x"20",  x"0c",  x"15",  x"66",  x"11",  x"33", -- 2A88
         x"ca",  x"3b",  x"d1",  x"e2",  x"03",  x"03",  x"7e",  x"02", -- 2A90
         x"0b",  x"0c",  x"64",  x"28",  x"23",  x"4e",  x"c9",  x"e6", -- 2A98
         x"4a",  x"c1",  x"f1",  x"b2",  x"bc",  x"1e",  x"21",  x"18", -- 2AA0
         x"90",  x"cd",  x"c5",  x"58",  x"46",  x"09",  x"28",  x"05", -- 2AA8
         x"6f",  x"54",  x"f2",  x"e1",  x"da",  x"61",  x"10",  x"fe", -- 2AB0
         x"34",  x"c9",  x"1e",  x"07",  x"ff",  x"c3",  x"0e",  x"e0", -- 2AB8
         x"ff",  x"00",  x"80",  x"c3",  x"d2",  x"e0",  x"d2",  x"9c", -- 2AC0
         x"02",  x"10",  x"57",  x"e1",  x"11",  x"04",  x"00",  x"e6", -- 2AC8
         x"c9",  x"00",  x"4e",  x"4b",  x"45",  x"59",  x"24",  x"ca", -- 2AD0
         x"4f",  x"59",  x"00",  x"53",  x"54",  x"d3",  x"54",  x"52", -- 2AD8
         x"49",  x"4e",  x"47",  x"48",  x"24",  x"11",  x"53",  x"08", -- 2AE0
         x"d2",  x"45",  x"00",  x"4e",  x"55",  x"4d",  x"c4",  x"45", -- 2AE8
         x"4c",  x"45",  x"54",  x"00",  x"45",  x"d0",  x"41",  x"55", -- 2AF0
         x"53",  x"45",  x"c2",  x"45",  x"10",  x"45",  x"50",  x"d7", -- 2AF8
         x"1d",  x"44",  x"4f",  x"57",  x"03",  x"c2",  x"4f",  x"52", -- 2B00
         x"44",  x"45",  x"52",  x"36",  x"24",  x"17",  x"50",  x"07", -- 2B08
         x"c1",  x"12",  x"54",  x"d0",  x"53",  x"23",  x"cc",  x"19", -- 2B10
         x"04",  x"45",  x"c3",  x"49",  x"52",  x"43",  x"2e",  x"a1", -- 2B18
         x"a8",  x"15",  x"0b",  x"0f",  x"41",  x"42",  x"81",  x"3a", -- 2B20
         x"d3",  x"49",  x"5a",  x"45",  x"da",  x"21",  x"04",  x"4f", -- 2B28
         x"c8",  x"4f",  x"4d",  x"16",  x"c7",  x"82",  x"1b",  x"53", -- 2B30
         x"d3",  x"43",  x"41",  x"20",  x"88",  x"04",  x"52",  x"45", -- 2B38
         x"5b",  x"d0",  x"4f",  x"c0",  x"25",  x"d8",  x"50",  x"4f", -- 2B40
         x"53",  x"30",  x"a1",  x"d9",  x"04",  x"80",  x"19",  x"00", -- 2B48
         x"e4",  x"f5",  x"e4",  x"3c",  x"e4",  x"c1",  x"e4",  x"f8", -- 2B50
         x"88",  x"b6",  x"e5",  x"a7",  x"00",  x"e3",  x"34",  x"e4", -- 2B58
         x"b5",  x"e1",  x"79",  x"e1",  x"7d",  x"00",  x"e1",  x"7e", -- 2B60
         x"e1",  x"17",  x"e5",  x"d6",  x"a7",  x"d9",  x"00",  x"a7", -- 2B68
         x"dc",  x"a7",  x"4a",  x"ca",  x"df",  x"a7",  x"e2",  x"43", -- 2B70
         x"a7",  x"1a",  x"e8",  x"a7",  x"eb",  x"0b",  x"00",  x"ee", -- 2B78
         x"a7",  x"f1",  x"a7",  x"f4",  x"a7",  x"18",  x"f7",  x"a7", -- 2B80
         x"fa",  x"0b",  x"fd",  x"17",  x"a7",  x"78",  x"d6",  x"e5", -- 2B88
         x"2f",  x"6d",  x"e9",  x"11",  x"07",  x"f1",  x"00",  x"e5", -- 2B90
         x"fe",  x"16",  x"30",  x"62",  x"07",  x"4f",  x"b8",  x"f9", -- 2B98
         x"eb",  x"21",  x"00",  x"9e",  x"e0",  x"09",  x"4e",  x"23", -- 2BA0
         x"46",  x"c5",  x"eb",  x"55",  x"c3",  x"8b",  x"d5",  x"34", -- 2BA8
         x"ec",  x"c0",  x"fe",  x"e2",  x"d0",  x"fe",  x"e1",  x"46", -- 2BB0
         x"ca",  x"4e",  x"3a",  x"fd",  x"cb",  x"05",  x"20",  x"3f", -- 2BB8
         x"bd",  x"53",  x"06",  x"3a",  x"fd",  x"e6",  x"f5",  x"19", -- 2BC0
         x"15",  x"28",  x"0d",  x"ad",  x"8a",  x"cd",  x"69",  x"0a", -- 2BC8
         x"06",  x"3b",  x"28",  x"35",  x"18",  x"25",  x"0c",  x"b8", -- 2BD0
         x"7d",  x"0c",  x"13",  x"28",  x"cd",  x"d6",  x"d2",  x"0e", -- 2BD8
         x"e0",  x"20",  x"13",  x"1e",  x"73",  x"ab",  x"56",  x"cd", -- 2BE0
         x"b2",  x"13",  x"f1",  x"32",  x"35",  x"c1",  x"97",  x"20", -- 2BE8
         x"e2",  x"d3",  x"b8",  x"c3",  x"ab",  x"e0",  x"06",  x"83", -- 2BF0
         x"67",  x"c9",  x"20",  x"2a",  x"90",  x"01",  x"79",  x"d6", -- 2BF8
         x"3e",  x"38",  x"e8",  x"fe",  x"07",  x"8a",  x"c4",  x"84", -- 2C00
         x"69",  x"32",  x"38",  x"ed",  x"40",  x"3b",  x"30",  x"d9", -- 2C08
         x"02",  x"eb",  x"01",  x"96",  x"e0",  x"e1",  x"6f",  x"86", -- 2C10
         x"30",  x"66",  x"69",  x"e2",  x"b1",  x"34",  x"06",  x"01", -- 2C18
         x"18",  x"02",  x"f6",  x"af",  x"b3",  x"45",  x"21",  x"d4", -- 2C20
         x"ab",  x"04",  x"38",  x"6e",  x"af",  x"40",  x"30",  x"6a", -- 2C28
         x"3d",  x"4f",  x"f1",  x"98",  x"ad",  x"0b",  x"cb",  x"68", -- 2C30
         x"21",  x"01",  x"3d",  x"28",  x"17",  x"88",  x"04",  x"41", -- 2C38
         x"b7",  x"94",  x"c2",  x"28",  x"0a",  x"d7",  x"e6",  x"b0", -- 2C40
         x"66",  x"00",  x"32",  x"28",  x"00",  x"c9",  x"e6",  x"70", -- 2C48
         x"18",  x"00",  x"f4",  x"79",  x"d3",  x"88",  x"c9",  x"0e", -- 2C50
         x"1d",  x"cd",  x"33",  x"05",  x"00",  x"f7",  x"01",  x"28", -- 2C58
         x"2d",  x"cd",  x"f7",  x"e7",  x"42",  x"77",  x"03",  x"4a", -- 2C60
         x"00",  x"3c",  x"3c",  x"57",  x"fe",  x"2a",  x"30",  x"20", -- 2C68
         x"12",  x"f1",  x"5f",  x"f1",  x"09",  x"47",  x"8d",  x"ab", -- 2C70
         x"9f",  x"80",  x"f1",  x"4f",  x"3c",  x"b8",  x"30",  x"10", -- 2C78
         x"05",  x"7b",  x"3c",  x"ba",  x"30",  x"0b",  x"f8",  x"d8", -- 2C80
         x"f3",  x"3a",  x"19",  x"a2",  x"00",  x"29",  x"c3",  x"e6", -- 2C88
         x"e7",  x"c3",  x"4b",  x"e1",  x"01",  x"00",  x"0a",  x"00", -- 2C90
         x"c5",  x"50",  x"58",  x"28",  x"27",  x"fe",  x"1e",  x"2c", -- 2C98
         x"28",  x"09",  x"98",  x"1c",  x"86",  x"c9",  x"9f",  x"08", -- 2CA0
         x"d1",  x"28",  x"1a",  x"e2",  x"cc",  x"0a",  x"b9",  x"a4", -- 2CA8
         x"f1",  x"08",  x"9a",  x"14",  x"c2",  x"00",  x"44",  x"e1", -- 2CB0
         x"7a",  x"b3",  x"28",  x"d1",  x"eb",  x"e3",  x"28",  x"eb", -- 2CB8
         x"d5",  x"bc",  x"1c",  x"bb",  x"c4",  x"d1",  x"05",  x"6c", -- 2CC0
         x"95",  x"d1",  x"ac",  x"91",  x"00",  x"eb",  x"38",  x"ba", -- 2CC8
         x"d1",  x"f1",  x"c1",  x"d5",  x"f5",  x"24",  x"18",  x"0e", -- 2CD0
         x"e9",  x"2c",  x"f4",  x"eb",  x"ec",  x"30",  x"f9",  x"ff", -- 2CD8
         x"14",  x"e1",  x"38",  x"04",  x"e9",  x"d5",  x"5e",  x"23", -- 2CE0
         x"56",  x"33",  x"eb",  x"97",  x"4c",  x"07",  x"90",  x"07", -- 2CE8
         x"b6",  x"2b",  x"eb",  x"20",  x"b4",  x"05",  x"0e",  x"80", -- 2CF0
         x"dd",  x"85",  x"c3",  x"af",  x"b0",  x"c3",  x"e2",  x"af", -- 2CF8
         x"3c",  x"04",  x"30",  x"dd",  x"e5",  x"43",  x"c1",  x"3d", -- 2D00
         x"73",  x"2a",  x"f0",  x"26",  x"5e",  x"37",  x"23",  x"a9", -- 2D08
         x"06",  x"eb",  x"09",  x"eb",  x"87",  x"06",  x"eb",  x"3d", -- 2D10
         x"23",  x"38",  x"01",  x"94",  x"00",  x"c5",  x"3e",  x"02", -- 2D18
         x"32",  x"4e",  x"03",  x"2a",  x"5f",  x"01",  x"03",  x"2b", -- 2D20
         x"c5",  x"c5",  x"23",  x"c1",  x"c1",  x"f0",  x"57",  x"2b", -- 2D28
         x"03",  x"c8",  x"c5",  x"d5",  x"af",  x"52",  x"df",  x"49", -- 2D30
         x"a6",  x"04",  x"eb",  x"4f",  x"3a",  x"1e",  x"b7",  x"17", -- 2D38
         x"79",  x"28",  x"5f",  x"b0",  x"0b",  x"20",  x"ee",  x"e5", -- 2D40
         x"bf",  x"33",  x"1e",  x"10",  x"24",  x"b5",  x"4b",  x"7e", -- 2D48
         x"02",  x"0e",  x"4d",  x"8f",  x"c2",  x"ed",  x"a0",  x"01", -- 2D50
         x"8b",  x"84",  x"f1",  x"a4",  x"18",  x"b3",  x"46",  x"eb", -- 2D58
         x"13",  x"98",  x"e6",  x"d5",  x"92",  x"42",  x"e1",  x"67", -- 2D60
         x"6d",  x"c5",  x"f9",  x"de",  x"98",  x"e5",  x"00",  x"c5", -- 2D68
         x"af",  x"06",  x"98",  x"cd",  x"ae",  x"d6",  x"cd",  x"2b", -- 2D70
         x"34",  x"d8",  x"0d",  x"ac",  x"08",  x"eb",  x"2b",  x"4f", -- 2D78
         x"aa",  x"23",  x"91",  x"1b",  x"e5",  x"81",  x"0e",  x"54", -- 2D80
         x"5d",  x"13",  x"9b",  x"d3",  x"1b",  x"2b",  x"b5",  x"c4", -- 2D88
         x"e1",  x"40",  x"c1",  x"00",  x"18",  x"e3",  x"fe",  x"88", -- 2D90
         x"28",  x"19",  x"fe",  x"8c",  x"00",  x"28",  x"15",  x"fe", -- 2D98
         x"8b",  x"28",  x"11",  x"fe",  x"d4",  x"88",  x"ab",  x"fe", -- 2DA0
         x"da",  x"90",  x"ae",  x"fe",  x"d3",  x"b0",  x"d3",  x"fe", -- 2DA8
         x"a9",  x"1b",  x"c2",  x"b2",  x"e2",  x"d2",  x"71",  x"c6", -- 2DB0
         x"cc",  x"18",  x"e1",  x"c9",  x"cb",  x"7e",  x"c6",  x"28", -- 2DB8
         x"f1",  x"9a",  x"6c",  x"eb",  x"0d",  x"23",  x"1d",  x"71", -- 2DC0
         x"23",  x"70",  x"d7",  x"57",  x"1d",  x"78",  x"77",  x"18", -- 2DC8
         x"f6",  x"03",  x"c1",  x"62",  x"6b",  x"1b",  x"1a",  x"20", -- 2DD0
         x"01",  x"10",  x"fe",  x"3a",  x"30",  x"0c",  x"a7",  x"d0", -- 2DD8
         x"2b",  x"e3",  x"f5",  x"8a",  x"c6",  x"87",  x"26",  x"d1", -- 2DE0
         x"ec",  x"1c",  x"6f",  x"67",  x"00",  x"72",  x"11",  x"71", -- 2DE8
         x"3e",  x"0d",  x"a6",  x"d8",  x"d1",  x"ed",  x"b3",  x"66", -- 2DF0
         x"e3",  x"14",  x"07",  x"49",  x"29",  x"d5",  x"5f",  x"93", -- 2DF8
         x"51",  x"84",  x"18",  x"9f",  x"ec",  x"e0",  x"20",  x"11", -- 2E00
         x"cd",  x"70",  x"f3",  x"a9",  x"fb",  x"cc",  x"89",  x"06", -- 2E08
         x"07",  x"fe",  x"1e",  x"20",  x"f3",  x"c2",  x"65",  x"ea", -- 2E10
         x"04",  x"5e",  x"c9",  x"94",  x"a4",  x"fc",  x"93",  x"d8", -- 2E18
         x"00",  x"dd",  x"21",  x"0b",  x"e4",  x"3e",  x"05",  x"0e", -- 2E20
         x"03",  x"8d",  x"06",  x"0a",  x"dd",  x"86",  x"00",  x"fc", -- 2E28
         x"a5",  x"0d",  x"ff",  x"ca",  x"3d",  x"85",  x"2c",  x"9c", -- 2E30
         x"86",  x"7e",  x"eb",  x"28",  x"1b",  x"6e",  x"6a",  x"39", -- 2E38
         x"08",  x"35",  x"8c",  x"bb",  x"80",  x"3d",  x"08",  x"d1", -- 2E40
         x"c1",  x"f1",  x"18",  x"cf",  x"cc",  x"3e",  x"07",  x"e1", -- 2E48
         x"f6",  x"c3",  x"f0",  x"97",  x"c3",  x"c1",  x"53",  x"49", -- 2E50
         x"43",  x"20",  x"00",  x"64",  x"e7",  x"8c",  x"3a",  x"c0", -- 2E58
         x"57",  x"0c",  x"e9",  x"9d",  x"e5",  x"33",  x"aa",  x"0f", -- 2E60
         x"a5",  x"9c",  x"cd",  x"a7",  x"60",  x"2b",  x"2a",  x"c2", -- 2E68
         x"03",  x"19",  x"77",  x"c3",  x"a9",  x"9f",  x"66",  x"0d", -- 2E70
         x"cb",  x"01",  x"0e",  x"02",  x"1e",  x"07",  x"80",  x"59", -- 2E78
         x"7e",  x"2a",  x"cc",  x"81",  x"a6",  x"f8",  x"08",  x"8e", -- 2E80
         x"e4",  x"03",  x"db",  x"c8",  x"88",  x"da",  x"44",  x"e5", -- 2E88
         x"e0",  x"f9",  x"4f",  x"af",  x"08",  x"b9",  x"28",  x"0c", -- 2E90
         x"b8",  x"69",  x"79",  x"05",  x"90",  x"a5",  x"81",  x"38", -- 2E98
         x"44",  x"29",  x"8b",  x"47",  x"54",  x"0e",  x"aa",  x"e1", -- 2EA0
         x"a6",  x"6b",  x"f6",  x"26",  x"7e",  x"d1",  x"81",  x"42", -- 2EA8
         x"7c",  x"02",  x"6f",  x"24",  x"25",  x"80",  x"64",  x"28", -- 2EB0
         x"40",  x"f2",  x"15",  x"d2",  x"c1",  x"e1",  x"ce",  x"51", -- 2EB8
         x"03",  x"5e",  x"02",  x"d3",  x"5a",  x"80",  x"1e",  x"1c", -- 2EC0
         x"c3",  x"56",  x"c3",  x"fc",  x"c8",  x"84",  x"77",  x"30", -- 2EC8
         x"d3",  x"23",  x"cf",  x"ec",  x"9b",  x"52",  x"ba",  x"02", -- 2ED0
         x"2b",  x"0d",  x"c5",  x"0c",  x"13",  x"48",  x"10",  x"11", -- 2ED8
         x"23",  x"0d",  x"50",  x"1a",  x"be",  x"28",  x"d1",  x"2d", -- 2EE0
         x"18",  x"2c",  x"e1",  x"36",  x"29",  x"31",  x"4a",  x"dc", -- 2EE8
         x"91",  x"a7",  x"dd",  x"08",  x"7d",  x"18",  x"2a",  x"84", -- 2EF0
         x"e2",  x"80",  x"2a",  x"89",  x"ab",  x"bc",  x"63",  x"88", -- 2EF8
         x"aa",  x"c9",  x"91",  x"4f",  x"03",  x"6d",  x"47",  x"ef", -- 2F00
         x"37",  x"df",  x"58",  x"35",  x"b8",  x"84",  x"3d",  x"20", -- 2F08
         x"f9",  x"af",  x"35",  x"11",  x"68",  x"f3",  x"9b",  x"18", -- 2F10
         x"48",  x"23",  x"dc",  x"18",  x"45",  x"f6",  x"8f",  x"66", -- 2F18
         x"68",  x"0d",  x"cd",  x"24",  x"d4",  x"12",  x"a7",  x"28", -- 2F20
         x"45",  x"93",  x"04",  x"30",  x"41",  x"0e",  x"06",  x"d0", -- 2F28
         x"61",  x"38",  x"3a",  x"8a",  x"70",  x"28",  x"01",  x"48", -- 2F30
         x"0c",  x"79",  x"c3",  x"c0",  x"d0",  x"97",  x"40",  x"cb", -- 2F38
         x"4f",  x"cb",  x"cf",  x"c4",  x"97",  x"63",  x"20",  x"83", -- 2F40
         x"11",  x"e9",  x"dd",  x"e2",  x"9b",  x"60",  x"fd",  x"7b", -- 2F48
         x"d9",  x"65",  x"d9",  x"c6",  x"47",  x"78",  x"fb",  x"db", -- 2F50
         x"e4",  x"02",  x"79",  x"fe",  x"28",  x"38",  x"03",  x"d2", -- 2F58
         x"d0",  x"2e",  x"00",  x"24",  x"65",  x"55",  x"e2",  x"44", -- 2F60
         x"04",  x"ae",  x"03",  x"0b",  x"19",  x"10",  x"fd",  x"59", -- 2F68
         x"ea",  x"42",  x"ec",  x"19",  x"df",  x"69",  x"9a",  x"ba", -- 2F70
         x"85",  x"98",  x"c6",  x"fe",  x"d5",  x"05",  x"38",  x"09", -- 2F78
         x"3a",  x"fc",  x"03",  x"6c",  x"cc",  x"b1",  x"06",  x"e0", -- 2F80
         x"e4",  x"1a",  x"3a",  x"55",  x"ae",  x"bd",  x"d4",  x"b8", -- 2F88
         x"34",  x"e0",  x"f5",  x"8a",  x"d1",  x"d8",  x"9f",  x"2a", -- 2F90
         x"e5",  x"00",  x"03",  x"34",  x"cd",  x"fe",  x"d2",  x"cd", -- 2F98
         x"ee",  x"d6",  x"05",  x"e1",  x"dd",  x"e1",  x"fd",  x"e1", -- 2FA0
         x"f5",  x"e0",  x"57",  x"1c",  x"1d",  x"01",  x"28",  x"13", -- 2FA8
         x"0a",  x"cd",  x"bf",  x"e5",  x"30",  x"e7",  x"f0",  x"77", -- 2FB0
         x"00",  x"fd",  x"4c",  x"72",  x"e0",  x"23",  x"1e",  x"fd", -- 2FB8
         x"23",  x"03",  x"96",  x"52",  x"87",  x"b0",  x"02",  x"f1", -- 2FC0
         x"8c",  x"eb",  x"03",  x"fd",  x"e5",  x"dd",  x"e5",  x"18", -- 2FC8
         x"a7",  x"04",  x"01",  x"e1",  x"d5",  x"11",  x"c0",  x"ef", -- 2FD0
         x"8b",  x"28",  x"d1",  x"92",  x"b0",  x"bd",  x"f4",  x"ca", -- 2FD8
         x"42",  x"5f",  x"c4",  x"bd",  x"44",  x"e1",  x"c0",  x"ff", -- 2FE0
         x"55",  x"90",  x"85",  x"d2",  x"4d",  x"b8",  x"d4",  x"82", -- 2FE8
         x"40",  x"38",  x"c4",  x"30",  x"f5",  x"c1",  x"c3",  x"00", -- 2FF0
         x"50",  x"c4",  x"47",  x"e5",  x"2a",  x"b0",  x"e0",  x"3e", -- 2FF8
         x"f8",  x"aa",  x"78",  x"e1",  x"2e",  x"c8",  x"c3",  x"de", -- 3000
         x"09",  x"ff",  x"cb",  x"6b",  x"c2",  x"eb",  x"94",  x"22", -- 3008
         x"62",  x"92",  x"c0",  x"21",  x"1e",  x"e6",  x"e5",  x"7b", -- 3010
         x"c1",  x"eb",  x"17",  x"ae",  x"a8",  x"21",  x"0c",  x"42", -- 3018
         x"e6",  x"09",  x"7e",  x"a6",  x"84",  x"6f",  x"e9",  x"c1", -- 3020
         x"53",  x"0a",  x"00",  x"0d",  x"56",  x"65",  x"72",  x"69", -- 3028
         x"66",  x"79",  x"20",  x"d0",  x"81",  x"59",  x"29",  x"00", -- 3030
         x"2f",  x"4e",  x"29",  x"3f",  x"3a",  x"00",  x"0a",  x"52", -- 3038
         x"00",  x"65",  x"77",  x"69",  x"6e",  x"64",  x"20",  x"3c", -- 3040
         x"3d",  x"40",  x"3d",  x"1d",  x"00",  x"52",  x"e6",  x"72", -- 3048
         x"e6",  x"01",  x"34",  x"e7",  x"85",  x"e6",  x"82",  x"dc", -- 3050
         x"6e",  x"03",  x"91",  x"01",  x"cb",  x"7b",  x"af",  x"31", -- 3058
         x"0e",  x"0b",  x"ce",  x"28",  x"b7",  x"b8",  x"8a",  x"cb", -- 3060
         x"bb",  x"30",  x"18",  x"0a",  x"a0",  x"c3",  x"0b",  x"0e", -- 3068
         x"01",  x"04",  x"19",  x"57",  x"b8",  x"32",  x"05",  x"f4", -- 3070
         x"a0",  x"bd",  x"d5",  x"5a",  x"c4",  x"0c",  x"d1",  x"1b", -- 3078
         x"c9",  x"00",  x"16",  x"0a",  x"18",  x"f1",  x"16",  x"0d", -- 3080
         x"18",  x"ed",  x"00",  x"d5",  x"cb",  x"5b",  x"28",  x"22", -- 3088
         x"d5",  x"0e",  x"0f",  x"c7",  x"16",  x"16",  x"9b",  x"d0", -- 3090
         x"4e",  x"01",  x"0b",  x"00",  x"44",  x"2a",  x"92",  x"23", -- 3098
         x"b8",  x"9a",  x"32",  x"75",  x"0b",  x"00",  x"11",  x"80", -- 30A0
         x"00",  x"ac",  x"40",  x"21",  x"6e",  x"00",  x"36",  x"25", -- 30A8
         x"0b",  x"21",  x"0a",  x"3a",  x"07",  x"9f",  x"18",  x"09", -- 30B0
         x"6d",  x"72",  x"b1",  x"08",  x"15",  x"cb",  x"73",  x"d3", -- 30B8
         x"60",  x"0f",  x"fe",  x"80",  x"c2",  x"14",  x"7d",  x"e7", -- 30C0
         x"3a",  x"28",  x"e3",  x"87",  x"20",  x"1a",  x"21",  x"26", -- 30C8
         x"47",  x"56",  x"43",  x"04",  x"23",  x"10",  x"f9",  x"21", -- 30D0
         x"d9",  x"55",  x"2b",  x"79",  x"9b",  x"23",  x"42",  x"a6", -- 30D8
         x"cc",  x"19",  x"26",  x"22",  x"1b",  x"0c",  x"15",  x"62", -- 30E0
         x"33",  x"af",  x"3b",  x"66",  x"88",  x"40",  x"28",  x"74", -- 30E8
         x"90",  x"0c",  x"5a",  x"62",  x"21",  x"e6",  x"cd",  x"56", -- 30F0
         x"62",  x"02",  x"10",  x"ea",  x"d0",  x"02",  x"81",  x"e6", -- 30F8
         x"fe",  x"07",  x"4e",  x"28",  x"66",  x"11",  x"34",  x"12", -- 3100
         x"1c",  x"0f",  x"14",  x"3a",  x"6b",  x"51",  x"26",  x"6c", -- 3108
         x"48",  x"00",  x"c3",  x"83",  x"21",  x"e7",  x"c1",  x"55", -- 3110
         x"18",  x"49",  x"d5",  x"79",  x"88",  x"44",  x"b2",  x"c6", -- 3118
         x"1b",  x"1f",  x"59",  x"a0",  x"19",  x"98",  x"18",  x"cd", -- 3120
         x"22",  x"9d",  x"e7",  x"a4",  x"08",  x"8b",  x"00",  x"56", -- 3128
         x"d5",  x"a9",  x"d1",  x"0c",  x"18",  x"1c",  x"ab",  x"1e", -- 3130
         x"2a",  x"d1",  x"13",  x"ad",  x"36",  x"a6",  x"23",  x"20", -- 3138
         x"10",  x"27",  x"36",  x"7c",  x"9d",  x"58",  x"bc",  x"89", -- 3140
         x"4a",  x"1d",  x"83",  x"08",  x"cb",  x"9b",  x"c9",  x"9a", -- 3148
         x"e9",  x"14",  x"14",  x"82",  x"d0",  x"cd",  x"67",  x"7e", -- 3150
         x"a9",  x"eb",  x"ed",  x"1c",  x"09",  x"20",  x"f5",  x"c3", -- 3158
         x"ca",  x"30",  x"19",  x"06",  x"0b",  x"8e",  x"cc",  x"a5", -- 3160
         x"90",  x"04",  x"0e",  x"0c",  x"09",  x"0e",  x"11",  x"2a", -- 3168
         x"8a",  x"00",  x"d3",  x"00",  x"1b",  x"20",  x"04",  x"2b", -- 3170
         x"10",  x"f8",  x"c9",  x"d6",  x"00",  x"04",  x"be",  x"20", -- 3178
         x"d8",  x"3e",  x"ff",  x"32",  x"5e",  x"a1",  x"99",  x"f0", -- 3180
         x"cf",  x"fe",  x"3f",  x"00",  x"16",  x"e1",  x"09",  x"3d", -- 3188
         x"c5",  x"00",  x"43",  x"3b",  x"00",  x"51",  x"14",  x"1c", -- 3190
         x"2f",  x"0e",  x"12",  x"ba",  x"8a",  x"c8",  x"d5",  x"d6", -- 3198
         x"a9",  x"8f",  x"c9",  x"00",  x"ff",  x"f8",  x"00",  x"c3", -- 31A0
         x"03",  x"80",  x"f3",  x"3e",  x"20",  x"21",  x"00",  x"00", -- 31A8
         x"e8",  x"11",  x"01",  x"e8",  x"01",  x"ff",  x"07",  x"77", -- 31B0
         x"00",  x"ed",  x"b0",  x"3e",  x"03",  x"d3",  x"8a",  x"3e", -- 31B8
         x"cf",  x"91",  x"03",  x"af",  x"02",  x"d3",  x"88",  x"18", -- 31C0
         x"00",  x"ec",  x"3e",  x"58",  x"77",  x"34",  x"7e",  x"fe", -- 31C8
         x"01",  x"59",  x"c2",  x"35",  x"81",  x"31",  x"bf",  x"ef", -- 31D0
         x"0f",  x"80",  x"11",  x"11",  x"81",  x"cd",  x"03",  x"00", -- 31D8
         x"81",  x"16",  x"00",  x"cd",  x"4b",  x"80",  x"cd",  x"5b", -- 31E0
         x"1c",  x"80",  x"16",  x"ff",  x"07",  x"88",  x"c3",  x"27", -- 31E8
         x"81",  x"1b",  x"00",  x"01",  x"00",  x"00",  x"40",  x"72", -- 31F0
         x"23",  x"0d",  x"79",  x"b7",  x"20",  x"0e",  x"f9",  x"10", -- 31F8
         x"f7",  x"c9",  x"0f",  x"40",  x"7e",  x"5f",  x"cd",  x"73", -- 3200
         x"80",  x"ba",  x"1c",  x"c2",  x"f6",  x"80",  x"17",  x"00", -- 3208
         x"f1",  x"10",  x"ef",  x"c9",  x"c5",  x"f5",  x"7c",  x"01", -- 3210
         x"e5",  x"21",  x"0a",  x"ec",  x"f5",  x"cb",  x"3f",  x"01", -- 3218
         x"c8",  x"fe",  x"0a",  x"38",  x"00",  x"02",  x"c6",  x"07", -- 3220
         x"c6",  x"30",  x"cd",  x"0b",  x"81",  x"1e",  x"f1",  x"e6", -- 3228
         x"0f",  x"0d",  x"40",  x"7d",  x"fe",  x"0e",  x"28",  x"08", -- 3230
         x"00",  x"e1",  x"e5",  x"7d",  x"21",  x"0c",  x"ec",  x"18", -- 3238
         x"d1",  x"27",  x"23",  x"7a",  x"3d",  x"0a",  x"16",  x"18", -- 3240
         x"02",  x"18",  x"01",  x"04",  x"3e",  x"46",  x"18",  x"f4", -- 3248
         x"23",  x"7b",  x"42",  x"f1",  x"3d",  x"7b",  x"42",  x"20", -- 3250
         x"22",  x"06",  x"08",  x"cb",  x"27",  x"10",  x"38",  x"0b", -- 3258
         x"0e",  x"0c",  x"0e",  x"81",  x"10",  x"00",  x"f5",  x"e1", -- 3260
         x"f1",  x"c1",  x"c9",  x"0e",  x"31",  x"18",  x"01",  x"f3", -- 3268
         x"21",  x"1f",  x"ec",  x"d5",  x"11",  x"20",  x"c7",  x"1a", -- 3270
         x"d1",  x"00",  x"18",  x"5f",  x"1a",  x"b7",  x"c8",  x"77", -- 3278
         x"23",  x"13",  x"22",  x"18",  x"f8",  x"04",  x"c9",  x"71", -- 3280
         x"02",  x"00",  x"52",  x"41",  x"4d",  x"54",  x"45",  x"53", -- 3288
         x"54",  x"00",  x"c0",  x"07",  x"20",  x"4f",  x"4b",  x"00", -- 3290
         x"01",  x"46",  x"45",  x"48",  x"4c",  x"45",  x"52",  x"00", -- 3298
         x"30",  x"86",  x"11",  x"19",  x"2f",  x"92",  x"3e",  x"40", -- 32A0
         x"94",  x"22",  x"76",  x"fc",  x"22",  x"18",  x"02",  x"f8", -- 32A8
         x"8f",  x"ef",  x"68",  x"ee",  x"ec",  x"ba",  x"20",  x"70", -- 32B0
         x"0d",  x"12",  x"f5",  x"01",  x"10",  x"f3",  x"ba",  x"28", -- 32B8
         x"d9",  x"18",  x"ce",  x"b7",  x"14",  x"83",  x"62",  x"20", -- 32C0
         x"85",  x"38",  x"08",  x"10",  x"fa",  x"18",  x"c8",  x"07", -- 32C8
         x"30",  x"03",  x"9a",  x"07",  x"76",  x"47",  x"18",  x"31", -- 32D0
         x"08",  x"af",  x"04",  x"03",  x"27",  x"09",  x"76",  x"08", -- 32D8
         x"d9",  x"fb",  x"1a",  x"ff",  x"34",  x"fb",  x"02",  x"10", -- 32E0
         x"f9",  x"d9",  x"08",  x"b7",  x"28",  x"ef",  x"20",  x"e5", -- 32E8
         x"ff",  x"28",  x"43",  x"0f",  x"29",  x"2d",  x"55",  x"5a", -- 32F0
         x"00",  x"ff",  x"f8",  x"00",  x"00",  x"00",  x"00",  x"00", -- 32F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3300
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3308
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3310
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3318
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3320
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3328
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3330
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3338
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3340
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3348
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3350
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3358
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3360
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3368
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3370
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3378
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3380
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3388
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3390
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3398
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 33A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 33A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 33B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 33B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 33C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 33C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 33D0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 33D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 33E0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 33E8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 33F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 33F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3400
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3408
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3410
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3418
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3420
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3428
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3430
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3438
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3440
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3448
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3450
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3458
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3460
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3468
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3470
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3478
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3480
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3488
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3490
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3498
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 34A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 34A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 34B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 34B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 34C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 34C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 34D0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 34D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 34E0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 34E8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 34F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 34F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3500
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3508
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3510
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3518
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3520
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3528
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3530
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3538
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3540
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3548
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3550
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3558
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3560
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3568
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3570
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3578
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3580
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3588
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3590
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3598
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 35A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 35A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 35B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 35B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 35C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 35C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 35D0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 35D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 35E0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 35E8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 35F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 35F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3600
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3608
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3610
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3618
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3620
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3628
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3630
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3638
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3640
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3648
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3650
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3658
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3660
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3668
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3670
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3678
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3680
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3688
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3690
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3698
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 36A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 36A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 36B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 36B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 36C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 36C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 36D0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 36D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 36E0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 36E8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 36F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 36F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3700
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3708
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3710
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3718
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3720
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3728
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3730
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3738
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3740
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3748
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3750
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3758
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3760
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3768
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3770
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3778
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3780
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3788
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3790
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3798
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 37A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 37A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 37B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 37B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 37C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 37C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 37D0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 37D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 37E0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 37E8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 37F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 37F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3800
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3808
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3810
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3818
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3820
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3828
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3830
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3838
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3840
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3848
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3850
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3858
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3860
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3868
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3870
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3878
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3880
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3888
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3890
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3898
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 38A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 38A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 38B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 38B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 38C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 38C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 38D0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 38D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 38E0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 38E8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 38F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 38F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3900
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3908
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3910
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3918
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3920
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3928
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3930
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3938
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3940
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3948
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3950
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3958
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3960
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3968
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3970
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3978
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3980
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3988
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3990
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3998
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 39A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 39A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 39B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 39B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 39C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 39C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 39D0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 39D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 39E0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 39E8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 39F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 39F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A10
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A28
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A30
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A38
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A40
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A48
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A50
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A58
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A60
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A68
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A70
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A78
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A80
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A88
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A90
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3AA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3AA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3AB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3AB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3AC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3AC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3AD0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3AD8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3AE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3AE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3AF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3AF8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B10
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B28
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B30
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B38
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B40
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B48
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B50
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B58
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B60
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B68
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B70
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B78
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B80
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B88
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B90
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3BA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3BA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3BB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3BB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3BC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3BC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3BD0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3BD8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3BE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3BE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3BF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3BF8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C10
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C28
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C30
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C38
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C40
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C48
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C50
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C58
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C60
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C68
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C70
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C78
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C80
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C88
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C90
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3CA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3CA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3CB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3CB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3CC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3CC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3CD0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3CD8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3CE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3CE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3CF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3CF8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D10
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D28
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D30
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D38
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D40
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D48
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D50
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D58
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D60
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D68
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D70
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D78
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D80
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D88
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D90
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3DA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3DA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3DB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3DB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3DC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3DC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3DD0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3DD8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3DE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3DE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3DF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3DF8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E10
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E28
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E30
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E38
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E40
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E48
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E50
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E58
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E60
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E68
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E70
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E78
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E80
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E88
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E90
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3EA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3EA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3EB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3EB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3EC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3EC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3ED0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3ED8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3EE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3EE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3EF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3EF8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F10
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F28
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F30
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F38
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F40
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F48
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F50
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F58
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F60
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F68
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F70
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F78
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F80
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F88
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F90
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3FA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3FA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3FB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3FB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3FC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3FC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3FD0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3FD8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3FE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3FE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3FF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00"  -- 3FF8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
