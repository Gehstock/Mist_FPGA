library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity pooyan_sound_prog is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of pooyan_sound_prog is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"21",X"00",X"30",X"06",X"00",X"C3",X"AC",X"00",X"32",X"00",X"50",X"3A",X"00",X"40",X"C9",X"FF",
		X"32",X"00",X"70",X"3A",X"00",X"60",X"C9",X"FF",X"78",X"CF",X"79",X"32",X"00",X"40",X"C9",X"FF",
		X"78",X"D7",X"79",X"32",X"00",X"60",X"C9",X"FF",X"87",X"85",X"6F",X"7C",X"CE",X"00",X"67",X"7E",
		X"23",X"66",X"6F",X"E9",X"FF",X"FF",X"FF",X"FF",X"D9",X"08",X"CD",X"40",X"00",X"08",X"D9",X"C9",
		X"3E",X"0E",X"CF",X"B7",X"28",X"40",X"57",X"E6",X"7F",X"FE",X"2B",X"D0",X"CB",X"7A",X"28",X"03",
		X"C3",X"A3",X"00",X"57",X"CD",X"91",X"00",X"28",X"04",X"23",X"36",X"00",X"C9",X"AF",X"CD",X"91",
		X"00",X"28",X"05",X"72",X"23",X"36",X"00",X"C9",X"21",X"00",X"30",X"1E",X"06",X"7E",X"1D",X"28",
		X"08",X"2C",X"2C",X"BE",X"38",X"F8",X"C3",X"6D",X"00",X"5F",X"7A",X"BB",X"D8",X"7B",X"CD",X"91",
		X"00",X"72",X"2C",X"36",X"00",X"C9",X"21",X"00",X"30",X"06",X"0C",X"AF",X"77",X"23",X"10",X"FC",
		X"C9",X"21",X"00",X"30",X"06",X"06",X"0E",X"07",X"BE",X"28",X"05",X"23",X"23",X"10",X"F9",X"41",
		X"79",X"90",X"C9",X"CD",X"91",X"00",X"C8",X"AF",X"77",X"23",X"77",X"C9",X"70",X"23",X"7C",X"FE",
		X"34",X"20",X"F9",X"F9",X"ED",X"56",X"21",X"00",X"80",X"22",X"0C",X"30",X"77",X"16",X"06",X"7A",
		X"CD",X"B0",X"01",X"15",X"20",X"F9",X"01",X"38",X"07",X"DF",X"E7",X"FB",X"3E",X"0F",X"CF",X"E6",
		X"80",X"20",X"F9",X"3E",X"0F",X"CF",X"E6",X"80",X"28",X"F9",X"F3",X"3E",X"01",X"32",X"0E",X"30",
		X"3A",X"01",X"30",X"B7",X"3A",X"00",X"30",X"CA",X"EF",X"00",X"CD",X"93",X"01",X"18",X"03",X"CD",
		X"7D",X"01",X"FB",X"00",X"00",X"F3",X"3E",X"02",X"32",X"0E",X"30",X"3A",X"03",X"30",X"B7",X"3A",
		X"02",X"30",X"CA",X"0A",X"01",X"CD",X"93",X"01",X"18",X"03",X"CD",X"7D",X"01",X"FB",X"00",X"00",
		X"F3",X"3E",X"03",X"32",X"0E",X"30",X"3A",X"05",X"30",X"B7",X"3A",X"04",X"30",X"CA",X"25",X"01",
		X"CD",X"93",X"01",X"18",X"03",X"CD",X"7D",X"01",X"FB",X"00",X"00",X"F3",X"3E",X"04",X"32",X"0E",
		X"30",X"3A",X"07",X"30",X"B7",X"3A",X"06",X"30",X"CA",X"40",X"01",X"CD",X"93",X"01",X"18",X"03",
		X"CD",X"7D",X"01",X"FB",X"00",X"00",X"F3",X"3E",X"05",X"32",X"0E",X"30",X"3A",X"09",X"30",X"B7",
		X"3A",X"08",X"30",X"CA",X"5B",X"01",X"CD",X"93",X"01",X"18",X"03",X"CD",X"7D",X"01",X"FB",X"00",
		X"00",X"F3",X"3E",X"06",X"32",X"0E",X"30",X"3A",X"0B",X"30",X"B7",X"3A",X"0A",X"30",X"CA",X"77",
		X"01",X"CD",X"93",X"01",X"C3",X"CB",X"00",X"CD",X"7D",X"01",X"C3",X"CB",X"00",X"21",X"D3",X"09",
		X"EF",X"B7",X"20",X"17",X"21",X"01",X"30",X"3A",X"0E",X"30",X"3D",X"87",X"5F",X"16",X"00",X"19",
		X"36",X"01",X"C9",X"B7",X"C8",X"21",X"29",X"0A",X"EF",X"B7",X"C8",X"21",X"00",X"30",X"3A",X"0E",
		X"30",X"3D",X"87",X"4F",X"06",X"00",X"09",X"70",X"23",X"70",X"C9",X"0E",X"00",X"3A",X"0E",X"30",
		X"FE",X"04",X"30",X"06",X"C6",X"07",X"47",X"C3",X"18",X"00",X"C6",X"04",X"47",X"C3",X"20",X"00",
		X"3A",X"0E",X"30",X"FE",X"04",X"30",X"0A",X"3D",X"87",X"47",X"4D",X"DF",X"4C",X"04",X"C3",X"18",
		X"00",X"D6",X"04",X"87",X"47",X"4D",X"E7",X"4C",X"04",X"C3",X"20",X"00",X"01",X"FC",X"FF",X"21",
		X"00",X"00",X"1F",X"CB",X"15",X"1F",X"CB",X"15",X"3A",X"0E",X"30",X"C6",X"02",X"FE",X"06",X"38",
		X"04",X"D6",X"06",X"28",X"0A",X"87",X"29",X"37",X"CB",X"11",X"CB",X"10",X"3D",X"20",X"F7",X"EB",
		X"2A",X"0C",X"30",X"7D",X"A1",X"B3",X"6F",X"7C",X"A0",X"B2",X"67",X"22",X"0C",X"30",X"77",X"C9",
		X"DD",X"35",X"01",X"20",X"20",X"DD",X"7E",X"08",X"DD",X"77",X"01",X"DD",X"35",X"00",X"28",X"38",
		X"DD",X"CB",X"00",X"46",X"C8",X"DD",X"7E",X"09",X"B7",X"C8",X"DD",X"86",X"07",X"F8",X"DD",X"77",
		X"07",X"4F",X"C3",X"AD",X"01",X"DD",X"7E",X"0A",X"FE",X"01",X"D8",X"DD",X"6E",X"0B",X"DD",X"66",
		X"0C",X"28",X"0B",X"DD",X"46",X"01",X"0E",X"9B",X"09",X"7C",X"AD",X"6F",X"26",X"01",X"23",X"DD",
		X"75",X"0B",X"DD",X"74",X"0C",X"C3",X"C0",X"01",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"7E",X"57",
		X"E6",X"1F",X"28",X"2A",X"FE",X"1F",X"28",X"3D",X"CD",X"8E",X"02",X"7A",X"E6",X"1F",X"3D",X"07",
		X"4F",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"09",X"5E",X"23",X"56",X"EB",X"DD",X"75",X"0B",X"DD",
		X"74",X"0C",X"CD",X"C0",X"01",X"DD",X"4E",X"06",X"DD",X"71",X"07",X"C3",X"AD",X"01",X"23",X"DD",
		X"75",X"02",X"DD",X"74",X"03",X"7A",X"E6",X"E0",X"07",X"07",X"07",X"47",X"3E",X"80",X"07",X"10",
		X"FD",X"DD",X"77",X"00",X"C9",X"7A",X"E6",X"E0",X"07",X"07",X"07",X"11",X"58",X"02",X"D5",X"23",
		X"5D",X"54",X"23",X"DD",X"75",X"02",X"DD",X"74",X"03",X"21",X"BF",X"02",X"C3",X"28",X"00",X"CF",
		X"02",X"E3",X"02",X"F3",X"02",X"F8",X"02",X"FD",X"02",X"02",X"03",X"0B",X"03",X"15",X"03",X"EB",
		X"4E",X"CB",X"21",X"06",X"00",X"21",X"1A",X"03",X"09",X"5E",X"23",X"56",X"DD",X"73",X"04",X"DD",
		X"72",X"05",X"C9",X"EB",X"4E",X"06",X"00",X"21",X"B2",X"03",X"09",X"7E",X"DD",X"77",X"08",X"DD",
		X"77",X"01",X"C9",X"1A",X"DD",X"77",X"06",X"C9",X"1A",X"DD",X"77",X"09",X"C9",X"1A",X"DD",X"77",
		X"0A",X"C9",X"1A",X"32",X"0A",X"30",X"AF",X"32",X"0B",X"30",X"C9",X"1A",X"DD",X"77",X"02",X"13",
		X"1A",X"DD",X"77",X"03",X"C9",X"E1",X"E1",X"3E",X"FF",X"C9",X"3A",X"03",X"3E",X"03",X"42",X"03",
		X"46",X"03",X"4A",X"03",X"4E",X"03",X"52",X"03",X"56",X"03",X"5A",X"03",X"5E",X"03",X"62",X"03",
		X"66",X"03",X"6A",X"03",X"6E",X"03",X"72",X"03",X"76",X"03",X"6B",X"08",X"F2",X"07",X"80",X"07",
		X"14",X"07",X"AE",X"06",X"4E",X"06",X"F3",X"05",X"9E",X"05",X"4E",X"05",X"01",X"05",X"B9",X"04",
		X"76",X"04",X"36",X"04",X"F9",X"03",X"C0",X"03",X"8A",X"03",X"57",X"03",X"27",X"03",X"FA",X"02",
		X"CF",X"02",X"A7",X"02",X"81",X"02",X"5D",X"02",X"3B",X"02",X"1B",X"02",X"FD",X"01",X"E0",X"01",
		X"C5",X"01",X"AC",X"01",X"94",X"01",X"7D",X"01",X"68",X"01",X"53",X"01",X"40",X"01",X"2E",X"01",
		X"1D",X"01",X"0D",X"01",X"FE",X"00",X"F0",X"00",X"E3",X"00",X"D6",X"00",X"CA",X"00",X"BE",X"00",
		X"B4",X"00",X"AA",X"00",X"A0",X"00",X"97",X"00",X"8F",X"00",X"87",X"00",X"7F",X"00",X"78",X"00",
		X"71",X"00",X"6B",X"00",X"65",X"00",X"5F",X"00",X"5A",X"00",X"55",X"00",X"50",X"00",X"4C",X"00",
		X"47",X"00",X"3C",X"38",X"34",X"30",X"2C",X"28",X"24",X"20",X"1E",X"1C",X"1A",X"18",X"16",X"14",
		X"12",X"10",X"0F",X"0E",X"0D",X"0C",X"0B",X"0A",X"09",X"08",X"07",X"06",X"05",X"04",X"21",X"FD",
		X"03",X"11",X"0F",X"30",X"01",X"27",X"00",X"ED",X"B0",X"07",X"4F",X"07",X"81",X"4F",X"06",X"00",
		X"21",X"DB",X"0A",X"09",X"11",X"11",X"30",X"CD",X"F3",X"03",X"11",X"1E",X"30",X"CD",X"F3",X"03",
		X"11",X"2B",X"30",X"7E",X"12",X"CD",X"FA",X"03",X"7E",X"12",X"23",X"13",X"C9",X"01",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"3E",X"01",X"CD",X"DC",X"01",X"21",X"3B",X"30",X"36",X"00",X"2C",X"36",
		X"03",X"2C",X"0E",X"06",X"71",X"CD",X"AD",X"01",X"21",X"18",X"00",X"22",X"39",X"30",X"CD",X"C0",
		X"01",X"AF",X"C9",X"21",X"3B",X"30",X"35",X"7E",X"57",X"E6",X"0F",X"20",X"1F",X"2C",X"7E",X"2C",
		X"86",X"FE",X"05",X"28",X"2D",X"77",X"FE",X"0F",X"20",X"0E",X"2D",X"36",X"FE",X"2A",X"39",X"30",
		X"01",X"F4",X"FF",X"09",X"22",X"39",X"30",X"3D",X"4F",X"CD",X"AD",X"01",X"2A",X"39",X"30",X"CB",
		X"62",X"01",X"02",X"00",X"20",X"03",X"01",X"FE",X"FF",X"09",X"22",X"39",X"30",X"CD",X"C0",X"01",
		X"AF",X"C9",X"3E",X"FF",X"C9",X"AF",X"CD",X"DC",X"01",X"0E",X"06",X"CD",X"AD",X"01",X"21",X"90",
		X"00",X"CD",X"C0",X"01",X"21",X"3E",X"30",X"36",X"00",X"2C",X"36",X"F4",X"2C",X"36",X"90",X"AF",
		X"C9",X"21",X"3E",X"30",X"35",X"7E",X"E6",X"07",X"20",X"1A",X"0E",X"00",X"CB",X"5E",X"20",X"11",
		X"2C",X"34",X"34",X"28",X"D4",X"7E",X"2C",X"86",X"77",X"6F",X"26",X"00",X"CD",X"C0",X"01",X"0E",
		X"06",X"CD",X"AD",X"01",X"AF",X"C9",X"3E",X"01",X"CD",X"DC",X"01",X"21",X"41",X"30",X"0E",X"0D",
		X"71",X"CD",X"AD",X"01",X"2C",X"36",X"80",X"2C",X"36",X"20",X"6E",X"26",X"03",X"CD",X"C0",X"01",
		X"AF",X"C9",X"21",X"42",X"30",X"35",X"7E",X"28",X"1E",X"E6",X"0F",X"20",X"07",X"2D",X"35",X"4E",
		X"CD",X"AD",X"01",X"2C",X"CB",X"5E",X"3E",X"08",X"20",X"02",X"ED",X"44",X"2C",X"86",X"77",X"6F",
		X"26",X"03",X"CD",X"C0",X"01",X"AF",X"C9",X"3D",X"C9",X"3E",X"01",X"CD",X"DC",X"01",X"0E",X"0B",
		X"CD",X"AD",X"01",X"21",X"B0",X"00",X"CD",X"C0",X"01",X"21",X"44",X"30",X"36",X"00",X"2C",X"36",
		X"B0",X"2C",X"36",X"84",X"2C",X"36",X"B0",X"AF",X"C9",X"21",X"44",X"30",X"35",X"7E",X"E6",X"01",
		X"20",X"0D",X"2C",X"35",X"7E",X"2C",X"BE",X"28",X"08",X"6F",X"26",X"00",X"CD",X"C0",X"01",X"AF",
		X"C9",X"2C",X"86",X"1F",X"FE",X"40",X"38",X"15",X"77",X"32",X"45",X"30",X"6F",X"26",X"00",X"CD",
		X"C0",X"01",X"7D",X"CB",X"3D",X"CB",X"3D",X"95",X"32",X"46",X"30",X"AF",X"C9",X"3E",X"FF",X"C9",
		X"AF",X"CD",X"DC",X"01",X"21",X"18",X"00",X"CD",X"C0",X"01",X"21",X"48",X"30",X"36",X"1E",X"2C",
		X"0E",X"0F",X"71",X"CD",X"AD",X"01",X"2C",X"36",X"53",X"2C",X"36",X"35",X"AF",X"C9",X"21",X"48",
		X"30",X"35",X"7E",X"28",X"1E",X"2C",X"E6",X"01",X"20",X"05",X"35",X"4E",X"CD",X"AD",X"01",X"2C",
		X"7E",X"C6",X"95",X"77",X"2C",X"AE",X"E6",X"7F",X"C6",X"30",X"77",X"6F",X"26",X"00",X"CD",X"C0",
		X"01",X"AF",X"C9",X"3D",X"C9",X"AF",X"CD",X"DC",X"01",X"21",X"4C",X"30",X"36",X"40",X"2C",X"36",
		X"A0",X"21",X"A0",X"00",X"CD",X"C0",X"01",X"0E",X"0B",X"CD",X"AD",X"01",X"AF",X"C9",X"21",X"4C",
		X"30",X"35",X"7E",X"28",X"26",X"FE",X"20",X"28",X"E5",X"57",X"E6",X"03",X"20",X"1B",X"7A",X"E6",
		X"07",X"20",X"0B",X"2C",X"7E",X"D6",X"20",X"77",X"6F",X"26",X"00",X"CD",X"C0",X"01",X"CB",X"52",
		X"0E",X"07",X"20",X"02",X"0E",X"0B",X"CD",X"AD",X"01",X"AF",X"C9",X"3D",X"C9",X"AF",X"CD",X"DC",
		X"01",X"0E",X"09",X"CD",X"AD",X"01",X"21",X"40",X"00",X"CD",X"C0",X"01",X"21",X"4E",X"30",X"36",
		X"80",X"2C",X"36",X"40",X"AF",X"C9",X"21",X"4E",X"30",X"35",X"7E",X"28",X"11",X"E6",X"1F",X"20",
		X"0B",X"2C",X"7E",X"D6",X"06",X"77",X"6F",X"26",X"00",X"CD",X"C0",X"01",X"AF",X"C9",X"3D",X"C9",
		X"AF",X"CD",X"DC",X"01",X"21",X"50",X"30",X"36",X"B6",X"2C",X"0E",X"00",X"71",X"CD",X"AD",X"01",
		X"2C",X"36",X"30",X"21",X"30",X"00",X"CD",X"C0",X"01",X"AF",X"C9",X"21",X"50",X"30",X"35",X"7E",
		X"28",X"35",X"2C",X"FE",X"80",X"38",X"15",X"FE",X"83",X"38",X"07",X"FE",X"B2",X"3E",X"00",X"D8",
		X"28",X"03",X"7E",X"C6",X"04",X"77",X"4F",X"CD",X"AD",X"01",X"AF",X"C9",X"57",X"E6",X"0F",X"20",
		X"05",X"35",X"4E",X"CD",X"AD",X"01",X"2C",X"35",X"CB",X"5A",X"28",X"03",X"34",X"34",X"34",X"6E",
		X"26",X"00",X"CD",X"C0",X"01",X"AF",X"C9",X"3D",X"C9",X"AF",X"CD",X"DC",X"01",X"0E",X"0C",X"CD",
		X"AD",X"01",X"21",X"0F",X"00",X"CD",X"C0",X"01",X"3E",X"10",X"32",X"53",X"30",X"AF",X"C9",X"21",
		X"53",X"30",X"35",X"7E",X"28",X"0E",X"E6",X"01",X"21",X"0E",X"00",X"20",X"02",X"2E",X"0F",X"CD",
		X"C0",X"01",X"AF",X"C9",X"3D",X"C9",X"AF",X"CD",X"DC",X"01",X"0E",X"09",X"CD",X"AD",X"01",X"21",
		X"40",X"00",X"CD",X"C0",X"01",X"21",X"54",X"30",X"36",X"80",X"2C",X"36",X"40",X"AF",X"C9",X"21",
		X"54",X"30",X"35",X"7E",X"28",X"18",X"57",X"E6",X"1F",X"20",X"11",X"2C",X"7E",X"D6",X"0C",X"CB",
		X"6A",X"20",X"02",X"C6",X"18",X"77",X"6F",X"26",X"00",X"CD",X"C0",X"01",X"AF",X"C9",X"3D",X"C9",
		X"3E",X"01",X"CD",X"DC",X"01",X"0E",X"0E",X"CD",X"AD",X"01",X"21",X"56",X"30",X"36",X"00",X"2C",
		X"36",X"60",X"6E",X"26",X"00",X"CD",X"C0",X"01",X"AF",X"C9",X"21",X"56",X"30",X"35",X"7E",X"28",
		X"0D",X"FE",X"80",X"38",X"04",X"E6",X"1F",X"28",X"E6",X"2C",X"34",X"C3",X"F2",X"06",X"3D",X"C9",
		X"3E",X"01",X"CD",X"DC",X"01",X"21",X"F8",X"00",X"22",X"58",X"30",X"CD",X"C0",X"01",X"0E",X"01",
		X"CD",X"AD",X"01",X"21",X"5A",X"30",X"36",X"00",X"2C",X"36",X"A0",X"AF",X"C9",X"21",X"5A",X"30",
		X"35",X"56",X"CB",X"46",X"20",X"2E",X"2C",X"35",X"7E",X"28",X"4B",X"2A",X"58",X"30",X"FE",X"0B",
		X"38",X"33",X"FE",X"90",X"38",X"38",X"01",X"10",X"00",X"28",X"15",X"FE",X"9B",X"38",X"0C",X"5F",
		X"C6",X"60",X"ED",X"44",X"87",X"3C",X"4F",X"CD",X"AD",X"01",X"7B",X"C6",X"60",X"4F",X"06",X"FF",
		X"09",X"22",X"58",X"30",X"2A",X"58",X"30",X"7A",X"B7",X"EA",X"70",X"07",X"01",X"06",X"00",X"09",
		X"CD",X"C0",X"01",X"AF",X"C9",X"4F",X"CD",X"AD",X"01",X"23",X"23",X"C3",X"61",X"07",X"E6",X"07",
		X"20",X"E5",X"23",X"C3",X"61",X"07",X"3D",X"C9",X"AF",X"CD",X"DC",X"01",X"21",X"40",X"00",X"CD",
		X"C0",X"01",X"0E",X"00",X"CD",X"AD",X"01",X"21",X"5C",X"30",X"36",X"20",X"AF",X"2C",X"77",X"2C",
		X"36",X"40",X"C9",X"21",X"5C",X"30",X"35",X"7E",X"28",X"18",X"E6",X"01",X"4F",X"28",X"0E",X"2C",
		X"34",X"7E",X"2C",X"86",X"77",X"6F",X"26",X"00",X"CD",X"C0",X"01",X"0E",X"0A",X"CD",X"AD",X"01",
		X"AF",X"C9",X"3D",X"C9",X"AF",X"CD",X"DC",X"01",X"0E",X"05",X"CD",X"AD",X"01",X"AF",X"21",X"5F",
		X"30",X"36",X"80",X"2C",X"77",X"2C",X"77",X"C9",X"21",X"5F",X"30",X"35",X"7E",X"28",X"1A",X"57",
		X"FE",X"08",X"38",X"23",X"FE",X"30",X"30",X"13",X"2C",X"7E",X"C6",X"C3",X"77",X"2C",X"AE",X"AA",
		X"77",X"6F",X"26",X"02",X"CD",X"C0",X"01",X"AF",X"C9",X"3D",X"C9",X"E6",X"07",X"20",X"E9",X"7A",
		X"0F",X"0F",X"0F",X"4F",X"3E",X"15",X"91",X"4F",X"CD",X"AD",X"01",X"AF",X"C9",X"3E",X"01",X"CD",
		X"DC",X"01",X"21",X"62",X"30",X"36",X"80",X"2C",X"0E",X"0F",X"71",X"CD",X"AD",X"01",X"2C",X"36",
		X"23",X"2C",X"36",X"D7",X"21",X"4C",X"01",X"CD",X"C0",X"01",X"AF",X"C9",X"21",X"62",X"30",X"35",
		X"7E",X"28",X"30",X"2C",X"FE",X"78",X"28",X"23",X"FE",X"70",X"28",X"1F",X"FE",X"68",X"28",X"1B",
		X"30",X"04",X"E6",X"07",X"20",X"05",X"35",X"4E",X"CD",X"AD",X"01",X"2C",X"7E",X"C6",X"5D",X"77",
		X"2C",X"AE",X"77",X"6F",X"26",X"01",X"CD",X"C0",X"01",X"AF",X"C9",X"0E",X"0F",X"71",X"CD",X"AD",
		X"01",X"AF",X"C9",X"3D",X"C9",X"AF",X"CD",X"DC",X"01",X"21",X"69",X"30",X"36",X"0C",X"4E",X"CD",
		X"AD",X"01",X"2D",X"36",X"00",X"21",X"80",X"00",X"22",X"66",X"30",X"CD",X"C0",X"01",X"AF",X"C9",
		X"21",X"68",X"30",X"34",X"7E",X"FE",X"59",X"28",X"0F",X"4F",X"06",X"00",X"2A",X"66",X"30",X"09",
		X"22",X"66",X"30",X"CD",X"C0",X"01",X"AF",X"C9",X"2C",X"7E",X"D6",X"04",X"28",X"04",X"77",X"C3",
		X"6E",X"08",X"3D",X"C9",X"AF",X"CD",X"DC",X"01",X"21",X"20",X"04",X"CD",X"C0",X"01",X"21",X"6A",
		X"30",X"36",X"00",X"2C",X"0E",X"0F",X"71",X"CD",X"AD",X"01",X"AF",X"C9",X"21",X"6A",X"30",X"35",
		X"7E",X"57",X"E6",X"0F",X"20",X"10",X"2C",X"7E",X"3C",X"CB",X"62",X"28",X"04",X"D6",X"03",X"28",
		X"07",X"77",X"4F",X"CD",X"AD",X"01",X"AF",X"C9",X"3D",X"C9",X"AF",X"CD",X"DC",X"01",X"21",X"50",
		X"00",X"CD",X"C0",X"01",X"21",X"6C",X"30",X"36",X"48",X"2C",X"0E",X"0F",X"71",X"CD",X"AD",X"01",
		X"AF",X"C9",X"21",X"6C",X"30",X"35",X"7E",X"28",X"13",X"57",X"E6",X"03",X"20",X"0C",X"2C",X"CB",
		X"52",X"0E",X"06",X"20",X"02",X"35",X"4E",X"CD",X"AD",X"01",X"AF",X"C9",X"3D",X"C9",X"AF",X"CD",
		X"DC",X"01",X"21",X"6E",X"30",X"36",X"09",X"2C",X"36",X"60",X"2C",X"0E",X"0C",X"71",X"CD",X"AD",
		X"01",X"2C",X"36",X"40",X"6E",X"26",X"00",X"CD",X"C0",X"01",X"AF",X"C9",X"21",X"6F",X"30",X"35",
		X"7E",X"28",X"24",X"FE",X"40",X"20",X"05",X"2D",X"35",X"20",X"DC",X"2C",X"57",X"E6",X"01",X"20",
		X"E9",X"2C",X"7A",X"E6",X"07",X"20",X"05",X"35",X"4E",X"CD",X"AD",X"01",X"2C",X"34",X"CB",X"52",
		X"20",X"D2",X"35",X"35",X"C3",X"24",X"09",X"3D",X"C9",X"3E",X"01",X"CD",X"DC",X"01",X"21",X"00",
		X"01",X"22",X"72",X"30",X"CD",X"C0",X"01",X"0E",X"05",X"CD",X"AD",X"01",X"21",X"74",X"30",X"36",
		X"00",X"2C",X"36",X"A0",X"AF",X"C9",X"21",X"74",X"30",X"35",X"7E",X"57",X"E6",X"03",X"20",X"2F",
		X"2C",X"35",X"7E",X"28",X"4C",X"2A",X"72",X"30",X"FE",X"0F",X"38",X"34",X"FE",X"90",X"38",X"39",
		X"01",X"10",X"00",X"28",X"16",X"FE",X"9B",X"38",X"0D",X"5F",X"C6",X"60",X"ED",X"44",X"87",X"C6",
		X"05",X"4F",X"CD",X"AD",X"01",X"7B",X"C6",X"60",X"4F",X"06",X"FF",X"09",X"22",X"72",X"30",X"2A",
		X"72",X"30",X"7A",X"B7",X"EA",X"BB",X"09",X"01",X"06",X"00",X"09",X"CD",X"C0",X"01",X"AF",X"C9",
		X"4F",X"CD",X"AD",X"01",X"23",X"23",X"C3",X"AC",X"09",X"E6",X"07",X"20",X"E5",X"23",X"C3",X"AC",
		X"09",X"3D",X"C9",X"AB",X"01",X"24",X"04",X"85",X"04",X"C6",X"04",X"09",X"05",X"60",X"05",X"A5",
		X"05",X"ED",X"05",X"20",X"06",X"79",X"06",X"A6",X"06",X"E0",X"06",X"10",X"07",X"88",X"07",X"C4",
		X"07",X"0D",X"08",X"65",X"08",X"A4",X"08",X"DA",X"08",X"0E",X"09",X"59",X"09",X"BA",X"0A",X"BA",
		X"0A",X"BA",X"0A",X"59",X"0A",X"5D",X"0A",X"62",X"0A",X"67",X"0A",X"6C",X"0A",X"71",X"0A",X"76",
		X"0A",X"7B",X"0A",X"80",X"0A",X"85",X"0A",X"8A",X"0A",X"8F",X"0A",X"94",X"0A",X"99",X"0A",X"9E",
		X"0A",X"A3",X"0A",X"A8",X"0A",X"AD",X"0A",X"B2",X"0A",X"00",X"00",X"43",X"04",X"A1",X"04",X"E2",
		X"04",X"29",X"05",X"7E",X"05",X"BE",X"05",X"06",X"06",X"3B",X"06",X"8F",X"06",X"BF",X"06",X"FA",
		X"06",X"2D",X"07",X"A3",X"07",X"D8",X"07",X"2C",X"08",X"80",X"08",X"BC",X"08",X"F2",X"08",X"2C",
		X"09",X"76",X"09",X"C0",X"0A",X"C9",X"0A",X"D2",X"0A",X"AF",X"C3",X"B4",X"0A",X"3E",X"01",X"C3",
		X"B4",X"0A",X"3E",X"02",X"C3",X"B4",X"0A",X"3E",X"03",X"C3",X"B4",X"0A",X"3E",X"04",X"C3",X"B4",
		X"0A",X"3E",X"05",X"C3",X"B4",X"0A",X"3E",X"06",X"C3",X"B4",X"0A",X"3E",X"07",X"C3",X"B4",X"0A",
		X"3E",X"08",X"C3",X"B4",X"0A",X"3E",X"09",X"C3",X"B4",X"0A",X"3E",X"0A",X"C3",X"B4",X"0A",X"3E",
		X"0B",X"C3",X"B4",X"0A",X"3E",X"0C",X"C3",X"B4",X"0A",X"3E",X"0D",X"C3",X"B4",X"0A",X"3E",X"0E",
		X"C3",X"B4",X"0A",X"3E",X"0F",X"C3",X"B4",X"0A",X"3E",X"10",X"C3",X"B4",X"0A",X"3E",X"11",X"C3",
		X"B4",X"0A",X"3E",X"12",X"CD",X"CE",X"03",X"3E",X"FF",X"C9",X"AF",X"CD",X"DC",X"01",X"AF",X"C9",
		X"DD",X"21",X"0F",X"30",X"CD",X"10",X"02",X"AF",X"C9",X"DD",X"21",X"1C",X"30",X"CD",X"10",X"02",
		X"AF",X"C9",X"DD",X"21",X"29",X"30",X"CD",X"10",X"02",X"AF",X"C9",X"4D",X"0B",X"5E",X"0B",X"5E",
		X"0B",X"5F",X"0B",X"72",X"0B",X"72",X"0B",X"73",X"0B",X"CD",X"0B",X"13",X"0C",X"3F",X"0C",X"8D",
		X"0C",X"C7",X"0C",X"01",X"0D",X"42",X"0D",X"6A",X"0D",X"91",X"0D",X"BB",X"0D",X"DD",X"0D",X"ED",
		X"0D",X"27",X"0E",X"27",X"0E",X"28",X"0E",X"65",X"0E",X"65",X"0E",X"66",X"0E",X"9C",X"0E",X"9C",
		X"0E",X"9D",X"0E",X"E6",X"0E",X"E6",X"0E",X"E7",X"0E",X"0C",X"0F",X"31",X"0F",X"75",X"0F",X"C2",
		X"0F",X"03",X"10",X"44",X"10",X"6E",X"10",X"9F",X"10",X"EE",X"10",X"37",X"11",X"7E",X"11",X"C5",
		X"11",X"F0",X"11",X"F0",X"11",X"F1",X"11",X"3A",X"12",X"3A",X"12",X"3B",X"12",X"79",X"12",X"B6",
		X"12",X"F1",X"12",X"81",X"13",X"AF",X"14",X"B0",X"15",X"B0",X"15",X"B0",X"15",X"1F",X"0F",X"3F",
		X"1B",X"5F",X"0A",X"9F",X"02",X"A1",X"81",X"81",X"A1",X"81",X"81",X"DF",X"55",X"0B",X"FF",X"1F",
		X"0F",X"3F",X"1B",X"5F",X"0A",X"9F",X"02",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"DF",
		X"67",X"0B",X"FF",X"1F",X"0C",X"3F",X"16",X"5F",X"06",X"8B",X"8D",X"8B",X"6D",X"6E",X"6F",X"92",
		X"60",X"94",X"92",X"97",X"60",X"76",X"79",X"97",X"96",X"99",X"60",X"97",X"94",X"92",X"72",X"72",
		X"74",X"92",X"97",X"60",X"76",X"77",X"74",X"72",X"8F",X"AD",X"60",X"71",X"74",X"77",X"76",X"77",
		X"76",X"74",X"72",X"70",X"6F",X"6D",X"8B",X"8D",X"8B",X"6D",X"6E",X"6F",X"6F",X"92",X"94",X"92",
		X"94",X"60",X"76",X"79",X"97",X"96",X"76",X"99",X"97",X"94",X"92",X"92",X"77",X"8B",X"AD",X"B2",
		X"60",X"7F",X"00",X"CB",X"7F",X"FF",X"8B",X"8B",X"8D",X"8E",X"DF",X"79",X"0B",X"1F",X"0C",X"3F",
		X"16",X"5F",X"06",X"86",X"86",X"86",X"86",X"86",X"86",X"86",X"86",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"86",X"86",X"86",X"86",X"88",X"88",X"88",X"88",X"85",X"85",X"85",X"85",X"86",
		X"86",X"86",X"86",X"86",X"86",X"86",X"86",X"86",X"86",X"86",X"86",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"86",X"86",X"86",X"86",X"86",X"86",X"86",X"86",X"86",X"86",X"86",X"86",X"C6",
		X"DF",X"D3",X"0B",X"1F",X"06",X"3F",X"16",X"5F",X"06",X"AB",X"A6",X"AB",X"8D",X"8F",X"B0",X"AB",
		X"B0",X"B0",X"AF",X"AF",X"A8",X"A8",X"AD",X"AD",X"A6",X"88",X"8A",X"AB",X"A6",X"AB",X"8D",X"8F",
		X"B0",X"AB",X"B0",X"B0",X"AF",X"AF",X"A6",X"88",X"8A",X"AB",X"A6",X"CB",X"DF",X"19",X"0C",X"1F",
		X"0F",X"3F",X"17",X"5F",X"07",X"8F",X"8B",X"8B",X"6D",X"6F",X"90",X"8D",X"8D",X"92",X"8F",X"8B",
		X"8B",X"8B",X"6D",X"6B",X"6A",X"68",X"A6",X"8F",X"8B",X"8B",X"6D",X"6F",X"90",X"8D",X"8D",X"92",
		X"8F",X"8B",X"8D",X"8A",X"8B",X"8B",X"AB",X"92",X"92",X"92",X"70",X"72",X"94",X"90",X"90",X"90",
		X"94",X"94",X"94",X"72",X"70",X"94",X"94",X"94",X"72",X"70",X"8F",X"8B",X"8B",X"6D",X"6F",X"90",
		X"8D",X"8D",X"92",X"8F",X"8B",X"8D",X"8A",X"8B",X"8B",X"AB",X"DF",X"45",X"0C",X"1F",X"05",X"3F",
		X"17",X"5F",X"06",X"87",X"97",X"B7",X"82",X"95",X"B5",X"87",X"97",X"B7",X"82",X"95",X"95",X"95",
		X"87",X"97",X"B7",X"82",X"95",X"B5",X"82",X"97",X"B8",X"97",X"97",X"B7",X"87",X"97",X"B7",X"8C",
		X"98",X"B8",X"8C",X"98",X"B8",X"87",X"97",X"B7",X"87",X"97",X"B7",X"82",X"95",X"B5",X"82",X"97",
		X"B8",X"97",X"97",X"B7",X"DF",X"93",X"0C",X"1F",X"05",X"3F",X"17",X"5F",X"06",X"87",X"8E",X"AE",
		X"82",X"8E",X"AE",X"87",X"8E",X"AE",X"82",X"8E",X"8E",X"8E",X"87",X"8E",X"AE",X"82",X"8E",X"AE",
		X"82",X"8E",X"AE",X"93",X"93",X"B3",X"87",X"8E",X"AE",X"8C",X"90",X"B0",X"8C",X"90",X"B0",X"87",
		X"8E",X"AE",X"87",X"8E",X"AE",X"82",X"8E",X"AE",X"82",X"8E",X"AE",X"93",X"93",X"B3",X"DF",X"CD",
		X"0C",X"1F",X"0E",X"3F",X"18",X"5F",X"09",X"88",X"87",X"88",X"85",X"94",X"93",X"94",X"91",X"85",
		X"84",X"85",X"81",X"91",X"90",X"91",X"8D",X"85",X"83",X"81",X"83",X"91",X"8F",X"8D",X"8F",X"88",
		X"8A",X"88",X"85",X"94",X"96",X"94",X"91",X"88",X"8A",X"8C",X"AD",X"A8",X"A5",X"A1",X"7F",X"00",
		X"CA",X"7F",X"FF",X"8A",X"8A",X"8C",X"8A",X"A8",X"A6",X"A5",X"A3",X"7F",X"00",X"C1",X"7F",X"FF",
		X"A1",X"FF",X"1F",X"0E",X"3F",X"18",X"5F",X"00",X"A1",X"A0",X"5F",X"09",X"A5",X"A5",X"80",X"A0",
		X"85",X"A5",X"A5",X"80",X"85",X"A5",X"A6",X"A6",X"A6",X"A6",X"A5",X"85",X"A5",X"A6",X"80",X"A5",
		X"C0",X"A5",X"A6",X"86",X"A6",X"C4",X"A8",X"A8",X"A8",X"FF",X"1F",X"08",X"3F",X"18",X"5F",X"00",
		X"A1",X"80",X"5F",X"08",X"AD",X"A8",X"AD",X"C8",X"A8",X"80",X"8D",X"A8",X"A3",X"A8",X"A3",X"A8",
		X"AD",X"C8",X"A8",X"AD",X"A8",X"AD",X"A5",X"A6",X"A1",X"A6",X"A7",X"A8",X"A8",X"AA",X"CC",X"C8",
		X"FF",X"1F",X"0E",X"3F",X"16",X"5F",X"09",X"69",X"89",X"69",X"86",X"89",X"A7",X"24",X"24",X"25",
		X"25",X"26",X"26",X"26",X"26",X"87",X"66",X"86",X"66",X"84",X"81",X"3F",X"10",X"22",X"23",X"24",
		X"25",X"26",X"27",X"28",X"29",X"2A",X"2B",X"2C",X"2D",X"AE",X"FF",X"1F",X"0E",X"3F",X"16",X"5F",
		X"09",X"66",X"86",X"66",X"82",X"86",X"A4",X"A0",X"62",X"82",X"62",X"81",X"80",X"3F",X"10",X"26",
		X"27",X"28",X"29",X"2A",X"2B",X"2C",X"2D",X"2E",X"2F",X"30",X"31",X"B2",X"FF",X"1F",X"08",X"3F",
		X"16",X"5F",X"08",X"A2",X"A0",X"A4",X"A0",X"A2",X"A1",X"3F",X"10",X"A2",X"FF",X"1F",X"0F",X"3F",
		X"1A",X"5F",X"0C",X"9F",X"02",X"81",X"81",X"A1",X"81",X"81",X"A1",X"81",X"81",X"81",X"81",X"A1",
		X"A1",X"81",X"81",X"A1",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"A1",X"A1",X"81",X"81",
		X"A1",X"81",X"81",X"A1",X"81",X"81",X"81",X"81",X"A1",X"A1",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"A1",X"81",X"81",X"A1",X"FF",X"FF",X"1F",X"0F",X"3F",X"1A",X"5F",X"0C",X"9F",X"02",
		X"81",X"81",X"A1",X"81",X"81",X"A1",X"A1",X"A1",X"61",X"61",X"61",X"61",X"81",X"81",X"81",X"81",
		X"A1",X"81",X"81",X"A1",X"A1",X"A1",X"61",X"61",X"61",X"61",X"81",X"81",X"81",X"81",X"A1",X"61",
		X"61",X"61",X"61",X"81",X"81",X"81",X"81",X"A1",X"61",X"61",X"61",X"61",X"81",X"81",X"81",X"81",
		X"81",X"81",X"A1",X"A1",X"A1",X"FF",X"1F",X"0F",X"3F",X"1A",X"5F",X"0C",X"9F",X"02",X"81",X"A1",
		X"A1",X"A1",X"80",X"81",X"A1",X"A1",X"A1",X"80",X"81",X"A1",X"61",X"61",X"61",X"61",X"61",X"61",
		X"81",X"A1",X"61",X"61",X"61",X"61",X"61",X"61",X"81",X"A1",X"A1",X"A1",X"80",X"81",X"A1",X"A1",
		X"A1",X"80",X"81",X"A1",X"81",X"81",X"A1",X"A1",X"A1",X"81",X"81",X"A1",X"FF",X"1F",X"0F",X"3F",
		X"1A",X"5F",X"0C",X"9F",X"02",X"A1",X"A1",X"61",X"61",X"61",X"61",X"61",X"61",X"61",X"61",X"A1",
		X"A1",X"61",X"61",X"61",X"61",X"61",X"61",X"61",X"61",X"A1",X"A1",X"81",X"A1",X"81",X"A1",X"A1",
		X"61",X"61",X"61",X"61",X"61",X"61",X"61",X"61",X"A1",X"A1",X"61",X"61",X"61",X"61",X"61",X"61",
		X"61",X"61",X"A1",X"A1",X"61",X"61",X"61",X"61",X"61",X"61",X"61",X"61",X"A1",X"A1",X"81",X"A1",
		X"81",X"81",X"81",X"81",X"81",X"A1",X"FF",X"1F",X"0E",X"3F",X"16",X"5F",X"09",X"95",X"97",X"99",
		X"9A",X"95",X"95",X"B5",X"93",X"92",X"B3",X"92",X"90",X"B2",X"90",X"AE",X"8B",X"8D",X"8E",X"AD",
		X"8E",X"B0",X"AE",X"E0",X"C0",X"A0",X"97",X"95",X"8B",X"8D",X"AE",X"FF",X"1F",X"0E",X"3F",X"16",
		X"5F",X"09",X"92",X"93",X"95",X"95",X"92",X"92",X"B2",X"90",X"8E",X"B0",X"8E",X"8D",X"AE",X"8D",
		X"AB",X"87",X"89",X"8B",X"A9",X"8B",X"AD",X"A9",X"E0",X"C0",X"A0",X"93",X"92",X"87",X"89",X"AB",
		X"FF",X"1F",X"02",X"3F",X"16",X"5F",X"00",X"A1",X"80",X"5F",X"09",X"8E",X"95",X"92",X"95",X"8E",
		X"90",X"92",X"B3",X"97",X"8E",X"B2",X"95",X"AE",X"93",X"97",X"8E",X"97",X"8D",X"95",X"90",X"5F",
		X"0B",X"7F",X"FE",X"9F",X"02",X"61",X"61",X"81",X"81",X"81",X"61",X"61",X"81",X"81",X"81",X"61",
		X"61",X"81",X"81",X"61",X"81",X"61",X"81",X"81",X"A1",X"5F",X"09",X"7F",X"FF",X"9F",X"00",X"97",
		X"95",X"8B",X"8D",X"AE",X"FF",X"1F",X"0F",X"3F",X"18",X"5F",X"09",X"66",X"68",X"8A",X"8D",X"8D",
		X"8F",X"8D",X"8A",X"86",X"66",X"68",X"8A",X"8A",X"88",X"86",X"A8",X"88",X"66",X"68",X"8A",X"8D",
		X"8D",X"6D",X"6F",X"8D",X"8A",X"86",X"66",X"68",X"8A",X"8A",X"88",X"88",X"A6",X"86",X"66",X"68",
		X"8A",X"8D",X"8D",X"6D",X"6F",X"8D",X"8A",X"86",X"66",X"68",X"8A",X"8A",X"88",X"86",X"A8",X"80",
		X"66",X"68",X"8A",X"8D",X"8D",X"8F",X"8D",X"8A",X"86",X"66",X"68",X"8A",X"8A",X"88",X"68",X"68",
		X"A6",X"FF",X"1F",X"0B",X"3F",X"18",X"5F",X"00",X"81",X"5F",X"08",X"82",X"92",X"92",X"92",X"82",
		X"92",X"92",X"92",X"82",X"92",X"84",X"94",X"89",X"93",X"B3",X"82",X"92",X"92",X"92",X"82",X"92",
		X"B4",X"82",X"92",X"89",X"93",X"82",X"92",X"B2",X"82",X"92",X"92",X"92",X"82",X"92",X"92",X"92",
		X"82",X"92",X"84",X"94",X"89",X"93",X"B3",X"82",X"92",X"92",X"92",X"82",X"92",X"92",X"92",X"B2",
		X"B3",X"B2",X"FF",X"1F",X"05",X"3F",X"18",X"5F",X"00",X"81",X"5F",X"09",X"82",X"8E",X"8E",X"8E",
		X"82",X"8E",X"8E",X"8E",X"82",X"8E",X"84",X"90",X"89",X"90",X"B0",X"82",X"8E",X"8E",X"8E",X"82",
		X"8E",X"B0",X"82",X"8E",X"89",X"90",X"82",X"8E",X"AE",X"82",X"8E",X"8E",X"8E",X"82",X"8E",X"8E",
		X"8E",X"82",X"8E",X"84",X"90",X"89",X"90",X"B0",X"82",X"8E",X"8E",X"8E",X"92",X"8E",X"8E",X"8E",
		X"AE",X"B0",X"CE",X"FF",X"1F",X"0E",X"3F",X"17",X"5F",X"09",X"92",X"93",X"B5",X"92",X"93",X"B5",
		X"97",X"99",X"99",X"97",X"97",X"96",X"B7",X"90",X"92",X"B3",X"90",X"92",X"B3",X"99",X"97",X"95",
		X"93",X"92",X"90",X"AE",X"E0",X"E0",X"A0",X"97",X"95",X"93",X"92",X"90",X"AE",X"FF",X"1F",X"08",
		X"3F",X"17",X"5F",X"08",X"8B",X"8D",X"8E",X"95",X"92",X"95",X"8E",X"95",X"92",X"95",X"93",X"97",
		X"8E",X"97",X"93",X"97",X"8E",X"97",X"8D",X"95",X"90",X"95",X"8D",X"95",X"90",X"95",X"8E",X"95",
		X"92",X"95",X"AE",X"E0",X"E0",X"A0",X"1F",X"0E",X"93",X"92",X"90",X"8E",X"8D",X"B2",X"FF",X"1F",
		X"08",X"3F",X"17",X"5F",X"00",X"A1",X"80",X"5F",X"09",X"9A",X"80",X"9A",X"80",X"9A",X"80",X"9A",
		X"80",X"9A",X"80",X"9A",X"80",X"9A",X"80",X"9A",X"80",X"99",X"80",X"99",X"80",X"99",X"80",X"99",
		X"80",X"9A",X"80",X"9A",X"B2",X"80",X"5F",X"0B",X"7F",X"FE",X"9F",X"02",X"61",X"61",X"81",X"81",
		X"81",X"61",X"61",X"81",X"81",X"81",X"61",X"61",X"81",X"81",X"81",X"81",X"81",X"81",X"A1",X"5F",
		X"09",X"7F",X"FF",X"9F",X"00",X"5F",X"08",X"97",X"95",X"93",X"92",X"90",X"AE",X"FF",X"1F",X"0F",
		X"3F",X"18",X"5F",X"09",X"86",X"83",X"86",X"86",X"86",X"84",X"88",X"88",X"68",X"68",X"6A",X"6A",
		X"8A",X"88",X"8A",X"8B",X"8D",X"AF",X"83",X"86",X"86",X"86",X"84",X"88",X"88",X"88",X"8A",X"6A",
		X"6A",X"88",X"8A",X"8B",X"86",X"AB",X"86",X"86",X"86",X"66",X"66",X"88",X"88",X"A8",X"6A",X"6A",
		X"8A",X"88",X"8A",X"8B",X"8D",X"AF",X"86",X"86",X"86",X"66",X"66",X"88",X"88",X"A8",X"6A",X"6A",
		X"8A",X"88",X"8A",X"8B",X"86",X"AB",X"FF",X"1F",X"0A",X"3F",X"18",X"5F",X"00",X"81",X"5F",X"08",
		X"89",X"99",X"8D",X"99",X"81",X"9A",X"89",X"9A",X"84",X"9A",X"88",X"9A",X"89",X"99",X"B9",X"89",
		X"99",X"8D",X"99",X"82",X"9A",X"89",X"9A",X"84",X"9A",X"88",X"9A",X"89",X"99",X"B9",X"89",X"99",
		X"8D",X"99",X"81",X"9A",X"89",X"9A",X"84",X"9A",X"88",X"9A",X"89",X"99",X"8D",X"99",X"89",X"99",
		X"8D",X"99",X"82",X"9A",X"89",X"9A",X"84",X"9A",X"88",X"9A",X"89",X"99",X"B9",X"FF",X"1F",X"04",
		X"3F",X"18",X"5F",X"00",X"81",X"5F",X"09",X"89",X"90",X"8D",X"90",X"81",X"92",X"89",X"92",X"84",
		X"90",X"88",X"90",X"89",X"90",X"B0",X"89",X"90",X"8D",X"90",X"82",X"92",X"89",X"92",X"84",X"92",
		X"88",X"92",X"89",X"90",X"B0",X"89",X"90",X"8D",X"90",X"81",X"92",X"89",X"92",X"84",X"92",X"88",
		X"92",X"89",X"90",X"8D",X"90",X"89",X"90",X"8D",X"90",X"82",X"92",X"89",X"92",X"84",X"90",X"88",
		X"90",X"89",X"90",X"B0",X"FF",X"3F",X"1A",X"5F",X"07",X"1F",X"0F",X"7E",X"7C",X"7A",X"78",X"77",
		X"75",X"73",X"72",X"70",X"6E",X"6C",X"6B",X"69",X"67",X"66",X"64",X"62",X"1F",X"00",X"7E",X"7D",
		X"7B",X"79",X"78",X"76",X"74",X"72",X"71",X"6F",X"6D",X"6C",X"6A",X"68",X"66",X"65",X"63",X"61",
		X"FF",X"1F",X"0F",X"3F",X"1A",X"5F",X"0A",X"9F",X"02",X"A1",X"A1",X"61",X"61",X"61",X"61",X"61",
		X"61",X"61",X"61",X"A1",X"A1",X"61",X"61",X"61",X"61",X"61",X"61",X"61",X"61",X"A1",X"A1",X"81",
		X"A1",X"81",X"A1",X"A1",X"61",X"61",X"61",X"61",X"61",X"61",X"61",X"61",X"A1",X"A1",X"61",X"61",
		X"61",X"61",X"61",X"61",X"61",X"61",X"A1",X"A1",X"61",X"61",X"61",X"61",X"61",X"61",X"61",X"61",
		X"A1",X"A1",X"81",X"A1",X"81",X"81",X"81",X"81",X"81",X"C1",X"FF",X"1F",X"0D",X"3F",X"18",X"5F",
		X"09",X"AD",X"AF",X"B2",X"8D",X"8F",X"92",X"8D",X"8F",X"92",X"8D",X"8F",X"92",X"8D",X"8F",X"B2",
		X"80",X"8F",X"92",X"94",X"8F",X"92",X"94",X"8F",X"92",X"94",X"8F",X"92",X"B4",X"80",X"94",X"96",
		X"99",X"94",X"96",X"99",X"94",X"96",X"99",X"94",X"96",X"B9",X"9B",X"B9",X"B7",X"92",X"B4",X"8F",
		X"B2",X"8D",X"AF",X"88",X"AD",X"A6",X"DF",X"44",X"12",X"3F",X"18",X"5F",X"00",X"C1",X"A0",X"5F",
		X"07",X"1F",X"0D",X"92",X"92",X"92",X"92",X"92",X"B2",X"B2",X"92",X"92",X"92",X"92",X"92",X"94",
		X"94",X"94",X"94",X"94",X"B4",X"B4",X"94",X"94",X"94",X"94",X"94",X"99",X"99",X"99",X"99",X"99",
		X"B9",X"B9",X"99",X"99",X"B9",X"80",X"A0",X"1F",X"07",X"B7",X"92",X"B4",X"8F",X"B2",X"8D",X"AF",
		X"88",X"AD",X"A6",X"DF",X"81",X"12",X"3F",X"18",X"5F",X"00",X"C1",X"A0",X"5F",X"08",X"1F",X"07",
		X"86",X"86",X"A3",X"81",X"A3",X"86",X"86",X"86",X"A3",X"86",X"85",X"88",X"88",X"A5",X"83",X"A5",
		X"88",X"88",X"88",X"A5",X"88",X"86",X"8D",X"8D",X"AA",X"88",X"AA",X"8D",X"8D",X"8D",X"8A",X"AA",
		X"80",X"A0",X"1F",X"01",X"B7",X"92",X"B4",X"8F",X"B2",X"8D",X"AF",X"88",X"AD",X"A6",X"DF",X"BE",
		X"12",X"3F",X"16",X"5F",X"08",X"1F",X"02",X"7F",X"00",X"CD",X"7F",X"FF",X"CC",X"7F",X"00",X"CD",
		X"7F",X"FF",X"CC",X"7F",X"00",X"CD",X"7F",X"FF",X"CC",X"7F",X"00",X"CD",X"7F",X"FF",X"CC",X"1F",
		X"0E",X"80",X"A8",X"A8",X"A8",X"A8",X"A8",X"A8",X"A8",X"A8",X"A8",X"A8",X"A8",X"A8",X"A8",X"8F",
		X"7F",X"00",X"88",X"7F",X"FF",X"C8",X"A8",X"A8",X"A8",X"A8",X"A8",X"A8",X"A8",X"A8",X"A8",X"A8",
		X"A8",X"A8",X"A8",X"8F",X"7F",X"00",X"88",X"7F",X"FF",X"A8",X"80",X"81",X"85",X"88",X"8D",X"86",
		X"8A",X"8D",X"92",X"88",X"8C",X"91",X"94",X"94",X"91",X"8C",X"88",X"86",X"8A",X"8D",X"92",X"81",
		X"85",X"88",X"8D",X"1F",X"08",X"8A",X"92",X"94",X"99",X"1F",X"0E",X"88",X"8C",X"8F",X"94",X"81",
		X"85",X"88",X"8D",X"86",X"8A",X"8D",X"92",X"88",X"8C",X"91",X"94",X"94",X"91",X"8C",X"88",X"86",
		X"8A",X"8D",X"92",X"81",X"85",X"88",X"8D",X"AD",X"B2",X"7F",X"00",X"88",X"7F",X"FF",X"A8",X"80",
		X"FF",X"3F",X"16",X"1F",X"08",X"5F",X"09",X"7F",X"00",X"CD",X"7F",X"FF",X"8C",X"BF",X"14",X"80",
		X"A0",X"7F",X"00",X"CD",X"7F",X"FF",X"CC",X"7F",X"00",X"CD",X"7F",X"FF",X"8C",X"BF",X"14",X"80",
		X"A0",X"7F",X"00",X"CD",X"1F",X"0E",X"5F",X"0A",X"9F",X"01",X"71",X"71",X"71",X"71",X"B1",X"5F",
		X"09",X"7F",X"FF",X"9F",X"00",X"88",X"88",X"86",X"86",X"85",X"85",X"83",X"83",X"A1",X"A3",X"7F",
		X"00",X"BF",X"01",X"85",X"BF",X"01",X"85",X"7F",X"FF",X"BF",X"01",X"A5",X"88",X"88",X"86",X"86",
		X"85",X"85",X"83",X"83",X"A1",X"A3",X"7F",X"00",X"BF",X"05",X"81",X"BF",X"05",X"81",X"7F",X"FF",
		X"BF",X"05",X"A1",X"88",X"88",X"86",X"86",X"85",X"85",X"83",X"83",X"A1",X"A3",X"BF",X"04",X"7F",
		X"00",X"85",X"7F",X"FF",X"A5",X"80",X"88",X"88",X"86",X"86",X"85",X"85",X"83",X"83",X"BF",X"04",
		X"81",X"1F",X"08",X"8C",X"1F",X"0E",X"81",X"83",X"BF",X"04",X"7F",X"00",X"A1",X"7F",X"FF",X"A1",
		X"7F",X"00",X"A8",X"7F",X"FF",X"A8",X"7F",X"00",X"AA",X"7F",X"FF",X"AA",X"BF",X"01",X"8C",X"BF",
		X"01",X"8A",X"BF",X"01",X"88",X"BF",X"01",X"8A",X"BF",X"01",X"7F",X"00",X"AC",X"7F",X"FF",X"AC",
		X"7F",X"00",X"B1",X"7F",X"FF",X"B1",X"7F",X"00",X"AC",X"7F",X"FF",X"AC",X"BF",X"09",X"8D",X"BF",
		X"09",X"8C",X"BF",X"09",X"8A",X"BF",X"09",X"88",X"BF",X"05",X"7F",X"00",X"A6",X"7F",X"FF",X"BF",
		X"03",X"A6",X"7F",X"00",X"A8",X"7F",X"FF",X"A8",X"7F",X"00",X"AA",X"7F",X"FF",X"AA",X"BF",X"0A",
		X"8C",X"8A",X"88",X"8A",X"BF",X"01",X"7F",X"00",X"AC",X"7F",X"FF",X"AC",X"BF",X"08",X"7F",X"00",
		X"B1",X"7F",X"FF",X"BF",X"03",X"B1",X"BF",X"08",X"7F",X"00",X"AD",X"7F",X"FF",X"BF",X"03",X"AD",
		X"BF",X"08",X"8A",X"88",X"BF",X"08",X"86",X"83",X"BF",X"03",X"7F",X"00",X"A5",X"7F",X"FF",X"BF",
		X"03",X"85",X"5F",X"0A",X"7F",X"FE",X"9F",X"02",X"61",X"61",X"81",X"81",X"81",X"61",X"61",X"81",
		X"81",X"81",X"61",X"61",X"81",X"81",X"61",X"81",X"61",X"81",X"81",X"BF",X"12",X"A1",X"FF",X"3F",
		X"16",X"1F",X"08",X"5F",X"09",X"7F",X"00",X"C7",X"7F",X"FF",X"C6",X"7F",X"00",X"C7",X"7F",X"FF",
		X"C6",X"7F",X"00",X"C7",X"7F",X"FF",X"C6",X"7F",X"00",X"C7",X"7F",X"FF",X"C6",X"1F",X"02",X"5F",
		X"08",X"8D",X"60",X"6D",X"2F",X"2F",X"2F",X"2F",X"91",X"74",X"8D",X"60",X"6D",X"2F",X"2F",X"2F",
		X"2F",X"91",X"74",X"8D",X"60",X"6D",X"2F",X"2F",X"2F",X"2F",X"91",X"74",X"94",X"88",X"8A",X"8C",
		X"8D",X"60",X"6D",X"2F",X"2F",X"2F",X"2F",X"91",X"74",X"8D",X"60",X"6D",X"2F",X"2F",X"2F",X"2F",
		X"91",X"74",X"8D",X"60",X"6D",X"2F",X"2F",X"2F",X"2F",X"91",X"74",X"94",X"92",X"91",X"8F",X"8D",
		X"60",X"6D",X"2F",X"2F",X"2F",X"2F",X"91",X"74",X"8D",X"60",X"6D",X"2F",X"2F",X"2F",X"2F",X"91",
		X"74",X"8D",X"60",X"6D",X"2F",X"2F",X"2F",X"2F",X"91",X"74",X"94",X"88",X"8A",X"8C",X"8D",X"60",
		X"6D",X"2F",X"2F",X"2F",X"2F",X"91",X"74",X"8D",X"60",X"6D",X"2F",X"2F",X"2F",X"2F",X"91",X"74",
		X"8D",X"60",X"6D",X"2F",X"2F",X"2F",X"2F",X"91",X"74",X"8D",X"8C",X"AD",X"1F",X"0E",X"5F",X"09",
		X"7F",X"00",X"A5",X"7F",X"FF",X"A5",X"7F",X"00",X"A6",X"7F",X"FF",X"A6",X"88",X"86",X"85",X"86",
		X"7F",X"00",X"88",X"7F",X"FF",X"A8",X"80",X"7F",X"00",X"AD",X"7F",X"FF",X"AD",X"7F",X"00",X"A8",
		X"7F",X"FF",X"A8",X"8A",X"88",X"86",X"85",X"7F",X"00",X"83",X"7F",X"FF",X"A3",X"80",X"7F",X"00",
		X"A5",X"7F",X"FF",X"A5",X"7F",X"00",X"A6",X"7F",X"FF",X"A6",X"88",X"86",X"85",X"86",X"7F",X"00",
		X"88",X"7F",X"FF",X"A8",X"80",X"7F",X"00",X"AD",X"7F",X"FF",X"AD",X"7F",X"00",X"A8",X"7F",X"FF",
		X"A8",X"86",X"85",X"83",X"1F",X"08",X"8C",X"1F",X"0E",X"7F",X"00",X"AD",X"7F",X"FF",X"AD",X"FF",
		X"FF",X"1F",X"0E",X"3F",X"15",X"5F",X"09",X"BA",X"D2",X"C6",X"D2",X"BF",X"C4",X"F3",X"F3",X"CC",
		X"BE",X"C5",X"CF",X"D2",X"C6",X"F3",X"F3",X"CA",X"CF",X"CE",X"C4",X"C5",X"F3",X"F3",X"D2",X"C1",
		X"D0",X"D2",X"CF",X"CA",X"D2",X"F3",X"F3",X"DA",X"DA",X"DA",X"F3",X"F3",X"D0",X"C4",X"C3",X"BA",
		X"C1",X"CA",X"CC",X"CB",X"BF",X"F3",X"C8",X"C4",X"C5",X"D2",X"C6",X"CA",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
