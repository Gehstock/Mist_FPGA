library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_PGM is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_PGM is
	type rom is array(0 to  24575) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"F3",X"C3",X"69",X"00",X"FF",X"FF",X"FF",X"C3",X"FF",X"04",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C3",X"E0",X"05",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"EC",X"05",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C3",X"FF",X"05",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C3",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"DA",X"0A",X"AF",X"21",X"00",X"A8",X"06",X"08",X"77",
		X"23",X"10",X"FC",X"3E",X"9B",X"32",X"03",X"98",X"3A",X"00",X"98",X"CB",X"47",X"CA",X"00",X"04",
		X"21",X"00",X"88",X"11",X"00",X"8C",X"FD",X"21",X"8D",X"00",X"C3",X"52",X"01",X"FD",X"21",X"94",
		X"00",X"C3",X"2F",X"02",X"21",X"9A",X"00",X"C3",X"62",X"02",X"52",X"41",X"4D",X"20",X"31",X"47",
		X"48",X"4A",X"4B",X"00",X"21",X"00",X"80",X"11",X"00",X"88",X"FD",X"21",X"B1",X"00",X"C3",X"52",
		X"01",X"21",X"B7",X"00",X"C3",X"62",X"02",X"32",X"43",X"20",X"52",X"4F",X"4D",X"20",X"20",X"20",
		X"00",X"21",X"00",X"00",X"DD",X"21",X"CB",X"00",X"C3",X"3A",X"01",X"21",X"D1",X"00",X"C3",X"62",
		X"02",X"32",X"45",X"00",X"21",X"00",X"10",X"DD",X"21",X"DE",X"00",X"C3",X"3A",X"01",X"21",X"E4",
		X"00",X"C3",X"62",X"02",X"32",X"46",X"00",X"21",X"00",X"20",X"DD",X"21",X"F1",X"00",X"C3",X"3A",
		X"01",X"21",X"F7",X"00",X"C3",X"62",X"02",X"32",X"48",X"00",X"21",X"00",X"30",X"DD",X"21",X"04",
		X"01",X"C3",X"3A",X"01",X"21",X"0A",X"01",X"C3",X"62",X"02",X"32",X"4A",X"00",X"21",X"00",X"40",
		X"DD",X"21",X"17",X"01",X"C3",X"3A",X"01",X"21",X"1D",X"01",X"C3",X"62",X"02",X"32",X"4C",X"00",
		X"21",X"00",X"50",X"DD",X"21",X"2A",X"01",X"C3",X"3A",X"01",X"21",X"30",X"01",X"C3",X"62",X"02",
		X"20",X"20",X"20",X"20",X"20",X"20",X"00",X"C3",X"E7",X"19",X"01",X"00",X"10",X"AF",X"86",X"23",
		X"0D",X"C2",X"3E",X"01",X"08",X"3A",X"00",X"70",X"08",X"10",X"F3",X"FE",X"FF",X"C2",X"83",X"02",
		X"DD",X"E9",X"DD",X"21",X"59",X"01",X"C3",X"99",X"01",X"44",X"4D",X"36",X"00",X"23",X"7D",X"BB",
		X"C2",X"5B",X"01",X"08",X"3A",X"00",X"B0",X"08",X"7C",X"BA",X"C2",X"5B",X"01",X"69",X"60",X"01",
		X"55",X"00",X"DD",X"21",X"79",X"01",X"C3",X"AA",X"01",X"01",X"AA",X"55",X"DD",X"21",X"83",X"01",
		X"C3",X"EC",X"01",X"01",X"FF",X"AA",X"DD",X"21",X"8D",X"01",X"C3",X"AA",X"01",X"01",X"00",X"FF",
		X"DD",X"21",X"97",X"01",X"C3",X"EC",X"01",X"FD",X"E9",X"06",X"00",X"70",X"7E",X"B8",X"C2",X"89",
		X"02",X"08",X"3A",X"00",X"B0",X"08",X"10",X"F3",X"DD",X"E9",X"08",X"3A",X"00",X"B0",X"08",X"7C",
		X"D9",X"67",X"D9",X"7D",X"D9",X"6F",X"D9",X"7B",X"D9",X"5F",X"D9",X"7A",X"D9",X"57",X"D9",X"7E",
		X"A8",X"C2",X"89",X"02",X"71",X"7E",X"A9",X"C2",X"89",X"02",X"23",X"7D",X"BB",X"C2",X"BF",X"01",
		X"08",X"3A",X"00",X"B0",X"08",X"7C",X"BA",X"C2",X"BF",X"01",X"D9",X"7C",X"D9",X"67",X"D9",X"7D",
		X"D9",X"6F",X"D9",X"7B",X"D9",X"5F",X"D9",X"7A",X"D9",X"57",X"DD",X"E9",X"08",X"3A",X"00",X"B0",
		X"08",X"7C",X"D9",X"67",X"D9",X"7D",X"D9",X"6F",X"D9",X"7B",X"D9",X"5F",X"D9",X"7A",X"D9",X"57",
		X"D9",X"EB",X"2B",X"7E",X"A8",X"C2",X"89",X"02",X"71",X"7E",X"A9",X"C2",X"89",X"02",X"08",X"3A",
		X"00",X"B0",X"08",X"7D",X"BB",X"C2",X"02",X"02",X"7C",X"BA",X"C2",X"02",X"02",X"D9",X"7C",X"D9",
		X"67",X"D9",X"7D",X"D9",X"6F",X"D9",X"7B",X"D9",X"5F",X"D9",X"7A",X"D9",X"57",X"DD",X"E9",X"21",
		X"00",X"88",X"11",X"00",X"8C",X"06",X"10",X"DD",X"21",X"3E",X"02",X"C3",X"4F",X"02",X"21",X"00",
		X"90",X"11",X"00",X"94",X"06",X"00",X"DD",X"21",X"4D",X"02",X"C3",X"4F",X"02",X"FD",X"E9",X"70",
		X"23",X"7D",X"BB",X"C2",X"4F",X"02",X"08",X"3A",X"00",X"B0",X"08",X"7C",X"BA",X"C2",X"4F",X"02",
		X"DD",X"E9",X"EB",X"21",X"6E",X"8B",X"1A",X"B7",X"CA",X"80",X"02",X"D6",X"30",X"F2",X"72",X"02",
		X"3E",X"10",X"77",X"08",X"3A",X"00",X"B0",X"08",X"01",X"E0",X"FF",X"09",X"13",X"C3",X"66",X"02",
		X"EB",X"23",X"E9",X"3A",X"00",X"B0",X"C3",X"83",X"02",X"3A",X"00",X"B0",X"C3",X"89",X"02",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"31",X"80",X"80",X"F5",X"3A",X"00",X"B0",X"F1",X"CD",X"82",X"05",X"F5",X"3A",X"00",X"B0",X"F1",
		X"D7",X"00",X"E7",X"04",X"04",X"01",X"E7",X"04",X"08",X"02",X"E7",X"04",X"0C",X"03",X"E7",X"04",
		X"10",X"04",X"3E",X"9B",X"32",X"03",X"98",X"3E",X"88",X"32",X"03",X"A0",X"F5",X"3A",X"00",X"B0",
		X"F1",X"3E",X"10",X"32",X"02",X"98",X"3E",X"00",X"32",X"02",X"98",X"CF",X"68",X"40",X"50",X"4F",
		X"52",X"54",X"20",X"41",X"00",X"21",X"50",X"40",X"CD",X"BF",X"04",X"3A",X"00",X"98",X"CD",X"A7",
		X"04",X"CF",X"68",X"60",X"50",X"4F",X"52",X"54",X"20",X"42",X"00",X"21",X"70",X"40",X"CD",X"BF",
		X"04",X"3A",X"01",X"98",X"CD",X"A7",X"04",X"CF",X"68",X"80",X"50",X"4F",X"52",X"54",X"20",X"43",
		X"00",X"21",X"90",X"40",X"CD",X"BF",X"04",X"3A",X"02",X"98",X"CD",X"A7",X"04",X"CF",X"40",X"A8",
		X"37",X"20",X"36",X"20",X"35",X"20",X"34",X"20",X"33",X"20",X"32",X"20",X"31",X"20",X"30",X"00",
		X"CF",X"50",X"B0",X"42",X"49",X"54",X"20",X"4E",X"55",X"4D",X"42",X"45",X"52",X"53",X"00",X"2E",
		X"00",X"2D",X"20",X"FD",X"C3",X"2C",X"04",X"06",X"08",X"07",X"F5",X"E6",X"01",X"F6",X"30",X"CD",
		X"6A",X"05",X"AF",X"CD",X"6A",X"05",X"F5",X"3A",X"00",X"B0",X"F1",X"F1",X"10",X"EB",X"C9",X"F5",
		X"AF",X"C3",X"C4",X"04",X"94",X"3D",X"67",X"CB",X"3C",X"CB",X"3C",X"CB",X"3C",X"CB",X"3C",X"CB",
		X"1D",X"CB",X"3C",X"CB",X"1D",X"CB",X"3C",X"CB",X"1D",X"D5",X"11",X"00",X"88",X"19",X"D1",X"F1",
		X"C9",X"D5",X"11",X"00",X"88",X"B7",X"ED",X"52",X"CB",X"25",X"CB",X"14",X"CB",X"25",X"CB",X"14",
		X"CB",X"25",X"CB",X"14",X"7C",X"2F",X"67",X"CB",X"24",X"CB",X"24",X"CB",X"24",X"D1",X"C9",X"E3",
		X"F5",X"C5",X"D5",X"56",X"23",X"5E",X"23",X"EB",X"CD",X"BF",X"04",X"1A",X"13",X"B7",X"CA",X"17",
		X"05",X"CD",X"6A",X"05",X"C3",X"0B",X"05",X"EB",X"D1",X"C1",X"F1",X"E3",X"C9",X"0E",X"03",X"C3",
		X"29",X"05",X"0E",X"00",X"C3",X"29",X"05",X"0E",X"01",X"F5",X"C5",X"D5",X"E5",X"CD",X"BF",X"04",
		X"78",X"3D",X"20",X"02",X"CB",X"81",X"1A",X"CB",X"40",X"20",X"05",X"07",X"07",X"07",X"07",X"1B",
		X"13",X"E6",X"0F",X"C2",X"55",X"05",X"CB",X"41",X"CA",X"57",X"05",X"3E",X"20",X"CB",X"49",X"C2",
		X"63",X"05",X"C3",X"60",X"05",X"CB",X"81",X"C6",X"30",X"FE",X"3A",X"DA",X"60",X"05",X"C6",X"07",
		X"CD",X"6A",X"05",X"10",X"CB",X"E1",X"D1",X"C1",X"F1",X"C9",X"C5",X"D6",X"30",X"F2",X"72",X"05",
		X"3E",X"10",X"77",X"01",X"E0",X"FF",X"09",X"7C",X"FE",X"88",X"30",X"04",X"01",X"00",X"04",X"09",
		X"C1",X"C9",X"F5",X"C5",X"E5",X"D5",X"3E",X"00",X"32",X"40",X"86",X"06",X"B4",X"21",X"79",X"85",
		X"36",X"00",X"23",X"10",X"FB",X"21",X"00",X"88",X"0E",X"04",X"3E",X"10",X"CD",X"B8",X"05",X"21",
		X"00",X"90",X"0E",X"01",X"CD",X"B7",X"05",X"3E",X"00",X"32",X"03",X"A8",X"32",X"05",X"A8",X"32",
		X"04",X"A8",X"D1",X"E1",X"C1",X"F1",X"C9",X"AF",X"06",X"00",X"77",X"23",X"10",X"FC",X"0D",X"20",
		X"F9",X"C9",X"F5",X"C5",X"D5",X"E5",X"50",X"E5",X"CD",X"BF",X"04",X"3E",X"20",X"CD",X"6A",X"05",
		X"10",X"F9",X"E1",X"7D",X"C6",X"08",X"6F",X"42",X"0D",X"20",X"EC",X"E1",X"D1",X"C1",X"F1",X"C9",
		X"E1",X"7E",X"23",X"E5",X"11",X"00",X"00",X"06",X"20",X"C3",X"09",X"06",X"E1",X"7E",X"23",X"E5",
		X"47",X"0F",X"0F",X"E6",X"3E",X"4F",X"78",X"06",X"00",X"21",X"01",X"90",X"09",X"77",X"C9",X"E1",
		X"46",X"23",X"5E",X"16",X"00",X"23",X"7E",X"23",X"E5",X"21",X"01",X"90",X"19",X"19",X"77",X"23",
		X"23",X"10",X"FB",X"C9",X"21",X"01",X"90",X"19",X"19",X"77",X"23",X"23",X"10",X"FB",X"C9",X"77",
		X"3C",X"23",X"77",X"3C",X"11",X"1F",X"00",X"19",X"77",X"3C",X"23",X"77",X"C9",X"DF",X"FC",X"CF",
		X"10",X"F8",X"3B",X"31",X"39",X"38",X"32",X"20",X"53",X"54",X"45",X"52",X"4E",X"20",X"45",X"4C",
		X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",X"43",X"00",X"C9",X"AF",
		X"32",X"54",X"85",X"3A",X"EE",X"80",X"B7",X"28",X"1E",X"DF",X"F2",X"CF",X"80",X"F0",X"20",X"43",
		X"52",X"45",X"44",X"49",X"54",X"53",X"5B",X"20",X"20",X"20",X"00",X"21",X"F0",X"C8",X"11",X"EE",
		X"80",X"06",X"02",X"CD",X"27",X"05",X"C9",X"DF",X"F6",X"CF",X"80",X"F0",X"49",X"4E",X"53",X"45",
		X"52",X"54",X"20",X"43",X"4F",X"49",X"4E",X"00",X"C9",X"AF",X"32",X"53",X"85",X"DF",X"0B",X"CF",
		X"20",X"00",X"31",X"53",X"54",X"00",X"21",X"08",X"10",X"11",X"2B",X"81",X"06",X"06",X"CD",X"27",
		X"05",X"CF",X"58",X"00",X"48",X"49",X"47",X"48",X"20",X"53",X"43",X"4F",X"52",X"45",X"00",X"21",
		X"08",X"68",X"11",X"EF",X"80",X"06",X"06",X"CD",X"27",X"05",X"3A",X"56",X"85",X"FE",X"02",X"C0",
		X"CF",X"D0",X"00",X"32",X"4E",X"44",X"00",X"21",X"08",X"C0",X"11",X"2E",X"81",X"06",X"06",X"CD",
		X"27",X"05",X"C9",X"DF",X"F9",X"3A",X"29",X"85",X"B7",X"C8",X"3D",X"C8",X"FE",X"08",X"38",X"02",
		X"3E",X"08",X"21",X"F8",X"18",X"E5",X"CD",X"BF",X"04",X"36",X"3C",X"E1",X"3D",X"C8",X"08",X"7C",
		X"C6",X"08",X"67",X"08",X"18",X"EF",X"C9",X"CF",X"58",X"D8",X"20",X"4C",X"45",X"56",X"45",X"4C",
		X"20",X"20",X"20",X"00",X"21",X"D8",X"88",X"11",X"2E",X"85",X"06",X"02",X"CD",X"27",X"05",X"C9",
		X"3A",X"EE",X"80",X"B7",X"C8",X"21",X"B8",X"00",X"01",X"05",X"20",X"CD",X"C2",X"05",X"E7",X"05",
		X"17",X"05",X"3A",X"EE",X"80",X"FE",X"01",X"20",X"41",X"CF",X"18",X"B8",X"50",X"55",X"53",X"48",
		X"20",X"31",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"53",X"54",X"41",X"52",X"54",X"20",
		X"42",X"55",X"54",X"54",X"4F",X"4E",X"00",X"CF",X"68",X"C8",X"5B",X"20",X"4F",X"52",X"20",X"5B",
		X"00",X"CF",X"30",X"D8",X"49",X"4E",X"53",X"45",X"52",X"54",X"20",X"41",X"4E",X"4F",X"54",X"48",
		X"45",X"52",X"20",X"43",X"4F",X"49",X"4E",X"00",X"18",X"34",X"CF",X"48",X"B8",X"50",X"55",X"53",
		X"48",X"20",X"31",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"00",X"CF",X"68",X"C8",X"5B",X"20",
		X"4F",X"52",X"20",X"5B",X"00",X"CF",X"28",X"D8",X"32",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",
		X"20",X"53",X"54",X"41",X"52",X"54",X"20",X"42",X"55",X"54",X"54",X"4F",X"4E",X"00",X"06",X"05",
		X"C5",X"E7",X"05",X"17",X"01",X"3E",X"02",X"CD",X"88",X"1A",X"E7",X"05",X"17",X"02",X"3E",X"02",
		X"CD",X"88",X"1A",X"E7",X"05",X"17",X"03",X"3E",X"02",X"CD",X"88",X"1A",X"E7",X"05",X"17",X"04",
		X"3E",X"02",X"CD",X"88",X"1A",X"E7",X"05",X"17",X"05",X"3E",X"02",X"CD",X"88",X"1A",X"E7",X"05",
		X"17",X"06",X"3E",X"02",X"CD",X"88",X"1A",X"E7",X"05",X"17",X"07",X"3E",X"02",X"CD",X"88",X"1A",
		X"E7",X"05",X"17",X"00",X"3E",X"02",X"CD",X"88",X"1A",X"C1",X"10",X"B4",X"C9",X"3A",X"2F",X"85",
		X"B7",X"28",X"1B",X"FE",X"08",X"38",X"02",X"3E",X"08",X"21",X"F8",X"60",X"E5",X"CD",X"BF",X"04",
		X"36",X"2C",X"E1",X"3D",X"28",X"0D",X"08",X"7C",X"C6",X"08",X"67",X"08",X"18",X"EE",X"21",X"F8",
		X"60",X"18",X"06",X"08",X"7C",X"C6",X"08",X"67",X"08",X"CD",X"BF",X"04",X"36",X"10",X"C9",X"F5",
		X"3A",X"55",X"85",X"B7",X"28",X"09",X"3A",X"01",X"98",X"E6",X"02",X"28",X"02",X"F1",X"C9",X"F1",
		X"F3",X"32",X"00",X"A0",X"AF",X"32",X"01",X"A0",X"E3",X"E3",X"3E",X"08",X"32",X"01",X"A0",X"FB",
		X"C9",X"61",X"D5",X"E5",X"ED",X"5B",X"4E",X"85",X"21",X"AA",X"AA",X"19",X"29",X"19",X"29",X"19",
		X"29",X"19",X"29",X"29",X"19",X"29",X"29",X"19",X"29",X"29",X"19",X"29",X"19",X"29",X"29",X"19",
		X"29",X"19",X"29",X"19",X"11",X"2F",X"6A",X"19",X"22",X"4E",X"85",X"7C",X"E1",X"D1",X"C9",X"FD",
		X"E1",X"DD",X"21",X"40",X"82",X"DD",X"CB",X"00",X"C6",X"DD",X"CB",X"00",X"CE",X"CD",X"80",X"09",
		X"31",X"90",X"80",X"FD",X"E9",X"FD",X"E1",X"DD",X"21",X"12",X"82",X"DD",X"CB",X"00",X"C6",X"DD",
		X"CB",X"00",X"CE",X"CD",X"80",X"09",X"31",X"B8",X"80",X"DD",X"21",X"9A",X"81",X"DD",X"CB",X"00",
		X"C6",X"CD",X"69",X"09",X"CD",X"94",X"09",X"FD",X"E9",X"C9",X"FD",X"E1",X"DD",X"21",X"12",X"82",
		X"DD",X"CB",X"00",X"C6",X"DD",X"CB",X"00",X"CE",X"CD",X"80",X"09",X"31",X"B8",X"80",X"DD",X"21",
		X"9A",X"81",X"DD",X"CB",X"00",X"C6",X"CD",X"69",X"09",X"CD",X"94",X"09",X"FD",X"E9",X"D9",X"21",
		X"A8",X"0A",X"CD",X"4E",X"09",X"D9",X"D0",X"CD",X"69",X"09",X"CD",X"94",X"09",X"37",X"C9",X"D9",
		X"21",X"B8",X"0A",X"CD",X"4E",X"09",X"D9",X"D0",X"CD",X"69",X"09",X"CD",X"94",X"09",X"37",X"C9",
		X"FD",X"E1",X"CD",X"3E",X"09",X"30",X"12",X"DD",X"CB",X"00",X"C6",X"DD",X"CB",X"00",X"CE",X"CD",
		X"80",X"09",X"CD",X"29",X"0A",X"CD",X"DF",X"08",X"37",X"FD",X"E9",X"FD",X"E1",X"CD",X"46",X"09",
		X"30",X"12",X"DD",X"CB",X"00",X"C6",X"DD",X"CB",X"00",X"CE",X"CD",X"80",X"09",X"CD",X"29",X"0A",
		X"CD",X"DF",X"08",X"37",X"FD",X"E9",X"E1",X"D9",X"21",X"C8",X"0A",X"CD",X"4E",X"09",X"D9",X"D2",
		X"3D",X"09",X"DD",X"22",X"DA",X"80",X"CD",X"80",X"09",X"CD",X"29",X"0A",X"37",X"E9",X"E1",X"D9",
		X"21",X"96",X"0A",X"C3",X"2B",X"09",X"E1",X"D9",X"21",X"A6",X"0A",X"C3",X"2B",X"09",X"E5",X"D1",
		X"7E",X"23",X"66",X"6F",X"B4",X"C8",X"7E",X"B7",X"28",X"06",X"13",X"13",X"D5",X"E1",X"18",X"F0",
		X"E5",X"DD",X"E1",X"DD",X"CB",X"00",X"C6",X"37",X"C9",X"D9",X"DD",X"E5",X"E1",X"DD",X"2A",X"DA",
		X"80",X"DD",X"75",X"01",X"DD",X"74",X"02",X"DD",X"CB",X"00",X"DE",X"E5",X"DD",X"E1",X"D9",X"C9",
		X"D9",X"DD",X"CB",X"00",X"CE",X"DD",X"E5",X"E1",X"22",X"DA",X"80",X"AF",X"06",X"0F",X"23",X"77",
		X"10",X"FC",X"D9",X"C9",X"D9",X"DD",X"E5",X"E1",X"22",X"D8",X"80",X"AF",X"06",X"0E",X"23",X"77",
		X"10",X"FC",X"D9",X"C9",X"21",X"00",X"00",X"39",X"31",X"68",X"80",X"FD",X"E5",X"FD",X"2A",X"DA",
		X"80",X"FD",X"22",X"DE",X"80",X"FD",X"75",X"0E",X"FD",X"74",X"0F",X"C9",X"21",X"00",X"00",X"39",
		X"31",X"68",X"80",X"DD",X"2A",X"DA",X"80",X"DD",X"75",X"0E",X"DD",X"74",X"0F",X"2A",X"DE",X"80",
		X"7C",X"B5",X"28",X"0C",X"DD",X"2A",X"DE",X"80",X"21",X"00",X"00",X"22",X"DE",X"80",X"18",X"04",
		X"DD",X"2A",X"DA",X"80",X"CD",X"F9",X"09",X"DD",X"CB",X"00",X"46",X"28",X"F7",X"DD",X"22",X"DA",
		X"80",X"DD",X"66",X"0F",X"DD",X"6E",X"0E",X"F9",X"C9",X"D9",X"01",X"2E",X"00",X"DD",X"09",X"DD",
		X"E5",X"E1",X"01",X"20",X"85",X"B7",X"ED",X"42",X"38",X"04",X"DD",X"21",X"12",X"82",X"D9",X"C9",
		X"DD",X"2A",X"DA",X"80",X"DD",X"77",X"03",X"DD",X"CB",X"00",X"EE",X"CD",X"BC",X"09",X"DD",X"2A",
		X"DA",X"80",X"DD",X"CB",X"00",X"6E",X"20",X"F3",X"C9",X"D9",X"D1",X"01",X"2E",X"00",X"DD",X"E5",
		X"E1",X"09",X"F9",X"D5",X"D9",X"C9",X"CD",X"46",X"0A",X"D9",X"2A",X"DA",X"80",X"06",X"10",X"AF",
		X"77",X"23",X"10",X"FC",X"D9",X"C9",X"DD",X"2A",X"DA",X"80",X"DD",X"CB",X"00",X"5E",X"C8",X"DD",
		X"CB",X"00",X"9E",X"D9",X"DD",X"6E",X"01",X"DD",X"66",X"02",X"06",X"0F",X"AF",X"77",X"23",X"10",
		X"FC",X"DD",X"77",X"01",X"DD",X"77",X"01",X"D9",X"C9",X"CD",X"FE",X"0B",X"DD",X"21",X"12",X"82",
		X"AF",X"DD",X"77",X"00",X"DD",X"21",X"6E",X"82",X"DD",X"77",X"00",X"CD",X"F9",X"09",X"30",X"02",
		X"18",X"F6",X"DD",X"21",X"31",X"81",X"11",X"0F",X"00",X"06",X"0F",X"DD",X"77",X"00",X"DD",X"19",
		X"10",X"F9",X"CD",X"04",X"0C",X"C9",X"DE",X"83",X"0C",X"84",X"3A",X"84",X"68",X"84",X"96",X"84",
		X"C4",X"84",X"F2",X"84",X"00",X"00",X"00",X"00",X"31",X"81",X"40",X"81",X"4F",X"81",X"5E",X"81",
		X"6D",X"81",X"7C",X"81",X"8B",X"81",X"00",X"00",X"A9",X"81",X"B8",X"81",X"C7",X"81",X"D6",X"81",
		X"E5",X"81",X"F4",X"81",X"03",X"82",X"00",X"00",X"6E",X"82",X"9C",X"82",X"CA",X"82",X"F8",X"82",
		X"26",X"83",X"54",X"83",X"82",X"83",X"B0",X"83",X"00",X"00",X"F5",X"3A",X"00",X"B0",X"AF",X"32",
		X"01",X"A8",X"3C",X"32",X"01",X"A8",X"3A",X"E2",X"80",X"CB",X"0F",X"32",X"E2",X"80",X"DA",X"D8",
		X"0B",X"3A",X"E3",X"80",X"B7",X"C2",X"D6",X"0B",X"3C",X"32",X"E3",X"80",X"ED",X"73",X"DC",X"80",
		X"31",X"40",X"80",X"08",X"F5",X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",X"D9",X"C5",X"D5",X"E5",
		X"21",X"38",X"86",X"34",X"3A",X"38",X"86",X"FE",X"1E",X"20",X"09",X"36",X"00",X"2A",X"39",X"86",
		X"23",X"22",X"39",X"86",X"21",X"31",X"81",X"11",X"40",X"90",X"06",X"08",X"C5",X"CB",X"46",X"CC",
		X"B3",X"0F",X"01",X"06",X"00",X"09",X"7E",X"12",X"23",X"13",X"7E",X"12",X"23",X"13",X"7E",X"12",
		X"23",X"23",X"23",X"23",X"13",X"7E",X"12",X"23",X"23",X"23",X"13",X"C1",X"10",X"DE",X"21",X"A9",
		X"81",X"11",X"61",X"90",X"06",X"07",X"C5",X"E5",X"DD",X"E1",X"CB",X"46",X"CC",X"B3",X"0F",X"01",
		X"06",X"00",X"09",X"3A",X"59",X"85",X"FE",X"02",X"20",X"16",X"3A",X"02",X"98",X"E6",X"08",X"20",
		X"0F",X"7E",X"C6",X"06",X"12",X"01",X"06",X"00",X"09",X"13",X"13",X"7E",X"C6",X"04",X"18",X"0E",
		X"7E",X"C6",X"08",X"12",X"01",X"06",X"00",X"09",X"13",X"13",X"7E",X"2F",X"C6",X"F1",X"12",X"13",
		X"13",X"23",X"23",X"23",X"C1",X"10",X"BF",X"CD",X"0A",X"32",X"CD",X"4E",X"12",X"21",X"12",X"82",
		X"06",X"11",X"C5",X"46",X"CB",X"40",X"C4",X"0A",X"0C",X"CB",X"58",X"C4",X"59",X"0C",X"11",X"2E",
		X"00",X"19",X"C1",X"10",X"ED",X"CD",X"D8",X"0E",X"CD",X"80",X"0F",X"CD",X"D2",X"0F",X"CD",X"F5",
		X"10",X"E1",X"D1",X"C1",X"D9",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"F1",X"08",X"ED",X"7B",
		X"DC",X"80",X"AF",X"32",X"E3",X"80",X"F1",X"C9",X"ED",X"73",X"E0",X"80",X"31",X"D8",X"80",X"C5",
		X"D5",X"E5",X"DD",X"E5",X"08",X"D9",X"F5",X"C5",X"D5",X"E5",X"CD",X"F5",X"10",X"E1",X"D1",X"C1",
		X"F1",X"D9",X"08",X"DD",X"E1",X"E1",X"D1",X"C1",X"ED",X"7B",X"E0",X"80",X"F1",X"C9",X"3E",X"FF",
		X"32",X"E2",X"80",X"C9",X"3E",X"55",X"32",X"E2",X"80",X"C9",X"E5",X"CB",X"48",X"CA",X"56",X"0C",
		X"23",X"5E",X"23",X"56",X"D5",X"FD",X"E1",X"23",X"CB",X"68",X"28",X"05",X"35",X"20",X"02",X"CB",
		X"A8",X"23",X"CB",X"60",X"28",X"2C",X"35",X"20",X"29",X"CB",X"F8",X"23",X"5E",X"23",X"56",X"13",
		X"13",X"13",X"13",X"13",X"1A",X"B7",X"C2",X"4A",X"0C",X"13",X"1A",X"B7",X"C2",X"43",X"0C",X"CB",
		X"A0",X"CB",X"B8",X"EB",X"23",X"7E",X"23",X"66",X"6F",X"EB",X"72",X"2B",X"73",X"13",X"13",X"1A",
		X"2B",X"77",X"CB",X"50",X"28",X"00",X"E1",X"70",X"C9",X"CB",X"48",X"C8",X"E5",X"DD",X"E1",X"E5",
		X"FD",X"CB",X"00",X"66",X"28",X"17",X"DD",X"7E",X"08",X"C6",X"08",X"67",X"DD",X"7E",X"0A",X"C6",
		X"08",X"6F",X"CD",X"BF",X"04",X"FD",X"7E",X"0E",X"77",X"FD",X"CB",X"00",X"A6",X"E1",X"CB",X"78",
		X"28",X"14",X"CB",X"BE",X"DD",X"66",X"06",X"DD",X"6E",X"05",X"23",X"23",X"23",X"7E",X"FD",X"77",
		X"07",X"23",X"7E",X"FD",X"77",X"08",X"FD",X"CB",X"00",X"4E",X"28",X"09",X"FD",X"35",X"01",X"20",
		X"04",X"FD",X"CB",X"00",X"8E",X"FD",X"CB",X"00",X"56",X"28",X"09",X"FD",X"35",X"02",X"20",X"04",
		X"FD",X"CB",X"00",X"96",X"CB",X"50",X"28",X"49",X"DD",X"7E",X"07",X"FD",X"77",X"05",X"DD",X"7E",
		X"08",X"FD",X"77",X"06",X"DD",X"7E",X"09",X"FD",X"77",X"0B",X"DD",X"7E",X"0A",X"FD",X"77",X"0C",
		X"FD",X"E5",X"E1",X"23",X"23",X"23",X"5E",X"23",X"56",X"23",X"4E",X"23",X"46",X"EB",X"09",X"EB",
		X"DD",X"72",X"08",X"DD",X"73",X"07",X"2B",X"73",X"23",X"72",X"23",X"23",X"23",X"5E",X"23",X"56",
		X"23",X"4E",X"23",X"46",X"EB",X"09",X"EB",X"DD",X"72",X"0A",X"DD",X"73",X"09",X"2B",X"73",X"23",
		X"72",X"DD",X"7E",X"08",X"C6",X"08",X"67",X"DD",X"7E",X"0A",X"C6",X"08",X"6F",X"CD",X"BF",X"04",
		X"7E",X"FD",X"77",X"0D",X"CD",X"1A",X"0D",X"C3",X"D4",X"0E",X"FD",X"CB",X"00",X"6E",X"C8",X"3A",
		X"32",X"85",X"B7",X"28",X"29",X"FE",X"01",X"28",X"0F",X"FE",X"02",X"28",X"16",X"FD",X"7E",X"0D",
		X"FE",X"70",X"D8",X"FE",X"74",X"D0",X"18",X"1F",X"FD",X"7E",X"0D",X"FE",X"88",X"D8",X"FE",X"8C",
		X"D0",X"18",X"14",X"FD",X"7E",X"0D",X"FE",X"60",X"D8",X"FE",X"64",X"D0",X"18",X"09",X"FD",X"7E",
		X"0D",X"FE",X"38",X"D8",X"FE",X"3C",X"D0",X"FD",X"7E",X"09",X"B7",X"20",X"15",X"FD",X"7E",X"0A",
		X"B7",X"20",X"0F",X"FD",X"7E",X"03",X"B7",X"C2",X"09",X"0E",X"FD",X"7E",X"04",X"B7",X"C2",X"09",
		X"0E",X"C9",X"E5",X"FD",X"CB",X"0A",X"7E",X"20",X"48",X"23",X"3A",X"32",X"85",X"B7",X"28",X"29",
		X"FE",X"01",X"28",X"0F",X"FE",X"02",X"28",X"16",X"7E",X"FE",X"70",X"38",X"27",X"FE",X"74",X"30",
		X"23",X"18",X"E6",X"7E",X"FE",X"88",X"38",X"1C",X"FE",X"8C",X"30",X"18",X"18",X"DB",X"7E",X"FE",
		X"60",X"38",X"11",X"FE",X"64",X"30",X"0D",X"18",X"D0",X"7E",X"FE",X"38",X"38",X"06",X"FE",X"3C",
		X"30",X"02",X"18",X"C5",X"FE",X"3D",X"DA",X"A4",X"0E",X"FE",X"44",X"D2",X"A4",X"0E",X"C3",X"D2",
		X"0E",X"2B",X"3A",X"32",X"85",X"B7",X"28",X"29",X"FE",X"01",X"28",X"1A",X"FE",X"02",X"28",X"0B",
		X"7E",X"FE",X"70",X"38",X"27",X"FE",X"74",X"30",X"23",X"18",X"E6",X"7E",X"FE",X"60",X"38",X"1C",
		X"FE",X"64",X"30",X"18",X"18",X"DB",X"7E",X"FE",X"88",X"38",X"11",X"FE",X"8C",X"30",X"0D",X"18",
		X"D0",X"7E",X"FE",X"38",X"38",X"06",X"FE",X"3C",X"30",X"02",X"18",X"C5",X"FE",X"3D",X"DA",X"A4",
		X"0E",X"FE",X"44",X"D2",X"A4",X"0E",X"C3",X"D2",X"0E",X"FD",X"CB",X"04",X"7E",X"28",X"49",X"11",
		X"20",X"00",X"E5",X"19",X"3A",X"32",X"85",X"B7",X"28",X"29",X"FE",X"01",X"28",X"1A",X"FE",X"02",
		X"28",X"0B",X"7E",X"FE",X"70",X"38",X"27",X"FE",X"74",X"30",X"23",X"18",X"E6",X"7E",X"FE",X"60",
		X"38",X"1C",X"FE",X"64",X"30",X"18",X"18",X"DB",X"7E",X"FE",X"88",X"38",X"11",X"FE",X"8C",X"30",
		X"0D",X"18",X"D0",X"7E",X"FE",X"38",X"38",X"06",X"FE",X"3C",X"30",X"02",X"18",X"C5",X"FE",X"3D",
		X"38",X"52",X"FE",X"44",X"30",X"4E",X"18",X"7A",X"11",X"20",X"00",X"E5",X"37",X"3F",X"ED",X"52",
		X"3A",X"32",X"85",X"B7",X"28",X"29",X"FE",X"01",X"28",X"0F",X"FE",X"02",X"28",X"16",X"7E",X"FE",
		X"70",X"38",X"27",X"FE",X"74",X"30",X"23",X"18",X"E3",X"7E",X"FE",X"88",X"38",X"1C",X"FE",X"8C",
		X"30",X"18",X"18",X"D8",X"7E",X"FE",X"60",X"38",X"11",X"FE",X"64",X"30",X"0D",X"18",X"CD",X"7E",
		X"FE",X"38",X"38",X"06",X"FE",X"3C",X"30",X"02",X"18",X"C2",X"FE",X"3D",X"38",X"06",X"FE",X"44",
		X"30",X"02",X"18",X"2E",X"3A",X"32",X"85",X"B7",X"28",X"20",X"FE",X"01",X"28",X"14",X"FE",X"02",
		X"28",X"08",X"3E",X"70",X"77",X"E1",X"3E",X"10",X"77",X"C9",X"3E",X"60",X"77",X"E1",X"3E",X"10",
		X"77",X"C9",X"3E",X"88",X"77",X"E1",X"3E",X"10",X"77",X"C9",X"3E",X"38",X"77",X"E1",X"3E",X"10",
		X"77",X"C9",X"E1",X"C9",X"DD",X"E5",X"E1",X"C9",X"DD",X"21",X"DE",X"83",X"06",X"07",X"DD",X"CB",
		X"00",X"46",X"C4",X"ED",X"0E",X"11",X"2E",X"00",X"DD",X"19",X"10",X"F2",X"C9",X"DD",X"7E",X"0D",
		X"B7",X"C0",X"DD",X"66",X"02",X"DD",X"6E",X"01",X"E5",X"FD",X"E1",X"3A",X"32",X"85",X"B7",X"28",
		X"32",X"FE",X"01",X"28",X"20",X"FE",X"02",X"28",X"0E",X"FD",X"7E",X"0D",X"D9",X"FE",X"70",X"38",
		X"6D",X"FE",X"74",X"30",X"69",X"18",X"28",X"FD",X"7E",X"0D",X"D9",X"FE",X"60",X"38",X"5F",X"FE",
		X"64",X"30",X"5B",X"18",X"1A",X"FD",X"7E",X"0D",X"D9",X"FE",X"88",X"38",X"51",X"FE",X"8C",X"30",
		X"4D",X"18",X"0C",X"FD",X"7E",X"0D",X"D9",X"FE",X"38",X"38",X"43",X"FE",X"3C",X"30",X"3F",X"DD",
		X"36",X"0D",X"FF",X"01",X"02",X"01",X"CD",X"57",X"1F",X"DD",X"7E",X"08",X"C6",X"08",X"67",X"DD",
		X"7E",X"0A",X"C6",X"08",X"6F",X"CD",X"BF",X"04",X"36",X"2E",X"EB",X"21",X"79",X"85",X"CD",X"42",
		X"08",X"E6",X"03",X"20",X"01",X"3C",X"CD",X"1F",X"08",X"06",X"59",X"4E",X"23",X"7E",X"23",X"B1",
		X"20",X"07",X"2B",X"2B",X"73",X"23",X"72",X"18",X"05",X"10",X"F0",X"EB",X"36",X"10",X"D9",X"C9",
		X"21",X"78",X"85",X"35",X"7E",X"B7",X"C0",X"36",X"05",X"21",X"79",X"85",X"06",X"5A",X"5E",X"23",
		X"56",X"23",X"7A",X"B3",X"28",X"1A",X"1A",X"FE",X"2E",X"38",X"0A",X"FE",X"37",X"28",X"06",X"30",
		X"04",X"3C",X"12",X"18",X"0B",X"3E",X"10",X"12",X"2B",X"2B",X"36",X"00",X"23",X"36",X"00",X"23",
		X"10",X"DC",X"C9",X"AF",X"E5",X"DD",X"E1",X"DD",X"77",X"06",X"DD",X"77",X"0C",X"C9",X"7A",X"2F",
		X"57",X"7B",X"2F",X"5F",X"13",X"C9",X"78",X"2F",X"47",X"79",X"2F",X"4F",X"03",X"C9",X"00",X"00",
		X"00",X"00",X"DD",X"21",X"12",X"82",X"FD",X"21",X"6E",X"82",X"3E",X"08",X"6F",X"DD",X"4E",X"0A",
		X"D9",X"3E",X"08",X"6F",X"DD",X"4E",X"08",X"06",X"08",X"FD",X"7E",X"00",X"E6",X"41",X"EE",X"41",
		X"20",X"3B",X"FD",X"56",X"06",X"FD",X"5E",X"05",X"1A",X"67",X"13",X"1A",X"D9",X"85",X"1F",X"67",
		X"FD",X"7E",X"0A",X"91",X"30",X"02",X"ED",X"44",X"BC",X"D9",X"30",X"21",X"7C",X"85",X"1F",X"67",
		X"FD",X"7E",X"08",X"91",X"30",X"02",X"ED",X"44",X"BC",X"30",X"12",X"DD",X"7E",X"0D",X"FD",X"B6",
		X"0C",X"DD",X"77",X"0D",X"FD",X"7E",X"0D",X"DD",X"B6",X"0C",X"FD",X"77",X"0D",X"11",X"2E",X"00",
		X"FD",X"19",X"10",X"B5",X"DD",X"21",X"DE",X"83",X"CD",X"5B",X"10",X"DD",X"21",X"0C",X"84",X"CD",
		X"5B",X"10",X"DD",X"21",X"3A",X"84",X"CD",X"5B",X"10",X"DD",X"21",X"68",X"84",X"CD",X"5B",X"10",
		X"DD",X"21",X"96",X"84",X"CD",X"5B",X"10",X"DD",X"21",X"C4",X"84",X"DD",X"7E",X"00",X"E6",X"41",
		X"EE",X"41",X"C0",X"FD",X"21",X"6E",X"82",X"3E",X"02",X"6F",X"DD",X"4E",X"0A",X"D9",X"3E",X"02",
		X"6F",X"DD",X"4E",X"08",X"06",X"08",X"FD",X"7E",X"00",X"E6",X"41",X"EE",X"41",X"20",X"6D",X"FD",
		X"56",X"06",X"FD",X"5E",X"05",X"1A",X"67",X"13",X"1A",X"D9",X"85",X"1F",X"67",X"FD",X"7E",X"0A",
		X"91",X"30",X"02",X"ED",X"44",X"BC",X"D9",X"30",X"53",X"7C",X"85",X"1F",X"67",X"FD",X"7E",X"08",
		X"91",X"30",X"02",X"ED",X"44",X"BC",X"30",X"44",X"DD",X"7E",X"0D",X"FD",X"B6",X"0C",X"DD",X"77",
		X"0D",X"FD",X"7E",X"0D",X"DD",X"B6",X"0C",X"FD",X"77",X"0D",X"DD",X"E5",X"FD",X"E5",X"DD",X"56",
		X"02",X"DD",X"5E",X"01",X"D5",X"DD",X"E1",X"FD",X"56",X"02",X"FD",X"5E",X"01",X"D5",X"FD",X"E1",
		X"DD",X"7E",X"03",X"FD",X"77",X"03",X"DD",X"7E",X"04",X"FD",X"77",X"04",X"DD",X"7E",X"09",X"FD",
		X"77",X"09",X"DD",X"7E",X"0A",X"FD",X"77",X"0A",X"FD",X"E1",X"DD",X"E1",X"11",X"2E",X"00",X"FD",
		X"19",X"10",X"83",X"D9",X"C9",X"21",X"E4",X"80",X"7E",X"23",X"46",X"A8",X"4F",X"3A",X"00",X"98",
		X"2F",X"77",X"2B",X"70",X"A1",X"E6",X"C0",X"23",X"23",X"CB",X"7F",X"28",X"01",X"34",X"23",X"CB",
		X"77",X"28",X"01",X"34",X"CD",X"42",X"11",X"CD",X"A9",X"11",X"C9",X"3A",X"EE",X"80",X"C6",X"99",
		X"27",X"32",X"EE",X"80",X"C9",X"47",X"B7",X"C8",X"3E",X"FF",X"32",X"54",X"85",X"3A",X"EE",X"80",
		X"FE",X"99",X"C8",X"80",X"27",X"30",X"02",X"3E",X"99",X"32",X"EE",X"80",X"3E",X"05",X"CD",X"1F",
		X"08",X"C9",X"D9",X"11",X"E6",X"80",X"3A",X"E8",X"80",X"4F",X"21",X"EE",X"11",X"CD",X"67",X"11",
		X"79",X"32",X"E8",X"80",X"11",X"E7",X"80",X"3A",X"E9",X"80",X"4F",X"21",X"1E",X"12",X"CD",X"67",
		X"11",X"79",X"32",X"E9",X"80",X"D9",X"C9",X"3A",X"02",X"98",X"2F",X"E6",X"06",X"CB",X"3F",X"47",
		X"28",X"08",X"D5",X"11",X"0C",X"00",X"19",X"10",X"FD",X"D1",X"1A",X"B7",X"C8",X"09",X"AF",X"86",
		X"08",X"79",X"FE",X"0B",X"20",X"0A",X"D5",X"11",X"0C",X"00",X"AF",X"ED",X"52",X"0E",X"FF",X"D1",
		X"0C",X"23",X"08",X"EB",X"35",X"CD",X"9F",X"11",X"EB",X"20",X"E4",X"CD",X"25",X"11",X"C9",X"F5",
		X"3A",X"EA",X"80",X"3C",X"32",X"EA",X"80",X"F1",X"C9",X"3A",X"ED",X"80",X"B7",X"28",X"25",X"3A",
		X"EC",X"80",X"B7",X"28",X"05",X"3D",X"32",X"EC",X"80",X"C9",X"3A",X"EB",X"80",X"B7",X"28",X"0E",
		X"3E",X"00",X"32",X"02",X"A8",X"32",X"EB",X"80",X"3E",X"0C",X"32",X"EC",X"80",X"C9",X"3E",X"00",
		X"32",X"ED",X"80",X"C9",X"3A",X"EA",X"80",X"B7",X"C8",X"3D",X"32",X"EA",X"80",X"3E",X"FF",X"32",
		X"ED",X"80",X"32",X"EB",X"80",X"32",X"02",X"A8",X"3E",X"04",X"32",X"EC",X"80",X"C9",X"04",X"04",
		X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"03",X"03",X"03",X"03",X"03",X"03",
		X"03",X"03",X"03",X"03",X"03",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"01",X"00",X"00",X"01",
		X"00",X"00",X"01",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"DD",X"21",
		X"20",X"85",X"21",X"00",X"98",X"CD",X"9B",X"12",X"DD",X"23",X"23",X"CD",X"9B",X"12",X"DD",X"23",
		X"23",X"CD",X"9B",X"12",X"3A",X"59",X"85",X"FE",X"02",X"C0",X"3A",X"02",X"98",X"E6",X"08",X"C0",
		X"3A",X"23",X"85",X"E6",X"C0",X"6F",X"3A",X"24",X"85",X"E6",X"3C",X"B5",X"32",X"23",X"85",X"3A",
		X"24",X"85",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"E6",X"03",
		X"6F",X"3A",X"23",X"85",X"E6",X"FC",X"B5",X"32",X"23",X"85",X"C9",X"DD",X"7E",X"00",X"DD",X"46",
		X"03",X"A8",X"57",X"7E",X"2F",X"4F",X"7A",X"A1",X"DD",X"77",X"06",X"DD",X"70",X"00",X"DD",X"71",
		X"03",X"C9",X"CD",X"26",X"09",X"D2",X"E0",X"09",X"CD",X"CE",X"08",X"D2",X"F9",X"14",X"FD",X"2A",
		X"DA",X"80",X"FD",X"66",X"02",X"FD",X"6E",X"01",X"E5",X"DD",X"E1",X"CD",X"07",X"17",X"CD",X"5F",
		X"15",X"FD",X"CB",X"00",X"F6",X"FD",X"CB",X"0C",X"D6",X"DD",X"CB",X"00",X"EE",X"FD",X"CB",X"00",
		X"D6",X"FD",X"36",X"0D",X"00",X"3E",X"0A",X"CD",X"1F",X"08",X"DD",X"E5",X"CD",X"BC",X"09",X"FD",
		X"E1",X"DD",X"CB",X"0D",X"4E",X"C2",X"E8",X"14",X"DD",X"7E",X"0D",X"B7",X"CA",X"0B",X"13",X"FD",
		X"36",X"01",X"04",X"FD",X"CB",X"00",X"CE",X"DD",X"36",X"0D",X"00",X"FD",X"7E",X"07",X"FE",X"35",
		X"20",X"06",X"DD",X"CB",X"00",X"96",X"18",X"04",X"DD",X"CB",X"00",X"D6",X"FD",X"CB",X"00",X"4E",
		X"20",X"0B",X"FD",X"36",X"01",X"14",X"FD",X"CB",X"00",X"CE",X"CD",X"37",X"13",X"CD",X"3D",X"14",
		X"FD",X"E5",X"CD",X"BC",X"09",X"18",X"B8",X"CD",X"06",X"19",X"CD",X"DC",X"14",X"DD",X"CB",X"00",
		X"A6",X"FE",X"01",X"20",X"17",X"21",X"40",X"02",X"FD",X"75",X"03",X"FD",X"74",X"04",X"FD",X"36",
		X"09",X"00",X"FD",X"36",X"0A",X"00",X"21",X"71",X"15",X"C3",X"2A",X"14",X"FE",X"03",X"20",X"18",
		X"21",X"40",X"02",X"FD",X"75",X"03",X"FD",X"74",X"04",X"21",X"C0",X"FD",X"FD",X"75",X"09",X"FD",
		X"74",X"0A",X"21",X"71",X"15",X"C3",X"2A",X"14",X"FE",X"02",X"20",X"17",X"FD",X"36",X"03",X"00",
		X"FD",X"36",X"04",X"00",X"21",X"C0",X"FD",X"FD",X"75",X"09",X"FD",X"74",X"0A",X"21",X"AB",X"15",
		X"C3",X"2A",X"14",X"FE",X"06",X"20",X"15",X"21",X"C0",X"FD",X"FD",X"75",X"03",X"FD",X"74",X"04",
		X"FD",X"75",X"09",X"FD",X"74",X"0A",X"21",X"AB",X"15",X"C3",X"2A",X"14",X"FE",X"04",X"20",X"17",
		X"21",X"C0",X"FD",X"FD",X"75",X"03",X"FD",X"74",X"04",X"FD",X"36",X"09",X"00",X"FD",X"36",X"0A",
		X"00",X"21",X"8E",X"15",X"C3",X"2A",X"14",X"FE",X"0C",X"20",X"18",X"21",X"C0",X"FD",X"FD",X"75",
		X"03",X"FD",X"74",X"04",X"21",X"40",X"02",X"FD",X"75",X"09",X"FD",X"74",X"0A",X"21",X"8E",X"15",
		X"C3",X"2A",X"14",X"FE",X"08",X"20",X"17",X"FD",X"36",X"03",X"00",X"FD",X"36",X"04",X"00",X"21",
		X"40",X"02",X"FD",X"75",X"09",X"FD",X"74",X"0A",X"21",X"C8",X"15",X"C3",X"2A",X"14",X"FE",X"09",
		X"20",X"15",X"21",X"40",X"02",X"FD",X"75",X"03",X"FD",X"74",X"04",X"FD",X"75",X"09",X"FD",X"74",
		X"0A",X"21",X"C8",X"15",X"C3",X"2A",X"14",X"FD",X"36",X"03",X"00",X"FD",X"36",X"04",X"00",X"FD",
		X"36",X"09",X"00",X"FD",X"36",X"0A",X"00",X"21",X"C8",X"15",X"DD",X"75",X"05",X"DD",X"74",X"06",
		X"DD",X"36",X"04",X"01",X"FD",X"CB",X"00",X"96",X"DD",X"CB",X"00",X"E6",X"C9",X"DD",X"7E",X"0A",
		X"FE",X"17",X"30",X"18",X"CD",X"BE",X"14",X"FD",X"56",X"0A",X"FD",X"5E",X"09",X"CD",X"BE",X"0F",
		X"FD",X"72",X"0A",X"FD",X"73",X"09",X"3E",X"18",X"DD",X"77",X"0A",X"C9",X"DD",X"7E",X"0A",X"FE",
		X"D8",X"38",X"18",X"CD",X"BE",X"14",X"FD",X"56",X"0A",X"FD",X"5E",X"09",X"CD",X"BE",X"0F",X"FD",
		X"72",X"0A",X"FD",X"73",X"09",X"3E",X"D6",X"DD",X"77",X"0A",X"C9",X"21",X"34",X"86",X"DD",X"7E",
		X"08",X"BE",X"38",X"19",X"CD",X"BE",X"14",X"FD",X"56",X"04",X"FD",X"5E",X"03",X"CD",X"BE",X"0F",
		X"FD",X"72",X"04",X"FD",X"73",X"03",X"7E",X"3D",X"3D",X"DD",X"77",X"08",X"C9",X"21",X"33",X"86",
		X"DD",X"7E",X"08",X"BE",X"D0",X"CD",X"BE",X"14",X"FD",X"56",X"04",X"FD",X"5E",X"03",X"CD",X"BE",
		X"0F",X"FD",X"72",X"04",X"FD",X"73",X"03",X"7E",X"3C",X"3C",X"DD",X"77",X"08",X"C9",X"FD",X"7E",
		X"04",X"B7",X"F2",X"C7",X"14",X"2F",X"3C",X"FE",X"04",X"30",X"0C",X"FD",X"7E",X"0A",X"B7",X"F2",
		X"D4",X"14",X"2F",X"3C",X"FE",X"04",X"D8",X"E1",X"E1",X"C3",X"E8",X"14",X"CD",X"42",X"08",X"FE",
		X"32",X"38",X"02",X"78",X"C9",X"E6",X"0F",X"C9",X"3E",X"05",X"CD",X"1F",X"08",X"01",X"02",X"02",
		X"CD",X"57",X"1F",X"CD",X"01",X"15",X"C3",X"BE",X"12",X"CD",X"36",X"0A",X"CD",X"BC",X"09",X"18",
		X"FB",X"AF",X"DD",X"77",X"0D",X"FD",X"77",X"04",X"FD",X"77",X"03",X"FD",X"77",X"0A",X"FD",X"77",
		X"09",X"DD",X"CB",X"0C",X"96",X"DD",X"CB",X"00",X"A6",X"DD",X"CB",X"00",X"B6",X"21",X"E5",X"15",
		X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",X"36",X"04",X"01",X"DD",X"CB",X"00",X"E6",X"CD",X"BC",
		X"09",X"DD",X"CB",X"00",X"66",X"20",X"F7",X"DD",X"36",X"0A",X"00",X"DD",X"36",X"08",X"00",X"DD",
		X"66",X"02",X"DD",X"6E",X"01",X"E5",X"FD",X"E1",X"FD",X"36",X"06",X"00",X"FD",X"36",X"0C",X"00",
		X"DD",X"CB",X"00",X"96",X"CD",X"42",X"08",X"F6",X"20",X"E6",X"7F",X"CD",X"10",X"0A",X"C9",X"21",
		X"71",X"15",X"FD",X"75",X"05",X"FD",X"74",X"06",X"FD",X"36",X"04",X"01",X"FD",X"CB",X"00",X"E6",
		X"C9",X"00",X"00",X"01",X"00",X"00",X"0C",X"0C",X"05",X"35",X"07",X"0C",X"0C",X"04",X"33",X"07",
		X"0C",X"0C",X"05",X"34",X"07",X"0C",X"0C",X"04",X"33",X"07",X"00",X"01",X"76",X"15",X"00",X"00",
		X"01",X"00",X"00",X"0C",X"0C",X"04",X"35",X"07",X"0C",X"0C",X"03",X"33",X"07",X"0C",X"0C",X"05",
		X"34",X"07",X"0C",X"0C",X"03",X"33",X"07",X"00",X"01",X"93",X"15",X"00",X"00",X"01",X"00",X"00",
		X"0C",X"0C",X"04",X"35",X"07",X"0C",X"0C",X"03",X"33",X"07",X"0C",X"0C",X"05",X"34",X"07",X"0C",
		X"0C",X"03",X"33",X"07",X"00",X"01",X"B0",X"15",X"00",X"00",X"01",X"00",X"00",X"0C",X"0C",X"04",
		X"35",X"07",X"0C",X"0C",X"03",X"33",X"07",X"0C",X"0C",X"05",X"34",X"07",X"0C",X"0C",X"03",X"33",
		X"07",X"00",X"01",X"CD",X"15",X"00",X"00",X"01",X"00",X"00",X"01",X"00",X"03",X"1B",X"02",X"01",
		X"00",X"03",X"9B",X"03",X"01",X"00",X"03",X"1A",X"04",X"01",X"00",X"03",X"9A",X"05",X"01",X"00",
		X"03",X"19",X"06",X"01",X"00",X"03",X"99",X"07",X"01",X"00",X"03",X"17",X"02",X"01",X"00",X"03",
		X"97",X"03",X"01",X"00",X"03",X"16",X"04",X"01",X"00",X"03",X"96",X"05",X"01",X"00",X"03",X"12",
		X"06",X"01",X"00",X"03",X"92",X"07",X"00",X"00",X"00",X"00",X"9D",X"CD",X"26",X"09",X"D2",X"E0",
		X"09",X"CD",X"CE",X"08",X"D2",X"FF",X"16",X"FD",X"2A",X"DA",X"80",X"FD",X"66",X"02",X"FD",X"6E",
		X"01",X"E5",X"DD",X"E1",X"CD",X"07",X"17",X"CD",X"F7",X"17",X"FD",X"CB",X"00",X"F6",X"FD",X"CB",
		X"0C",X"D6",X"DD",X"CB",X"00",X"EE",X"FD",X"CB",X"00",X"D6",X"FD",X"36",X"0D",X"00",X"3E",X"0A",
		X"CD",X"1F",X"08",X"DD",X"E5",X"CD",X"BC",X"09",X"FD",X"E1",X"DD",X"7E",X"0D",X"B7",X"C2",X"EE",
		X"16",X"CD",X"7B",X"16",X"FD",X"E5",X"CD",X"BC",X"09",X"18",X"ED",X"DD",X"7E",X"0A",X"FE",X"17",
		X"30",X"15",X"FD",X"56",X"0A",X"FD",X"5E",X"09",X"CD",X"BE",X"0F",X"FD",X"72",X"0A",X"FD",X"73",
		X"09",X"3E",X"17",X"DD",X"77",X"0A",X"C9",X"DD",X"7E",X"0A",X"FE",X"D8",X"38",X"15",X"FD",X"56",
		X"0A",X"FD",X"5E",X"09",X"CD",X"BE",X"0F",X"FD",X"72",X"0A",X"FD",X"73",X"09",X"3E",X"D7",X"DD",
		X"77",X"0A",X"C9",X"21",X"34",X"86",X"DD",X"7E",X"08",X"BE",X"38",X"15",X"FD",X"56",X"04",X"FD",
		X"5E",X"03",X"CD",X"BE",X"0F",X"FD",X"72",X"04",X"FD",X"73",X"03",X"7E",X"3D",X"DD",X"77",X"08",
		X"C9",X"21",X"33",X"86",X"DD",X"7E",X"08",X"BE",X"D0",X"FD",X"56",X"04",X"FD",X"5E",X"03",X"CD",
		X"BE",X"0F",X"FD",X"72",X"04",X"FD",X"73",X"03",X"7E",X"3C",X"DD",X"77",X"08",X"C9",X"3E",X"05",
		X"CD",X"1F",X"08",X"01",X"05",X"01",X"CD",X"57",X"1F",X"CD",X"01",X"15",X"C3",X"37",X"16",X"CD",
		X"36",X"0A",X"CD",X"BC",X"09",X"18",X"FB",X"CD",X"42",X"08",X"E6",X"03",X"28",X"0C",X"FE",X"01",
		X"28",X"3C",X"FE",X"02",X"CA",X"85",X"17",X"C3",X"BE",X"17",X"3A",X"1A",X"82",X"FE",X"AA",X"30",
		X"07",X"3A",X"1C",X"82",X"FE",X"78",X"38",X"DF",X"21",X"33",X"86",X"7E",X"3C",X"3C",X"FD",X"77",
		X"08",X"FD",X"36",X"0A",X"18",X"11",X"60",X"03",X"DD",X"72",X"04",X"DD",X"73",X"03",X"DD",X"72",
		X"0A",X"DD",X"73",X"09",X"3E",X"0A",X"DD",X"77",X"01",X"DD",X"CB",X"00",X"CE",X"C9",X"3A",X"1A",
		X"82",X"FE",X"AA",X"30",X"07",X"3A",X"1C",X"82",X"FE",X"78",X"30",X"AB",X"21",X"33",X"86",X"7E",
		X"3C",X"3C",X"FD",X"77",X"08",X"FD",X"36",X"0A",X"D6",X"11",X"60",X"03",X"DD",X"72",X"04",X"DD",
		X"73",X"03",X"CD",X"BE",X"0F",X"DD",X"72",X"0A",X"DD",X"73",X"09",X"3E",X"0A",X"DD",X"77",X"01",
		X"DD",X"CB",X"00",X"CE",X"C9",X"3A",X"1A",X"82",X"FE",X"46",X"DA",X"95",X"17",X"3A",X"1C",X"82",
		X"FE",X"78",X"D2",X"07",X"17",X"21",X"34",X"86",X"7E",X"3D",X"3D",X"FD",X"77",X"08",X"FD",X"36",
		X"0A",X"D6",X"11",X"60",X"03",X"CD",X"BE",X"0F",X"DD",X"72",X"04",X"DD",X"73",X"03",X"DD",X"72",
		X"0A",X"DD",X"73",X"09",X"3E",X"0A",X"DD",X"77",X"01",X"DD",X"CB",X"00",X"CE",X"C9",X"3A",X"1A",
		X"82",X"FE",X"46",X"DA",X"CE",X"17",X"3A",X"1C",X"82",X"FE",X"78",X"DA",X"07",X"17",X"21",X"34",
		X"86",X"7E",X"3D",X"3D",X"FD",X"77",X"08",X"FD",X"36",X"0A",X"18",X"11",X"60",X"03",X"DD",X"72",
		X"0A",X"DD",X"73",X"09",X"CD",X"BE",X"0F",X"DD",X"72",X"04",X"DD",X"73",X"03",X"3E",X"0A",X"DD",
		X"77",X"01",X"DD",X"CB",X"00",X"CE",X"C9",X"21",X"09",X"18",X"FD",X"75",X"05",X"FD",X"74",X"06",
		X"FD",X"36",X"04",X"01",X"FD",X"CB",X"00",X"E6",X"C9",X"00",X"00",X"01",X"00",X"00",X"0C",X"0C",
		X"04",X"2E",X"01",X"0C",X"0C",X"04",X"2D",X"01",X"0C",X"0C",X"04",X"2C",X"01",X"0C",X"0C",X"04",
		X"2B",X"01",X"0C",X"0C",X"04",X"2C",X"01",X"0C",X"0C",X"04",X"2D",X"01",X"00",X"01",X"0E",X"18",
		X"CD",X"26",X"09",X"D2",X"E0",X"09",X"CD",X"CE",X"08",X"D2",X"47",X"19",X"FD",X"2A",X"DA",X"80",
		X"FD",X"66",X"02",X"FD",X"6E",X"01",X"E5",X"DD",X"E1",X"CD",X"07",X"17",X"CD",X"4F",X"19",X"FD",
		X"36",X"0D",X"00",X"FD",X"CB",X"00",X"F6",X"FD",X"CB",X"0C",X"D6",X"DD",X"CB",X"00",X"EE",X"FD",
		X"CB",X"00",X"D6",X"3E",X"0A",X"CD",X"1F",X"08",X"DD",X"E5",X"CD",X"BC",X"09",X"FD",X"E1",X"DD",
		X"7E",X"0D",X"B7",X"C2",X"36",X"19",X"FD",X"CB",X"00",X"4E",X"20",X"11",X"CD",X"42",X"08",X"E6",
		X"1F",X"F6",X"08",X"FD",X"77",X"01",X"FD",X"CB",X"00",X"CE",X"CD",X"97",X"18",X"CD",X"7B",X"16",
		X"FD",X"E5",X"CD",X"BC",X"09",X"18",X"D6",X"CD",X"06",X"19",X"CD",X"27",X"19",X"CB",X"57",X"28",
		X"12",X"21",X"20",X"FE",X"FD",X"75",X"03",X"FD",X"74",X"04",X"FD",X"36",X"09",X"00",X"FD",X"36",
		X"0A",X"00",X"C9",X"CB",X"4F",X"28",X"12",X"FD",X"36",X"03",X"00",X"FD",X"36",X"04",X"00",X"21",
		X"20",X"FE",X"FD",X"75",X"09",X"FD",X"74",X"0A",X"C9",X"CB",X"47",X"28",X"12",X"21",X"E0",X"01",
		X"FD",X"75",X"03",X"FD",X"74",X"04",X"FD",X"36",X"09",X"00",X"FD",X"36",X"0A",X"00",X"C9",X"CB",
		X"5F",X"28",X"12",X"FD",X"36",X"03",X"00",X"FD",X"36",X"04",X"00",X"21",X"E0",X"01",X"FD",X"75",
		X"09",X"FD",X"74",X"0A",X"C9",X"FD",X"36",X"03",X"00",X"FD",X"36",X"04",X"00",X"FD",X"36",X"09",
		X"00",X"FD",X"36",X"0A",X"00",X"C9",X"06",X"00",X"3A",X"A6",X"81",X"FD",X"BE",X"0C",X"38",X"04",
		X"CB",X"D8",X"18",X"04",X"28",X"02",X"CB",X"C8",X"3A",X"A0",X"81",X"FD",X"BE",X"06",X"38",X"03",
		X"CB",X"C0",X"C9",X"C8",X"CB",X"D0",X"C9",X"CD",X"42",X"08",X"CB",X"77",X"28",X"04",X"78",X"E6",
		X"0A",X"C9",X"78",X"E6",X"05",X"C9",X"3E",X"05",X"CD",X"1F",X"08",X"01",X"05",X"01",X"CD",X"57",
		X"1F",X"CD",X"01",X"15",X"C3",X"3C",X"18",X"CD",X"36",X"0A",X"CD",X"BC",X"09",X"18",X"FB",X"21",
		X"61",X"19",X"FD",X"75",X"05",X"FD",X"74",X"06",X"FD",X"36",X"04",X"01",X"FD",X"CB",X"00",X"E6",
		X"C9",X"00",X"00",X"01",X"00",X"00",X"0E",X"0E",X"04",X"2A",X"03",X"0E",X"0E",X"04",X"29",X"03",
		X"0E",X"0E",X"04",X"28",X"03",X"0E",X"0E",X"04",X"27",X"03",X"0E",X"0E",X"04",X"28",X"03",X"0E",
		X"0E",X"04",X"29",X"03",X"00",X"01",X"66",X"19",X"21",X"44",X"86",X"35",X"C0",X"3E",X"04",X"77",
		X"21",X"45",X"86",X"34",X"3E",X"10",X"21",X"42",X"88",X"11",X"20",X"00",X"06",X"1C",X"77",X"19",
		X"10",X"FC",X"21",X"42",X"88",X"11",X"1B",X"00",X"19",X"11",X"20",X"00",X"06",X"1C",X"77",X"19",
		X"10",X"FC",X"CF",X"48",X"10",X"5B",X"5B",X"5B",X"5B",X"20",X"45",X"58",X"49",X"54",X"20",X"5B",
		X"5B",X"5B",X"5B",X"00",X"CF",X"48",X"E8",X"5B",X"5B",X"5B",X"5B",X"20",X"45",X"58",X"49",X"54",
		X"20",X"5B",X"5B",X"5B",X"5B",X"00",X"21",X"05",X"90",X"34",X"21",X"3B",X"90",X"34",X"DD",X"36",
		X"0B",X"00",X"FD",X"CB",X"00",X"FE",X"C9",X"3E",X"00",X"32",X"01",X"A8",X"32",X"02",X"A8",X"32",
		X"03",X"A8",X"32",X"04",X"A8",X"32",X"07",X"A8",X"32",X"06",X"A8",X"3E",X"9B",X"32",X"03",X"98",
		X"3E",X"88",X"32",X"03",X"A0",X"31",X"68",X"80",X"21",X"68",X"80",X"0E",X"08",X"CD",X"B7",X"05",
		X"3E",X"FF",X"32",X"E4",X"80",X"32",X"E5",X"80",X"21",X"B0",X"1A",X"11",X"EF",X"80",X"01",X"3C",
		X"00",X"ED",X"B0",X"31",X"68",X"80",X"21",X"00",X"90",X"0E",X"01",X"CD",X"B7",X"05",X"3E",X"01",
		X"32",X"59",X"85",X"CD",X"60",X"1A",X"CD",X"C2",X"1C",X"FD",X"21",X"EC",X"1A",X"CD",X"A4",X"09",
		X"CD",X"BC",X"09",X"DD",X"21",X"12",X"82",X"DD",X"CB",X"0B",X"46",X"28",X"F3",X"CD",X"69",X"0A",
		X"21",X"12",X"82",X"CB",X"F6",X"CD",X"DB",X"1F",X"3E",X"02",X"CD",X"7D",X"1A",X"C3",X"2E",X"1A",
		X"E1",X"22",X"50",X"85",X"32",X"52",X"85",X"CD",X"69",X"0A",X"CD",X"6F",X"08",X"AF",X"32",X"E3",
		X"80",X"3E",X"FF",X"32",X"01",X"A8",X"2A",X"50",X"85",X"3A",X"52",X"85",X"E9",X"F5",X"3E",X"1E",
		X"CD",X"88",X"1A",X"F1",X"3D",X"20",X"F6",X"C9",X"F5",X"D5",X"E5",X"C5",X"DD",X"2A",X"DA",X"80",
		X"DD",X"CB",X"00",X"EE",X"DD",X"36",X"03",X"01",X"CD",X"89",X"2D",X"3A",X"54",X"85",X"B7",X"C4",
		X"4F",X"06",X"DD",X"CB",X"00",X"6E",X"20",X"F0",X"C1",X"E1",X"D1",X"F1",X"3D",X"20",X"D9",X"C9",
		X"01",X"04",X"80",X"4F",X"42",X"45",X"01",X"01",X"00",X"47",X"4A",X"4C",X"00",X"39",X"10",X"52",
		X"41",X"51",X"00",X"28",X"70",X"4A",X"56",X"43",X"00",X"18",X"30",X"45",X"4C",X"50",X"00",X"17",
		X"70",X"4A",X"49",X"4D",X"00",X"16",X"40",X"4A",X"4D",X"48",X"00",X"15",X"90",X"44",X"41",X"4E",
		X"00",X"14",X"10",X"41",X"50",X"48",X"00",X"12",X"00",X"42",X"49",X"4C",X"3E",X"FF",X"32",X"55",
		X"85",X"CD",X"85",X"08",X"3E",X"14",X"32",X"33",X"86",X"3E",X"E6",X"32",X"34",X"86",X"3E",X"00",
		X"32",X"36",X"86",X"32",X"37",X"86",X"DD",X"21",X"12",X"82",X"DD",X"CB",X"00",X"F6",X"DD",X"21",
		X"12",X"82",X"FD",X"21",X"9A",X"81",X"21",X"2A",X"85",X"36",X"00",X"21",X"2B",X"85",X"36",X"00",
		X"CD",X"63",X"1C",X"DD",X"CB",X"00",X"D6",X"AF",X"DD",X"77",X"0D",X"DD",X"CB",X"0C",X"C6",X"DD",
		X"36",X"08",X"0A",X"DD",X"36",X"0A",X"CF",X"DD",X"CB",X"00",X"F6",X"3E",X"05",X"32",X"78",X"85",
		X"21",X"E7",X"1B",X"E5",X"FD",X"21",X"9A",X"81",X"FD",X"CB",X"00",X"56",X"20",X"0F",X"3E",X"03",
		X"FD",X"77",X"02",X"FD",X"CB",X"00",X"D6",X"3E",X"FE",X"21",X"40",X"86",X"77",X"3A",X"36",X"86",
		X"CB",X"4F",X"C2",X"77",X"1B",X"3A",X"36",X"86",X"E6",X"3C",X"21",X"2B",X"85",X"46",X"77",X"A8",
		X"C4",X"80",X"1C",X"DD",X"CB",X"00",X"E6",X"01",X"00",X"00",X"11",X"00",X"00",X"3A",X"36",X"86",
		X"CB",X"4F",X"C2",X"95",X"1B",X"3A",X"36",X"86",X"67",X"CD",X"41",X"1C",X"CD",X"4B",X"1C",X"CD",
		X"52",X"1C",X"CD",X"59",X"1C",X"FD",X"70",X"04",X"FD",X"71",X"03",X"FD",X"72",X"0A",X"FD",X"73",
		X"09",X"3A",X"36",X"86",X"CB",X"4F",X"C4",X"F3",X"1B",X"FD",X"CB",X"00",X"4E",X"C2",X"C9",X"1B",
		X"E1",X"7E",X"B7",X"CA",X"D9",X"1B",X"FD",X"77",X"01",X"FD",X"CB",X"00",X"CE",X"23",X"7E",X"32",
		X"36",X"86",X"23",X"7E",X"32",X"37",X"86",X"23",X"E5",X"CD",X"89",X"2D",X"CD",X"BC",X"09",X"3A",
		X"54",X"85",X"B7",X"C4",X"4F",X"06",X"C3",X"44",X"1B",X"DD",X"CB",X"0B",X"C6",X"3E",X"00",X"32",
		X"55",X"85",X"CD",X"BC",X"09",X"18",X"FB",X"21",X"10",X"00",X"30",X"06",X"00",X"50",X"10",X"00",
		X"00",X"00",X"00",X"3A",X"36",X"86",X"E6",X"3C",X"C8",X"DD",X"CB",X"00",X"A6",X"06",X"00",X"CB",
		X"3F",X"CB",X"3F",X"4F",X"21",X"31",X"1C",X"09",X"7E",X"FD",X"77",X"07",X"3A",X"2A",X"85",X"FE",
		X"07",X"C8",X"D0",X"DD",X"CB",X"00",X"6E",X"C0",X"DD",X"36",X"03",X"02",X"DD",X"CB",X"00",X"EE",
		X"FD",X"21",X"DD",X"3D",X"CD",X"A4",X"09",X"FD",X"21",X"9A",X"81",X"3E",X"04",X"CD",X"1F",X"08",
		X"C9",X"00",X"3E",X"3F",X"00",X"95",X"94",X"93",X"00",X"15",X"14",X"13",X"00",X"00",X"00",X"00",
		X"00",X"CB",X"54",X"C8",X"11",X"00",X"02",X"CD",X"BE",X"0F",X"C9",X"CB",X"5C",X"C8",X"11",X"00",
		X"02",X"C9",X"CB",X"64",X"C8",X"01",X"00",X"02",X"C9",X"CB",X"6C",X"C8",X"01",X"00",X"02",X"CD",
		X"C6",X"0F",X"C9",X"21",X"42",X"38",X"11",X"5A",X"85",X"01",X"1E",X"00",X"ED",X"B0",X"21",X"5A",
		X"85",X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",X"36",X"04",X"01",X"DD",X"CB",X"00",X"E6",X"C9",
		X"21",X"2F",X"3D",X"06",X"00",X"3A",X"2B",X"85",X"CB",X"3F",X"CB",X"3F",X"4F",X"09",X"09",X"09",
		X"09",X"7E",X"B7",X"C8",X"DD",X"CB",X"00",X"A6",X"DD",X"E5",X"DD",X"21",X"5A",X"85",X"11",X"05",
		X"00",X"DD",X"19",X"DD",X"77",X"03",X"DD",X"19",X"23",X"7E",X"DD",X"77",X"03",X"DD",X"19",X"23",
		X"7E",X"DD",X"77",X"03",X"DD",X"19",X"23",X"7E",X"DD",X"77",X"03",X"DD",X"E1",X"DD",X"36",X"04",
		X"01",X"C9",X"CD",X"82",X"05",X"CD",X"5F",X"22",X"CD",X"2D",X"06",X"CD",X"4F",X"06",X"CF",X"28",
		X"00",X"53",X"54",X"45",X"52",X"4E",X"20",X"50",X"52",X"4F",X"55",X"44",X"4C",X"59",X"20",X"50",
		X"52",X"45",X"53",X"45",X"4E",X"54",X"53",X"00",X"CF",X"50",X"18",X"54",X"41",X"5A",X"5A",X"20",
		X"5B",X"20",X"4D",X"41",X"4E",X"49",X"41",X"00",X"CF",X"10",X"E0",X"50",X"55",X"4C",X"4C",X"20",
		X"53",X"54",X"49",X"43",X"4B",X"20",X"46",X"4F",X"52",X"20",X"49",X"4E",X"53",X"54",X"52",X"55",
		X"43",X"54",X"49",X"4F",X"4E",X"53",X"00",X"E7",X"06",X"07",X"05",X"E7",X"06",X"0D",X"02",X"E7",
		X"07",X"13",X"07",X"DF",X"28",X"CF",X"40",X"28",X"20",X"54",X"4F",X"50",X"20",X"31",X"30",X"20",
		X"53",X"43",X"4F",X"52",X"45",X"53",X"20",X"00",X"3E",X"38",X"32",X"05",X"89",X"32",X"05",X"8B",
		X"06",X"0A",X"21",X"A7",X"8A",X"36",X"38",X"23",X"23",X"10",X"FA",X"21",X"12",X"82",X"CB",X"F6",
		X"11",X"EF",X"80",X"21",X"38",X"38",X"3E",X"01",X"08",X"D5",X"EB",X"7E",X"23",X"B6",X"23",X"B6",
		X"EB",X"D1",X"C8",X"E5",X"D5",X"08",X"32",X"00",X"80",X"08",X"06",X"02",X"11",X"00",X"80",X"CD",
		X"27",X"05",X"01",X"00",X"20",X"09",X"D1",X"06",X"06",X"CD",X"27",X"05",X"13",X"13",X"13",X"01",
		X"00",X"30",X"09",X"CD",X"BF",X"04",X"06",X"03",X"3E",X"20",X"CD",X"6A",X"05",X"10",X"F9",X"06",
		X"03",X"1A",X"13",X"CD",X"6A",X"05",X"10",X"F9",X"E1",X"01",X"10",X"00",X"09",X"08",X"C6",X"01",
		X"27",X"FE",X"11",X"DA",X"58",X"1D",X"3E",X"01",X"CD",X"7D",X"1A",X"C9",X"3A",X"59",X"85",X"B7",
		X"C8",X"CD",X"4A",X"1F",X"0E",X"0A",X"11",X"EF",X"80",X"E5",X"D5",X"06",X"03",X"1A",X"BE",X"38",
		X"11",X"20",X"04",X"13",X"23",X"10",X"F6",X"D1",X"21",X"06",X"00",X"19",X"EB",X"E1",X"0D",X"20",
		X"E8",X"C9",X"D1",X"D5",X"0D",X"28",X"16",X"06",X"00",X"21",X"00",X"00",X"09",X"29",X"09",X"29",
		X"E5",X"19",X"2B",X"54",X"5D",X"01",X"06",X"00",X"09",X"EB",X"C1",X"ED",X"B8",X"D1",X"E1",X"01",
		X"03",X"00",X"ED",X"B0",X"D5",X"CD",X"82",X"05",X"CD",X"07",X"2F",X"CD",X"89",X"06",X"DF",X"1A",
		X"CF",X"20",X"28",X"43",X"4F",X"4E",X"47",X"52",X"41",X"54",X"55",X"4C",X"41",X"54",X"49",X"4F",
		X"4E",X"53",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"00",X"21",X"28",X"D8",X"11",X"59",X"85",
		X"06",X"01",X"CD",X"27",X"05",X"E7",X"0A",X"07",X"06",X"DF",X"4C",X"CF",X"50",X"38",X"59",X"4F",
		X"55",X"20",X"4D",X"41",X"44",X"45",X"20",X"54",X"48",X"45",X"00",X"CF",X"48",X"48",X"54",X"41",
		X"5A",X"5A",X"20",X"5B",X"20",X"4D",X"41",X"4E",X"49",X"41",X"43",X"53",X"00",X"CF",X"50",X"58",
		X"48",X"41",X"4C",X"4C",X"20",X"4F",X"46",X"20",X"46",X"41",X"4D",X"45",X"00",X"E7",X"03",X"0F",
		X"05",X"CF",X"20",X"78",X"5B",X"20",X"45",X"4E",X"54",X"45",X"52",X"20",X"59",X"4F",X"55",X"52",
		X"20",X"49",X"4E",X"49",X"54",X"49",X"41",X"4C",X"53",X"20",X"5B",X"00",X"CF",X"70",X"88",X"5B",
		X"5B",X"5B",X"00",X"E7",X"03",X"16",X"07",X"CF",X"20",X"B0",X"4D",X"4F",X"56",X"45",X"20",X"53",
		X"54",X"49",X"43",X"4B",X"20",X"4C",X"45",X"46",X"54",X"20",X"4F",X"52",X"20",X"52",X"49",X"47",
		X"48",X"54",X"00",X"CF",X"30",X"C0",X"54",X"4F",X"20",X"43",X"48",X"41",X"4E",X"47",X"45",X"20",
		X"54",X"48",X"45",X"20",X"4C",X"45",X"54",X"54",X"45",X"52",X"00",X"CF",X"20",X"D0",X"50",X"55",
		X"4C",X"4C",X"20",X"53",X"54",X"49",X"43",X"4B",X"20",X"44",X"4F",X"57",X"4E",X"20",X"54",X"4F",
		X"20",X"45",X"4E",X"54",X"45",X"52",X"00",X"E1",X"E5",X"06",X"03",X"36",X"20",X"23",X"10",X"FB",
		X"21",X"88",X"70",X"CD",X"BF",X"04",X"D1",X"06",X"03",X"0E",X"41",X"3E",X"FA",X"32",X"50",X"85",
		X"CD",X"1F",X"1F",X"20",X"FB",X"79",X"E5",X"CD",X"6A",X"05",X"C5",X"D5",X"3E",X"05",X"CD",X"88",
		X"1A",X"D1",X"C1",X"E1",X"3A",X"50",X"85",X"3D",X"32",X"50",X"85",X"C8",X"CD",X"1F",X"1F",X"20",
		X"05",X"CD",X"25",X"1F",X"18",X"DA",X"79",X"12",X"13",X"CD",X"6A",X"05",X"10",X"CD",X"C9",X"3A",
		X"23",X"85",X"E6",X"08",X"C9",X"F5",X"D5",X"3A",X"23",X"85",X"57",X"79",X"CB",X"62",X"28",X"0A",
		X"C6",X"01",X"FE",X"5B",X"38",X"10",X"3E",X"40",X"18",X"0C",X"CB",X"6A",X"28",X"08",X"D6",X"01",
		X"FE",X"40",X"30",X"02",X"3E",X"5A",X"4F",X"D1",X"F1",X"C9",X"21",X"2B",X"81",X"3A",X"59",X"85",
		X"FE",X"01",X"C8",X"21",X"2E",X"81",X"C9",X"3A",X"55",X"85",X"B7",X"C0",X"3E",X"FF",X"32",X"53",
		X"85",X"3E",X"01",X"F5",X"CD",X"6F",X"1F",X"F1",X"3D",X"20",X"F8",X"CD",X"96",X"1F",X"C9",X"CD",
		X"4A",X"1F",X"1E",X"04",X"23",X"23",X"23",X"CB",X"38",X"08",X"04",X"2B",X"1D",X"10",X"FC",X"08",
		X"30",X"08",X"CB",X"21",X"CB",X"21",X"CB",X"21",X"CB",X"21",X"79",X"86",X"27",X"77",X"D0",X"2B",
		X"1D",X"C8",X"0E",X"01",X"18",X"F4",X"CD",X"D3",X"1F",X"EB",X"2A",X"30",X"85",X"7A",X"BC",X"D8",
		X"7B",X"BD",X"D8",X"3A",X"29",X"85",X"C6",X"01",X"27",X"32",X"29",X"85",X"3E",X"0F",X"CD",X"1F",
		X"08",X"CD",X"B8",X"1F",X"CD",X"D3",X"06",X"C9",X"2A",X"30",X"85",X"1E",X"10",X"16",X"00",X"06",
		X"04",X"CB",X"23",X"CB",X"12",X"10",X"FA",X"7D",X"83",X"27",X"6F",X"7C",X"8A",X"27",X"67",X"22",
		X"30",X"85",X"C9",X"CD",X"4A",X"1F",X"7E",X"23",X"6E",X"67",X"C9",X"CD",X"82",X"05",X"3E",X"00",
		X"32",X"07",X"A8",X"32",X"06",X"A8",X"3E",X"01",X"32",X"59",X"85",X"CD",X"5F",X"22",X"CD",X"2D",
		X"06",X"CD",X"4F",X"06",X"DF",X"02",X"CF",X"28",X"00",X"53",X"54",X"45",X"52",X"4E",X"20",X"50",
		X"52",X"4F",X"55",X"44",X"4C",X"59",X"20",X"50",X"52",X"45",X"53",X"45",X"4E",X"54",X"53",X"00",
		X"CF",X"10",X"E0",X"50",X"55",X"4C",X"4C",X"20",X"53",X"54",X"49",X"43",X"4B",X"20",X"46",X"4F",
		X"52",X"20",X"49",X"4E",X"53",X"54",X"52",X"55",X"43",X"54",X"49",X"4F",X"4E",X"53",X"00",X"CD",
		X"C3",X"20",X"DF",X"B7",X"DF",X"C3",X"CF",X"10",X"B0",X"5B",X"44",X"45",X"53",X"49",X"47",X"4E",
		X"45",X"44",X"20",X"41",X"4E",X"44",X"20",X"50",X"52",X"4F",X"47",X"52",X"41",X"4D",X"4D",X"45",
		X"44",X"20",X"42",X"59",X"5B",X"00",X"CF",X"10",X"C0",X"47",X"55",X"4E",X"41",X"52",X"53",X"20",
		X"4C",X"49",X"43",X"49",X"54",X"49",X"53",X"5B",X"5B",X"43",X"48",X"52",X"49",X"53",X"20",X"4F",
		X"42",X"45",X"52",X"54",X"48",X"00",X"CF",X"10",X"D0",X"45",X"58",X"54",X"52",X"41",X"20",X"4D",
		X"41",X"4E",X"20",X"45",X"56",X"45",X"52",X"59",X"20",X"31",X"30",X"30",X"30",X"30",X"20",X"50",
		X"4F",X"49",X"4E",X"54",X"53",X"00",X"3E",X"02",X"CD",X"7D",X"1A",X"FD",X"21",X"D6",X"43",X"CD",
		X"A4",X"09",X"CD",X"BC",X"09",X"DD",X"21",X"12",X"82",X"DD",X"CB",X"0B",X"46",X"28",X"F3",X"CD",
		X"69",X"0A",X"21",X"12",X"82",X"CB",X"F6",X"21",X"A8",X"10",X"01",X"08",X"1C",X"CD",X"C2",X"05",
		X"C3",X"10",X"07",X"11",X"63",X"8B",X"21",X"0F",X"21",X"06",X"17",X"C5",X"01",X"07",X"00",X"ED",
		X"B0",X"E5",X"EB",X"11",X"27",X"00",X"AF",X"ED",X"52",X"EB",X"E1",X"C1",X"10",X"ED",X"11",X"8D",
		X"8B",X"21",X"B0",X"21",X"06",X"19",X"C5",X"01",X"07",X"00",X"ED",X"B0",X"E5",X"EB",X"11",X"27",
		X"00",X"AF",X"ED",X"52",X"EB",X"E1",X"C1",X"10",X"ED",X"21",X"07",X"90",X"CD",X"06",X"21",X"21",
		X"1B",X"90",X"CD",X"06",X"21",X"C9",X"06",X"07",X"36",X"06",X"23",X"23",X"10",X"FA",X"C9",X"38",
		X"10",X"10",X"10",X"10",X"10",X"10",X"39",X"10",X"10",X"10",X"10",X"10",X"10",X"3A",X"3A",X"3A",
		X"3A",X"3A",X"3A",X"3A",X"3B",X"10",X"10",X"10",X"10",X"10",X"10",X"38",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"39",X"39",X"39",X"39",X"39",
		X"10",X"3A",X"10",X"10",X"3A",X"10",X"10",X"3B",X"10",X"10",X"10",X"3B",X"10",X"10",X"10",X"38",
		X"10",X"10",X"38",X"10",X"10",X"10",X"10",X"39",X"39",X"39",X"39",X"39",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"3A",X"10",X"10",X"10",X"10",X"3A",X"3A",X"3B",X"10",X"10",X"10",X"3B",X"10",
		X"3B",X"38",X"10",X"10",X"38",X"10",X"10",X"38",X"39",X"10",X"39",X"10",X"10",X"10",X"39",X"3A",
		X"3A",X"10",X"10",X"10",X"10",X"3A",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"3B",X"10",X"10",
		X"10",X"10",X"3B",X"3B",X"38",X"10",X"10",X"10",X"38",X"10",X"38",X"39",X"10",X"10",X"39",X"10",
		X"10",X"39",X"3A",X"10",X"3A",X"10",X"10",X"10",X"3A",X"3B",X"3B",X"10",X"10",X"10",X"10",X"3B",
		X"38",X"38",X"38",X"38",X"38",X"38",X"38",X"10",X"39",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"3A",X"10",X"10",X"10",X"10",X"10",X"3B",X"10",X"10",X"10",X"10",X"10",X"38",X"38",X"38",X"38",
		X"38",X"38",X"38",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"39",X"39",X"39",X"39",
		X"39",X"10",X"3A",X"10",X"10",X"3A",X"10",X"10",X"3B",X"10",X"10",X"10",X"3B",X"10",X"10",X"10",
		X"38",X"10",X"10",X"38",X"10",X"10",X"10",X"10",X"39",X"39",X"39",X"39",X"39",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"10",X"10",X"3B",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"38",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"39",X"10",X"10",
		X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"3B",X"3B",
		X"3B",X"3B",X"3B",X"3B",X"3B",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"38",X"38",
		X"38",X"38",X"38",X"10",X"39",X"10",X"10",X"39",X"10",X"10",X"3A",X"10",X"10",X"10",X"3A",X"10",
		X"10",X"10",X"3B",X"10",X"10",X"3B",X"10",X"10",X"10",X"10",X"38",X"38",X"38",X"38",X"38",X"3A",
		X"23",X"85",X"CB",X"57",X"C8",X"3A",X"23",X"85",X"CB",X"4F",X"C8",X"CB",X"47",X"C8",X"21",X"81",
		X"88",X"11",X"20",X"00",X"3A",X"3B",X"86",X"E6",X"0F",X"CD",X"D3",X"22",X"3A",X"3B",X"86",X"CB",
		X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CD",X"D3",X"22",X"3A",X"3C",X"86",X"E6",X"0F",X"CD",
		X"D3",X"22",X"3A",X"3C",X"86",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CD",X"D3",X"22",
		X"21",X"01",X"8B",X"11",X"20",X"00",X"3A",X"3D",X"86",X"E6",X"0F",X"CD",X"D3",X"22",X"3A",X"3D",
		X"86",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CD",X"D3",X"22",X"3A",X"3E",X"86",X"E6",
		X"0F",X"CD",X"D3",X"22",X"3A",X"3E",X"86",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CD",
		X"D3",X"22",X"C9",X"01",X"DC",X"22",X"81",X"4F",X"0A",X"77",X"19",X"C9",X"00",X"01",X"02",X"03",
		X"04",X"05",X"06",X"07",X"08",X"09",X"11",X"12",X"13",X"14",X"15",X"16",X"17",X"18",X"CD",X"26",
		X"09",X"D2",X"E0",X"09",X"CD",X"CE",X"08",X"D2",X"3F",X"24",X"FD",X"2A",X"DA",X"80",X"FD",X"66",
		X"02",X"FD",X"6E",X"01",X"E5",X"DD",X"E1",X"CD",X"07",X"17",X"CD",X"47",X"24",X"FD",X"36",X"0D",
		X"00",X"FD",X"CB",X"00",X"F6",X"FD",X"CB",X"0C",X"D6",X"DD",X"CB",X"00",X"EE",X"FD",X"CB",X"00",
		X"D6",X"3E",X"0A",X"CD",X"1F",X"08",X"DD",X"E5",X"CD",X"BC",X"09",X"FD",X"E1",X"DD",X"7E",X"0D",
		X"B7",X"C2",X"2E",X"24",X"FD",X"CB",X"00",X"4E",X"20",X"03",X"CD",X"47",X"23",X"CD",X"7B",X"16",
		X"FD",X"E5",X"CD",X"BC",X"09",X"18",X"E4",X"CD",X"06",X"19",X"CD",X"DF",X"23",X"CB",X"57",X"28",
		X"17",X"21",X"20",X"FD",X"FD",X"75",X"03",X"FD",X"74",X"04",X"FD",X"36",X"09",X"00",X"FD",X"36",
		X"0A",X"00",X"21",X"8A",X"24",X"C3",X"CC",X"23",X"CB",X"4F",X"28",X"17",X"FD",X"36",X"03",X"00",
		X"FD",X"36",X"04",X"00",X"21",X"20",X"FD",X"FD",X"75",X"09",X"FD",X"74",X"0A",X"21",X"8A",X"24",
		X"C3",X"CC",X"23",X"CB",X"47",X"28",X"17",X"21",X"E0",X"02",X"FD",X"75",X"03",X"FD",X"74",X"04",
		X"FD",X"36",X"09",X"00",X"FD",X"36",X"0A",X"00",X"21",X"8A",X"24",X"C3",X"CC",X"23",X"CB",X"5F",
		X"28",X"17",X"FD",X"36",X"03",X"00",X"FD",X"36",X"04",X"00",X"21",X"E0",X"02",X"FD",X"75",X"09",
		X"FD",X"74",X"0A",X"21",X"8A",X"24",X"C3",X"CC",X"23",X"FD",X"36",X"03",X"00",X"FD",X"36",X"04",
		X"00",X"FD",X"36",X"09",X"00",X"FD",X"36",X"0A",X"00",X"21",X"59",X"24",X"DD",X"75",X"05",X"DD",
		X"74",X"06",X"DD",X"36",X"04",X"01",X"FD",X"CB",X"00",X"96",X"DD",X"CB",X"00",X"E6",X"C9",X"CD",
		X"42",X"08",X"CB",X"77",X"28",X"2F",X"FD",X"7E",X"04",X"B7",X"20",X"18",X"FD",X"7E",X"0A",X"B7",
		X"20",X"12",X"CD",X"42",X"08",X"F6",X"08",X"E6",X"3F",X"FD",X"77",X"01",X"FD",X"CB",X"00",X"CE",
		X"78",X"E6",X"0A",X"C9",X"CD",X"42",X"08",X"F6",X"10",X"E6",X"3F",X"FD",X"77",X"01",X"FD",X"CB",
		X"00",X"CE",X"3E",X"00",X"C9",X"FD",X"7E",X"04",X"B7",X"20",X"E9",X"FD",X"7E",X"0A",X"B7",X"20",
		X"E3",X"3E",X"19",X"FD",X"77",X"01",X"FD",X"CB",X"00",X"CE",X"78",X"E6",X"05",X"C9",X"3E",X"05",
		X"CD",X"1F",X"08",X"01",X"07",X"01",X"CD",X"57",X"1F",X"CD",X"01",X"15",X"C3",X"FA",X"22",X"CD",
		X"36",X"0A",X"CD",X"BC",X"09",X"18",X"FB",X"21",X"8A",X"24",X"FD",X"75",X"05",X"FD",X"74",X"06",
		X"FD",X"36",X"04",X"01",X"FD",X"CB",X"00",X"E6",X"C9",X"00",X"00",X"01",X"00",X"00",X"05",X"05",
		X"03",X"32",X"00",X"05",X"05",X"03",X"32",X"01",X"05",X"05",X"03",X"32",X"02",X"05",X"05",X"03",
		X"32",X"03",X"05",X"05",X"03",X"32",X"04",X"05",X"05",X"03",X"32",X"05",X"05",X"05",X"03",X"32",
		X"06",X"05",X"05",X"03",X"32",X"07",X"00",X"01",X"5E",X"24",X"00",X"00",X"01",X"00",X"00",X"0E",
		X"0E",X"01",X"20",X"01",X"0E",X"0E",X"01",X"A0",X"01",X"0E",X"0E",X"01",X"21",X"01",X"0E",X"0E",
		X"01",X"A1",X"01",X"0E",X"0E",X"01",X"60",X"01",X"0E",X"0E",X"01",X"61",X"01",X"0E",X"0E",X"01",
		X"E0",X"01",X"0E",X"0E",X"01",X"E1",X"01",X"00",X"01",X"8F",X"24",X"2F",X"CD",X"26",X"09",X"D2",
		X"E0",X"09",X"CD",X"CE",X"08",X"D2",X"E2",X"25",X"FD",X"2A",X"DA",X"80",X"FD",X"66",X"02",X"FD",
		X"6E",X"01",X"E5",X"DD",X"E1",X"CD",X"EA",X"25",X"FD",X"36",X"0D",X"00",X"FD",X"CB",X"00",X"F6",
		X"FD",X"CB",X"0C",X"D6",X"DD",X"CB",X"00",X"EE",X"FD",X"CB",X"00",X"D6",X"FD",X"36",X"0B",X"00",
		X"3E",X"0A",X"CD",X"1F",X"08",X"DD",X"E5",X"CD",X"BC",X"09",X"FD",X"E1",X"DD",X"7E",X"0B",X"FE",
		X"06",X"38",X"03",X"C3",X"22",X"27",X"DD",X"7E",X"0D",X"B7",X"C2",X"D1",X"25",X"CD",X"18",X"25",
		X"FD",X"E5",X"CD",X"BC",X"09",X"C3",X"FA",X"24",X"DD",X"7E",X"0A",X"FE",X"16",X"30",X"1F",X"11",
		X"80",X"04",X"FD",X"72",X"04",X"FD",X"73",X"03",X"FD",X"36",X"0A",X"00",X"FD",X"36",X"09",X"00",
		X"3E",X"16",X"DD",X"77",X"0A",X"DD",X"34",X"0B",X"21",X"56",X"28",X"C3",X"BE",X"25",X"DD",X"7E",
		X"08",X"21",X"34",X"86",X"BE",X"38",X"20",X"11",X"80",X"04",X"FD",X"72",X"0A",X"FD",X"73",X"09",
		X"FD",X"36",X"04",X"00",X"FD",X"36",X"03",X"00",X"7E",X"3D",X"3D",X"DD",X"77",X"08",X"DD",X"34",
		X"0B",X"21",X"7C",X"28",X"C3",X"BE",X"25",X"DD",X"7E",X"0A",X"FE",X"D9",X"38",X"22",X"11",X"80",
		X"04",X"CD",X"BE",X"0F",X"FD",X"72",X"04",X"FD",X"73",X"03",X"FD",X"36",X"0A",X"00",X"FD",X"36",
		X"09",X"00",X"3E",X"D8",X"DD",X"77",X"0A",X"DD",X"34",X"0B",X"21",X"43",X"28",X"C3",X"BE",X"25",
		X"DD",X"7E",X"08",X"21",X"33",X"86",X"BE",X"30",X"24",X"11",X"80",X"04",X"CD",X"BE",X"0F",X"FD",
		X"72",X"0A",X"FD",X"73",X"09",X"FD",X"36",X"04",X"00",X"FD",X"36",X"03",X"00",X"7E",X"3C",X"3C",
		X"3C",X"DD",X"77",X"08",X"DD",X"34",X"0B",X"21",X"69",X"28",X"C3",X"BE",X"25",X"C9",X"DD",X"75",
		X"05",X"DD",X"74",X"06",X"DD",X"36",X"04",X"01",X"FD",X"CB",X"00",X"96",X"DD",X"CB",X"00",X"E6",
		X"C9",X"3E",X"05",X"CD",X"1F",X"08",X"01",X"05",X"01",X"CD",X"57",X"1F",X"CD",X"01",X"15",X"C3",
		X"C8",X"24",X"CD",X"36",X"0A",X"CD",X"BC",X"09",X"18",X"FB",X"CD",X"42",X"08",X"E6",X"03",X"28",
		X"0C",X"FE",X"01",X"28",X"4F",X"FE",X"02",X"CA",X"8C",X"26",X"C3",X"D7",X"26",X"3A",X"1A",X"82",
		X"FE",X"78",X"30",X"07",X"3A",X"1C",X"82",X"FE",X"78",X"38",X"DF",X"21",X"33",X"86",X"7E",X"3C",
		X"3C",X"FD",X"77",X"08",X"FD",X"36",X"0A",X"16",X"11",X"80",X"04",X"DD",X"72",X"04",X"DD",X"73",
		X"03",X"DD",X"36",X"0A",X"00",X"DD",X"36",X"09",X"00",X"21",X"56",X"28",X"FD",X"75",X"05",X"FD",
		X"74",X"06",X"FD",X"36",X"04",X"01",X"FD",X"CB",X"00",X"E6",X"3E",X"0A",X"DD",X"77",X"01",X"DD",
		X"CB",X"00",X"CE",X"C9",X"3A",X"1A",X"82",X"FE",X"78",X"38",X"08",X"3A",X"1C",X"82",X"FE",X"78",
		X"DA",X"EA",X"25",X"21",X"34",X"86",X"7E",X"3D",X"3D",X"FD",X"77",X"08",X"FD",X"36",X"0A",X"16",
		X"11",X"80",X"04",X"DD",X"72",X"0A",X"DD",X"73",X"09",X"DD",X"36",X"04",X"00",X"DD",X"36",X"03",
		X"00",X"21",X"7C",X"28",X"FD",X"75",X"05",X"FD",X"74",X"06",X"FD",X"36",X"04",X"01",X"FD",X"CB",
		X"00",X"E6",X"3E",X"0A",X"DD",X"77",X"01",X"DD",X"CB",X"00",X"CE",X"C9",X"3A",X"1A",X"82",X"FE",
		X"78",X"38",X"08",X"3A",X"1C",X"82",X"FE",X"78",X"D2",X"EA",X"25",X"21",X"34",X"86",X"7E",X"3D",
		X"3D",X"FD",X"77",X"08",X"FD",X"36",X"0A",X"D8",X"11",X"80",X"04",X"CD",X"BE",X"0F",X"DD",X"72",
		X"04",X"DD",X"73",X"03",X"DD",X"36",X"0A",X"00",X"DD",X"36",X"09",X"00",X"21",X"43",X"28",X"FD",
		X"75",X"05",X"FD",X"74",X"06",X"FD",X"36",X"04",X"01",X"FD",X"CB",X"00",X"E6",X"3E",X"0A",X"DD",
		X"77",X"01",X"DD",X"CB",X"00",X"CE",X"C9",X"3A",X"1A",X"82",X"FE",X"78",X"30",X"08",X"3A",X"1C",
		X"82",X"FE",X"78",X"D2",X"EA",X"25",X"21",X"33",X"86",X"7E",X"3C",X"3C",X"FD",X"77",X"08",X"FD",
		X"36",X"0A",X"D8",X"11",X"80",X"04",X"DD",X"36",X"04",X"00",X"DD",X"36",X"03",X"00",X"CD",X"BE",
		X"0F",X"DD",X"72",X"0A",X"DD",X"73",X"09",X"21",X"69",X"28",X"FD",X"75",X"05",X"FD",X"74",X"06",
		X"FD",X"36",X"04",X"01",X"FD",X"CB",X"00",X"E6",X"3E",X"0A",X"DD",X"77",X"01",X"DD",X"CB",X"00",
		X"CE",X"C9",X"CD",X"20",X"28",X"3E",X"0B",X"CD",X"1F",X"08",X"DD",X"7E",X"0D",X"B7",X"C2",X"32",
		X"28",X"FD",X"CB",X"00",X"4E",X"20",X"0B",X"FD",X"36",X"01",X"05",X"FD",X"CB",X"00",X"CE",X"CD",
		X"4F",X"27",X"CD",X"7B",X"16",X"FD",X"E5",X"CD",X"BC",X"09",X"FD",X"E1",X"C3",X"2A",X"27",X"CD",
		X"06",X"19",X"CD",X"14",X"28",X"FE",X"01",X"20",X"12",X"21",X"80",X"03",X"FD",X"75",X"03",X"FD",
		X"74",X"04",X"FD",X"36",X"09",X"00",X"FD",X"36",X"0A",X"00",X"C9",X"FE",X"03",X"20",X"13",X"21",
		X"80",X"03",X"FD",X"75",X"03",X"FD",X"74",X"04",X"21",X"80",X"FC",X"FD",X"75",X"09",X"FD",X"74",
		X"0A",X"C9",X"FE",X"02",X"20",X"12",X"FD",X"36",X"03",X"00",X"FD",X"36",X"04",X"00",X"21",X"80",
		X"FC",X"FD",X"75",X"09",X"FD",X"74",X"0A",X"C9",X"FE",X"06",X"20",X"10",X"21",X"80",X"FC",X"FD",
		X"75",X"03",X"FD",X"74",X"04",X"FD",X"75",X"09",X"FD",X"74",X"0A",X"C9",X"FE",X"04",X"20",X"12",
		X"21",X"80",X"FC",X"FD",X"75",X"03",X"FD",X"74",X"04",X"FD",X"36",X"09",X"00",X"FD",X"36",X"0A",
		X"00",X"C9",X"FE",X"0C",X"20",X"13",X"21",X"80",X"FC",X"FD",X"75",X"03",X"FD",X"74",X"04",X"21",
		X"80",X"03",X"FD",X"75",X"09",X"FD",X"74",X"0A",X"C9",X"FE",X"08",X"20",X"12",X"FD",X"36",X"03",
		X"00",X"FD",X"36",X"04",X"00",X"21",X"80",X"03",X"FD",X"75",X"09",X"FD",X"74",X"0A",X"C9",X"FE",
		X"09",X"20",X"10",X"21",X"80",X"03",X"FD",X"75",X"03",X"FD",X"74",X"04",X"FD",X"75",X"09",X"FD",
		X"74",X"0A",X"C9",X"FD",X"36",X"03",X"00",X"FD",X"36",X"04",X"00",X"FD",X"36",X"09",X"00",X"FD",
		X"36",X"0A",X"00",X"C9",X"CD",X"42",X"08",X"FE",X"7F",X"38",X"02",X"78",X"C9",X"E6",X"0F",X"C9",
		X"21",X"8F",X"28",X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",X"36",X"04",X"01",X"DD",X"CB",X"00",
		X"E6",X"C9",X"3E",X"05",X"CD",X"1F",X"08",X"01",X"01",X"02",X"CD",X"57",X"1F",X"CD",X"01",X"15",
		X"C3",X"C8",X"24",X"00",X"00",X"01",X"00",X"00",X"0E",X"09",X"03",X"26",X"04",X"0E",X"09",X"03",
		X"25",X"04",X"00",X"01",X"48",X"28",X"00",X"00",X"01",X"00",X"00",X"0E",X"09",X"04",X"E6",X"04",
		X"0E",X"09",X"04",X"E5",X"04",X"00",X"01",X"5B",X"28",X"00",X"00",X"01",X"00",X"00",X"09",X"0E",
		X"04",X"E3",X"04",X"09",X"0E",X"04",X"E4",X"04",X"00",X"01",X"6E",X"28",X"00",X"00",X"01",X"00",
		X"00",X"09",X"0E",X"04",X"23",X"04",X"09",X"0E",X"04",X"24",X"04",X"00",X"01",X"81",X"28",X"00",
		X"00",X"01",X"00",X"00",X"0C",X"0C",X"02",X"1F",X"00",X"0C",X"0C",X"02",X"1E",X"01",X"0C",X"0C",
		X"02",X"1D",X"02",X"0C",X"0C",X"02",X"1E",X"03",X"0C",X"0C",X"02",X"1F",X"04",X"0C",X"0C",X"02",
		X"1E",X"05",X"0C",X"0C",X"02",X"1D",X"06",X"0C",X"0C",X"02",X"1E",X"07",X"00",X"01",X"94",X"28",
		X"CD",X"26",X"09",X"D2",X"E0",X"09",X"CD",X"CE",X"08",X"D2",X"32",X"2A",X"FD",X"2A",X"DA",X"80",
		X"FD",X"66",X"02",X"FD",X"6E",X"01",X"E5",X"DD",X"E1",X"CD",X"07",X"17",X"CD",X"3A",X"2A",X"FD",
		X"36",X"0D",X"00",X"FD",X"CB",X"00",X"F6",X"FD",X"CB",X"0C",X"D6",X"DD",X"CB",X"00",X"EE",X"FD",
		X"CB",X"00",X"D6",X"3E",X"0A",X"CD",X"1F",X"08",X"DD",X"E5",X"CD",X"BC",X"09",X"FD",X"E1",X"DD",
		X"CB",X"0D",X"4E",X"C2",X"21",X"2A",X"DD",X"CB",X"0D",X"76",X"C4",X"20",X"29",X"FD",X"CB",X"00",
		X"4E",X"20",X"03",X"CD",X"63",X"29",X"CD",X"7B",X"16",X"FD",X"E5",X"CD",X"BC",X"09",X"18",X"DD",
		X"3E",X"0C",X"CD",X"1F",X"08",X"01",X"01",X"01",X"CD",X"57",X"1F",X"DD",X"36",X"0D",X"00",X"CD",
		X"42",X"08",X"F6",X"40",X"E6",X"7F",X"FD",X"77",X"01",X"FD",X"CB",X"00",X"CE",X"FD",X"36",X"03",
		X"00",X"FD",X"36",X"04",X"00",X"FD",X"36",X"09",X"00",X"FD",X"36",X"0A",X"00",X"21",X"4C",X"2A",
		X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",X"36",X"04",X"01",X"FD",X"CB",X"00",X"96",X"DD",X"CB",
		X"00",X"E6",X"C9",X"CD",X"06",X"19",X"CD",X"FB",X"29",X"CB",X"57",X"28",X"17",X"21",X"10",X"FE",
		X"FD",X"75",X"03",X"FD",X"74",X"04",X"FD",X"36",X"09",X"00",X"FD",X"36",X"0A",X"00",X"21",X"7D",
		X"2A",X"C3",X"E8",X"29",X"CB",X"4F",X"28",X"17",X"FD",X"36",X"03",X"00",X"FD",X"36",X"04",X"00",
		X"21",X"10",X"FE",X"FD",X"75",X"09",X"FD",X"74",X"0A",X"21",X"7D",X"2A",X"C3",X"E8",X"29",X"CB",
		X"47",X"28",X"17",X"21",X"F0",X"01",X"FD",X"75",X"03",X"FD",X"74",X"04",X"FD",X"36",X"09",X"00",
		X"FD",X"36",X"0A",X"00",X"21",X"7D",X"2A",X"C3",X"E8",X"29",X"CB",X"5F",X"28",X"17",X"21",X"F0",
		X"01",X"FD",X"36",X"03",X"00",X"FD",X"36",X"04",X"00",X"FD",X"75",X"09",X"FD",X"74",X"0A",X"21",
		X"7D",X"2A",X"C3",X"E8",X"29",X"FD",X"36",X"03",X"00",X"FD",X"36",X"04",X"00",X"FD",X"36",X"09",
		X"00",X"FD",X"36",X"0A",X"00",X"21",X"4C",X"2A",X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",X"36",
		X"04",X"01",X"FD",X"CB",X"00",X"96",X"DD",X"CB",X"00",X"E6",X"C9",X"CD",X"42",X"08",X"CB",X"77",
		X"28",X"12",X"CD",X"42",X"08",X"E6",X"08",X"F6",X"3F",X"FD",X"77",X"01",X"FD",X"CB",X"00",X"CE",
		X"78",X"E6",X"0A",X"C9",X"3E",X"19",X"FD",X"77",X"01",X"FD",X"CB",X"00",X"CE",X"78",X"E6",X"05",
		X"C9",X"3E",X"05",X"CD",X"1F",X"08",X"01",X"04",X"01",X"CD",X"57",X"1F",X"CD",X"01",X"15",X"C3",
		X"CC",X"28",X"CD",X"36",X"0A",X"CD",X"BC",X"09",X"18",X"FB",X"21",X"7D",X"2A",X"FD",X"75",X"05",
		X"FD",X"74",X"06",X"FD",X"36",X"04",X"01",X"FD",X"CB",X"00",X"E6",X"C9",X"00",X"00",X"01",X"00",
		X"00",X"05",X"05",X"04",X"32",X"00",X"05",X"05",X"04",X"32",X"01",X"05",X"05",X"04",X"32",X"02",
		X"05",X"05",X"04",X"32",X"03",X"05",X"05",X"04",X"32",X"04",X"05",X"05",X"04",X"32",X"05",X"05",
		X"05",X"04",X"32",X"06",X"05",X"05",X"04",X"32",X"07",X"00",X"01",X"51",X"2A",X"00",X"00",X"01",
		X"00",X"00",X"0E",X"0E",X"01",X"31",X"02",X"0E",X"0E",X"01",X"30",X"02",X"0E",X"0E",X"01",X"2F",
		X"02",X"0E",X"0E",X"01",X"70",X"02",X"00",X"01",X"82",X"2A",X"CD",X"65",X"34",X"CD",X"D3",X"06",
		X"CD",X"89",X"06",X"CF",X"58",X"80",X"42",X"4F",X"4E",X"55",X"53",X"20",X"52",X"4F",X"4F",X"4D",
		X"00",X"CF",X"40",X"F8",X"41",X"4C",X"4C",X"20",X"4E",X"55",X"4D",X"42",X"45",X"52",X"53",X"20",
		X"58",X"20",X"31",X"30",X"30",X"00",X"CD",X"85",X"08",X"DD",X"21",X"12",X"82",X"FD",X"21",X"9A",
		X"81",X"21",X"2A",X"85",X"36",X"00",X"21",X"2B",X"85",X"36",X"00",X"CD",X"C2",X"3C",X"DD",X"CB",
		X"00",X"D6",X"AF",X"DD",X"77",X"0D",X"DD",X"CB",X"0C",X"C6",X"CD",X"7B",X"2C",X"CD",X"F0",X"2C",
		X"DD",X"CB",X"00",X"F6",X"3E",X"01",X"32",X"44",X"86",X"FD",X"21",X"9A",X"81",X"DD",X"CB",X"00",
		X"6E",X"20",X"29",X"3A",X"67",X"85",X"FE",X"3D",X"28",X"22",X"DD",X"36",X"03",X"05",X"DD",X"CB",
		X"00",X"EE",X"FD",X"CB",X"00",X"7E",X"28",X"0B",X"3E",X"08",X"CD",X"1F",X"08",X"FD",X"CB",X"00",
		X"BE",X"18",X"09",X"3E",X"09",X"CD",X"1F",X"08",X"FD",X"CB",X"00",X"FE",X"DD",X"7E",X"0D",X"CB",
		X"57",X"C2",X"0E",X"2C",X"FD",X"CB",X"00",X"4E",X"20",X"14",X"FD",X"CB",X"00",X"F6",X"FD",X"36",
		X"01",X"05",X"FD",X"CB",X"00",X"CE",X"3E",X"01",X"32",X"44",X"86",X"CD",X"88",X"19",X"3A",X"23",
		X"85",X"E6",X"3C",X"21",X"2B",X"85",X"46",X"77",X"A8",X"C4",X"DF",X"3C",X"DD",X"CB",X"00",X"E6",
		X"FD",X"7E",X"0D",X"FE",X"2C",X"20",X"0B",X"21",X"2F",X"85",X"34",X"3E",X"0E",X"CD",X"1F",X"08",
		X"18",X"16",X"FE",X"01",X"38",X"2F",X"FE",X"09",X"30",X"2B",X"4F",X"06",X"02",X"CD",X"57",X"1F",
		X"CD",X"89",X"06",X"3E",X"06",X"CD",X"1F",X"08",X"FD",X"36",X"0D",X"00",X"DD",X"7E",X"08",X"C6",
		X"08",X"67",X"DD",X"7E",X"0A",X"C6",X"08",X"6F",X"CD",X"BF",X"04",X"36",X"10",X"FD",X"36",X"02",
		X"05",X"FD",X"CB",X"00",X"D6",X"01",X"00",X"00",X"11",X"00",X"00",X"3A",X"23",X"85",X"67",X"CD",
		X"7B",X"3C",X"CD",X"8C",X"3C",X"CD",X"9A",X"3C",X"CD",X"AC",X"3C",X"FD",X"70",X"04",X"FD",X"71",
		X"03",X"FD",X"72",X"0A",X"FD",X"73",X"09",X"FD",X"CB",X"00",X"56",X"28",X"13",X"FD",X"CB",X"02",
		X"56",X"28",X"08",X"3E",X"FF",X"32",X"04",X"A8",X"C3",X"E0",X"2B",X"3E",X"00",X"32",X"04",X"A8",
		X"3A",X"34",X"86",X"47",X"DD",X"7E",X"08",X"B8",X"38",X"03",X"DD",X"70",X"08",X"3A",X"33",X"86",
		X"47",X"DD",X"7E",X"08",X"B8",X"30",X"03",X"DD",X"70",X"08",X"DD",X"7E",X"0A",X"FE",X"17",X"38",
		X"04",X"FE",X"D7",X"38",X"06",X"CD",X"36",X"0A",X"CD",X"BC",X"09",X"C3",X"F9",X"2A",X"DD",X"CB",
		X"0C",X"86",X"3A",X"29",X"85",X"C6",X"99",X"27",X"32",X"29",X"85",X"3E",X"05",X"CD",X"1F",X"08",
		X"AF",X"FD",X"77",X"03",X"FD",X"77",X"04",X"FD",X"77",X"09",X"FD",X"77",X"0A",X"DD",X"21",X"12",
		X"82",X"DD",X"CB",X"00",X"B6",X"DD",X"CB",X"00",X"A6",X"21",X"E5",X"15",X"DD",X"75",X"05",X"DD",
		X"74",X"06",X"DD",X"36",X"04",X"01",X"DD",X"CB",X"00",X"E6",X"DD",X"CB",X"00",X"66",X"28",X"02",
		X"18",X"F8",X"AF",X"FD",X"77",X"03",X"FD",X"77",X"04",X"FD",X"77",X"09",X"FD",X"77",X"0A",X"DD",
		X"77",X"08",X"DD",X"77",X"0A",X"FD",X"77",X"06",X"FD",X"77",X"0C",X"CD",X"36",X"0A",X"DD",X"21",
		X"12",X"82",X"DD",X"36",X"0B",X"FF",X"CD",X"BC",X"09",X"18",X"FB",X"DD",X"36",X"08",X"7A",X"DD",
		X"36",X"0A",X"D7",X"01",X"00",X"00",X"11",X"00",X"02",X"CD",X"BE",X"0F",X"FD",X"70",X"04",X"FD",
		X"71",X"03",X"FD",X"72",X"0A",X"FD",X"73",X"09",X"3A",X"2B",X"85",X"CB",X"D7",X"32",X"2B",X"85",
		X"CD",X"DF",X"3C",X"DD",X"CB",X"00",X"E6",X"FD",X"36",X"01",X"05",X"FD",X"CB",X"00",X"CE",X"3E",
		X"08",X"CD",X"1F",X"08",X"FD",X"CB",X"00",X"4E",X"28",X"0A",X"DD",X"7E",X"0A",X"FE",X"7D",X"30",
		X"F3",X"C3",X"DE",X"2C",X"FD",X"36",X"01",X"05",X"FD",X"CB",X"00",X"CE",X"3E",X"09",X"CD",X"1F",
		X"08",X"FD",X"CB",X"00",X"4E",X"28",X"D0",X"DD",X"7E",X"0A",X"FE",X"7D",X"30",X"F3",X"11",X"00",
		X"00",X"FD",X"72",X"0A",X"FD",X"73",X"09",X"FD",X"36",X"07",X"3D",X"DD",X"CB",X"00",X"A6",X"C9",
		X"E7",X"1D",X"02",X"01",X"3E",X"1E",X"B7",X"C8",X"47",X"CD",X"27",X"2D",X"CD",X"42",X"08",X"E6",
		X"07",X"FE",X"01",X"28",X"01",X"3C",X"77",X"C5",X"06",X"14",X"C5",X"06",X"FF",X"10",X"FE",X"C1",
		X"10",X"F8",X"3E",X"06",X"CD",X"1F",X"08",X"C1",X"10",X"DF",X"CD",X"27",X"2D",X"3E",X"2C",X"77",
		X"CD",X"27",X"2D",X"3E",X"2C",X"77",X"C9",X"CD",X"42",X"08",X"FE",X"3A",X"38",X"F9",X"FE",X"C8",
		X"30",X"F5",X"67",X"CD",X"42",X"08",X"FE",X"3A",X"38",X"F9",X"FE",X"C8",X"30",X"F5",X"6F",X"3E",
		X"5B",X"BC",X"30",X"12",X"3E",X"98",X"BC",X"38",X"0D",X"3E",X"6B",X"BD",X"30",X"08",X"3E",X"A8",
		X"BD",X"38",X"03",X"C3",X"27",X"2D",X"CD",X"BF",X"04",X"7E",X"FE",X"10",X"20",X"C9",X"E5",X"23",
		X"7E",X"FE",X"10",X"C2",X"85",X"2D",X"2B",X"2B",X"7E",X"FE",X"10",X"C2",X"85",X"2D",X"23",X"11",
		X"20",X"00",X"19",X"7E",X"FE",X"10",X"C2",X"85",X"2D",X"E1",X"E5",X"ED",X"52",X"7E",X"FE",X"10",
		X"C2",X"85",X"2D",X"E1",X"C9",X"E1",X"C3",X"27",X"2D",X"3A",X"46",X"86",X"B7",X"20",X"08",X"3A",
		X"00",X"98",X"CB",X"5F",X"CA",X"D1",X"4F",X"3A",X"EE",X"80",X"B7",X"C8",X"FE",X"01",X"28",X"07",
		X"3A",X"28",X"85",X"CB",X"77",X"20",X"08",X"3A",X"28",X"85",X"CB",X"47",X"20",X"12",X"C9",X"CD",
		X"1B",X"11",X"3E",X"02",X"32",X"56",X"85",X"21",X"39",X"85",X"CD",X"27",X"2F",X"C3",X"C5",X"2D",
		X"3E",X"01",X"32",X"56",X"85",X"3E",X"0A",X"CD",X"1B",X"11",X"21",X"29",X"85",X"CD",X"27",X"2F",
		X"CD",X"60",X"1A",X"21",X"00",X"00",X"22",X"2B",X"81",X"22",X"2D",X"81",X"22",X"2F",X"81",X"22",
		X"E6",X"80",X"21",X"00",X"01",X"22",X"30",X"85",X"CD",X"E5",X"2E",X"21",X"00",X"01",X"22",X"30",
		X"85",X"CD",X"E5",X"2E",X"AF",X"32",X"55",X"85",X"3E",X"01",X"32",X"59",X"85",X"AF",X"32",X"38",
		X"86",X"32",X"39",X"86",X"32",X"3A",X"86",X"CD",X"82",X"05",X"CD",X"07",X"2F",X"CD",X"47",X"2F",
		X"3E",X"0A",X"CD",X"10",X"0A",X"CD",X"69",X"0A",X"AF",X"CD",X"1F",X"08",X"3A",X"29",X"85",X"B7",
		X"CC",X"65",X"2E",X"CD",X"E5",X"2E",X"3A",X"29",X"85",X"B7",X"C2",X"07",X"2E",X"CD",X"E5",X"2E",
		X"3A",X"29",X"85",X"B7",X"20",X"D1",X"2A",X"39",X"86",X"ED",X"4B",X"3B",X"86",X"09",X"22",X"3B",
		X"86",X"2A",X"3D",X"86",X"23",X"3A",X"56",X"85",X"FE",X"02",X"20",X"01",X"23",X"22",X"3D",X"86",
		X"3E",X"01",X"32",X"46",X"86",X"CD",X"AC",X"1D",X"CD",X"E5",X"2E",X"CD",X"AC",X"1D",X"AF",X"32",
		X"46",X"86",X"C3",X"2E",X"1A",X"3E",X"05",X"CD",X"10",X"0A",X"3E",X"00",X"32",X"32",X"85",X"CF",
		X"28",X"68",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"00",X"CF",X"28",X"70",X"20",X"20",X"50",X"4C",
		X"41",X"59",X"45",X"52",X"20",X"20",X"20",X"47",X"41",X"4D",X"45",X"20",X"4F",X"56",X"45",X"52",
		X"20",X"20",X"00",X"CF",X"28",X"78",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"00",X"21",X"70",X"70",
		X"11",X"59",X"85",X"06",X"01",X"CD",X"27",X"05",X"06",X"32",X"3E",X"FD",X"32",X"40",X"86",X"3E",
		X"03",X"CD",X"10",X"0A",X"10",X"F4",X"C9",X"3A",X"01",X"98",X"2F",X"E6",X"01",X"28",X"03",X"36",
		X"05",X"C9",X"36",X"03",X"C9",X"D9",X"3A",X"59",X"85",X"3C",X"FE",X"02",X"28",X"02",X"3E",X"01",
		X"32",X"59",X"85",X"21",X"29",X"85",X"11",X"39",X"85",X"06",X"10",X"1A",X"4E",X"EB",X"12",X"71",
		X"EB",X"23",X"13",X"10",X"F6",X"D9",X"C9",X"3A",X"59",X"85",X"FE",X"02",X"20",X"10",X"3A",X"02",
		X"98",X"E6",X"08",X"20",X"09",X"3E",X"FF",X"32",X"07",X"A8",X"32",X"06",X"A8",X"C9",X"3E",X"00",
		X"32",X"07",X"A8",X"32",X"06",X"A8",X"C9",X"CD",X"D7",X"2E",X"23",X"36",X"00",X"23",X"36",X"00",
		X"23",X"36",X"0F",X"23",X"36",X"0F",X"23",X"36",X"01",X"23",X"36",X"02",X"21",X"32",X"85",X"36",
		X"00",X"3E",X"00",X"32",X"46",X"86",X"C9",X"AF",X"32",X"57",X"85",X"32",X"53",X"85",X"32",X"58",
		X"85",X"3E",X"05",X"32",X"78",X"85",X"CD",X"65",X"34",X"CD",X"89",X"06",X"FD",X"21",X"6D",X"38",
		X"CD",X"A4",X"09",X"3E",X"28",X"CD",X"10",X"0A",X"CD",X"90",X"2F",X"DD",X"21",X"12",X"82",X"DD",
		X"7E",X"00",X"B7",X"C8",X"3A",X"55",X"85",X"B7",X"C4",X"89",X"2D",X"3A",X"53",X"85",X"B7",X"C4",
		X"89",X"06",X"3A",X"58",X"85",X"FE",X"02",X"CA",X"61",X"3F",X"CD",X"BC",X"09",X"C3",X"6B",X"2F",
		X"CD",X"83",X"30",X"E5",X"7E",X"B7",X"28",X"11",X"47",X"C5",X"FD",X"21",X"B2",X"12",X"CD",X"A4",
		X"09",X"3E",X"0A",X"CD",X"10",X"0A",X"C1",X"10",X"F0",X"E1",X"23",X"E5",X"7E",X"B7",X"28",X"11",
		X"47",X"C5",X"FD",X"21",X"2B",X"16",X"CD",X"A4",X"09",X"3E",X"0A",X"CD",X"10",X"0A",X"C1",X"10",
		X"F0",X"E1",X"23",X"E5",X"7E",X"B7",X"28",X"11",X"47",X"C5",X"FD",X"21",X"30",X"18",X"CD",X"A4",
		X"09",X"3E",X"0A",X"CD",X"10",X"0A",X"C1",X"10",X"F0",X"E1",X"23",X"E5",X"7E",X"B7",X"28",X"11",
		X"47",X"C5",X"FD",X"21",X"EE",X"22",X"CD",X"A4",X"09",X"3E",X"0A",X"CD",X"10",X"0A",X"C1",X"10",
		X"F0",X"E1",X"23",X"E5",X"7E",X"B7",X"28",X"11",X"47",X"C5",X"FD",X"21",X"BC",X"24",X"CD",X"A4",
		X"09",X"3E",X"0A",X"CD",X"10",X"0A",X"C1",X"10",X"F0",X"E1",X"23",X"E5",X"7E",X"B7",X"28",X"11",
		X"47",X"C5",X"FD",X"21",X"C0",X"28",X"CD",X"A4",X"09",X"3E",X"0A",X"CD",X"10",X"0A",X"C1",X"10",
		X"F0",X"E1",X"23",X"E5",X"7E",X"B7",X"28",X"11",X"47",X"C5",X"FD",X"21",X"AE",X"45",X"CD",X"A4",
		X"09",X"3E",X"0A",X"CD",X"10",X"0A",X"C1",X"10",X"F0",X"E1",X"23",X"E5",X"7E",X"B7",X"28",X"11",
		X"47",X"C5",X"FD",X"21",X"50",X"47",X"CD",X"A4",X"09",X"3E",X"0A",X"CD",X"10",X"0A",X"C1",X"10",
		X"F0",X"E1",X"23",X"E5",X"7E",X"B7",X"28",X"11",X"47",X"C5",X"FD",X"21",X"EA",X"48",X"CD",X"A4",
		X"09",X"3E",X"0A",X"CD",X"10",X"0A",X"C1",X"10",X"F0",X"E1",X"23",X"E5",X"7E",X"B7",X"28",X"11",
		X"47",X"C5",X"FD",X"21",X"ED",X"4C",X"CD",X"A4",X"09",X"3E",X"0A",X"CD",X"10",X"0A",X"C1",X"10",
		X"F0",X"E1",X"C9",X"21",X"A2",X"30",X"3A",X"2E",X"85",X"BE",X"28",X"14",X"38",X"0C",X"3E",X"FF",
		X"BE",X"28",X"07",X"11",X"0B",X"00",X"19",X"C3",X"86",X"30",X"11",X"0B",X"00",X"B7",X"ED",X"52",
		X"23",X"C9",X"01",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"03",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"05",X"00",
		X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"04",
		X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"09",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0B",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"03",X"00",X"0F",X"00",X"00",X"00",
		X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",
		X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"12",X"07",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"13",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"00",X"00",X"00",X"14",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"15",X"01",
		X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"16",X"01",X"01",X"00",X"01",X"01",X"01",
		X"01",X"01",X"00",X"00",X"17",X"01",X"01",X"01",X"00",X"01",X"01",X"01",X"01",X"00",X"00",X"18",
		X"01",X"01",X"01",X"01",X"00",X"01",X"01",X"01",X"00",X"00",X"19",X"01",X"01",X"01",X"01",X"01",
		X"00",X"01",X"01",X"00",X"00",X"1A",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"01",X"00",X"00",
		X"1B",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"1C",X"00",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"00",X"00",X"1D",X"01",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"00",
		X"00",X"1E",X"01",X"01",X"00",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"1F",X"01",X"01",X"01",
		X"00",X"01",X"01",X"01",X"01",X"00",X"00",X"20",X"01",X"01",X"01",X"01",X"00",X"01",X"01",X"01",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"64",X"3A",X"40",X"86",X"FE",X"FF",X"28",
		X"0B",X"FE",X"FE",X"28",X"2F",X"FE",X"FD",X"28",X"48",X"C3",X"86",X"32",X"AF",X"32",X"40",X"86",
		X"21",X"41",X"86",X"34",X"3A",X"41",X"86",X"21",X"07",X"90",X"06",X"07",X"CD",X"76",X"32",X"21",
		X"39",X"90",X"06",X"01",X"CD",X"76",X"32",X"3A",X"41",X"86",X"21",X"1B",X"90",X"06",X"07",X"CD",
		X"76",X"32",X"18",X"42",X"AF",X"32",X"40",X"86",X"21",X"41",X"86",X"34",X"3A",X"41",X"86",X"21",
		X"07",X"90",X"06",X"0C",X"CD",X"7D",X"32",X"21",X"39",X"90",X"06",X"01",X"CD",X"76",X"32",X"18",
		X"25",X"AF",X"32",X"40",X"86",X"21",X"41",X"86",X"34",X"3A",X"41",X"86",X"21",X"05",X"90",X"06",
		X"1C",X"CD",X"76",X"32",X"18",X"10",X"77",X"23",X"23",X"3C",X"10",X"FA",X"C9",X"77",X"23",X"23",
		X"23",X"23",X"3C",X"10",X"F8",X"C9",X"21",X"9A",X"81",X"CB",X"76",X"CA",X"6A",X"33",X"CB",X"B6",
		X"21",X"33",X"86",X"34",X"34",X"7E",X"FE",X"78",X"38",X"08",X"DD",X"21",X"12",X"82",X"DD",X"CB",
		X"0D",X"D6",X"21",X"2E",X"86",X"34",X"7E",X"2A",X"2F",X"86",X"E6",X"03",X"20",X"09",X"11",X"20",
		X"00",X"B7",X"ED",X"52",X"22",X"2F",X"86",X"06",X"1A",X"C6",X"3D",X"4F",X"3A",X"32",X"85",X"B7",
		X"28",X"32",X"FE",X"01",X"28",X"20",X"FE",X"02",X"28",X"0E",X"7E",X"FE",X"70",X"38",X"31",X"FE",
		X"74",X"30",X"2D",X"CD",X"58",X"0E",X"18",X"28",X"7E",X"FE",X"60",X"38",X"23",X"FE",X"64",X"30",
		X"1F",X"CD",X"58",X"0E",X"18",X"1A",X"7E",X"FE",X"88",X"38",X"15",X"FE",X"8C",X"30",X"11",X"CD",
		X"58",X"0E",X"18",X"0C",X"7E",X"FE",X"38",X"38",X"07",X"FE",X"3C",X"30",X"03",X"CD",X"58",X"0E",
		X"71",X"23",X"10",X"B8",X"21",X"34",X"86",X"35",X"35",X"21",X"2E",X"86",X"7E",X"2A",X"31",X"86",
		X"E6",X"03",X"20",X"07",X"11",X"20",X"00",X"19",X"22",X"31",X"86",X"06",X"1A",X"4F",X"3E",X"43",
		X"99",X"4F",X"3A",X"32",X"85",X"B7",X"28",X"32",X"FE",X"01",X"28",X"20",X"FE",X"02",X"28",X"0E",
		X"7E",X"FE",X"70",X"38",X"31",X"FE",X"74",X"30",X"2D",X"CD",X"0F",X"0E",X"18",X"28",X"7E",X"FE",
		X"60",X"38",X"23",X"FE",X"64",X"30",X"1F",X"CD",X"0F",X"0E",X"18",X"1A",X"7E",X"FE",X"88",X"38",
		X"15",X"FE",X"8C",X"30",X"11",X"CD",X"0F",X"0E",X"18",X"0C",X"7E",X"FE",X"38",X"38",X"07",X"FE",
		X"3C",X"30",X"03",X"CD",X"0F",X"0E",X"71",X"23",X"10",X"B8",X"3A",X"12",X"82",X"CB",X"77",X"C8",
		X"21",X"2D",X"86",X"34",X"7E",X"E6",X"03",X"CA",X"87",X"33",X"FE",X"01",X"CA",X"A1",X"33",X"FE",
		X"02",X"CA",X"E2",X"33",X"C3",X"B6",X"33",X"21",X"60",X"88",X"3E",X"00",X"32",X"35",X"86",X"06",
		X"5F",X"CD",X"F7",X"33",X"10",X"FB",X"21",X"C0",X"88",X"06",X"5F",X"CD",X"F7",X"33",X"10",X"FB",
		X"C9",X"21",X"20",X"89",X"06",X"7F",X"CD",X"F7",X"33",X"10",X"FB",X"21",X"A0",X"89",X"06",X"5F",
		X"CD",X"F7",X"33",X"10",X"FB",X"C9",X"21",X"00",X"8A",X"06",X"5F",X"CD",X"F7",X"33",X"10",X"FB",
		X"21",X"60",X"8A",X"06",X"7F",X"CD",X"F7",X"33",X"10",X"FB",X"3A",X"35",X"86",X"32",X"2C",X"85",
		X"B7",X"C0",X"21",X"3F",X"86",X"3E",X"FF",X"BE",X"C8",X"34",X"3E",X"05",X"BE",X"C0",X"3E",X"FF",
		X"77",X"C9",X"21",X"E0",X"8A",X"06",X"5F",X"CD",X"F7",X"33",X"10",X"FB",X"21",X"40",X"8B",X"06",
		X"5F",X"CD",X"F7",X"33",X"10",X"FB",X"C9",X"3A",X"32",X"85",X"B7",X"28",X"20",X"FE",X"01",X"28",
		X"34",X"FE",X"02",X"28",X"48",X"23",X"7E",X"FE",X"70",X"D8",X"FE",X"74",X"D0",X"3C",X"FE",X"74",
		X"20",X"02",X"3E",X"70",X"77",X"3A",X"35",X"86",X"3C",X"32",X"35",X"86",X"C9",X"23",X"7E",X"FE",
		X"38",X"D8",X"FE",X"3C",X"D0",X"3C",X"FE",X"3C",X"20",X"02",X"3E",X"38",X"77",X"3A",X"35",X"86",
		X"3C",X"32",X"35",X"86",X"C9",X"23",X"7E",X"FE",X"88",X"D8",X"FE",X"8C",X"D0",X"3C",X"FE",X"8C",
		X"20",X"02",X"3E",X"88",X"77",X"3A",X"35",X"86",X"3C",X"32",X"35",X"86",X"C9",X"23",X"7E",X"FE",
		X"60",X"D8",X"FE",X"64",X"D0",X"3C",X"FE",X"64",X"20",X"02",X"3E",X"60",X"77",X"3A",X"35",X"86",
		X"3C",X"32",X"35",X"86",X"C9",X"3E",X"00",X"32",X"3F",X"86",X"32",X"35",X"86",X"3E",X"14",X"32",
		X"33",X"86",X"3E",X"DC",X"32",X"34",X"86",X"21",X"A3",X"8B",X"22",X"2F",X"86",X"21",X"43",X"88",
		X"22",X"31",X"86",X"3E",X"FF",X"32",X"2E",X"86",X"21",X"48",X"86",X"3A",X"2E",X"85",X"E6",X"07",
		X"28",X"1A",X"FE",X"01",X"28",X"1E",X"FE",X"02",X"28",X"22",X"FE",X"03",X"28",X"26",X"FE",X"04",
		X"28",X"2A",X"FE",X"05",X"28",X"2E",X"FE",X"06",X"28",X"32",X"18",X"38",X"36",X"00",X"E7",X"1D",
		X"02",X"00",X"18",X"38",X"36",X"01",X"E7",X"1D",X"02",X"01",X"18",X"30",X"36",X"02",X"E7",X"1D",
		X"02",X"02",X"18",X"28",X"36",X"03",X"E7",X"1D",X"02",X"03",X"18",X"20",X"36",X"04",X"E7",X"1D",
		X"02",X"04",X"18",X"18",X"36",X"05",X"E7",X"1D",X"02",X"05",X"18",X"10",X"36",X"06",X"E7",X"1D",
		X"02",X"06",X"18",X"08",X"36",X"07",X"E7",X"1D",X"02",X"07",X"18",X"00",X"AF",X"32",X"58",X"85",
		X"CD",X"9F",X"35",X"3E",X"40",X"21",X"42",X"88",X"06",X"1B",X"77",X"23",X"10",X"FC",X"21",X"A2",
		X"8B",X"06",X"1B",X"77",X"23",X"10",X"FC",X"3E",X"40",X"21",X"42",X"88",X"11",X"20",X"00",X"06",
		X"1C",X"77",X"19",X"10",X"FC",X"21",X"42",X"88",X"11",X"1B",X"00",X"19",X"11",X"20",X"00",X"06",
		X"1C",X"77",X"19",X"10",X"FC",X"C9",X"3A",X"2C",X"85",X"B7",X"C8",X"47",X"CD",X"67",X"35",X"CD",
		X"42",X"08",X"E6",X"03",X"4F",X"3A",X"32",X"85",X"B7",X"28",X"0C",X"FE",X"01",X"28",X"0C",X"FE",
		X"02",X"28",X"0C",X"3E",X"70",X"18",X"0A",X"3E",X"38",X"18",X"06",X"3E",X"88",X"18",X"02",X"3E",
		X"60",X"81",X"77",X"C5",X"06",X"14",X"C5",X"06",X"FF",X"10",X"FE",X"C1",X"10",X"F8",X"3E",X"06",
		X"CD",X"1F",X"08",X"C1",X"10",X"C6",X"C9",X"CD",X"42",X"08",X"FE",X"26",X"38",X"F9",X"FE",X"DC",
		X"30",X"F5",X"67",X"CD",X"42",X"08",X"FE",X"26",X"38",X"F9",X"FE",X"DC",X"30",X"F5",X"6F",X"3E",
		X"5B",X"BC",X"30",X"12",X"3E",X"98",X"BC",X"38",X"0D",X"3E",X"6B",X"BD",X"30",X"08",X"3E",X"A8",
		X"BD",X"38",X"03",X"C3",X"67",X"35",X"CD",X"BF",X"04",X"7E",X"FE",X"10",X"C8",X"18",X"C8",X"3A",
		X"55",X"85",X"B7",X"C0",X"21",X"CB",X"35",X"3A",X"2E",X"85",X"BE",X"28",X"14",X"38",X"0C",X"3E",
		X"FF",X"BE",X"28",X"07",X"11",X"04",X"00",X"19",X"C3",X"A7",X"35",X"11",X"04",X"00",X"B7",X"ED",
		X"52",X"23",X"01",X"03",X"00",X"11",X"49",X"85",X"ED",X"B0",X"C9",X"01",X"07",X"00",X"02",X"02",
		X"07",X"00",X"02",X"03",X"07",X"00",X"02",X"04",X"07",X"00",X"02",X"05",X"07",X"00",X"02",X"06",
		X"07",X"00",X"02",X"07",X"07",X"00",X"02",X"08",X"07",X"00",X"02",X"09",X"07",X"00",X"02",X"0A",
		X"07",X"00",X"02",X"0B",X"07",X"00",X"02",X"0C",X"07",X"00",X"02",X"0D",X"07",X"00",X"02",X"0E",
		X"07",X"00",X"02",X"0F",X"07",X"00",X"02",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3A",X"2E",
		X"85",X"FE",X"14",X"38",X"02",X"3E",X"13",X"CB",X"27",X"4F",X"06",X"00",X"21",X"25",X"36",X"09",
		X"5E",X"23",X"56",X"EB",X"E9",X"4D",X"36",X"4D",X"36",X"61",X"36",X"7D",X"36",X"92",X"36",X"A8",
		X"36",X"C3",X"36",X"DC",X"36",X"F5",X"36",X"09",X"37",X"1F",X"37",X"39",X"37",X"5B",X"37",X"76",
		X"37",X"92",X"37",X"B3",X"37",X"D2",X"37",X"F1",X"37",X"0B",X"38",X"27",X"38",X"CF",X"48",X"F0",
		X"54",X"48",X"45",X"20",X"46",X"41",X"43",X"45",X"20",X"52",X"4F",X"4F",X"4D",X"00",X"DF",X"F0",
		X"C9",X"CF",X"28",X"F0",X"54",X"48",X"45",X"20",X"45",X"56",X"49",X"4C",X"20",X"45",X"59",X"45",
		X"42",X"41",X"4C",X"4C",X"20",X"52",X"4F",X"4F",X"4D",X"00",X"DF",X"F1",X"C9",X"CF",X"48",X"F0",
		X"54",X"48",X"45",X"20",X"53",X"51",X"55",X"49",X"44",X"20",X"52",X"4F",X"4F",X"4D",X"00",X"DF",
		X"F7",X"C9",X"CF",X"40",X"F0",X"54",X"48",X"45",X"20",X"53",X"49",X"43",X"4B",X"4C",X"45",X"20",
		X"52",X"4F",X"4F",X"4D",X"00",X"DF",X"F1",X"C9",X"CF",X"30",X"F0",X"54",X"48",X"45",X"20",X"43",
		X"41",X"54",X"45",X"52",X"50",X"49",X"4C",X"4C",X"41",X"52",X"20",X"52",X"4F",X"4F",X"4D",X"00",
		X"DF",X"F3",X"C9",X"CF",X"38",X"F0",X"54",X"48",X"45",X"20",X"50",X"52",X"4F",X"50",X"45",X"4C",
		X"4C",X"45",X"52",X"20",X"52",X"4F",X"4F",X"4D",X"00",X"DF",X"F7",X"C9",X"CF",X"38",X"F0",X"54",
		X"48",X"45",X"20",X"43",X"59",X"43",X"4C",X"4F",X"54",X"52",X"4F",X"4E",X"20",X"52",X"4F",X"4F",
		X"4D",X"00",X"DF",X"F3",X"C9",X"CF",X"48",X"F0",X"54",X"48",X"45",X"20",X"54",X"41",X"5A",X"5A",
		X"20",X"52",X"4F",X"4F",X"4D",X"00",X"DF",X"F1",X"C9",X"CF",X"40",X"F0",X"54",X"48",X"45",X"20",
		X"48",X"4F",X"50",X"50",X"45",X"52",X"20",X"52",X"4F",X"4F",X"4D",X"00",X"DF",X"F0",X"C9",X"CF",
		X"30",X"F0",X"54",X"48",X"45",X"20",X"53",X"55",X"50",X"45",X"52",X"20",X"46",X"41",X"43",X"45",
		X"20",X"52",X"4F",X"4F",X"4D",X"00",X"DF",X"F1",X"C9",X"CF",X"10",X"F0",X"54",X"48",X"45",X"20",
		X"45",X"56",X"49",X"4C",X"20",X"53",X"55",X"50",X"45",X"52",X"20",X"45",X"59",X"45",X"42",X"41",
		X"4C",X"4C",X"20",X"52",X"4F",X"4F",X"4D",X"00",X"DF",X"F7",X"C9",X"CF",X"30",X"F0",X"54",X"48",
		X"45",X"20",X"53",X"55",X"50",X"45",X"52",X"20",X"53",X"51",X"55",X"49",X"44",X"20",X"52",X"4F",
		X"4F",X"4D",X"00",X"DF",X"F1",X"C9",X"CF",X"28",X"F0",X"54",X"48",X"45",X"20",X"53",X"55",X"50",
		X"45",X"52",X"20",X"53",X"49",X"43",X"4B",X"4C",X"45",X"20",X"52",X"4F",X"4F",X"4D",X"00",X"DF",
		X"F3",X"C9",X"CF",X"18",X"F0",X"54",X"48",X"45",X"20",X"53",X"55",X"50",X"45",X"52",X"20",X"43",
		X"41",X"54",X"45",X"52",X"50",X"49",X"4C",X"4C",X"41",X"52",X"20",X"52",X"4F",X"4F",X"4D",X"00",
		X"DF",X"F7",X"C9",X"CF",X"20",X"F0",X"54",X"48",X"45",X"20",X"53",X"55",X"50",X"45",X"52",X"20",
		X"50",X"52",X"4F",X"50",X"45",X"4C",X"4C",X"45",X"52",X"20",X"52",X"4F",X"4F",X"4D",X"00",X"DF",
		X"F3",X"C9",X"CF",X"20",X"F0",X"54",X"48",X"45",X"20",X"53",X"55",X"50",X"45",X"52",X"20",X"43",
		X"59",X"43",X"4C",X"4F",X"54",X"52",X"4F",X"4E",X"20",X"52",X"4F",X"4F",X"4D",X"00",X"DF",X"F1",
		X"C9",X"CF",X"30",X"F0",X"54",X"48",X"45",X"20",X"53",X"55",X"50",X"45",X"52",X"20",X"54",X"41",
		X"5A",X"5A",X"20",X"52",X"4F",X"4F",X"4D",X"00",X"DF",X"F0",X"C9",X"CF",X"28",X"F0",X"54",X"48",
		X"45",X"20",X"53",X"55",X"50",X"45",X"52",X"20",X"48",X"4F",X"50",X"50",X"45",X"52",X"20",X"52",
		X"4F",X"4F",X"4D",X"00",X"DF",X"F1",X"C9",X"CF",X"30",X"F0",X"54",X"48",X"45",X"20",X"53",X"55",
		X"50",X"45",X"52",X"20",X"4D",X"49",X"58",X"45",X"44",X"20",X"52",X"4F",X"4F",X"4D",X"00",X"DF",
		X"F7",X"C9",X"00",X"00",X"01",X"00",X"00",X"06",X"06",X"02",X"3D",X"02",X"06",X"06",X"02",X"3D",
		X"02",X"06",X"06",X"02",X"3D",X"02",X"06",X"06",X"02",X"3D",X"02",X"00",X"01",X"5F",X"85",X"00",
		X"00",X"01",X"00",X"00",X"0A",X"0A",X"02",X"37",X"01",X"00",X"01",X"64",X"38",X"CD",X"0E",X"36",
		X"CD",X"D3",X"06",X"CD",X"ED",X"07",X"21",X"6F",X"3D",X"06",X"00",X"3A",X"2E",X"85",X"F5",X"4F",
		X"09",X"7E",X"32",X"2E",X"85",X"CF",X"A8",X"F8",X"4C",X"45",X"56",X"45",X"4C",X"20",X"00",X"21",
		X"F8",X"D8",X"11",X"2E",X"85",X"06",X"02",X"CD",X"27",X"05",X"F1",X"32",X"2E",X"85",X"CD",X"85",
		X"08",X"DD",X"21",X"12",X"82",X"FD",X"21",X"9A",X"81",X"21",X"2A",X"85",X"36",X"00",X"21",X"2B",
		X"85",X"36",X"00",X"CD",X"C2",X"3C",X"DD",X"CB",X"00",X"D6",X"AF",X"DD",X"77",X"0D",X"DD",X"CB",
		X"0C",X"C6",X"CD",X"DA",X"3B",X"DD",X"CB",X"00",X"F6",X"FD",X"36",X"01",X"14",X"FD",X"CB",X"00",
		X"CE",X"3E",X"01",X"32",X"44",X"86",X"CD",X"BC",X"09",X"FD",X"21",X"9A",X"81",X"3A",X"25",X"85",
		X"E6",X"08",X"20",X"0A",X"3A",X"24",X"85",X"E6",X"3C",X"28",X"03",X"C3",X"B8",X"3A",X"21",X"43",
		X"86",X"7E",X"B7",X"28",X"01",X"35",X"3A",X"59",X"85",X"FE",X"02",X"20",X"11",X"3A",X"02",X"98",
		X"E6",X"08",X"20",X"0A",X"3A",X"27",X"85",X"CB",X"77",X"C4",X"21",X"3B",X"18",X"08",X"3A",X"26",
		X"85",X"CB",X"47",X"C4",X"21",X"3B",X"DD",X"7E",X"0D",X"CB",X"57",X"C2",X"6D",X"3B",X"FD",X"CB",
		X"00",X"4E",X"20",X"1E",X"FD",X"CB",X"00",X"F6",X"3A",X"2C",X"85",X"FE",X"05",X"FD",X"36",X"01",
		X"1E",X"30",X"0B",X"FD",X"36",X"01",X"0A",X"B7",X"20",X"04",X"FD",X"36",X"01",X"05",X"FD",X"CB",
		X"00",X"CE",X"3A",X"23",X"85",X"CB",X"4F",X"C2",X"5C",X"39",X"3A",X"23",X"85",X"E6",X"3C",X"21",
		X"2B",X"85",X"46",X"77",X"A8",X"C4",X"DF",X"3C",X"DD",X"CB",X"00",X"E6",X"3A",X"32",X"85",X"E6",
		X"03",X"28",X"35",X"FE",X"01",X"28",X"22",X"FE",X"02",X"28",X"0F",X"FD",X"7E",X"0D",X"FE",X"70",
		X"DA",X"A5",X"39",X"FE",X"74",X"DA",X"6D",X"3B",X"18",X"2B",X"FD",X"7E",X"0D",X"FE",X"60",X"DA",
		X"A5",X"39",X"FE",X"64",X"DA",X"6D",X"3B",X"18",X"1C",X"FD",X"7E",X"0D",X"FE",X"88",X"DA",X"A5",
		X"39",X"FE",X"8C",X"DA",X"6D",X"3B",X"18",X"0D",X"FD",X"7E",X"0D",X"FE",X"38",X"DA",X"A5",X"39",
		X"FE",X"3C",X"DA",X"6D",X"3B",X"01",X"00",X"00",X"11",X"00",X"00",X"3A",X"23",X"85",X"CB",X"4F",
		X"C2",X"C3",X"39",X"3A",X"23",X"85",X"67",X"CD",X"7B",X"3C",X"CD",X"8C",X"3C",X"CD",X"9A",X"3C",
		X"CD",X"AC",X"3C",X"FD",X"70",X"04",X"FD",X"71",X"03",X"FD",X"72",X"0A",X"FD",X"73",X"09",X"3A",
		X"23",X"85",X"CB",X"4F",X"C4",X"D6",X"3A",X"FD",X"CB",X"00",X"56",X"28",X"3F",X"21",X"40",X"86",
		X"36",X"FD",X"FD",X"CB",X"02",X"56",X"28",X"0B",X"3E",X"FF",X"32",X"03",X"A8",X"32",X"04",X"A8",
		X"C3",X"1C",X"3A",X"3E",X"00",X"32",X"03",X"A8",X"32",X"04",X"A8",X"3E",X"01",X"CD",X"10",X"0A",
		X"CD",X"21",X"3D",X"11",X"2E",X"00",X"06",X"07",X"DD",X"E5",X"FD",X"E5",X"DD",X"21",X"6E",X"82",
		X"DD",X"CB",X"0D",X"CE",X"DD",X"19",X"10",X"F8",X"FD",X"E1",X"DD",X"E1",X"3A",X"34",X"86",X"47",
		X"DD",X"7E",X"08",X"B8",X"38",X"03",X"DD",X"70",X"08",X"3A",X"33",X"86",X"47",X"DD",X"7E",X"08",
		X"B8",X"30",X"03",X"DD",X"70",X"08",X"3A",X"3F",X"86",X"CB",X"7F",X"CA",X"53",X"3A",X"CD",X"88",
		X"19",X"3E",X"01",X"32",X"58",X"85",X"DD",X"7E",X"0A",X"FE",X"17",X"38",X"0E",X"FE",X"D7",X"38",
		X"02",X"18",X"39",X"3E",X"01",X"CD",X"10",X"0A",X"C3",X"D9",X"38",X"CD",X"88",X"19",X"01",X"00",
		X"00",X"11",X"00",X"02",X"CD",X"BE",X"0F",X"FD",X"21",X"9A",X"81",X"FD",X"70",X"04",X"FD",X"71",
		X"03",X"FD",X"72",X"0A",X"FD",X"73",X"09",X"3E",X"00",X"CB",X"D7",X"32",X"2B",X"85",X"CD",X"DF",
		X"3C",X"DD",X"CB",X"00",X"E6",X"3E",X"0B",X"CD",X"10",X"0A",X"18",X"2C",X"CD",X"88",X"19",X"01",
		X"00",X"00",X"11",X"00",X"02",X"FD",X"21",X"9A",X"81",X"FD",X"70",X"04",X"FD",X"71",X"03",X"FD",
		X"72",X"0A",X"FD",X"73",X"09",X"3E",X"00",X"CB",X"DF",X"32",X"2B",X"85",X"CD",X"DF",X"3C",X"DD",
		X"CB",X"00",X"E6",X"3E",X"10",X"CD",X"10",X"0A",X"3E",X"02",X"32",X"58",X"85",X"FD",X"21",X"9A",
		X"81",X"FD",X"36",X"03",X"00",X"FD",X"36",X"04",X"00",X"FD",X"36",X"09",X"00",X"FD",X"36",X"0A",
		X"00",X"CD",X"BC",X"09",X"18",X"FB",X"3A",X"23",X"85",X"E6",X"3C",X"C8",X"DD",X"CB",X"00",X"A6",
		X"06",X"00",X"CB",X"3F",X"CB",X"3F",X"4F",X"21",X"11",X"3B",X"09",X"7E",X"FD",X"77",X"07",X"3A",
		X"2A",X"85",X"FE",X"07",X"C8",X"D0",X"3A",X"43",X"86",X"B7",X"C0",X"3E",X"02",X"32",X"43",X"86",
		X"FD",X"21",X"DD",X"3D",X"CD",X"A4",X"09",X"FD",X"21",X"9A",X"81",X"3E",X"04",X"CD",X"1F",X"08",
		X"C9",X"00",X"3E",X"3F",X"00",X"95",X"94",X"93",X"00",X"15",X"14",X"13",X"00",X"00",X"00",X"00",
		X"00",X"CB",X"87",X"32",X"26",X"85",X"FD",X"7E",X"02",X"B7",X"C0",X"3A",X"2F",X"85",X"B7",X"C8",
		X"3D",X"32",X"2F",X"85",X"FD",X"36",X"01",X"FA",X"FD",X"CB",X"00",X"CE",X"FD",X"36",X"02",X"23",
		X"FD",X"CB",X"00",X"D6",X"11",X"2E",X"00",X"06",X"07",X"DD",X"E5",X"FD",X"E5",X"DD",X"21",X"6E",
		X"82",X"DD",X"CB",X"0D",X"CE",X"DD",X"19",X"10",X"F8",X"CD",X"ED",X"07",X"CD",X"58",X"0F",X"3E",
		X"07",X"CD",X"1F",X"08",X"FD",X"E1",X"DD",X"E1",X"DD",X"36",X"0D",X"00",X"C9",X"DD",X"CB",X"0C",
		X"86",X"3A",X"29",X"85",X"C6",X"99",X"27",X"32",X"29",X"85",X"3E",X"05",X"CD",X"1F",X"08",X"AF",
		X"FD",X"77",X"03",X"FD",X"77",X"04",X"FD",X"77",X"09",X"FD",X"77",X"0A",X"DD",X"21",X"12",X"82",
		X"DD",X"CB",X"00",X"B6",X"DD",X"CB",X"00",X"A6",X"21",X"E5",X"15",X"DD",X"75",X"05",X"DD",X"74",
		X"06",X"DD",X"36",X"04",X"01",X"DD",X"CB",X"00",X"E6",X"DD",X"CB",X"00",X"66",X"28",X"05",X"CD",
		X"BC",X"09",X"18",X"F5",X"AF",X"FD",X"77",X"03",X"FD",X"77",X"04",X"FD",X"77",X"09",X"FD",X"77",
		X"0A",X"DD",X"77",X"08",X"DD",X"77",X"0A",X"FD",X"77",X"06",X"FD",X"77",X"0C",X"3E",X"0A",X"CD",
		X"10",X"0A",X"CD",X"36",X"0A",X"CD",X"BC",X"09",X"18",X"FB",X"CF",X"50",X"78",X"50",X"4C",X"41",
		X"59",X"45",X"52",X"20",X"20",X"20",X"55",X"50",X"00",X"21",X"78",X"88",X"11",X"59",X"85",X"06",
		X"01",X"CD",X"27",X"05",X"DD",X"36",X"08",X"7A",X"DD",X"36",X"0A",X"D7",X"01",X"00",X"00",X"11",
		X"00",X"02",X"CD",X"BE",X"0F",X"FD",X"70",X"04",X"FD",X"71",X"03",X"FD",X"72",X"0A",X"FD",X"73",
		X"09",X"3A",X"2B",X"85",X"CB",X"D7",X"32",X"2B",X"85",X"CD",X"DF",X"3C",X"DD",X"CB",X"00",X"E6",
		X"FD",X"36",X"01",X"05",X"FD",X"CB",X"00",X"CE",X"3E",X"08",X"CD",X"1F",X"08",X"FD",X"CB",X"00",
		X"4E",X"28",X"0A",X"DD",X"7E",X"0A",X"FE",X"7D",X"30",X"F3",X"C3",X"57",X"3C",X"FD",X"36",X"01",
		X"05",X"FD",X"CB",X"00",X"CE",X"3E",X"09",X"CD",X"1F",X"08",X"FD",X"CB",X"00",X"4E",X"28",X"D0",
		X"DD",X"7E",X"0A",X"FE",X"7D",X"30",X"F3",X"11",X"00",X"00",X"FD",X"72",X"0A",X"FD",X"73",X"09",
		X"FD",X"36",X"07",X"3D",X"DD",X"CB",X"00",X"A6",X"CF",X"50",X"78",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"00",X"CD",X"26",X"35",X"C9",X"CB",X"54",X"C8",X"FD",X"7E",
		X"0C",X"FE",X"16",X"D8",X"ED",X"5B",X"4A",X"85",X"CD",X"BE",X"0F",X"C9",X"CB",X"5C",X"C8",X"FD",
		X"7E",X"0C",X"FE",X"D8",X"D0",X"ED",X"5B",X"4A",X"85",X"C9",X"CB",X"64",X"C8",X"FD",X"7E",X"06",
		X"E5",X"21",X"34",X"86",X"BE",X"E1",X"D0",X"ED",X"4B",X"4A",X"85",X"C9",X"CB",X"6C",X"C8",X"FD",
		X"7E",X"06",X"E5",X"21",X"33",X"86",X"BE",X"E1",X"D8",X"C8",X"ED",X"4B",X"4A",X"85",X"CD",X"C6",
		X"0F",X"C9",X"21",X"42",X"38",X"11",X"5A",X"85",X"01",X"1E",X"00",X"ED",X"B0",X"21",X"5A",X"85",
		X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",X"36",X"04",X"01",X"DD",X"CB",X"00",X"E6",X"C9",X"21",
		X"2F",X"3D",X"06",X"00",X"3A",X"2B",X"85",X"CB",X"3F",X"CB",X"3F",X"4F",X"09",X"09",X"09",X"09",
		X"7E",X"B7",X"C8",X"DD",X"CB",X"00",X"A6",X"DD",X"E5",X"DD",X"21",X"5A",X"85",X"11",X"05",X"00",
		X"DD",X"19",X"DD",X"77",X"03",X"DD",X"19",X"23",X"7E",X"DD",X"77",X"03",X"DD",X"19",X"23",X"7E",
		X"DD",X"77",X"03",X"DD",X"19",X"23",X"7E",X"DD",X"77",X"03",X"DD",X"E1",X"DD",X"36",X"04",X"01",
		X"C9",X"21",X"05",X"90",X"06",X"1C",X"3A",X"48",X"86",X"77",X"23",X"23",X"10",X"FB",X"C9",X"3D",
		X"3D",X"3D",X"3D",X"3B",X"3A",X"BB",X"BA",X"3D",X"3C",X"BD",X"BC",X"00",X"00",X"00",X"00",X"B9",
		X"B8",X"B6",X"B7",X"B9",X"B8",X"B6",X"B7",X"B9",X"B8",X"B6",X"B7",X"00",X"00",X"00",X"00",X"39",
		X"38",X"36",X"37",X"39",X"38",X"36",X"37",X"39",X"38",X"36",X"37",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"02",X"03",X"04",X"05",X"06",X"07",X"08",X"09",X"10",X"11",X"12",X"13",X"14",X"15",X"16",
		X"17",X"18",X"19",X"20",X"21",X"22",X"23",X"24",X"25",X"26",X"27",X"28",X"29",X"30",X"31",X"32",
		X"33",X"34",X"35",X"36",X"37",X"38",X"39",X"40",X"41",X"42",X"43",X"44",X"45",X"46",X"47",X"48",
		X"49",X"50",X"51",X"52",X"53",X"54",X"55",X"56",X"57",X"58",X"59",X"60",X"61",X"62",X"63",X"64",
		X"65",X"66",X"67",X"68",X"69",X"70",X"71",X"72",X"73",X"74",X"75",X"76",X"77",X"78",X"79",X"80",
		X"81",X"82",X"83",X"84",X"85",X"86",X"87",X"88",X"89",X"90",X"91",X"92",X"93",X"94",X"95",X"96",
		X"97",X"98",X"99",X"00",X"00",X"01",X"00",X"00",X"04",X"04",X"00",X"00",X"00",X"CD",X"F0",X"08",
		X"D2",X"3A",X"3E",X"DD",X"E5",X"FD",X"E1",X"DD",X"2A",X"DA",X"80",X"21",X"2A",X"85",X"34",X"CD",
		X"C2",X"3E",X"CD",X"F0",X"3E",X"DD",X"CB",X"0C",X"F6",X"21",X"D3",X"3D",X"DD",X"75",X"05",X"DD",
		X"74",X"06",X"3E",X"0C",X"DD",X"77",X"03",X"DD",X"CB",X"00",X"EE",X"DD",X"CB",X"00",X"D6",X"DD",
		X"CB",X"00",X"F6",X"FD",X"E5",X"CD",X"BC",X"09",X"FD",X"E1",X"CD",X"46",X"3E",X"CD",X"61",X"3E",
		X"CD",X"9F",X"3E",X"CD",X"7C",X"3E",X"DD",X"7E",X"0D",X"CB",X"57",X"20",X"0D",X"DD",X"CB",X"00",
		X"6E",X"28",X"07",X"FD",X"E5",X"CD",X"BC",X"09",X"18",X"DE",X"21",X"2A",X"85",X"35",X"CD",X"36",
		X"0A",X"CD",X"BC",X"09",X"18",X"FB",X"DD",X"7E",X"0A",X"FE",X"14",X"D0",X"FD",X"46",X"0A",X"FD",
		X"4E",X"09",X"CD",X"C6",X"0F",X"FD",X"70",X"0A",X"FD",X"71",X"09",X"3E",X"16",X"DD",X"77",X"0A",
		X"C9",X"DD",X"7E",X"0A",X"FE",X"DA",X"D8",X"FD",X"46",X"0A",X"FD",X"4E",X"09",X"CD",X"C6",X"0F",
		X"FD",X"70",X"0A",X"FD",X"71",X"09",X"3E",X"D8",X"DD",X"77",X"0A",X"C9",X"3A",X"34",X"86",X"47",
		X"DD",X"7E",X"08",X"04",X"04",X"B8",X"D8",X"FD",X"46",X"04",X"FD",X"4E",X"03",X"CD",X"C6",X"0F",
		X"FD",X"70",X"04",X"FD",X"71",X"03",X"3A",X"34",X"86",X"3D",X"3D",X"DD",X"77",X"08",X"C9",X"3A",
		X"33",X"86",X"47",X"DD",X"7E",X"08",X"05",X"05",X"B8",X"D0",X"FD",X"46",X"04",X"FD",X"4E",X"03",
		X"CD",X"C6",X"0F",X"FD",X"70",X"04",X"FD",X"71",X"03",X"3A",X"33",X"86",X"3C",X"3C",X"DD",X"77",
		X"08",X"C9",X"FD",X"E5",X"FD",X"21",X"12",X"82",X"FD",X"46",X"08",X"05",X"05",X"CD",X"42",X"08",
		X"E6",X"07",X"FE",X"06",X"30",X"F7",X"80",X"DD",X"77",X"08",X"FD",X"46",X"0A",X"05",X"05",X"05",
		X"CD",X"42",X"08",X"E6",X"07",X"FE",X"06",X"30",X"F7",X"80",X"DD",X"77",X"0A",X"FD",X"E1",X"C9",
		X"3A",X"55",X"85",X"B7",X"3A",X"36",X"86",X"20",X"03",X"3A",X"23",X"85",X"E6",X"3C",X"C8",X"CB",
		X"3F",X"CB",X"3F",X"5F",X"16",X"00",X"21",X"21",X"3F",X"19",X"19",X"19",X"19",X"5E",X"23",X"56",
		X"23",X"4E",X"23",X"46",X"FD",X"73",X"03",X"FD",X"72",X"04",X"FD",X"71",X"09",X"FD",X"70",X"0A",
		X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"F8",X"00",X"00",X"F0",X"07",X"00",X"00",X"00",
		X"00",X"F0",X"07",X"00",X"00",X"60",X"06",X"A0",X"F9",X"60",X"06",X"60",X"06",X"00",X"00",X"00",
		X"00",X"10",X"F8",X"00",X"00",X"A0",X"F9",X"A0",X"F9",X"A0",X"F9",X"60",X"06",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"CD",X"69",X"0A",X"CD",X"82",X"05",X"21",X"2E",X"85",X"34",X"3E",X"00",X"32",X"58",X"85",
		X"3A",X"2E",X"85",X"E6",X"0F",X"FE",X"03",X"28",X"12",X"FE",X"06",X"28",X"0E",X"FE",X"09",X"28",
		X"0A",X"FE",X"0C",X"28",X"06",X"FE",X"0F",X"28",X"02",X"18",X"12",X"FD",X"21",X"9A",X"2A",X"CD",
		X"A4",X"09",X"21",X"32",X"85",X"7E",X"3C",X"E6",X"03",X"77",X"C3",X"7D",X"41",X"D7",X"00",X"3E",
		X"05",X"CD",X"10",X"0A",X"CD",X"82",X"05",X"CD",X"89",X"06",X"CD",X"D3",X"06",X"CD",X"ED",X"07",
		X"21",X"6F",X"3D",X"06",X"00",X"3A",X"2E",X"85",X"F5",X"4F",X"09",X"7E",X"32",X"2E",X"85",X"CF",
		X"A8",X"F8",X"4C",X"45",X"56",X"45",X"4C",X"20",X"00",X"21",X"F8",X"D8",X"11",X"2E",X"85",X"06",
		X"02",X"CD",X"27",X"05",X"F1",X"32",X"2E",X"85",X"CF",X"20",X"48",X"43",X"4F",X"4E",X"47",X"52",
		X"41",X"54",X"55",X"4C",X"41",X"54",X"49",X"4F",X"4E",X"53",X"20",X"59",X"4F",X"55",X"20",X"48",
		X"41",X"56",X"45",X"00",X"CF",X"30",X"60",X"43",X"4C",X"45",X"41",X"52",X"45",X"44",X"20",X"41",
		X"4E",X"4F",X"54",X"48",X"45",X"52",X"20",X"52",X"4F",X"4F",X"4D",X"00",X"CF",X"20",X"90",X"53",
		X"4F",X"20",X"50",X"52",X"45",X"50",X"41",X"52",X"45",X"20",X"59",X"4F",X"55",X"52",X"53",X"45",
		X"4C",X"46",X"20",X"46",X"4F",X"52",X"00",X"E7",X"12",X"05",X"02",X"CD",X"A2",X"41",X"FD",X"21",
		X"E4",X"40",X"CD",X"A4",X"09",X"FD",X"21",X"48",X"40",X"CD",X"A4",X"09",X"CD",X"BC",X"09",X"3A",
		X"12",X"82",X"B7",X"CA",X"7D",X"41",X"18",X"F4",X"CD",X"85",X"08",X"DD",X"21",X"12",X"82",X"FD",
		X"21",X"9A",X"81",X"CD",X"C2",X"3C",X"DD",X"CB",X"00",X"D6",X"DD",X"CB",X"0C",X"C6",X"DD",X"36",
		X"08",X"7A",X"DD",X"36",X"0A",X"00",X"01",X"00",X"00",X"11",X"00",X"03",X"1E",X"00",X"FD",X"70",
		X"04",X"FD",X"71",X"03",X"FD",X"72",X"0A",X"FD",X"73",X"09",X"3E",X"00",X"CB",X"DF",X"32",X"2B",
		X"85",X"CD",X"DF",X"3C",X"DD",X"CB",X"00",X"E6",X"FD",X"36",X"01",X"0A",X"FD",X"CB",X"00",X"CE",
		X"FD",X"36",X"02",X"05",X"FD",X"CB",X"00",X"D6",X"FD",X"CB",X"00",X"4E",X"20",X"0D",X"3E",X"08",
		X"CD",X"1F",X"08",X"FD",X"36",X"01",X"0A",X"FD",X"CB",X"00",X"CE",X"FD",X"CB",X"00",X"56",X"20",
		X"0D",X"3E",X"09",X"CD",X"1F",X"08",X"FD",X"36",X"02",X"0A",X"FD",X"CB",X"00",X"D6",X"DD",X"7E",
		X"0A",X"FE",X"FD",X"30",X"09",X"FD",X"E5",X"CD",X"BC",X"09",X"FD",X"E1",X"18",X"CA",X"11",X"00",
		X"00",X"FD",X"72",X"0A",X"FD",X"73",X"09",X"3E",X"14",X"CD",X"10",X"0A",X"CD",X"36",X"0A",X"CD",
		X"BC",X"09",X"18",X"FB",X"CD",X"26",X"09",X"D2",X"CE",X"40",X"CD",X"CE",X"08",X"D2",X"CE",X"40",
		X"FD",X"2A",X"DA",X"80",X"FD",X"E5",X"3E",X"04",X"CD",X"10",X"0A",X"FD",X"E1",X"FD",X"66",X"02",
		X"FD",X"6E",X"01",X"E5",X"DD",X"E1",X"FD",X"36",X"08",X"7A",X"FD",X"36",X"0A",X"00",X"01",X"00",
		X"00",X"11",X"00",X"02",X"DD",X"70",X"04",X"DD",X"71",X"03",X"DD",X"72",X"0A",X"DD",X"73",X"09",
		X"CD",X"4E",X"41",X"FD",X"CB",X"0C",X"D6",X"FD",X"CB",X"00",X"D6",X"FD",X"36",X"0D",X"00",X"DD",
		X"E5",X"CD",X"BC",X"09",X"FD",X"E1",X"FD",X"7E",X"07",X"FE",X"35",X"20",X"06",X"DD",X"CB",X"00",
		X"96",X"18",X"04",X"DD",X"CB",X"00",X"D6",X"FD",X"E5",X"CD",X"BC",X"09",X"18",X"E6",X"21",X"60",
		X"41",X"FD",X"75",X"05",X"FD",X"74",X"06",X"FD",X"36",X"04",X"01",X"FD",X"CB",X"00",X"E6",X"C9",
		X"00",X"00",X"01",X"00",X"00",X"0C",X"0C",X"05",X"35",X"06",X"0C",X"0C",X"04",X"33",X"06",X"0C",
		X"0C",X"05",X"34",X"06",X"0C",X"0C",X"04",X"33",X"06",X"00",X"01",X"65",X"41",X"CD",X"69",X"0A",
		X"3A",X"2D",X"85",X"C6",X"0A",X"FE",X"F5",X"38",X"02",X"3E",X"F5",X"32",X"2D",X"85",X"32",X"2C",
		X"85",X"CD",X"82",X"05",X"DD",X"21",X"12",X"82",X"DD",X"CB",X"0B",X"7E",X"C2",X"6B",X"2F",X"C3",
		X"47",X"2F",X"3A",X"2E",X"85",X"FE",X"14",X"38",X"02",X"3E",X"13",X"CB",X"27",X"4F",X"06",X"00",
		X"21",X"B9",X"41",X"09",X"5E",X"23",X"56",X"EB",X"E9",X"E1",X"41",X"E1",X"41",X"F5",X"41",X"11",
		X"42",X"26",X"42",X"3C",X"42",X"57",X"42",X"70",X"42",X"89",X"42",X"9D",X"42",X"B3",X"42",X"CD",
		X"42",X"EF",X"42",X"0A",X"43",X"26",X"43",X"47",X"43",X"66",X"43",X"85",X"43",X"9F",X"43",X"BB",
		X"43",X"CF",X"48",X"A8",X"54",X"48",X"45",X"20",X"46",X"41",X"43",X"45",X"20",X"52",X"4F",X"4F",
		X"4D",X"00",X"DF",X"AD",X"C9",X"CF",X"28",X"A8",X"54",X"48",X"45",X"20",X"45",X"56",X"49",X"4C",
		X"20",X"45",X"59",X"45",X"42",X"41",X"4C",X"4C",X"20",X"52",X"4F",X"4F",X"4D",X"00",X"DF",X"AD",
		X"C9",X"CF",X"48",X"A8",X"54",X"48",X"45",X"20",X"53",X"51",X"55",X"49",X"44",X"20",X"52",X"4F",
		X"4F",X"4D",X"00",X"DF",X"AD",X"C9",X"CF",X"40",X"A8",X"54",X"48",X"45",X"20",X"53",X"49",X"43",
		X"4B",X"4C",X"45",X"20",X"52",X"4F",X"4F",X"4D",X"00",X"DF",X"AD",X"C9",X"CF",X"30",X"A8",X"54",
		X"48",X"45",X"20",X"43",X"41",X"54",X"45",X"52",X"50",X"49",X"4C",X"4C",X"41",X"52",X"20",X"52",
		X"4F",X"4F",X"4D",X"00",X"DF",X"AD",X"C9",X"CF",X"38",X"A8",X"54",X"48",X"45",X"20",X"50",X"52",
		X"4F",X"50",X"45",X"4C",X"4C",X"45",X"52",X"20",X"52",X"4F",X"4F",X"4D",X"00",X"DF",X"AD",X"C9",
		X"CF",X"38",X"A8",X"54",X"48",X"45",X"20",X"43",X"59",X"43",X"4C",X"4F",X"54",X"52",X"4F",X"4E",
		X"20",X"52",X"4F",X"4F",X"4D",X"00",X"DF",X"AD",X"C9",X"CF",X"48",X"A8",X"54",X"48",X"45",X"20",
		X"54",X"41",X"5A",X"5A",X"20",X"52",X"4F",X"4F",X"4D",X"00",X"DF",X"AD",X"C9",X"CF",X"40",X"A8",
		X"54",X"48",X"45",X"20",X"48",X"4F",X"50",X"50",X"45",X"52",X"20",X"52",X"4F",X"4F",X"4D",X"00",
		X"DF",X"AD",X"C9",X"CF",X"30",X"A8",X"54",X"48",X"45",X"20",X"53",X"55",X"50",X"45",X"52",X"20",
		X"46",X"41",X"43",X"45",X"20",X"52",X"4F",X"4F",X"4D",X"00",X"DF",X"AD",X"C9",X"CF",X"10",X"A8",
		X"54",X"48",X"45",X"20",X"53",X"55",X"50",X"45",X"52",X"20",X"45",X"56",X"49",X"4C",X"20",X"45",
		X"59",X"45",X"42",X"41",X"4C",X"4C",X"20",X"52",X"4F",X"4F",X"4D",X"00",X"DF",X"AD",X"C9",X"CF",
		X"30",X"A8",X"54",X"48",X"45",X"20",X"53",X"55",X"50",X"45",X"52",X"20",X"53",X"51",X"55",X"49",
		X"44",X"20",X"52",X"4F",X"4F",X"4D",X"00",X"DF",X"AD",X"C9",X"CF",X"28",X"A8",X"54",X"48",X"45",
		X"20",X"53",X"55",X"50",X"45",X"52",X"20",X"53",X"49",X"43",X"4B",X"4C",X"45",X"20",X"52",X"4F",
		X"4F",X"4D",X"00",X"DF",X"AD",X"C9",X"CF",X"18",X"A8",X"54",X"48",X"45",X"20",X"53",X"55",X"50",
		X"45",X"52",X"20",X"43",X"41",X"54",X"45",X"52",X"50",X"49",X"4C",X"4C",X"41",X"52",X"20",X"52",
		X"4F",X"4F",X"4D",X"00",X"DF",X"AD",X"C9",X"CF",X"20",X"A8",X"54",X"48",X"45",X"20",X"53",X"55",
		X"50",X"45",X"52",X"20",X"50",X"52",X"4F",X"50",X"45",X"4C",X"4C",X"45",X"52",X"20",X"52",X"4F",
		X"4F",X"4D",X"00",X"DF",X"AD",X"C9",X"CF",X"20",X"A8",X"54",X"48",X"45",X"20",X"53",X"55",X"50",
		X"45",X"52",X"20",X"43",X"59",X"43",X"4C",X"4F",X"54",X"52",X"4F",X"4E",X"20",X"52",X"4F",X"4F",
		X"4D",X"00",X"DF",X"AD",X"C9",X"CF",X"30",X"A8",X"54",X"48",X"45",X"20",X"53",X"55",X"50",X"45",
		X"52",X"20",X"54",X"41",X"5A",X"5A",X"20",X"52",X"4F",X"4F",X"4D",X"00",X"DF",X"AD",X"C9",X"CF",
		X"28",X"A8",X"54",X"48",X"45",X"20",X"53",X"55",X"50",X"45",X"52",X"20",X"48",X"4F",X"50",X"50",
		X"45",X"52",X"20",X"52",X"4F",X"4F",X"4D",X"00",X"DF",X"AD",X"C9",X"CF",X"30",X"A8",X"54",X"48",
		X"45",X"20",X"53",X"55",X"50",X"45",X"52",X"20",X"4D",X"49",X"58",X"45",X"44",X"20",X"52",X"4F",
		X"4F",X"4D",X"00",X"DF",X"AD",X"C9",X"3E",X"FF",X"32",X"55",X"85",X"CD",X"5F",X"22",X"CD",X"85",
		X"08",X"3E",X"14",X"32",X"33",X"86",X"3E",X"FA",X"32",X"34",X"86",X"3E",X"00",X"32",X"36",X"86",
		X"32",X"37",X"86",X"DD",X"21",X"12",X"82",X"DD",X"CB",X"00",X"F6",X"DD",X"21",X"12",X"82",X"FD",
		X"21",X"9A",X"81",X"21",X"2A",X"85",X"36",X"00",X"21",X"2B",X"85",X"36",X"00",X"CD",X"C2",X"3C",
		X"DD",X"CB",X"00",X"D6",X"AF",X"DD",X"77",X"0D",X"DD",X"CB",X"0C",X"C6",X"DD",X"36",X"08",X"0A",
		X"DD",X"36",X"0A",X"52",X"DD",X"CB",X"00",X"F6",X"3E",X"05",X"32",X"78",X"85",X"21",X"D4",X"44",
		X"E5",X"FD",X"21",X"9A",X"81",X"3A",X"36",X"86",X"CB",X"4F",X"C2",X"4F",X"44",X"3A",X"36",X"86",
		X"E6",X"3C",X"21",X"2B",X"85",X"46",X"77",X"A8",X"C4",X"DF",X"3C",X"DD",X"CB",X"00",X"E6",X"01",
		X"00",X"00",X"11",X"00",X"00",X"3A",X"36",X"86",X"CB",X"4F",X"C2",X"6D",X"44",X"3A",X"36",X"86",
		X"67",X"CD",X"8B",X"45",X"CD",X"95",X"45",X"CD",X"9C",X"45",X"CD",X"A3",X"45",X"FD",X"70",X"04",
		X"FD",X"71",X"03",X"FD",X"72",X"0A",X"FD",X"73",X"09",X"3A",X"36",X"86",X"CB",X"4F",X"C4",X"3D",
		X"45",X"FD",X"CB",X"00",X"4E",X"C2",X"A1",X"44",X"E1",X"7E",X"B7",X"CA",X"C6",X"44",X"FD",X"77",
		X"01",X"FD",X"CB",X"00",X"CE",X"23",X"7E",X"32",X"36",X"86",X"23",X"7E",X"32",X"37",X"86",X"23",
		X"E5",X"CD",X"89",X"2D",X"FD",X"CB",X"00",X"56",X"C2",X"B9",X"44",X"3E",X"03",X"FD",X"77",X"02",
		X"FD",X"CB",X"00",X"D6",X"3E",X"FF",X"32",X"40",X"86",X"CD",X"BC",X"09",X"3A",X"54",X"85",X"B7",
		X"C4",X"4F",X"06",X"C3",X"31",X"44",X"DD",X"CB",X"0B",X"C6",X"3E",X"00",X"32",X"55",X"85",X"CD",
		X"BC",X"09",X"18",X"FB",X"11",X"10",X"00",X"16",X"16",X"00",X"16",X"06",X"00",X"16",X"0A",X"00",
		X"16",X"0A",X"00",X"16",X"2A",X"00",X"11",X"10",X"00",X"16",X"16",X"00",X"16",X"0A",X"00",X"16",
		X"2A",X"00",X"16",X"06",X"00",X"16",X"1A",X"00",X"11",X"10",X"00",X"16",X"06",X"00",X"16",X"16",
		X"00",X"16",X"0A",X"00",X"16",X"1A",X"00",X"16",X"26",X"00",X"16",X"2A",X"00",X"10",X"10",X"00",
		X"16",X"06",X"00",X"16",X"1A",X"00",X"16",X"26",X"00",X"16",X"0A",X"00",X"16",X"2A",X"00",X"16",
		X"16",X"00",X"11",X"10",X"00",X"16",X"16",X"00",X"16",X"06",X"00",X"16",X"26",X"00",X"16",X"1A",
		X"00",X"16",X"0A",X"00",X"16",X"2A",X"00",X"1F",X"10",X"00",X"00",X"00",X"00",X"3A",X"36",X"86",
		X"E6",X"3C",X"C8",X"DD",X"CB",X"00",X"A6",X"06",X"00",X"CB",X"3F",X"CB",X"3F",X"4F",X"21",X"7B",
		X"45",X"09",X"7E",X"FD",X"77",X"07",X"3A",X"2A",X"85",X"FE",X"07",X"C8",X"D0",X"DD",X"CB",X"00",
		X"6E",X"C0",X"DD",X"36",X"03",X"02",X"DD",X"CB",X"00",X"EE",X"FD",X"21",X"DD",X"3D",X"CD",X"A4",
		X"09",X"FD",X"21",X"9A",X"81",X"3E",X"04",X"CD",X"1F",X"08",X"C9",X"00",X"3E",X"3F",X"00",X"95",
		X"94",X"93",X"00",X"15",X"14",X"13",X"00",X"00",X"00",X"00",X"00",X"CB",X"54",X"C8",X"11",X"00",
		X"02",X"CD",X"BE",X"0F",X"C9",X"CB",X"5C",X"C8",X"11",X"00",X"02",X"C9",X"CB",X"64",X"C8",X"01",
		X"00",X"02",X"C9",X"CB",X"6C",X"C8",X"01",X"00",X"02",X"CD",X"C6",X"0F",X"C9",X"18",X"CD",X"26",
		X"09",X"D2",X"E0",X"09",X"CD",X"CE",X"08",X"D2",X"05",X"47",X"FD",X"2A",X"DA",X"80",X"FD",X"66",
		X"02",X"FD",X"6E",X"01",X"E5",X"DD",X"E1",X"CD",X"07",X"17",X"21",X"00",X"00",X"DD",X"75",X"03",
		X"DD",X"74",X"04",X"DD",X"75",X"09",X"DD",X"74",X"0A",X"CD",X"0D",X"47",X"FD",X"CB",X"00",X"F6",
		X"FD",X"CB",X"0C",X"D6",X"DD",X"CB",X"00",X"EE",X"FD",X"CB",X"00",X"D6",X"FD",X"36",X"0D",X"00",
		X"3E",X"0A",X"CD",X"1F",X"08",X"DD",X"E5",X"CD",X"BC",X"09",X"FD",X"E1",X"DD",X"7E",X"0D",X"B7",
		X"C2",X"F4",X"46",X"FD",X"CB",X"00",X"4E",X"20",X"08",X"3A",X"23",X"85",X"CB",X"4F",X"C4",X"1B",
		X"46",X"CD",X"7B",X"16",X"FD",X"E5",X"CD",X"BC",X"09",X"18",X"DF",X"FD",X"36",X"01",X"0A",X"FD",
		X"CB",X"00",X"CE",X"CD",X"06",X"19",X"CD",X"E8",X"46",X"FE",X"01",X"20",X"12",X"21",X"C0",X"02",
		X"FD",X"75",X"03",X"FD",X"74",X"04",X"FD",X"36",X"09",X"00",X"FD",X"36",X"0A",X"00",X"C9",X"FE",
		X"03",X"20",X"13",X"21",X"C0",X"02",X"FD",X"75",X"03",X"FD",X"74",X"04",X"21",X"40",X"FD",X"FD",
		X"75",X"09",X"FD",X"74",X"0A",X"C9",X"FE",X"02",X"20",X"12",X"21",X"40",X"FD",X"FD",X"36",X"03",
		X"00",X"FD",X"36",X"04",X"00",X"FD",X"75",X"09",X"FD",X"74",X"0A",X"C9",X"FE",X"06",X"20",X"10",
		X"21",X"40",X"FD",X"FD",X"75",X"03",X"FD",X"74",X"04",X"FD",X"75",X"09",X"FD",X"74",X"0A",X"C9",
		X"FE",X"04",X"20",X"12",X"21",X"40",X"FD",X"FD",X"75",X"03",X"FD",X"74",X"04",X"FD",X"36",X"09",
		X"00",X"FD",X"36",X"0A",X"00",X"C9",X"FE",X"0C",X"20",X"13",X"21",X"40",X"FD",X"FD",X"75",X"03",
		X"FD",X"74",X"04",X"21",X"C0",X"02",X"FD",X"75",X"09",X"FD",X"74",X"0A",X"C9",X"FE",X"08",X"20",
		X"12",X"FD",X"36",X"03",X"00",X"FD",X"36",X"04",X"00",X"21",X"C0",X"02",X"FD",X"75",X"09",X"FD",
		X"74",X"0A",X"C9",X"FE",X"09",X"20",X"10",X"21",X"C0",X"02",X"FD",X"75",X"03",X"FD",X"74",X"04",
		X"FD",X"75",X"09",X"FD",X"74",X"0A",X"C9",X"FD",X"36",X"03",X"00",X"FD",X"36",X"04",X"00",X"FD",
		X"36",X"09",X"00",X"FD",X"36",X"0A",X"00",X"C9",X"CD",X"42",X"08",X"FE",X"64",X"38",X"02",X"78",
		X"C9",X"E6",X"0F",X"C9",X"3E",X"05",X"CD",X"1F",X"08",X"01",X"06",X"01",X"CD",X"57",X"1F",X"CD",
		X"01",X"15",X"C3",X"BA",X"45",X"CD",X"36",X"0A",X"CD",X"BC",X"09",X"18",X"FB",X"21",X"1F",X"47",
		X"FD",X"75",X"05",X"FD",X"74",X"06",X"FD",X"36",X"04",X"01",X"FD",X"CB",X"00",X"E6",X"C9",X"00",
		X"00",X"01",X"00",X"00",X"0C",X"0C",X"03",X"11",X"00",X"0C",X"0C",X"03",X"91",X"01",X"0C",X"0C",
		X"03",X"D1",X"02",X"0C",X"0C",X"03",X"51",X"03",X"0C",X"0C",X"03",X"11",X"04",X"0C",X"0C",X"03",
		X"91",X"05",X"0C",X"0C",X"03",X"D1",X"06",X"0C",X"0C",X"03",X"51",X"07",X"00",X"01",X"24",X"47",
		X"CD",X"26",X"09",X"D2",X"E0",X"09",X"CD",X"CE",X"08",X"D2",X"B3",X"48",X"FD",X"2A",X"DA",X"80",
		X"FD",X"66",X"02",X"FD",X"6E",X"01",X"E5",X"DD",X"E1",X"CD",X"07",X"17",X"21",X"00",X"00",X"DD",
		X"75",X"03",X"DD",X"74",X"04",X"DD",X"75",X"09",X"DD",X"74",X"0A",X"CD",X"BB",X"48",X"FD",X"CB",
		X"00",X"F6",X"FD",X"CB",X"0C",X"D6",X"DD",X"CB",X"00",X"EE",X"FD",X"CB",X"00",X"D6",X"FD",X"36",
		X"0D",X"00",X"3E",X"0A",X"CD",X"1F",X"08",X"DD",X"E5",X"CD",X"BC",X"09",X"FD",X"E1",X"DD",X"7E",
		X"0D",X"B7",X"C2",X"A2",X"48",X"3A",X"59",X"85",X"FE",X"02",X"20",X"0C",X"3A",X"02",X"98",X"E6",
		X"08",X"20",X"05",X"3A",X"27",X"85",X"18",X"03",X"3A",X"26",X"85",X"E6",X"3C",X"28",X"08",X"3A",
		X"23",X"85",X"CB",X"4F",X"CC",X"D1",X"47",X"CD",X"7B",X"16",X"FD",X"E5",X"CD",X"BC",X"09",X"18",
		X"CB",X"CD",X"06",X"19",X"CD",X"96",X"48",X"FE",X"01",X"20",X"12",X"21",X"C0",X"02",X"FD",X"75",
		X"03",X"FD",X"74",X"04",X"FD",X"36",X"09",X"00",X"FD",X"36",X"0A",X"00",X"C9",X"FE",X"03",X"20",
		X"13",X"21",X"C0",X"02",X"FD",X"75",X"03",X"FD",X"74",X"04",X"21",X"40",X"FD",X"FD",X"75",X"09",
		X"FD",X"74",X"0A",X"C9",X"FE",X"02",X"20",X"12",X"FD",X"36",X"03",X"00",X"FD",X"36",X"04",X"00",
		X"21",X"40",X"FD",X"FD",X"75",X"09",X"FD",X"74",X"0A",X"C9",X"FE",X"06",X"20",X"10",X"21",X"40",
		X"FD",X"FD",X"75",X"03",X"FD",X"74",X"04",X"FD",X"75",X"09",X"FD",X"74",X"0A",X"C9",X"FE",X"04",
		X"20",X"12",X"21",X"40",X"FD",X"FD",X"75",X"03",X"FD",X"74",X"04",X"FD",X"36",X"09",X"00",X"FD",
		X"36",X"0A",X"00",X"C9",X"FE",X"0C",X"20",X"13",X"21",X"40",X"FD",X"FD",X"75",X"03",X"FD",X"74",
		X"04",X"21",X"C0",X"02",X"FD",X"75",X"09",X"FD",X"74",X"0A",X"C9",X"FE",X"08",X"20",X"12",X"FD",
		X"36",X"03",X"00",X"FD",X"36",X"04",X"00",X"21",X"C0",X"02",X"FD",X"75",X"09",X"FD",X"74",X"0A",
		X"C9",X"FE",X"09",X"20",X"10",X"21",X"C0",X"02",X"FD",X"75",X"03",X"FD",X"74",X"04",X"FD",X"75",
		X"09",X"FD",X"74",X"0A",X"C9",X"FD",X"36",X"03",X"00",X"FD",X"36",X"04",X"00",X"FD",X"36",X"09",
		X"00",X"FD",X"36",X"0A",X"00",X"C9",X"CD",X"42",X"08",X"FE",X"4B",X"38",X"02",X"78",X"C9",X"E6",
		X"0F",X"C9",X"3E",X"05",X"CD",X"1F",X"08",X"01",X"06",X"01",X"CD",X"57",X"1F",X"CD",X"01",X"15",
		X"C3",X"5C",X"47",X"CD",X"36",X"0A",X"CD",X"BC",X"09",X"18",X"FB",X"21",X"CD",X"48",X"FD",X"75",
		X"05",X"FD",X"74",X"06",X"FD",X"36",X"04",X"01",X"FD",X"CB",X"00",X"E6",X"C9",X"00",X"00",X"01",
		X"00",X"00",X"0C",X"0C",X"03",X"03",X"03",X"0C",X"0C",X"03",X"83",X"03",X"0C",X"0C",X"03",X"C3",
		X"03",X"0C",X"0C",X"03",X"43",X"03",X"00",X"01",X"D2",X"48",X"CD",X"26",X"09",X"D2",X"E0",X"09",
		X"CD",X"CE",X"08",X"D2",X"0A",X"4A",X"FD",X"2A",X"DA",X"80",X"FD",X"66",X"02",X"FD",X"6E",X"01",
		X"E5",X"DD",X"E1",X"CD",X"12",X"4A",X"FD",X"36",X"0D",X"00",X"FD",X"CB",X"00",X"F6",X"FD",X"CB",
		X"0C",X"D6",X"DD",X"CB",X"00",X"EE",X"FD",X"CB",X"00",X"D6",X"FD",X"36",X"0B",X"00",X"3E",X"0A",
		X"CD",X"1F",X"08",X"DD",X"E5",X"CD",X"BC",X"09",X"FD",X"E1",X"DD",X"7E",X"0B",X"FE",X"06",X"38",
		X"03",X"C3",X"47",X"4B",X"DD",X"7E",X"0D",X"B7",X"C2",X"F9",X"49",X"CD",X"46",X"49",X"FD",X"E5",
		X"CD",X"BC",X"09",X"C3",X"28",X"49",X"DD",X"7E",X"0A",X"FE",X"16",X"30",X"1F",X"11",X"80",X"FB",
		X"FD",X"72",X"04",X"FD",X"73",X"03",X"FD",X"36",X"0A",X"00",X"FD",X"36",X"09",X"00",X"3E",X"16",
		X"DD",X"77",X"0A",X"DD",X"34",X"0B",X"21",X"70",X"4C",X"C3",X"E6",X"49",X"DD",X"7E",X"08",X"21",
		X"34",X"86",X"BE",X"38",X"20",X"11",X"80",X"FB",X"FD",X"72",X"0A",X"FD",X"73",X"09",X"FD",X"36",
		X"04",X"00",X"FD",X"36",X"03",X"00",X"7E",X"3D",X"3D",X"DD",X"77",X"08",X"DD",X"34",X"0B",X"21",
		X"96",X"4C",X"C3",X"E6",X"49",X"DD",X"7E",X"0A",X"FE",X"D9",X"38",X"1F",X"11",X"80",X"04",X"FD",
		X"72",X"04",X"FD",X"73",X"03",X"FD",X"36",X"0A",X"00",X"FD",X"36",X"09",X"00",X"3E",X"D8",X"DD",
		X"77",X"0A",X"DD",X"34",X"0B",X"21",X"83",X"4C",X"C3",X"E6",X"49",X"DD",X"7E",X"08",X"21",X"33",
		X"86",X"BE",X"30",X"21",X"11",X"80",X"04",X"FD",X"72",X"0A",X"FD",X"73",X"09",X"FD",X"36",X"04",
		X"00",X"FD",X"36",X"03",X"00",X"7E",X"3C",X"3C",X"3C",X"DD",X"77",X"08",X"DD",X"34",X"0B",X"21",
		X"A9",X"4C",X"C3",X"E6",X"49",X"C9",X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",X"36",X"04",X"01",
		X"FD",X"CB",X"00",X"96",X"DD",X"CB",X"00",X"E6",X"C9",X"3E",X"05",X"CD",X"1F",X"08",X"01",X"05",
		X"01",X"CD",X"57",X"1F",X"CD",X"01",X"15",X"C3",X"F6",X"48",X"CD",X"36",X"0A",X"CD",X"BC",X"09",
		X"18",X"FB",X"CD",X"42",X"08",X"E6",X"03",X"28",X"0C",X"FE",X"01",X"28",X"4F",X"FE",X"02",X"CA",
		X"B4",X"4A",X"C3",X"FF",X"4A",X"3A",X"1A",X"82",X"FE",X"78",X"30",X"07",X"3A",X"1C",X"82",X"FE",
		X"78",X"38",X"DF",X"21",X"33",X"86",X"7E",X"3C",X"3C",X"FD",X"77",X"08",X"FD",X"36",X"0A",X"16",
		X"11",X"80",X"04",X"DD",X"72",X"0A",X"DD",X"73",X"09",X"DD",X"36",X"04",X"00",X"DD",X"36",X"03",
		X"00",X"21",X"A9",X"4C",X"FD",X"75",X"05",X"FD",X"74",X"06",X"FD",X"36",X"04",X"01",X"FD",X"CB",
		X"00",X"E6",X"3E",X"0A",X"DD",X"77",X"01",X"DD",X"CB",X"00",X"CE",X"C9",X"3A",X"1A",X"82",X"FE",
		X"78",X"38",X"08",X"3A",X"1C",X"82",X"FE",X"78",X"DA",X"12",X"4A",X"21",X"34",X"86",X"7E",X"3D",
		X"3D",X"FD",X"77",X"08",X"FD",X"36",X"0A",X"16",X"11",X"80",X"FB",X"DD",X"72",X"0A",X"DD",X"73",
		X"09",X"DD",X"36",X"04",X"00",X"DD",X"36",X"03",X"00",X"21",X"70",X"4C",X"FD",X"75",X"05",X"FD",
		X"74",X"06",X"FD",X"36",X"04",X"01",X"FD",X"CB",X"00",X"E6",X"3E",X"0A",X"DD",X"77",X"01",X"DD",
		X"CB",X"00",X"CE",X"C9",X"3A",X"1A",X"82",X"FE",X"78",X"38",X"08",X"3A",X"1C",X"82",X"FE",X"78",
		X"D2",X"12",X"4A",X"21",X"34",X"86",X"7E",X"3D",X"3D",X"FD",X"77",X"08",X"FD",X"36",X"0A",X"D8",
		X"11",X"80",X"04",X"CD",X"BE",X"0F",X"DD",X"72",X"0A",X"DD",X"73",X"09",X"DD",X"36",X"04",X"00",
		X"DD",X"36",X"03",X"00",X"21",X"96",X"4C",X"FD",X"75",X"05",X"FD",X"74",X"06",X"FD",X"36",X"04",
		X"01",X"FD",X"CB",X"00",X"E6",X"3E",X"0A",X"DD",X"77",X"01",X"DD",X"CB",X"00",X"CE",X"C9",X"3A",
		X"1A",X"82",X"FE",X"78",X"30",X"08",X"3A",X"1C",X"82",X"FE",X"78",X"D2",X"12",X"4A",X"21",X"33",
		X"86",X"7E",X"3C",X"3C",X"FD",X"77",X"08",X"FD",X"36",X"0A",X"D8",X"11",X"80",X"04",X"DD",X"36",
		X"04",X"00",X"DD",X"36",X"03",X"00",X"DD",X"72",X"0A",X"DD",X"73",X"09",X"21",X"83",X"4C",X"FD",
		X"75",X"05",X"FD",X"74",X"06",X"FD",X"36",X"04",X"01",X"FD",X"CB",X"00",X"E6",X"3E",X"0A",X"DD",
		X"77",X"01",X"DD",X"CB",X"00",X"CE",X"C9",X"CD",X"4D",X"4C",X"3E",X"0B",X"CD",X"1F",X"08",X"DD",
		X"7E",X"0D",X"B7",X"C2",X"5F",X"4C",X"FD",X"CB",X"00",X"4E",X"20",X"0B",X"FD",X"36",X"01",X"05",
		X"FD",X"CB",X"00",X"CE",X"CD",X"74",X"4B",X"CD",X"7B",X"16",X"FD",X"E5",X"CD",X"BC",X"09",X"FD",
		X"E1",X"C3",X"4F",X"4B",X"CD",X"06",X"19",X"CD",X"39",X"4C",X"FE",X"01",X"20",X"12",X"21",X"80",
		X"03",X"FD",X"75",X"03",X"FD",X"74",X"04",X"FD",X"36",X"09",X"00",X"FD",X"36",X"0A",X"00",X"C9",
		X"FE",X"03",X"20",X"13",X"21",X"80",X"03",X"FD",X"75",X"03",X"FD",X"74",X"04",X"21",X"80",X"FC",
		X"FD",X"75",X"09",X"FD",X"74",X"0A",X"C9",X"FE",X"02",X"20",X"12",X"FD",X"36",X"03",X"00",X"FD",
		X"36",X"04",X"00",X"21",X"80",X"FC",X"FD",X"75",X"09",X"FD",X"74",X"0A",X"C9",X"FE",X"06",X"20",
		X"10",X"21",X"80",X"FC",X"FD",X"75",X"03",X"FD",X"74",X"04",X"FD",X"75",X"09",X"FD",X"74",X"0A",
		X"C9",X"FE",X"04",X"20",X"12",X"21",X"80",X"FC",X"FD",X"75",X"03",X"FD",X"74",X"04",X"FD",X"36",
		X"09",X"00",X"FD",X"36",X"0A",X"00",X"C9",X"FE",X"0C",X"20",X"13",X"21",X"80",X"FC",X"FD",X"75",
		X"03",X"FD",X"74",X"04",X"21",X"80",X"03",X"FD",X"75",X"09",X"FD",X"74",X"0A",X"C9",X"FE",X"08",
		X"20",X"12",X"FD",X"36",X"03",X"00",X"FD",X"36",X"04",X"00",X"21",X"80",X"03",X"FD",X"75",X"09",
		X"FD",X"74",X"0A",X"C9",X"FE",X"09",X"20",X"10",X"21",X"80",X"03",X"FD",X"75",X"03",X"FD",X"74",
		X"04",X"FD",X"75",X"09",X"FD",X"74",X"0A",X"C9",X"FD",X"36",X"03",X"00",X"FD",X"36",X"04",X"00",
		X"FD",X"36",X"09",X"00",X"FD",X"36",X"0A",X"00",X"C9",X"CD",X"42",X"08",X"FE",X"7F",X"38",X"02",
		X"78",X"C9",X"E6",X"0F",X"C9",X"CD",X"36",X"0A",X"CD",X"BC",X"09",X"18",X"FB",X"21",X"BC",X"4C",
		X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",X"36",X"04",X"01",X"DD",X"CB",X"00",X"E6",X"C9",X"3E",
		X"05",X"CD",X"1F",X"08",X"01",X"01",X"02",X"CD",X"57",X"1F",X"CD",X"01",X"15",X"C3",X"F6",X"48",
		X"00",X"00",X"01",X"00",X"00",X"0E",X"09",X"03",X"66",X"04",X"0E",X"09",X"03",X"65",X"04",X"00",
		X"01",X"75",X"4C",X"00",X"00",X"01",X"00",X"00",X"0E",X"09",X"04",X"A6",X"04",X"0E",X"09",X"04",
		X"A5",X"04",X"00",X"01",X"88",X"4C",X"00",X"00",X"01",X"00",X"00",X"09",X"0E",X"04",X"63",X"04",
		X"09",X"0E",X"04",X"64",X"04",X"00",X"01",X"9B",X"4C",X"00",X"00",X"01",X"00",X"00",X"09",X"0E",
		X"04",X"A3",X"04",X"09",X"0E",X"04",X"A4",X"04",X"00",X"01",X"AE",X"4C",X"00",X"00",X"01",X"00",
		X"00",X"0C",X"0C",X"02",X"1F",X"00",X"0C",X"0C",X"02",X"1E",X"01",X"0C",X"0C",X"02",X"1D",X"02",
		X"0C",X"0C",X"02",X"1E",X"03",X"0C",X"0C",X"02",X"1F",X"04",X"0C",X"0C",X"02",X"1E",X"05",X"0C",
		X"0C",X"02",X"1D",X"06",X"0C",X"0C",X"02",X"1E",X"07",X"00",X"01",X"C1",X"4C",X"CD",X"26",X"09",
		X"D2",X"E0",X"09",X"CD",X"CE",X"08",X"D2",X"43",X"4F",X"FD",X"2A",X"DA",X"80",X"FD",X"66",X"02",
		X"FD",X"6E",X"01",X"E5",X"DD",X"E1",X"CD",X"07",X"17",X"CD",X"4B",X"4F",X"FD",X"CB",X"00",X"F6",
		X"FD",X"CB",X"0C",X"D6",X"DD",X"CB",X"00",X"EE",X"FD",X"CB",X"00",X"D6",X"FD",X"36",X"0D",X"00",
		X"3E",X"0A",X"CD",X"1F",X"08",X"DD",X"E5",X"CD",X"BC",X"09",X"FD",X"E1",X"DD",X"7E",X"0D",X"B7",
		X"C2",X"32",X"4F",X"FD",X"CB",X"00",X"4E",X"20",X"0B",X"FD",X"36",X"01",X"0A",X"FD",X"CB",X"00",
		X"CE",X"CD",X"4E",X"4D",X"CD",X"54",X"4E",X"FD",X"E5",X"CD",X"BC",X"09",X"18",X"DC",X"CD",X"06",
		X"19",X"CD",X"1D",X"4F",X"DD",X"CB",X"00",X"A6",X"FE",X"01",X"20",X"17",X"21",X"50",X"02",X"FD",
		X"75",X"03",X"FD",X"74",X"04",X"FD",X"36",X"09",X"00",X"FD",X"36",X"0A",X"00",X"21",X"7A",X"4F",
		X"C3",X"41",X"4E",X"FE",X"03",X"20",X"18",X"21",X"50",X"02",X"FD",X"75",X"03",X"FD",X"74",X"04",
		X"21",X"B0",X"FD",X"FD",X"75",X"09",X"FD",X"74",X"0A",X"21",X"7A",X"4F",X"C3",X"41",X"4E",X"FE",
		X"02",X"20",X"17",X"FD",X"36",X"03",X"00",X"FD",X"36",X"04",X"00",X"21",X"B0",X"FD",X"FD",X"75",
		X"09",X"FD",X"74",X"0A",X"21",X"97",X"4F",X"C3",X"41",X"4E",X"FE",X"06",X"20",X"15",X"21",X"B0",
		X"FD",X"FD",X"75",X"03",X"FD",X"74",X"04",X"FD",X"75",X"09",X"FD",X"74",X"0A",X"21",X"5D",X"4F",
		X"C3",X"41",X"4E",X"FE",X"04",X"20",X"17",X"21",X"B0",X"FD",X"FD",X"75",X"03",X"FD",X"74",X"04",
		X"FD",X"36",X"09",X"00",X"FD",X"36",X"0A",X"00",X"21",X"5D",X"4F",X"C3",X"41",X"4E",X"FE",X"0C",
		X"20",X"18",X"21",X"B0",X"FD",X"FD",X"75",X"03",X"FD",X"74",X"04",X"21",X"50",X"02",X"FD",X"75",
		X"09",X"FD",X"74",X"0A",X"21",X"5D",X"4F",X"C3",X"41",X"4E",X"FE",X"08",X"20",X"17",X"FD",X"36",
		X"03",X"00",X"FD",X"36",X"04",X"00",X"21",X"50",X"02",X"FD",X"75",X"09",X"FD",X"74",X"0A",X"21",
		X"B4",X"4F",X"C3",X"41",X"4E",X"FE",X"09",X"20",X"15",X"21",X"50",X"02",X"FD",X"75",X"03",X"FD",
		X"74",X"04",X"FD",X"75",X"09",X"FD",X"74",X"0A",X"21",X"7A",X"4F",X"C3",X"41",X"4E",X"FD",X"36",
		X"03",X"00",X"FD",X"36",X"04",X"00",X"FD",X"36",X"09",X"00",X"FD",X"36",X"0A",X"00",X"21",X"B4",
		X"4F",X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",X"36",X"04",X"01",X"FD",X"CB",X"00",X"96",X"DD",
		X"CB",X"00",X"E6",X"C9",X"DD",X"7E",X"0A",X"FE",X"17",X"30",X"2A",X"FD",X"56",X"0A",X"FD",X"5E",
		X"09",X"CD",X"BE",X"0F",X"FD",X"72",X"0A",X"FD",X"73",X"09",X"3E",X"18",X"DD",X"77",X"0A",X"21",
		X"B4",X"4F",X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",X"36",X"04",X"01",X"FD",X"CB",X"00",X"96",
		X"DD",X"CB",X"00",X"E6",X"C9",X"DD",X"7E",X"0A",X"FE",X"D8",X"38",X"2A",X"FD",X"56",X"0A",X"FD",
		X"5E",X"09",X"CD",X"BE",X"0F",X"FD",X"72",X"0A",X"FD",X"73",X"09",X"3E",X"D6",X"DD",X"77",X"0A",
		X"21",X"97",X"4F",X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",X"36",X"04",X"01",X"FD",X"CB",X"00",
		X"96",X"DD",X"CB",X"00",X"E6",X"C9",X"21",X"34",X"86",X"DD",X"7E",X"08",X"BE",X"38",X"2B",X"FD",
		X"56",X"04",X"FD",X"5E",X"03",X"CD",X"BE",X"0F",X"FD",X"72",X"04",X"FD",X"73",X"03",X"7E",X"3D",
		X"3D",X"DD",X"77",X"08",X"21",X"5D",X"4F",X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",X"36",X"04",
		X"01",X"FD",X"CB",X"00",X"96",X"DD",X"CB",X"00",X"E6",X"C9",X"21",X"33",X"86",X"DD",X"7E",X"08",
		X"BE",X"D0",X"FD",X"56",X"04",X"FD",X"5E",X"03",X"CD",X"BE",X"0F",X"FD",X"72",X"04",X"FD",X"73",
		X"03",X"7E",X"3C",X"3C",X"DD",X"77",X"08",X"21",X"7A",X"4F",X"DD",X"75",X"05",X"DD",X"74",X"06",
		X"DD",X"36",X"04",X"01",X"FD",X"CB",X"00",X"96",X"DD",X"CB",X"00",X"E6",X"C9",X"CD",X"42",X"08",
		X"FE",X"4B",X"30",X"04",X"78",X"E6",X"0A",X"C9",X"FE",X"AF",X"30",X"02",X"78",X"C9",X"78",X"E6",
		X"05",X"C9",X"3E",X"05",X"CD",X"1F",X"08",X"01",X"01",X"02",X"CD",X"57",X"1F",X"CD",X"01",X"15",
		X"C3",X"F9",X"4C",X"CD",X"36",X"0A",X"CD",X"BC",X"09",X"18",X"FB",X"21",X"5D",X"4F",X"FD",X"75",
		X"05",X"FD",X"74",X"06",X"FD",X"36",X"04",X"01",X"FD",X"CB",X"00",X"E6",X"C9",X"00",X"00",X"01",
		X"00",X"00",X"0C",X"0C",X"02",X"39",X"07",X"0C",X"0C",X"02",X"38",X"07",X"0C",X"0C",X"02",X"36",
		X"07",X"0C",X"0C",X"02",X"37",X"07",X"00",X"01",X"62",X"4F",X"00",X"00",X"01",X"00",X"00",X"0C",
		X"0C",X"02",X"B9",X"07",X"0C",X"0C",X"02",X"B8",X"07",X"0C",X"0C",X"02",X"B6",X"07",X"0C",X"0C",
		X"02",X"B7",X"07",X"00",X"01",X"7F",X"4F",X"00",X"00",X"01",X"00",X"00",X"0C",X"0C",X"02",X"3B",
		X"07",X"0C",X"0C",X"02",X"3A",X"07",X"0C",X"0C",X"02",X"BB",X"07",X"0C",X"0C",X"02",X"BA",X"07",
		X"00",X"01",X"9C",X"4F",X"00",X"00",X"01",X"00",X"00",X"0C",X"0C",X"02",X"3D",X"07",X"0C",X"0C",
		X"02",X"3C",X"07",X"0C",X"0C",X"02",X"BD",X"07",X"0C",X"0C",X"02",X"BC",X"07",X"00",X"01",X"B9",
		X"4F",X"3E",X"FF",X"32",X"55",X"85",X"3E",X"01",X"32",X"46",X"86",X"CD",X"69",X"0A",X"CD",X"60",
		X"1A",X"CD",X"82",X"05",X"CF",X"18",X"18",X"5B",X"53",X"43",X"4F",X"52",X"49",X"4E",X"47",X"20",
		X"47",X"4F",X"45",X"53",X"20",X"41",X"53",X"20",X"46",X"4F",X"4C",X"4C",X"4F",X"57",X"53",X"5B",
		X"00",X"CF",X"10",X"28",X"46",X"41",X"43",X"45",X"20",X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",
		X"5D",X"5D",X"5D",X"5D",X"5D",X"20",X"20",X"35",X"30",X"20",X"50",X"4F",X"49",X"4E",X"54",X"53",
		X"00",X"CF",X"10",X"38",X"45",X"59",X"45",X"42",X"41",X"4C",X"4C",X"20",X"5D",X"5D",X"5D",X"5D",
		X"5D",X"5D",X"5D",X"5D",X"5D",X"20",X"20",X"35",X"30",X"20",X"50",X"4F",X"49",X"4E",X"54",X"53",
		X"00",X"CF",X"10",X"48",X"53",X"51",X"55",X"49",X"44",X"20",X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",
		X"5D",X"5D",X"5D",X"5D",X"5D",X"20",X"20",X"37",X"30",X"20",X"50",X"4F",X"49",X"4E",X"54",X"53",
		X"00",X"CF",X"10",X"58",X"53",X"49",X"43",X"4B",X"4C",X"45",X"20",X"5D",X"5D",X"5D",X"5D",X"5D",
		X"5D",X"5D",X"5D",X"5D",X"5D",X"20",X"20",X"36",X"30",X"20",X"50",X"4F",X"49",X"4E",X"54",X"53",
		X"00",X"CF",X"10",X"68",X"43",X"41",X"54",X"45",X"52",X"50",X"49",X"4C",X"4C",X"41",X"52",X"20",
		X"5D",X"5D",X"5D",X"5D",X"5D",X"20",X"20",X"35",X"30",X"20",X"50",X"4F",X"49",X"4E",X"54",X"53",
		X"00",X"CF",X"10",X"78",X"42",X"55",X"54",X"54",X"45",X"52",X"46",X"4C",X"59",X"20",X"5D",X"5D",
		X"5D",X"5D",X"5D",X"5D",X"5D",X"20",X"31",X"30",X"30",X"20",X"50",X"4F",X"49",X"4E",X"54",X"53",
		X"00",X"CF",X"10",X"88",X"50",X"52",X"4F",X"50",X"45",X"4C",X"4C",X"45",X"52",X"20",X"5D",X"5D",
		X"5D",X"5D",X"5D",X"5D",X"5D",X"20",X"20",X"34",X"30",X"20",X"50",X"4F",X"49",X"4E",X"54",X"53",
		X"00",X"CF",X"10",X"98",X"43",X"59",X"43",X"4C",X"4F",X"54",X"52",X"4F",X"4E",X"20",X"5D",X"5D",
		X"5D",X"5D",X"5D",X"5D",X"5D",X"20",X"20",X"36",X"30",X"20",X"50",X"4F",X"49",X"4E",X"54",X"53",
		X"00",X"CF",X"10",X"A8",X"54",X"41",X"5A",X"5A",X"20",X"4D",X"45",X"4E",X"20",X"5D",X"5D",X"5D",
		X"5D",X"5D",X"5D",X"5D",X"5D",X"20",X"31",X"30",X"30",X"20",X"50",X"4F",X"49",X"4E",X"54",X"53",
		X"00",X"CF",X"10",X"B8",X"48",X"4F",X"50",X"50",X"45",X"52",X"53",X"20",X"5D",X"5D",X"5D",X"5D",
		X"5D",X"5D",X"5D",X"5D",X"5D",X"20",X"32",X"30",X"30",X"20",X"50",X"4F",X"49",X"4E",X"54",X"53",
		X"00",X"CF",X"10",X"C8",X"4C",X"49",X"54",X"54",X"4C",X"45",X"20",X"48",X"4F",X"50",X"50",X"45",
		X"52",X"53",X"20",X"5D",X"5D",X"20",X"20",X"32",X"30",X"20",X"50",X"4F",X"49",X"4E",X"54",X"53",
		X"00",X"06",X"32",X"CD",X"E3",X"53",X"CD",X"82",X"05",X"CF",X"20",X"28",X"55",X"53",X"45",X"20",
		X"54",X"48",X"45",X"20",X"4A",X"4F",X"59",X"53",X"54",X"49",X"43",X"4B",X"20",X"54",X"4F",X"20",
		X"52",X"55",X"4E",X"00",X"CF",X"40",X"38",X"41",X"52",X"4F",X"55",X"4E",X"44",X"20",X"54",X"48",
		X"45",X"20",X"52",X"4F",X"4F",X"4D",X"5D",X"00",X"CF",X"20",X"48",X"54",X"4F",X"20",X"53",X"48",
		X"4F",X"4F",X"54",X"20",X"50",X"52",X"45",X"53",X"53",X"20",X"54",X"48",X"45",X"20",X"46",X"49",
		X"52",X"45",X"00",X"CF",X"20",X"58",X"42",X"55",X"54",X"54",X"4F",X"4E",X"20",X"41",X"4E",X"44",
		X"20",X"41",X"49",X"4D",X"20",X"57",X"49",X"54",X"48",X"20",X"54",X"48",X"45",X"00",X"CF",X"10",
		X"68",X"4A",X"4F",X"59",X"53",X"54",X"49",X"43",X"4B",X"5D",X"20",X"48",X"4F",X"4C",X"44",X"20",
		X"44",X"4F",X"57",X"4E",X"20",X"54",X"48",X"45",X"20",X"46",X"49",X"52",X"45",X"00",X"CF",X"28",
		X"78",X"42",X"55",X"54",X"54",X"4F",X"4E",X"20",X"46",X"4F",X"52",X"20",X"52",X"41",X"50",X"49",
		X"44",X"20",X"46",X"49",X"52",X"45",X"5D",X"00",X"CF",X"10",X"88",X"57",X"48",X"45",X"4E",X"20",
		X"41",X"4C",X"4C",X"20",X"54",X"48",X"45",X"20",X"4C",X"49",X"54",X"54",X"4C",X"45",X"20",X"48",
		X"4F",X"50",X"50",X"45",X"52",X"53",X"00",X"CF",X"18",X"98",X"41",X"52",X"45",X"20",X"47",X"4F",
		X"4E",X"45",X"20",X"54",X"48",X"45",X"20",X"44",X"4F",X"4F",X"52",X"53",X"20",X"41",X"54",X"20",
		X"54",X"48",X"45",X"00",X"CF",X"18",X"A8",X"54",X"4F",X"50",X"20",X"41",X"4E",X"44",X"20",X"54",
		X"48",X"45",X"20",X"42",X"4F",X"54",X"54",X"4F",X"4D",X"20",X"4F",X"46",X"20",X"54",X"48",X"45",
		X"00",X"CF",X"40",X"B8",X"52",X"4F",X"4F",X"4D",X"20",X"57",X"49",X"4C",X"4C",X"20",X"4F",X"50",
		X"45",X"4E",X"5D",X"00",X"06",X"32",X"CD",X"E3",X"53",X"CD",X"F0",X"53",X"CD",X"82",X"05",X"CF",
		X"18",X"28",X"45",X"56",X"45",X"52",X"59",X"20",X"43",X"4F",X"55",X"50",X"4C",X"45",X"20",X"4F",
		X"46",X"20",X"52",X"4F",X"4F",X"4D",X"53",X"20",X"49",X"53",X"20",X"41",X"00",X"CF",X"30",X"38",
		X"42",X"4F",X"4E",X"55",X"53",X"20",X"52",X"4F",X"4F",X"4D",X"5D",X"20",X"52",X"55",X"4E",X"20",
		X"4F",X"56",X"45",X"52",X"00",X"CF",X"20",X"48",X"41",X"4C",X"4C",X"20",X"54",X"48",X"45",X"20",
		X"50",X"4F",X"49",X"4E",X"54",X"53",X"20",X"59",X"4F",X"55",X"20",X"43",X"41",X"4E",X"5D",X"00",
		X"CF",X"30",X"58",X"41",X"4C",X"53",X"4F",X"20",X"49",X"4E",X"20",X"54",X"48",X"45",X"20",X"52",
		X"4F",X"4F",X"4D",X"20",X"41",X"52",X"45",X"00",X"CF",X"20",X"68",X"54",X"57",X"4F",X"20",X"42",
		X"4F",X"4D",X"42",X"53",X"5D",X"20",X"52",X"55",X"4E",X"20",X"4F",X"56",X"45",X"52",X"20",X"54",
		X"48",X"45",X"00",X"CF",X"28",X"78",X"42",X"4F",X"4D",X"42",X"53",X"20",X"54",X"4F",X"20",X"50",
		X"49",X"43",X"4B",X"20",X"54",X"48",X"45",X"4D",X"20",X"55",X"50",X"5D",X"00",X"CF",X"10",X"88",
		X"59",X"4F",X"55",X"20",X"43",X"41",X"4E",X"20",X"55",X"53",X"45",X"20",X"54",X"48",X"45",X"20",
		X"42",X"4F",X"4D",X"42",X"53",X"20",X"49",X"4E",X"20",X"41",X"4E",X"59",X"00",X"CF",X"30",X"98",
		X"4F",X"46",X"20",X"54",X"48",X"45",X"20",X"4F",X"54",X"48",X"45",X"52",X"20",X"52",X"4F",X"4F",
		X"4D",X"53",X"5D",X"00",X"06",X"28",X"CD",X"E3",X"53",X"CD",X"46",X"54",X"CD",X"82",X"05",X"CF",
		X"20",X"28",X"54",X"48",X"45",X"20",X"42",X"4F",X"4D",X"42",X"53",X"20",X"44",X"4F",X"20",X"54",
		X"57",X"4F",X"20",X"54",X"48",X"49",X"4E",X"47",X"53",X"00",X"CF",X"20",X"38",X"46",X"49",X"52",
		X"53",X"54",X"20",X"54",X"48",X"45",X"59",X"20",X"4B",X"49",X"4C",X"4C",X"20",X"41",X"4C",X"4C",
		X"20",X"54",X"48",X"45",X"00",X"CF",X"40",X"48",X"41",X"54",X"54",X"41",X"43",X"4B",X"49",X"4E",
		X"47",X"20",X"45",X"4E",X"45",X"4D",X"59",X"5D",X"00",X"CF",X"30",X"58",X"53",X"45",X"43",X"4F",
		X"4E",X"44",X"20",X"54",X"48",X"45",X"59",X"20",X"53",X"54",X"4F",X"50",X"20",X"54",X"48",X"45",
		X"00",X"CF",X"40",X"68",X"43",X"52",X"55",X"53",X"48",X"49",X"4E",X"47",X"20",X"57",X"41",X"4C",
		X"4C",X"53",X"5D",X"00",X"06",X"1E",X"CD",X"E3",X"53",X"CD",X"8C",X"54",X"AF",X"32",X"46",X"86",
		X"C3",X"2E",X"1A",X"3E",X"FE",X"32",X"40",X"86",X"3E",X"04",X"CD",X"88",X"1A",X"10",X"F4",X"C9",
		X"21",X"65",X"8B",X"06",X"17",X"CD",X"BA",X"54",X"21",X"E7",X"8A",X"06",X"10",X"CD",X"BA",X"54",
		X"21",X"69",X"8B",X"06",X"17",X"CD",X"BA",X"54",X"21",X"6B",X"8B",X"06",X"17",X"CD",X"BA",X"54",
		X"21",X"AD",X"8B",X"06",X"1C",X"CD",X"BA",X"54",X"21",X"4F",X"8B",X"06",X"16",X"CD",X"BA",X"54",
		X"21",X"B1",X"8B",X"06",X"1B",X"CD",X"BA",X"54",X"21",X"93",X"8B",X"06",X"19",X"CD",X"BA",X"54",
		X"21",X"95",X"8B",X"06",X"19",X"CD",X"BA",X"54",X"21",X"F7",X"8A",X"06",X"0F",X"CD",X"BA",X"54",
		X"3E",X"02",X"CD",X"7D",X"1A",X"C9",X"21",X"85",X"8B",X"06",X"1A",X"CD",X"BA",X"54",X"21",X"27",
		X"8B",X"06",X"14",X"CD",X"BA",X"54",X"21",X"69",X"8B",X"06",X"17",X"CD",X"BA",X"54",X"21",X"2B",
		X"8B",X"06",X"14",X"CD",X"BA",X"54",X"21",X"6D",X"8B",X"06",X"17",X"CD",X"BA",X"54",X"21",X"4F",
		X"8B",X"06",X"16",X"CD",X"BA",X"54",X"21",X"B1",X"8B",X"06",X"1C",X"CD",X"BA",X"54",X"21",X"33",
		X"8B",X"06",X"13",X"CD",X"BA",X"54",X"3E",X"02",X"CD",X"7D",X"1A",X"C9",X"21",X"65",X"8B",X"06",
		X"17",X"CD",X"BA",X"54",X"21",X"67",X"8B",X"06",X"17",X"CD",X"BA",X"54",X"21",X"E9",X"8A",X"06",
		X"10",X"CD",X"BA",X"54",X"21",X"2B",X"8B",X"06",X"14",X"CD",X"BA",X"54",X"21",X"ED",X"8A",X"06",
		X"0F",X"CD",X"BA",X"54",X"3E",X"02",X"CD",X"7D",X"1A",X"C9",X"11",X"20",X"00",X"D5",X"E5",X"C5",
		X"CD",X"58",X"0F",X"21",X"47",X"86",X"34",X"7E",X"E6",X"03",X"20",X"05",X"3E",X"FE",X"32",X"40",
		X"86",X"3E",X"01",X"CD",X"88",X"1A",X"C1",X"E1",X"D1",X"AF",X"ED",X"52",X"10",X"DF",X"C9",X"6D",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
