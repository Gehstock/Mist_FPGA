library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity GALAXIAN_1H is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of GALAXIAN_1H is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",X"00",X"02",X"02",X"FE",X"FE",X"42",X"02",X"00",X"00",
		X"62",X"F2",X"BA",X"9A",X"9E",X"CE",X"46",X"00",X"8C",X"DE",X"F2",X"B2",X"92",X"86",X"04",X"00",
		X"08",X"FE",X"FE",X"C8",X"68",X"38",X"18",X"00",X"1C",X"BE",X"A2",X"A2",X"A2",X"E6",X"E4",X"00",
		X"0C",X"9E",X"92",X"92",X"D2",X"7E",X"3C",X"00",X"C0",X"E0",X"B0",X"9E",X"8E",X"C0",X"C0",X"00",
		X"0C",X"6E",X"9A",X"9A",X"B2",X"F2",X"6C",X"00",X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",X"00",
		X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",
		X"44",X"C6",X"82",X"82",X"C6",X"7C",X"38",X"00",X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",
		X"82",X"92",X"92",X"92",X"FE",X"FE",X"00",X"00",X"80",X"90",X"90",X"90",X"90",X"FE",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",
		X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",X"44",X"C6",X"82",X"82",X"C6",X"7C",X"38",X"00",
		X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",X"82",X"92",X"92",X"92",X"FE",X"FE",X"00",X"00",
		X"80",X"90",X"90",X"90",X"90",X"FE",X"FE",X"00",X"9E",X"9E",X"92",X"82",X"C6",X"7C",X"38",X"00",
		X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",X"82",X"82",X"FE",X"FE",X"82",X"82",X"00",X"00",
		X"FC",X"FE",X"02",X"02",X"02",X"06",X"04",X"00",X"82",X"C6",X"6E",X"3C",X"18",X"FE",X"FE",X"00",
		X"02",X"02",X"02",X"02",X"FE",X"FE",X"00",X"00",X"FE",X"FE",X"70",X"38",X"70",X"FE",X"FE",X"00",
		X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",X"00",
		X"70",X"F8",X"88",X"88",X"88",X"FE",X"FE",X"00",X"7A",X"FC",X"8E",X"8A",X"82",X"FE",X"7C",X"00",
		X"72",X"F6",X"9E",X"8C",X"88",X"FE",X"FE",X"00",X"0C",X"5E",X"D2",X"92",X"92",X"F6",X"64",X"00",
		X"80",X"80",X"FE",X"FE",X"80",X"80",X"00",X"00",X"FC",X"FE",X"02",X"02",X"02",X"FE",X"FC",X"00",
		X"F0",X"F8",X"1C",X"0E",X"1C",X"F8",X"F0",X"00",X"F8",X"FE",X"1C",X"38",X"1C",X"FE",X"F8",X"00",
		X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",X"C0",X"F0",X"1E",X"1E",X"F0",X"C0",X"00",X"00",
		X"C2",X"E2",X"F2",X"BA",X"9E",X"8E",X"86",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"00",
		X"FF",X"FF",X"F7",X"FF",X"FF",X"FE",X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",X"FF",X"DF",X"FF",X"FD",
		X"BF",X"F7",X"FF",X"FF",X"FF",X"FF",X"DF",X"FF",X"FF",X"FF",X"FF",X"DF",X"FF",X"FF",X"FB",X"FF",
		X"B0",X"C0",X"82",X"C3",X"C2",X"81",X"83",X"81",X"03",X"07",X"1F",X"77",X"EB",X"ED",X"36",X"DB",
		X"C3",X"82",X"C1",X"81",X"82",X"C3",X"A0",X"F0",X"67",X"36",X"6D",X"E3",X"7F",X"DF",X"07",X"03",
		X"FF",X"FF",X"DF",X"AF",X"A1",X"BE",X"A9",X"D4",X"F7",X"FF",X"E7",X"DB",X"A1",X"40",X"C0",X"18",
		X"FA",X"FD",X"FE",X"FF",X"FF",X"FD",X"DF",X"FF",X"21",X"C0",X"40",X"00",X"81",X"C3",X"E7",X"FF",
		X"F0",X"EF",X"DF",X"BF",X"BF",X"BF",X"BF",X"3F",X"0F",X"E7",X"E3",X"F1",X"F8",X"F0",X"F0",X"F8",
		X"0F",X"BF",X"BF",X"BF",X"BF",X"DF",X"EF",X"F0",X"F0",X"E0",X"F8",X"F0",X"F1",X"E3",X"E7",X"1F",
		X"FF",X"FD",X"F2",X"F2",X"E9",X"CF",X"C9",X"D5",X"F7",X"FF",X"FF",X"7F",X"3F",X"9F",X"CF",X"F5",
		X"9F",X"C9",X"C7",X"E1",X"F6",X"FA",X"DD",X"FF",X"F7",X"CF",X"9F",X"3F",X"7F",X"FF",X"FB",X"FF",
		X"F8",X"C0",X"B0",X"78",X"48",X"48",X"B0",X"C0",X"00",X"00",X"60",X"20",X"21",X"61",X"40",X"40",
		X"C0",X"B0",X"48",X"48",X"78",X"B0",X"C0",X"F8",X"40",X"40",X"61",X"21",X"20",X"60",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"FF",X"FF",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"7F",X"37",X"3F",X"7F",X"7E",X"7F",X"3F",X"F4",X"FC",X"FC",X"FC",X"F8",X"DC",X"FC",X"FC",
		X"1F",X"17",X"3F",X"3F",X"3F",X"0F",X"1F",X"3F",X"F8",X"F8",X"FC",X"DC",X"FC",X"FE",X"FA",X"FE",
		X"00",X"00",X"04",X"0C",X"1C",X"3C",X"7C",X"7A",X"00",X"C0",X"C0",X"D8",X"D8",X"F8",X"78",X"FC",
		X"7F",X"79",X"3F",X"06",X"00",X"00",X"00",X"00",X"FE",X"FE",X"74",X"34",X"30",X"30",X"00",X"00",
		X"00",X"00",X"08",X"18",X"3C",X"7C",X"7C",X"7A",X"00",X"00",X"00",X"18",X"3C",X"7C",X"7E",X"FE",
		X"7F",X"79",X"3F",X"06",X"00",X"00",X"00",X"00",X"FE",X"FC",X"78",X"30",X"30",X"30",X"00",X"00",
		X"00",X"00",X"10",X"18",X"3C",X"3C",X"7C",X"7A",X"00",X"30",X"30",X"30",X"70",X"FC",X"7C",X"FC",
		X"7F",X"79",X"3F",X"06",X"00",X"00",X"00",X"00",X"F8",X"F8",X"F0",X"D0",X"C0",X"C0",X"00",X"00",
		X"00",X"03",X"0F",X"03",X"3F",X"3F",X"07",X"03",X"00",X"00",X"80",X"F8",X"F8",X"E0",X"FE",X"BE",
		X"07",X"0D",X"0D",X"07",X"07",X"07",X"03",X"00",X"00",X"80",X"7C",X"F8",X"F0",X"E0",X"C0",X"00",
		X"00",X"01",X"03",X"07",X"3F",X"3F",X"07",X"03",X"00",X"C0",X"F0",X"F8",X"F8",X"F0",X"80",X"80",
		X"07",X"0D",X"0D",X"07",X"07",X"07",X"03",X"00",X"00",X"80",X"70",X"FC",X"F8",X"F0",X"E0",X"00",
		X"00",X"00",X"00",X"03",X"0F",X"07",X"3F",X"3F",X"00",X"00",X"E0",X"E0",X"FE",X"FE",X"F0",X"A0",
		X"07",X"0D",X"0D",X"07",X"07",X"07",X"03",X"00",X"00",X"80",X"70",X"F8",X"FC",X"F0",X"C0",X"00",
		X"FF",X"1F",X"17",X"1F",X"3F",X"FE",X"1F",X"1F",X"F7",X"F8",X"F8",X"F8",X"F8",X"DF",X"FC",X"F8",
		X"1F",X"17",X"FF",X"1F",X"1F",X"1F",X"1F",X"FF",X"F8",X"F8",X"FF",X"D8",X"F8",X"FC",X"F8",X"FF",
		X"FF",X"FE",X"FA",X"F1",X"E4",X"F0",X"F9",X"F1",X"1F",X"AF",X"97",X"4B",X"BC",X"C7",X"3F",X"E0",
		X"AE",X"F0",X"FB",X"F0",X"E5",X"F0",X"DB",X"FF",X"0F",X"E8",X"97",X"69",X"8A",X"15",X"C5",X"EB",
		X"FF",X"FF",X"F7",X"FD",X"F8",X"F2",X"F9",X"FC",X"CF",X"B7",X"7B",X"7D",X"BE",X"0E",X"C7",X"3F",
		X"BE",X"F9",X"F2",X"E4",X"F1",X"FB",X"DF",X"FF",X"D3",X"2E",X"DE",X"BD",X"7B",X"77",X"0F",X"FF",
		X"00",X"00",X"19",X"35",X"35",X"3D",X"19",X"01",X"00",X"00",X"40",X"40",X"40",X"40",X"40",X"40",
		X"19",X"35",X"35",X"3C",X"18",X"00",X"00",X"00",X"40",X"40",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"32",X"4A",X"4A",X"7A",X"32",X"02",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"10",
		X"32",X"4A",X"4B",X"79",X"30",X"00",X"00",X"00",X"10",X"10",X"30",X"E0",X"00",X"00",X"00",X"00",
		X"7F",X"3F",X"0F",X"03",X"00",X"00",X"00",X"00",X"FC",X"7F",X"3F",X"7F",X"FC",X"F0",X"F0",X"FC",
		X"1F",X"1F",X"3F",X"7F",X"FF",X"FC",X"F0",X"F0",X"1C",X"1E",X"0F",X"0F",X"1F",X"1C",X"1C",X"1C",
		X"F0",X"F0",X"F8",X"7F",X"3F",X"1F",X"1E",X"1C",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"7C",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"01",X"03",X"07",X"0F",X"1F",X"3E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"30",
		X"3F",X"00",X"1C",X"26",X"3E",X"1C",X"00",X"00",X"E0",X"00",X"70",X"98",X"F8",X"70",X"00",X"00",
		X"00",X"00",X"00",X"00",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"30",X"10",X"10",
		X"00",X"3F",X"00",X"1C",X"26",X"26",X"1C",X"00",X"30",X"E0",X"00",X"70",X"98",X"98",X"70",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"04",X"08",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",
		X"08",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"20",X"20",X"40",X"80",X"00",X"00",X"00",X"00",
		X"03",X"03",X"0B",X"1F",X"73",X"7F",X"7F",X"73",X"00",X"00",X"00",X"9C",X"FE",X"FE",X"F8",X"F0",
		X"1F",X"0B",X"03",X"7B",X"79",X"7D",X"3C",X"1E",X"F0",X"F8",X"7C",X"B8",X"98",X"80",X"00",X"00",
		X"00",X"01",X"07",X"1E",X"3C",X"7F",X"7F",X"3F",X"00",X"80",X"C0",X"40",X"E0",X"98",X"FC",X"FC",
		X"7F",X"7C",X"3E",X"3D",X"1E",X"1E",X"0C",X"00",X"94",X"E0",X"60",X"F0",X"78",X"38",X"00",X"00",
		X"00",X"00",X"1C",X"1E",X"1F",X"0F",X"07",X"07",X"0C",X"0C",X"0C",X"0C",X"CC",X"9C",X"F2",X"FE",
		X"1F",X"3F",X"3F",X"07",X"00",X"00",X"00",X"00",X"FE",X"F2",X"9C",X"CC",X"0C",X"0C",X"0C",X"0C",
		X"00",X"00",X"00",X"00",X"01",X"73",X"53",X"51",X"0C",X"CC",X"CC",X"CC",X"CC",X"9C",X"F2",X"FE",
		X"51",X"53",X"73",X"01",X"00",X"00",X"00",X"00",X"FE",X"F2",X"9C",X"CC",X"CC",X"CC",X"CC",X"0C",
		X"BD",X"40",X"80",X"00",X"80",X"80",X"80",X"00",X"78",X"70",X"70",X"79",X"3F",X"1F",X"0F",X"03",
		X"00",X"00",X"00",X"00",X"03",X"0F",X"1F",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"83",
		X"00",X"E0",X"F8",X"FE",X"FF",X"3F",X"0F",X"03",X"00",X"00",X"C0",X"00",X"01",X"07",X"0F",X"07",
		X"FE",X"FE",X"F8",X"E0",X"01",X"07",X"0F",X"07",X"3F",X"7F",X"7F",X"3F",X"1F",X"00",X"00",X"00",
		X"1F",X"3F",X"FF",X"FF",X"FF",X"FF",X"3F",X"3F",X"7F",X"7F",X"3F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"07",X"1F",X"3F",X"3F",X"7F",X"F0",X"F0",X"F8",X"FC",X"FE",X"FC",X"C0",X"00",
		X"F0",X"E0",X"E1",X"E1",X"E1",X"E1",X"E1",X"E0",X"FF",X"3F",X"FF",X"FF",X"FF",X"FC",X"F8",X"F0",
		X"E1",X"E1",X"E1",X"E0",X"E0",X"E0",X"F0",X"F8",X"0F",X"1F",X"3F",X"7F",X"F8",X"F0",X"E0",X"E0",
		X"F8",X"78",X"78",X"78",X"F8",X"F8",X"F0",X"E0",X"F8",X"78",X"78",X"78",X"F8",X"F0",X"E0",X"F0",
		X"F8",X"78",X"78",X"78",X"F8",X"F0",X"E0",X"F0",X"FF",X"FF",X"FF",X"F8",X"F8",X"78",X"78",X"78",
		X"F8",X"FC",X"FE",X"FE",X"FE",X"1E",X"1F",X"1F",X"FC",X"FC",X"FC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"E0",X"F0",X"F8",X"FC",X"FC",X"7C",X"00",X"00",X"00",X"00",X"01",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"F0",X"F8",X"FC",X"FE",X"1F",X"0F",X"07",X"07",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"80",X"80",X"80",X"80",X"80",X"80",X"82",X"82",X"01",X"01",X"01",X"01",X"01",X"01",X"21",X"A1",
		X"82",X"83",X"80",X"80",X"80",X"80",X"80",X"FF",X"A1",X"E1",X"01",X"01",X"01",X"01",X"01",X"FF",
		X"80",X"80",X"80",X"80",X"80",X"80",X"83",X"80",X"01",X"01",X"01",X"01",X"01",X"01",X"61",X"81",
		X"80",X"83",X"80",X"80",X"80",X"80",X"80",X"80",X"81",X"61",X"01",X"01",X"01",X"01",X"01",X"01",
		X"80",X"80",X"80",X"80",X"80",X"80",X"82",X"82",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"83",X"82",X"82",X"80",X"80",X"80",X"80",X"80",X"E1",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"80",X"80",X"80",X"80",X"80",X"80",X"81",X"82",X"01",X"01",X"01",X"01",X"01",X"01",X"21",X"A1",
		X"82",X"83",X"80",X"80",X"80",X"80",X"80",X"80",X"C1",X"E1",X"01",X"01",X"01",X"01",X"01",X"01",
		X"FF",X"80",X"80",X"80",X"80",X"80",X"81",X"82",X"FF",X"01",X"01",X"01",X"01",X"01",X"E1",X"81",
		X"82",X"81",X"80",X"80",X"80",X"80",X"80",X"80",X"81",X"E1",X"01",X"01",X"01",X"01",X"01",X"01",
		X"00",X"0F",X"3F",X"7F",X"4F",X"4C",X"48",X"78",X"00",X"E0",X"F0",X"F8",X"F8",X"18",X"00",X"00",
		X"78",X"48",X"4C",X"4F",X"7F",X"3F",X"0F",X"00",X"00",X"00",X"18",X"F8",X"F8",X"F0",X"E0",X"00",
		X"00",X"0F",X"3F",X"7F",X"4F",X"4C",X"48",X"7B",X"00",X"E0",X"F0",X"F8",X"F8",X"F8",X"78",X"28",
		X"7B",X"49",X"4D",X"4F",X"7F",X"3F",X"0F",X"00",X"20",X"F0",X"F8",X"F8",X"F8",X"F0",X"E0",X"00",
		X"00",X"0F",X"3F",X"7F",X"4F",X"4C",X"48",X"7B",X"00",X"E0",X"F0",X"F8",X"F8",X"F8",X"70",X"20",
		X"7B",X"49",X"4D",X"4F",X"7F",X"3F",X"0F",X"00",X"28",X"F8",X"F8",X"F8",X"F8",X"F0",X"E0",X"00",
		X"7C",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"C7",X"00",X"00",X"00",X"00",
		X"E3",X"E7",X"E7",X"C7",X"07",X"07",X"0F",X"1F",X"CF",X"FF",X"FF",X"FF",X"F0",X"E0",X"E0",X"E0",
		X"FE",X"FC",X"F8",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"1E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0E",X"1E",X"1C",X"3C",X"78",X"F8",X"FC",X"3E",X"0E",X"0F",X"0F",X"07",X"07",X"07",X"0F",X"0F",
		X"FE",X"FC",X"F8",X"F0",X"F8",X"3C",X"1C",X"1E",X"07",X"87",X"87",X"87",X"07",X"07",X"0F",X"1F",
		X"B0",X"C0",X"82",X"C3",X"C2",X"80",X"83",X"80",X"07",X"03",X"01",X"E1",X"03",X"01",X"E0",X"01",
		X"C3",X"80",X"C3",X"80",X"82",X"C3",X"A0",X"F0",X"61",X"82",X"61",X"01",X"A3",X"E1",X"01",X"03",
		X"00",X"10",X"70",X"E0",X"80",X"80",X"80",X"E0",X"00",X"08",X"08",X"04",X"04",X"04",X"04",X"04",
		X"E0",X"80",X"80",X"80",X"E0",X"70",X"10",X"00",X"04",X"04",X"04",X"04",X"04",X"08",X"08",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
