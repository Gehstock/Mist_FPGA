library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity spr_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of spr_rom is
	type rom is array(0 to  32767) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"ED",X"C0",X"00",X"FF",X"00",X"00",X"05",X"33",X"30",X"00",X"FF",X"00",X"00",
		X"55",X"66",X"65",X"00",X"FF",X"00",X"05",X"51",X"44",X"44",X"50",X"FF",X"00",X"03",X"55",X"67",
		X"88",X"70",X"FF",X"00",X"44",X"35",X"67",X"99",X"85",X"FF",X"04",X"56",X"7A",X"55",X"55",X"55",
		X"FF",X"04",X"58",X"6A",X"58",X"98",X"86",X"FF",X"0A",X"45",X"A3",X"55",X"56",X"66",X"FF",X"AA",
		X"AA",X"43",X"55",X"56",X"6A",X"FF",X"0A",X"A4",X"41",X"4A",X"AA",X"50",X"FF",X"00",X"AA",X"33",
		X"55",X"55",X"A0",X"FF",X"00",X"0A",X"A3",X"33",X"3A",X"00",X"FF",X"00",X"00",X"AA",X"ED",X"CA",
		X"00",X"FF",X"00",X"00",X"A0",X"00",X"00",X"00",X"FF",X"00",X"0A",X"A3",X"30",X"00",X"00",X"FF",
		X"00",X"AA",X"34",X"63",X"00",X"00",X"FF",X"0A",X"A3",X"46",X"85",X"30",X"00",X"FF",X"AA",X"35",
		X"A5",X"73",X"53",X"00",X"FF",X"A3",X"45",X"5A",X"A5",X"55",X"30",X"FF",X"A4",X"51",X"55",X"55",
		X"15",X"40",X"FF",X"E4",X"64",X"58",X"58",X"46",X"4E",X"FF",X"D4",X"6A",X"58",X"59",X"46",X"4D",
		X"FF",X"D3",X"6A",X"58",X"59",X"46",X"4D",X"FF",X"C3",X"5A",X"57",X"58",X"46",X"4C",X"FF",X"0A",
		X"45",X"57",X"57",X"66",X"00",X"FF",X"00",X"34",X"56",X"46",X"60",X"00",X"FF",X"00",X"0A",X"45",
		X"35",X"00",X"00",X"FF",X"00",X"00",X"00",X"33",X"34",X"43",X"FF",X"00",X"0E",X"35",X"4A",X"89",
		X"64",X"FF",X"00",X"D4",X"55",X"5A",X"88",X"74",X"FF",X"0C",X"46",X"41",X"5C",X"66",X"54",X"FF",
		X"04",X"53",X"44",X"5C",X"45",X"44",X"FF",X"A4",X"3A",X"87",X"55",X"55",X"54",X"FF",X"A4",X"A7",
		X"85",X"78",X"41",X"53",X"FF",X"A3",X"67",X"57",X"89",X"44",X"53",X"FF",X"AA",X"55",X"68",X"83",
		X"56",X"3E",X"FF",X"0A",X"35",X"67",X"35",X"63",X"E0",X"FF",X"0A",X"A3",X"65",X"55",X"3D",X"00",
		X"FF",X"00",X"AA",X"33",X"A3",X"C0",X"00",X"FF",X"00",X"0A",X"AA",X"AA",X"00",X"00",X"FF",X"00",
		X"00",X"ED",X"C0",X"00",X"FF",X"00",X"05",X"33",X"30",X"00",X"FF",X"00",X"55",X"66",X"65",X"00",
		X"FF",X"05",X"51",X"44",X"44",X"50",X"FF",X"03",X"55",X"67",X"88",X"70",X"FF",X"04",X"35",X"67",
		X"99",X"85",X"FF",X"36",X"7A",X"55",X"55",X"55",X"FF",X"36",X"6A",X"58",X"98",X"86",X"FF",X"04",
		X"A3",X"55",X"56",X"66",X"FF",X"AA",X"43",X"55",X"56",X"6A",X"FF",X"A3",X"41",X"4A",X"AA",X"50",
		X"FF",X"AA",X"33",X"55",X"55",X"A0",X"FF",X"0A",X"A3",X"33",X"3A",X"00",X"FF",X"00",X"AA",X"ED",
		X"CA",X"00",X"FF",X"00",X"00",X"ED",X"C0",X"00",X"FF",X"00",X"05",X"33",X"30",X"00",X"FF",X"00",
		X"55",X"66",X"65",X"00",X"FF",X"05",X"51",X"44",X"44",X"50",X"FF",X"03",X"55",X"67",X"88",X"70",
		X"FF",X"A3",X"35",X"67",X"99",X"85",X"FF",X"AA",X"3A",X"55",X"55",X"55",X"FF",X"0A",X"3A",X"58",
		X"98",X"86",X"FF",X"00",X"A3",X"55",X"56",X"66",X"FF",X"03",X"43",X"55",X"56",X"6A",X"FF",X"03",
		X"41",X"4A",X"AA",X"50",X"FF",X"AA",X"33",X"55",X"55",X"A0",X"FF",X"AA",X"A3",X"33",X"3A",X"00",
		X"FF",X"00",X"AA",X"ED",X"CA",X"00",X"FF",X"00",X"00",X"00",X"ED",X"C0",X"00",X"FF",X"00",X"00",
		X"05",X"33",X"30",X"00",X"FF",X"00",X"00",X"55",X"66",X"65",X"00",X"FF",X"00",X"05",X"51",X"44",
		X"44",X"50",X"FF",X"00",X"03",X"55",X"67",X"88",X"70",X"FF",X"00",X"A3",X"35",X"67",X"99",X"85",
		X"FF",X"00",X"BB",X"1A",X"55",X"55",X"55",X"FF",X"BB",X"B1",X"2A",X"58",X"98",X"86",X"FF",X"00",
		X"BB",X"33",X"55",X"56",X"66",X"FF",X"00",X"03",X"43",X"55",X"56",X"6A",X"FF",X"00",X"03",X"41",
		X"4A",X"AA",X"50",X"FF",X"00",X"AA",X"33",X"55",X"55",X"A0",X"FF",X"00",X"AA",X"A3",X"33",X"3A",
		X"00",X"FF",X"00",X"00",X"AA",X"ED",X"CA",X"00",X"FF",X"00",X"AA",X"00",X"A0",X"00",X"00",X"FF",
		X"0A",X"A3",X"A3",X"3A",X"30",X"00",X"FF",X"AA",X"35",X"37",X"73",X"53",X"00",X"FF",X"A3",X"45",
		X"5A",X"A5",X"55",X"30",X"FF",X"A4",X"51",X"55",X"55",X"15",X"50",X"FF",X"E4",X"64",X"57",X"58",
		X"46",X"4E",X"FF",X"D4",X"6A",X"58",X"59",X"46",X"4D",X"FF",X"D3",X"6A",X"58",X"59",X"46",X"4D",
		X"FF",X"C3",X"5A",X"57",X"58",X"46",X"4C",X"FF",X"0A",X"45",X"57",X"57",X"66",X"00",X"FF",X"00",
		X"34",X"56",X"56",X"50",X"00",X"FF",X"00",X"03",X"45",X"45",X"00",X"00",X"FF",X"00",X"A0",X"00",
		X"0A",X"00",X"00",X"FF",X"0A",X"AA",X"00",X"AA",X"30",X"00",X"FF",X"AA",X"35",X"AA",X"A3",X"53",
		X"00",X"FF",X"A3",X"45",X"5A",X"A5",X"55",X"30",X"FF",X"A4",X"51",X"55",X"55",X"15",X"50",X"FF",
		X"E4",X"64",X"57",X"58",X"46",X"4E",X"FF",X"D4",X"6A",X"58",X"59",X"46",X"4D",X"FF",X"D3",X"6A",
		X"58",X"59",X"46",X"4D",X"FF",X"C3",X"5A",X"57",X"58",X"46",X"4C",X"FF",X"0A",X"45",X"57",X"57",
		X"66",X"00",X"FF",X"00",X"34",X"56",X"56",X"50",X"00",X"FF",X"00",X"03",X"45",X"45",X"00",X"00",
		X"FF",X"00",X"00",X"0B",X"00",X"00",X"00",X"FF",X"00",X"00",X"0B",X"B0",X"00",X"00",X"FF",X"00",
		X"A0",X"B1",X"1B",X"00",X"00",X"FF",X"0A",X"A3",X"11",X"11",X"30",X"00",X"FF",X"AA",X"35",X"32",
		X"23",X"53",X"00",X"FF",X"A3",X"45",X"5A",X"A5",X"55",X"30",X"FF",X"A4",X"51",X"55",X"55",X"15",
		X"40",X"FF",X"E4",X"64",X"69",X"58",X"46",X"4E",X"FF",X"D4",X"6A",X"69",X"59",X"46",X"4D",X"FF",
		X"D3",X"6A",X"68",X"59",X"46",X"4D",X"FF",X"C3",X"5A",X"68",X"58",X"46",X"4C",X"FF",X"AA",X"45",
		X"67",X"57",X"65",X"00",X"FF",X"0A",X"34",X"56",X"56",X"50",X"00",X"FF",X"00",X"A3",X"45",X"45",
		X"00",X"00",X"FF",X"00",X"00",X"03",X"33",X"00",X"00",X"FF",X"00",X"0E",X"35",X"4A",X"33",X"30",
		X"FF",X"00",X"D4",X"55",X"5A",X"69",X"30",X"FF",X"0C",X"46",X"41",X"5C",X"67",X"30",X"FF",X"04",
		X"53",X"44",X"5C",X"45",X"44",X"FF",X"A3",X"3A",X"87",X"55",X"55",X"54",X"FF",X"A3",X"A8",X"86",
		X"58",X"41",X"53",X"FF",X"A3",X"67",X"65",X"89",X"44",X"53",X"FF",X"AA",X"55",X"57",X"83",X"65",
		X"3E",X"FF",X"0A",X"35",X"67",X"36",X"53",X"E0",X"FF",X"0A",X"A3",X"65",X"55",X"3D",X"00",X"FF",
		X"00",X"AA",X"33",X"A3",X"C0",X"00",X"FF",X"00",X"0A",X"AA",X"AA",X"00",X"00",X"FF",X"00",X"00",
		X"03",X"33",X"00",X"00",X"FF",X"00",X"0E",X"35",X"4A",X"00",X"00",X"FF",X"00",X"D4",X"55",X"5A",
		X"40",X"00",X"FF",X"0C",X"46",X"41",X"5C",X"74",X"00",X"FF",X"04",X"53",X"44",X"5C",X"45",X"44",
		X"FF",X"A3",X"3A",X"87",X"55",X"55",X"54",X"FF",X"A3",X"A8",X"85",X"78",X"41",X"53",X"FF",X"A3",
		X"67",X"57",X"89",X"44",X"53",X"FF",X"AA",X"55",X"68",X"93",X"65",X"3E",X"FF",X"0A",X"35",X"69",
		X"36",X"53",X"E0",X"FF",X"0A",X"A3",X"65",X"55",X"3D",X"00",X"FF",X"00",X"AA",X"33",X"A3",X"C0",
		X"00",X"FF",X"00",X"0A",X"AA",X"AA",X"00",X"00",X"FF",X"00",X"0A",X"AA",X"00",X"00",X"BB",X"FF",
		X"00",X"AA",X"33",X"30",X"BB",X"B0",X"FF",X"0A",X"E3",X"54",X"AB",X"11",X"B0",X"FF",X"AD",X"45",
		X"55",X"A2",X"21",X"B0",X"FF",X"C4",X"64",X"15",X"32",X"2B",X"00",X"FF",X"45",X"34",X"45",X"C4",
		X"54",X"40",X"FF",X"33",X"A8",X"75",X"55",X"55",X"40",X"FF",X"3A",X"88",X"57",X"84",X"15",X"30",
		X"FF",X"36",X"75",X"78",X"94",X"45",X"30",X"FF",X"A5",X"56",X"89",X"36",X"53",X"E0",X"FF",X"A3",
		X"56",X"93",X"65",X"3E",X"00",X"FF",X"0A",X"36",X"55",X"53",X"D0",X"00",X"FF",X"00",X"03",X"3A",
		X"3C",X"00",X"00",X"FF",X"00",X"0A",X"00",X"FF",X"00",X"5A",X"A0",X"FF",X"05",X"AB",X"AA",X"FF",
		X"05",X"BC",X"DB",X"FF",X"00",X"AB",X"A0",X"FF",X"00",X"0A",X"00",X"FF",X"00",X"0C",X"00",X"FF",
		X"00",X"DB",X"A0",X"FF",X"0C",X"BA",X"AB",X"FF",X"0A",X"AA",X"BC",X"FF",X"00",X"BB",X"C0",X"FF",
		X"00",X"0B",X"00",X"FF",X"00",X"0B",X"00",X"FF",X"00",X"AB",X"A0",X"FF",X"0A",X"DC",X"BA",X"FF",
		X"0A",X"BB",X"A5",X"FF",X"00",X"AA",X"50",X"FF",X"00",X"05",X"00",X"FF",X"00",X"0A",X"00",X"FF",
		X"00",X"AB",X"B0",X"FF",X"0A",X"BB",X"AA",X"FF",X"0A",X"BB",X"AA",X"FF",X"00",X"AA",X"A0",X"FF",
		X"00",X"0A",X"00",X"FF",X"08",X"88",X"77",X"67",X"78",X"00",X"FF",X"98",X"81",X"62",X"6A",X"69",
		X"00",X"FF",X"99",X"89",X"86",X"69",X"80",X"00",X"FF",X"99",X"88",X"55",X"35",X"68",X"3B",X"FF",
		X"09",X"96",X"66",X"56",X"76",X"76",X"FF",X"09",X"8E",X"ED",X"DC",X"C9",X"88",X"FF",X"09",X"8E",
		X"ED",X"DC",X"C9",X"88",X"FF",X"09",X"96",X"66",X"56",X"78",X"86",X"FF",X"09",X"88",X"55",X"36",
		X"68",X"3B",X"FF",X"09",X"89",X"86",X"69",X"80",X"00",X"FF",X"98",X"81",X"62",X"6A",X"69",X"00",
		X"FF",X"98",X"87",X"76",X"67",X"88",X"00",X"FF",X"99",X"99",X"99",X"99",X"00",X"00",X"FF",X"00",
		X"40",X"B8",X"8B",X"04",X"00",X"FF",X"00",X"05",X"87",X"78",X"50",X"00",X"FF",X"06",X"88",X"89",
		X"98",X"88",X"60",X"FF",X"98",X"A6",X"7C",X"C7",X"6A",X"80",X"FF",X"97",X"75",X"6C",X"C7",X"57",
		X"70",X"FF",X"96",X"64",X"5C",X"C4",X"34",X"60",X"FF",X"97",X"15",X"6D",X"D6",X"31",X"70",X"FF",
		X"97",X"66",X"7D",X"D7",X"56",X"70",X"FF",X"97",X"77",X"7D",X"D7",X"67",X"70",X"FF",X"97",X"27",
		X"7E",X"E7",X"62",X"70",X"FF",X"98",X"77",X"7E",X"E7",X"77",X"80",X"FF",X"98",X"88",X"98",X"89",
		X"88",X"80",X"FF",X"98",X"88",X"99",X"99",X"88",X"80",X"FF",X"99",X"90",X"00",X"09",X"99",X"00",
		X"FF",X"00",X"00",X"00",X"88",X"80",X"B6",X"00",X"FF",X"00",X"00",X"07",X"7A",X"88",X"48",X"80",
		X"FF",X"00",X"00",X"76",X"56",X"69",X"77",X"86",X"FF",X"00",X"07",X"62",X"44",X"7C",X"97",X"4B",
		X"FF",X"00",X"87",X"65",X"47",X"CC",X"C9",X"80",X"FF",X"08",X"81",X"66",X"7C",X"C6",X"55",X"78",
		X"FF",X"08",X"88",X"68",X"DD",X"64",X"3A",X"68",X"FF",X"98",X"88",X"8E",X"D6",X"53",X"45",X"78",
		X"FF",X"99",X"89",X"8E",X"76",X"62",X"55",X"79",X"FF",X"09",X"99",X"98",X"76",X"66",X"67",X"90",
		X"FF",X"00",X"00",X"09",X"71",X"77",X"79",X"00",X"FF",X"00",X"00",X"08",X"88",X"88",X"90",X"00",
		X"FF",X"00",X"00",X"08",X"88",X"89",X"00",X"00",X"FF",X"00",X"00",X"09",X"88",X"90",X"00",X"00",
		X"FF",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"FF",X"FF",X"00",X"AB",X"B0",X"FF",X"0A",X"BB",
		X"AA",X"FF",X"0A",X"BB",X"AA",X"FF",X"00",X"AA",X"A0",X"FF",X"00",X"0A",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"76",X"67",X"00",X"FF",X"00",X"00",
		X"00",X"27",X"65",X"55",X"70",X"FF",X"00",X"00",X"00",X"02",X"72",X"54",X"EE",X"FF",X"00",X"02",
		X"33",X"27",X"AA",X"24",X"57",X"FF",X"03",X"3E",X"EE",X"EA",X"99",X"A7",X"45",X"FF",X"23",X"EE",
		X"11",X"E9",X"88",X"92",X"44",X"FF",X"03",X"3E",X"EE",X"EA",X"99",X"A2",X"44",X"FF",X"0C",X"C2",
		X"33",X"27",X"AA",X"77",X"47",X"FF",X"00",X"00",X"CC",X"C2",X"66",X"54",X"EE",X"FF",X"00",X"00",
		X"00",X"27",X"65",X"44",X"70",X"FF",X"00",X"00",X"00",X"00",X"77",X"77",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"77",X"77",X"00",X"FF",X"00",X"00",X"33",X"27",X"65",X"56",X"70",X"FF",X"00",X"02",
		X"EE",X"32",X"62",X"54",X"11",X"FF",X"00",X"03",X"E1",X"E6",X"AA",X"24",X"57",X"FF",X"00",X"3E",
		X"11",X"EA",X"99",X"A6",X"45",X"FF",X"00",X"21",X"11",X"E9",X"88",X"92",X"44",X"FF",X"00",X"3E",
		X"11",X"EA",X"99",X"A2",X"44",X"FF",X"00",X"03",X"11",X"E6",X"AA",X"66",X"46",X"FF",X"00",X"02",
		X"EE",X"32",X"66",X"64",X"11",X"FF",X"00",X"00",X"33",X"27",X"66",X"54",X"60",X"FF",X"00",X"00",
		X"0C",X"CC",X"77",X"77",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"77",X"77",X"00",X"FF",X"00",X"00",
		X"03",X"27",X"65",X"56",X"70",X"FF",X"00",X"00",X"2E",X"32",X"62",X"54",X"EE",X"FF",X"00",X"00",
		X"31",X"E6",X"AA",X"24",X"57",X"FF",X"00",X"03",X"E1",X"EA",X"99",X"A6",X"45",X"FF",X"00",X"02",
		X"E1",X"E9",X"88",X"92",X"44",X"FF",X"00",X"03",X"E1",X"EA",X"99",X"A2",X"44",X"FF",X"00",X"00",
		X"31",X"E6",X"AA",X"66",X"46",X"FF",X"00",X"00",X"2E",X"32",X"66",X"64",X"EE",X"FF",X"00",X"00",
		X"03",X"27",X"66",X"54",X"60",X"FF",X"00",X"00",X"00",X"CC",X"77",X"77",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"0E",X"64",X"6E",X"00",X"FF",X"00",X"6E",X"44",X"4E",
		X"60",X"FF",X"06",X"44",X"72",X"64",X"47",X"FF",X"07",X"45",X"A9",X"A5",X"47",X"FF",X"07",X"5A",
		X"98",X"9A",X"57",X"FF",X"07",X"6A",X"98",X"9A",X"67",X"FF",X"06",X"67",X"A9",X"A7",X"66",X"FF",
		X"02",X"26",X"EA",X"E6",X"22",X"FF",X"02",X"03",X"EE",X"E3",X"02",X"FF",X"00",X"03",X"E1",X"E3",
		X"00",X"FF",X"00",X"03",X"E1",X"E3",X"00",X"FF",X"00",X"02",X"E1",X"E2",X"00",X"FF",X"00",X"00",
		X"3E",X"30",X"00",X"FF",X"00",X"00",X"3E",X"30",X"00",X"FF",X"00",X"00",X"02",X"00",X"00",X"FF",
		X"00",X"01",X"64",X"51",X"00",X"FF",X"00",X"61",X"44",X"41",X"60",X"FF",X"06",X"44",X"72",X"64",
		X"47",X"FF",X"07",X"45",X"A9",X"A5",X"47",X"FF",X"07",X"5A",X"98",X"9A",X"57",X"FF",X"07",X"6A",
		X"98",X"9A",X"67",X"FF",X"06",X"67",X"A9",X"A7",X"66",X"FF",X"02",X"27",X"3A",X"36",X"22",X"FF",
		X"02",X"03",X"EE",X"E3",X"02",X"FF",X"00",X"3E",X"11",X"1E",X"30",X"FF",X"00",X"23",X"E1",X"E3",
		X"20",X"FF",X"00",X"02",X"3E",X"32",X"00",X"FF",X"00",X"00",X"32",X"30",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"0E",X"64",X"6E",X"00",X"FF",
		X"00",X"6E",X"44",X"4E",X"60",X"FF",X"06",X"44",X"72",X"64",X"47",X"FF",X"07",X"45",X"A9",X"A5",
		X"47",X"FF",X"07",X"5A",X"98",X"9A",X"57",X"FF",X"07",X"6A",X"98",X"9A",X"67",X"FF",X"06",X"67",
		X"A9",X"A7",X"66",X"FF",X"02",X"27",X"3A",X"36",X"22",X"FF",X"02",X"33",X"EE",X"E3",X"32",X"FF",
		X"00",X"31",X"11",X"11",X"30",X"FF",X"00",X"23",X"EE",X"E3",X"20",X"FF",X"00",X"02",X"32",X"32",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"06",X"66",X"E6",X"00",X"FF",X"00",X"00",X"65",X"5E",X"55",
		X"60",X"FF",X"00",X"06",X"65",X"56",X"44",X"56",X"FF",X"00",X"07",X"7A",X"99",X"64",X"4E",X"FF",
		X"00",X"22",X"A9",X"98",X"95",X"E6",X"FF",X"00",X"07",X"A9",X"89",X"96",X"56",X"FF",X"00",X"03",
		X"E9",X"99",X"A5",X"56",X"FF",X"00",X"3E",X"EE",X"AA",X"76",X"67",X"FF",X"03",X"E1",X"EE",X"3C",
		X"77",X"70",X"FF",X"2E",X"11",X"E3",X"C0",X"27",X"00",X"FF",X"3E",X"1E",X"3C",X"00",X"00",X"00",
		X"FF",X"3E",X"E2",X"00",X"00",X"00",X"00",X"FF",X"23",X"30",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"06",X"66",X"16",X"00",X"FF",X"00",X"00",X"65",X"51",X"E5",X"60",X"FF",X"00",X"06",X"65",
		X"56",X"44",X"56",X"FF",X"00",X"07",X"7A",X"A9",X"64",X"E1",X"FF",X"00",X"22",X"A9",X"98",X"95",
		X"16",X"FF",X"00",X"07",X"A9",X"89",X"A6",X"56",X"FF",X"00",X"C3",X"E9",X"99",X"A5",X"56",X"FF",
		X"00",X"3E",X"1E",X"AA",X"76",X"67",X"FF",X"00",X"31",X"11",X"33",X"77",X"70",X"FF",X"00",X"3E",
		X"1E",X"30",X"27",X"00",X"FF",X"00",X"C3",X"3C",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"06",X"66",X"E6",X"00",
		X"FF",X"00",X"00",X"65",X"5E",X"55",X"60",X"FF",X"00",X"06",X"65",X"56",X"44",X"56",X"FF",X"00",
		X"07",X"7A",X"A9",X"64",X"5E",X"FF",X"00",X"22",X"A9",X"98",X"95",X"E6",X"FF",X"00",X"07",X"A9",
		X"89",X"A6",X"56",X"FF",X"00",X"23",X"E9",X"99",X"A5",X"56",X"FF",X"00",X"31",X"1E",X"AA",X"76",
		X"67",X"FF",X"00",X"3E",X"11",X"33",X"77",X"70",X"FF",X"00",X"02",X"E1",X"30",X"27",X"00",X"FF",
		X"00",X"00",X"33",X"20",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"0E",X"E0",X"FF",X"EB",X"CE",X"FF",X"EC",X"BE",X"FF",X"0E",X"E0",
		X"FF",X"0E",X"EE",X"00",X"FF",X"EB",X"CB",X"E0",X"FF",X"EC",X"8C",X"E0",X"FF",X"EB",X"CB",X"E0",
		X"FF",X"0E",X"EE",X"00",X"FF",X"00",X"DD",X"D0",X"00",X"FF",X"0D",X"CB",X"BD",X"00",X"FF",X"EC",
		X"9A",X"8B",X"D0",X"FF",X"EC",X"A1",X"AB",X"D0",X"FF",X"EC",X"8A",X"9C",X"D0",X"FF",X"0E",X"CC",
		X"CE",X"00",X"FF",X"00",X"EE",X"E0",X"00",X"FF",X"11",X"FF",X"11",X"FF",X"11",X"FF",X"22",X"44",
		X"FF",X"77",X"77",X"FF",X"22",X"44",X"FF",X"44",X"66",X"88",X"FF",X"77",X"77",X"77",X"FF",X"44",
		X"66",X"88",X"FF",X"66",X"88",X"AA",X"CC",X"FF",X"77",X"77",X"77",X"77",X"FF",X"66",X"88",X"AA",
		X"CC",X"FF",X"88",X"AA",X"CC",X"EE",X"11",X"FF",X"87",X"77",X"77",X"77",X"77",X"FF",X"88",X"AA",
		X"CC",X"EE",X"11",X"FF",X"AA",X"CC",X"EE",X"11",X"22",X"44",X"FF",X"77",X"77",X"77",X"77",X"77",
		X"77",X"FF",X"AA",X"CC",X"EE",X"11",X"22",X"44",X"FF",X"CC",X"EE",X"11",X"22",X"44",X"66",X"88",
		X"FF",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"FF",X"CC",X"EE",X"11",X"22",X"44",X"66",X"88",
		X"FF",X"EE",X"11",X"22",X"44",X"66",X"88",X"AA",X"CC",X"FF",X"77",X"77",X"77",X"77",X"77",X"77",
		X"77",X"77",X"FF",X"EE",X"11",X"22",X"44",X"66",X"88",X"AA",X"CC",X"FF",X"11",X"10",X"FF",X"11",
		X"10",X"FF",X"27",X"20",X"FF",X"27",X"20",X"FF",X"47",X"40",X"FF",X"47",X"40",X"FF",X"47",X"40",
		X"FF",X"47",X"40",X"FF",X"67",X"60",X"FF",X"67",X"60",X"FF",X"87",X"80",X"FF",X"87",X"80",X"FF",
		X"67",X"60",X"FF",X"67",X"60",X"FF",X"87",X"80",X"FF",X"87",X"80",X"FF",X"A7",X"A0",X"FF",X"A7",
		X"A0",X"FF",X"C7",X"C0",X"FF",X"C7",X"C0",X"FF",X"88",X"80",X"FF",X"87",X"80",X"FF",X"A7",X"A0",
		X"FF",X"A7",X"A0",X"FF",X"C7",X"C0",X"FF",X"C7",X"C0",X"FF",X"E7",X"E0",X"FF",X"E7",X"E0",X"FF",
		X"17",X"10",X"FF",X"17",X"10",X"FF",X"A7",X"A0",X"FF",X"A7",X"A0",X"FF",X"C7",X"C0",X"FF",X"C7",
		X"C0",X"FF",X"E7",X"E0",X"FF",X"E7",X"E0",X"FF",X"17",X"10",X"FF",X"17",X"10",X"FF",X"27",X"20",
		X"FF",X"27",X"20",X"FF",X"47",X"40",X"FF",X"47",X"40",X"FF",X"C7",X"C0",X"FF",X"C7",X"C0",X"FF",
		X"E7",X"E0",X"FF",X"E7",X"E0",X"FF",X"17",X"10",X"FF",X"17",X"10",X"FF",X"27",X"20",X"FF",X"27",
		X"20",X"FF",X"47",X"40",X"FF",X"47",X"40",X"FF",X"67",X"60",X"FF",X"67",X"60",X"FF",X"87",X"80",
		X"FF",X"87",X"80",X"FF",X"E7",X"E0",X"FF",X"E7",X"E0",X"FF",X"17",X"10",X"FF",X"17",X"10",X"FF",
		X"27",X"20",X"FF",X"27",X"20",X"FF",X"47",X"40",X"FF",X"47",X"40",X"FF",X"67",X"60",X"FF",X"67",
		X"60",X"FF",X"87",X"80",X"FF",X"87",X"80",X"FF",X"A7",X"A0",X"FF",X"A7",X"A0",X"FF",X"C7",X"C0",
		X"FF",X"C7",X"C0",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"9A",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"0A",X"9A",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"0A",X"89",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"08",X"AA",X"A0",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"0A",X"A9",X"A0",X"00",X"00",X"00",X"FF",X"00",X"00",X"EE",X"88",X"A0",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"0A",X"A9",X"88",X"00",X"CC",X"00",X"FF",X"00",X"00",X"0A",
		X"9A",X"AA",X"00",X"C0",X"00",X"FF",X"00",X"00",X"0A",X"99",X"AA",X"DD",X"D0",X"00",X"FF",X"00",
		X"00",X"0A",X"99",X"AA",X"DD",X"DC",X"00",X"FF",X"00",X"B4",X"DB",X"89",X"9A",X"A0",X"00",X"00",
		X"FF",X"CB",X"BA",X"CB",X"88",X"99",X"9A",X"AA",X"BB",X"FF",X"DD",X"BC",X"DD",X"CC",X"CC",X"CB",
		X"BB",X"BC",X"FF",X"00",X"C4",X"DD",X"CC",X"BB",X"C0",X"00",X"00",X"FF",X"00",X"00",X"0D",X"CB",
		X"BB",X"DD",X"DC",X"00",X"FF",X"00",X"00",X"0C",X"BB",X"BB",X"DD",X"D0",X"00",X"FF",X"00",X"00",
		X"0B",X"BA",X"AB",X"00",X"C0",X"00",X"FF",X"00",X"00",X"0B",X"AA",X"AA",X"00",X"CC",X"00",X"FF",
		X"00",X"00",X"EE",X"BB",X"C0",X"00",X"00",X"00",X"FF",X"00",X"00",X"0C",X"AB",X"B0",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"0B",X"CA",X"B0",X"00",X"00",X"00",X"FF",X"00",X"00",X"0B",X"BC",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"0C",X"BB",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"CB",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"AA",X"A0",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"AA",X"AA",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"09",X"99",X"AA",X"00",X"00",X"00",X"FF",X"00",X"00",X"09",X"99",X"99",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"DD",X"BB",X"BB",X"00",X"CC",X"00",X"FF",X"00",X"00",X"0B",X"BB",
		X"BB",X"BD",X"D0",X"00",X"FF",X"00",X"00",X"0B",X"BB",X"BB",X"BD",X"DC",X"0A",X"FF",X"00",X"BD",
		X"DB",X"AA",X"AB",X"BB",X"0A",X"AB",X"FF",X"CB",X"BA",X"CA",X"99",X"AA",X"AA",X"AB",X"B0",X"FF",
		X"CC",X"CB",X"DC",X"CC",X"CC",X"BB",X"BC",X"00",X"FF",X"00",X"CD",X"DC",X"BB",X"BB",X"BB",X"00",
		X"00",X"FF",X"00",X"00",X"0C",X"BA",X"AA",X"BD",X"DC",X"00",X"FF",X"00",X"00",X"0C",X"AA",X"AA",
		X"BD",X"D0",X"00",X"FF",X"00",X"00",X"DD",X"CC",X"CC",X"00",X"CC",X"00",X"FF",X"00",X"00",X"0C",
		X"CC",X"BB",X"00",X"00",X"00",X"FF",X"00",X"00",X"0B",X"BB",X"BB",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"BB",X"BB",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"BB",X"B0",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"BB",X"A0",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"0E",X"ED",X"CA",X"00",X"00",X"00",X"FF",X"00",X"00",X"0D",X"DD",
		X"DC",X"00",X"CC",X"00",X"FF",X"00",X"00",X"EE",X"DD",X"DD",X"CD",X"DC",X"00",X"FF",X"00",X"00",
		X"0D",X"DD",X"CC",X"CD",X"D0",X"00",X"FF",X"00",X"B4",X"DD",X"CB",X"BB",X"CC",X"00",X"00",X"FF",
		X"CB",X"BA",X"CC",X"A9",X"AA",X"AB",X"BB",X"BB",X"FF",X"CC",X"CB",X"DE",X"DD",X"DD",X"CC",X"CC",
		X"CC",X"FF",X"00",X"C4",X"DD",X"DD",X"DC",X"CC",X"00",X"00",X"FF",X"00",X"00",X"0D",X"CC",X"CC",
		X"CD",X"D0",X"00",X"FF",X"00",X"00",X"EE",X"CC",X"BB",X"BD",X"DC",X"00",X"FF",X"00",X"00",X"0B",
		X"BB",X"BB",X"00",X"CC",X"00",X"FF",X"00",X"00",X"0A",X"BB",X"BA",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"AA",X"A0",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"AA",X"A0",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"AA",X"9A",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"0A",X"99",X"AA",X"00",X"00",X"00",X"FF",X"00",X"00",X"0A",X"9A",
		X"A9",X"00",X"00",X"00",X"FF",X"00",X"00",X"DD",X"BA",X"99",X"00",X"CC",X"00",X"FF",X"00",X"00",
		X"0B",X"AA",X"AA",X"BD",X"D0",X"00",X"FF",X"00",X"00",X"0B",X"A8",X"AA",X"BD",X"DC",X"00",X"FF",
		X"00",X"BE",X"DB",X"A8",X"8A",X"AB",X"00",X"00",X"FF",X"CB",X"BA",X"CA",X"88",X"88",X"AA",X"AB",
		X"00",X"FF",X"CC",X"CB",X"DD",X"CC",X"CC",X"CC",X"CA",X"A0",X"FF",X"00",X"CE",X"DD",X"CC",X"CB",
		X"BC",X"00",X"BA",X"FF",X"00",X"00",X"0D",X"CB",X"BB",X"CD",X"DC",X"00",X"FF",X"00",X"00",X"0D",
		X"CB",X"BC",X"CD",X"D0",X"00",X"FF",X"00",X"00",X"EE",X"CC",X"BB",X"00",X"CC",X"00",X"FF",X"00",
		X"00",X"0D",X"DB",X"BB",X"00",X"00",X"00",X"FF",X"00",X"00",X"0D",X"CD",X"CC",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"DC",X"DD",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"DC",X"C0",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"BA",
		X"A0",X"00",X"00",X"00",X"FF",X"00",X"00",X"0B",X"AA",X"9A",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"0B",X"A9",X"AA",X"00",X"CC",X"00",X"FF",X"00",X"00",X"EE",X"89",X"99",X"9D",X"DC",X"00",X"FF",
		X"00",X"00",X"0C",X"A9",X"AA",X"BD",X"E0",X"00",X"FF",X"00",X"B4",X"DC",X"B8",X"89",X"AB",X"00",
		X"00",X"FF",X"CB",X"BA",X"CB",X"A8",X"88",X"9A",X"AA",X"AA",X"FF",X"CC",X"CB",X"DE",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"FF",X"00",X"C4",X"DD",X"CC",X"CC",X"CC",X"00",X"00",X"FF",X"00",X"00",X"0D",
		X"CC",X"CC",X"CD",X"D0",X"00",X"FF",X"00",X"00",X"EE",X"BC",X"BB",X"BD",X"DC",X"00",X"FF",X"00",
		X"00",X"0D",X"CB",X"CC",X"00",X"CC",X"00",X"FF",X"00",X"00",X"0D",X"DC",X"BC",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"DD",X"D0",X"00",X"00",X"00",X"FF",X"08",X"80",X"FF",X"08",X"80",X"FF",
		X"08",X"80",X"FF",X"08",X"80",X"FF",X"00",X"90",X"FF",X"09",X"99",X"FF",X"99",X"90",X"FF",X"09",
		X"00",X"FF",X"00",X"00",X"FF",X"88",X"88",X"FF",X"88",X"88",X"FF",X"00",X"00",X"FF",X"08",X"00",
		X"FF",X"88",X"80",X"FF",X"08",X"88",X"FF",X"00",X"80",X"FF",X"09",X"00",X"07",X"00",X"09",X"00",
		X"FF",X"00",X"90",X"65",X"50",X"90",X"00",X"FF",X"09",X"08",X"65",X"58",X"09",X"00",X"FF",X"00",
		X"06",X"54",X"56",X"00",X"00",X"FF",X"0E",X"EE",X"52",X"5E",X"EE",X"00",X"FF",X"B1",X"91",X"65",
		X"61",X"91",X"E0",X"FF",X"BB",X"BB",X"B4",X"BB",X"B0",X"00",X"FF",X"00",X"CB",X"62",X"50",X"00",
		X"00",X"FF",X"0B",X"4B",X"69",X"40",X"00",X"00",X"FF",X"00",X"BB",X"49",X"40",X"C0",X"00",X"FF",
		X"00",X"0B",X"63",X"5B",X"40",X"00",X"FF",X"00",X"00",X"B3",X"0B",X"00",X"00",X"FF",X"00",X"00",
		X"BC",X"00",X"00",X"00",X"FF",X"00",X"00",X"BC",X"00",X"00",X"00",X"FF",X"00",X"00",X"B3",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"0B",X"30",X"00",X"00",X"FF",X"01",X"00",X"07",X"00",X"01",X"00",
		X"FF",X"00",X"10",X"65",X"50",X"10",X"00",X"FF",X"01",X"0B",X"65",X"5B",X"01",X"00",X"FF",X"00",
		X"06",X"54",X"56",X"00",X"00",X"FF",X"0E",X"EE",X"52",X"5E",X"EE",X"00",X"FF",X"B1",X"91",X"E5",
		X"E1",X"91",X"E0",X"FF",X"BB",X"BB",X"B4",X"BB",X"B0",X"00",X"FF",X"00",X"0B",X"62",X"60",X"C0",
		X"00",X"FF",X"00",X"0B",X"69",X"4B",X"40",X"00",X"FF",X"00",X"CB",X"49",X"4B",X"00",X"00",X"FF",
		X"0B",X"4B",X"63",X"60",X"00",X"00",X"FF",X"00",X"BB",X"B3",X"30",X"00",X"00",X"FF",X"00",X"00",
		X"BB",X"BC",X"00",X"00",X"FF",X"00",X"0B",X"33",X"33",X"00",X"00",X"FF",X"00",X"00",X"BB",X"B0",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"01",X"01",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"FF",X"00",X"70",X"0B",X"60",X"00",X"00",
		X"00",X"FF",X"00",X"06",X"55",X"66",X"EE",X"00",X"00",X"FF",X"10",X"66",X"44",X"5E",X"E9",X"00",
		X"00",X"FF",X"01",X"B6",X"52",X"5E",X"9B",X"00",X"00",X"FF",X"10",X"66",X"5E",X"55",X"B0",X"C0",
		X"00",X"FF",X"00",X"06",X"EE",X"64",X"45",X"B4",X"00",X"FF",X"00",X"0E",X"E9",X"B5",X"99",X"5B",
		X"00",X"FF",X"00",X"0B",X"9B",X"06",X"49",X"4B",X"00",X"FF",X"00",X"00",X"B0",X"0B",X"65",X"4B",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"BB",X"B3",X"00",X"FF",X"00",X"00",X"00",X"0C",X"00",X"0B",
		X"C0",X"FF",X"00",X"00",X"00",X"0B",X"40",X"0B",X"C0",X"FF",X"00",X"00",X"00",X"00",X"B0",X"00",
		X"BC",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"B3",X"FF",X"00",X"00",X"09",X"09",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"FF",X"00",X"70",X"08",X"60",X"00",X"00",
		X"00",X"FF",X"00",X"06",X"55",X"56",X"EE",X"00",X"00",X"FF",X"90",X"66",X"44",X"5E",X"E9",X"00",
		X"00",X"FF",X"09",X"86",X"52",X"6E",X"9B",X"00",X"00",X"FF",X"90",X"66",X"5E",X"65",X"B0",X"00",
		X"00",X"FF",X"00",X"06",X"EE",X"64",X"65",X"00",X"00",X"FF",X"00",X"0E",X"E9",X"B5",X"99",X"60",
		X"00",X"FF",X"00",X"0B",X"9B",X"B5",X"59",X"4B",X"C0",X"FF",X"00",X"00",X"BB",X"CB",X"55",X"4B",
		X"B4",X"FF",X"00",X"00",X"00",X"B4",X"BB",X"33",X"3B",X"FF",X"00",X"00",X"00",X"0B",X"00",X"BB",
		X"C0",X"FF",X"00",X"00",X"00",X"00",X"B3",X"3C",X"00",X"FF",X"00",X"00",X"00",X"00",X"0B",X"B0",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"E0",X"00",X"00",X"00",
		X"00",X"FF",X"90",X"9E",X"10",X"00",X"00",X"00",X"00",X"FF",X"09",X"6E",X"90",X"00",X"0C",X"40",
		X"00",X"FF",X"08",X"6E",X"10",X"06",X"5B",X"B0",X"00",X"FF",X"06",X"55",X"E0",X"54",X"95",X"00",
		X"03",X"FF",X"75",X"42",X"45",X"49",X"94",X"1C",X"CB",X"FF",X"06",X"55",X"EB",X"64",X"56",X"BB",
		X"B0",X"FF",X"08",X"6E",X"1B",X"B6",X"6B",X"00",X"00",X"FF",X"09",X"6E",X"9B",X"0B",X"B0",X"00",
		X"00",X"FF",X"90",X"9E",X"1B",X"C4",X"00",X"00",X"00",X"FF",X"00",X"0B",X"B0",X"BB",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"FF",X"10",X"1E",X"10",X"C4",X"00",X"00",
		X"00",X"FF",X"01",X"5E",X"90",X"0B",X"B0",X"00",X"00",X"FF",X"0B",X"5E",X"10",X"06",X"50",X"03",
		X"C0",X"FF",X"05",X"55",X"E0",X"54",X"95",X"3B",X"30",X"FF",X"75",X"42",X"45",X"49",X"94",X"1B",
		X"30",X"FF",X"06",X"55",X"EB",X"64",X"56",X"BB",X"30",X"FF",X"0B",X"6E",X"1B",X"B6",X"6B",X"0B",
		X"C0",X"FF",X"01",X"6E",X"9B",X"0B",X"BC",X"4B",X"00",X"FF",X"10",X"1E",X"1B",X"00",X"0B",X"B0",
		X"00",X"FF",X"00",X"0B",X"B0",X"00",X"00",X"00",X"00",X"FF",X"00",X"0C",X"60",X"FF",X"00",X"CC",
		X"C6",X"FF",X"00",X"CC",X"BB",X"FF",X"06",X"CB",X"B0",X"FF",X"06",X"6B",X"00",X"FF",X"CC",X"B0",
		X"00",X"FF",X"00",X"6C",X"FF",X"00",X"66",X"FF",X"0C",X"CB",X"FF",X"0C",X"CB",X"FF",X"06",X"6B",
		X"FF",X"EC",X"6B",X"FF",X"EC",X"CB",X"FF",X"0C",X"CB",X"FF",X"00",X"60",X"FF",X"00",X"C0",X"FF",
		X"0B",X"66",X"66",X"A0",X"FF",X"C6",X"BB",X"BB",X"6B",X"FF",X"6C",X"CC",X"CC",X"C6",X"FF",X"CC",
		X"C6",X"6C",X"CB",X"FF",X"0E",X"CC",X"6C",X"E0",X"FF",X"00",X"EC",X"60",X"00",X"FF",X"0C",X"FF",
		X"6C",X"FF",X"6C",X"FF",X"C0",X"FF",X"B0",X"C6",X"FF",X"0E",X"EC",X"FF",X"6C",X"CB",X"FF",X"66",
		X"B6",X"FF",X"0B",X"FF",X"BB",X"FF",X"EB",X"FF",X"0E",X"FF",X"88",X"FF",X"88",X"FF",X"80",X"00",
		X"00",X"00",X"FF",X"80",X"08",X"00",X"00",X"FF",X"88",X"80",X"00",X"00",X"FF",X"88",X"00",X"00",
		X"00",X"FF",X"88",X"80",X"80",X"88",X"FF",X"88",X"80",X"80",X"88",X"FF",X"88",X"00",X"00",X"00",
		X"FF",X"88",X"80",X"00",X"00",X"FF",X"80",X"08",X"00",X"00",X"FF",X"80",X"00",X"00",X"00",X"FF",
		X"B0",X"00",X"00",X"00",X"FF",X"B0",X"00",X"0B",X"00",X"FF",X"B0",X"00",X"B0",X"00",X"FF",X"BB",
		X"0B",X"B0",X"00",X"FF",X"BB",X"BB",X"00",X"00",X"FF",X"BB",X"B0",X"00",X"00",X"FF",X"BB",X"BB",
		X"B0",X"00",X"FF",X"BB",X"BB",X"BB",X"BB",X"FF",X"BB",X"BB",X"00",X"00",X"FF",X"BB",X"B0",X"00",
		X"00",X"FF",X"BB",X"BB",X"00",X"00",X"FF",X"B0",X"0B",X"B0",X"00",X"FF",X"B0",X"00",X"0B",X"00",
		X"FF",X"B0",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"80",X"FF",X"00",X"00",X"88",X"00",X"FF",
		X"00",X"88",X"80",X"00",X"FF",X"00",X"88",X"80",X"00",X"FF",X"08",X"88",X"00",X"00",X"FF",X"08",
		X"88",X"00",X"00",X"FF",X"88",X"88",X"80",X"00",X"FF",X"88",X"88",X"80",X"00",X"FF",X"08",X"88",
		X"00",X"00",X"FF",X"08",X"88",X"00",X"00",X"FF",X"00",X"88",X"80",X"00",X"FF",X"00",X"88",X"80",
		X"00",X"FF",X"00",X"00",X"88",X"00",X"FF",X"00",X"00",X"00",X"80",X"FF",X"60",X"00",X"80",X"FF",
		X"68",X"08",X"00",X"FF",X"66",X"88",X"00",X"FF",X"68",X"88",X"00",X"FF",X"86",X"86",X"00",X"FF",
		X"86",X"86",X"00",X"FF",X"68",X"88",X"00",X"FF",X"66",X"88",X"00",X"FF",X"68",X"08",X"00",X"FF",
		X"60",X"00",X"80",X"FF",X"08",X"80",X"00",X"00",X"FF",X"08",X"80",X"00",X"00",X"FF",X"00",X"80",
		X"00",X"00",X"FF",X"08",X"00",X"00",X"80",X"FF",X"80",X"08",X"88",X"08",X"FF",X"88",X"88",X"80",
		X"00",X"FF",X"08",X"00",X"00",X"00",X"FF",X"08",X"80",X"00",X"00",X"FF",X"00",X"88",X"00",X"00",
		X"FF",X"00",X"88",X"00",X"00",X"FF",X"00",X"88",X"80",X"00",X"FF",X"08",X"08",X"80",X"00",X"FF",
		X"00",X"88",X"80",X"00",X"FF",X"08",X"88",X"00",X"00",X"FF",X"08",X"88",X"00",X"00",X"FF",X"00",
		X"80",X"00",X"00",X"FF",X"08",X"00",X"00",X"80",X"FF",X"80",X"08",X"08",X"08",X"FF",X"88",X"08",
		X"00",X"00",X"FF",X"08",X"00",X"00",X"00",X"FF",X"08",X"80",X"00",X"00",X"FF",X"00",X"88",X"00",
		X"00",X"FF",X"00",X"88",X"00",X"00",X"FF",X"08",X"00",X"80",X"00",X"FF",X"08",X"88",X"88",X"00",
		X"FF",X"00",X"88",X"88",X"00",X"FF",X"00",X"88",X"80",X"00",X"FF",X"08",X"08",X"88",X"00",X"FF",
		X"00",X"88",X"88",X"80",X"FF",X"08",X"88",X"88",X"80",X"FF",X"08",X"88",X"88",X"00",X"FF",X"00",
		X"88",X"00",X"00",X"FF",X"08",X"00",X"00",X"00",X"FF",X"80",X"80",X"80",X"00",X"FF",X"88",X"08",
		X"00",X"80",X"FF",X"08",X"00",X"00",X"00",X"FF",X"08",X"88",X"00",X"00",X"FF",X"00",X"88",X"88",
		X"00",X"FF",X"00",X"88",X"88",X"80",X"FF",X"00",X"08",X"88",X"00",X"FF",X"00",X"88",X"88",X"00",
		X"FF",X"00",X"08",X"80",X"00",X"FF",X"00",X"08",X"80",X"FF",X"00",X"00",X"00",X"FF",X"00",X"80",
		X"80",X"FF",X"00",X"00",X"80",X"FF",X"00",X"80",X"08",X"FF",X"00",X"80",X"80",X"FF",X"08",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"FF",X"80",X"08",X"00",X"FF",X"08",X"00",X"00",X"FF",X"00",X"88",
		X"00",X"FF",X"00",X"80",X"08",X"FF",X"00",X"88",X"80",X"FF",X"08",X"00",X"08",X"FF",X"00",X"00",
		X"00",X"FF",X"00",X"80",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"80",X"FF",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"80",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"80",X"80",
		X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"10",X"FF",X"11",X"11",X"FF",X"01",X"10",X"FF",X"01",
		X"10",X"FF",X"01",X"00",X"FF",X"11",X"10",X"FF",X"01",X"11",X"FF",X"11",X"10",X"FF",X"01",X"11",
		X"FF",X"00",X"10",X"FF",X"00",X"01",X"00",X"FF",X"01",X"11",X"00",X"FF",X"01",X"A1",X"11",X"FF",
		X"01",X"A1",X"10",X"FF",X"11",X"11",X"10",X"FF",X"01",X"1A",X"A1",X"FF",X"01",X"1A",X"10",X"FF",
		X"00",X"01",X"00",X"FF",X"00",X"11",X"01",X"00",X"FF",X"00",X"11",X"11",X"00",X"FF",X"01",X"1D",
		X"11",X"00",X"FF",X"11",X"1D",X"D1",X"10",X"FF",X"01",X"11",X"DD",X"11",X"FF",X"11",X"D1",X"D1",
		X"10",X"FF",X"11",X"D1",X"11",X"00",X"FF",X"01",X"DD",X"1D",X"10",X"FF",X"01",X"DD",X"11",X"00",
		X"FF",X"00",X"11",X"10",X"00",X"FF",X"00",X"00",X"01",X"00",X"FF",X"00",X"10",X"11",X"00",X"FF",
		X"00",X"11",X"B1",X"00",X"FF",X"00",X"1B",X"11",X"00",X"FF",X"01",X"1B",X"B1",X"00",X"FF",X"11",
		X"11",X"11",X"11",X"FF",X"11",X"11",X"11",X"11",X"FF",X"01",X"1B",X"B1",X"10",X"FF",X"00",X"1B",
		X"11",X"00",X"FF",X"00",X"11",X"11",X"00",X"FF",X"00",X"11",X"11",X"00",X"FF",X"00",X"10",X"01",
		X"00",X"FF",X"00",X"00",X"10",X"00",X"00",X"FF",X"00",X"01",X"10",X"01",X"00",X"FF",X"00",X"11",
		X"10",X"11",X"00",X"FF",X"01",X"11",X"11",X"11",X"00",X"FF",X"00",X"1A",X"11",X"A1",X"10",X"FF",
		X"00",X"01",X"11",X"11",X"11",X"FF",X"00",X"1A",X"1A",X"A1",X"00",X"FF",X"01",X"1A",X"11",X"A1",
		X"10",X"FF",X"1A",X"11",X"1A",X"11",X"11",X"FF",X"01",X"1A",X"11",X"A1",X"00",X"FF",X"00",X"1A",
		X"11",X"11",X"00",X"FF",X"00",X"01",X"1A",X"01",X"00",X"FF",X"00",X"00",X"11",X"00",X"00",X"FF",
		X"00",X"00",X"01",X"00",X"00",X"FF",X"00",X"00",X"00",X"01",X"00",X"00",X"FF",X"00",X"01",X"00",
		X"01",X"10",X"00",X"FF",X"00",X"01",X"10",X"11",X"D1",X"00",X"FF",X"00",X"01",X"11",X"D1",X"DD",
		X"10",X"FF",X"00",X"01",X"1D",X"11",X"D1",X"00",X"FF",X"00",X"01",X"DD",X"D1",X"10",X"00",X"FF",
		X"00",X"11",X"DD",X"11",X"10",X"00",X"FF",X"01",X"D1",X"D1",X"D1",X"D1",X"00",X"FF",X"1D",X"D1",
		X"1D",X"D1",X"DD",X"10",X"FF",X"01",X"D1",X"DD",X"D1",X"DD",X"D1",X"FF",X"00",X"11",X"DD",X"D1",
		X"DD",X"10",X"FF",X"01",X"D1",X"DD",X"D1",X"D1",X"00",X"FF",X"00",X"11",X"1D",X"D1",X"10",X"00",
		X"FF",X"00",X"01",X"D1",X"D1",X"00",X"00",X"FF",X"00",X"01",X"1D",X"11",X"00",X"00",X"FF",X"00",
		X"00",X"01",X"01",X"00",X"00",X"FF",X"43",X"FF",X"24",X"44",X"42",X"FF",X"33",X"44",X"22",X"FF",
		X"02",X"22",X"20",X"FF",X"00",X"22",X"00",X"FF",X"00",X"33",X"30",X"00",X"FF",X"04",X"55",X"43",
		X"00",X"FF",X"25",X"77",X"54",X"30",X"FF",X"33",X"44",X"42",X"21",X"FF",X"34",X"55",X"43",X"21",
		X"FF",X"23",X"44",X"32",X"10",X"FF",X"02",X"32",X"21",X"00",X"FF",X"00",X"11",X"10",X"00",X"FF",
		X"00",X"33",X"33",X"20",X"00",X"FF",X"03",X"45",X"44",X"22",X"00",X"FF",X"34",X"56",X"75",X"42",
		X"30",X"FF",X"22",X"24",X"44",X"22",X"21",X"FF",X"33",X"45",X"55",X"33",X"10",X"FF",X"13",X"34",
		X"43",X"22",X"10",X"FF",X"03",X"22",X"32",X"11",X"00",X"FF",X"00",X"11",X"21",X"10",X"00",X"FF",
		X"00",X"01",X"AA",X"AA",X"A3",X"02",X"00",X"00",X"FF",X"00",X"10",X"11",X"AA",X"01",X"22",X"00",
		X"00",X"FF",X"11",X"11",X"05",X"65",X"55",X"12",X"50",X"00",X"FF",X"44",X"40",X"53",X"33",X"33",
		X"51",X"55",X"E0",X"FF",X"55",X"05",X"33",X"34",X"43",X"35",X"12",X"50",X"FF",X"E0",X"63",X"34",
		X"55",X"75",X"42",X"11",X"20",X"FF",X"44",X"23",X"45",X"77",X"65",X"52",X"14",X"12",X"FF",X"65",
		X"21",X"22",X"44",X"42",X"21",X"6D",X"41",X"FF",X"44",X"23",X"45",X"65",X"43",X"11",X"6D",X"21",
		X"FF",X"33",X"21",X"33",X"43",X"33",X"21",X"22",X"11",X"FF",X"11",X"12",X"13",X"33",X"22",X"16",
		X"41",X"15",X"FF",X"11",X"01",X"21",X"22",X"11",X"44",X"10",X"00",X"FF",X"10",X"01",X"13",X"44",
		X"44",X"45",X"1E",X"E0",X"FF",X"00",X"00",X"14",X"44",X"41",X"11",X"40",X"00",X"FF",X"00",X"00",
		X"1A",X"0A",X"A1",X"E0",X"00",X"00",X"FF",X"00",X"01",X"99",X"99",X"91",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"01",X"11",X"11",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"18",X"88",X"88",X"10",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"11",X"E5",X"A9",X"8E",X"00",X"00",X"00",X"FF",X"0E",X"EE",
		X"EE",X"76",X"55",X"22",X"E0",X"00",X"00",X"FF",X"16",X"66",X"37",X"43",X"33",X"35",X"9E",X"EE",
		X"10",X"FF",X"15",X"53",X"64",X"34",X"54",X"43",X"59",X"99",X"10",X"FF",X"0E",X"E6",X"43",X"45",
		X"65",X"55",X"25",X"E1",X"10",X"FF",X"14",X"47",X"34",X"44",X"67",X"75",X"22",X"55",X"10",X"FF",
		X"16",X"57",X"22",X"33",X"33",X"33",X"31",X"5C",X"50",X"FF",X"14",X"46",X"22",X"44",X"67",X"65",
		X"11",X"4C",X"40",X"FF",X"13",X"36",X"12",X"45",X"55",X"33",X"22",X"44",X"E0",X"FF",X"1E",X"E6",
		X"41",X"24",X"43",X"31",X"14",X"EE",X"10",X"FF",X"15",X"52",X"54",X"12",X"33",X"11",X"4A",X"AA",
		X"10",X"FF",X"14",X"44",X"25",X"33",X"11",X"44",X"AE",X"EE",X"00",X"FF",X"1E",X"EE",X"EE",X"44",
		X"44",X"11",X"E1",X"00",X"00",X"FF",X"11",X"11",X"11",X"E4",X"BA",X"8E",X"10",X"00",X"00",X"FF",
		X"00",X"00",X"08",X"88",X"88",X"10",X"00",X"00",X"00",X"FF",X"00",X"00",X"01",X"11",X"11",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"88",X"00",X"FF",X"08",X"77",X"80",X"FF",X"87",X"55",X"78",X"FF",
		X"85",X"44",X"58",X"FF",X"85",X"44",X"58",X"FF",X"77",X"55",X"78",X"FF",X"07",X"77",X"80",X"FF",
		X"00",X"77",X"00",X"FF",X"00",X"99",X"00",X"FF",X"09",X"88",X"90",X"FF",X"98",X"77",X"89",X"FF",
		X"98",X"66",X"89",X"FF",X"98",X"77",X"89",X"FF",X"09",X"88",X"90",X"FF",X"00",X"99",X"00",X"FF",
		X"00",X"9A",X"00",X"FF",X"0A",X"88",X"90",X"FF",X"A9",X"77",X"9A",X"FF",X"A9",X"77",X"9A",X"FF",
		X"0A",X"88",X"A0",X"FF",X"00",X"AA",X"00",X"FF",X"0A",X"A0",X"FF",X"A9",X"9A",X"FF",X"A8",X"8A",
		X"FF",X"A9",X"9A",X"FF",X"0A",X"A0",X"FF",X"0A",X"A0",X"FF",X"A9",X"AA",X"FF",X"A9",X"9A",X"FF",
		X"AA",X"9A",X"FF",X"0A",X"A0",X"FF",X"05",X"50",X"FF",X"52",X"25",X"FF",X"52",X"25",X"FF",X"05",
		X"50",X"FF",X"00",X"80",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"90",X"00",
		X"08",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"80",X"00",X"00",X"FF",X"00",X"09",
		X"00",X"FF",X"00",X"66",X"00",X"FF",X"04",X"22",X"40",X"FF",X"62",X"11",X"26",X"FF",X"41",X"11",
		X"14",X"FF",X"43",X"11",X"34",X"FF",X"74",X"22",X"47",X"FF",X"05",X"44",X"50",X"FF",X"00",X"77",
		X"00",X"FF",X"00",X"A9",X"00",X"FF",X"09",X"84",X"40",X"FF",X"97",X"43",X"34",X"FF",X"94",X"33",
		X"24",X"FF",X"94",X"32",X"24",X"FF",X"A4",X"33",X"24",X"FF",X"0A",X"43",X"40",X"FF",X"00",X"AA",
		X"00",X"FF",X"00",X"9A",X"00",X"FF",X"09",X"99",X"A0",X"FF",X"99",X"95",X"6A",X"FF",X"A8",X"65",
		X"59",X"FF",X"A9",X"55",X"54",X"FF",X"A9",X"55",X"44",X"FF",X"0A",X"A4",X"40",X"FF",X"00",X"AA",
		X"00",X"FF",X"00",X"BB",X"00",X"FF",X"0B",X"AA",X"A0",X"FF",X"B3",X"3A",X"9A",X"FF",X"B3",X"3B",
		X"88",X"FF",X"BA",X"B8",X"85",X"FF",X"BA",X"98",X"75",X"FF",X"0B",X"AA",X"50",X"FF",X"00",X"BB",
		X"00",X"FF",X"00",X"77",X"00",X"FF",X"07",X"88",X"80",X"FF",X"78",X"88",X"A8",X"FF",X"78",X"81",
		X"18",X"FF",X"11",X"81",X"18",X"FF",X"11",X"88",X"87",X"FF",X"07",X"88",X"70",X"FF",X"00",X"77",
		X"00",X"FF",X"00",X"77",X"00",X"FF",X"07",X"77",X"70",X"FF",X"71",X"17",X"7A",X"FF",X"71",X"17",
		X"82",X"FF",X"77",X"77",X"71",X"FF",X"77",X"77",X"77",X"FF",X"07",X"88",X"70",X"FF",X"00",X"22",
		X"00",X"FF",X"00",X"22",X"00",X"FF",X"08",X"22",X"70",X"FF",X"77",X"77",X"72",X"FF",X"22",X"77",
		X"72",X"FF",X"22",X"72",X"27",X"FF",X"77",X"72",X"27",X"FF",X"07",X"77",X"70",X"FF",X"00",X"22",
		X"00",X"FF",X"00",X"AA",X"00",X"FF",X"03",X"33",X"30",X"FF",X"33",X"88",X"33",X"FF",X"33",X"58",
		X"33",X"FF",X"88",X"83",X"58",X"FF",X"33",X"38",X"83",X"FF",X"03",X"38",X"30",X"FF",X"00",X"58",
		X"00",X"FF",X"00",X"77",X"00",X"FF",X"02",X"92",X"20",X"FF",X"15",X"85",X"52",X"FF",X"19",X"18",
		X"55",X"FF",X"88",X"11",X"89",X"FF",X"56",X"88",X"25",X"FF",X"08",X"55",X"20",X"FF",X"00",X"11",
		X"00",X"FF",X"00",X"11",X"00",X"FF",X"09",X"33",X"90",X"FF",X"39",X"99",X"13",X"FF",X"91",X"18",
		X"13",X"FF",X"91",X"19",X"99",X"FF",X"19",X"91",X"19",X"FF",X"01",X"91",X"30",X"FF",X"00",X"39",
		X"00",X"FF",X"00",X"55",X"00",X"FF",X"02",X"42",X"20",X"FF",X"74",X"14",X"52",X"FF",X"21",X"51",
		X"74",X"FF",X"42",X"71",X"44",X"FF",X"74",X"14",X"17",X"FF",X"02",X"77",X"20",X"FF",X"00",X"44",
		X"00",X"FF",X"00",X"01",X"10",X"00",X"FF",X"00",X"04",X"40",X"00",X"FF",X"11",X"AA",X"AA",X"10",
		X"FF",X"04",X"B1",X"B4",X"A0",X"FF",X"0A",X"11",X"1A",X"A0",X"FF",X"0A",X"B1",X"BB",X"A0",X"FF",
		X"04",X"BB",X"BA",X"40",X"FF",X"10",X"A6",X"6A",X"01",X"FF",X"00",X"04",X"40",X"00",X"FF",X"00",
		X"01",X"10",X"00",X"FF",X"00",X"00",X"02",X"20",X"00",X"00",X"FF",X"00",X"00",X"07",X"70",X"00",
		X"00",X"FF",X"02",X"20",X"0A",X"A0",X"22",X"00",X"FF",X"02",X"77",X"00",X"00",X"52",X"00",X"FF",
		X"00",X"0A",X"02",X"00",X"00",X"00",X"FF",X"00",X"00",X"21",X"20",X"00",X"72",X"FF",X"00",X"00",
		X"02",X"00",X"00",X"72",X"FF",X"00",X"00",X"00",X"00",X"A0",X"00",X"FF",X"25",X"70",X"00",X"00",
		X"07",X"00",X"FF",X"25",X"50",X"00",X"00",X"00",X"52",X"FF",X"00",X"00",X"0B",X"B0",X"00",X"22",
		X"FF",X"00",X"00",X"08",X"90",X"00",X"00",X"FF",X"00",X"00",X"08",X"70",X"00",X"00",X"FF",X"00",
		X"00",X"05",X"50",X"00",X"00",X"FF",X"00",X"00",X"02",X"20",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"04",X"40",X"00",X"00",X"00",X"04",X"40",X"00",X"FF",X"00",
		X"04",X"50",X"00",X"00",X"00",X"54",X"40",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"95",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"33",X"00",X"00",X"00",X"FF",X"00",X"00",X"03",X"30",X"00",X"34",X"00",X"00",X"00",
		X"FF",X"45",X"90",X"03",X"40",X"00",X"00",X"00",X"09",X"54",X"FF",X"45",X"90",X"00",X"00",X"00",
		X"00",X"00",X"09",X"44",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"05",X"30",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"35",X"00",X"03",X"30",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"33",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"45",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"FF",X"00",X"44",X"00",X"00",X"00",
		X"00",X"05",X"40",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"40",X"00",X"FF",X"00",
		X"00",X"00",X"09",X"90",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"05",X"50",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"04",X"40",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"33",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"FF",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",
		X"00",X"33",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"33",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"FF",
		X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"33",X"00",X"00",
		X"02",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"33",X"00",X"00",X"02",X"20",X"00",
		X"00",X"40",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"20",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"20",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"30",X"00",X"FF",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"30",
		X"00",X"FF",X"00",X"03",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"03",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"03",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"30",X"04",X"03",X"04",X"00",X"00",X"FF",X"00",X"03",X"00",
		X"3F",X"30",X"04",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"43",X"00",X"31",
		X"01",X"01",X"43",X"00",X"FF",X"00",X"00",X"10",X"02",X"00",X"00",X"30",X"FF",X"21",X"00",X"20",
		X"10",X"00",X"00",X"00",X"FF",X"00",X"10",X"01",X"00",X"10",X"01",X"42",X"FF",X"10",X"01",X"00",
		X"00",X"00",X"10",X"00",X"FF",X"10",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"00",X"01",X"01",
		X"00",X"00",X"12",X"10",X"FF",X"01",X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"00",X"20",X"01",
		X"02",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"10",X"34",X"00",X"FF",X"00",X"00",X"30",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"FF",X"00",X"00",X"01",
		X"10",X"01",X"10",X"00",X"00",X"00",X"FF",X"00",X"00",X"01",X"10",X"01",X"10",X"11",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"22",X"00",X"11",X"01",X"10",X"FF",X"00",X"11",X"03",X"00",X"22",
		X"30",X"00",X"01",X"10",X"FF",X"00",X"11",X"00",X"00",X"00",X"00",X"02",X"20",X"00",X"FF",X"00",
		X"02",X"21",X"10",X"00",X"00",X"02",X"20",X"11",X"FF",X"11",X"02",X"21",X"10",X"30",X"30",X"30",
		X"00",X"11",X"FF",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"FF",X"00",X"02",X"20",
		X"02",X"20",X"00",X"00",X"22",X"00",X"FF",X"00",X"02",X"23",X"02",X"20",X"00",X"00",X"22",X"00",
		X"FF",X"00",X"03",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"FF",X"00",X"00",X"02",X"20",X"00",
		X"30",X"00",X"00",X"11",X"FF",X"01",X"10",X"02",X"20",X"30",X"00",X"03",X"03",X"11",X"FF",X"01",
		X"10",X"30",X"00",X"00",X"02",X"20",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"30",X"02",X"20",
		X"22",X"00",X"FF",X"00",X"01",X"10",X"02",X"20",X"03",X"00",X"22",X"00",X"FF",X"00",X"01",X"10",
		X"02",X"20",X"00",X"01",X"10",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"10",X"00",
		X"FF",X"00",X"00",X"01",X"10",X"11",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"01",X"10",X"11",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"01",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"11",
		X"00",X"00",X"FF",X"00",X"00",X"01",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"30",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"10",X"03",X"00",X"03",X"00",X"00",X"FF",X"00",X"00",X"00",X"03",X"00",X"11",X"01",
		X"10",X"00",X"01",X"10",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"01",X"10",X"00",X"00",X"FF",X"00",X"00",X"00",X"01",X"10",X"00",X"00",X"01",X"10",X"00",X"00",
		X"30",X"00",X"FF",X"11",X"00",X"03",X"01",X"10",X"00",X"00",X"01",X"10",X"00",X"00",X"00",X"00",
		X"FF",X"11",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"01",X"10",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"30",X"00",X"11",X"00",X"00",X"00",X"01",X"10",X"00",X"11",X"FF",X"00",X"00",X"00",
		X"01",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"FF",X"00",X"00",X"00",X"01",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"10",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"01",X"10",X"00",X"00",X"00",
		X"01",X"10",X"03",X"00",X"FF",X"00",X"00",X"00",X"30",X"01",X"10",X"01",X"10",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"10",X"11",X"01",X"10",X"00",X"00",
		X"FF",X"00",X"01",X"10",X"00",X"00",X"00",X"00",X"00",X"11",X"01",X"10",X"00",X"00",X"FF",X"00",
		X"01",X"10",X"00",X"30",X"01",X"10",X"00",X"03",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"01",X"10",X"01",X"10",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"10",X"00",X"30",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"30",
		X"00",X"00",X"00",X"00",X"01",X"10",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",
		X"00",X"00",X"01",X"10",X"FF",X"00",X"00",X"00",X"00",X"01",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"01",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"22",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"00",
		X"00",X"FF",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"22",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"FF",X"00",
		X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"20",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"20",X"03",X"00",X"FF",
		X"30",X"02",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"02",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"02",X"20",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"02",X"20",X"00",X"02",X"20",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"20",
		X"00",X"FF",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"02",X"20",X"30",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"02",X"20",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"01",X"10",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"01",X"10",X"00",X"03",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"FF",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"FF",X"11",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"00",X"FF",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"10",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"10",X"FF",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"07",X"50",X"00",X"00",
		X"00",X"FF",X"00",X"E7",X"50",X"EA",X"E0",X"00",X"FF",X"00",X"5D",X"10",X"4A",X"E0",X"00",X"FF",
		X"EE",X"06",X"10",X"11",X"04",X"00",X"FF",X"EE",X"10",X"10",X"10",X"13",X"40",X"FF",X"E1",X"81",
		X"00",X"11",X"11",X"36",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"E1",X"81",X"00",X"11",
		X"11",X"36",X"FF",X"EE",X"10",X"10",X"10",X"13",X"40",X"FF",X"EE",X"06",X"10",X"11",X"05",X"E0",
		X"FF",X"E0",X"5D",X"10",X"4A",X"E0",X"00",X"FF",X"0E",X"E7",X"50",X"EA",X"E0",X"00",X"FF",X"00",
		X"E7",X"00",X"EE",X"00",X"00",X"FF",X"00",X"0E",X"E0",X"00",X"00",X"00",X"FF",X"00",X"00",X"01",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"00",X"00",X"11",X"10",X"00",
		X"00",X"FF",X"00",X"00",X"11",X"10",X"00",X"00",X"FF",X"00",X"01",X"11",X"11",X"00",X"00",X"FF",
		X"00",X"11",X"11",X"11",X"10",X"00",X"FF",X"11",X"11",X"11",X"11",X"11",X"10",X"FF",X"00",X"11",
		X"11",X"11",X"10",X"00",X"FF",X"00",X"01",X"11",X"11",X"00",X"00",X"FF",X"00",X"00",X"11",X"10",
		X"00",X"00",X"FF",X"00",X"00",X"11",X"10",X"00",X"00",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"65",X"00",X"00",X"00",X"00",X"FF",X"00",X"0E",X"7E",X"00",X"EB",X"E0",X"06",X"FF",
		X"06",X"00",X"DE",X"00",X"EB",X"E0",X"60",X"FF",X"00",X"60",X"0E",X"00",X"EB",X"66",X"00",X"FF",
		X"EE",X"06",X"60",X"06",X"66",X"60",X"00",X"FF",X"EE",X"E6",X"66",X"66",X"66",X"6E",X"E0",X"FF",
		X"EE",X"80",X"66",X"66",X"66",X"E4",X"56",X"FF",X"00",X"00",X"66",X"66",X"66",X"00",X"00",X"FF",
		X"EE",X"80",X"66",X"66",X"66",X"E4",X"56",X"FF",X"EE",X"06",X"66",X"66",X"66",X"E4",X"E0",X"FF",
		X"E0",X"06",X"66",X"66",X"66",X"6E",X"00",X"FF",X"00",X"66",X"DE",X"00",X"E6",X"60",X"00",X"FF",
		X"00",X"6E",X"DE",X"00",X"EB",X"06",X"00",X"FF",X"06",X"EE",X"7E",X"00",X"EB",X"E0",X"00",X"FF",
		X"60",X"0E",X"6E",X"00",X"EB",X"E0",X"00",X"FF",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"01",X"50",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"01",X"10",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"05",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"51",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"10",X"00",
		X"00",X"00",X"10",X"05",X"50",X"00",X"00",X"FF",X"00",X"00",X"00",X"01",X"00",X"01",X"11",X"01",
		X"50",X"00",X"00",X"FF",X"00",X"00",X"00",X"11",X"15",X"51",X"11",X"11",X"00",X"01",X"50",X"FF",
		X"00",X"00",X"55",X"01",X"15",X"51",X"11",X"10",X"00",X"11",X"50",X"FF",X"00",X"00",X"51",X"10",
		X"11",X"11",X"11",X"11",X"00",X"11",X"00",X"FF",X"00",X"00",X"00",X"11",X"11",X"11",X"11",X"11",
		X"00",X"00",X"00",X"FF",X"55",X"01",X"11",X"11",X"11",X"11",X"11",X"11",X"10",X"00",X"00",X"FF",
		X"55",X"01",X"11",X"11",X"11",X"11",X"11",X"10",X"00",X"11",X"15",X"FF",X"00",X"01",X"11",X"55",
		X"11",X"11",X"11",X"11",X"00",X"01",X"15",X"FF",X"00",X"00",X"11",X"55",X"11",X"11",X"11",X"01",
		X"15",X"00",X"00",X"FF",X"00",X"00",X"01",X"11",X"11",X"11",X"11",X"10",X"55",X"00",X"00",X"FF",
		X"00",X"00",X"11",X"11",X"11",X"11",X"11",X"10",X"00",X"00",X"00",X"FF",X"00",X"00",X"11",X"01",
		X"11",X"11",X"11",X"11",X"00",X"00",X"00",X"FF",X"00",X"00",X"10",X"01",X"11",X"11",X"11",X"10",
		X"00",X"00",X"00",X"FF",X"00",X"51",X"00",X"51",X"01",X"11",X"00",X"00",X"11",X"00",X"00",X"FF",
		X"00",X"05",X"00",X"55",X"01",X"10",X"00",X"00",X"01",X"50",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"05",X"50",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"01",X"10",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"10",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"05",X"50",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"01",X"11",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"05",X"11",X"55",X"55",X"00",X"00",X"00",X"FF",X"00",X"01",X"15",X"11",
		X"51",X"15",X"11",X"00",X"00",X"FF",X"00",X"55",X"55",X"11",X"77",X"71",X"55",X"50",X"00",X"FF",
		X"05",X"51",X"15",X"77",X"66",X"67",X"71",X"15",X"00",X"FF",X"05",X"51",X"17",X"66",X"67",X"76",
		X"77",X"15",X"00",X"FF",X"15",X"15",X"76",X"77",X"77",X"22",X"66",X"75",X"10",X"FF",X"55",X"11",
		X"73",X"73",X"23",X"23",X"36",X"65",X"10",X"FF",X"51",X"17",X"67",X"72",X"23",X"32",X"23",X"67",
		X"11",X"FF",X"51",X"17",X"77",X"22",X"22",X"23",X"23",X"67",X"51",X"FF",X"51",X"16",X"73",X"22",
		X"22",X"23",X"22",X"76",X"51",X"FF",X"15",X"17",X"63",X"32",X"22",X"33",X"22",X"76",X"51",X"FF",
		X"15",X"17",X"66",X"32",X"33",X"32",X"77",X"66",X"51",X"FF",X"51",X"11",X"76",X"63",X"33",X"27",
		X"76",X"75",X"51",X"FF",X"05",X"15",X"77",X"66",X"36",X"76",X"67",X"21",X"10",X"FF",X"05",X"15",
		X"17",X"77",X"77",X"66",X"67",X"51",X"10",X"FF",X"05",X"55",X"11",X"27",X"76",X"66",X"71",X"51",
		X"00",X"FF",X"00",X"15",X"11",X"11",X"77",X"75",X"15",X"51",X"00",X"FF",X"00",X"05",X"51",X"11",
		X"51",X"11",X"55",X"10",X"00",X"FF",X"00",X"00",X"11",X"15",X"55",X"11",X"11",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"11",X"11",X"11",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"01",X"11",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"01",X"00",X"00",
		X"00",X"00",X"00",X"01",X"00",X"FF",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"FF",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"10",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"FF",X"00",X"10",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"FF",X"00",X"00",
		X"01",X"00",X"01",X"00",X"00",X"10",X"00",X"FF",X"00",X"00",X"01",X"10",X"00",X"11",X"00",X"00",
		X"00",X"FF",X"10",X"FF",X"51",X"10",X"00",X"00",X"00",X"00",X"00",X"05",X"10",X"FF",X"51",X"10",
		X"00",X"00",X"00",X"00",X"00",X"01",X"50",X"FF",X"51",X"10",X"00",X"00",X"00",X"00",X"00",X"01",
		X"50",X"FF",X"15",X"10",X"00",X"00",X"00",X"00",X"00",X"01",X"50",X"FF",X"15",X"10",X"00",X"00",
		X"00",X"00",X"00",X"01",X"50",X"FF",X"51",X"11",X"00",X"00",X"00",X"00",X"00",X"15",X"50",X"FF",
		X"15",X"15",X"00",X"00",X"00",X"00",X"00",X"11",X"10",X"FF",X"05",X"15",X"10",X"00",X"00",X"00",
		X"01",X"51",X"00",X"FF",X"05",X"55",X"11",X"10",X"00",X"01",X"11",X"51",X"00",X"FF",X"00",X"15",
		X"11",X"11",X"11",X"15",X"15",X"50",X"00",X"FF",X"00",X"05",X"51",X"11",X"51",X"11",X"55",X"00",
		X"00",X"FF",X"00",X"00",X"01",X"15",X"55",X"11",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"01",
		X"11",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"FF",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"FF",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"10",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"FF",X"00",X"10",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"FF",
		X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"10",X"00",X"FF",X"00",X"00",X"01",X"10",X"00",X"11",
		X"00",X"00",X"00",X"FF",X"55",X"00",X"00",X"00",X"00",X"FF",X"53",X"55",X"57",X"70",X"00",X"FF",
		X"05",X"23",X"55",X"57",X"00",X"FF",X"05",X"32",X"23",X"55",X"70",X"FF",X"05",X"52",X"11",X"35",
		X"70",X"FF",X"07",X"53",X"11",X"25",X"50",X"FF",X"07",X"55",X"32",X"23",X"50",X"FF",X"00",X"75",
		X"55",X"32",X"50",X"FF",X"00",X"07",X"75",X"55",X"35",X"FF",X"00",X"00",X"00",X"00",X"55",X"FF",
		X"00",X"00",X"00",X"00",X"55",X"FF",X"00",X"07",X"75",X"55",X"35",X"FF",X"00",X"75",X"55",X"32",
		X"50",X"FF",X"07",X"55",X"32",X"23",X"50",X"FF",X"07",X"53",X"11",X"25",X"50",X"FF",X"05",X"52",
		X"11",X"35",X"70",X"FF",X"05",X"32",X"23",X"55",X"70",X"FF",X"05",X"23",X"55",X"57",X"00",X"FF",
		X"53",X"55",X"57",X"70",X"00",X"FF",X"55",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"55",X"00",
		X"00",X"FF",X"00",X"05",X"33",X"50",X"00",X"FF",X"00",X"75",X"22",X"57",X"00",X"FF",X"07",X"53",
		X"22",X"35",X"70",X"FF",X"07",X"53",X"11",X"35",X"70",X"FF",X"77",X"32",X"11",X"23",X"77",X"FF",
		X"77",X"32",X"11",X"23",X"77",X"FF",X"07",X"53",X"11",X"35",X"70",X"FF",X"07",X"53",X"22",X"35",
		X"70",X"FF",X"00",X"75",X"22",X"57",X"00",X"FF",X"00",X"05",X"33",X"50",X"00",X"FF",X"00",X"00",
		X"55",X"00",X"00",X"FF",X"00",X"00",X"77",X"77",X"00",X"00",X"FF",X"00",X"07",X"55",X"55",X"70",
		X"00",X"FF",X"00",X"75",X"33",X"33",X"57",X"00",X"FF",X"05",X"53",X"22",X"22",X"35",X"50",X"FF",
		X"53",X"22",X"11",X"11",X"22",X"35",X"FF",X"53",X"22",X"11",X"11",X"22",X"35",X"FF",X"05",X"53",
		X"22",X"22",X"35",X"50",X"FF",X"00",X"75",X"33",X"33",X"57",X"00",X"FF",X"00",X"07",X"55",X"55",
		X"70",X"00",X"FF",X"00",X"00",X"77",X"77",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"0C",X"CC",
		X"CC",X"C0",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0C",X"CB",X"BB",X"BB",X"BC",X"C0",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"CB",X"BB",X"BB",X"BB",X"BB",X"BC",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"0C",X"BB",X"BA",X"AA",X"AA",X"AB",X"BB",X"C0",X"00",X"00",X"FF",X"00",X"00",
		X"CB",X"BA",X"AA",X"AA",X"AA",X"AA",X"AB",X"BC",X"00",X"00",X"FF",X"00",X"0C",X"BB",X"AA",X"A9",
		X"99",X"99",X"9A",X"AA",X"BB",X"C0",X"00",X"FF",X"00",X"CB",X"BA",X"A9",X"99",X"99",X"99",X"99",
		X"9A",X"AB",X"BC",X"00",X"FF",X"00",X"CB",X"AA",X"99",X"99",X"88",X"88",X"99",X"99",X"AA",X"BC",
		X"00",X"FF",X"0C",X"BB",X"A9",X"99",X"88",X"87",X"78",X"88",X"99",X"9A",X"BB",X"C0",X"FF",X"0C",
		X"BA",X"A9",X"98",X"87",X"77",X"77",X"78",X"89",X"9A",X"AB",X"C0",X"FF",X"0C",X"BA",X"99",X"88",
		X"77",X"76",X"67",X"77",X"88",X"99",X"AB",X"C0",X"FF",X"CB",X"BA",X"99",X"87",X"76",X"65",X"56",
		X"67",X"78",X"99",X"AB",X"BC",X"FF",X"CB",X"A9",X"98",X"87",X"65",X"54",X"45",X"56",X"78",X"89",
		X"9A",X"BC",X"FF",X"CB",X"A9",X"98",X"77",X"65",X"43",X"34",X"56",X"77",X"89",X"9A",X"BC",X"FF",
		X"CB",X"A9",X"98",X"76",X"54",X"32",X"23",X"45",X"67",X"89",X"9A",X"BC",X"FF",X"CB",X"A9",X"98",
		X"76",X"54",X"21",X"12",X"45",X"67",X"89",X"9A",X"BC",X"FF",X"CB",X"A9",X"98",X"76",X"54",X"21",
		X"12",X"45",X"67",X"89",X"9A",X"BC",X"FF",X"CB",X"A9",X"98",X"76",X"54",X"32",X"23",X"45",X"67",
		X"89",X"9A",X"BC",X"FF",X"CB",X"A9",X"98",X"77",X"65",X"43",X"34",X"56",X"77",X"89",X"9A",X"BC",
		X"FF",X"CB",X"A9",X"98",X"87",X"65",X"54",X"45",X"56",X"78",X"89",X"9A",X"BC",X"FF",X"CB",X"BA",
		X"99",X"87",X"76",X"65",X"56",X"67",X"78",X"99",X"AB",X"BC",X"FF",X"0C",X"BA",X"99",X"88",X"77",
		X"76",X"67",X"77",X"88",X"99",X"AB",X"C0",X"FF",X"0C",X"BA",X"A9",X"98",X"87",X"77",X"77",X"78",
		X"89",X"9A",X"AB",X"C0",X"FF",X"0C",X"BB",X"A9",X"99",X"88",X"87",X"78",X"88",X"99",X"9A",X"BB",
		X"C0",X"FF",X"00",X"CB",X"AA",X"99",X"99",X"88",X"88",X"99",X"99",X"AA",X"BC",X"00",X"FF",X"00",
		X"CB",X"BA",X"A9",X"99",X"99",X"99",X"99",X"9A",X"AB",X"BC",X"00",X"FF",X"00",X"0C",X"BB",X"AA",
		X"A9",X"99",X"99",X"9A",X"AA",X"BB",X"C0",X"00",X"FF",X"00",X"00",X"CB",X"BA",X"AA",X"AA",X"AA",
		X"AA",X"AB",X"BC",X"00",X"00",X"FF",X"00",X"00",X"0C",X"BB",X"BA",X"AA",X"AA",X"AB",X"BB",X"C0",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"CB",X"BB",X"BB",X"BB",X"BB",X"BC",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"0C",X"CB",X"BB",X"BB",X"BC",X"C0",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"0C",X"CC",X"CC",X"C0",X"00",X"00",X"00",X"00",X"FF",X"56",X"A8",X"8A",X"77",X"76",X"54",
		X"32",X"11",X"FF",X"00",X"00",X"33",X"59",X"88",X"AA",X"75",X"50",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"33",X"77",X"66",X"AA",X"95",X"33",X"00",X"00",X"00",X"FF",X"00",X"00",X"06",X"64",X"46",
		X"99",X"0A",X"33",X"00",X"00",X"00",X"FF",X"00",X"00",X"55",X"64",X"49",X"77",X"00",X"65",X"50",
		X"00",X"00",X"FF",X"00",X"04",X"45",X"00",X"08",X"85",X"50",X"05",X"44",X"00",X"00",X"FF",X"00",
		X"33",X"40",X"00",X"07",X"70",X"33",X"00",X"43",X"30",X"00",X"FF",X"02",X"23",X"00",X"00",X"06",
		X"60",X"33",X"00",X"03",X"22",X"00",X"FF",X"11",X"20",X"00",X"00",X"05",X"50",X"00",X"00",X"00",
		X"21",X"10",X"FF",X"11",X"00",X"00",X"00",X"04",X"40",X"00",X"00",X"00",X"01",X"10",X"FF",X"00",
		X"00",X"00",X"00",X"03",X"30",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"02",
		X"20",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"01",X"10",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"01",X"10",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"FF",X"02",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"11",X"FF",X"02",X"23",X"00",X"00",X"02",X"20",X"00",X"00",X"32",X"20",X"FF",
		X"00",X"33",X"40",X"00",X"03",X"30",X"00",X"04",X"33",X"00",X"FF",X"00",X"04",X"45",X"02",X"24",
		X"40",X"00",X"54",X"40",X"00",X"FF",X"00",X"00",X"55",X"62",X"25",X"50",X"06",X"55",X"00",X"00",
		X"FF",X"00",X"00",X"06",X"63",X"36",X"60",X"06",X"60",X"00",X"00",X"FF",X"02",X"30",X"22",X"77",
		X"44",X"70",X"73",X"30",X"32",X"00",X"FF",X"03",X"34",X"22",X"38",X"85",X"88",X"43",X"34",X"43",
		X"00",X"FF",X"00",X"44",X"53",X"34",X"95",X"57",X"44",X"54",X"40",X"00",X"FF",X"22",X"05",X"56",
		X"44",X"57",X"59",X"77",X"55",X"33",X"00",X"FF",X"22",X"45",X"66",X"75",X"58",X"A9",X"91",X"14",
		X"33",X"00",X"FF",X"00",X"45",X"67",X"78",X"88",X"B7",X"41",X"14",X"40",X"00",X"FF",X"00",X"00",
		X"77",X"9A",X"94",X"47",X"44",X"66",X"00",X"00",X"FF",X"00",X"02",X"34",X"5A",X"A4",X"48",X"78",
		X"76",X"54",X"32",X"FF",X"00",X"02",X"36",X"7A",X"A8",X"8A",X"77",X"76",X"54",X"32",X"FF",X"00",
		X"04",X"56",X"79",X"88",X"AA",X"75",X"50",X"00",X"00",X"FF",X"03",X"34",X"50",X"77",X"66",X"AA",
		X"95",X"44",X"00",X"00",X"FF",X"22",X"30",X"06",X"65",X"55",X"99",X"0A",X"43",X"30",X"00",X"FF",
		X"22",X"00",X"55",X"64",X"49",X"88",X"00",X"63",X"22",X"00",X"FF",X"00",X"04",X"45",X"33",X"48",
		X"87",X"70",X"05",X"22",X"00",X"FF",X"00",X"33",X"40",X"33",X"07",X"70",X"66",X"00",X"43",X"30",
		X"FF",X"00",X"23",X"00",X"00",X"06",X"60",X"55",X"00",X"03",X"20",X"FF",X"00",X"00",X"00",X"00",
		X"05",X"50",X"44",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"04",X"40",X"03",X"30",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"03",X"30",X"03",X"22",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"02",X"20",X"00",X"22",X"00",X"00",X"FF",X"01",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"01",X"12",X"00",X"00",X"00",X"01",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"22",X"30",X"00",X"00",X"01",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"03",X"34",X"00",X"00",X"02",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"44",X"50",X"00",X"03",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"05",X"56",X"00",X"04",X"40",X"00",X"00",X"00",X"32",X"00",X"00",X"FF",X"00",X"00",X"11",X"66",
		X"70",X"00",X"55",X"00",X"00",X"04",X"33",X"00",X"00",X"FF",X"00",X"00",X"11",X"27",X"78",X"00",
		X"66",X"00",X"00",X"54",X"22",X"00",X"00",X"FF",X"00",X"00",X"02",X"23",X"88",X"90",X"77",X"50",
		X"06",X"53",X"22",X"00",X"00",X"FF",X"00",X"00",X"00",X"33",X"49",X"9A",X"55",X"60",X"06",X"43",
		X"30",X"00",X"00",X"FF",X"00",X"00",X"00",X"04",X"45",X"AA",X"66",X"60",X"75",X"44",X"32",X"00",
		X"00",X"FF",X"11",X"30",X"00",X"00",X"55",X"68",X"87",X"88",X"65",X"54",X"43",X"00",X"22",X"FF",
		X"11",X"34",X"50",X"04",X"56",X"67",X"95",X"57",X"66",X"54",X"40",X"03",X"22",X"FF",X"00",X"44",
		X"56",X"05",X"56",X"77",X"87",X"59",X"77",X"55",X"65",X"43",X"00",X"FF",X"00",X"00",X"66",X"78",
		X"9A",X"78",X"89",X"A9",X"97",X"97",X"65",X"40",X"00",X"FF",X"00",X"00",X"00",X"78",X"9A",X"78",
		X"99",X"A7",X"55",X"97",X"40",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"77",X"9A",X"97",X"77",
		X"55",X"66",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"04",X"5A",X"A7",X"7A",X"A8",X"76",
		X"50",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"09",X"AA",X"A8",X"8A",X"99",X"76",X"50",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"67",X"89",X"A9",X"88",X"AA",X"98",X"80",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"45",X"67",X"80",X"77",X"99",X"AA",X"98",X"77",X"00",X"00",X"00",X"FF",X"00",X"33",
		X"45",X"00",X"06",X"65",X"77",X"AA",X"0A",X"76",X"60",X"00",X"00",X"FF",X"01",X"13",X"00",X"00",
		X"55",X"66",X"69",X"AA",X"00",X"66",X"55",X"00",X"00",X"FF",X"01",X"10",X"00",X"00",X"45",X"77",
		X"78",X"8A",X"A0",X"05",X"54",X"40",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"66",X"07",X"70",
		X"99",X"00",X"04",X"33",X"00",X"FF",X"00",X"00",X"00",X"00",X"05",X"50",X"06",X"60",X"88",X"00",
		X"00",X"32",X"20",X"FF",X"00",X"00",X"00",X"00",X"04",X"40",X"05",X"50",X"77",X"00",X"00",X"02",
		X"11",X"FF",X"00",X"00",X"00",X"00",X"33",X"30",X"00",X"00",X"06",X"60",X"00",X"00",X"11",X"FF",
		X"00",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"05",X"52",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"01",X"10",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"01",
		X"10",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"21",X"10",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"10",X"00",X"00",X"FF",X"12",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"22",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"03",X"34",X"00",X"00",X"02",X"20",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",
		X"FF",X"00",X"44",X"50",X"00",X"03",X"30",X"00",X"00",X"00",X"00",X"02",X"11",X"00",X"00",X"FF",
		X"00",X"05",X"56",X"00",X"04",X"40",X"00",X"00",X"00",X"00",X"32",X"20",X"00",X"00",X"FF",X"00",
		X"00",X"66",X"70",X"00",X"55",X"00",X"00",X"00",X"04",X"33",X"00",X"00",X"00",X"FF",X"00",X"01",
		X"27",X"78",X"00",X"66",X"00",X"00",X"00",X"54",X"40",X"00",X"00",X"00",X"FF",X"00",X"02",X"23",
		X"88",X"90",X"77",X"50",X"00",X"06",X"55",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"33",X"49",
		X"9A",X"55",X"60",X"06",X"76",X"60",X"00",X"00",X"00",X"11",X"FF",X"00",X"00",X"04",X"45",X"AA",
		X"66",X"60",X"78",X"77",X"00",X"00",X"00",X"02",X"11",X"FF",X"00",X"00",X"00",X"55",X"68",X"87",
		X"88",X"98",X"84",X"00",X"00",X"54",X"32",X"20",X"FF",X"34",X"50",X"00",X"06",X"67",X"95",X"5A",
		X"99",X"54",X"40",X"06",X"54",X"30",X"00",X"FF",X"44",X"56",X"00",X"06",X"77",X"87",X"59",X"A7",
		X"55",X"68",X"76",X"00",X"00",X"00",X"FF",X"00",X"66",X"78",X"9A",X"78",X"89",X"A9",X"97",X"97",
		X"98",X"70",X"00",X"00",X"00",X"FF",X"00",X"00",X"78",X"9A",X"78",X"99",X"A7",X"55",X"97",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"77",X"9A",X"97",X"77",X"55",X"60",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"33",X"A7",X"7A",X"A8",X"76",X"54",X"40",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"09",X"33",X"A8",X"8A",X"99",X"76",X"54",X"40",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"67",X"89",X"A9",X"88",X"A4",X"48",X"80",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"45",X"67",X"80",X"77",X"99",X"A4",X"48",X"77",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"33",X"45",X"00",X"00",X"05",X"77",X"AA",X"0A",X"76",X"60",X"00",X"00",X"00",X"00",X"FF",X"13",
		X"00",X"00",X"00",X"06",X"69",X"AA",X"00",X"66",X"55",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"77",X"78",X"8A",X"A0",X"05",X"54",X"40",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"66",X"07",X"70",X"99",X"00",X"04",X"33",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"05",
		X"50",X"00",X"00",X"88",X"00",X"00",X"32",X"20",X"00",X"00",X"FF",X"00",X"00",X"00",X"04",X"40",
		X"00",X"00",X"77",X"00",X"00",X"02",X"10",X"00",X"00",X"FF",X"00",X"00",X"00",X"33",X"30",X"00",
		X"00",X"06",X"60",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"22",X"00",X"00",X"00",
		X"05",X"52",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"34",X"00",X"00",X"02",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"44",X"50",X"00",X"03",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"05",X"56",X"00",X"04",X"40",X"00",X"00",X"00",X"00",X"32",X"00",X"00",X"FF",X"00",X"00",
		X"66",X"70",X"00",X"55",X"00",X"00",X"00",X"04",X"33",X"00",X"00",X"FF",X"00",X"00",X"07",X"70",
		X"00",X"66",X"00",X"00",X"00",X"54",X"40",X"00",X"00",X"FF",X"00",X"00",X"23",X"00",X"00",X"77",
		X"50",X"00",X"06",X"55",X"00",X"00",X"00",X"FF",X"00",X"00",X"33",X"40",X"00",X"55",X"60",X"06",
		X"76",X"60",X"00",X"00",X"00",X"FF",X"00",X"00",X"04",X"45",X"00",X"66",X"60",X"70",X"77",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"55",X"60",X"07",X"00",X"00",X"04",X"00",X"00",X"54",
		X"32",X"FF",X"34",X"50",X"00",X"06",X"67",X"05",X"50",X"00",X"54",X"40",X"06",X"54",X"30",X"FF",
		X"44",X"56",X"00",X"06",X"77",X"07",X"50",X"07",X"55",X"60",X"76",X"00",X"00",X"FF",X"00",X"66",
		X"70",X"00",X"70",X"00",X"00",X"07",X"07",X"00",X"70",X"00",X"00",X"FF",X"00",X"00",X"70",X"00",
		X"70",X"00",X"07",X"55",X"07",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"77",X"00",X"07",
		X"77",X"55",X"60",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"33",X"07",X"70",X"00",
		X"76",X"54",X"40",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"76",X"54",
		X"40",X"00",X"00",X"FF",X"00",X"00",X"67",X"00",X"00",X"00",X"04",X"40",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"45",X"67",X"00",X"77",X"00",X"04",X"40",X"77",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"45",X"00",X"00",X"05",X"77",X"00",X"00",X"76",X"60",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"06",X"60",X"00",X"00",X"66",X"55",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"77",X"70",X"00",X"00",X"05",X"54",X"40",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"66",X"07",
		X"70",X"00",X"00",X"04",X"33",X"00",X"00",X"FF",X"00",X"00",X"00",X"05",X"50",X"00",X"00",X"00",
		X"00",X"00",X"32",X"00",X"00",X"FF",X"00",X"00",X"00",X"04",X"40",X"00",X"00",X"77",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"03",X"30",X"00",X"00",X"06",X"60",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"55",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"00",X"FF",X"01",X"10",X"00",X"01",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"01",X"16",X"00",X"01",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"00",X"66",X"00",X"00",X"55",X"00",X"00",X"00",X"01",X"10",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"51",X"10",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"50",X"00",X"06",X"55",X"00",X"00",X"FF",X"00",X"01",X"10",X"00",X"00",X"60",X"00",X"06",
		X"60",X"00",X"00",X"FF",X"00",X"01",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"55",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"FF",X"00",X"00",X"06",X"60",
		X"05",X"50",X"00",X"00",X"00",X"06",X"11",X"FF",X"11",X"00",X"00",X"00",X"00",X"50",X"00",X"00",
		X"00",X"06",X"00",X"FF",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"06",
		X"51",X"10",X"00",X"FF",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"06",X"51",X"10",X"00",X"FF",
		X"00",X"11",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"FF",X"00",X"11",X"00",X"00",
		X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"06",X"60",X"00",X"00",X"06",X"11",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"FF",X"00",X"00",X"00",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"01",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"01",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"60",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"05",X"11",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"FF",X"00",X"B0",X"00",X"05",X"30",X"00",X"FF",X"00",X"05",X"30",X"55",X"04",
		X"BB",X"FF",X"0E",X"B2",X"22",X"22",X"20",X"00",X"FF",X"E5",X"D8",X"86",X"66",X"00",X"00",X"FF",
		X"6E",X"BC",X"CC",X"CC",X"C0",X"00",X"FF",X"06",X"6B",X"46",X"5B",X"05",X"BB",X"FF",X"00",X"B0",
		X"00",X"65",X"40",X"00",X"FF",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"20",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"02",X"05",X"5B",X"44",X"BB",X"B0",X"FF",
		X"00",X"EB",X"23",X"33",X"00",X"00",X"00",X"00",X"FF",X"0B",X"BB",X"88",X"44",X"40",X"00",X"00",
		X"00",X"FF",X"66",X"EB",X"CE",X"EE",X"60",X"00",X"00",X"00",X"FF",X"06",X"66",X"6C",X"65",X"BB",
		X"44",X"BB",X"B0",X"FF",X"00",X"00",X"60",X"C6",X"60",X"00",X"00",X"00",X"FF",X"00",X"00",X"06",
		X"0C",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"06",X"20",X"20",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"06",X"22",X"20",X"00",X"00",X"00",X"00",X"FF",X"00",X"06",X"22",X"05",X"5B",X"40",
		X"00",X"00",X"FF",X"00",X"EB",X"23",X"33",X"00",X"04",X"BB",X"B0",X"FF",X"0B",X"BB",X"88",X"44",
		X"40",X"00",X"00",X"00",X"FF",X"00",X"EB",X"CE",X"EE",X"60",X"04",X"BB",X"B0",X"FF",X"06",X"66",
		X"CC",X"75",X"BB",X"40",X"00",X"00",X"FF",X"66",X"66",X"CC",X"C7",X"60",X"00",X"00",X"00",X"FF",
		X"06",X"66",X"C7",X"C0",X"00",X"00",X"00",X"00",X"FF",X"00",X"06",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"06",X"66",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"06",X"06",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"02",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"02",X"20",X"02",X"00",X"00",X"00",X"FF",X"00",X"00",X"20",
		X"20",X"00",X"00",X"00",X"FF",X"00",X"60",X"22",X"05",X"50",X"00",X"00",X"FF",X"00",X"EB",X"23",
		X"33",X"04",X"00",X"00",X"FF",X"0B",X"BB",X"88",X"44",X"40",X"45",X"BB",X"FF",X"00",X"EB",X"CE",
		X"EE",X"64",X"00",X"00",X"FF",X"06",X"66",X"CC",X"65",X"B0",X"00",X"00",X"FF",X"66",X"66",X"C6",
		X"C6",X"60",X"00",X"00",X"FF",X"06",X"6C",X"C6",X"6C",X"00",X"00",X"00",X"FF",X"00",X"0C",X"66",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"06",X"06",X"60",X"00",X"00",X"00",X"FF",X"00",X"66",X"00",
		X"60",X"00",X"00",X"00",X"FF",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"FF",X"0C",X"66",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"06",X"06",X"60",X"00",X"00",X"00",X"00",X"FF",X"00",X"66",
		X"00",X"60",X"00",X"00",X"00",X"00",X"FF",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"11",X"00",X"00",X"FF",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"0B",X"B0",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"0B",X"B0",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"01",X"10",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"01",X"10",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"07",X"50",X"00",X"00",X"00",
		X"FF",X"00",X"E7",X"55",X"EA",X"E0",X"00",X"FF",X"0E",X"5D",X"44",X"4A",X"EC",X"00",X"FF",X"EE",
		X"56",X"32",X"22",X"44",X"00",X"FF",X"EE",X"E6",X"21",X"11",X"23",X"40",X"FF",X"EE",X"8E",X"EE",
		X"11",X"12",X"36",X"FF",X"EE",X"81",X"1E",X"66",X"EE",X"E0",X"FF",X"EE",X"8E",X"EE",X"22",X"23",
		X"36",X"FF",X"EE",X"E6",X"23",X"33",X"33",X"40",X"FF",X"EE",X"46",X"33",X"34",X"45",X"E0",X"FF",
		X"EE",X"5D",X"44",X"4A",X"EC",X"00",X"FF",X"0E",X"E7",X"55",X"EA",X"E0",X"00",X"FF",X"00",X"E7",
		X"5E",X"EE",X"00",X"00",X"FF",X"00",X"0E",X"EE",X"00",X"00",X"00",X"FF",X"00",X"05",X"50",X"00",
		X"00",X"00",X"FF",X"00",X"E7",X"55",X"AE",X"B0",X"00",X"FF",X"0E",X"57",X"44",X"4E",X"BE",X"00",
		X"FF",X"EE",X"56",X"32",X"24",X"44",X"00",X"FF",X"EE",X"E6",X"21",X"11",X"23",X"40",X"FF",X"EE",
		X"8E",X"EE",X"11",X"12",X"36",X"FF",X"EE",X"81",X"1E",X"66",X"EE",X"E0",X"FF",X"EE",X"8E",X"EE",
		X"22",X"23",X"36",X"FF",X"EE",X"E6",X"23",X"33",X"33",X"40",X"FF",X"EE",X"46",X"33",X"34",X"45",
		X"E0",X"FF",X"EE",X"57",X"44",X"5E",X"BE",X"00",X"FF",X"0E",X"E7",X"55",X"AE",X"B0",X"00",X"FF",
		X"00",X"E5",X"5E",X"EE",X"E0",X"00",X"FF",X"00",X"0E",X"EE",X"E0",X"00",X"00",X"FF",X"00",X"00",
		X"0C",X"C0",X"00",X"60",X"FF",X"00",X"00",X"EE",X"44",X"42",X"E0",X"FF",X"00",X"55",X"44",X"32",
		X"1E",X"E6",X"FF",X"0E",X"77",X"43",X"21",X"EE",X"30",X"FF",X"EE",X"46",X"11",X"16",X"62",X"30",
		X"FF",X"EE",X"52",X"EE",X"E6",X"12",X"30",X"FF",X"EE",X"EE",X"11",X"E1",X"23",X"40",X"FF",X"EE",
		X"E8",X"11",X"E1",X"34",X"C0",X"FF",X"0E",X"E8",X"8E",X"14",X"45",X"C0",X"FF",X"0E",X"EE",X"8E",
		X"64",X"4E",X"00",X"FF",X"00",X"EE",X"EE",X"57",X"50",X"00",X"FF",X"00",X"0E",X"EE",X"57",X"50",
		X"00",X"FF",X"00",X"00",X"0E",X"EE",X"00",X"00",X"FF",X"00",X"00",X"0E",X"E0",X"00",X"60",X"FF",
		X"00",X"00",X"BB",X"44",X"42",X"E0",X"FF",X"00",X"55",X"44",X"32",X"1E",X"E6",X"FF",X"0E",X"7D",
		X"43",X"21",X"EE",X"30",X"FF",X"EE",X"46",X"11",X"16",X"62",X"30",X"FF",X"EE",X"52",X"EE",X"E6",
		X"12",X"30",X"FF",X"EE",X"EE",X"11",X"E1",X"23",X"40",X"FF",X"EE",X"E8",X"11",X"E1",X"34",X"E0",
		X"FF",X"0E",X"E8",X"8E",X"14",X"44",X"E0",X"FF",X"0E",X"EE",X"8E",X"64",X"4B",X"00",X"FF",X"00",
		X"EE",X"EE",X"5D",X"50",X"00",X"FF",X"00",X"0E",X"EE",X"57",X"50",X"00",X"FF",X"00",X"00",X"0E",
		X"EE",X"00",X"00",X"FF",X"00",X"00",X"E6",X"06",X"00",X"00",X"FF",X"00",X"00",X"E3",X"E3",X"00",
		X"00",X"FF",X"00",X"0E",X"53",X"E3",X"40",X"00",X"FF",X"00",X"EE",X"43",X"E3",X"40",X"00",X"FF",
		X"0E",X"EC",X"42",X"E1",X"3C",X"00",X"FF",X"0E",X"EE",X"42",X"E1",X"3E",X"E0",X"FF",X"EE",X"B5",
		X"32",X"61",X"24",X"B0",X"FF",X"EE",X"E4",X"32",X"61",X"24",X"E0",X"FF",X"EE",X"54",X"2E",X"EE",
		X"24",X"40",X"FF",X"EE",X"54",X"2E",X"1E",X"24",X"40",X"FF",X"EE",X"D7",X"6E",X"1E",X"67",X"D0",
		X"FF",X"EE",X"54",X"4E",X"8E",X"45",X"50",X"FF",X"0E",X"E5",X"E8",X"88",X"E5",X"E0",X"FF",X"00",
		X"EE",X"EE",X"EE",X"EE",X"00",X"FF",X"00",X"0E",X"EE",X"EE",X"E0",X"00",X"FF",X"00",X"00",X"E6",
		X"06",X"00",X"00",X"FF",X"00",X"00",X"E3",X"E3",X"00",X"00",X"FF",X"00",X"0E",X"53",X"E3",X"40",
		X"00",X"FF",X"00",X"EE",X"43",X"E3",X"40",X"00",X"FF",X"0E",X"EE",X"42",X"E1",X"3E",X"00",X"FF",
		X"0E",X"BB",X"42",X"E1",X"3B",X"B0",X"FF",X"EE",X"E5",X"32",X"61",X"24",X"E0",X"FF",X"EE",X"A4",
		X"32",X"61",X"24",X"A0",X"FF",X"EE",X"54",X"2E",X"EE",X"24",X"40",X"FF",X"EE",X"54",X"2E",X"1E",
		X"24",X"40",X"FF",X"EE",X"D7",X"6E",X"1E",X"67",X"D0",X"FF",X"EE",X"54",X"4E",X"8E",X"45",X"50",
		X"FF",X"0E",X"E5",X"E8",X"88",X"E5",X"E0",X"FF",X"00",X"EE",X"EE",X"EE",X"EE",X"00",X"FF",X"00",
		X"0E",X"EE",X"EE",X"E0",X"00",X"FF",X"0E",X"54",X"00",X"00",X"00",X"FF",X"EC",X"74",X"EA",X"00",
		X"00",X"FF",X"EC",X"73",X"44",X"00",X"00",X"FF",X"EE",X"74",X"34",X"54",X"00",X"FF",X"0E",X"E6",
		X"43",X"45",X"50",X"FF",X"E8",X"8E",X"6E",X"E3",X"55",X"FF",X"E8",X"88",X"E1",X"1E",X"E0",X"FF",
		X"E8",X"8E",X"6E",X"E3",X"55",X"FF",X"EE",X"E6",X"54",X"45",X"50",X"FF",X"0E",X"75",X"44",X"54",
		X"00",X"FF",X"EC",X"75",X"44",X"00",X"00",X"FF",X"EC",X"75",X"EA",X"00",X"00",X"FF",X"EE",X"55",
		X"00",X"00",X"00",X"FF",X"0E",X"E0",X"00",X"00",X"00",X"FF",X"00",X"EE",X"40",X"00",X"FF",X"EB",
		X"EC",X"43",X"00",X"FF",X"EB",X"EC",X"43",X"40",X"FF",X"EE",X"EE",X"E3",X"40",X"FF",X"00",X"EE",
		X"EE",X"34",X"FF",X"0E",X"E8",X"8E",X"E3",X"FF",X"0E",X"E8",X"88",X"E1",X"FF",X"0E",X"E8",X"8E",
		X"E4",X"FF",X"0E",X"EE",X"EE",X"55",X"FF",X"00",X"EE",X"E5",X"50",X"FF",X"EB",X"EC",X"55",X"50",
		X"FF",X"EB",X"EC",X"55",X"00",X"FF",X"EE",X"EE",X"50",X"00",X"FF",X"B5",X"00",X"FF",X"B5",X"00",
		X"FF",X"0E",X"50",X"FF",X"E8",X"E5",X"FF",X"E8",X"E4",X"FF",X"0E",X"50",X"FF",X"B5",X"00",X"FF",
		X"B5",X"00",X"FF",X"00",X"00",X"00",X"55",X"00",X"FF",X"05",X"7E",X"55",X"55",X"00",X"FF",X"CE",
		X"46",X"44",X"4E",X"05",X"FF",X"CE",X"E4",X"45",X"EE",X"45",X"FF",X"EE",X"EE",X"11",X"E3",X"45",
		X"FF",X"0E",X"E8",X"E1",X"23",X"40",X"FF",X"0E",X"E8",X"8E",X"23",X"40",X"FF",X"0E",X"EE",X"8E",
		X"64",X"E0",X"FF",X"00",X"EE",X"EE",X"64",X"E0",X"FF",X"00",X"0E",X"EE",X"54",X"00",X"FF",X"00",
		X"00",X"0C",X"C0",X"00",X"FF",X"05",X"50",X"00",X"00",X"FF",X"E5",X"55",X"52",X"00",X"FF",X"EE",
		X"54",X"55",X"20",X"FF",X"0E",X"8E",X"E5",X"30",X"FF",X"00",X"E8",X"E5",X"30",X"FF",X"00",X"EE",
		X"85",X"40",X"FF",X"00",X"0E",X"E5",X"40",X"FF",X"00",X"00",X"E5",X"55",X"FF",X"00",X"00",X"EE",
		X"50",X"FF",X"55",X"00",X"FF",X"E5",X"50",X"FF",X"E8",X"55",X"FF",X"0E",X"85",X"FF",X"00",X"E5",
		X"FF",X"00",X"00",X"05",X"04",X"00",X"00",X"FF",X"00",X"00",X"54",X"E4",X"40",X"00",X"FF",X"00",
		X"EE",X"43",X"E3",X"4E",X"00",X"FF",X"0E",X"A5",X"43",X"32",X"34",X"A0",X"FF",X"0E",X"E5",X"4E",
		X"1E",X"34",X"E0",X"FF",X"0E",X"55",X"6E",X"1E",X"64",X"50",X"FF",X"EE",X"57",X"EE",X"8E",X"E7",
		X"50",X"FF",X"EE",X"7E",X"E8",X"88",X"EE",X"70",X"FF",X"EE",X"EE",X"58",X"88",X"5E",X"E0",X"FF",
		X"0E",X"CC",X"EE",X"EE",X"EC",X"C0",X"FF",X"00",X"EE",X"EE",X"EE",X"EE",X"E0",X"FF",X"00",X"04",
		X"13",X"00",X"00",X"FF",X"00",X"45",X"E3",X"30",X"00",X"FF",X"04",X"5E",X"EE",X"33",X"00",X"FF",
		X"55",X"EE",X"8E",X"E4",X"40",X"FF",X"CC",X"E8",X"88",X"EC",X"C0",X"FF",X"EE",X"E8",X"88",X"EE",
		X"E0",X"FF",X"BB",X"EE",X"EE",X"EB",X"B0",X"FF",X"EE",X"00",X"00",X"0E",X"E0",X"FF",X"00",X"05",
		X"50",X"00",X"FF",X"00",X"5E",X"E5",X"00",X"FF",X"55",X"E8",X"8E",X"55",X"FF",X"BB",X"0E",X"E0",
		X"BB",X"FF",X"00",X"00",X"02",X"34",X"67",X"90",X"FF",X"00",X"00",X"01",X"33",X"58",X"70",X"FF",
		X"00",X"00",X"09",X"90",X"00",X"90",X"FF",X"00",X"0E",X"E7",X"B6",X"00",X"00",X"FF",X"00",X"ED",
		X"D4",X"B5",X"00",X"00",X"FF",X"00",X"ED",X"D4",X"B6",X"00",X"00",X"FF",X"00",X"0B",X"BB",X"B7",
		X"00",X"00",X"FF",X"8C",X"00",X"09",X"90",X"00",X"00",X"FF",X"CC",X"A9",X"87",X"43",X"00",X"00",
		X"FF",X"8B",X"06",X"97",X"63",X"00",X"00",X"FF",X"00",X"21",X"24",X"60",X"00",X"FF",X"00",X"21",
		X"24",X"60",X"00",X"FF",X"00",X"09",X"90",X"00",X"00",X"FF",X"00",X"07",X"B6",X"00",X"00",X"FF",
		X"0D",X"D4",X"B5",X"00",X"00",X"FF",X"ED",X"D4",X"B6",X"00",X"00",X"FF",X"EE",X"EB",X"B7",X"00",
		X"00",X"FF",X"8E",X"E9",X"90",X"00",X"00",X"FF",X"BC",X"98",X"23",X"00",X"00",X"FF",X"89",X"68",
		X"23",X"00",X"00",X"FF",X"00",X"07",X"32",X"40",X"00",X"00",X"FF",X"00",X"08",X"32",X"40",X"00",
		X"00",X"FF",X"00",X"0A",X"99",X"00",X"00",X"00",X"FF",X"0E",X"E6",X"7B",X"60",X"00",X"00",X"FF",
		X"EE",X"D6",X"4B",X"50",X"00",X"00",X"FF",X"EE",X"D6",X"4B",X"60",X"00",X"00",X"FF",X"0C",X"BB",
		X"BB",X"70",X"00",X"00",X"FF",X"00",X"0A",X"99",X"00",X"00",X"00",X"FF",X"00",X"08",X"32",X"40",
		X"00",X"00",X"FF",X"00",X"07",X"32",X"40",X"00",X"00",X"FF",X"8B",X"06",X"97",X"63",X"00",X"00",
		X"FF",X"CC",X"A9",X"87",X"43",X"00",X"00",X"FF",X"8C",X"00",X"09",X"90",X"00",X"00",X"FF",X"00",
		X"0D",X"D7",X"B7",X"00",X"00",X"FF",X"00",X"ED",X"D4",X"B6",X"00",X"00",X"FF",X"00",X"EE",X"E4",
		X"B5",X"00",X"00",X"FF",X"00",X"0C",X"CC",X"B6",X"00",X"00",X"FF",X"00",X"00",X"09",X"90",X"00",
		X"90",X"FF",X"00",X"00",X"01",X"33",X"58",X"70",X"FF",X"00",X"00",X"02",X"34",X"67",X"90",X"FF",
		X"89",X"68",X"23",X"00",X"00",X"FF",X"BC",X"98",X"23",X"00",X"00",X"FF",X"8E",X"E9",X"90",X"00",
		X"00",X"FF",X"ED",X"D7",X"B7",X"00",X"00",X"FF",X"ED",X"D4",X"B6",X"00",X"00",X"FF",X"0C",X"C4",
		X"B5",X"00",X"00",X"FF",X"00",X"0C",X"B6",X"00",X"00",X"FF",X"00",X"09",X"90",X"00",X"00",X"FF",
		X"00",X"21",X"24",X"60",X"00",X"FF",X"00",X"21",X"24",X"60",X"00",X"FF",X"8C",X"80",X"00",X"00",
		X"00",X"FF",X"CC",X"C0",X"00",X"00",X"00",X"FF",X"0C",X"00",X"00",X"00",X"00",X"FF",X"7A",X"00",
		X"E0",X"00",X"00",X"FF",X"89",X"0B",X"DD",X"00",X"00",X"FF",X"98",X"0B",X"DD",X"00",X"00",X"FF",
		X"77",X"9B",X"44",X"91",X"20",X"FF",X"64",X"9B",X"BB",X"93",X"30",X"FF",X"33",X"07",X"55",X"03",
		X"40",X"FF",X"00",X"00",X"00",X"06",X"70",X"FF",X"00",X"00",X"00",X"07",X"80",X"FF",X"00",X"00",
		X"00",X"08",X"70",X"FF",X"00",X"00",X"00",X"97",X"90",X"FF",X"8B",X"8E",X"00",X"00",X"00",X"FF",
		X"9C",X"ED",X"D0",X"00",X"00",X"FF",X"69",X"ED",X"D0",X"02",X"20",X"FF",X"88",X"96",X"47",X"91",
		X"10",X"FF",X"22",X"9B",X"BB",X"92",X"20",X"FF",X"33",X"07",X"65",X"04",X"40",X"FF",X"00",X"00",
		X"00",X"05",X"60",X"FF",X"00",X"00",X"00",X"06",X"60",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"E0",X"00",X"00",X"FF",X"00",X"0C",X"DD",X"00",X"00",X"FF",X"00",X"0B",X"DD",X"00",
		X"00",X"FF",X"77",X"AB",X"66",X"A7",X"70",X"FF",X"33",X"9B",X"44",X"93",X"30",X"FF",X"21",X"9B",
		X"BB",X"92",X"10",X"FF",X"33",X"07",X"65",X"03",X"30",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"8C",
		X"80",X"FF",X"00",X"00",X"00",X"CC",X"C0",X"FF",X"00",X"00",X"00",X"0C",X"00",X"FF",X"00",X"00",
		X"E0",X"0A",X"60",X"FF",X"00",X"0C",X"DD",X"09",X"70",X"FF",X"00",X"0C",X"DD",X"08",X"90",X"FF",
		X"21",X"9C",X"43",X"97",X"70",X"FF",X"33",X"9B",X"BB",X"94",X"50",X"FF",X"43",X"06",X"45",X"03",
		X"30",X"FF",X"65",X"00",X"00",X"00",X"00",X"FF",X"87",X"00",X"00",X"00",X"00",X"FF",X"68",X"00",
		X"00",X"00",X"00",X"FF",X"97",X"90",X"00",X"00",X"00",X"FF",X"00",X"00",X"0D",X"8C",X"80",X"FF",
		X"00",X"00",X"CD",X"DC",X"90",X"FF",X"22",X"00",X"CD",X"D9",X"60",X"FF",X"11",X"9C",X"44",X"97",
		X"80",X"FF",X"22",X"9B",X"BB",X"92",X"20",X"FF",X"44",X"06",X"56",X"03",X"30",X"FF",X"66",X"00",
		X"00",X"00",X"00",X"FF",X"66",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"53",X"33",X"35",X"00",X"FF",X"00",X"53",X"32",X"22",X"22",X"30",X"FF",X"05",X"33",
		X"22",X"21",X"12",X"25",X"FF",X"75",X"33",X"22",X"11",X"11",X"23",X"FF",X"75",X"33",X"22",X"11",
		X"11",X"23",X"FF",X"75",X"33",X"22",X"21",X"12",X"25",X"FF",X"75",X"53",X"32",X"22",X"22",X"35",
		X"FF",X"07",X"55",X"33",X"33",X"33",X"57",X"FF",X"00",X"75",X"55",X"55",X"55",X"70",X"FF",X"00",
		X"00",X"77",X"77",X"77",X"00",X"FF",X"00",X"53",X"33",X"35",X"00",X"FF",X"05",X"32",X"22",X"23",
		X"30",X"FF",X"53",X"22",X"11",X"12",X"35",X"FF",X"53",X"22",X"11",X"12",X"35",X"FF",X"53",X"22",
		X"11",X"12",X"35",X"FF",X"53",X"32",X"22",X"23",X"35",X"FF",X"75",X"33",X"33",X"33",X"57",X"FF",
		X"07",X"55",X"55",X"55",X"70",X"FF",X"00",X"77",X"77",X"77",X"00",X"FF",X"00",X"53",X"33",X"50",
		X"FF",X"05",X"33",X"22",X"35",X"FF",X"53",X"32",X"11",X"13",X"FF",X"53",X"22",X"11",X"13",X"FF",
		X"53",X"22",X"22",X"23",X"FF",X"53",X"32",X"22",X"35",X"FF",X"55",X"33",X"33",X"57",X"FF",X"05",
		X"55",X"55",X"50",X"FF",X"00",X"55",X"55",X"00",X"FF",X"00",X"00",X"00",X"05",X"33",X"50",X"FF",
		X"00",X"00",X"00",X"53",X"22",X"35",X"FF",X"00",X"00",X"00",X"32",X"21",X"23",X"FF",X"00",X"00",
		X"00",X"32",X"11",X"13",X"FF",X"00",X"00",X"00",X"32",X"21",X"23",X"FF",X"00",X"00",X"00",X"33",
		X"22",X"33",X"FF",X"00",X"00",X"00",X"53",X"33",X"35",X"FF",X"00",X"00",X"00",X"75",X"55",X"57",
		X"FF",X"04",X"40",X"00",X"07",X"77",X"70",X"FF",X"4E",X"E4",X"00",X"00",X"00",X"00",X"FF",X"EE",
		X"EE",X"00",X"00",X"00",X"00",X"FF",X"EE",X"EE",X"00",X"00",X"00",X"00",X"FF",X"4E",X"E4",X"00",
		X"00",X"00",X"00",X"FF",X"04",X"40",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"05",X"32",X"30",
		X"FF",X"00",X"00",X"53",X"22",X"23",X"FF",X"00",X"00",X"32",X"21",X"12",X"FF",X"00",X"00",X"32",
		X"21",X"12",X"FF",X"00",X"00",X"33",X"22",X"23",X"FF",X"00",X"00",X"53",X"33",X"33",X"FF",X"0E",
		X"EE",X"05",X"33",X"30",X"FF",X"EE",X"EE",X"E0",X"00",X"00",X"FF",X"EE",X"EE",X"E0",X"00",X"00",
		X"FF",X"EE",X"EE",X"E0",X"00",X"00",X"FF",X"0E",X"EE",X"00",X"00",X"00",X"FF",X"00",X"03",X"23",
		X"00",X"FF",X"00",X"32",X"21",X"30",X"FF",X"0E",X"32",X"21",X"20",X"FF",X"EE",X"33",X"22",X"30",
		X"FF",X"EE",X"33",X"33",X"30",X"FF",X"EE",X"E3",X"33",X"00",X"FF",X"EE",X"EE",X"E0",X"00",X"FF",
		X"0E",X"EE",X"00",X"00",X"FF",X"00",X"33",X"00",X"FF",X"03",X"32",X"30",X"FF",X"E3",X"32",X"30",
		X"FF",X"E5",X"33",X"50",X"FF",X"EE",X"55",X"00",X"FF",X"0E",X"E0",X"00",X"FF",X"03",X"02",X"00",
		X"FF",X"53",X"2C",X"20",X"FF",X"23",X"93",X"23",X"FF",X"53",X"02",X"50",X"FF",X"00",X"55",X"00",
		X"FF",X"00",X"20",X"20",X"FF",X"30",X"00",X"32",X"FF",X"30",X"91",X"03",X"FF",X"00",X"6C",X"00",
		X"FF",X"33",X"50",X"03",X"FF",X"03",X"05",X"22",X"FF",X"00",X"00",X"30",X"FF",X"00",X"00",X"10",
		X"00",X"FF",X"00",X"03",X"20",X"00",X"FF",X"00",X"00",X"00",X"31",X"FF",X"03",X"0A",X"A0",X"01",
		X"FF",X"33",X"0C",X"60",X"33",X"FF",X"30",X"01",X"90",X"21",X"FF",X"03",X"00",X"00",X"00",X"FF",
		X"35",X"30",X"33",X"30",X"FF",X"03",X"30",X"55",X"00",X"FF",X"00",X"00",X"00",X"11",X"00",X"FF",
		X"00",X"00",X"00",X"02",X"00",X"FF",X"03",X"30",X"00",X"00",X"00",X"FF",X"33",X"00",X"AA",X"00",
		X"22",X"FF",X"00",X"0D",X"69",X"D0",X"03",X"FF",X"00",X"0D",X"C1",X"D0",X"00",X"FF",X"33",X"00",
		X"BB",X"00",X"01",X"FF",X"35",X"50",X"00",X"00",X"32",X"FF",X"05",X"00",X"30",X"00",X"20",X"FF",
		X"00",X"05",X"50",X"00",X"00",X"FF",X"00",X"00",X"30",X"00",X"00",X"FF",X"00",X"20",X"00",X"02",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"20",X"08",
		X"AA",X"00",X"00",X"FF",X"00",X"08",X"11",X"B0",X"20",X"FF",X"50",X"0D",X"11",X"D0",X"00",X"FF",
		X"00",X"00",X"BB",X"D0",X"00",X"FF",X"00",X"50",X"00",X"00",X"00",X"FF",X"05",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"05",X"00",X"50",X"00",X"FF",X"12",X"3E",X"FF",X"45",X"67",X"FF",X"89",X"AB",
		X"FF",X"EC",X"D1",X"FF",X"88",X"88",X"80",X"FF",X"00",X"00",X"00",X"FF",X"88",X"88",X"80",X"FF",
		X"80",X"00",X"80",X"FF",X"88",X"88",X"80",X"FF",X"00",X"00",X"00",X"FF",X"88",X"88",X"80",X"FF",
		X"80",X"00",X"80",X"FF",X"88",X"88",X"80",X"FF",X"00",X"00",X"00",X"FF",X"88",X"88",X"80",X"FF",
		X"80",X"00",X"80",X"FF",X"88",X"88",X"80",X"FF",X"00",X"00",X"00",X"FF",X"88",X"88",X"80",X"FF",
		X"80",X"00",X"80",X"FF",X"88",X"88",X"80",X"FF",X"88",X"88",X"80",X"FF",X"00",X"00",X"00",X"FF",
		X"88",X"88",X"80",X"FF",X"80",X"00",X"80",X"FF",X"88",X"88",X"80",X"FF",X"00",X"00",X"00",X"FF",
		X"88",X"88",X"80",X"FF",X"80",X"00",X"80",X"FF",X"88",X"88",X"80",X"FF",X"88",X"80",X"80",X"FF",
		X"80",X"88",X"80",X"FF",X"00",X"00",X"00",X"FF",X"88",X"88",X"80",X"FF",X"80",X"00",X"80",X"FF",
		X"88",X"88",X"80",X"FF",X"00",X"00",X"00",X"FF",X"88",X"88",X"80",X"FF",X"80",X"00",X"80",X"FF",
		X"88",X"88",X"80",X"FF",X"80",X"80",X"80",X"FF",X"88",X"88",X"80",X"FF",X"00",X"00",X"00",X"FF",
		X"88",X"88",X"80",X"FF",X"80",X"00",X"80",X"FF",X"88",X"88",X"80",X"FF",X"00",X"00",X"00",X"FF",
		X"88",X"88",X"80",X"FF",X"80",X"00",X"80",X"FF",X"88",X"88",X"80",X"FF",X"08",X"88",X"80",X"FF",
		X"08",X"00",X"00",X"FF",X"88",X"88",X"80",X"FF",X"00",X"00",X"00",X"FF",X"88",X"88",X"80",X"FF",
		X"80",X"00",X"80",X"FF",X"88",X"88",X"80",X"FF",X"00",X"00",X"00",X"FF",X"88",X"88",X"80",X"FF",
		X"80",X"00",X"80",X"FF",X"88",X"88",X"80",X"FF",X"80",X"88",X"80",X"FF",X"88",X"80",X"80",X"FF",
		X"00",X"00",X"00",X"FF",X"88",X"88",X"80",X"FF",X"80",X"00",X"80",X"FF",X"88",X"88",X"80",X"FF",
		X"00",X"00",X"00",X"FF",X"88",X"88",X"80",X"FF",X"80",X"00",X"80",X"FF",X"88",X"88",X"80",X"FF",
		X"88",X"88",X"80",X"FF",X"80",X"80",X"80",X"FF",X"88",X"80",X"80",X"FF",X"00",X"00",X"00",X"FF",
		X"88",X"88",X"80",X"FF",X"80",X"00",X"80",X"FF",X"88",X"88",X"80",X"FF",X"00",X"00",X"00",X"FF",
		X"88",X"88",X"80",X"FF",X"80",X"00",X"80",X"FF",X"88",X"88",X"80",X"FF",X"88",X"88",X"80",X"FF",
		X"80",X"80",X"80",X"FF",X"88",X"88",X"80",X"FF",X"00",X"00",X"00",X"FF",X"88",X"88",X"80",X"FF",
		X"80",X"00",X"80",X"FF",X"88",X"88",X"80",X"FF",X"00",X"00",X"00",X"FF",X"88",X"88",X"80",X"FF",
		X"80",X"00",X"80",X"FF",X"88",X"88",X"80",X"FF",X"88",X"88",X"80",X"FF",X"00",X"00",X"00",X"FF",
		X"88",X"88",X"80",X"FF",X"80",X"00",X"80",X"FF",X"88",X"88",X"80",X"FF",X"00",X"00",X"00",X"FF",
		X"88",X"88",X"80",X"FF",X"80",X"00",X"80",X"FF",X"88",X"88",X"80",X"FF",X"00",X"00",X"00",X"FF",
		X"88",X"88",X"80",X"FF",X"80",X"00",X"80",X"FF",X"88",X"88",X"80",X"FF",X"88",X"88",X"80",X"FF",
		X"00",X"00",X"00",X"FF",X"88",X"80",X"80",X"FF",X"80",X"88",X"80",X"FF",X"00",X"00",X"00",X"FF",
		X"88",X"88",X"80",X"FF",X"80",X"00",X"80",X"FF",X"88",X"88",X"80",X"FF",X"00",X"00",X"00",X"FF",
		X"88",X"88",X"80",X"FF",X"80",X"00",X"80",X"FF",X"88",X"88",X"80",X"FF",X"88",X"88",X"80",X"FF",
		X"00",X"00",X"00",X"FF",X"80",X"88",X"80",X"FF",X"88",X"80",X"80",X"FF",X"00",X"00",X"00",X"FF",
		X"88",X"88",X"80",X"FF",X"80",X"00",X"80",X"FF",X"88",X"88",X"80",X"FF",X"00",X"00",X"00",X"FF",
		X"88",X"88",X"80",X"FF",X"80",X"00",X"80",X"FF",X"88",X"88",X"80",X"FF",X"88",X"88",X"80",X"FF",
		X"00",X"00",X"00",X"FF",X"88",X"88",X"80",X"FF",X"80",X"80",X"80",X"FF",X"88",X"80",X"80",X"FF",
		X"00",X"00",X"00",X"FF",X"88",X"88",X"80",X"FF",X"80",X"00",X"80",X"FF",X"88",X"88",X"80",X"FF",
		X"00",X"00",X"00",X"FF",X"88",X"88",X"80",X"FF",X"80",X"00",X"80",X"FF",X"88",X"88",X"80",X"FF",
		X"88",X"80",X"80",X"FF",X"80",X"88",X"80",X"FF",X"00",X"00",X"00",X"FF",X"88",X"88",X"80",X"FF",
		X"80",X"00",X"80",X"FF",X"88",X"88",X"80",X"FF",X"00",X"00",X"00",X"FF",X"88",X"88",X"80",X"FF",
		X"80",X"00",X"80",X"FF",X"88",X"88",X"80",X"FF",X"00",X"00",X"00",X"FF",X"88",X"88",X"80",X"FF",
		X"80",X"00",X"80",X"FF",X"88",X"88",X"80",X"FF",X"88",X"80",X"80",X"FF",X"80",X"88",X"80",X"FF",
		X"00",X"00",X"00",X"FF",X"08",X"88",X"80",X"FF",X"08",X"00",X"00",X"FF",X"88",X"88",X"80",X"FF",
		X"00",X"00",X"00",X"FF",X"88",X"88",X"80",X"FF",X"80",X"00",X"80",X"FF",X"88",X"88",X"80",X"FF",
		X"00",X"00",X"00",X"FF",X"88",X"88",X"80",X"FF",X"80",X"00",X"80",X"FF",X"88",X"88",X"80",X"FF",
		X"80",X"80",X"80",X"FF",X"88",X"88",X"80",X"FF",X"00",X"00",X"00",X"FF",X"88",X"88",X"80",X"FF",
		X"80",X"00",X"80",X"FF",X"88",X"88",X"80",X"FF",X"00",X"00",X"00",X"FF",X"88",X"88",X"80",X"FF",
		X"80",X"00",X"80",X"FF",X"88",X"88",X"80",X"FF",X"00",X"00",X"00",X"FF",X"88",X"88",X"80",X"FF",
		X"80",X"00",X"80",X"FF",X"88",X"88",X"80",X"FF",X"80",X"80",X"80",X"FF",X"88",X"88",X"80",X"FF",
		X"00",X"00",X"00",X"FF",X"88",X"80",X"80",X"FF",X"80",X"88",X"80",X"FF",X"00",X"00",X"00",X"FF",
		X"88",X"88",X"80",X"FF",X"80",X"00",X"80",X"FF",X"88",X"88",X"80",X"FF",X"00",X"00",X"00",X"FF",
		X"88",X"88",X"80",X"FF",X"80",X"00",X"80",X"FF",X"88",X"88",X"80",X"FF",X"80",X"88",X"80",X"FF",
		X"88",X"80",X"80",X"FF",X"00",X"00",X"00",X"FF",X"88",X"88",X"80",X"FF",X"80",X"00",X"80",X"FF",
		X"88",X"88",X"80",X"FF",X"00",X"00",X"00",X"FF",X"88",X"88",X"80",X"FF",X"80",X"00",X"80",X"FF",
		X"88",X"88",X"80",X"FF",X"00",X"00",X"00",X"FF",X"88",X"88",X"80",X"FF",X"80",X"00",X"80",X"FF",
		X"88",X"88",X"80",X"FF",X"88",X"88",X"80",X"FF",X"80",X"80",X"80",X"FF",X"88",X"80",X"80",X"FF",
		X"00",X"00",X"00",X"FF",X"08",X"88",X"80",X"FF",X"08",X"00",X"00",X"FF",X"88",X"88",X"80",X"FF",
		X"00",X"00",X"00",X"FF",X"88",X"88",X"80",X"FF",X"80",X"00",X"80",X"FF",X"88",X"88",X"80",X"FF",
		X"00",X"00",X"00",X"FF",X"88",X"88",X"80",X"FF",X"80",X"00",X"80",X"FF",X"88",X"88",X"80",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"10",X"00",X"FF",X"00",X"00",X"00",X"10",
		X"00",X"11",X"01",X"00",X"11",X"00",X"00",X"FF",X"00",X"00",X"10",X"11",X"10",X"11",X"00",X"00",
		X"11",X"00",X"00",X"FF",X"00",X"00",X"10",X"11",X"10",X"00",X"10",X"00",X"10",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"02",X"20",X"00",X"00",X"FF",X"00",X"01",X"02",X"00",
		X"10",X"01",X"10",X"13",X"10",X"01",X"00",X"FF",X"11",X"00",X"00",X"20",X"01",X"00",X"11",X"33",
		X"01",X"00",X"10",X"FF",X"11",X"00",X"00",X"12",X"10",X"11",X"11",X"14",X"00",X"00",X"01",X"FF",
		X"00",X"11",X"10",X"10",X"21",X"12",X"11",X"41",X"00",X"11",X"00",X"FF",X"00",X"01",X"20",X"11",
		X"00",X"11",X"11",X"01",X"22",X"10",X"40",X"FF",X"11",X"01",X"02",X"11",X"21",X"14",X"41",X"11",
		X"31",X"21",X"00",X"FF",X"00",X"00",X"00",X"31",X"21",X"11",X"50",X"11",X"41",X"55",X"13",X"FF",
		X"00",X"11",X"00",X"00",X"11",X"16",X"11",X"51",X"11",X"05",X"10",X"FF",X"0D",X"D0",X"01",X"D1",
		X"01",X"4B",X"11",X"15",X"0D",X"50",X"00",X"FF",X"00",X"00",X"1D",X"11",X"1B",X"10",X"10",X"61",
		X"00",X"01",X"00",X"FF",X"00",X"00",X"00",X"01",X"10",X"01",X"15",X"03",X"11",X"00",X"00",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"09",X"00",X"FF",X"75",X"A0",X"FF",X"09",X"00",X"FF",X"09",X"00",X"FF",X"79",X"A0",X"FF",X"64",
		X"90",X"FF",X"56",X"70",X"FF",X"06",X"00",X"FF",X"09",X"AA",X"00",X"FF",X"99",X"A9",X"90",X"FF",
		X"79",X"A9",X"90",X"FF",X"77",X"47",X"70",X"FF",X"66",X"56",X"70",X"FF",X"66",X"56",X"60",X"FF",
		X"05",X"56",X"00",X"FF",X"00",X"A9",X"9E",X"00",X"FF",X"0A",X"A9",X"99",X"E0",X"FF",X"0A",X"A9",
		X"97",X"E0",X"FF",X"9A",X"A9",X"77",X"7E",X"FF",X"99",X"93",X"66",X"6E",X"FF",X"99",X"76",X"56",
		X"6E",X"FF",X"07",X"76",X"55",X"E0",X"FF",X"07",X"76",X"55",X"E0",X"FF",X"00",X"66",X"5E",X"00",
		X"FF",X"00",X"09",X"97",X"EE",X"00",X"FF",X"00",X"99",X"77",X"7E",X"E0",X"FF",X"0A",X"99",X"77",
		X"77",X"EB",X"FF",X"0A",X"99",X"77",X"77",X"AE",X"FF",X"AA",X"A9",X"76",X"66",X"6E",X"FF",X"AA",
		X"AA",X"15",X"56",X"6E",X"FF",X"99",X"99",X"75",X"55",X"9E",X"FF",X"09",X"97",X"76",X"55",X"E0",
		X"FF",X"09",X"77",X"76",X"69",X"E0",X"FF",X"00",X"77",X"76",X"6E",X"00",X"FF",X"00",X"07",X"76",
		X"E0",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"0C",X"CC",X"EE",X"00",X"00",X"FF",X"00",X"09",X"77",X"6E",X"E0",X"00",X"FF",X"00",
		X"97",X"76",X"66",X"EE",X"00",X"FF",X"09",X"97",X"76",X"66",X"6E",X"B0",X"FF",X"09",X"97",X"76",
		X"66",X"6A",X"E0",X"FF",X"99",X"99",X"76",X"55",X"55",X"E0",X"FF",X"99",X"99",X"91",X"66",X"55",
		X"E0",X"FF",X"99",X"99",X"A9",X"66",X"65",X"E0",X"FF",X"0A",X"AA",X"99",X"76",X"6B",X"00",X"FF",
		X"0A",X"A9",X"99",X"77",X"6E",X"00",X"FF",X"00",X"99",X"99",X"77",X"E0",X"00",X"FF",X"00",X"09",
		X"97",X"7E",X"00",X"00",X"FF",X"00",X"0D",X"DD",X"E0",X"00",X"00",X"FF",X"00",X"00",X"CC",X"CE",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"0C",X"CC",X"E0",X"00",X"00",X"FF",X"00",X"00",X"00",X"DD",X"DE",X"00",
		X"00",X"FF",X"00",X"0A",X"E9",X"66",X"5E",X"E0",X"00",X"FF",X"00",X"AE",X"76",X"65",X"55",X"EE",
		X"00",X"FF",X"0A",X"E7",X"76",X"65",X"55",X"9E",X"B0",X"FF",X"AA",X"E7",X"76",X"65",X"56",X"6E",
		X"E0",X"FF",X"AE",X"77",X"77",X"65",X"66",X"6A",X"E0",X"FF",X"0E",X"97",X"77",X"71",X"77",X"69",
		X"E0",X"FF",X"AE",X"99",X"99",X"9A",X"97",X"7A",X"E0",X"FF",X"AA",X"E9",X"99",X"AA",X"99",X"9E",
		X"00",X"FF",X"0A",X"E9",X"9A",X"AA",X"99",X"AE",X"00",X"FF",X"00",X"AE",X"AA",X"AA",X"99",X"E0",
		X"00",X"FF",X"00",X"0A",X"EA",X"A9",X"9E",X"00",X"00",X"FF",X"00",X"00",X"0D",X"DD",X"E0",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"DD",X"DE",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"CE",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"0C",X"CC",X"CE",X"00",X"00",X"FF",X"00",X"09",X"E6",X"55",X"6B",X"E0",
		X"00",X"FF",X"00",X"9E",X"65",X"56",X"66",X"BE",X"00",X"FF",X"09",X"E6",X"65",X"56",X"66",X"6E",
		X"00",X"FF",X"99",X"E6",X"65",X"56",X"67",X"7E",X"E0",X"FF",X"9E",X"66",X"66",X"56",X"77",X"7B",
		X"E0",X"FF",X"0E",X"76",X"66",X"61",X"99",X"7A",X"E0",X"FF",X"9E",X"77",X"77",X"79",X"A9",X"9B",
		X"E0",X"FF",X"99",X"E7",X"77",X"99",X"AA",X"9E",X"00",X"FF",X"09",X"E7",X"79",X"99",X"AA",X"BE",
		X"00",X"FF",X"00",X"AE",X"99",X"99",X"AB",X"E0",X"00",X"FF",X"00",X"09",X"E9",X"9A",X"BE",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"DD",X"E0",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"CC",X"CE",X"00",X"00",X"FF",X"00",X"00",X"0D",X"DD",X"EE",X"00",
		X"00",X"FF",X"00",X"09",X"E6",X"55",X"6B",X"E0",X"00",X"FF",X"00",X"9E",X"65",X"56",X"66",X"BE",
		X"00",X"FF",X"09",X"E6",X"65",X"56",X"66",X"6E",X"00",X"FF",X"99",X"E6",X"65",X"56",X"67",X"7E",
		X"E0",X"FF",X"9E",X"66",X"66",X"56",X"77",X"7B",X"E0",X"FF",X"0E",X"76",X"66",X"61",X"99",X"7A",
		X"E0",X"FF",X"9E",X"77",X"77",X"79",X"A9",X"9B",X"E0",X"FF",X"99",X"E7",X"77",X"99",X"AA",X"9E",
		X"00",X"FF",X"09",X"E7",X"79",X"99",X"AA",X"BE",X"00",X"FF",X"00",X"AE",X"99",X"99",X"AB",X"E0",
		X"00",X"FF",X"00",X"09",X"E9",X"9A",X"BE",X"00",X"00",X"FF",X"00",X"00",X"0D",X"DD",X"E0",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"DD",X"DE",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"CC",X"CE",X"00",X"00",X"FF",X"00",X"00",X"00",X"DD",X"DE",X"00",
		X"00",X"FF",X"00",X"00",X"0D",X"DD",X"EE",X"00",X"00",X"FF",X"00",X"06",X"E6",X"77",X"9E",X"E0",
		X"00",X"FF",X"00",X"6E",X"67",X"77",X"99",X"EB",X"00",X"FF",X"06",X"E6",X"67",X"79",X"99",X"AE",
		X"00",X"FF",X"66",X"E6",X"67",X"79",X"99",X"9B",X"E0",X"FF",X"6E",X"66",X"66",X"79",X"AA",X"AB",
		X"E0",X"FF",X"0E",X"56",X"66",X"61",X"99",X"9A",X"E0",X"FF",X"6E",X"55",X"55",X"56",X"79",X"9B",
		X"E0",X"FF",X"66",X"E5",X"55",X"66",X"77",X"9E",X"00",X"FF",X"06",X"E5",X"56",X"66",X"77",X"BE",
		X"00",X"FF",X"00",X"6E",X"66",X"66",X"79",X"E0",X"00",X"FF",X"00",X"06",X"E6",X"67",X"9E",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"DD",X"DE",X"E0",X"00",X"FF",X"00",X"00",X"00",X"0D",X"DC",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"CC",X"E0",X"00",
		X"00",X"FF",X"00",X"00",X"0D",X"DD",X"E0",X"00",X"00",X"FF",X"00",X"00",X"0D",X"DD",X"EE",X"00",
		X"00",X"FF",X"00",X"07",X"E7",X"99",X"9E",X"E0",X"00",X"FF",X"00",X"7E",X"79",X"99",X"AA",X"EB",
		X"00",X"FF",X"07",X"E7",X"79",X"9A",X"AA",X"BE",X"00",X"FF",X"77",X"E7",X"79",X"9A",X"AA",X"AB",
		X"E0",X"FF",X"7E",X"77",X"77",X"9A",X"99",X"9B",X"E0",X"FF",X"0E",X"67",X"77",X"71",X"77",X"9A",
		X"E0",X"FF",X"7E",X"66",X"66",X"65",X"67",X"7B",X"E0",X"FF",X"77",X"E6",X"66",X"55",X"66",X"7E",
		X"00",X"FF",X"07",X"E6",X"65",X"55",X"66",X"AE",X"00",X"FF",X"00",X"7E",X"55",X"55",X"66",X"E0",
		X"00",X"FF",X"00",X"07",X"E5",X"56",X"6E",X"00",X"00",X"FF",X"00",X"00",X"0D",X"CC",X"E0",X"00",
		X"00",X"FF",X"00",X"00",X"0D",X"CC",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"FF",X"00",X"00",X"00",X"0D",X"DE",X"00",
		X"00",X"FF",X"00",X"00",X"0D",X"DD",X"EE",X"00",X"00",X"FF",X"00",X"09",X"E6",X"55",X"6B",X"E0",
		X"00",X"FF",X"00",X"9E",X"65",X"56",X"66",X"BE",X"00",X"FF",X"09",X"E6",X"65",X"56",X"66",X"6E",
		X"00",X"FF",X"99",X"E6",X"65",X"56",X"67",X"7E",X"E0",X"FF",X"9E",X"66",X"66",X"56",X"77",X"7B",
		X"E0",X"FF",X"0E",X"76",X"66",X"61",X"99",X"7A",X"E0",X"FF",X"9E",X"77",X"77",X"79",X"A9",X"9B",
		X"E0",X"FF",X"99",X"E7",X"77",X"99",X"AA",X"9E",X"00",X"FF",X"09",X"E7",X"79",X"99",X"AA",X"BE",
		X"00",X"FF",X"00",X"AE",X"99",X"99",X"AB",X"E0",X"00",X"FF",X"00",X"09",X"E9",X"9A",X"BE",X"00",
		X"00",X"FF",X"00",X"00",X"0D",X"DD",X"E0",X"00",X"00",X"FF",X"00",X"00",X"0C",X"CC",X"E0",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"DC",X"CE",X"00",X"00",X"FF",X"00",X"0E",X"DD",X"E0",X"00",X"00",X"FF",X"00",
		X"0E",X"DD",X"EE",X"00",X"00",X"FF",X"00",X"9A",X"DB",X"9E",X"00",X"00",X"FF",X"09",X"7E",X"75",
		X"3B",X"00",X"00",X"FF",X"77",X"E7",X"75",X"97",X"90",X"00",X"FF",X"68",X"E7",X"59",X"77",X"3B",
		X"00",X"FF",X"EE",X"E7",X"59",X"75",X"99",X"10",X"FF",X"75",X"E7",X"59",X"75",X"99",X"00",X"FF",
		X"97",X"EB",X"59",X"99",X"6E",X"E0",X"FF",X"09",X"7E",X"B6",X"9A",X"EE",X"00",X"FF",X"00",X"AA",
		X"DB",X"BE",X"E0",X"00",X"FF",X"00",X"0E",X"DD",X"EE",X"E0",X"00",X"FF",X"00",X"0E",X"DD",X"DE",
		X"00",X"00",X"FF",X"00",X"00",X"0C",X"CE",X"E0",X"00",X"FF",X"00",X"00",X"0C",X"0E",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"0C",X"CD",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"08",X"E4",X"EC",X"7D",X"D0",X"00",X"00",X"00",X"00",X"FF",X"08",
		X"E4",X"E7",X"ED",X"D0",X"00",X"00",X"00",X"00",X"FF",X"08",X"EA",X"A9",X"AD",X"59",X"00",X"00",
		X"00",X"00",X"FF",X"0E",X"A9",X"99",X"9E",X"97",X"57",X"00",X"00",X"00",X"FF",X"EA",X"97",X"75",
		X"5E",X"75",X"77",X"75",X"00",X"00",X"FF",X"EA",X"97",X"44",X"5E",X"47",X"97",X"57",X"70",X"00",
		X"FF",X"EE",X"EE",X"EE",X"EE",X"49",X"95",X"97",X"9A",X"10",X"FF",X"EA",X"96",X"55",X"5E",X"59",
		X"7A",X"99",X"A0",X"00",X"FF",X"EA",X"97",X"66",X"7E",X"97",X"A9",X"9A",X"E0",X"00",X"FF",X"EE",
		X"A9",X"99",X"9E",X"99",X"AA",X"EE",X"EE",X"00",X"FF",X"EE",X"8A",X"AA",X"AD",X"AA",X"EE",X"EE",
		X"E0",X"00",X"FF",X"EE",X"8E",X"4E",X"7D",X"EE",X"CE",X"E0",X"00",X"00",X"FF",X"EE",X"8E",X"4E",
		X"7D",X"DC",X"C0",X"00",X"00",X"00",X"FF",X"EE",X"EE",X"EE",X"EE",X"DE",X"00",X"00",X"00",X"00",
		X"FF",X"0E",X"EE",X"EE",X"EE",X"E0",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0C",X"C0",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0E",X"C0",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"ED",X"D0",X"00",X"00",X"00",X"00",X"FF",X"00",X"8E",X"7E",X"4D",X"D0",X"00",X"00",
		X"00",X"00",X"FF",X"0E",X"8E",X"7E",X"4D",X"D0",X"00",X"00",X"00",X"00",X"FF",X"0E",X"8B",X"AA",
		X"AD",X"B7",X"00",X"00",X"00",X"00",X"FF",X"0E",X"A9",X"99",X"9E",X"59",X"77",X"00",X"00",X"00",
		X"FF",X"0A",X"97",X"75",X"5E",X"95",X"57",X"75",X"00",X"00",X"FF",X"E9",X"75",X"43",X"2E",X"44",
		X"75",X"59",X"70",X"00",X"FF",X"EE",X"EE",X"EE",X"EE",X"47",X"44",X"75",X"57",X"10",X"FF",X"E9",
		X"76",X"55",X"5E",X"97",X"47",X"44",X"70",X"00",X"FF",X"EA",X"97",X"66",X"5E",X"75",X"97",X"47",
		X"E0",X"00",X"FF",X"EE",X"A9",X"99",X"9E",X"59",X"95",X"EE",X"EE",X"00",X"FF",X"E5",X"EB",X"AA",
		X"AD",X"BA",X"EE",X"EE",X"E0",X"00",X"FF",X"E5",X"E7",X"E8",X"ED",X"DE",X"EE",X"E0",X"00",X"00",
		X"FF",X"E5",X"E7",X"E8",X"ED",X"DD",X"CC",X"00",X"00",X"00",X"FF",X"EE",X"EE",X"EE",X"EE",X"DD",
		X"C0",X"00",X"00",X"00",X"FF",X"0E",X"EE",X"EE",X"E0",X"EE",X"EE",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"D0",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0D",X"DD",X"00",X"00",X"00",X"00",
		X"FF",X"07",X"E8",X"E4",X"ED",X"DD",X"C0",X"00",X"00",X"00",X"FF",X"07",X"E8",X"E4",X"ED",X"D0",
		X"CC",X"00",X"00",X"00",X"FF",X"07",X"EB",X"AA",X"AE",X"B7",X"00",X"00",X"00",X"00",X"FF",X"0E",
		X"A9",X"99",X"9E",X"7A",X"9A",X"00",X"00",X"00",X"FF",X"0A",X"97",X"75",X"5E",X"99",X"75",X"AA",
		X"00",X"00",X"FF",X"EA",X"95",X"52",X"4E",X"75",X"59",X"A9",X"70",X"00",X"FF",X"EE",X"EE",X"EE",
		X"EE",X"54",X"79",X"75",X"99",X"10",X"FF",X"EA",X"96",X"64",X"6E",X"47",X"77",X"57",X"90",X"00",
		X"FF",X"EA",X"97",X"66",X"7E",X"97",X"54",X"79",X"E0",X"00",X"FF",X"EE",X"A9",X"99",X"9E",X"75",
		X"49",X"EE",X"EE",X"00",X"FF",X"EE",X"7B",X"AA",X"AE",X"B5",X"EE",X"EE",X"E0",X"00",X"FF",X"EE",
		X"7E",X"8E",X"DD",X"EE",X"EE",X"E0",X"00",X"00",X"FF",X"EE",X"7E",X"8E",X"DD",X"EE",X"E0",X"00",
		X"00",X"00",X"FF",X"0E",X"EE",X"EE",X"DE",X"E0",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"0E",
		X"DD",X"C0",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"0E",X"ED",X"C0",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"DD",X"DC",X"00",X"00",X"00",X"FF",X"0A",
		X"EC",X"E4",X"ED",X"DD",X"DC",X"C0",X"00",X"00",X"FF",X"0A",X"EC",X"E4",X"ED",X"D0",X"00",X"00",
		X"00",X"00",X"FF",X"0A",X"EB",X"AA",X"AD",X"B9",X"00",X"00",X"00",X"00",X"FF",X"00",X"A9",X"99",
		X"9E",X"A9",X"A9",X"00",X"00",X"00",X"FF",X"0A",X"97",X"76",X"5E",X"9A",X"AA",X"9A",X"00",X"00",
		X"FF",X"EA",X"93",X"34",X"5E",X"AA",X"A7",X"AA",X"A0",X"00",X"FF",X"EE",X"EE",X"EE",X"EE",X"AA",
		X"7A",X"AA",X"7A",X"10",X"FF",X"EA",X"75",X"56",X"6E",X"AA",X"7A",X"A7",X"A0",X"00",X"FF",X"EA",
		X"97",X"76",X"6E",X"A7",X"6A",X"A6",X"E0",X"00",X"FF",X"EE",X"A9",X"99",X"9E",X"A6",X"A9",X"EE",
		X"EE",X"00",X"FF",X"EA",X"EB",X"AA",X"AD",X"BB",X"EE",X"EE",X"E0",X"00",X"FF",X"EA",X"E8",X"E4",
		X"DD",X"EE",X"EE",X"E0",X"00",X"00",X"FF",X"EA",X"E8",X"E4",X"DD",X"EE",X"E0",X"00",X"00",X"00",
		X"FF",X"EE",X"EE",X"EC",X"DD",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"EE",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"90",X"70",X"00",X"00",X"FF",X"00",X"00",X"09",
		X"6E",X"57",X"00",X"00",X"FF",X"00",X"00",X"99",X"4E",X"14",X"70",X"00",X"FF",X"00",X"EE",X"AE",
		X"EE",X"EE",X"AE",X"E0",X"FF",X"00",X"ED",X"DB",X"99",X"7B",X"DD",X"D0",X"FF",X"0D",X"DD",X"B9",
		X"99",X"57",X"BD",X"DD",X"FF",X"EC",X"CE",X"A9",X"AA",X"A5",X"9E",X"DD",X"FF",X"ED",X"CE",X"AB",
		X"99",X"A5",X"9E",X"C0",X"FF",X"EE",X"CE",X"E9",X"99",X"7A",X"00",X"00",X"FF",X"0E",X"00",X"EB",
		X"AA",X"5A",X"00",X"00",X"FF",X"00",X"00",X"EE",X"A9",X"B0",X"00",X"00",X"FF",X"00",X"00",X"0E",
		X"08",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0E",X"EE",X"E0",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"EE",X"EE",X"9E",X"9E",X"E0",X"00",X"00",X"FF",X"00",X"0E",X"88",X"E9",X"7E",X"7A",X"E8",
		X"80",X"00",X"FF",X"00",X"0E",X"EE",X"B9",X"6E",X"57",X"BE",X"E0",X"00",X"FF",X"00",X"0E",X"44",
		X"97",X"6E",X"57",X"A4",X"40",X"00",X"FF",X"00",X"0E",X"EE",X"96",X"5E",X"45",X"AE",X"EE",X"E0",
		X"FF",X"00",X"0E",X"77",X"95",X"5E",X"45",X"A7",X"CC",X"C0",X"FF",X"0E",X"EE",X"EE",X"95",X"5E",
		X"34",X"AE",X"EC",X"C0",X"FF",X"EE",X"DE",X"DD",X"EE",X"EE",X"EE",X"DD",X"ED",X"C0",X"FF",X"ED",
		X"DE",X"DD",X"BA",X"A5",X"7A",X"BD",X"DD",X"00",X"FF",X"0E",X"DD",X"EE",X"A9",X"9A",X"55",X"A0",
		X"00",X"00",X"FF",X"00",X"EC",X"CE",X"9A",X"77",X"A4",X"50",X"00",X"00",X"FF",X"00",X"0E",X"CE",
		X"A7",X"A5",X"5A",X"50",X"00",X"00",X"FF",X"00",X"00",X"0E",X"EA",X"7A",X"45",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"0E",X"EA",X"75",X"A5",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"E9",X"A4",
		X"5A",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"EE",X"7A",X"50",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"0E",X"96",X"A0",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0E",X"03",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"EE",X"E0",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0E",X"AE",X"A0",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"0E",X"EE",X"EA",X"9E",X"9A",X"E4",X"40",X"00",X"00",X"FF",X"00",X"0E",
		X"44",X"A9",X"7E",X"77",X"AE",X"E0",X"00",X"00",X"FF",X"00",X"0E",X"EE",X"A9",X"7E",X"77",X"A7",
		X"70",X"00",X"00",X"FF",X"00",X"0E",X"77",X"A9",X"5E",X"56",X"AE",X"E0",X"00",X"00",X"FF",X"00",
		X"0E",X"EE",X"A7",X"5E",X"46",X"A8",X"80",X"00",X"00",X"FF",X"00",X"EE",X"88",X"A7",X"5E",X"45",
		X"AE",X"EE",X"EE",X"00",X"FF",X"0E",X"ED",X"DD",X"DE",X"EE",X"EE",X"DD",X"DD",X"DD",X"E0",X"FF",
		X"0E",X"DD",X"DD",X"B7",X"53",X"59",X"BD",X"DD",X"DC",X"C0",X"FF",X"0E",X"DD",X"0E",X"96",X"77",
		X"35",X"90",X"00",X"EC",X"00",X"FF",X"0E",X"DD",X"0E",X"A9",X"55",X"75",X"70",X"00",X"00",X"00",
		X"FF",X"0E",X"CC",X"0E",X"E7",X"73",X"57",X"00",X"00",X"00",X"00",X"FF",X"00",X"EC",X"00",X"E6",
		X"57",X"37",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"E7",X"55",X"95",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"EE",X"73",X"50",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"0E",X"57",X"50",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0E",X"05",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"0E",X"EE",X"EA",X"EA",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"E7",X"7E",X"AA",X"EA",X"AE",X"EE",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"EE",X"EA",X"A9",X"E9",X"AA",X"77",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"E8",X"8A",X"97",X"E5",X"7A",X"EE",X"00",X"00",X"00",X"FF",X"00",X"00",X"EE",X"EA",X"65",X"E4",
		X"6A",X"88",X"00",X"00",X"00",X"FF",X"00",X"EE",X"E4",X"4A",X"65",X"E3",X"6A",X"EE",X"00",X"00",
		X"00",X"FF",X"EE",X"ED",X"DD",X"DA",X"75",X"E4",X"5A",X"44",X"EE",X"00",X"00",X"FF",X"EC",X"DD",
		X"DD",X"DD",X"EE",X"EE",X"ED",X"DD",X"DD",X"E0",X"00",X"FF",X"0C",X"C0",X"00",X"EB",X"54",X"97",
		X"AB",X"DD",X"DD",X"D0",X"00",X"FF",X"00",X"00",X"00",X"E9",X"A4",X"59",X"9A",X"EE",X"DD",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"E7",X"79",X"56",X"99",X"EC",X"C0",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"EE",X"57",X"95",X"70",X"0C",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0E",X"55",X"9A",
		X"70",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0E",X"A5",X"79",X"A0",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"0E",X"EA",X"5A",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"E9",X"A7",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"E0",X"90",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"FF",X"00",X"0E",X"EE",X"EA",X"EA",
		X"E0",X"00",X"00",X"FF",X"00",X"E9",X"9E",X"AA",X"EA",X"AE",X"99",X"00",X"FF",X"00",X"EE",X"EA",
		X"A9",X"E9",X"AA",X"EE",X"00",X"FF",X"00",X"EC",X"CA",X"97",X"E5",X"9A",X"CC",X"00",X"FF",X"EE",
		X"EE",X"EA",X"75",X"E3",X"6A",X"EE",X"00",X"FF",X"EC",X"E4",X"4A",X"65",X"E4",X"6A",X"44",X"00",
		X"FF",X"ED",X"DD",X"DA",X"65",X"E5",X"6A",X"EE",X"E0",X"FF",X"0E",X"DD",X"DD",X"EE",X"EE",X"ED",
		X"DD",X"DE",X"FF",X"00",X"00",X"EA",X"AA",X"AA",X"9A",X"DD",X"DD",X"FF",X"00",X"00",X"E9",X"7A",
		X"AA",X"A9",X"0E",X"DD",X"FF",X"00",X"00",X"EA",X"77",X"7A",X"AA",X"0E",X"DD",X"FF",X"00",X"00",
		X"EE",X"AA",X"A7",X"A0",X"0E",X"CC",X"FF",X"00",X"00",X"0E",X"AA",X"AA",X"90",X"00",X"C0",X"FF",
		X"00",X"00",X"0E",X"77",X"AA",X"A0",X"00",X"00",X"FF",X"00",X"00",X"0E",X"EA",X"7A",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"EA",X"A9",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"E0",X"A0",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"FF",X"00",X"00",X"77",
		X"00",X"00",X"00",X"FF",X"00",X"09",X"41",X"70",X"00",X"00",X"FF",X"00",X"4E",X"EE",X"EE",X"DD",
		X"00",X"FF",X"07",X"5E",X"E7",X"6B",X"DD",X"D0",X"FF",X"07",X"5E",X"79",X"9A",X"AD",X"D0",X"FF",
		X"0A",X"EB",X"99",X"76",X"4E",X"C0",X"FF",X"0A",X"EA",X"97",X"99",X"A0",X"00",X"FF",X"0A",X"EA",
		X"99",X"96",X"40",X"00",X"FF",X"0D",X"EB",X"9A",X"79",X"A0",X"00",X"FF",X"ED",X"DC",X"CA",X"79",
		X"10",X"00",X"FF",X"ED",X"DD",X"CE",X"EE",X"00",X"00",X"FF",X"0E",X"EE",X"E0",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"0E",X"08",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"0E",X"EE",X"88",
		X"EC",X"C0",X"00",X"00",X"FF",X"00",X"00",X"EA",X"AA",X"EE",X"EE",X"CD",X"00",X"00",X"FF",X"00",
		X"0E",X"BE",X"77",X"AA",X"4E",X"DD",X"D0",X"00",X"FF",X"00",X"0E",X"AE",X"E5",X"5A",X"AE",X"7D",
		X"D0",X"00",X"FF",X"0E",X"EE",X"A7",X"EE",X"34",X"AA",X"ED",X"D0",X"00",X"FF",X"EE",X"8E",X"A6",
		X"6E",X"E2",X"EE",X"ED",X"00",X"00",X"FF",X"E8",X"8E",X"B7",X"55",X"EE",X"99",X"A0",X"00",X"00",
		X"FF",X"EE",X"E4",X"B9",X"75",X"E5",X"54",X"60",X"00",X"00",X"FF",X"EE",X"44",X"EB",X"9E",X"79",
		X"99",X"90",X"00",X"00",X"FF",X"0E",X"EE",X"7E",X"EA",X"A9",X"55",X"46",X"00",X"00",X"FF",X"0E",
		X"E7",X"7E",X"DA",X"99",X"99",X"99",X"00",X"00",X"FF",X"00",X"EE",X"ED",X"EA",X"AA",X"A5",X"54",
		X"00",X"00",X"FF",X"00",X"0E",X"ED",X"EE",X"AA",X"99",X"77",X"00",X"00",X"FF",X"00",X"00",X"EC",
		X"CC",X"EE",X"AA",X"A9",X"90",X"00",X"FF",X"00",X"00",X"EE",X"CC",X"EE",X"EE",X"AA",X"10",X"00",
		X"FF",X"00",X"00",X"0E",X"0C",X"0E",X"EE",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"E0",X"00",X"00",X"FF",X"00",X"00",X"00",X"0E",X"04",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"0E",X"EE",X"44",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"EA",X"AA",X"EE",X"E7",X"00",
		X"00",X"00",X"FF",X"00",X"0E",X"BE",X"77",X"AA",X"77",X"EE",X"EC",X"00",X"FF",X"00",X"0E",X"AE",
		X"E5",X"7A",X"AE",X"8D",X"DC",X"C0",X"FF",X"0E",X"EE",X"A7",X"EE",X"47",X"AA",X"ED",X"D0",X"00",
		X"FF",X"EE",X"4E",X"A5",X"5E",X"E3",X"EE",X"ED",X"00",X"00",X"FF",X"E4",X"4E",X"B7",X"44",X"EE",
		X"99",X"A0",X"00",X"00",X"FF",X"EE",X"E7",X"B7",X"73",X"E1",X"45",X"60",X"00",X"00",X"FF",X"EE",
		X"77",X"E9",X"9E",X"57",X"79",X"90",X"00",X"00",X"FF",X"0E",X"EE",X"8E",X"DA",X"79",X"14",X"56",
		X"00",X"00",X"FF",X"0E",X"E8",X"8D",X"DA",X"95",X"77",X"99",X"00",X"00",X"FF",X"00",X"EE",X"DD",
		X"EA",X"A7",X"A1",X"46",X"00",X"00",X"FF",X"00",X"0E",X"DD",X"EE",X"AA",X"57",X"77",X"00",X"00",
		X"FF",X"00",X"0E",X"CC",X"EE",X"EE",X"AA",X"14",X"60",X"00",X"FF",X"00",X"00",X"EC",X"0E",X"EE",
		X"EE",X"AA",X"10",X"00",X"FF",X"00",X"00",X"00",X"00",X"0E",X"EE",X"E0",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"E0",X"00",X"00",X"FF",X"00",X"00",X"00",X"0E",X"07",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"0E",X"EE",X"77",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"EA",
		X"AA",X"EE",X"E8",X"00",X"00",X"00",X"FF",X"00",X"0E",X"BE",X"77",X"AA",X"88",X"00",X"00",X"00",
		X"FF",X"00",X"0E",X"AE",X"E5",X"5A",X"AE",X"40",X"00",X"00",X"FF",X"0E",X"EE",X"A7",X"EE",X"44",
		X"AA",X"ED",X"D0",X"00",X"FF",X"EE",X"7E",X"A6",X"6E",X"E3",X"EE",X"DD",X"DD",X"00",X"FF",X"E7",
		X"7E",X"B7",X"55",X"EE",X"99",X"A0",X"DD",X"00",X"FF",X"EE",X"E8",X"B7",X"74",X"E6",X"7A",X"A0",
		X"DD",X"00",X"FF",X"EE",X"88",X"E9",X"9E",X"99",X"99",X"90",X"CC",X"00",X"FF",X"0E",X"EE",X"4E",
		X"D5",X"45",X"67",X"AA",X"C0",X"00",X"FF",X"0E",X"E4",X"4D",X"DA",X"99",X"99",X"99",X"00",X"00",
		X"FF",X"0E",X"EE",X"DD",X"EA",X"64",X"56",X"7A",X"00",X"00",X"FF",X"0E",X"CC",X"DD",X"EE",X"AA",
		X"99",X"AA",X"00",X"00",X"FF",X"0E",X"CC",X"CE",X"EE",X"EE",X"64",X"56",X"70",X"00",X"FF",X"00",
		X"00",X"00",X"0E",X"EE",X"EE",X"AA",X"10",X"00",X"FF",X"00",X"00",X"00",X"00",X"0E",X"EE",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"0E",X"E0",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"E9",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"0E",X"EE",X"99",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"EA",X"AA",X"EE",X"EC",X"00",X"00",X"00",X"FF",X"00",X"0E",X"BE",X"77",X"AA",
		X"CC",X"00",X"00",X"00",X"FF",X"00",X"0E",X"AE",X"E5",X"7A",X"AE",X"40",X"00",X"00",X"FF",X"00",
		X"EE",X"A7",X"EE",X"47",X"AA",X"4D",X"D0",X"00",X"FF",X"0E",X"9E",X"A5",X"5E",X"E3",X"EE",X"DD",
		X"DD",X"00",X"FF",X"E9",X"9E",X"B7",X"55",X"EE",X"BA",X"9E",X"DD",X"DC",X"FF",X"EE",X"EC",X"B7",
		X"75",X"E7",X"77",X"70",X"ED",X"CC",X"FF",X"EE",X"CC",X"E9",X"9E",X"9A",X"BA",X"A0",X"00",X"00",
		X"FF",X"0E",X"ED",X"4E",X"E7",X"77",X"77",X"77",X"00",X"00",X"FF",X"0E",X"ED",X"DD",X"D7",X"99",
		X"AB",X"A9",X"00",X"00",X"FF",X"00",X"EE",X"DD",X"E7",X"77",X"77",X"77",X"00",X"00",X"FF",X"00",
		X"EE",X"EE",X"EE",X"79",X"9A",X"BA",X"00",X"00",X"FF",X"00",X"00",X"EE",X"EE",X"EE",X"77",X"77",
		X"70",X"00",X"FF",X"00",X"00",X"00",X"0E",X"EE",X"EE",X"9A",X"10",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"0E",X"EE",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"0E",X"E0",X"00",X"00",
		X"FF",X"00",X"0E",X"EE",X"66",X"EE",X"66",X"EE",X"66",X"EE",X"EE",X"EC",X"FF",X"00",X"CC",X"CC",
		X"CC",X"BC",X"CC",X"CC",X"BB",X"CC",X"DD",X"CB",X"FF",X"0C",X"CC",X"CC",X"BA",X"A9",X"95",X"74",
		X"CC",X"CD",X"DC",X"BE",X"FF",X"EC",X"CD",X"7D",X"CC",X"CA",X"57",X"4D",X"DD",X"DD",X"BB",X"DE",
		X"FF",X"EC",X"CD",X"7D",X"B7",X"7C",X"CC",X"DD",X"66",X"6B",X"BD",X"DE",X"FF",X"EC",X"CB",X"CB",
		X"B7",X"74",X"45",X"7D",X"D6",X"BA",X"DD",X"CE",X"FF",X"EC",X"CD",X"7E",X"B7",X"DD",X"B7",X"77",
		X"DB",X"AD",X"6D",X"CE",X"FF",X"EC",X"CD",X"7E",X"BD",X"CC",X"B7",X"32",X"11",X"D6",X"6D",X"BE",
		X"FF",X"EC",X"CC",X"CC",X"CC",X"CC",X"B5",X"73",X"21",X"DD",X"6D",X"CE",X"FF",X"EB",X"BB",X"BB",
		X"BB",X"BB",X"C5",X"57",X"32",X"DD",X"D7",X"C6",X"FF",X"EC",X"BB",X"BC",X"BB",X"BC",X"CB",X"55",
		X"73",X"5D",X"77",X"C6",X"FF",X"EC",X"CC",X"CD",X"B3",X"1C",X"CB",X"B5",X"57",X"BC",X"75",X"BE",
		X"FF",X"ED",X"CC",X"DC",X"31",X"7C",X"CB",X"BB",X"55",X"4C",X"55",X"CE",X"FF",X"0E",X"ED",X"C3",
		X"17",X"5C",X"BC",X"BB",X"BA",X"4C",X"59",X"C6",X"FF",X"00",X"EB",X"31",X"75",X"CC",X"BB",X"BB",
		X"BA",X"7C",X"A9",X"C6",X"FF",X"00",X"B3",X"17",X"5C",X"DB",X"BB",X"BB",X"A7",X"77",X"CA",X"BE",
		X"FF",X"00",X"01",X"75",X"CD",X"CD",X"B3",X"2B",X"AB",X"BB",X"C9",X"CE",X"FF",X"00",X"00",X"5C",
		X"ED",X"DB",X"31",X"7B",X"AE",X"EE",X"C9",X"C6",X"FF",X"00",X"00",X"00",X"0D",X"B3",X"17",X"5B",
		X"77",X"77",X"C9",X"C6",X"FF",X"00",X"00",X"00",X"DB",X"31",X"75",X"BB",X"77",X"77",X"CA",X"BE",
		X"FF",X"00",X"00",X"00",X"B3",X"17",X"5C",X"BB",X"BB",X"BB",X"BA",X"BE",X"FF",X"00",X"00",X"00",
		X"31",X"75",X"CC",X"BB",X"DD",X"BD",X"DC",X"BE",X"FF",X"00",X"00",X"00",X"07",X"5C",X"EC",X"BB",
		X"77",X"C7",X"7C",X"CE",X"FF",X"00",X"00",X"00",X"00",X"00",X"0E",X"CB",X"DD",X"BD",X"DC",X"B0",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"EB",X"CC",X"CC",X"CC",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0E",X"EE",X"EE",X"E0",X"00",X"FF",X"00",X"00",X"00",X"EE",X"CC",X"CC",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"0E",X"EC",X"CC",X"BB",X"CE",X"E0",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"EE",X"77",X"DC",X"CB",X"CE",X"E6",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"0E",X"EC",X"77",X"D7",X"CB",X"BC",X"EE",X"00",X"00",X"00",X"00",X"FF",X"00",X"EE",X"77",
		X"DD",X"77",X"7C",X"AA",X"CE",X"E0",X"00",X"00",X"00",X"FF",X"00",X"EC",X"77",X"DC",X"7D",X"7C",
		X"99",X"CE",X"E6",X"00",X"00",X"00",X"FF",X"00",X"EC",X"BB",X"BC",X"CD",X"44",X"C5",X"5C",X"EE",
		X"00",X"00",X"00",X"FF",X"0D",X"DD",X"DD",X"BB",X"CC",X"D4",X"4C",X"77",X"CE",X"E0",X"00",X"00",
		X"FF",X"A3",X"33",X"33",X"3B",X"BC",X"CD",X"44",X"C4",X"CD",X"E6",X"00",X"00",X"FF",X"71",X"11",
		X"11",X"11",X"CB",X"CC",X"73",X"3D",X"DC",X"DE",X"00",X"00",X"FF",X"55",X"55",X"55",X"55",X"CB",
		X"B7",X"33",X"2D",X"6D",X"CD",X"E0",X"00",X"FF",X"CB",X"BB",X"BB",X"BC",X"BB",X"57",X"32",X"2D",
		X"66",X"DC",X"DE",X"00",X"FF",X"0D",X"DD",X"DD",X"CB",X"BB",X"57",X"32",X"1D",X"DD",X"DD",X"DD",
		X"E0",X"FF",X"00",X"ED",X"CC",X"BB",X"BB",X"57",X"32",X"11",X"BB",X"BB",X"CC",X"CC",X"FF",X"00",
		X"ED",X"CC",X"BB",X"BB",X"57",X"32",X"11",X"BB",X"BB",X"CC",X"CC",X"FF",X"0D",X"DD",X"DD",X"CB",
		X"BB",X"57",X"32",X"1D",X"DD",X"DD",X"DD",X"E0",X"FF",X"A3",X"33",X"33",X"3B",X"BB",X"57",X"32",
		X"2D",X"66",X"DC",X"DE",X"00",X"FF",X"71",X"11",X"11",X"11",X"CA",X"A7",X"33",X"2D",X"6D",X"CD",
		X"E0",X"00",X"FF",X"55",X"55",X"55",X"55",X"CA",X"AA",X"73",X"3D",X"DC",X"DE",X"00",X"00",X"FF",
		X"CB",X"BB",X"BB",X"BC",X"CA",X"AA",X"BB",X"C4",X"CD",X"E6",X"00",X"00",X"FF",X"0D",X"DD",X"DD",
		X"CC",X"AA",X"AA",X"4C",X"77",X"CE",X"E0",X"00",X"00",X"FF",X"00",X"DC",X"CB",X"BA",X"AE",X"74",
		X"C5",X"5C",X"EE",X"00",X"00",X"00",X"FF",X"00",X"EC",X"BD",X"E7",X"7D",X"E7",X"99",X"CE",X"E6",
		X"00",X"00",X"00",X"FF",X"00",X"EE",X"B7",X"DE",X"77",X"DE",X"AA",X"CE",X"E0",X"00",X"00",X"00",
		X"FF",X"00",X"0E",X"E7",X"7D",X"E7",X"7C",X"BB",X"EE",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"EE",X"C7",X"DE",X"7B",X"BE",X"E6",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"0E",X"E7",X"7D",
		X"CB",X"BE",X"E0",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"EE",X"CC",X"CC",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"EE",X"9C",X"7C",X"90",X"FF",X"00",X"00",X"00",
		X"00",X"EE",X"E7",X"DD",X"00",X"FF",X"EE",X"EE",X"E0",X"EE",X"EE",X"E0",X"FF",X"EE",X"AD",X"DA",
		X"EA",X"DD",X"A0",X"FF",X"EE",X"A7",X"DA",X"EA",X"D7",X"A0",X"FF",X"EE",X"97",X"79",X"E9",X"77",
		X"90",X"FF",X"EE",X"87",X"E8",X"E8",X"7E",X"80",X"FF",X"EE",X"66",X"66",X"E6",X"66",X"60",X"FF",
		X"EE",X"BB",X"BB",X"EB",X"BB",X"B0",X"FF",X"0E",X"EE",X"BC",X"AC",X"BE",X"00",X"FF",X"0E",X"CC",
		X"BC",X"9C",X"BC",X"C0",X"FF",X"0E",X"BC",X"BC",X"8C",X"BB",X"C0",X"FF",X"0E",X"EE",X"AC",X"4C",
		X"AE",X"00",X"FF",X"0E",X"CB",X"AE",X"2E",X"AB",X"C0",X"FF",X"0E",X"BB",X"EE",X"1E",X"EB",X"C0",
		X"FF",X"0E",X"EE",X"66",X"26",X"6E",X"00",X"FF",X"0E",X"CC",X"B9",X"49",X"BC",X"C0",X"FF",X"00",
		X"BC",X"DC",X"6C",X"DB",X"B0",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"EE",X"EE",
		X"E0",X"EE",X"EE",X"E0",X"00",X"FF",X"EE",X"EE",X"E0",X"EE",X"EE",X"E0",X"00",X"FF",X"EE",X"EE",
		X"E0",X"EE",X"EE",X"E0",X"00",X"FF",X"EE",X"8D",X"DD",X"8E",X"87",X"DD",X"80",X"FF",X"EE",X"65",
		X"7D",X"6E",X"67",X"7D",X"60",X"FF",X"EE",X"47",X"5E",X"4E",X"45",X"57",X"40",X"FF",X"EE",X"35",
		X"7E",X"3E",X"35",X"57",X"30",X"FF",X"EE",X"2E",X"EE",X"2C",X"2E",X"EE",X"20",X"FF",X"EE",X"11",
		X"11",X"16",X"11",X"11",X"10",X"FF",X"00",X"EE",X"CA",X"C4",X"CA",X"4B",X"00",X"FF",X"00",X"EB",
		X"CA",X"E2",X"EA",X"4C",X"00",X"FF",X"00",X"EC",X"BE",X"E1",X"EE",X"B0",X"00",X"FF",X"00",X"EE",
		X"B6",X"62",X"66",X"9B",X"00",X"FF",X"00",X"EB",X"BB",X"94",X"99",X"CC",X"00",X"FF",X"00",X"0C",
		X"CE",X"B6",X"B0",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"E0",X"00",X"00",X"E0",
		X"00",X"00",X"00",X"FF",X"00",X"0E",X"EE",X"00",X"0E",X"EE",X"00",X"00",X"00",X"FF",X"00",X"0E",
		X"EE",X"30",X"EE",X"3E",X"E0",X"00",X"00",X"FF",X"00",X"04",X"EE",X"E6",X"E6",X"EE",X"E4",X"00",
		X"00",X"FF",X"00",X"DD",X"3E",X"E6",X"E6",X"EE",X"37",X"70",X"00",X"FF",X"05",X"7D",X"E2",X"BB",
		X"6B",X"B2",X"E7",X"75",X"00",X"FF",X"47",X"7D",X"EE",X"1B",X"4B",X"1E",X"ED",X"D7",X"40",X"FF",
		X"03",X"ED",X"E1",X"BB",X"2B",X"B1",X"ED",X"E3",X"00",X"FF",X"00",X"2E",X"1A",X"AE",X"4E",X"BA",
		X"1E",X"20",X"00",X"FF",X"00",X"01",X"CC",X"AE",X"4E",X"AA",X"B1",X"00",X"00",X"FF",X"00",X"0E",
		X"EB",X"EA",X"4A",X"EB",X"B0",X"00",X"00",X"FF",X"00",X"0E",X"CB",X"A8",X"48",X"AE",X"00",X"00",
		X"00",X"FF",X"00",X"0E",X"BB",X"BA",X"4A",X"BC",X"C0",X"00",X"00",X"FF",X"00",X"00",X"00",X"0B",
		X"4B",X"EB",X"B0",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"EE",X"0E",X"E0",X"00",X"FF",X"EE",X"EE",X"66",X"E6",X"6E",X"E0",X"FF",
		X"EE",X"EE",X"E6",X"E6",X"EE",X"E0",X"FF",X"EE",X"EE",X"EB",X"CB",X"EE",X"E0",X"FF",X"E6",X"32",
		X"1B",X"BB",X"12",X"36",X"FF",X"E7",X"7E",X"1B",X"4B",X"1E",X"57",X"FF",X"E7",X"DE",X"19",X"49",
		X"1E",X"77",X"FF",X"E5",X"7E",X"18",X"48",X"1E",X"75",X"FF",X"E7",X"DE",X"18",X"48",X"1E",X"DD",
		X"FF",X"06",X"32",X"19",X"49",X"12",X"36",X"FF",X"0E",X"BB",X"BB",X"4B",X"CC",X"C0",X"FF",X"0E",
		X"CC",X"EB",X"4B",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"03",X"00",X"03",X"00",X"00",X"FF",X"00",X"00",
		X"E0",X"60",X"60",X"00",X"00",X"FF",X"00",X"00",X"0E",X"6E",X"60",X"00",X"00",X"FF",X"00",X"00",
		X"0E",X"CB",X"C0",X"00",X"00",X"FF",X"EE",X"EE",X"0E",X"B6",X"BE",X"EE",X"E0",X"FF",X"E6",X"6C",
		X"CE",X"B6",X"BE",X"BC",X"66",X"FF",X"E7",X"6B",X"CE",X"94",X"9E",X"BC",X"65",X"FF",X"E7",X"6B",
		X"CE",X"92",X"9E",X"BC",X"65",X"FF",X"E7",X"6B",X"CE",X"91",X"9E",X"BC",X"65",X"FF",X"E7",X"6B",
		X"CA",X"94",X"9B",X"CB",X"65",X"FF",X"08",X"6B",X"CC",X"B9",X"BC",X"BC",X"68",X"FF",X"00",X"00",
		X"00",X"C9",X"C0",X"BB",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9B",X"BB",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"8C",X"CC",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"66",X"66",X"6B",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"BB",X"BB",X"BB",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"CC",X"CC",X"CB",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"00",X"EE",X"EE",X"EB",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0E",X"66",X"B9",X"64",X"46",X"9B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"EE",X"44",X"44",X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"B9",X"64",X"46",X"9B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",
		X"EE",X"EE",X"EE",X"EB",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",
		X"0E",X"CC",X"CC",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",
		X"BB",X"BB",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"66",
		X"66",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"8C",X"CC",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"9C",X"CC",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"EE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"11",X"00",X"00",X"00",X"01",X"10",X"FF",
		X"00",X"11",X"01",X"01",X"10",X"00",X"FF",X"00",X"00",X"13",X"10",X"00",X"00",X"FF",X"00",X"00",
		X"03",X"00",X"00",X"00",X"FF",X"22",X"00",X"00",X"00",X"02",X"20",X"FF",X"00",X"22",X"02",X"02",
		X"20",X"00",X"FF",X"00",X"00",X"21",X"20",X"00",X"00",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"33",X"00",X"00",X"00",X"03",X"30",X"FF",X"00",X"33",X"03",X"03",X"30",X"00",X"FF",X"00",
		X"00",X"32",X"30",X"00",X"00",X"FF",X"00",X"00",X"02",X"00",X"00",X"00",X"FF",X"10",X"00",X"00",
		X"00",X"10",X"FF",X"10",X"00",X"00",X"00",X"10",X"FF",X"01",X"00",X"10",X"01",X"00",X"FF",X"00",
		X"11",X"11",X"10",X"00",X"FF",X"00",X"01",X"31",X"00",X"00",X"FF",X"00",X"00",X"30",X"00",X"00",
		X"FF",X"20",X"00",X"00",X"00",X"20",X"FF",X"20",X"00",X"00",X"00",X"20",X"FF",X"02",X"00",X"20",
		X"02",X"00",X"FF",X"00",X"22",X"22",X"20",X"00",X"FF",X"00",X"02",X"12",X"00",X"00",X"FF",X"00",
		X"00",X"10",X"00",X"00",X"FF",X"30",X"00",X"00",X"00",X"30",X"FF",X"30",X"00",X"00",X"00",X"30",
		X"FF",X"03",X"00",X"30",X"03",X"00",X"FF",X"00",X"33",X"33",X"30",X"00",X"FF",X"00",X"03",X"23",
		X"00",X"00",X"FF",X"00",X"00",X"20",X"00",X"00",X"FF",X"DD",X"DD",X"00",X"FF",X"D9",X"DD",X"CE",
		X"00",X"FF",X"09",X"DE",X"CE",X"00",X"FF",X"CC",X"C9",X"80",X"FF",X"98",X"86",X"7D",X"D6",X"55",
		X"78",X"FF",X"99",X"88",X"ED",X"65",X"5A",X"68",X"FF",X"09",X"98",X"E6",X"55",X"57",X"88",X"FF",
		X"00",X"99",X"86",X"66",X"27",X"89",X"FF",X"00",X"09",X"98",X"17",X"68",X"90",X"FF",X"00",X"00",
		X"98",X"88",X"89",X"00",X"FF",X"00",X"00",X"09",X"88",X"90",X"00",X"FF",X"00",X"00",X"00",X"99",
		X"00",X"00",X"FF",X"00",X"00",X"A0",X"00",X"00",X"FF",X"00",X"0E",X"90",X"00",X"00",X"FF",X"00",
		X"0E",X"60",X"00",X"00",X"FF",X"00",X"06",X"16",X"00",X"00",X"FF",X"BB",X"52",X"12",X"9A",X"B0",
		X"FF",X"EE",X"E6",X"26",X"0E",X"00",X"FF",X"0E",X"EE",X"6E",X"E0",X"00",X"FF",X"00",X"EE",X"BE",
		X"00",X"00",X"FF",X"00",X"0E",X"C0",X"00",X"00",X"FF",X"00",X"09",X"60",X"00",X"FF",X"00",X"E9",
		X"50",X"00",X"FF",X"00",X"E5",X"40",X"00",X"FF",X"09",X"21",X"34",X"60",X"FF",X"EA",X"22",X"35",
		X"70",X"FF",X"EE",X"E8",X"6E",X"00",X"FF",X"00",X"E9",X"80",X"00",X"FF",X"00",X"EA",X"90",X"00",
		X"FF",X"00",X"09",X"60",X"00",X"FF",X"00",X"E9",X"50",X"00",X"FF",X"00",X"E5",X"40",X"00",X"FF",
		X"09",X"75",X"21",X"60",X"FF",X"EA",X"85",X"22",X"70",X"FF",X"0E",X"E8",X"6E",X"00",X"FF",X"00",
		X"E9",X"8E",X"00",X"FF",X"00",X"EA",X"90",X"00",X"FF",X"00",X"09",X"60",X"00",X"FF",X"00",X"E9",
		X"50",X"00",X"FF",X"00",X"E6",X"60",X"00",X"FF",X"09",X"75",X"54",X"60",X"FF",X"EA",X"92",X"15",
		X"70",X"FF",X"0E",X"E2",X"2E",X"00",X"FF",X"0E",X"E9",X"80",X"00",X"FF",X"0E",X"EA",X"90",X"00",
		X"FF",X"00",X"EE",X"00",X"00",X"FF",X"00",X"09",X"60",X"00",X"FF",X"0E",X"E9",X"50",X"00",X"FF",
		X"0E",X"E2",X"10",X"00",X"FF",X"09",X"72",X"24",X"60",X"FF",X"EA",X"95",X"55",X"70",X"FF",X"0E",
		X"E8",X"6E",X"00",X"FF",X"00",X"E9",X"80",X"00",X"FF",X"00",X"EA",X"90",X"00",X"FF",X"00",X"0B",
		X"A0",X"00",X"FF",X"00",X"74",X"36",X"00",X"FF",X"0A",X"42",X"13",X"90",X"FF",X"0B",X"42",X"24",
		X"A0",X"FF",X"EE",X"84",X"46",X"00",X"FF",X"EE",X"EB",X"A0",X"00",X"FF",X"0E",X"E0",X"00",X"00",
		X"FF",X"00",X"00",X"09",X"40",X"00",X"FF",X"00",X"00",X"96",X"38",X"00",X"FF",X"00",X"09",X"64",
		X"24",X"80",X"FF",X"00",X"A4",X"32",X"13",X"49",X"FF",X"00",X"A6",X"55",X"24",X"69",X"FF",X"0C",
		X"C9",X"65",X"36",X"80",X"FF",X"BC",X"DD",X"96",X"48",X"00",X"FF",X"BC",X"DD",X"CA",X"80",X"00",
		X"FF",X"0C",X"CC",X"C0",X"00",X"00",X"FF",X"00",X"BB",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"09",X"50",X"00",X"FF",X"00",X"00",X"00",X"88",X"47",X"00",X"FF",X"00",X"00",X"09",X"88",X"37",
		X"90",X"FF",X"00",X"00",X"08",X"78",X"27",X"70",X"FF",X"00",X"00",X"54",X"32",X"12",X"34",X"FF",
		X"00",X"00",X"98",X"83",X"27",X"78",X"FF",X"00",X"00",X"08",X"78",X"37",X"70",X"FF",X"00",X"00",
		X"09",X"88",X"47",X"90",X"FF",X"00",X"00",X"00",X"88",X"57",X"00",X"FF",X"00",X"CC",X"00",X"A9",
		X"60",X"00",X"FF",X"0C",X"CC",X"C0",X"00",X"00",X"00",X"FF",X"BC",X"EE",X"CB",X"00",X"00",X"00",
		X"FF",X"BC",X"EE",X"CB",X"00",X"00",X"00",X"FF",X"0C",X"CC",X"C0",X"00",X"00",X"00",X"FF",X"00",
		X"CC",X"00",X"00",X"00",X"00",X"FF",X"08",X"77",X"E5",X"57",X"8B",X"00",X"FF",X"9B",X"71",X"3E",
		X"44",X"89",X"00",X"FF",X"99",X"89",X"73",X"34",X"50",X"00",X"FF",X"99",X"BB",X"BB",X"B4",X"48",
		X"44",X"FF",X"09",X"9B",X"BC",X"CB",X"B8",X"80",X"FF",X"00",X"BC",X"CD",X"DD",X"C9",X"78",X"FF",
		X"09",X"BC",X"CD",X"DD",X"C9",X"78",X"FF",X"09",X"9B",X"BC",X"CB",X"B8",X"80",X"FF",X"00",X"BB",
		X"BB",X"B4",X"48",X"44",X"FF",X"09",X"89",X"73",X"34",X"50",X"00",X"FF",X"9B",X"81",X"34",X"45",
		X"89",X"00",X"FF",X"98",X"77",X"E5",X"67",X"8B",X"00",X"FF",X"99",X"99",X"99",X"99",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"B6",X"00",X"FF",X"00",X"00",X"99",X"00",X"86",X"40",X"FF",X"00",
		X"00",X"99",X"90",X"75",X"E0",X"FF",X"0B",X"87",X"66",X"66",X"74",X"E0",X"FF",X"9B",X"8A",X"61",
		X"62",X"86",X"40",X"FF",X"99",X"89",X"79",X"79",X"86",X"00",X"FF",X"99",X"BB",X"BB",X"BB",X"B8",
		X"54",X"FF",X"00",X"9B",X"BD",X"EB",X"BB",X"80",X"FF",X"09",X"BC",X"DE",X"EE",X"D9",X"78",X"FF",
		X"09",X"BC",X"DE",X"3E",X"D9",X"78",X"FF",X"09",X"9B",X"BD",X"DB",X"BB",X"80",X"FF",X"00",X"BB",
		X"BB",X"BB",X"B8",X"54",X"FF",X"09",X"89",X"79",X"79",X"86",X"00",X"FF",X"9B",X"8A",X"61",X"62",
		X"86",X"40",X"FF",X"9B",X"88",X"66",X"66",X"74",X"E0",X"FF",X"99",X"99",X"99",X"99",X"75",X"E0",
		X"FF",X"00",X"00",X"99",X"90",X"85",X"40",X"FF",X"00",X"00",X"99",X"00",X"B6",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"E0",X"00",X"FF",X"00",X"00",X"90",X"00",X"86",X"00",X"FF",X"00",X"00",X"99",
		X"00",X"86",X"60",X"FF",X"00",X"00",X"99",X"90",X"75",X"40",X"FF",X"00",X"00",X"99",X"90",X"65",
		X"30",X"FF",X"00",X"00",X"99",X"90",X"65",X"40",X"FF",X"0B",X"87",X"66",X"68",X"76",X"50",X"FF",
		X"9B",X"82",X"6A",X"61",X"86",X"60",X"FF",X"99",X"89",X"79",X"79",X"86",X"00",X"FF",X"99",X"BB",
		X"BB",X"BB",X"B8",X"55",X"FF",X"00",X"9B",X"BC",X"CB",X"BB",X"80",X"FF",X"09",X"BC",X"DE",X"ED",
		X"C9",X"78",X"FF",X"09",X"BC",X"DE",X"ED",X"C9",X"78",X"FF",X"09",X"9B",X"BC",X"CB",X"BB",X"80",
		X"FF",X"00",X"BB",X"BB",X"BB",X"B8",X"55",X"FF",X"09",X"89",X"79",X"79",X"86",X"00",X"FF",X"9B",
		X"82",X"6A",X"61",X"86",X"60",X"FF",X"9B",X"88",X"66",X"67",X"86",X"50",X"FF",X"99",X"99",X"99",
		X"99",X"75",X"40",X"FF",X"00",X"00",X"99",X"90",X"65",X"30",X"FF",X"00",X"00",X"99",X"90",X"65",
		X"40",X"FF",X"00",X"00",X"99",X"90",X"76",X"50",X"FF",X"00",X"00",X"99",X"90",X"86",X"60",X"FF",
		X"00",X"00",X"99",X"00",X"86",X"00",X"FF",X"00",X"00",X"90",X"00",X"E0",X"00",X"FF",X"00",X"05",
		X"08",X"80",X"50",X"00",X"FF",X"00",X"05",X"87",X"78",X"50",X"00",X"FF",X"08",X"88",X"89",X"98",
		X"88",X"80",X"FF",X"97",X"45",X"39",X"93",X"54",X"70",X"FF",X"94",X"43",X"BC",X"CB",X"34",X"40",
		X"FF",X"55",X"3B",X"CC",X"CC",X"B3",X"55",X"FF",X"53",X"2B",X"CD",X"DC",X"B2",X"35",X"FF",X"37",
		X"7B",X"CD",X"DC",X"B7",X"73",X"FF",X"96",X"1B",X"CD",X"DC",X"B1",X"60",X"FF",X"97",X"7B",X"CC",
		X"CC",X"B7",X"70",X"FF",X"98",X"AB",X"9C",X"C9",X"BA",X"80",X"FF",X"98",X"8B",X"9B",X"B9",X"B8",
		X"80",X"FF",X"98",X"80",X"99",X"99",X"98",X"80",X"FF",X"99",X"00",X"00",X"00",X"99",X"00",X"FF",
		X"00",X"00",X"05",X"08",X"80",X"50",X"00",X"00",X"FF",X"00",X"00",X"05",X"87",X"78",X"50",X"00",
		X"00",X"FF",X"00",X"64",X"68",X"89",X"98",X"86",X"45",X"00",X"FF",X"66",X"43",X"46",X"6C",X"C6",
		X"64",X"34",X"46",X"FF",X"B8",X"77",X"78",X"BD",X"DB",X"87",X"77",X"8B",X"FF",X"00",X"96",X"6B",
		X"DE",X"3D",X"B6",X"60",X"00",X"FF",X"00",X"96",X"1B",X"DE",X"ED",X"B1",X"69",X"00",X"FF",X"99",
		X"96",X"6B",X"CE",X"EC",X"B6",X"69",X"99",X"FF",X"99",X"97",X"AB",X"CD",X"DC",X"BA",X"79",X"99",
		X"FF",X"00",X"97",X"6B",X"CC",X"CC",X"B6",X"70",X"00",X"FF",X"00",X"97",X"2B",X"9C",X"C9",X"B2",
		X"70",X"00",X"FF",X"00",X"98",X"8B",X"9B",X"B9",X"B8",X"80",X"00",X"FF",X"00",X"98",X"80",X"99",
		X"99",X"98",X"80",X"00",X"FF",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"05",X"08",X"80",X"50",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"05",
		X"87",X"78",X"50",X"00",X"00",X"00",X"00",X"FF",X"00",X"66",X"54",X"35",X"68",X"89",X"98",X"86",
		X"55",X"34",X"56",X"00",X"FF",X"66",X"65",X"44",X"44",X"56",X"6C",X"C6",X"65",X"54",X"44",X"55",
		X"66",X"FF",X"E8",X"88",X"76",X"67",X"88",X"BD",X"DB",X"88",X"87",X"66",X"78",X"8E",X"FF",X"00",
		X"00",X"00",X"96",X"6B",X"CE",X"EC",X"B6",X"60",X"00",X"00",X"00",X"FF",X"00",X"99",X"99",X"96",
		X"AB",X"CE",X"EC",X"BA",X"69",X"99",X"99",X"00",X"FF",X"99",X"99",X"99",X"96",X"6B",X"CD",X"DC",
		X"B6",X"69",X"99",X"99",X"99",X"FF",X"99",X"99",X"99",X"97",X"2B",X"CD",X"DC",X"B2",X"79",X"99",
		X"99",X"99",X"FF",X"00",X"00",X"00",X"97",X"6B",X"CC",X"CC",X"B6",X"70",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"98",X"1B",X"9C",X"C9",X"B1",X"80",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"98",X"80",X"9B",X"B9",X"98",X"80",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"98",X"80",X"99",
		X"99",X"98",X"80",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"07",X"88",X"00",X"50",X"00",X"FF",X"00",X"00",X"74",X"A7",
		X"85",X"78",X"00",X"FF",X"00",X"04",X"44",X"45",X"99",X"77",X"50",X"FF",X"00",X"65",X"66",X"66",
		X"C9",X"95",X"00",X"FF",X"00",X"72",X"7B",X"DD",X"EC",X"98",X"00",X"FF",X"07",X"87",X"6B",X"DE",
		X"D4",X"38",X"80",X"FF",X"81",X"78",X"BC",X"ED",X"B4",X"37",X"80",X"FF",X"88",X"8B",X"CC",X"CB",
		X"B4",X"47",X"80",X"FF",X"98",X"9B",X"CC",X"B6",X"64",X"68",X"90",X"FF",X"09",X"99",X"BB",X"82",
		X"66",X"69",X"00",X"FF",X"00",X"00",X"98",X"88",X"76",X"90",X"00",X"FF",X"00",X"00",X"81",X"88",
		X"89",X"00",X"00",X"FF",X"00",X"00",X"88",X"88",X"90",X"00",X"00",X"FF",X"00",X"00",X"98",X"89",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"09",X"90",X"00",X"00",X"00",X"FF",X"00",X"00",X"66",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"0B",X"55",X"60",X"00",X"00",X"00",X"00",X"FF",X"09",X"90",
		X"75",X"36",X"00",X"40",X"00",X"00",X"FF",X"99",X"99",X"67",X"44",X"74",X"78",X"00",X"00",X"FF",
		X"09",X"96",X"28",X"85",X"99",X"77",X"40",X"00",X"FF",X"00",X"76",X"6B",X"8B",X"D9",X"94",X"00",
		X"00",X"FF",X"0B",X"81",X"6B",X"EE",X"3D",X"97",X"00",X"00",X"FF",X"08",X"88",X"BD",X"E3",X"E8",
		X"65",X"60",X"00",X"FF",X"8A",X"88",X"BD",X"3E",X"EB",X"85",X"55",X"00",X"FF",X"88",X"8B",X"CD",
		X"DB",X"BB",X"77",X"53",X"50",X"FF",X"98",X"9B",X"CC",X"BB",X"66",X"67",X"75",X"50",X"FF",X"09",
		X"99",X"BB",X"88",X"16",X"69",X"0B",X"60",X"FF",X"00",X"00",X"99",X"87",X"76",X"99",X"90",X"00",
		X"FF",X"00",X"00",X"08",X"A8",X"79",X"99",X"99",X"00",X"FF",X"00",X"00",X"88",X"88",X"90",X"09",
		X"99",X"00",X"FF",X"00",X"00",X"98",X"89",X"00",X"00",X"99",X"00",X"FF",X"00",X"00",X"09",X"90",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"E6",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"08",X"55",X"60",X"00",X"00",X"00",X"00",X"00",X"FF",X"99",X"90",X"74",X"35",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"09",X"99",X"07",X"44",X"60",X"04",X"00",X"00",X"00",X"FF",X"00",X"99",X"96",
		X"75",X"67",X"47",X"80",X"00",X"00",X"FF",X"00",X"09",X"61",X"68",X"B9",X"97",X"74",X"00",X"00",
		X"FF",X"00",X"07",X"68",X"B8",X"BC",X"99",X"40",X"00",X"00",X"FF",X"00",X"97",X"A6",X"BD",X"EE",
		X"C9",X"70",X"00",X"00",X"FF",X"00",X"88",X"8B",X"CD",X"EE",X"86",X"56",X"00",X"00",X"FF",X"08",
		X"28",X"8B",X"CD",X"DD",X"B8",X"55",X"40",X"00",X"FF",X"08",X"88",X"BC",X"CC",X"BB",X"B7",X"74",
		X"34",X"00",X"FF",X"09",X"89",X"BC",X"CB",X"B6",X"16",X"77",X"44",X"60",X"FF",X"00",X"99",X"9B",
		X"B8",X"A6",X"66",X"90",X"75",X"50",X"FF",X"00",X"00",X"09",X"88",X"77",X"69",X"99",X"07",X"56",
		X"FF",X"00",X"00",X"08",X"28",X"87",X"90",X"99",X"90",X"86",X"FF",X"00",X"00",X"08",X"88",X"89",
		X"00",X"09",X"99",X"0E",X"FF",X"00",X"00",X"09",X"88",X"90",X"00",X"00",X"99",X"90",X"FF",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"90",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"90",X"FF",X"11",X"17",X"80",X"FF",X"07",X"AA",X"AA",X"00",X"00",X"00",X"AA",X"AA",X"80",
		X"FF",X"00",X"00",X"00",X"06",X"00",X"00",X"08",X"00",X"80",X"00",X"FF",X"00",X"AE",X"8C",X"CC",
		X"C0",X"FF",X"09",X"EE",X"CC",X"CC",X"CC",X"FF",X"E9",X"7A",X"E6",X"E6",X"E6",X"FF",X"E9",X"AA",
		X"DD",X"DD",X"DD",X"FF",X"EE",X"9A",X"8D",X"DD",X"D0",X"FF",X"0E",X"E8",X"EA",X"8E",X"00",X"FF",
		X"00",X"00",X"00",X"0C",X"C0",X"00",X"FF",X"00",X"00",X"00",X"CC",X"00",X"00",X"FF",X"00",X"AA",
		X"0C",X"C2",X"A0",X"00",X"FF",X"09",X"EE",X"CC",X"A2",X"A2",X"00",X"FF",X"E9",X"7A",X"AB",X"EB",
		X"A4",X"A0",X"FF",X"E9",X"AA",X"DD",X"A4",X"A4",X"00",X"FF",X"EE",X"9A",X"ED",X"D4",X"A0",X"00",
		X"FF",X"0E",X"E0",X"EE",X"DD",X"00",X"00",X"FF",X"00",X"00",X"0E",X"ED",X"D0",X"00",X"FF",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"FF",X"00",X"00",X"0C",X"C0",X"00",X"FF",X"00",X"00",X"0C",X"C0",
		X"00",X"FF",X"00",X"00",X"CC",X"33",X"00",X"FF",X"00",X"00",X"CC",X"30",X"00",X"FF",X"0A",X"AC",
		X"C3",X"3E",X"00",X"FF",X"AA",X"AC",X"CA",X"2E",X"20",X"FF",X"A7",X"E5",X"BE",X"BE",X"4E",X"FF",
		X"AE",X"EC",X"CE",X"4E",X"40",X"FF",X"0A",X"AC",X"C3",X"4E",X"00",X"FF",X"00",X"00",X"CC",X"30",
		X"00",X"FF",X"00",X"00",X"CC",X"33",X"00",X"FF",X"00",X"00",X"0C",X"C0",X"00",X"FF",X"00",X"00",
		X"0C",X"C0",X"00",X"FF",X"00",X"00",X"C3",X"00",X"00",X"FF",X"00",X"0C",X"C3",X"00",X"00",X"FF",
		X"00",X"0C",X"C3",X"00",X"00",X"FF",X"00",X"0C",X"C3",X"00",X"00",X"FF",X"0E",X"EC",X"C0",X"2E",
		X"00",X"FF",X"EA",X"AC",X"4A",X"2E",X"20",X"FF",X"E7",X"E5",X"BE",X"BE",X"4E",X"FF",X"EE",X"EC",
		X"4E",X"4E",X"40",X"FF",X"0A",X"AC",X"C0",X"4E",X"00",X"FF",X"00",X"0C",X"C4",X"00",X"00",X"FF",
		X"00",X"0C",X"C4",X"00",X"00",X"FF",X"00",X"0C",X"C4",X"00",X"00",X"FF",X"00",X"00",X"C4",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"22",X"00",X"FF",X"00",X"00",X"00",X"02",X"20",X"00",X"FF",
		X"00",X"00",X"00",X"22",X"E0",X"00",X"FF",X"00",X"0E",X"E2",X"24",X"E3",X"00",X"FF",X"00",X"EE",
		X"72",X"EB",X"E2",X"E0",X"FF",X"00",X"EA",X"72",X"E4",X"E5",X"E0",X"FF",X"00",X"EA",X"A2",X"25",
		X"E6",X"00",X"FF",X"0E",X"EE",X"E0",X"22",X"E0",X"00",X"FF",X"EE",X"EE",X"EE",X"02",X"20",X"00",
		X"FF",X"0E",X"EE",X"E0",X"00",X"22",X"00",X"FF",X"00",X"EE",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"0E",X"E0",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"20",X"00",X"FF",X"00",X"00",X"02",X"33",
		X"00",X"FF",X"00",X"00",X"02",X"30",X"00",X"FF",X"00",X"0E",X"23",X"5E",X"00",X"FF",X"00",X"AE",
		X"2E",X"4E",X"40",X"FF",X"00",X"A7",X"8E",X"CE",X"CE",X"FF",X"0E",X"A9",X"2E",X"4E",X"40",X"FF",
		X"EE",X"EA",X"23",X"5E",X"00",X"FF",X"EE",X"EE",X"E2",X"3E",X"00",X"FF",X"0E",X"EE",X"02",X"33",
		X"00",X"FF",X"00",X"EE",X"00",X"20",X"00",X"FF",X"00",X"0E",X"E0",X"00",X"00",X"FF",X"00",X"00",
		X"03",X"00",X"00",X"FF",X"00",X"00",X"34",X"40",X"00",X"FF",X"00",X"E3",X"45",X"E0",X"00",X"FF",
		X"0E",X"E4",X"E5",X"E6",X"00",X"FF",X"EE",X"76",X"E4",X"E5",X"E0",X"FF",X"EA",X"94",X"E6",X"E6",
		X"00",X"FF",X"EE",X"A3",X"46",X"E0",X"00",X"FF",X"0E",X"EE",X"34",X"40",X"00",X"FF",X"0E",X"EE",
		X"E3",X"00",X"00",X"FF",X"00",X"EE",X"E0",X"00",X"00",X"FF",X"00",X"0E",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"03",X"30",X"FF",X"00",X"00",X"33",X"00",X"FF",X"00",X"E3",X"3E",X"50",X"FF",X"0A",
		X"73",X"4E",X"3E",X"FF",X"EE",X"A3",X"5E",X"5E",X"FF",X"EE",X"E3",X"3E",X"50",X"FF",X"0E",X"EE",
		X"33",X"00",X"FF",X"00",X"0E",X"E3",X"30",X"FF",X"00",X"00",X"EE",X"00",X"FF",X"00",X"00",X"30",
		X"00",X"FF",X"00",X"03",X"90",X"00",X"FF",X"5E",X"39",X"E6",X"00",X"FF",X"E7",X"E5",X"E3",X"E0",
		X"FF",X"5E",X"3D",X"E8",X"00",X"FF",X"00",X"E3",X"D0",X"00",X"FF",X"00",X"0E",X"30",X"00",X"FF",
		X"0E",X"E0",X"00",X"00",X"00",X"FF",X"E7",X"EE",X"CC",X"CC",X"CC",X"FF",X"EE",X"EC",X"CC",X"CC",
		X"C0",X"FF",X"0E",X"C5",X"4E",X"33",X"30",X"FF",X"0C",X"C4",X"EC",X"E0",X"00",X"FF",X"0C",X"CE",
		X"53",X"E5",X"00",X"FF",X"0C",X"C6",X"5E",X"2D",X"00",X"FF",X"0C",X"C3",X"E5",X"45",X"00",X"FF",
		X"0C",X"C3",X"06",X"5E",X"00",X"FF",X"0C",X"C3",X"00",X"00",X"00",X"FF",X"0C",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"0C",X"C0",X"FF",X"00",X"EE",X"00",X"CC",X"C3",X"FF",X"0E",X"7E",
		X"EC",X"CC",X"33",X"FF",X"0E",X"EE",X"CC",X"C3",X"30",X"FF",X"00",X"EC",X"54",X"E5",X"00",X"FF",
		X"00",X"CC",X"4E",X"BE",X"00",X"FF",X"0C",X"CC",X"E5",X"CE",X"50",X"FF",X"CC",X"C3",X"65",X"EC",
		X"50",X"FF",X"CC",X"33",X"AE",X"D2",X"50",X"FF",X"03",X"30",X"00",X"65",X"E0",X"FF",X"00",X"00",
		X"0E",X"E0",X"00",X"00",X"FF",X"00",X"00",X"EE",X"EE",X"00",X"00",X"FF",X"00",X"00",X"EE",X"7E",
		X"00",X"00",X"FF",X"00",X"00",X"C5",X"6C",X"00",X"00",X"FF",X"00",X"0C",X"C5",X"5C",X"C0",X"00",
		X"FF",X"00",X"CC",X"34",X"B3",X"CC",X"00",X"FF",X"0C",X"C3",X"EE",X"EE",X"3C",X"C0",X"FF",X"CC",
		X"33",X"54",X"B4",X"33",X"CC",X"FF",X"00",X"30",X"EE",X"EE",X"03",X"00",X"FF",X"00",X"00",X"04",
		X"B0",X"00",X"00",X"FF",X"00",X"00",X"0E",X"E0",X"00",X"00",X"FF",X"00",X"00",X"0E",X"E0",X"00",
		X"00",X"FF",X"00",X"00",X"EE",X"EE",X"00",X"00",X"FF",X"00",X"00",X"EE",X"7E",X"00",X"00",X"FF",
		X"CC",X"CC",X"C5",X"5C",X"CC",X"CC",X"FF",X"4C",X"CC",X"C6",X"6C",X"CC",X"C4",X"FF",X"43",X"33",
		X"54",X"B4",X"33",X"34",X"FF",X"33",X"30",X"EE",X"EE",X"03",X"33",X"FF",X"00",X"00",X"54",X"B3",
		X"00",X"00",X"FF",X"00",X"00",X"EE",X"EE",X"00",X"00",X"FF",X"00",X"00",X"04",X"30",X"00",X"00",
		X"FF",X"00",X"00",X"0E",X"E0",X"00",X"00",X"FF",X"00",X"00",X"10",X"00",X"FF",X"00",X"03",X"20",
		X"00",X"FF",X"00",X"00",X"00",X"31",X"FF",X"03",X"09",X"80",X"01",X"FF",X"33",X"08",X"88",X"33",
		X"FF",X"30",X"09",X"80",X"21",X"FF",X"03",X"00",X"00",X"00",X"FF",X"35",X"30",X"33",X"30",X"FF",
		X"03",X"30",X"55",X"00",X"FF",X"00",X"00",X"00",X"11",X"00",X"FF",X"00",X"00",X"00",X"02",X"00",
		X"FF",X"03",X"30",X"00",X"00",X"00",X"FF",X"33",X"00",X"98",X"CE",X"22",X"FF",X"00",X"08",X"98",
		X"88",X"03",X"FF",X"00",X"0B",X"88",X"A8",X"80",X"FF",X"33",X"0D",X"9D",X"DD",X"01",X"FF",X"35",
		X"50",X"9D",X"CE",X"32",X"FF",X"05",X"00",X"30",X"00",X"20",X"FF",X"00",X"05",X"50",X"00",X"00",
		X"FF",X"00",X"00",X"30",X"00",X"00",X"FF",X"00",X"20",X"00",X"02",X"00",X"FF",X"00",X"08",X"00",
		X"00",X"00",X"FF",X"00",X"98",X"10",X"00",X"00",X"FF",X"21",X"98",X"88",X"10",X"00",X"FF",X"0B",
		X"88",X"AA",X"88",X"20",X"FF",X"5D",X"9D",X"DD",X"D0",X"00",X"FF",X"00",X"9D",X"D0",X"00",X"00",
		X"FF",X"00",X"0D",X"00",X"00",X"00",X"FF",X"05",X"00",X"00",X"00",X"00",X"FF",X"00",X"05",X"00",
		X"50",X"00",X"FF",X"09",X"8E",X"CE",X"00",X"FF",X"89",X"88",X"CE",X"00",X"FF",X"89",X"88",X"88",
		X"00",X"FF",X"B8",X"AA",X"88",X"88",X"FF",X"D9",X"DD",X"DD",X"00",X"FF",X"D9",X"DD",X"CE",X"00",
		X"FF",X"09",X"DE",X"CE",X"00",X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",X"76",X"11",X"8D",X"84",
		X"48",X"D8",X"11",X"78",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"76",X"11",X"18",
		X"85",X"58",X"81",X"11",X"78",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"76",X"BB",
		X"B8",X"86",X"68",X"8B",X"BB",X"78",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"86",
		X"CC",X"C0",X"00",X"00",X"0C",X"CC",X"78",X"00",X"00",X"00",X"00",X"FF",X"00",X"77",X"00",X"FF",
		X"07",X"88",X"70",X"FF",X"78",X"88",X"87",X"FF",X"78",X"91",X"87",X"FF",X"78",X"59",X"87",X"FF",
		X"78",X"88",X"87",X"FF",X"07",X"88",X"70",X"FF",X"00",X"77",X"00",X"FF",X"00",X"00",X"07",X"70",
		X"00",X"00",X"FF",X"00",X"07",X"7E",X"E7",X"70",X"00",X"FF",X"00",X"7E",X"E8",X"8E",X"E7",X"00",
		X"FF",X"07",X"E8",X"88",X"88",X"8E",X"70",X"FF",X"07",X"E8",X"88",X"88",X"8E",X"70",X"FF",X"7E",
		X"88",X"88",X"88",X"88",X"E7",X"FF",X"7E",X"88",X"85",X"58",X"88",X"E7",X"FF",X"7E",X"88",X"85",
		X"58",X"88",X"E7",X"FF",X"7E",X"88",X"88",X"88",X"88",X"E7",X"FF",X"07",X"E8",X"88",X"88",X"8E",
		X"70",X"FF",X"07",X"E8",X"88",X"88",X"8E",X"70",X"FF",X"00",X"7E",X"E8",X"8E",X"E7",X"00",X"FF",
		X"00",X"07",X"7E",X"E7",X"70",X"00",X"FF",X"00",X"00",X"07",X"70",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"77",X"77",X"00",X"00",X"00",X"FF",X"00",X"00",X"77",X"EE",X"CC",X"77",X"00",X"00",X"FF",
		X"00",X"07",X"DE",X"EE",X"CC",X"CD",X"70",X"00",X"FF",X"00",X"7D",X"55",X"22",X"22",X"5D",X"D7",
		X"00",X"FF",X"07",X"D5",X"52",X"88",X"88",X"2D",X"DD",X"70",X"FF",X"07",X"CC",X"28",X"88",X"88",
		X"82",X"DE",X"70",X"FF",X"7C",X"CC",X"28",X"88",X"88",X"82",X"EE",X"E7",X"FF",X"7C",X"C2",X"88",
		X"89",X"B8",X"88",X"2E",X"E7",X"FF",X"7C",X"C2",X"88",X"94",X"4B",X"88",X"2E",X"E7",X"FF",X"7E",
		X"E2",X"88",X"94",X"1B",X"88",X"2C",X"C7",X"FF",X"7E",X"E2",X"88",X"89",X"B8",X"88",X"2C",X"C7",
		X"FF",X"7E",X"EE",X"28",X"88",X"88",X"82",X"CC",X"C7",X"FF",X"07",X"ED",X"28",X"88",X"88",X"82",
		X"CC",X"70",X"FF",X"07",X"D5",X"52",X"88",X"88",X"25",X"55",X"70",X"FF",X"00",X"7D",X"55",X"22",
		X"22",X"55",X"D7",X"00",X"FF",X"00",X"07",X"DC",X"CC",X"EE",X"ED",X"70",X"00",X"FF",X"00",X"00",
		X"77",X"CC",X"EE",X"77",X"00",X"00",X"FF",X"00",X"00",X"00",X"77",X"77",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"FF",X"00",X"00",X"08",X"87",X"99",
		X"99",X"78",X"80",X"00",X"00",X"FF",X"00",X"00",X"87",X"99",X"EE",X"CC",X"99",X"78",X"00",X"00",
		X"FF",X"00",X"08",X"79",X"EE",X"EE",X"CC",X"CC",X"97",X"80",X"00",X"FF",X"00",X"87",X"9D",X"EE",
		X"E9",X"9C",X"CC",X"D9",X"78",X"00",X"FF",X"08",X"79",X"DD",X"D2",X"88",X"88",X"8D",X"DD",X"97",
		X"80",X"FF",X"08",X"9D",X"DD",X"28",X"88",X"88",X"88",X"DD",X"D9",X"80",X"FF",X"87",X"9C",X"D2",
		X"88",X"88",X"88",X"88",X"8D",X"E9",X"78",X"FF",X"89",X"CC",X"C2",X"88",X"88",X"88",X"88",X"8E",
		X"EE",X"98",X"FF",X"79",X"CC",X"28",X"88",X"88",X"88",X"88",X"88",X"EE",X"97",X"FF",X"7C",X"CC",
		X"28",X"88",X"69",X"B8",X"88",X"88",X"EE",X"E7",X"FF",X"7C",X"C9",X"88",X"86",X"94",X"4B",X"88",
		X"88",X"9E",X"E7",X"FF",X"7E",X"E9",X"88",X"86",X"94",X"41",X"88",X"88",X"9C",X"C7",X"FF",X"7E",
		X"EE",X"28",X"86",X"69",X"B8",X"88",X"88",X"CC",X"C7",X"FF",X"79",X"EE",X"28",X"88",X"66",X"68",
		X"88",X"88",X"CC",X"97",X"FF",X"89",X"EE",X"E2",X"88",X"88",X"88",X"88",X"8C",X"CC",X"98",X"FF",
		X"87",X"9E",X"D2",X"88",X"88",X"88",X"88",X"8D",X"C9",X"78",X"FF",X"08",X"9D",X"DD",X"28",X"88",
		X"88",X"88",X"DD",X"D9",X"80",X"FF",X"08",X"79",X"DD",X"D2",X"88",X"88",X"8D",X"DD",X"97",X"80",
		X"FF",X"00",X"87",X"9D",X"CC",X"C9",X"9E",X"EE",X"D9",X"78",X"00",X"FF",X"00",X"08",X"79",X"CC",
		X"CC",X"EE",X"EE",X"97",X"80",X"00",X"FF",X"00",X"00",X"87",X"99",X"CC",X"EE",X"99",X"78",X"00",
		X"00",X"FF",X"00",X"00",X"08",X"87",X"99",X"99",X"78",X"80",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"88",X"88",X"88",X"88",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"08",X"87",X"99",X"99",X"78",X"80",X"00",X"00",X"FF",X"00",X"00",
		X"87",X"99",X"EE",X"CC",X"99",X"78",X"00",X"00",X"FF",X"00",X"08",X"79",X"EE",X"EE",X"CC",X"CC",
		X"97",X"80",X"00",X"FF",X"00",X"87",X"9D",X"EE",X"E9",X"9C",X"CC",X"D9",X"78",X"00",X"FF",X"08",
		X"79",X"DD",X"D2",X"88",X"88",X"8D",X"DD",X"97",X"80",X"FF",X"08",X"9D",X"DD",X"28",X"88",X"88",
		X"88",X"DD",X"D9",X"80",X"FF",X"87",X"9C",X"D2",X"88",X"88",X"88",X"88",X"8D",X"E9",X"78",X"FF",
		X"89",X"CC",X"C2",X"88",X"66",X"68",X"88",X"8E",X"EE",X"98",X"FF",X"79",X"CC",X"28",X"86",X"BB",
		X"BB",X"88",X"88",X"EE",X"97",X"FF",X"7C",X"CC",X"28",X"6B",X"B3",X"3B",X"B8",X"88",X"EE",X"E7",
		X"FF",X"7C",X"C9",X"86",X"69",X"94",X"93",X"B8",X"88",X"9E",X"E7",X"FF",X"7E",X"E9",X"86",X"69",
		X"94",X"91",X"38",X"88",X"9C",X"C7",X"FF",X"7E",X"EE",X"26",X"6B",X"33",X"33",X"B8",X"88",X"CC",
		X"C7",X"FF",X"79",X"EE",X"26",X"66",X"B3",X"3B",X"88",X"88",X"CC",X"97",X"FF",X"89",X"EE",X"E2",
		X"66",X"66",X"68",X"88",X"8C",X"CC",X"98",X"FF",X"87",X"9E",X"D2",X"86",X"66",X"88",X"88",X"8D",
		X"C9",X"78",X"FF",X"08",X"9D",X"DD",X"28",X"88",X"88",X"88",X"DD",X"D9",X"80",X"FF",X"08",X"79",
		X"DD",X"D2",X"88",X"88",X"8D",X"DD",X"97",X"80",X"FF",X"00",X"87",X"9D",X"CC",X"C9",X"9E",X"EE",
		X"D9",X"78",X"00",X"FF",X"00",X"08",X"79",X"CC",X"CC",X"EE",X"EE",X"97",X"80",X"00",X"FF",X"00",
		X"00",X"87",X"99",X"CC",X"EE",X"99",X"78",X"00",X"00",X"FF",X"00",X"00",X"08",X"87",X"99",X"99",
		X"78",X"80",X"00",X"00",X"FF",X"00",X"00",X"00",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"FF",X"00",X"00",X"08",X"87",X"99",
		X"99",X"78",X"80",X"00",X"00",X"FF",X"00",X"00",X"87",X"99",X"EE",X"CC",X"99",X"78",X"00",X"00",
		X"FF",X"00",X"08",X"79",X"EE",X"EE",X"CC",X"CC",X"97",X"80",X"00",X"FF",X"00",X"87",X"9D",X"EE",
		X"E9",X"9C",X"CC",X"D9",X"78",X"00",X"FF",X"08",X"79",X"DD",X"D2",X"88",X"88",X"8D",X"DD",X"97",
		X"80",X"FF",X"08",X"9D",X"DD",X"28",X"88",X"88",X"88",X"DD",X"D9",X"80",X"FF",X"87",X"9C",X"D2",
		X"86",X"BB",X"BB",X"88",X"8D",X"E9",X"78",X"FF",X"89",X"CC",X"C8",X"6B",X"BB",X"BB",X"B8",X"8E",
		X"EE",X"98",X"FF",X"79",X"CC",X"86",X"6B",X"B3",X"13",X"B8",X"88",X"EE",X"97",X"FF",X"7C",X"CC",
		X"86",X"BB",X"34",X"44",X"3B",X"88",X"EE",X"E7",X"FF",X"7C",X"C9",X"66",X"99",X"95",X"94",X"3B",
		X"88",X"9E",X"E7",X"FF",X"7E",X"E9",X"66",X"99",X"94",X"94",X"1B",X"88",X"9C",X"C7",X"FF",X"7E",
		X"EE",X"86",X"B3",X"44",X"45",X"4B",X"88",X"CC",X"C7",X"FF",X"79",X"EE",X"86",X"6B",X"34",X"14",
		X"B8",X"88",X"CC",X"97",X"FF",X"89",X"EE",X"E8",X"6B",X"33",X"33",X"B8",X"8C",X"CC",X"98",X"FF",
		X"87",X"9E",X"D8",X"66",X"BB",X"BB",X"88",X"8D",X"C9",X"78",X"FF",X"08",X"9D",X"DD",X"86",X"66",
		X"68",X"88",X"DD",X"D9",X"80",X"FF",X"08",X"79",X"DD",X"D8",X"88",X"88",X"8D",X"DD",X"97",X"80",
		X"FF",X"00",X"87",X"9D",X"CC",X"C9",X"9E",X"EE",X"D9",X"78",X"00",X"FF",X"00",X"08",X"79",X"CC",
		X"CC",X"EE",X"EE",X"97",X"80",X"00",X"FF",X"00",X"00",X"87",X"99",X"CC",X"EE",X"99",X"78",X"00",
		X"00",X"FF",X"00",X"00",X"08",X"87",X"99",X"99",X"78",X"80",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"88",X"88",X"88",X"88",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"08",X"87",X"99",X"99",X"78",X"80",X"00",X"00",X"FF",X"00",X"00",
		X"87",X"99",X"EE",X"CC",X"99",X"78",X"00",X"00",X"FF",X"00",X"08",X"79",X"EE",X"EE",X"CC",X"CC",
		X"97",X"80",X"00",X"FF",X"00",X"87",X"9D",X"EE",X"E9",X"9C",X"CC",X"D9",X"78",X"00",X"FF",X"08",
		X"79",X"DD",X"D8",X"88",X"88",X"8D",X"DD",X"97",X"80",X"FF",X"08",X"9D",X"DD",X"88",X"BB",X"BB",
		X"88",X"DD",X"D9",X"80",X"FF",X"87",X"9C",X"D8",X"6B",X"33",X"44",X"B8",X"8D",X"E9",X"78",X"FF",
		X"89",X"CC",X"C6",X"BB",X"44",X"14",X"3B",X"8E",X"EE",X"98",X"FF",X"79",X"CC",X"86",X"B3",X"45",
		X"55",X"4B",X"88",X"EE",X"97",X"FF",X"7C",X"CC",X"6B",X"B4",X"59",X"95",X"53",X"B8",X"EE",X"E7",
		X"FF",X"7C",X"C9",X"69",X"99",X"90",X"59",X"54",X"B8",X"9E",X"E7",X"FF",X"7E",X"E9",X"69",X"99",
		X"90",X"59",X"51",X"B8",X"9C",X"C7",X"FF",X"7E",X"EE",X"6B",X"B4",X"59",X"95",X"54",X"B8",X"CC",
		X"C7",X"FF",X"79",X"EE",X"86",X"B4",X"45",X"55",X"4B",X"88",X"CC",X"97",X"FF",X"89",X"EE",X"E6",
		X"B3",X"44",X"14",X"4B",X"8C",X"CC",X"98",X"FF",X"87",X"9E",X"D8",X"6B",X"44",X"44",X"B8",X"8D",
		X"C9",X"78",X"FF",X"08",X"9D",X"DD",X"86",X"BB",X"BB",X"88",X"DD",X"D9",X"80",X"FF",X"08",X"79",
		X"DD",X"D8",X"66",X"68",X"8D",X"DD",X"97",X"80",X"FF",X"00",X"87",X"9D",X"CC",X"C9",X"9E",X"EE",
		X"D9",X"78",X"00",X"FF",X"00",X"08",X"79",X"CC",X"CC",X"EE",X"EE",X"97",X"80",X"00",X"FF",X"00",
		X"00",X"87",X"99",X"CC",X"EE",X"99",X"78",X"00",X"00",X"FF",X"00",X"00",X"08",X"87",X"99",X"99",
		X"78",X"80",X"00",X"00",X"FF",X"00",X"00",X"00",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"FF",X"00",X"00",X"08",X"87",X"99",
		X"99",X"78",X"80",X"00",X"00",X"FF",X"00",X"00",X"87",X"99",X"EE",X"CC",X"99",X"78",X"00",X"00",
		X"FF",X"00",X"08",X"79",X"EE",X"EE",X"CC",X"CC",X"97",X"80",X"00",X"FF",X"00",X"87",X"9D",X"EE",
		X"E9",X"9C",X"CC",X"D9",X"78",X"00",X"FF",X"08",X"79",X"DD",X"D6",X"33",X"33",X"8D",X"DD",X"97",
		X"80",X"FF",X"08",X"9D",X"DD",X"6B",X"BB",X"BB",X"33",X"DD",X"D9",X"80",X"FF",X"87",X"9C",X"D6",
		X"BB",X"33",X"13",X"BB",X"3D",X"E9",X"78",X"FF",X"89",X"CC",X"C6",X"B3",X"34",X"43",X"3B",X"BE",
		X"EE",X"98",X"FF",X"79",X"CC",X"6B",X"B3",X"44",X"44",X"43",X"B3",X"EE",X"97",X"FF",X"7C",X"CC",
		X"69",X"B3",X"49",X"94",X"44",X"B3",X"EE",X"E7",X"FF",X"7C",X"C9",X"69",X"99",X"90",X"D9",X"45",
		X"B3",X"9E",X"E7",X"FF",X"7E",X"E9",X"69",X"99",X"90",X"D9",X"54",X"13",X"9C",X"C7",X"FF",X"7E",
		X"EE",X"69",X"B3",X"49",X"94",X"54",X"B3",X"CC",X"C7",X"FF",X"79",X"EE",X"6B",X"B3",X"44",X"55",
		X"43",X"B3",X"CC",X"97",X"FF",X"89",X"EE",X"E6",X"B3",X"34",X"44",X"3B",X"BC",X"CC",X"98",X"FF",
		X"87",X"9E",X"D6",X"BB",X"33",X"13",X"BB",X"3D",X"C9",X"78",X"FF",X"08",X"9D",X"DD",X"6B",X"BB",
		X"BB",X"B3",X"DD",X"D9",X"80",X"FF",X"08",X"79",X"DD",X"D6",X"33",X"33",X"3D",X"DD",X"97",X"80",
		X"FF",X"00",X"87",X"9D",X"CC",X"C9",X"9E",X"EE",X"D9",X"78",X"00",X"FF",X"00",X"08",X"79",X"CC",
		X"CC",X"EE",X"EE",X"97",X"80",X"00",X"FF",X"00",X"00",X"87",X"99",X"CC",X"EE",X"99",X"78",X"00",
		X"00",X"FF",X"00",X"00",X"08",X"87",X"99",X"99",X"78",X"80",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"88",X"88",X"88",X"88",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"08",X"87",X"99",X"99",X"78",X"80",X"00",X"00",X"FF",X"00",X"00",
		X"87",X"99",X"EE",X"CC",X"99",X"78",X"00",X"00",X"FF",X"00",X"08",X"79",X"EE",X"E3",X"3C",X"CC",
		X"97",X"80",X"00",X"FF",X"00",X"87",X"9D",X"EB",X"BB",X"BB",X"BC",X"D9",X"78",X"00",X"FF",X"08",
		X"79",X"DD",X"BB",X"B3",X"33",X"3B",X"DD",X"97",X"80",X"FF",X"08",X"9D",X"DB",X"B3",X"41",X"14",
		X"33",X"BD",X"D9",X"80",X"FF",X"87",X"9C",X"DB",X"34",X"45",X"55",X"43",X"BD",X"E9",X"78",X"FF",
		X"89",X"CC",X"B3",X"44",X"55",X"55",X"54",X"3B",X"EE",X"98",X"FF",X"79",X"CC",X"B3",X"45",X"99",
		X"99",X"55",X"4B",X"EE",X"97",X"FF",X"7C",X"C9",X"99",X"99",X"99",X"49",X"95",X"4B",X"3E",X"E7",
		X"FF",X"7C",X"C9",X"99",X"99",X"90",X"59",X"95",X"1B",X"3E",X"E7",X"FF",X"7E",X"E9",X"99",X"99",
		X"90",X"59",X"95",X"1B",X"3C",X"C7",X"FF",X"7E",X"E9",X"99",X"99",X"99",X"49",X"95",X"4B",X"3C",
		X"C7",X"FF",X"79",X"EE",X"BB",X"34",X"99",X"99",X"54",X"3B",X"CC",X"97",X"FF",X"89",X"EE",X"BB",
		X"34",X"45",X"55",X"43",X"3B",X"CC",X"98",X"FF",X"87",X"9E",X"DB",X"33",X"44",X"44",X"33",X"BD",
		X"C9",X"78",X"FF",X"08",X"9D",X"DB",X"B3",X"31",X"13",X"3B",X"BD",X"D9",X"80",X"FF",X"08",X"79",
		X"DD",X"BB",X"B3",X"3B",X"BB",X"DD",X"97",X"80",X"FF",X"00",X"87",X"9D",X"CB",X"BB",X"BB",X"BE",
		X"D9",X"78",X"00",X"FF",X"00",X"08",X"79",X"CC",X"C3",X"3E",X"EE",X"97",X"80",X"00",X"FF",X"00",
		X"00",X"87",X"99",X"CC",X"EE",X"99",X"78",X"00",X"00",X"FF",X"00",X"00",X"08",X"87",X"99",X"99",
		X"78",X"80",X"00",X"00",X"FF",X"00",X"00",X"00",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"FF",X"00",X"00",X"08",X"87",X"99",
		X"99",X"78",X"80",X"00",X"00",X"FF",X"00",X"00",X"87",X"99",X"EE",X"CC",X"99",X"78",X"00",X"00",
		X"FF",X"00",X"08",X"79",X"EE",X"E3",X"3C",X"CC",X"97",X"80",X"00",X"FF",X"00",X"87",X"9D",X"EB",
		X"BB",X"BB",X"BC",X"D9",X"78",X"00",X"FF",X"08",X"79",X"DD",X"BB",X"BB",X"BB",X"BB",X"DD",X"97",
		X"80",X"FF",X"08",X"9D",X"DB",X"BB",X"31",X"13",X"3B",X"BD",X"D9",X"80",X"FF",X"87",X"9C",X"DB",
		X"33",X"34",X"44",X"33",X"BD",X"E9",X"78",X"FF",X"89",X"CC",X"B3",X"34",X"55",X"55",X"43",X"BB",
		X"EE",X"98",X"FF",X"79",X"CC",X"B3",X"45",X"99",X"99",X"54",X"3B",X"EE",X"97",X"FF",X"7C",X"C3",
		X"B4",X"59",X"99",X"99",X"95",X"4B",X"3E",X"E7",X"FF",X"7C",X"C3",X"B1",X"59",X"45",X"54",X"95",
		X"1B",X"3E",X"E7",X"FF",X"7E",X"E3",X"B1",X"59",X"90",X"09",X"95",X"1B",X"3C",X"C7",X"FF",X"7E",
		X"E3",X"B5",X"59",X"99",X"99",X"95",X"5B",X"3C",X"C7",X"FF",X"79",X"EE",X"B4",X"55",X"99",X"99",
		X"55",X"3B",X"CC",X"97",X"FF",X"89",X"EE",X"B3",X"45",X"99",X"99",X"54",X"3B",X"CC",X"98",X"FF",
		X"87",X"9E",X"DB",X"34",X"99",X"99",X"44",X"BD",X"C9",X"78",X"FF",X"08",X"9D",X"DB",X"B3",X"99",
		X"99",X"3B",X"BD",X"D9",X"80",X"FF",X"08",X"79",X"DD",X"BB",X"99",X"99",X"BB",X"DD",X"97",X"80",
		X"FF",X"00",X"87",X"9D",X"CB",X"99",X"99",X"BE",X"D9",X"78",X"00",X"FF",X"00",X"08",X"79",X"CC",
		X"C9",X"9E",X"EE",X"97",X"80",X"00",X"FF",X"00",X"00",X"87",X"99",X"CC",X"EE",X"99",X"78",X"00",
		X"00",X"FF",X"00",X"00",X"08",X"87",X"99",X"99",X"78",X"80",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"88",X"88",X"88",X"88",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"08",X"87",X"99",X"99",X"78",X"80",X"00",X"00",X"FF",X"00",X"00",
		X"87",X"99",X"EE",X"CC",X"99",X"78",X"00",X"00",X"FF",X"00",X"08",X"79",X"EE",X"E3",X"3C",X"CC",
		X"97",X"80",X"00",X"FF",X"00",X"87",X"9D",X"EB",X"BB",X"BB",X"BC",X"D9",X"78",X"00",X"FF",X"08",
		X"79",X"DD",X"BB",X"33",X"3B",X"BB",X"DD",X"97",X"80",X"FF",X"08",X"9D",X"DB",X"B4",X"44",X"44",
		X"3B",X"BD",X"D9",X"80",X"FF",X"87",X"9C",X"DB",X"34",X"55",X"54",X"13",X"BD",X"E9",X"78",X"FF",
		X"89",X"CC",X"B3",X"41",X"55",X"55",X"41",X"3B",X"EE",X"98",X"FF",X"79",X"CC",X"B4",X"15",X"59",
		X"99",X"54",X"3B",X"EE",X"97",X"FF",X"7C",X"C3",X"B4",X"55",X"94",X"99",X"95",X"4B",X"3E",X"E7",
		X"FF",X"7C",X"C3",X"B4",X"59",X"90",X"59",X"95",X"4B",X"3E",X"E7",X"FF",X"7E",X"E3",X"B3",X"49",
		X"99",X"04",X"95",X"4B",X"3C",X"C7",X"FF",X"7E",X"E3",X"B4",X"99",X"99",X"99",X"55",X"4B",X"3C",
		X"C7",X"FF",X"79",X"EE",X"B9",X"99",X"99",X"95",X"54",X"3B",X"CC",X"97",X"FF",X"89",X"EE",X"99",
		X"99",X"99",X"54",X"41",X"BB",X"CC",X"98",X"FF",X"87",X"9E",X"D9",X"99",X"94",X"44",X"13",X"BD",
		X"C9",X"78",X"FF",X"08",X"9D",X"D9",X"99",X"33",X"33",X"3B",X"BD",X"D9",X"80",X"FF",X"08",X"79",
		X"DD",X"9B",X"B3",X"3B",X"BB",X"DD",X"97",X"80",X"FF",X"00",X"87",X"9D",X"C9",X"BB",X"BB",X"BE",
		X"D9",X"78",X"00",X"FF",X"00",X"08",X"79",X"CC",X"C3",X"3E",X"EE",X"97",X"80",X"00",X"FF",X"00",
		X"00",X"87",X"99",X"CC",X"EE",X"99",X"78",X"00",X"00",X"FF",X"00",X"00",X"08",X"87",X"99",X"99",
		X"78",X"80",X"00",X"00",X"FF",X"00",X"00",X"00",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"01",X"11",X"11",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"18",X"88",X"88",X"10",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"11",X"E5",X"A9",X"8E",X"00",X"00",X"00",X"FF",X"0E",X"EE",
		X"EE",X"76",X"55",X"22",X"E0",X"00",X"00",X"FF",X"16",X"66",X"37",X"43",X"13",X"35",X"9E",X"EE",
		X"10",X"FF",X"15",X"53",X"64",X"36",X"14",X"43",X"59",X"99",X"10",X"FF",X"0E",X"E6",X"43",X"46",
		X"15",X"55",X"25",X"E1",X"10",X"FF",X"14",X"47",X"34",X"44",X"17",X"75",X"22",X"55",X"10",X"FF",
		X"16",X"57",X"11",X"11",X"11",X"11",X"11",X"5D",X"50",X"FF",X"14",X"46",X"22",X"44",X"17",X"65",
		X"11",X"4D",X"40",X"FF",X"13",X"36",X"12",X"45",X"15",X"33",X"22",X"44",X"E0",X"FF",X"1E",X"E6",
		X"41",X"26",X"13",X"31",X"14",X"EE",X"10",X"FF",X"15",X"52",X"54",X"12",X"13",X"11",X"4A",X"AA",
		X"10",X"FF",X"14",X"44",X"25",X"33",X"11",X"44",X"AE",X"EE",X"00",X"FF",X"1E",X"EE",X"EE",X"44",
		X"44",X"11",X"E1",X"00",X"00",X"FF",X"11",X"11",X"11",X"E4",X"BA",X"8E",X"10",X"00",X"00",X"FF",
		X"00",X"00",X"08",X"88",X"88",X"10",X"00",X"00",X"00",X"FF",X"00",X"00",X"01",X"11",X"11",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"01",X"11",X"11",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"18",X"88",X"88",X"10",X"00",X"00",X"00",X"FF",X"00",X"00",X"11",X"E5",X"A9",X"8E",X"00",X"00",
		X"00",X"FF",X"0E",X"EE",X"EE",X"76",X"45",X"22",X"E0",X"00",X"00",X"FF",X"16",X"66",X"37",X"43",
		X"E3",X"35",X"9E",X"EE",X"10",X"FF",X"15",X"53",X"64",X"35",X"14",X"43",X"59",X"99",X"10",X"FF",
		X"0E",X"E6",X"43",X"45",X"15",X"55",X"25",X"E1",X"10",X"FF",X"14",X"47",X"34",X"51",X"ED",X"77",
		X"22",X"55",X"10",X"FF",X"16",X"57",X"EE",X"11",X"DD",X"EE",X"11",X"5D",X"50",X"FF",X"14",X"46",
		X"22",X"41",X"ED",X"74",X"11",X"4D",X"40",X"FF",X"13",X"36",X"12",X"45",X"15",X"33",X"22",X"44",
		X"E0",X"FF",X"1E",X"E6",X"41",X"26",X"E3",X"31",X"14",X"EE",X"10",X"FF",X"15",X"52",X"54",X"12",
		X"E3",X"11",X"4A",X"AA",X"10",X"FF",X"14",X"44",X"25",X"33",X"E1",X"44",X"AE",X"EE",X"00",X"FF",
		X"1E",X"EE",X"EE",X"44",X"44",X"11",X"E1",X"00",X"00",X"FF",X"11",X"11",X"11",X"E4",X"BA",X"8E",
		X"10",X"00",X"00",X"FF",X"00",X"00",X"08",X"88",X"88",X"10",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"01",X"11",X"11",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"01",X"11",X"11",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"18",X"88",X"88",X"10",X"00",X"00",X"00",X"FF",X"00",X"00",X"11",X"E5",
		X"99",X"8E",X"00",X"00",X"00",X"FF",X"0E",X"EE",X"EE",X"76",X"45",X"22",X"E0",X"00",X"00",X"FF",
		X"16",X"66",X"37",X"23",X"E3",X"35",X"9E",X"EE",X"10",X"FF",X"15",X"53",X"42",X"35",X"E4",X"74",
		X"59",X"98",X"10",X"FF",X"0E",X"E6",X"23",X"4D",X"CD",X"47",X"55",X"E1",X"10",X"FF",X"14",X"47",
		X"34",X"DC",X"BC",X"D4",X"42",X"55",X"10",X"FF",X"16",X"57",X"ED",X"CB",X"AB",X"CD",X"E1",X"5B",
		X"50",X"FF",X"14",X"46",X"ED",X"CB",X"AB",X"CD",X"E1",X"4B",X"40",X"FF",X"13",X"36",X"24",X"DC",
		X"BC",X"D4",X"22",X"44",X"E0",X"FF",X"1E",X"E6",X"42",X"4D",X"CD",X"43",X"14",X"EE",X"10",X"FF",
		X"15",X"52",X"54",X"22",X"E4",X"21",X"49",X"98",X"10",X"FF",X"14",X"44",X"25",X"33",X"E1",X"44",
		X"9E",X"EE",X"00",X"FF",X"1E",X"EE",X"EE",X"44",X"44",X"11",X"E1",X"00",X"00",X"FF",X"11",X"11",
		X"11",X"E4",X"99",X"8E",X"10",X"00",X"00",X"FF",X"00",X"00",X"08",X"88",X"88",X"10",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"01",X"11",X"11",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"22",X"20",X"12",X"00",X"00",X"00",X"00",X"FF",X"01",X"20",X"02",X"10",X"01",X"12",X"11",X"10",
		X"11",X"00",X"10",X"FF",X"02",X"01",X"11",X"11",X"11",X"11",X"11",X"11",X"20",X"11",X"00",X"FF",
		X"00",X"11",X"11",X"11",X"22",X"31",X"33",X"11",X"11",X"13",X"10",X"FF",X"02",X"11",X"11",X"31",
		X"22",X"11",X"31",X"13",X"31",X"13",X"11",X"FF",X"21",X"13",X"33",X"33",X"33",X"44",X"42",X"11",
		X"11",X"11",X"00",X"FF",X"01",X"23",X"33",X"24",X"33",X"33",X"43",X"44",X"33",X"11",X"20",X"FF",
		X"02",X"31",X"32",X"24",X"34",X"44",X"44",X"43",X"33",X"31",X"10",X"FF",X"21",X"13",X"44",X"44",
		X"44",X"44",X"44",X"43",X"33",X"11",X"10",X"FF",X"11",X"43",X"33",X"44",X"45",X"55",X"54",X"44",
		X"44",X"33",X"12",X"FF",X"31",X"43",X"35",X"55",X"55",X"55",X"55",X"54",X"43",X"43",X"12",X"FF",
		X"31",X"44",X"55",X"55",X"56",X"66",X"55",X"55",X"44",X"43",X"31",X"FF",X"44",X"45",X"55",X"56",
		X"66",X"66",X"66",X"65",X"54",X"44",X"33",X"FF",X"45",X"45",X"56",X"66",X"66",X"00",X"66",X"66",
		X"65",X"44",X"33",X"FF",X"36",X"66",X"66",X"60",X"00",X"00",X"00",X"06",X"66",X"55",X"63",X"FF",
		X"66",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"FF",X"1D",X"DE",X"11",X"11",
		X"00",X"FF",X"00",X"00",X"0D",X"4E",X"10",X"00",X"00",X"FF",X"00",X"00",X"00",X"31",X"10",X"00",
		X"00",X"FF",X"00",X"00",X"06",X"36",X"11",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"D0",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"06",X"AC",X"00",X"6A",X"FF",X"00",X"00",X"00",X"06",X"9B",X"6C",
		X"A6",X"FF",X"00",X"00",X"00",X"66",X"49",X"C6",X"C6",X"FF",X"00",X"00",X"06",X"66",X"26",X"A6",
		X"60",X"FF",X"00",X"8D",X"DD",X"D6",X"14",X"AA",X"00",X"FF",X"53",X"13",X"99",X"96",X"22",X"38",
		X"3A",X"FF",X"CB",X"8B",X"DA",X"D6",X"36",X"49",X"9B",X"FF",X"06",X"BB",X"BB",X"B6",X"88",X"9B",
		X"66",X"FF",X"66",X"66",X"66",X"66",X"89",X"A6",X"66",X"FF",X"66",X"66",X"66",X"E6",X"96",X"B6",
		X"E0",X"FF",X"06",X"66",X"66",X"6D",X"9A",X"66",X"BE",X"FF",X"00",X"00",X"66",X"6C",X"AC",X"66",
		X"EB",X"FF",X"00",X"00",X"06",X"66",X"C6",X"60",X"66",X"FF",X"00",X"00",X"06",X"66",X"66",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"66",X"60",X"00",X"00",X"FF",X"00",X"00",X"00",X"06",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"CA",X"00",X"00",X"00",X"FF",X"00",X"00",X"06",X"AD",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"66",X"EE",X"00",X"00",X"00",X"FF",X"0B",X"AA",X"AA",X"66",X"BA",X"00",
		X"00",X"FF",X"0B",X"A9",X"99",X"BC",X"A9",X"A0",X"00",X"FF",X"00",X"A9",X"76",X"84",X"9A",X"C0",
		X"00",X"FF",X"66",X"6B",X"21",X"37",X"9C",X"E0",X"00",X"FF",X"66",X"66",X"B2",X"16",X"9B",X"6D",
		X"A0",X"FF",X"66",X"66",X"C6",X"28",X"9A",X"CA",X"D0",X"FF",X"66",X"6C",X"7B",X"B7",X"96",X"C6",
		X"60",X"FF",X"D6",X"CB",X"7C",X"AB",X"9A",X"B6",X"00",X"FF",X"C6",X"B4",X"AB",X"66",X"B9",X"B0",
		X"00",X"FF",X"0B",X"17",X"CB",X"66",X"6C",X"C0",X"00",X"FF",X"09",X"1D",X"B6",X"66",X"66",X"00",
		X"00",X"FF",X"08",X"9B",X"66",X"66",X"66",X"00",X"00",X"FF",X"65",X"A6",X"66",X"66",X"00",X"00",
		X"00",X"FF",X"65",X"B6",X"60",X"00",X"00",X"00",X"00",X"FF",X"66",X"66",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"66",X"60",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0C",X"BB",X"A0",
		X"00",X"00",X"FF",X"00",X"00",X"B6",X"6D",X"A9",X"A0",X"6B",X"00",X"FF",X"00",X"00",X"6B",X"6D",
		X"A9",X"A6",X"B6",X"00",X"FF",X"00",X"00",X"06",X"6B",X"B7",X"A6",X"60",X"00",X"FF",X"00",X"06",
		X"CB",X"AA",X"98",X"3A",X"A0",X"00",X"FF",X"00",X"6C",X"B6",X"99",X"68",X"36",X"8A",X"00",X"FF",
		X"06",X"CA",X"99",X"88",X"83",X"22",X"88",X"A0",X"FF",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"00",X"FF",X"06",X"66",X"66",X"6B",X"D9",X"C6",X"60",X"00",X"FF",X"00",X"66",X"66",X"6B",X"D9",
		X"C6",X"00",X"00",X"FF",X"00",X"00",X"66",X"6B",X"C9",X"C0",X"00",X"00",X"FF",X"00",X"00",X"06",
		X"6B",X"D9",X"C0",X"00",X"00",X"FF",X"00",X"00",X"06",X"6B",X"D4",X"A0",X"00",X"00",X"FF",X"00",
		X"00",X"06",X"6B",X"91",X"80",X"00",X"00",X"FF",X"00",X"00",X"06",X"6C",X"94",X"90",X"00",X"00",
		X"FF",X"00",X"00",X"06",X"6C",X"C5",X"90",X"00",X"00",X"FF",X"00",X"00",X"06",X"66",X"C5",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"88",X"80",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"66",X"AA",X"A0",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"66",X"66",X"00",X"CC",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"6E",X"AA",X"AA",X"A0",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"06",X"CC",X"E9",X"99",X"EA",X"0C",X"0C",X"00",X"FF",X"00",X"11",
		X"11",X"1C",X"BE",X"7E",X"27",X"EB",X"0B",X"00",X"FF",X"66",X"99",X"44",X"CC",X"55",X"E1",X"27",
		X"DA",X"DA",X"D0",X"FF",X"66",X"66",X"6D",X"CC",X"55",X"B1",X"27",X"69",X"69",X"B0",X"FF",X"00",
		X"11",X"11",X"CC",X"55",X"E2",X"37",X"DA",X"DA",X"D0",X"FF",X"66",X"99",X"44",X"7C",X"BE",X"8E",
		X"37",X"EB",X"6B",X"00",X"FF",X"66",X"66",X"66",X"DC",X"E9",X"99",X"EA",X"6C",X"6C",X"00",X"FF",
		X"00",X"00",X"66",X"6E",X"AA",X"AA",X"A6",X"66",X"00",X"00",X"FF",X"00",X"00",X"06",X"66",X"CC",
		X"CC",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"66",X"66",X"60",X"EE",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"99",X"96",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"66",
		X"BB",X"B0",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"66",X"60",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"FF",X"00",X"00",X"98",X"0C",X"C0",
		X"0B",X"A9",X"60",X"FF",X"00",X"09",X"8B",X"0D",X"00",X"BA",X"6A",X"A0",X"FF",X"00",X"98",X"B0",
		X"CA",X"E8",X"6B",X"86",X"B0",X"FF",X"00",X"0B",X"0D",X"A9",X"E4",X"86",X"BA",X"B0",X"FF",X"00",
		X"00",X"CA",X"98",X"E2",X"28",X"6B",X"00",X"FF",X"00",X"00",X"EE",X"EE",X"E1",X"14",X"8B",X"00",
		X"FF",X"00",X"06",X"CC",X"C5",X"5E",X"EE",X"E0",X"00",X"FF",X"00",X"66",X"C9",X"C5",X"5E",X"89",
		X"A0",X"00",X"FF",X"00",X"66",X"8A",X"C5",X"5E",X"9A",X"B0",X"D0",X"FF",X"00",X"61",X"8A",X"EC",
		X"CE",X"AB",X"CE",X"D0",X"FF",X"00",X"18",X"9E",X"8A",X"DE",X"BC",X"60",X"00",X"FF",X"01",X"89",
		X"61",X"8A",X"DE",X"C6",X"69",X"00",X"FF",X"08",X"96",X"18",X"9E",X"EE",X"66",X"9A",X"00",X"FF",
		X"66",X"61",X"89",X"66",X"66",X"69",X"AC",X"00",X"FF",X"66",X"08",X"96",X"66",X"66",X"0A",X"C0",
		X"00",X"FF",X"00",X"66",X"60",X"00",X"00",X"0C",X"00",X"00",X"FF",X"00",X"66",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"06",X"EC",X"E0",X"00",X"00",X"FF",X"00",X"00",X"6B",X"A9",
		X"AB",X"00",X"00",X"FF",X"00",X"00",X"06",X"EC",X"E0",X"00",X"00",X"FF",X"00",X"00",X"6B",X"A9",
		X"AB",X"00",X"00",X"FF",X"00",X"00",X"6E",X"CE",X"CE",X"00",X"00",X"FF",X"06",X"C0",X"6E",X"AA",
		X"AE",X"06",X"C0",X"FF",X"06",X"C6",X"CE",X"99",X"9E",X"96",X"C0",X"FF",X"06",X"6C",X"AE",X"88",
		X"8E",X"39",X"00",X"FF",X"0B",X"6B",X"A9",X"EE",X"E1",X"24",X"67",X"FF",X"6B",X"6B",X"99",X"EB",
		X"E1",X"14",X"67",X"FF",X"6B",X"6A",X"9E",X"55",X"5E",X"14",X"67",X"FF",X"6B",X"6A",X"EB",X"55",
		X"5B",X"E4",X"67",X"FF",X"06",X"6E",X"CC",X"CC",X"CC",X"CE",X"00",X"FF",X"00",X"66",X"C8",X"CC",
		X"C2",X"C0",X"00",X"FF",X"00",X"06",X"68",X"2D",X"82",X"00",X"00",X"FF",X"00",X"06",X"68",X"16",
		X"81",X"00",X"00",X"FF",X"00",X"06",X"69",X"16",X"91",X"00",X"00",X"FF",X"00",X"06",X"69",X"16",
		X"91",X"00",X"00",X"FF",X"00",X"06",X"69",X"16",X"91",X"00",X"00",X"FF",X"0A",X"A0",X"FF",X"A9",
		X"9A",X"FF",X"A8",X"8A",X"FF",X"A9",X"9A",X"FF",X"0A",X"A0",X"FF",X"00",X"99",X"00",X"FF",X"09",
		X"88",X"90",X"FF",X"09",X"55",X"90",X"FF",X"95",X"55",X"59",X"FF",X"09",X"55",X"90",X"FF",X"09",
		X"88",X"90",X"FF",X"00",X"99",X"00",X"FF",X"00",X"77",X"70",X"00",X"FF",X"07",X"66",X"67",X"00",
		X"FF",X"07",X"43",X"47",X"00",X"FF",X"76",X"21",X"26",X"70",X"FF",X"76",X"21",X"26",X"70",X"FF",
		X"05",X"43",X"47",X"00",X"FF",X"07",X"66",X"67",X"00",X"FF",X"00",X"77",X"70",X"00",X"FF",X"00",
		X"88",X"80",X"00",X"FF",X"08",X"55",X"58",X"00",X"FF",X"05",X"33",X"35",X"00",X"FF",X"83",X"22",
		X"23",X"80",X"FF",X"82",X"11",X"12",X"80",X"FF",X"82",X"11",X"12",X"80",X"FF",X"83",X"22",X"23",
		X"80",X"FF",X"05",X"33",X"35",X"00",X"FF",X"08",X"55",X"58",X"00",X"FF",X"00",X"88",X"80",X"00",
		X"FF",X"0E",X"E0",X"FF",X"EE",X"EE",X"FF",X"EE",X"EE",X"FF",X"EE",X"EE",X"FF",X"0E",X"E0",X"FF",
		X"01",X"10",X"FF",X"11",X"11",X"FF",X"11",X"11",X"FF",X"11",X"11",X"FF",X"01",X"10",X"FF",X"00",
		X"10",X"00",X"FF",X"00",X"20",X"00",X"FF",X"00",X"4A",X"01",X"FF",X"1A",X"AA",X"A0",X"FF",X"0A",
		X"A2",X"10",X"FF",X"02",X"AA",X"A0",X"FF",X"10",X"A4",X"01",X"FF",X"00",X"02",X"00",X"FF",X"00",
		X"01",X"00",X"FF",X"00",X"00",X"01",X"10",X"00",X"00",X"FF",X"00",X"00",X"04",X"40",X"00",X"00",
		X"FF",X"00",X"00",X"07",X"70",X"01",X"10",X"FF",X"00",X"00",X"00",X"00",X"08",X"10",X"FF",X"11",
		X"04",X"40",X"44",X"00",X"00",X"FF",X"14",X"04",X"A0",X"A4",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0A",X"40",X"41",X"FF",X"00",X"04",X"A0",X"04",X"40",
		X"41",X"FF",X"00",X"04",X"40",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"A4",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"44",X"00",X"00",X"FF",X"18",X"00",X"00",X"00",X"08",X"10",X"FF",X"11",X"00",
		X"00",X"00",X"01",X"10",X"FF",X"00",X"00",X"00",X"77",X"00",X"00",X"FF",X"00",X"00",X"00",X"44",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"11",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"04",X"40",X"00",X"00",X"00",X"04",X"40",X"00",X"FF",X"00",X"04",X"50",X"00",
		X"00",X"00",X"54",X"40",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"95",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"01",X"10",X"00",X"14",X"00",X"00",X"00",X"FF",X"45",X"90",
		X"01",X"40",X"00",X"00",X"00",X"09",X"54",X"FF",X"45",X"90",X"00",X"00",X"00",X"00",X"00",X"09",
		X"44",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"05",X"10",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"15",X"00",X"01",X"10",X"00",X"00",X"FF",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"45",
		X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"FF",X"00",X"44",X"00",X"00",X"00",X"00",X"05",X"40",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"40",X"00",X"FF",X"00",X"00",X"00",X"09",
		X"90",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"05",X"50",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"04",X"40",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"0E",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"0C",X"B0",X"00",X"00",X"00",X"00",X"CE",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"BC",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"EB",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"EB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BE",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"CB",
		X"00",X"00",X"00",X"00",X"0B",X"C0",X"00",X"FF",X"00",X"EC",X"00",X"00",X"00",X"00",X"0C",X"E0",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"FF",X"0D",X"AA",X"FF",X"ED",X"CC",X"FF",
		X"ED",X"CC",X"FF",X"EE",X"E0",X"FF",X"00",X"D0",X"FF",X"0D",X"DA",X"FF",X"ED",X"CA",X"FF",X"EC",
		X"CC",X"FF",X"EE",X"C0",X"FF",X"00",X"A0",X"FF",X"0A",X"AA",X"FF",X"0D",X"AC",X"FF",X"ED",X"DC",
		X"FF",X"EE",X"D0",X"FF",X"0D",X"AA",X"FF",X"0D",X"AA",X"FF",X"ED",X"CC",X"FF",X"EE",X"CC",X"FF",
		X"EE",X"E0",X"FF",X"00",X"D0",X"FF",X"0D",X"DA",X"FF",X"0D",X"CA",X"FF",X"EC",X"CC",X"FF",X"EC",
		X"CC",X"FF",X"EE",X"C0",X"FF",X"00",X"A0",X"FF",X"0A",X"AA",X"FF",X"0A",X"AA",X"FF",X"ED",X"AC",
		X"FF",X"ED",X"CC",X"FF",X"EE",X"C0",X"FF",X"0D",X"AA",X"A0",X"FF",X"0D",X"CC",X"C0",X"FF",X"0D",
		X"CC",X"C0",X"FF",X"ED",X"CC",X"C0",X"FF",X"EE",X"CC",X"C0",X"FF",X"EE",X"EE",X"00",X"FF",X"00",
		X"00",X"B0",X"00",X"FF",X"00",X"0B",X"BB",X"00",X"FF",X"00",X"BB",X"BB",X"B0",X"FF",X"00",X"DA",
		X"BB",X"C0",X"FF",X"0E",X"DD",X"AC",X"C0",X"FF",X"EE",X"DD",X"CC",X"C0",X"FF",X"0E",X"ED",X"CC",
		X"00",X"FF",X"00",X"EE",X"C0",X"00",X"FF",X"00",X"00",X"D0",X"00",X"FF",X"00",X"0D",X"DA",X"00",
		X"FF",X"00",X"DD",X"CA",X"A0",X"FF",X"0E",X"DC",X"CC",X"A0",X"FF",X"EE",X"CC",X"CC",X"C0",X"FF",
		X"EE",X"EC",X"CC",X"00",X"FF",X"0E",X"EE",X"C0",X"00",X"FF",X"00",X"0D",X"00",X"00",X"FF",X"00",
		X"DD",X"A0",X"00",X"FF",X"0D",X"DD",X"AA",X"00",X"FF",X"DD",X"DC",X"AA",X"A0",X"FF",X"DD",X"CC",
		X"CA",X"A0",X"FF",X"DC",X"CC",X"CC",X"A0",X"FF",X"CC",X"CC",X"CC",X"C0",X"FF",X"0C",X"CC",X"CC",
		X"00",X"FF",X"00",X"CC",X"C0",X"00",X"FF",X"00",X"0C",X"00",X"00",X"FF",X"00",X"0A",X"00",X"00",
		X"FF",X"00",X"AA",X"A0",X"00",X"FF",X"0A",X"AA",X"AA",X"00",X"FF",X"BA",X"AA",X"AA",X"B0",X"FF",
		X"DB",X"AA",X"AB",X"C0",X"FF",X"DD",X"BA",X"BC",X"C0",X"FF",X"DD",X"DB",X"CC",X"C0",X"FF",X"DD",
		X"DC",X"CC",X"C0",X"FF",X"0D",X"DC",X"CC",X"00",X"FF",X"00",X"DC",X"C0",X"00",X"FF",X"00",X"0C",
		X"00",X"00",X"FF",X"AA",X"AA",X"80",X"FF",X"DA",X"AA",X"A8",X"FF",X"DD",X"CC",X"CC",X"FF",X"DD",
		X"CC",X"CC",X"FF",X"DD",X"CC",X"CC",X"FF",X"DD",X"CC",X"CC",X"FF",X"0D",X"CC",X"CC",X"FF",X"AA",
		X"AA",X"AA",X"00",X"FF",X"DA",X"AA",X"AA",X"A0",X"FF",X"DD",X"AA",X"AA",X"AA",X"FF",X"DD",X"CC",
		X"CC",X"CC",X"FF",X"DD",X"CC",X"CC",X"CC",X"FF",X"DD",X"CC",X"CC",X"CC",X"FF",X"DD",X"CC",X"CC",
		X"CC",X"FF",X"DD",X"CC",X"CC",X"CC",X"FF",X"0D",X"CC",X"CC",X"CC",X"FF",X"00",X"CC",X"CC",X"CC",
		X"FF",X"00",X"00",X"A0",X"00",X"00",X"FF",X"00",X"0A",X"AA",X"00",X"00",X"FF",X"00",X"AA",X"AA",
		X"A0",X"00",X"FF",X"0A",X"AA",X"AA",X"AA",X"00",X"FF",X"BA",X"AA",X"AA",X"AA",X"B0",X"FF",X"DB",
		X"AA",X"AA",X"AB",X"C0",X"FF",X"DD",X"BA",X"AA",X"BC",X"C0",X"FF",X"DD",X"DB",X"AB",X"CC",X"C0",
		X"FF",X"DD",X"DD",X"BC",X"CC",X"C0",X"FF",X"DD",X"DD",X"CC",X"CC",X"C0",X"FF",X"DD",X"DD",X"CC",
		X"CC",X"C0",X"FF",X"0D",X"DD",X"CC",X"CC",X"00",X"FF",X"00",X"DD",X"CC",X"C0",X"00",X"FF",X"00",
		X"0D",X"CC",X"00",X"00",X"FF",X"00",X"00",X"C0",X"00",X"00",X"FF",X"00",X"00",X"D0",X"00",X"00",
		X"FF",X"00",X"0D",X"DA",X"00",X"00",X"FF",X"00",X"DD",X"DA",X"A0",X"00",X"FF",X"0D",X"DD",X"DA",
		X"AA",X"00",X"FF",X"DD",X"DD",X"CA",X"AA",X"A0",X"FF",X"DD",X"DC",X"CC",X"AA",X"A0",X"FF",X"DD",
		X"CC",X"CC",X"CA",X"A0",X"FF",X"DC",X"CC",X"CC",X"CC",X"A0",X"FF",X"CC",X"CC",X"CC",X"CC",X"C0",
		X"FF",X"0C",X"CC",X"CC",X"CC",X"00",X"FF",X"00",X"CC",X"CC",X"C0",X"00",X"FF",X"00",X"0C",X"CC",
		X"00",X"00",X"FF",X"00",X"00",X"C0",X"00",X"00",X"FF",X"AA",X"AA",X"AA",X"AA",X"BB",X"FF",X"01",
		X"11",X"11",X"11",X"B8",X"FF",X"00",X"00",X"99",X"99",X"40",X"FF",X"00",X"00",X"99",X"94",X"40",
		X"FF",X"00",X"09",X"99",X"94",X"00",X"FF",X"00",X"09",X"99",X"94",X"40",X"FF",X"00",X"00",X"99",
		X"99",X"40",X"FF",X"00",X"09",X"99",X"94",X"40",X"FF",X"AA",X"AA",X"AA",X"AA",X"BB",X"FF",X"01",
		X"11",X"11",X"11",X"BA",X"FF",X"00",X"00",X"99",X"99",X"40",X"FF",X"00",X"00",X"99",X"99",X"44",
		X"FF",X"00",X"00",X"99",X"94",X"44",X"FF",X"00",X"09",X"99",X"94",X"00",X"FF",X"00",X"09",X"99",
		X"94",X"40",X"FF",X"00",X"00",X"99",X"99",X"40",X"FF",X"AA",X"AA",X"AA",X"AA",X"BB",X"FF",X"01",
		X"11",X"11",X"11",X"BA",X"FF",X"00",X"00",X"99",X"99",X"40",X"FF",X"00",X"00",X"99",X"99",X"44",
		X"FF",X"00",X"00",X"09",X"99",X"94",X"FF",X"00",X"00",X"09",X"99",X"44",X"FF",X"00",X"00",X"99",
		X"99",X"40",X"FF",X"00",X"00",X"09",X"99",X"44",X"FF",X"6F",X"FF",X"FF",X"00",X"04",X"32",X"22",
		X"26",X"FF",X"FF",X"00",X"03",X"22",X"22",X"00",X"00",X"99",X"00",X"00",X"FF",X"00",X"00",X"11",
		X"00",X"00",X"FF",X"00",X"00",X"CC",X"00",X"00",X"FF",X"00",X"00",X"11",X"00",X"00",X"FF",X"00",
		X"00",X"CC",X"00",X"00",X"FF",X"91",X"C1",X"00",X"1C",X"19",X"FF",X"91",X"C1",X"00",X"1C",X"19",
		X"FF",X"00",X"00",X"CC",X"00",X"00",X"FF",X"00",X"00",X"11",X"00",X"00",X"FF",X"00",X"00",X"CC",
		X"00",X"00",X"FF",X"00",X"00",X"11",X"00",X"00",X"FF",X"00",X"00",X"99",X"00",X"00",X"FF",X"10",
		X"00",X"FF",X"11",X"00",X"FF",X"01",X"00",X"FF",X"01",X"10",X"FF",X"00",X"10",X"FF",X"01",X"33",
		X"FF",X"00",X"10",X"FF",X"01",X"10",X"FF",X"01",X"00",X"FF",X"11",X"00",X"FF",X"10",X"00",X"FF",
		X"20",X"00",X"FF",X"22",X"00",X"FF",X"02",X"00",X"FF",X"02",X"20",X"FF",X"00",X"20",X"FF",X"02",
		X"11",X"FF",X"00",X"20",X"FF",X"02",X"20",X"FF",X"02",X"00",X"FF",X"22",X"00",X"FF",X"20",X"00",
		X"FF",X"30",X"00",X"FF",X"33",X"00",X"FF",X"03",X"00",X"FF",X"03",X"30",X"FF",X"00",X"30",X"FF",
		X"03",X"22",X"FF",X"00",X"30",X"FF",X"03",X"30",X"FF",X"03",X"00",X"FF",X"33",X"00",X"FF",X"30",
		X"00",X"FF",X"11",X"00",X"00",X"FF",X"00",X"11",X"00",X"FF",X"00",X"01",X"00",X"FF",X"00",X"01",
		X"10",X"FF",X"00",X"00",X"13",X"FF",X"00",X"01",X"10",X"FF",X"00",X"01",X"00",X"FF",X"00",X"11",
		X"00",X"FF",X"11",X"00",X"00",X"FF",X"22",X"00",X"00",X"FF",X"00",X"22",X"00",X"FF",X"00",X"02",
		X"00",X"FF",X"00",X"02",X"20",X"FF",X"00",X"00",X"21",X"FF",X"00",X"02",X"20",X"FF",X"00",X"02",
		X"00",X"FF",X"00",X"22",X"00",X"FF",X"22",X"00",X"00",X"FF",X"33",X"00",X"00",X"FF",X"00",X"33",
		X"00",X"FF",X"00",X"03",X"00",X"FF",X"00",X"03",X"30",X"FF",X"00",X"00",X"32",X"FF",X"00",X"03",
		X"30",X"FF",X"00",X"03",X"00",X"FF",X"00",X"33",X"00",X"FF",X"33",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"01",X"FF",X"00",X"00",X"00",X"01",X"FF",X"00",X"00",X"00",X"11",X"FF",X"00",X"00",X"00",
		X"10",X"FF",X"00",X"00",X"01",X"10",X"FF",X"00",X"01",X"13",X"00",X"FF",X"11",X"10",X"03",X"00",
		X"FF",X"00",X"00",X"00",X"02",X"FF",X"00",X"00",X"00",X"02",X"FF",X"00",X"00",X"00",X"22",X"FF",
		X"00",X"00",X"00",X"20",X"FF",X"00",X"00",X"02",X"20",X"FF",X"00",X"02",X"21",X"00",X"FF",X"22",
		X"20",X"01",X"00",X"FF",X"00",X"00",X"00",X"03",X"FF",X"00",X"00",X"00",X"03",X"FF",X"00",X"00",
		X"00",X"33",X"FF",X"00",X"00",X"00",X"30",X"FF",X"00",X"00",X"03",X"30",X"FF",X"00",X"03",X"32",
		X"00",X"FF",X"33",X"30",X"02",X"00",X"FF",X"00",X"00",X"01",X"FF",X"00",X"00",X"01",X"FF",X"00",
		X"00",X"11",X"FF",X"00",X"00",X"10",X"FF",X"00",X"00",X"10",X"FF",X"00",X"11",X"30",X"FF",X"11",
		X"10",X"30",X"FF",X"00",X"00",X"02",X"FF",X"00",X"00",X"02",X"FF",X"00",X"00",X"22",X"FF",X"00",
		X"00",X"20",X"FF",X"00",X"00",X"20",X"FF",X"00",X"22",X"10",X"FF",X"22",X"20",X"10",X"FF",X"00",
		X"00",X"03",X"FF",X"00",X"00",X"03",X"FF",X"00",X"00",X"33",X"FF",X"00",X"00",X"30",X"FF",X"00",
		X"00",X"30",X"FF",X"00",X"33",X"20",X"FF",X"33",X"30",X"20",X"FF",X"00",X"00",X"12",X"FF",X"05",
		X"50",X"FF",X"54",X"45",X"FF",X"43",X"34",X"FF",X"43",X"34",X"FF",X"54",X"45",X"FF",X"05",X"50",
		X"FF",X"00",X"07",X"70",X"00",X"FF",X"00",X"75",X"57",X"00",X"FF",X"07",X"54",X"45",X"70",X"FF",
		X"B7",X"43",X"34",X"70",X"FF",X"B7",X"43",X"34",X"70",X"FF",X"B7",X"54",X"45",X"70",X"FF",X"BB",
		X"75",X"57",X"00",X"FF",X"0B",X"B7",X"70",X"00",X"FF",X"00",X"BB",X"00",X"00",X"FF",X"00",X"06",
		X"60",X"00",X"FF",X"00",X"64",X"46",X"00",X"FF",X"06",X"43",X"34",X"60",X"FF",X"B6",X"31",X"13",
		X"60",X"FF",X"B6",X"31",X"13",X"60",X"FF",X"B6",X"43",X"34",X"60",X"FF",X"BB",X"64",X"46",X"00",
		X"FF",X"0B",X"B6",X"60",X"00",X"FF",X"00",X"BB",X"00",X"00",X"FF",X"00",X"05",X"50",X"00",X"FF",
		X"00",X"75",X"44",X"00",X"FF",X"07",X"74",X"34",X"40",X"FF",X"C7",X"54",X"23",X"40",X"FF",X"C9",
		X"55",X"35",X"50",X"FF",X"C9",X"95",X"55",X"60",X"FF",X"CC",X"99",X"56",X"00",X"FF",X"0C",X"C9",
		X"60",X"00",X"FF",X"00",X"CC",X"00",X"00",X"FF",X"00",X"73",X"00",X"00",X"FF",X"0D",X"77",X"00",
		X"73",X"FF",X"0D",X"D0",X"0D",X"77",X"FF",X"00",X"0A",X"6D",X"D0",X"FF",X"00",X"AA",X"66",X"00",
		X"FF",X"0A",X"A9",X"56",X"60",X"FF",X"DA",X"99",X"55",X"60",X"FF",X"DA",X"AA",X"77",X"80",X"FF",
		X"DA",X"AA",X"78",X"80",X"FF",X"DD",X"AA",X"88",X"00",X"FF",X"0D",X"DA",X"80",X"00",X"FF",X"00",
		X"DD",X"00",X"00",X"FF",X"00",X"00",X"00",X"09",X"30",X"FF",X"00",X"09",X"50",X"E9",X"90",X"FF",
		X"00",X"99",X"55",X"EE",X"00",X"FF",X"09",X"9E",X"E5",X"50",X"00",X"FF",X"E9",X"99",X"55",X"50",
		X"93",X"FF",X"EB",X"BB",X"77",X"7E",X"99",X"FF",X"EB",X"BE",X"E7",X"7E",X"E0",X"FF",X"EE",X"BB",
		X"77",X"00",X"00",X"FF",X"0E",X"EB",X"70",X"09",X"30",X"FF",X"00",X"EE",X"00",X"E9",X"90",X"FF",
		X"00",X"09",X"30",X"EE",X"00",X"FF",X"00",X"E9",X"90",X"00",X"00",X"FF",X"00",X"EE",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"95",X"00",X"0B",X"40",X"FF",X"00",X"00",X"0E",X"95",X"50",X"EB",
		X"B0",X"FF",X"0B",X"40",X"99",X"EE",X"E5",X"EE",X"00",X"FF",X"EB",X"BE",X"99",X"95",X"55",X"00",
		X"00",X"FF",X"EE",X"0E",X"BB",X"B7",X"77",X"0B",X"40",X"FF",X"00",X"0E",X"BB",X"EE",X"E7",X"EB",
		X"B0",X"FF",X"0B",X"4E",X"EE",X"B7",X"70",X"EE",X"00",X"FF",X"EB",X"B0",X"EE",X"B7",X"00",X"00",
		X"00",X"FF",X"EE",X"00",X"0E",X"E0",X"0B",X"40",X"00",X"FF",X"00",X"00",X"0B",X"40",X"EB",X"B0",
		X"00",X"FF",X"00",X"00",X"EB",X"B0",X"EE",X"00",X"00",X"FF",X"00",X"00",X"EE",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"B4",X"00",X"B4",X"00",X"00",X"FF",X"00",X"0E",X"BB",X"0E",X"BB",X"00",
		X"00",X"FF",X"00",X"0E",X"E0",X"0E",X"E0",X"00",X"00",X"FF",X"00",X"00",X"00",X"95",X"00",X"00",
		X"00",X"FF",X"0B",X"40",X"0E",X"95",X"E0",X"0B",X"20",X"FF",X"EB",X"B0",X"99",X"EE",X"E5",X"EB",
		X"B0",X"FF",X"EE",X"0E",X"99",X"9E",X"44",X"EE",X"00",X"FF",X"00",X"0E",X"BB",X"BE",X"77",X"00",
		X"00",X"FF",X"0B",X"4E",X"BB",X"EE",X"E7",X"0B",X"40",X"FF",X"EB",X"BE",X"EE",X"B7",X"E0",X"EB",
		X"B0",X"FF",X"EE",X"00",X"EE",X"B7",X"00",X"EE",X"00",X"FF",X"00",X"00",X"0E",X"E0",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"B4",X"00",X"B4",X"00",X"00",X"FF",X"00",X"0E",X"BB",X"0E",X"BB",X"00",
		X"00",X"FF",X"00",X"0E",X"E0",X"0E",X"E0",X"00",X"00",X"FF",X"00",X"00",X"0B",X"40",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"EB",X"B0",X"0B",X"40",X"00",X"FF",X"00",X"00",X"EE",X"00",X"EB",X"B0",
		X"00",X"FF",X"00",X"B4",X"00",X"95",X"EE",X"00",X"00",X"FF",X"0E",X"BB",X"0E",X"95",X"E0",X"00",
		X"00",X"FF",X"0E",X"E0",X"99",X"EE",X"E5",X"0B",X"40",X"FF",X"00",X"0E",X"99",X"9E",X"44",X"EB",
		X"B0",X"FF",X"0B",X"4E",X"BB",X"BE",X"77",X"EE",X"00",X"FF",X"EB",X"BE",X"BB",X"EE",X"E7",X"00",
		X"00",X"FF",X"EE",X"0E",X"EE",X"BB",X"E0",X"B4",X"00",X"FF",X"00",X"00",X"EE",X"BB",X"0E",X"BB",
		X"00",X"FF",X"00",X"0B",X"4E",X"E0",X"0E",X"E0",X"00",X"FF",X"00",X"EB",X"B0",X"0B",X"40",X"00",
		X"00",X"FF",X"00",X"EE",X"00",X"EB",X"B0",X"00",X"00",X"FF",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"B1",X"00",X"00",X"00",X"FF",X"00",X"00",X"0E",X"BB",X"00",X"00",
		X"00",X"FF",X"00",X"B4",X"0E",X"E0",X"00",X"B4",X"00",X"FF",X"0E",X"BB",X"00",X"95",X"0E",X"BB",
		X"00",X"FF",X"0E",X"E0",X"0E",X"95",X"EE",X"E0",X"00",X"FF",X"00",X"00",X"99",X"EE",X"E5",X"00",
		X"00",X"FF",X"0B",X"4E",X"99",X"9E",X"55",X"0B",X"40",X"FF",X"EB",X"BE",X"BB",X"BE",X"77",X"EB",
		X"B0",X"FF",X"EE",X"EE",X"BB",X"EE",X"E7",X"EE",X"00",X"FF",X"00",X"0E",X"EE",X"B7",X"E0",X"00",
		X"00",X"FF",X"00",X"B4",X"EE",X"B7",X"00",X"B4",X"00",X"FF",X"0E",X"BB",X"0E",X"E0",X"0E",X"BB",
		X"00",X"FF",X"0E",X"E0",X"00",X"B4",X"0E",X"E0",X"00",X"FF",X"00",X"00",X"0E",X"BB",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"0E",X"E0",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0B",X"40",X"00",
		X"00",X"FF",X"00",X"0B",X"40",X"EB",X"B0",X"00",X"00",X"FF",X"00",X"EB",X"B0",X"EE",X"00",X"00",
		X"00",X"FF",X"00",X"EE",X"00",X"95",X"00",X"0B",X"10",X"FF",X"00",X"00",X"0E",X"95",X"E0",X"EB",
		X"B0",X"FF",X"0B",X"40",X"99",X"EE",X"E5",X"EE",X"00",X"FF",X"EB",X"BE",X"99",X"9E",X"55",X"00",
		X"00",X"FF",X"EE",X"0E",X"BB",X"BE",X"77",X"0B",X"40",X"FF",X"00",X"0E",X"BB",X"EE",X"E7",X"EB",
		X"B0",X"FF",X"0B",X"4E",X"EE",X"B7",X"E0",X"EE",X"00",X"FF",X"EB",X"B0",X"EE",X"B7",X"00",X"00",
		X"00",X"FF",X"EE",X"00",X"0E",X"E0",X"0B",X"40",X"00",X"FF",X"00",X"00",X"0B",X"40",X"EB",X"B0",
		X"00",X"FF",X"00",X"00",X"EB",X"B0",X"EE",X"00",X"00",X"FF",X"00",X"00",X"EE",X"00",X"00",X"00",
		X"00",X"FF",X"16",X"FF",X"BA",X"FF",X"B1",X"FF",X"85",X"FF",X"8B",X"FF",X"51",X"FF",X"58",X"FF",
		X"1B",X"FF",X"11",X"50",X"FF",X"11",X"55",X"FF",X"BB",X"88",X"FF",X"0B",X"80",X"FF",X"0B",X"11",
		X"FF",X"BB",X"11",X"FF",X"88",X"55",X"FF",X"08",X"50",X"FF",X"08",X"B0",X"FF",X"88",X"BB",X"FF",
		X"55",X"11",X"FF",X"05",X"11",X"FF",X"05",X"80",X"FF",X"55",X"88",X"FF",X"11",X"BB",X"FF",X"11",
		X"B0",X"FF",X"07",X"70",X"FF",X"72",X"27",X"FF",X"72",X"27",X"FF",X"07",X"70",X"FF",X"02",X"20",
		X"FF",X"20",X"02",X"FF",X"20",X"02",X"FF",X"20",X"02",X"FF",X"02",X"20",X"FF",X"00",X"44",X"42",
		X"FF",X"04",X"00",X"04",X"FF",X"40",X"00",X"04",X"FF",X"40",X"00",X"40",X"FF",X"44",X"44",X"00",
		X"FF",X"00",X"00",X"55",X"40",X"FF",X"00",X"07",X"00",X"30",X"FF",X"00",X"70",X"05",X"50",X"FF",
		X"07",X"00",X"55",X"00",X"FF",X"70",X"07",X"50",X"00",X"FF",X"70",X"77",X"00",X"00",X"FF",X"77",
		X"70",X"00",X"00",X"FF",X"00",X"00",X"04",X"70",X"FF",X"00",X"00",X"21",X"40",X"FF",X"00",X"04",
		X"22",X"00",X"FF",X"00",X"64",X"40",X"00",X"FF",X"07",X"66",X"00",X"00",X"FF",X"77",X"70",X"00",
		X"00",X"FF",X"77",X"00",X"00",X"00",X"FF",X"00",X"07",X"77",X"FF",X"00",X"77",X"07",X"FF",X"07",
		X"77",X"07",X"FF",X"06",X"60",X"07",X"FF",X"44",X"50",X"77",X"FF",X"12",X"00",X"77",X"FF",X"25",
		X"07",X"70",X"FF",X"45",X"07",X"70",X"FF",X"65",X"77",X"00",X"FF",X"77",X"70",X"00",X"FF",X"00",
		X"77",X"77",X"00",X"FF",X"06",X"77",X"77",X"70",X"FF",X"56",X"55",X"07",X"77",X"FF",X"55",X"50",
		X"00",X"77",X"FF",X"44",X"40",X"00",X"77",X"FF",X"33",X"30",X"00",X"77",X"FF",X"44",X"40",X"00",
		X"77",X"FF",X"05",X"55",X"07",X"77",X"FF",X"06",X"77",X"77",X"70",X"FF",X"00",X"77",X"77",X"00",
		X"FF",X"00",X"07",X"77",X"70",X"00",X"FF",X"00",X"77",X"77",X"77",X"00",X"FF",X"07",X"77",X"77",
		X"77",X"70",X"FF",X"77",X"77",X"00",X"77",X"77",X"FF",X"77",X"70",X"00",X"07",X"77",X"FF",X"77",
		X"70",X"00",X"07",X"77",X"FF",X"77",X"70",X"00",X"07",X"77",X"FF",X"77",X"70",X"00",X"07",X"77",
		X"FF",X"77",X"65",X"00",X"77",X"77",X"FF",X"07",X"66",X"34",X"57",X"70",X"FF",X"00",X"55",X"34",
		X"66",X"00",X"FF",X"00",X"05",X"34",X"50",X"00",X"FF",X"07",X"77",X"77",X"00",X"00",X"FF",X"00",
		X"03",X"40",X"04",X"40",X"00",X"FF",X"00",X"00",X"04",X"40",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"03",X"33",X"33",X"33",X"33",X"33",X"33",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"07",X"23",X"33",X"33",X"33",X"33",X"33",X"33",X"30",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"02",X"77",X"22",X"33",X"33",X"33",X"33",X"33",X"33",X"63",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"22",X"77",X"72",X"33",X"33",X"33",X"33",X"33",X"33",
		X"63",X"30",X"00",X"00",X"00",X"FF",X"00",X"00",X"02",X"22",X"77",X"72",X"23",X"33",X"33",X"33",
		X"33",X"36",X"63",X"33",X"00",X"00",X"00",X"FF",X"00",X"00",X"72",X"22",X"27",X"77",X"23",X"33",
		X"33",X"33",X"33",X"36",X"33",X"36",X"00",X"00",X"00",X"FF",X"00",X"07",X"77",X"22",X"27",X"77",
		X"22",X"33",X"33",X"33",X"33",X"66",X"33",X"36",X"60",X"00",X"00",X"FF",X"00",X"07",X"77",X"72",
		X"22",X"77",X"72",X"33",X"33",X"33",X"33",X"63",X"33",X"66",X"60",X"00",X"00",X"FF",X"00",X"CC",
		X"BB",X"BB",X"22",X"77",X"72",X"23",X"33",X"33",X"36",X"63",X"33",X"66",X"66",X"00",X"00",X"FF",
		X"00",X"CC",X"BB",X"BB",X"22",X"27",X"77",X"23",X"33",X"33",X"36",X"33",X"36",X"66",X"62",X"20",
		X"00",X"FF",X"0C",X"CC",X"CB",X"BB",X"72",X"27",X"77",X"75",X"55",X"55",X"56",X"33",X"36",X"66",
		X"22",X"70",X"00",X"FF",X"0C",X"CC",X"CB",X"BB",X"72",X"22",X"77",X"55",X"55",X"55",X"55",X"33",
		X"66",X"62",X"22",X"77",X"00",X"FF",X"CC",X"CC",X"CC",X"BB",X"77",X"22",X"75",X"55",X"55",X"55",
		X"55",X"53",X"66",X"22",X"27",X"73",X"00",X"FF",X"DC",X"CC",X"CC",X"BB",X"77",X"22",X"55",X"55",
		X"55",X"55",X"55",X"56",X"62",X"22",X"27",X"73",X"30",X"FF",X"DC",X"CC",X"CC",X"CB",X"77",X"72",
		X"55",X"55",X"55",X"55",X"55",X"56",X"22",X"22",X"77",X"33",X"30",X"FF",X"DD",X"CC",X"CC",X"CB",
		X"77",X"76",X"55",X"55",X"55",X"55",X"55",X"54",X"22",X"22",X"77",X"33",X"30",X"FF",X"DD",X"CC",
		X"CC",X"CB",X"77",X"76",X"55",X"55",X"55",X"55",X"55",X"54",X"22",X"27",X"77",X"33",X"30",X"FF",
		X"DD",X"DC",X"CC",X"CB",X"77",X"72",X"55",X"55",X"55",X"55",X"55",X"56",X"22",X"27",X"73",X"33",
		X"30",X"FF",X"DD",X"DC",X"CC",X"CC",X"77",X"72",X"55",X"55",X"55",X"55",X"55",X"56",X"22",X"77",
		X"73",X"33",X"30",X"FF",X"DD",X"DD",X"CC",X"CC",X"77",X"72",X"55",X"55",X"55",X"55",X"55",X"56",
		X"22",X"77",X"33",X"33",X"30",X"FF",X"DD",X"DD",X"CC",X"CC",X"77",X"72",X"55",X"55",X"55",X"55",
		X"55",X"56",X"22",X"77",X"33",X"33",X"30",X"FF",X"DD",X"DD",X"DC",X"CC",X"77",X"72",X"55",X"55",
		X"55",X"55",X"55",X"56",X"22",X"73",X"33",X"33",X"30",X"FF",X"DD",X"DD",X"DC",X"CC",X"77",X"72",
		X"55",X"55",X"55",X"55",X"55",X"56",X"22",X"73",X"33",X"33",X"30",X"FF",X"DD",X"DD",X"DD",X"CC",
		X"77",X"72",X"55",X"55",X"55",X"55",X"55",X"54",X"22",X"73",X"33",X"33",X"30",X"FF",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"10",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"20",X"33",X"33",
		X"33",X"33",X"33",X"33",X"33",X"30",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"40",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"50",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"60",X"77",X"77",
		X"77",X"77",X"77",X"77",X"77",X"70",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"80",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"90",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
