library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_1M is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_1M is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"CD",X"E4",X"42",X"06",X"00",X"3A",X"77",X"80",X"B7",X"CA",X"28",X"40",X"04",X"3A",X"74",X"80",
		X"B7",X"C2",X"28",X"40",X"04",X"3A",X"80",X"80",X"B7",X"C2",X"28",X"40",X"04",X"3A",X"9B",X"81",
		X"3D",X"32",X"9B",X"81",X"F2",X"28",X"40",X"04",X"78",X"21",X"2F",X"40",X"C3",X"EA",X"00",X"5C",
		X"40",X"AD",X"40",X"87",X"41",X"BA",X"41",X"75",X"42",X"E6",X"42",X"E6",X"42",X"CD",X"55",X"44",
		X"3E",X"00",X"32",X"4E",X"82",X"3E",X"00",X"32",X"4F",X"82",X"3E",X"00",X"32",X"49",X"82",X"3E",
		X"00",X"32",X"77",X"82",X"3E",X"01",X"32",X"03",X"80",X"C3",X"C0",X"00",X"CD",X"E8",X"42",X"CD",
		X"3D",X"43",X"3E",X"00",X"32",X"4B",X"82",X"3A",X"17",X"80",X"B7",X"CA",X"8C",X"40",X"3E",X"A0",
		X"CD",X"FC",X"00",X"AF",X"CD",X"D9",X"4B",X"CD",X"67",X"4B",X"3E",X"01",X"32",X"70",X"80",X"CD",
		X"FD",X"43",X"3E",X"00",X"32",X"70",X"80",X"CD",X"69",X"43",X"18",X"03",X"CD",X"CF",X"45",X"CD",
		X"95",X"44",X"CD",X"55",X"44",X"3E",X"00",X"32",X"81",X"80",X"3E",X"01",X"32",X"70",X"80",X"01",
		X"1E",X"00",X"CD",X"E1",X"00",X"3E",X"01",X"32",X"03",X"80",X"C3",X"C0",X"00",X"3E",X"00",X"32",
		X"28",X"80",X"32",X"77",X"80",X"32",X"74",X"80",X"32",X"88",X"80",X"00",X"CD",X"F8",X"5F",X"CD",
		X"30",X"60",X"3E",X"01",X"CD",X"FC",X"00",X"3E",X"25",X"CD",X"FC",X"00",X"3E",X"01",X"32",X"8D",
		X"80",X"01",X"F0",X"00",X"3E",X"01",X"32",X"6E",X"80",X"3A",X"6E",X"80",X"B7",X"C2",X"D9",X"40",
		X"C5",X"CD",X"33",X"60",X"CD",X"00",X"20",X"CD",X"10",X"30",X"C1",X"0B",X"78",X"B1",X"20",X"E4",
		X"21",X"48",X"0D",X"22",X"51",X"88",X"3E",X"00",X"32",X"8D",X"80",X"CD",X"20",X"4E",X"3E",X"00",
		X"32",X"AC",X"81",X"CD",X"67",X"4B",X"AF",X"CD",X"D9",X"4B",X"CD",X"F5",X"5F",X"CD",X"E0",X"2F",
		X"CD",X"E6",X"2F",X"CD",X"20",X"4E",X"21",X"A2",X"81",X"01",X"05",X"00",X"CD",X"CC",X"00",X"3E",
		X"00",X"32",X"AB",X"81",X"32",X"AC",X"81",X"32",X"B0",X"81",X"3A",X"A0",X"81",X"3C",X"32",X"A0",
		X"81",X"3A",X"A0",X"81",X"FE",X"41",X"DA",X"3E",X"41",X"3E",X"20",X"32",X"A0",X"81",X"3A",X"AF",
		X"81",X"FE",X"99",X"28",X"05",X"C6",X"01",X"27",X"18",X"02",X"3E",X"00",X"32",X"AF",X"81",X"3A",
		X"27",X"80",X"CD",X"40",X"44",X"3E",X"01",X"32",X"48",X"82",X"CD",X"CE",X"4E",X"CD",X"F4",X"4B",
		X"3E",X"18",X"32",X"A2",X"81",X"CD",X"0C",X"60",X"CD",X"E9",X"5F",X"CD",X"E8",X"42",X"CD",X"3D",
		X"43",X"CD",X"1F",X"44",X"C3",X"A0",X"4F",X"CD",X"E0",X"5F",X"3E",X"00",X"32",X"53",X"84",X"3E",
		X"01",X"32",X"54",X"84",X"C3",X"3D",X"40",X"3E",X"00",X"32",X"77",X"80",X"3E",X"00",X"32",X"80",
		X"80",X"3E",X"00",X"32",X"88",X"80",X"3E",X"00",X"32",X"8E",X"80",X"CD",X"20",X"4E",X"AF",X"CD",
		X"D9",X"4B",X"CD",X"F0",X"00",X"DD",X"21",X"4A",X"D2",X"CD",X"D2",X"00",X"3E",X"0D",X"CD",X"18",
		X"60",X"CD",X"FB",X"5F",X"CD",X"F8",X"5F",X"C3",X"F0",X"40",X"3E",X"00",X"32",X"77",X"80",X"3E",
		X"00",X"32",X"88",X"80",X"3E",X"00",X"32",X"95",X"80",X"3A",X"28",X"80",X"CB",X"97",X"32",X"28",
		X"80",X"3E",X"01",X"32",X"8D",X"80",X"06",X"7E",X"3E",X"01",X"32",X"6E",X"80",X"3A",X"6E",X"80",
		X"B7",X"C2",X"DD",X"41",X"C5",X"CD",X"00",X"20",X"CD",X"10",X"30",X"C1",X"78",X"FE",X"78",X"C2",
		X"F7",X"41",X"3E",X"01",X"CD",X"FC",X"00",X"10",X"DF",X"21",X"48",X"0D",X"22",X"51",X"88",X"3E",
		X"00",X"32",X"8D",X"80",X"3E",X"00",X"CD",X"D9",X"4B",X"CD",X"67",X"4B",X"3E",X"00",X"32",X"B0",
		X"81",X"CD",X"20",X"4E",X"CD",X"EF",X"5F",X"3A",X"27",X"80",X"CD",X"40",X"44",X"CD",X"87",X"45",
		X"3A",X"27",X"80",X"CD",X"2B",X"44",X"3A",X"AC",X"81",X"FE",X"00",X"28",X"05",X"CD",X"E3",X"2F",
		X"18",X"03",X"CD",X"E0",X"2F",X"CD",X"E6",X"2F",X"CD",X"0C",X"60",X"CD",X"EC",X"5F",X"3E",X"00",
		X"32",X"48",X"82",X"CD",X"CE",X"4E",X"CD",X"20",X"4E",X"CD",X"F4",X"4B",X"CD",X"E6",X"2F",X"CD",
		X"E9",X"5F",X"CD",X"E8",X"42",X"CD",X"1F",X"44",X"CD",X"C9",X"47",X"3A",X"9B",X"81",X"3C",X"32",
		X"9B",X"81",X"CD",X"3D",X"43",X"CD",X"E0",X"5F",X"3A",X"9B",X"81",X"3D",X"32",X"9B",X"81",X"CD",
		X"3D",X"43",X"C3",X"3D",X"40",X"3E",X"00",X"32",X"77",X"80",X"3E",X"00",X"32",X"88",X"80",X"3E",
		X"00",X"32",X"8D",X"80",X"3E",X"00",X"32",X"4B",X"82",X"3E",X"01",X"CD",X"FC",X"00",X"3E",X"26",
		X"CD",X"FC",X"00",X"3E",X"01",X"CD",X"D9",X"4B",X"3A",X"27",X"80",X"CD",X"40",X"44",X"CD",X"E3",
		X"5F",X"CD",X"20",X"4E",X"CD",X"67",X"4B",X"CD",X"00",X"48",X"3E",X"01",X"CD",X"FC",X"00",X"CD",
		X"20",X"4E",X"3A",X"8B",X"80",X"B7",X"C2",X"D3",X"42",X"3A",X"26",X"80",X"B7",X"CA",X"D3",X"42",
		X"3A",X"27",X"80",X"B7",X"C2",X"CC",X"42",X"3A",X"CD",X"81",X"18",X"03",X"3A",X"B4",X"81",X"B7",
		X"F2",X"11",X"42",X"CD",X"39",X"4B",X"3E",X"00",X"32",X"70",X"80",X"3E",X"01",X"32",X"03",X"80",
		X"C3",X"C6",X"00",X"C9",X"00",X"C9",X"00",X"C9",X"3A",X"70",X"80",X"B7",X"CA",X"14",X"43",X"3A",
		X"27",X"80",X"B7",X"CA",X"FE",X"42",X"CD",X"CF",X"00",X"91",X"CA",X"03",X"18",X"2A",X"3A",X"26",
		X"80",X"B7",X"20",X"08",X"CD",X"CF",X"00",X"89",X"CA",X"04",X"18",X"1C",X"CD",X"CF",X"00",X"83",
		X"CA",X"03",X"18",X"14",X"3A",X"26",X"80",X"B7",X"20",X"08",X"CD",X"CF",X"00",X"6D",X"CA",X"04",
		X"18",X"06",X"CD",X"CF",X"00",X"67",X"CA",X"03",X"3A",X"26",X"80",X"B7",X"20",X"08",X"CD",X"D8",
		X"00",X"7B",X"CA",X"02",X"18",X"06",X"CD",X"D8",X"00",X"75",X"CA",X"03",X"C9",X"CD",X"AC",X"44",
		X"DD",X"21",X"A7",X"CA",X"CD",X"D2",X"00",X"DD",X"21",X"C1",X"CA",X"CD",X"D5",X"00",X"DD",X"21",
		X"C7",X"CA",X"3A",X"AF",X"81",X"FE",X"10",X"DA",X"5E",X"43",X"DD",X"21",X"CF",X"CA",X"CD",X"D2",
		X"00",X"DD",X"21",X"D5",X"CA",X"CD",X"D2",X"00",X"C9",X"CD",X"E8",X"42",X"CD",X"3D",X"43",X"CD",
		X"E0",X"2F",X"CD",X"20",X"4E",X"3A",X"17",X"80",X"B7",X"CA",X"C8",X"43",X"3A",X"8B",X"80",X"B7",
		X"C2",X"8B",X"43",X"CD",X"DF",X"4C",X"3E",X"01",X"32",X"81",X"80",X"CD",X"0B",X"45",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"01",X"32",X"70",X"80",
		X"CD",X"20",X"4E",X"CD",X"2A",X"60",X"21",X"B4",X"81",X"01",X"32",X"00",X"CD",X"CC",X"00",X"CD",
		X"CC",X"43",X"AF",X"CD",X"40",X"44",X"3E",X"01",X"CD",X"40",X"44",X"3E",X"00",X"32",X"E5",X"81",
		X"3A",X"CD",X"81",X"32",X"75",X"80",X"18",X"03",X"CD",X"CC",X"43",X"C9",X"CD",X"20",X"4E",X"3E",
		X"00",X"32",X"48",X"82",X"CD",X"CE",X"4E",X"CD",X"F4",X"4B",X"CD",X"0C",X"60",X"CD",X"E9",X"5F",
		X"CD",X"C9",X"47",X"3A",X"17",X"80",X"B7",X"28",X"00",X"CD",X"E8",X"42",X"3A",X"9B",X"81",X"3D",
		X"32",X"9B",X"81",X"CD",X"1F",X"44",X"CD",X"E0",X"5F",X"CD",X"3D",X"43",X"C9",X"21",X"9B",X"81",
		X"01",X"19",X"00",X"CD",X"CC",X"00",X"3A",X"71",X"80",X"32",X"9B",X"81",X"3E",X"01",X"32",X"A0",
		X"81",X"3E",X"18",X"32",X"A2",X"81",X"3E",X"01",X"32",X"AF",X"81",X"CD",X"15",X"60",X"C9",X"CD",
		X"E7",X"00",X"CD",X"27",X"4E",X"3E",X"01",X"32",X"8C",X"80",X"C9",X"B7",X"C2",X"34",X"44",X"21",
		X"B4",X"81",X"18",X"03",X"21",X"CD",X"81",X"11",X"9B",X"81",X"01",X"19",X"00",X"ED",X"B0",X"C9",
		X"B7",X"C2",X"49",X"44",X"11",X"B4",X"81",X"18",X"03",X"11",X"CD",X"81",X"21",X"9B",X"81",X"01",
		X"19",X"00",X"ED",X"B0",X"C9",X"DD",X"21",X"28",X"80",X"DD",X"36",X"00",X"00",X"DD",X"36",X"01",
		X"18",X"DD",X"36",X"02",X"00",X"DD",X"36",X"03",X"78",X"DD",X"36",X"04",X"78",X"DD",X"36",X"05",
		X"00",X"DD",X"36",X"06",X"00",X"DD",X"36",X"09",X"80",X"DD",X"36",X"0B",X"FF",X"DD",X"36",X"0E",
		X"00",X"DD",X"36",X"0E",X"00",X"DD",X"36",X"12",X"FF",X"21",X"29",X"80",X"01",X"04",X"00",X"11",
		X"00",X"85",X"ED",X"B0",X"C9",X"3E",X"00",X"32",X"53",X"84",X"3E",X"01",X"32",X"54",X"84",X"21",
		X"E0",X"00",X"22",X"5B",X"84",X"21",X"E0",X"FE",X"22",X"5D",X"84",X"C9",X"3A",X"9B",X"81",X"B7",
		X"CA",X"D3",X"44",X"FE",X"01",X"CA",X"DA",X"44",X"FE",X"02",X"CA",X"E1",X"44",X"FE",X"03",X"CA",
		X"E8",X"44",X"FE",X"04",X"CA",X"EF",X"44",X"FE",X"05",X"CA",X"F6",X"44",X"FE",X"06",X"CA",X"FD",
		X"44",X"18",X"31",X"CD",X"CF",X"00",X"DB",X"CA",X"02",X"C9",X"CD",X"CF",X"00",X"DF",X"CA",X"02",
		X"C9",X"CD",X"CF",X"00",X"E3",X"CA",X"02",X"C9",X"CD",X"CF",X"00",X"E7",X"CA",X"02",X"C9",X"CD",
		X"CF",X"00",X"EB",X"CA",X"02",X"C9",X"CD",X"CF",X"00",X"EF",X"CA",X"02",X"C9",X"CD",X"CF",X"00",
		X"F3",X"CA",X"02",X"C9",X"CD",X"CF",X"00",X"F7",X"CA",X"02",X"C9",X"3E",X"02",X"32",X"8C",X"80",
		X"3A",X"8B",X"80",X"F5",X"3E",X"00",X"32",X"8B",X"80",X"F1",X"FE",X"02",X"CA",X"3E",X"45",X"FE",
		X"01",X"CA",X"68",X"45",X"3A",X"02",X"B0",X"E6",X"08",X"C2",X"36",X"45",X"3A",X"02",X"B0",X"E6",
		X"04",X"C2",X"68",X"45",X"18",X"D5",X"3A",X"17",X"80",X"FE",X"02",X"DA",X"0B",X"45",X"3E",X"01",
		X"32",X"26",X"80",X"3A",X"87",X"80",X"B7",X"CA",X"5D",X"45",X"3A",X"87",X"80",X"3D",X"32",X"87",
		X"80",X"CA",X"7D",X"45",X"3A",X"87",X"80",X"3D",X"32",X"87",X"80",X"18",X"29",X"3A",X"17",X"80",
		X"C6",X"98",X"27",X"32",X"17",X"80",X"18",X"1E",X"3E",X"00",X"32",X"26",X"80",X"3A",X"87",X"80",
		X"B7",X"CA",X"7D",X"45",X"3A",X"87",X"80",X"3D",X"32",X"87",X"80",X"18",X"09",X"3A",X"17",X"80",
		X"C6",X"99",X"27",X"32",X"17",X"80",X"C9",X"3A",X"26",X"80",X"B7",X"CA",X"CE",X"45",X"3A",X"75",
		X"80",X"B7",X"FA",X"CE",X"45",X"3A",X"27",X"80",X"3C",X"E6",X"01",X"32",X"27",X"80",X"3A",X"13",
		X"80",X"E6",X"40",X"C2",X"B9",X"45",X"3A",X"27",X"80",X"B7",X"CA",X"B4",X"45",X"3E",X"01",X"32",
		X"04",X"B0",X"18",X"05",X"3E",X"00",X"32",X"04",X"B0",X"3A",X"27",X"80",X"B7",X"C2",X"C8",X"45",
		X"3A",X"CD",X"81",X"32",X"75",X"80",X"18",X"06",X"3A",X"B4",X"81",X"32",X"75",X"80",X"C9",X"3E",
		X"00",X"32",X"88",X"80",X"3E",X"00",X"32",X"8D",X"80",X"3E",X"01",X"CD",X"FC",X"00",X"CD",X"20",
		X"4E",X"AF",X"CD",X"D9",X"4B",X"CD",X"E4",X"42",X"CD",X"67",X"4B",X"3A",X"AB",X"81",X"F5",X"CD",
		X"FD",X"43",X"F1",X"32",X"AB",X"81",X"CD",X"3D",X"43",X"3A",X"79",X"80",X"21",X"22",X"46",X"CD",
		X"EA",X"00",X"3A",X"79",X"80",X"3C",X"32",X"79",X"80",X"3A",X"79",X"80",X"FE",X"04",X"DA",X"16",
		X"46",X"3E",X"00",X"32",X"79",X"80",X"3E",X"00",X"32",X"78",X"80",X"3E",X"00",X"32",X"4B",X"82",
		X"18",X"AD",X"32",X"46",X"5A",X"46",X"50",X"47",X"C5",X"46",X"E6",X"42",X"E6",X"42",X"E6",X"42",
		X"E6",X"42",X"CD",X"CF",X"00",X"00",X"C0",X"0C",X"00",X"CD",X"D8",X"00",X"96",X"C1",X"0A",X"CD",
		X"CF",X"00",X"E6",X"C1",X"0A",X"CD",X"D8",X"00",X"FA",X"C1",X"0A",X"CD",X"9B",X"47",X"3E",X"0D",
		X"CD",X"18",X"60",X"01",X"2C",X"01",X"CD",X"E1",X"00",X"C9",X"CD",X"FD",X"43",X"CD",X"69",X"43",
		X"CD",X"95",X"44",X"CD",X"55",X"44",X"3E",X"00",X"32",X"7A",X"80",X"3E",X"00",X"32",X"7B",X"80",
		X"3A",X"E8",X"80",X"FE",X"00",X"20",X"05",X"2A",X"F8",X"CD",X"18",X"03",X"2A",X"FA",X"CD",X"22",
		X"7C",X"80",X"22",X"7E",X"80",X"01",X"1E",X"00",X"CD",X"E1",X"00",X"18",X"00",X"21",X"01",X"00",
		X"22",X"6E",X"80",X"CD",X"59",X"47",X"CD",X"00",X"10",X"3A",X"6E",X"80",X"B7",X"28",X"EE",X"CD",
		X"00",X"20",X"3A",X"6E",X"80",X"B7",X"28",X"E5",X"CD",X"00",X"30",X"3A",X"6E",X"80",X"B7",X"28",
		X"DC",X"CD",X"00",X"50",X"3A",X"78",X"80",X"B7",X"C2",X"C4",X"46",X"3A",X"6E",X"80",X"B7",X"CA",
		X"8D",X"46",X"18",X"F7",X"C9",X"3A",X"AB",X"81",X"FE",X"17",X"20",X"11",X"3E",X"3C",X"32",X"B3",
		X"81",X"21",X"E0",X"00",X"22",X"5B",X"84",X"21",X"E0",X"FE",X"22",X"5D",X"84",X"3E",X"00",X"32",
		X"AB",X"81",X"3E",X"02",X"32",X"A0",X"81",X"3E",X"18",X"32",X"A2",X"81",X"3E",X"02",X"32",X"AF",
		X"81",X"3A",X"71",X"80",X"32",X"9B",X"81",X"3A",X"E8",X"80",X"FE",X"00",X"20",X"0A",X"2A",X"FC",
		X"CD",X"3E",X"01",X"32",X"E8",X"80",X"18",X"08",X"2A",X"FE",X"CD",X"3E",X"00",X"32",X"E8",X"80",
		X"22",X"7C",X"80",X"22",X"7E",X"80",X"3E",X"01",X"32",X"48",X"82",X"3E",X"00",X"32",X"A7",X"81",
		X"18",X"00",X"CD",X"E0",X"2F",X"CD",X"CE",X"4E",X"CD",X"F4",X"4B",X"CD",X"0C",X"60",X"CD",X"E9",
		X"5F",X"3E",X"00",X"32",X"7A",X"80",X"3E",X"00",X"32",X"7B",X"80",X"CD",X"3D",X"43",X"CD",X"E8",
		X"42",X"CD",X"1F",X"44",X"CD",X"C9",X"47",X"CD",X"E0",X"5F",X"CD",X"55",X"44",X"C3",X"8D",X"46",
		X"3E",X"0D",X"CD",X"18",X"60",X"CD",X"21",X"60",X"C9",X"DD",X"21",X"7A",X"80",X"DD",X"7E",X"01",
		X"FE",X"00",X"C2",X"97",X"47",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"7E",X"DD",X"77",X"01",X"FE",
		X"FF",X"C2",X"8A",X"47",X"DD",X"36",X"00",X"00",X"DD",X"36",X"01",X"01",X"DD",X"7E",X"04",X"DD",
		X"77",X"02",X"DD",X"7E",X"05",X"DD",X"77",X"03",X"18",X"0C",X"23",X"7E",X"DD",X"77",X"00",X"23",
		X"DD",X"75",X"02",X"DD",X"74",X"03",X"C9",X"DD",X"35",X"01",X"C9",X"21",X"28",X"81",X"DD",X"21",
		X"87",X"94",X"06",X"0A",X"4E",X"DD",X"22",X"E6",X"80",X"7E",X"B9",X"38",X"07",X"28",X"05",X"DD",
		X"22",X"E6",X"80",X"4F",X"23",X"DD",X"23",X"DD",X"23",X"10",X"EE",X"2A",X"E6",X"80",X"36",X"0F",
		X"B7",X"11",X"20",X"00",X"ED",X"52",X"36",X"0F",X"C9",X"3E",X"21",X"CD",X"FC",X"00",X"21",X"3D",
		X"DE",X"01",X"06",X"00",X"3A",X"A0",X"81",X"CD",X"F6",X"00",X"7E",X"C6",X"22",X"CD",X"FC",X"00",
		X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DD",X"21",X"00",X"81",X"06",X"0A",X"0E",X"00",X"FD",X"21",X"9C",X"81",X"FD",X"7E",X"03",X"DD",
		X"96",X"03",X"38",X"22",X"20",X"2D",X"FD",X"7E",X"02",X"DD",X"96",X"02",X"38",X"18",X"20",X"23",
		X"FD",X"7E",X"01",X"DD",X"96",X"01",X"38",X"0E",X"20",X"19",X"FD",X"7E",X"00",X"DD",X"96",X"00",
		X"38",X"04",X"28",X"02",X"18",X"0D",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"0C",X"10",
		X"CB",X"18",X"07",X"79",X"32",X"96",X"81",X"CD",X"4B",X"48",X"C9",X"CD",X"20",X"4E",X"21",X"00",
		X"85",X"01",X"60",X"00",X"CD",X"CC",X"00",X"CD",X"FC",X"48",X"CD",X"7C",X"49",X"CD",X"20",X"4B",
		X"3E",X"A6",X"CD",X"FC",X"00",X"3A",X"96",X"81",X"B7",X"C2",X"79",X"48",X"3E",X"29",X"CD",X"FC",
		X"00",X"3E",X"0D",X"CD",X"18",X"60",X"C3",X"83",X"48",X"3E",X"2A",X"CD",X"FC",X"00",X"3E",X"0D",
		X"CD",X"18",X"60",X"CD",X"9B",X"47",X"2A",X"E6",X"80",X"E5",X"DD",X"E1",X"DD",X"36",X"00",X"02",
		X"DD",X"36",X"E0",X"02",X"DD",X"21",X"87",X"96",X"DD",X"36",X"A0",X"02",X"DD",X"36",X"C0",X"02",
		X"DD",X"36",X"E0",X"02",X"DD",X"36",X"00",X"02",X"DD",X"36",X"20",X"02",X"DD",X"36",X"40",X"02",
		X"DD",X"36",X"60",X"02",X"DD",X"36",X"80",X"02",X"DD",X"21",X"1C",X"96",X"DD",X"36",X"80",X"01",
		X"DD",X"36",X"A0",X"01",X"DD",X"36",X"C0",X"01",X"DD",X"36",X"E0",X"01",X"DD",X"36",X"00",X"01",
		X"DD",X"36",X"20",X"01",X"3A",X"96",X"81",X"DD",X"21",X"07",X"94",X"FE",X"00",X"28",X"07",X"DD",
		X"23",X"DD",X"23",X"3D",X"18",X"F5",X"3E",X"20",X"11",X"20",X"00",X"FE",X"00",X"28",X"09",X"DD",
		X"36",X"00",X"0F",X"DD",X"19",X"3D",X"18",X"F3",X"CD",X"93",X"49",X"C9",X"3A",X"96",X"81",X"21",
		X"31",X"81",X"11",X"30",X"81",X"F5",X"47",X"3E",X"09",X"90",X"47",X"B7",X"28",X"06",X"1A",X"77",
		X"2B",X"1B",X"10",X"FA",X"3A",X"AF",X"81",X"77",X"F1",X"F5",X"47",X"3E",X"09",X"90",X"47",X"B7",
		X"28",X"41",X"21",X"20",X"81",X"11",X"24",X"81",X"0E",X"04",X"7E",X"12",X"23",X"13",X"0D",X"20",
		X"F9",X"C5",X"01",X"F8",X"FF",X"09",X"E5",X"EB",X"09",X"EB",X"E1",X"C1",X"10",X"EA",X"F1",X"F5",
		X"47",X"3E",X"09",X"90",X"47",X"21",X"84",X"81",X"11",X"8E",X"81",X"0E",X"03",X"7E",X"12",X"23",
		X"23",X"13",X"13",X"0D",X"20",X"F7",X"C5",X"01",X"F0",X"FF",X"09",X"E5",X"EB",X"09",X"EB",X"E1",
		X"C1",X"10",X"E8",X"F1",X"47",X"00",X"21",X"FC",X"80",X"11",X"04",X"00",X"04",X"19",X"10",X"FD",
		X"11",X"9C",X"81",X"06",X"04",X"1A",X"77",X"13",X"23",X"10",X"FA",X"C9",X"3A",X"96",X"81",X"3C",
		X"21",X"2A",X"81",X"11",X"0A",X"00",X"19",X"3D",X"20",X"FC",X"06",X"03",X"36",X"00",X"23",X"23",
		X"10",X"FA",X"C9",X"01",X"10",X"0E",X"ED",X"43",X"6E",X"80",X"3E",X"01",X"32",X"97",X"81",X"CD",
		X"41",X"4A",X"CD",X"CD",X"4A",X"CD",X"B4",X"4A",X"36",X"41",X"CD",X"CD",X"4A",X"3A",X"1B",X"80",
		X"CB",X"67",X"C2",X"05",X"4A",X"3A",X"19",X"80",X"CB",X"67",X"C2",X"DE",X"49",X"3A",X"20",X"80",
		X"FE",X"03",X"28",X"69",X"CD",X"83",X"4E",X"B7",X"C2",X"DD",X"49",X"ED",X"4B",X"6E",X"80",X"79",
		X"B0",X"20",X"DA",X"AF",X"CD",X"41",X"4A",X"01",X"B4",X"00",X"CD",X"E1",X"00",X"C9",X"3E",X"00",
		X"32",X"19",X"80",X"CD",X"B4",X"4A",X"7E",X"FE",X"00",X"20",X"04",X"36",X"41",X"18",X"11",X"FE",
		X"5A",X"20",X"04",X"36",X"2E",X"18",X"09",X"FE",X"2E",X"20",X"04",X"36",X"00",X"18",X"01",X"34",
		X"CD",X"CD",X"4A",X"18",X"BF",X"3E",X"00",X"32",X"1B",X"80",X"CD",X"B4",X"4A",X"7E",X"FE",X"00",
		X"20",X"04",X"36",X"2E",X"18",X"11",X"FE",X"41",X"20",X"04",X"36",X"00",X"18",X"09",X"FE",X"2E",
		X"20",X"04",X"36",X"5A",X"18",X"01",X"35",X"CD",X"CD",X"4A",X"C3",X"C4",X"49",X"3C",X"3C",X"32",
		X"20",X"80",X"3A",X"97",X"81",X"3C",X"FE",X"04",X"32",X"97",X"81",X"DA",X"A5",X"49",X"D2",X"D3",
		X"49",X"F5",X"11",X"00",X"00",X"21",X"82",X"4A",X"3A",X"96",X"81",X"87",X"5F",X"19",X"5E",X"23",
		X"56",X"EB",X"F1",X"11",X"96",X"4A",X"B7",X"28",X"03",X"11",X"A5",X"4A",X"06",X"05",X"0E",X"03",
		X"D5",X"E5",X"1A",X"FE",X"FF",X"28",X"01",X"77",X"FE",X"00",X"28",X"06",X"11",X"00",X"04",X"19",
		X"36",X"0F",X"E1",X"D1",X"23",X"13",X"0D",X"20",X"E7",X"D5",X"11",X"1D",X"00",X"19",X"D1",X"10",
		X"DD",X"C9",X"66",X"91",X"68",X"91",X"6A",X"91",X"6C",X"91",X"6E",X"91",X"70",X"91",X"72",X"91",
		X"74",X"91",X"76",X"91",X"78",X"91",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"FF",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"F2",X"F4",X"F7",X"F1",X"00",X"F6",X"F1",X"00",X"F6",X"F1",X"00",
		X"F6",X"F0",X"F3",X"F5",X"3A",X"96",X"81",X"21",X"32",X"81",X"11",X"0A",X"00",X"B7",X"28",X"04",
		X"19",X"3D",X"18",X"F9",X"3A",X"97",X"81",X"87",X"16",X"00",X"5F",X"19",X"C9",X"3A",X"96",X"81",
		X"21",X"32",X"81",X"11",X"0A",X"00",X"B7",X"28",X"05",X"19",X"3D",X"C3",X"D6",X"4A",X"E5",X"DD",
		X"E1",X"DD",X"7E",X"03",X"F5",X"DD",X"7E",X"05",X"F5",X"DD",X"7E",X"07",X"F5",X"DD",X"36",X"03",
		X"06",X"DD",X"36",X"05",X"06",X"DD",X"36",X"07",X"06",X"3A",X"97",X"81",X"FE",X"03",X"28",X"0C",
		X"FE",X"02",X"28",X"04",X"DD",X"36",X"03",X"03",X"DD",X"36",X"05",X"03",X"DD",X"36",X"07",X"03",
		X"CD",X"D2",X"00",X"F1",X"DD",X"77",X"07",X"F1",X"DD",X"77",X"05",X"F1",X"DD",X"77",X"03",X"C9",
		X"CD",X"CF",X"00",X"4A",X"C2",X"0D",X"CD",X"D8",X"00",X"96",X"C1",X"0A",X"CD",X"CF",X"00",X"E6",
		X"C1",X"0A",X"CD",X"D8",X"00",X"FA",X"C1",X"0A",X"C9",X"CD",X"67",X"4B",X"21",X"9B",X"81",X"01",
		X"19",X"00",X"CD",X"CC",X"00",X"21",X"B9",X"81",X"01",X"14",X"00",X"CD",X"CC",X"00",X"21",X"D2",
		X"81",X"01",X"14",X"00",X"CD",X"CC",X"00",X"3E",X"00",X"32",X"79",X"80",X"3E",X"00",X"32",X"04",
		X"B0",X"3E",X"00",X"32",X"27",X"80",X"C9",X"2A",X"5B",X"84",X"E5",X"2A",X"5D",X"84",X"E5",X"21",
		X"28",X"80",X"01",X"46",X"00",X"CD",X"CC",X"00",X"21",X"78",X"82",X"01",X"F4",X"01",X"CD",X"CC",
		X"00",X"21",X"D2",X"80",X"01",X"10",X"00",X"CD",X"CC",X"00",X"21",X"C0",X"80",X"01",X"12",X"00",
		X"CD",X"CC",X"00",X"21",X"00",X"89",X"01",X"14",X"00",X"CD",X"CC",X"00",X"E1",X"22",X"5D",X"84",
		X"E1",X"22",X"5B",X"84",X"C9",X"21",X"00",X"90",X"01",X"00",X"04",X"36",X"00",X"23",X"0B",X"78",
		X"B1",X"C2",X"AB",X"4B",X"21",X"00",X"98",X"01",X"00",X"04",X"36",X"00",X"23",X"0B",X"78",X"B1",
		X"C2",X"BA",X"4B",X"C9",X"F5",X"C5",X"E5",X"21",X"28",X"80",X"01",X"20",X"00",X"36",X"00",X"23",
		X"0B",X"78",X"B1",X"20",X"F8",X"E1",X"C1",X"F1",X"C9",X"C5",X"E5",X"B7",X"CA",X"E7",X"4B",X"21",
		X"08",X"85",X"06",X"58",X"C3",X"EC",X"4B",X"21",X"00",X"85",X"06",X"60",X"36",X"00",X"23",X"10",
		X"FB",X"E1",X"C1",X"C9",X"3E",X"01",X"32",X"8F",X"80",X"3A",X"A0",X"81",X"3D",X"01",X"06",X"00",
		X"21",X"38",X"DE",X"CD",X"F6",X"00",X"7E",X"32",X"A1",X"81",X"21",X"74",X"7C",X"CD",X"EA",X"00",
		X"3E",X"00",X"32",X"8F",X"80",X"21",X"3A",X"DE",X"01",X"06",X"00",X"3A",X"A0",X"81",X"3D",X"CD",
		X"F6",X"00",X"7E",X"E6",X"07",X"CD",X"18",X"60",X"C9",X"C5",X"D5",X"E5",X"57",X"3E",X"01",X"32",
		X"8F",X"80",X"1E",X"66",X"CD",X"D3",X"5F",X"06",X"0D",X"21",X"43",X"90",X"73",X"23",X"73",X"34",
		X"23",X"10",X"F9",X"21",X"A3",X"93",X"06",X"0D",X"73",X"23",X"73",X"34",X"23",X"10",X"F9",X"7A",
		X"21",X"43",X"94",X"06",X"1A",X"4F",X"77",X"23",X"10",X"FC",X"21",X"A3",X"97",X"06",X"1A",X"79",
		X"77",X"23",X"10",X"FC",X"11",X"80",X"87",X"21",X"A3",X"4C",X"01",X"3C",X"00",X"ED",X"B0",X"4F",
		X"CD",X"98",X"4C",X"DD",X"21",X"80",X"87",X"CD",X"D2",X"00",X"3E",X"1D",X"32",X"80",X"87",X"3E",
		X"6A",X"32",X"82",X"87",X"3E",X"6B",X"32",X"B8",X"87",X"79",X"CD",X"98",X"4C",X"DD",X"21",X"80",
		X"87",X"CD",X"D2",X"00",X"E1",X"D1",X"C1",X"C9",X"06",X"1C",X"21",X"83",X"87",X"77",X"23",X"23",
		X"10",X"FB",X"C9",X"02",X"02",X"68",X"01",X"62",X"01",X"63",X"01",X"62",X"01",X"63",X"01",X"62",
		X"01",X"63",X"01",X"62",X"01",X"63",X"01",X"62",X"01",X"63",X"01",X"62",X"01",X"63",X"01",X"62",
		X"01",X"63",X"01",X"62",X"01",X"63",X"01",X"62",X"01",X"63",X"01",X"62",X"01",X"63",X"01",X"62",
		X"01",X"63",X"01",X"62",X"01",X"63",X"01",X"62",X"01",X"63",X"01",X"69",X"01",X"FF",X"FF",X"3E",
		X"0D",X"CD",X"18",X"60",X"CD",X"27",X"60",X"CD",X"24",X"60",X"CD",X"CF",X"00",X"00",X"D0",X"04",
		X"DD",X"21",X"14",X"D0",X"3A",X"17",X"80",X"FE",X"01",X"CA",X"00",X"4D",X"DD",X"21",X"40",X"D0",
		X"CD",X"D2",X"00",X"CD",X"F0",X"00",X"C3",X"63",X"4D",X"E6",X"07",X"21",X"11",X"4D",X"C3",X"EA",
		X"00",X"21",X"4D",X"24",X"4D",X"2D",X"4D",X"36",X"4D",X"3F",X"4D",X"48",X"4D",X"51",X"4D",X"5A",
		X"4D",X"C3",X"68",X"4D",X"CD",X"CF",X"00",X"AA",X"D0",X"02",X"C3",X"68",X"4D",X"CD",X"CF",X"00",
		X"AE",X"D0",X"02",X"C3",X"68",X"4D",X"CD",X"CF",X"00",X"B2",X"D0",X"02",X"C3",X"68",X"4D",X"CD",
		X"CF",X"00",X"B6",X"D0",X"02",X"C3",X"68",X"4D",X"CD",X"CF",X"00",X"BA",X"D0",X"04",X"C3",X"68",
		X"4D",X"CD",X"CF",X"00",X"C2",X"D0",X"04",X"C3",X"68",X"4D",X"CD",X"CF",X"00",X"CA",X"D0",X"06",
		X"C3",X"68",X"4D",X"3E",X"0D",X"CD",X"18",X"60",X"C9",X"3A",X"70",X"80",X"FE",X"00",X"28",X"08",
		X"3A",X"14",X"80",X"E6",X"18",X"0F",X"0F",X"0F",X"21",X"7E",X"4D",X"C3",X"EA",X"00",X"86",X"4D",
		X"90",X"4D",X"9B",X"4D",X"A6",X"4D",X"3A",X"A8",X"81",X"3C",X"32",X"A8",X"81",X"C3",X"B1",X"4D",
		X"3A",X"A8",X"81",X"C6",X"02",X"32",X"A8",X"81",X"C3",X"B1",X"4D",X"3A",X"A8",X"81",X"C6",X"04",
		X"32",X"A8",X"81",X"C3",X"B1",X"4D",X"3A",X"A8",X"81",X"C6",X"08",X"32",X"A8",X"81",X"C3",X"B1",
		X"4D",X"3A",X"A8",X"81",X"FE",X"20",X"DA",X"BE",X"4D",X"3E",X"1F",X"32",X"A8",X"81",X"C9",X"3A",
		X"70",X"80",X"FE",X"00",X"28",X"08",X"3A",X"14",X"80",X"E6",X"60",X"07",X"07",X"07",X"21",X"D4",
		X"4D",X"C3",X"EA",X"00",X"DC",X"4D",X"E6",X"4D",X"FC",X"4D",X"07",X"4E",X"3A",X"A9",X"81",X"3C",
		X"32",X"A9",X"81",X"C3",X"12",X"4E",X"3A",X"AA",X"81",X"3C",X"E6",X"01",X"32",X"AA",X"81",X"C2",
		X"12",X"4E",X"3A",X"A9",X"81",X"3C",X"32",X"A9",X"81",X"C3",X"12",X"4E",X"3A",X"A9",X"81",X"C6",
		X"02",X"32",X"A9",X"81",X"C3",X"12",X"4E",X"3A",X"A9",X"81",X"C6",X"04",X"32",X"A9",X"81",X"C3",
		X"12",X"4E",X"3A",X"A9",X"81",X"FE",X"20",X"DA",X"1F",X"4E",X"3E",X"13",X"32",X"A9",X"81",X"C9",
		X"01",X"1C",X"02",X"CD",X"ED",X"00",X"C9",X"21",X"39",X"DE",X"01",X"06",X"00",X"3A",X"A0",X"81",
		X"3D",X"CD",X"F6",X"00",X"23",X"7E",X"F5",X"2B",X"7E",X"21",X"00",X"D6",X"01",X"10",X"00",X"CD",
		X"F6",X"00",X"11",X"90",X"8C",X"ED",X"B0",X"F1",X"F5",X"21",X"00",X"D7",X"01",X"10",X"00",X"CD",
		X"F6",X"00",X"11",X"A0",X"8C",X"ED",X"B0",X"F1",X"21",X"80",X"D7",X"01",X"10",X"00",X"CD",X"F6",
		X"00",X"11",X"80",X"8C",X"ED",X"B0",X"21",X"3C",X"DE",X"01",X"06",X"00",X"3A",X"A0",X"81",X"3D",
		X"CD",X"F6",X"00",X"7E",X"21",X"80",X"D6",X"01",X"10",X"00",X"CD",X"F6",X"00",X"11",X"50",X"8C",
		X"ED",X"B0",X"C9",X"3A",X"17",X"80",X"B7",X"CA",X"B4",X"4E",X"3A",X"26",X"80",X"B7",X"CA",X"A4",
		X"4E",X"3A",X"27",X"80",X"B7",X"C2",X"9D",X"4E",X"3A",X"CD",X"81",X"18",X"03",X"3A",X"B4",X"81",
		X"B7",X"F2",X"B4",X"4E",X"3A",X"02",X"B0",X"E6",X"08",X"C2",X"BE",X"4E",X"3A",X"02",X"B0",X"E6",
		X"04",X"C2",X"B7",X"4E",X"3E",X"00",X"C9",X"3E",X"01",X"32",X"8B",X"80",X"18",X"0D",X"3A",X"17",
		X"80",X"FE",X"02",X"DA",X"B4",X"4E",X"3E",X"02",X"32",X"8B",X"80",X"3E",X"01",X"C9",X"00",X"21",
		X"D0",X"D8",X"3A",X"A0",X"81",X"3D",X"FE",X"20",X"DA",X"DD",X"4E",X"3E",X"1F",X"01",X"08",X"00",
		X"CD",X"F6",X"00",X"11",X"D2",X"80",X"ED",X"B0",X"11",X"01",X"00",X"ED",X"53",X"DA",X"80",X"2A",
		X"D8",X"80",X"22",X"DC",X"80",X"3A",X"48",X"82",X"FE",X"01",X"CA",X"02",X"4F",X"3A",X"A9",X"81",
		X"18",X"03",X"CD",X"BF",X"4D",X"21",X"B8",X"DB",X"01",X"14",X"00",X"CD",X"F6",X"00",X"11",X"5C",
		X"82",X"ED",X"B0",X"2A",X"5E",X"82",X"22",X"70",X"82",X"2A",X"62",X"82",X"22",X"72",X"82",X"2A",
		X"66",X"82",X"22",X"74",X"82",X"3A",X"48",X"82",X"FE",X"01",X"CA",X"32",X"4F",X"3A",X"A8",X"81",
		X"18",X"03",X"CD",X"69",X"4D",X"21",X"D8",X"D9",X"01",X"0C",X"00",X"CD",X"F6",X"00",X"11",X"C0",
		X"80",X"ED",X"B0",X"2A",X"C6",X"80",X"22",X"CC",X"80",X"2A",X"C8",X"80",X"22",X"CD",X"80",X"2A",
		X"CA",X"80",X"22",X"CF",X"80",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CD",X"C9",X"47",X"C3",X"77",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C3",X"29",X"4C",X"C3",X"3D",X"43",X"C3",X"D9",X"4B",X"C3",X"E6",X"42",X"C3",X"E6",X"42",X"00",
		X"CD",X"09",X"50",X"00",X"00",X"00",X"C3",X"C3",X"00",X"3A",X"70",X"80",X"B7",X"CA",X"30",X"50",
		X"CD",X"31",X"50",X"B7",X"CA",X"30",X"50",X"DD",X"21",X"21",X"CA",X"CD",X"D2",X"00",X"11",X"E2",
		X"80",X"21",X"9C",X"81",X"01",X"04",X"00",X"ED",X"B0",X"DD",X"21",X"55",X"CA",X"CD",X"D5",X"00",
		X"C9",X"DD",X"21",X"9F",X"81",X"21",X"E5",X"80",X"01",X"04",X"00",X"7E",X"DD",X"BE",X"00",X"DA",
		X"4D",X"50",X"C2",X"52",X"50",X"DD",X"2B",X"2B",X"10",X"F1",X"C3",X"52",X"50",X"3E",X"01",X"C3",
		X"53",X"50",X"AF",X"C9",X"0F",X"0F",X"0F",X"0F",X"C9",X"3A",X"00",X"B0",X"E6",X"40",X"CA",X"6B",
		X"50",X"3E",X"01",X"32",X"74",X"80",X"3E",X"01",X"32",X"77",X"80",X"C9",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3E",X"00",X"32",X"95",X"80",X"32",X"8D",X"80",X"32",X"88",X"80",X"3A",X"70",X"80",X"FE",X"00",
		X"20",X"15",X"DD",X"21",X"40",X"83",X"DD",X"36",X"02",X"AC",X"DD",X"36",X"03",X"2F",X"DD",X"36",
		X"04",X"70",X"DD",X"36",X"05",X"73",X"C9",X"3E",X"FF",X"32",X"94",X"80",X"3E",X"00",X"32",X"6C",
		X"84",X"3E",X"01",X"32",X"6E",X"80",X"3A",X"6E",X"80",X"FE",X"00",X"28",X"03",X"00",X"18",X"F6",
		X"DD",X"21",X"6C",X"84",X"DD",X"7E",X"00",X"E6",X"07",X"FE",X"05",X"28",X"63",X"06",X"00",X"3E",
		X"14",X"FE",X"00",X"28",X"08",X"DD",X"70",X"00",X"DD",X"23",X"3D",X"18",X"F4",X"DD",X"21",X"6C",
		X"84",X"3E",X"8B",X"32",X"14",X"88",X"FD",X"21",X"00",X"88",X"FD",X"36",X"00",X"0B",X"21",X"48",
		X"0D",X"22",X"01",X"88",X"FD",X"36",X"03",X"02",X"FD",X"36",X"04",X"01",X"FD",X"36",X"05",X"01",
		X"FD",X"36",X"06",X"01",X"FD",X"36",X"07",X"02",X"FD",X"36",X"08",X"00",X"21",X"00",X"00",X"22",
		X"B4",X"8C",X"DD",X"CB",X"00",X"D6",X"DD",X"CB",X"00",X"8E",X"DD",X"CB",X"00",X"C6",X"DD",X"36",
		X"06",X"03",X"DD",X"36",X"08",X"EE",X"DD",X"36",X"0A",X"03",X"CD",X"43",X"52",X"C3",X"31",X"51",
		X"DD",X"7E",X"0B",X"FE",X"84",X"DA",X"D6",X"51",X"DD",X"CB",X"00",X"CE",X"DD",X"36",X"01",X"00",
		X"FD",X"21",X"00",X"85",X"3E",X"40",X"FE",X"00",X"28",X"09",X"FD",X"36",X"00",X"00",X"FD",X"23",
		X"3D",X"18",X"F3",X"C3",X"1E",X"52",X"DD",X"7E",X"0B",X"FE",X"48",X"DA",X"E1",X"51",X"C3",X"15",
		X"52",X"DD",X"7E",X"0B",X"FE",X"10",X"DA",X"F4",X"51",X"2A",X"75",X"84",X"11",X"0C",X"00",X"ED",
		X"52",X"22",X"75",X"84",X"2A",X"71",X"84",X"ED",X"5B",X"75",X"84",X"19",X"22",X"71",X"84",X"2A",
		X"73",X"84",X"ED",X"52",X"22",X"73",X"84",X"DD",X"7E",X"0C",X"FE",X"50",X"D2",X"15",X"52",X"DD",
		X"86",X"0A",X"DD",X"77",X"0C",X"CD",X"43",X"52",X"DD",X"34",X"0B",X"C3",X"31",X"51",X"3E",X"00",
		X"32",X"94",X"80",X"3E",X"89",X"32",X"00",X"88",X"3E",X"8B",X"32",X"14",X"88",X"3A",X"A0",X"81",
		X"FE",X"06",X"30",X"0E",X"3D",X"87",X"47",X"3E",X"0A",X"90",X"47",X"3A",X"B3",X"81",X"80",X"32",
		X"B3",X"81",X"C9",X"FD",X"E5",X"DD",X"36",X"02",X"0B",X"DD",X"7E",X"0B",X"FE",X"48",X"20",X"11",
		X"21",X"00",X"0D",X"22",X"01",X"88",X"3E",X"02",X"32",X"05",X"88",X"21",X"C0",X"00",X"22",X"B2",
		X"8C",X"DD",X"7E",X"0B",X"FE",X"48",X"38",X"10",X"CB",X"4F",X"28",X"0C",X"3A",X"B2",X"8C",X"FE",
		X"00",X"28",X"05",X"D6",X"10",X"32",X"B2",X"8C",X"DD",X"36",X"04",X"7A",X"DD",X"7E",X"0C",X"FE",
		X"10",X"DA",X"00",X"53",X"FE",X"20",X"DA",X"DA",X"52",X"FE",X"30",X"DA",X"B4",X"52",X"DD",X"36",
		X"01",X"40",X"DD",X"7E",X"06",X"D6",X"30",X"DD",X"77",X"03",X"FD",X"21",X"00",X"85",X"CD",X"25",
		X"53",X"DD",X"36",X"01",X"47",X"DD",X"7E",X"08",X"C6",X"30",X"DD",X"77",X"03",X"FD",X"21",X"38",
		X"85",X"CD",X"25",X"53",X"DD",X"36",X"01",X"41",X"DD",X"7E",X"06",X"D6",X"20",X"DD",X"77",X"03",
		X"FD",X"21",X"08",X"85",X"CD",X"25",X"53",X"DD",X"36",X"01",X"46",X"DD",X"7E",X"08",X"C6",X"20",
		X"DD",X"77",X"03",X"FD",X"21",X"30",X"85",X"CD",X"25",X"53",X"DD",X"36",X"01",X"42",X"DD",X"7E",
		X"06",X"D6",X"10",X"DD",X"77",X"03",X"FD",X"21",X"10",X"85",X"CD",X"25",X"53",X"DD",X"36",X"01",
		X"45",X"DD",X"7E",X"08",X"C6",X"10",X"DD",X"77",X"03",X"FD",X"21",X"28",X"85",X"CD",X"25",X"53",
		X"DD",X"36",X"01",X"43",X"DD",X"7E",X"06",X"DD",X"77",X"03",X"FD",X"21",X"18",X"85",X"CD",X"25",
		X"53",X"DD",X"36",X"01",X"44",X"DD",X"7E",X"08",X"DD",X"77",X"03",X"FD",X"21",X"20",X"85",X"CD",
		X"25",X"53",X"FD",X"E1",X"C9",X"DD",X"7E",X"01",X"FD",X"77",X"00",X"DD",X"7E",X"02",X"FD",X"77",
		X"01",X"DD",X"7E",X"03",X"FD",X"77",X"02",X"DD",X"7E",X"04",X"FD",X"77",X"03",X"C9",X"3E",X"FF",
		X"32",X"94",X"80",X"3E",X"01",X"32",X"6E",X"80",X"3A",X"6E",X"80",X"FE",X"00",X"28",X"03",X"00",
		X"18",X"F6",X"DD",X"21",X"6C",X"84",X"DD",X"7E",X"00",X"E6",X"0F",X"FE",X"05",X"28",X"77",X"DD",
		X"36",X"00",X"05",X"DD",X"36",X"01",X"AC",X"DD",X"36",X"02",X"2B",X"3A",X"02",X"85",X"DD",X"77",
		X"03",X"3A",X"03",X"85",X"DD",X"77",X"04",X"21",X"00",X"00",X"22",X"71",X"84",X"22",X"77",X"84",
		X"21",X"FF",X"0F",X"22",X"BE",X"8C",X"3E",X"8B",X"32",X"14",X"88",X"DD",X"7E",X"03",X"21",X"80",
		X"01",X"FE",X"71",X"38",X"03",X"CD",X"F3",X"1F",X"22",X"73",X"84",X"DD",X"7E",X"04",X"21",X"80",
		X"01",X"FE",X"73",X"38",X"03",X"CD",X"F3",X"1F",X"22",X"75",X"84",X"11",X"71",X"00",X"21",X"00",
		X"00",X"DD",X"6E",X"03",X"ED",X"52",X"CD",X"F0",X"1F",X"4D",X"21",X"00",X"00",X"DD",X"6E",X"04",
		X"11",X"73",X"00",X"ED",X"52",X"CD",X"F0",X"1F",X"7D",X"B9",X"38",X"04",X"DD",X"CB",X"00",X"F6",
		X"CD",X"C2",X"54",X"C3",X"3E",X"53",X"DD",X"7E",X"0B",X"FE",X"10",X"30",X"09",X"CD",X"96",X"54",
		X"DD",X"34",X"0B",X"C3",X"3E",X"53",X"DD",X"7E",X"00",X"E6",X"30",X"FE",X"30",X"28",X"0F",X"CD",
		X"96",X"54",X"DD",X"34",X"0B",X"CD",X"24",X"54",X"CD",X"C2",X"54",X"C3",X"3E",X"53",X"DD",X"7E",
		X"0B",X"FE",X"FE",X"30",X"16",X"3E",X"01",X"32",X"6E",X"80",X"3A",X"6E",X"80",X"FE",X"00",X"28",
		X"02",X"18",X"F7",X"CD",X"96",X"54",X"DD",X"34",X"0B",X"18",X"E3",X"3E",X"00",X"32",X"94",X"80",
		X"32",X"00",X"85",X"C9",X"DD",X"CB",X"00",X"76",X"C2",X"61",X"54",X"21",X"00",X"00",X"DD",X"6E",
		X"03",X"11",X"71",X"00",X"ED",X"52",X"CD",X"F0",X"1F",X"7D",X"FE",X"02",X"28",X"02",X"30",X"0E",
		X"DD",X"CB",X"00",X"E6",X"DD",X"CB",X"00",X"F6",X"DD",X"36",X"03",X"71",X"18",X"D6",X"DD",X"66",
		X"03",X"DD",X"6E",X"05",X"ED",X"5B",X"73",X"84",X"19",X"DD",X"74",X"03",X"DD",X"75",X"05",X"18",
		X"34",X"21",X"00",X"00",X"DD",X"6E",X"04",X"11",X"73",X"00",X"ED",X"52",X"CD",X"F0",X"1F",X"7D",
		X"FE",X"02",X"28",X"02",X"30",X"0E",X"DD",X"CB",X"00",X"EE",X"DD",X"CB",X"00",X"B6",X"DD",X"36",
		X"04",X"73",X"18",X"11",X"DD",X"66",X"04",X"DD",X"6E",X"06",X"ED",X"5B",X"75",X"84",X"19",X"DD",
		X"74",X"04",X"DD",X"75",X"06",X"C9",X"3A",X"77",X"84",X"E6",X"07",X"FE",X"00",X"20",X"22",X"DD",
		X"34",X"0C",X"DD",X"7E",X"0C",X"FE",X"07",X"38",X"05",X"3E",X"00",X"32",X"78",X"84",X"87",X"16",
		X"00",X"5F",X"FD",X"21",X"DB",X"54",X"FD",X"19",X"FD",X"66",X"01",X"FD",X"6E",X"00",X"22",X"BE",
		X"8C",X"C9",X"DD",X"7E",X"01",X"32",X"00",X"85",X"DD",X"7E",X"02",X"32",X"01",X"85",X"DD",X"7E",
		X"03",X"32",X"02",X"85",X"DD",X"7E",X"04",X"32",X"03",X"85",X"C9",X"FF",X"0F",X"AF",X"0A",X"5F",
		X"05",X"0F",X"00",X"0F",X"00",X"5F",X"05",X"AF",X"0A",X"C9",X"E5",X"DD",X"E5",X"C5",X"FD",X"E5",
		X"3E",X"00",X"32",X"A6",X"81",X"3A",X"A2",X"81",X"FE",X"00",X"CA",X"69",X"55",X"3A",X"A0",X"81",
		X"3D",X"26",X"00",X"6F",X"06",X"00",X"4F",X"29",X"29",X"09",X"09",X"01",X"38",X"DE",X"09",X"23",
		X"23",X"23",X"23",X"7E",X"26",X"00",X"6F",X"29",X"44",X"4D",X"29",X"29",X"09",X"01",X"80",X"D8",
		X"09",X"E5",X"FD",X"E1",X"FD",X"7E",X"05",X"32",X"A0",X"85",X"FD",X"7E",X"06",X"32",X"A1",X"85",
		X"FD",X"7E",X"07",X"32",X"A2",X"85",X"FD",X"7E",X"08",X"32",X"A3",X"85",X"FD",X"7E",X"09",X"32",
		X"A4",X"85",X"DD",X"21",X"80",X"84",X"DD",X"7E",X"00",X"FE",X"FF",X"CA",X"69",X"55",X"DD",X"CB",
		X"00",X"76",X"C2",X"61",X"55",X"DD",X"46",X"01",X"DD",X"4E",X"02",X"CD",X"DE",X"00",X"CD",X"70",
		X"55",X"01",X"05",X"00",X"DD",X"09",X"C3",X"46",X"55",X"FD",X"E1",X"C1",X"DD",X"E1",X"E1",X"C9",
		X"E5",X"D5",X"DD",X"E5",X"E5",X"DD",X"E1",X"11",X"00",X"04",X"DD",X"19",X"FD",X"46",X"04",X"FD",
		X"7E",X"02",X"77",X"DD",X"70",X"00",X"DD",X"23",X"23",X"FD",X"7E",X"03",X"77",X"DD",X"70",X"00",
		X"11",X"DF",X"FF",X"ED",X"5A",X"DD",X"19",X"FD",X"7E",X"00",X"77",X"DD",X"70",X"00",X"DD",X"23",
		X"23",X"FD",X"7E",X"01",X"77",X"DD",X"70",X"00",X"DD",X"E1",X"D1",X"E1",X"C9",X"C5",X"D5",X"DD",
		X"E5",X"FD",X"E5",X"DD",X"21",X"A3",X"81",X"FD",X"21",X"80",X"84",X"DD",X"46",X"00",X"0E",X"08",
		X"FD",X"7E",X"00",X"FE",X"FF",X"CA",X"E8",X"55",X"CB",X"40",X"28",X"04",X"FD",X"CB",X"00",X"F6",
		X"11",X"05",X"00",X"FD",X"19",X"0D",X"79",X"FE",X"00",X"28",X"05",X"CB",X"38",X"C3",X"C0",X"55",
		X"11",X"01",X"00",X"DD",X"19",X"C3",X"BB",X"55",X"FD",X"E1",X"DD",X"E1",X"D1",X"C1",X"C9",X"C5",
		X"D5",X"DD",X"E5",X"FD",X"E5",X"DD",X"21",X"A3",X"81",X"FD",X"21",X"80",X"84",X"06",X"00",X"0E",
		X"08",X"FD",X"7E",X"00",X"FE",X"FF",X"CA",X"2A",X"56",X"CB",X"38",X"FD",X"CB",X"00",X"76",X"28",
		X"02",X"CB",X"F8",X"11",X"05",X"00",X"FD",X"19",X"0D",X"79",X"FE",X"00",X"C2",X"01",X"56",X"DD",
		X"70",X"00",X"11",X"01",X"00",X"DD",X"19",X"C3",X"FD",X"55",X"FD",X"E1",X"DD",X"E1",X"D1",X"C1",
		X"C9",X"C5",X"D5",X"E5",X"FD",X"E5",X"21",X"00",X"70",X"DD",X"7E",X"01",X"FE",X"02",X"38",X"08",
		X"FD",X"23",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"87",X"16",X"00",X"5F",X"19",X"FD",X"7E",X"02",
		X"56",X"82",X"47",X"FD",X"7E",X"03",X"23",X"56",X"82",X"4F",X"CD",X"DE",X"00",X"E5",X"FD",X"E1",
		X"11",X"00",X"00",X"DD",X"7E",X"01",X"FE",X"01",X"28",X"24",X"DD",X"CB",X"0B",X"7E",X"28",X"0C",
		X"FD",X"7E",X"FF",X"CD",X"FC",X"56",X"FE",X"00",X"28",X"02",X"CB",X"DB",X"DD",X"CB",X"0B",X"7E",
		X"20",X"0C",X"FD",X"7E",X"01",X"CD",X"FC",X"56",X"FE",X"00",X"28",X"02",X"CB",X"D3",X"DD",X"CB",
		X"09",X"7E",X"28",X"0C",X"FD",X"7E",X"20",X"CD",X"FC",X"56",X"FE",X"00",X"28",X"02",X"CB",X"CB",
		X"DD",X"CB",X"09",X"7E",X"20",X"0C",X"FD",X"7E",X"E0",X"CD",X"FC",X"56",X"FE",X"00",X"28",X"02",
		X"CB",X"C3",X"DD",X"7E",X"01",X"FE",X"01",X"C2",X"F5",X"56",X"FD",X"E1",X"FD",X"E5",X"FD",X"7E",
		X"02",X"C6",X"01",X"47",X"FD",X"7E",X"03",X"C6",X"08",X"4F",X"CD",X"DE",X"00",X"23",X"7E",X"CD",
		X"FC",X"56",X"FE",X"00",X"28",X"04",X"CB",X"D3",X"18",X"1B",X"FD",X"7E",X"02",X"C6",X"0E",X"47",
		X"FD",X"7E",X"03",X"C6",X"08",X"4F",X"CD",X"DE",X"00",X"23",X"7E",X"CD",X"FC",X"56",X"FE",X"00",
		X"CA",X"F5",X"56",X"CB",X"D3",X"7B",X"FD",X"E1",X"E1",X"D1",X"C1",X"C9",X"FE",X"60",X"38",X"0C",
		X"FE",X"80",X"38",X"0A",X"FE",X"A0",X"38",X"04",X"FE",X"C0",X"38",X"02",X"3E",X"00",X"C9",X"3A",
		X"AB",X"81",X"FE",X"14",X"DA",X"09",X"58",X"3E",X"2B",X"CD",X"FC",X"00",X"3E",X"00",X"32",X"82",
		X"89",X"32",X"83",X"89",X"32",X"84",X"89",X"3E",X"00",X"32",X"AC",X"81",X"CD",X"CF",X"00",X"0E",
		X"70",X"0F",X"3A",X"AB",X"81",X"FE",X"14",X"20",X"14",X"3E",X"0F",X"CD",X"18",X"60",X"CD",X"CF",
		X"00",X"D4",X"71",X"02",X"16",X"0A",X"3E",X"01",X"32",X"84",X"89",X"18",X"49",X"F5",X"3E",X"0F",
		X"CD",X"18",X"60",X"F1",X"FE",X"15",X"20",X"14",X"3E",X"0F",X"CD",X"18",X"60",X"CD",X"CF",X"00",
		X"D8",X"71",X"02",X"16",X"14",X"3E",X"02",X"32",X"84",X"89",X"18",X"2A",X"FE",X"16",X"20",X"14",
		X"3E",X"0F",X"CD",X"18",X"60",X"CD",X"CF",X"00",X"DC",X"71",X"02",X"16",X"1E",X"3E",X"03",X"32",
		X"84",X"89",X"18",X"12",X"3E",X"0E",X"CD",X"18",X"60",X"CD",X"CF",X"00",X"E0",X"71",X"02",X"16",
		X"32",X"3E",X"05",X"32",X"84",X"89",X"06",X"00",X"3E",X"01",X"32",X"6E",X"80",X"3A",X"6E",X"80",
		X"FE",X"00",X"20",X"F9",X"04",X"78",X"FE",X"78",X"20",X"EE",X"1E",X"00",X"3E",X"01",X"32",X"6E",
		X"80",X"3A",X"6E",X"80",X"FE",X"00",X"20",X"F9",X"7A",X"FE",X"00",X"28",X"28",X"1C",X"7B",X"E6",
		X"03",X"20",X"E9",X"01",X"00",X"10",X"CD",X"E4",X"00",X"3A",X"83",X"89",X"D6",X"0A",X"27",X"32",
		X"83",X"89",X"3A",X"84",X"89",X"DE",X"00",X"27",X"32",X"84",X"89",X"DD",X"21",X"44",X"72",X"CD",
		X"D5",X"00",X"15",X"18",X"C7",X"3E",X"00",X"32",X"F3",X"91",X"32",X"B3",X"91",X"32",X"93",X"91",
		X"06",X"00",X"3E",X"01",X"32",X"6E",X"80",X"3A",X"6E",X"80",X"FE",X"00",X"20",X"F9",X"04",X"78",
		X"FE",X"3C",X"20",X"EE",X"3E",X"AB",X"CD",X"FC",X"00",X"3E",X"00",X"32",X"AB",X"81",X"32",X"00",
		X"89",X"32",X"01",X"89",X"C9",X"DD",X"21",X"28",X"80",X"DD",X"36",X"02",X"00",X"DD",X"36",X"03",
		X"00",X"DD",X"36",X"04",X"00",X"DD",X"36",X"05",X"00",X"DD",X"36",X"06",X"14",X"DD",X"36",X"07",
		X"15",X"FD",X"21",X"18",X"85",X"FD",X"36",X"00",X"14",X"FD",X"36",X"01",X"0C",X"FD",X"36",X"02",
		X"78",X"FD",X"36",X"03",X"78",X"FD",X"36",X"08",X"AE",X"FD",X"36",X"09",X"2B",X"FD",X"36",X"0A",
		X"60",X"FD",X"36",X"0B",X"60",X"FD",X"36",X"10",X"AF",X"FD",X"36",X"11",X"2B",X"FD",X"36",X"12",
		X"80",X"FD",X"36",X"13",X"60",X"FD",X"36",X"18",X"B0",X"FD",X"36",X"19",X"2B",X"FD",X"36",X"1A",
		X"60",X"FD",X"36",X"1B",X"80",X"FD",X"36",X"20",X"B1",X"FD",X"36",X"21",X"2B",X"FD",X"36",X"22",
		X"80",X"FD",X"36",X"23",X"80",X"3E",X"01",X"32",X"6E",X"80",X"3A",X"6E",X"80",X"FE",X"00",X"28",
		X"03",X"00",X"18",X"F6",X"DD",X"34",X"02",X"3A",X"2A",X"80",X"FE",X"3C",X"38",X"07",X"DD",X"36",
		X"02",X"00",X"DD",X"34",X"03",X"DD",X"34",X"04",X"3A",X"2C",X"80",X"FE",X"04",X"38",X"07",X"CD",
		X"DB",X"59",X"DD",X"36",X"04",X"00",X"DD",X"34",X"05",X"3A",X"2D",X"80",X"FE",X"04",X"38",X"67",
		X"DD",X"36",X"05",X"00",X"3A",X"2E",X"80",X"FE",X"FF",X"28",X"06",X"CD",X"30",X"59",X"DD",X"35",
		X"06",X"3A",X"2F",X"80",X"FE",X"FF",X"28",X"06",X"CD",X"86",X"59",X"DD",X"35",X"07",X"3A",X"2B",
		X"80",X"FE",X"03",X"20",X"42",X"3A",X"2A",X"80",X"FE",X"10",X"20",X"0C",X"3E",X"00",X"32",X"40",
		X"85",X"3E",X"0A",X"32",X"41",X"85",X"18",X"2F",X"3A",X"2A",X"80",X"FE",X"0C",X"28",X"02",X"30",
		X"26",X"FE",X"00",X"20",X"1F",X"3A",X"17",X"80",X"FE",X"99",X"30",X"08",X"C6",X"01",X"27",X"32",
		X"17",X"80",X"18",X"09",X"3A",X"87",X"80",X"C6",X"01",X"27",X"32",X"87",X"80",X"CD",X"F0",X"00",
		X"DD",X"21",X"28",X"80",X"CD",X"F2",X"59",X"3A",X"2B",X"80",X"FE",X"0B",X"DA",X"85",X"58",X"C9",
		X"DD",X"E5",X"DD",X"21",X"B6",X"92",X"FD",X"21",X"B6",X"96",X"21",X"68",X"D2",X"01",X"00",X"00",
		X"79",X"FE",X"14",X"28",X"03",X"D2",X"83",X"59",X"DD",X"36",X"00",X"00",X"FD",X"36",X"00",X"0A",
		X"78",X"FE",X"00",X"20",X"1B",X"3A",X"2E",X"80",X"B9",X"28",X"02",X"30",X"13",X"7E",X"FE",X"FF",
		X"20",X"04",X"06",X"01",X"18",X"0A",X"7E",X"DD",X"77",X"00",X"23",X"7E",X"FD",X"77",X"00",X"23",
		X"79",X"FE",X"0E",X"38",X"04",X"DD",X"2B",X"FD",X"2B",X"11",X"E0",X"FF",X"DD",X"19",X"FD",X"19",
		X"0C",X"18",X"BD",X"DD",X"E1",X"C9",X"DD",X"E5",X"DD",X"21",X"37",X"91",X"FD",X"21",X"37",X"95",
		X"21",X"83",X"D2",X"01",X"00",X"00",X"79",X"FE",X"15",X"28",X"02",X"30",X"3B",X"DD",X"36",X"00",
		X"00",X"FD",X"36",X"00",X"0A",X"78",X"FE",X"00",X"20",X"1B",X"3A",X"2F",X"80",X"B9",X"28",X"02",
		X"30",X"13",X"7E",X"FE",X"FF",X"20",X"04",X"06",X"01",X"18",X"0A",X"7E",X"DD",X"77",X"00",X"23",
		X"7E",X"FD",X"77",X"00",X"23",X"79",X"FE",X"0D",X"38",X"04",X"DD",X"2B",X"FD",X"2B",X"11",X"20",
		X"00",X"DD",X"19",X"FD",X"19",X"0C",X"18",X"BE",X"DD",X"E1",X"C9",X"C5",X"3A",X"18",X"85",X"4F",
		X"E6",X"03",X"FE",X"03",X"20",X"05",X"79",X"E6",X"FC",X"18",X"02",X"0C",X"79",X"32",X"18",X"85",
		X"C1",X"C9",X"3E",X"AD",X"32",X"40",X"85",X"3E",X"3B",X"32",X"41",X"85",X"3E",X"8C",X"32",X"42",
		X"85",X"3E",X"D4",X"32",X"43",X"85",X"C9",X"C9",X"C5",X"D5",X"3A",X"AE",X"81",X"FE",X"FF",X"CA",
		X"E3",X"5A",X"3A",X"14",X"80",X"E6",X"07",X"FE",X"00",X"20",X"03",X"C3",X"E3",X"5A",X"FE",X"01",
		X"20",X"05",X"06",X"0A",X"C3",X"59",X"5A",X"FE",X"02",X"20",X"05",X"06",X"03",X"C3",X"59",X"5A",
		X"FE",X"03",X"20",X"05",X"06",X"05",X"C3",X"69",X"5A",X"FE",X"04",X"20",X"05",X"06",X"0A",X"C3",
		X"69",X"5A",X"FE",X"05",X"20",X"07",X"06",X"05",X"0E",X"0A",X"C3",X"7A",X"5A",X"FE",X"06",X"C2",
		X"9F",X"5A",X"06",X"0A",X"0E",X"1E",X"C3",X"7A",X"5A",X"16",X"00",X"3A",X"AD",X"81",X"B8",X"DA",
		X"D4",X"5A",X"14",X"90",X"32",X"AD",X"81",X"18",X"F2",X"3A",X"AD",X"81",X"B8",X"DA",X"E3",X"5A",
		X"16",X"01",X"3E",X"FF",X"32",X"AE",X"81",X"C3",X"D4",X"5A",X"16",X"00",X"3A",X"AE",X"81",X"FE",
		X"01",X"28",X"0D",X"3A",X"AD",X"81",X"B8",X"DA",X"E3",X"5A",X"14",X"3E",X"01",X"32",X"AE",X"81",
		X"3A",X"AD",X"81",X"B9",X"38",X"3E",X"14",X"3E",X"FF",X"32",X"AE",X"81",X"C3",X"D4",X"5A",X"16",
		X"00",X"3A",X"AE",X"81",X"FE",X"01",X"28",X"12",X"FE",X"02",X"28",X"1B",X"3A",X"AD",X"81",X"FE",
		X"05",X"DA",X"E3",X"5A",X"14",X"3E",X"01",X"32",X"AE",X"81",X"3A",X"AD",X"81",X"FE",X"0A",X"38",
		X"13",X"14",X"3E",X"02",X"32",X"AE",X"81",X"3A",X"AD",X"81",X"FE",X"1E",X"38",X"06",X"14",X"3E",
		X"FF",X"32",X"AE",X"81",X"7A",X"FE",X"00",X"28",X"0A",X"3A",X"9B",X"81",X"82",X"32",X"9B",X"81",
		X"CD",X"F3",X"4F",X"D1",X"C1",X"F1",X"C9",X"3A",X"04",X"B0",X"E6",X"03",X"FE",X"03",X"28",X"03",
		X"3C",X"18",X"02",X"3E",X"06",X"32",X"16",X"80",X"3A",X"04",X"B0",X"E6",X"0C",X"CB",X"3F",X"CB",
		X"3F",X"FE",X"01",X"20",X"0E",X"3E",X"FF",X"32",X"84",X"80",X"3E",X"00",X"32",X"85",X"80",X"3E",
		X"01",X"18",X"06",X"FE",X"00",X"20",X"02",X"3E",X"01",X"32",X"83",X"80",X"3A",X"04",X"B0",X"E6",
		X"30",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"FE",X"03",X"28",X"04",X"C6",X"03",X"18",
		X"02",X"3E",X"02",X"32",X"71",X"80",X"3A",X"04",X"B0",X"E6",X"40",X"28",X"02",X"3E",X"01",X"32",
		X"72",X"80",X"3A",X"04",X"B0",X"E6",X"80",X"28",X"02",X"3E",X"01",X"32",X"73",X"80",X"C9",X"DD",
		X"E5",X"DD",X"21",X"00",X"89",X"DD",X"CB",X"00",X"46",X"28",X"0F",X"CD",X"EC",X"2F",X"DD",X"7E",
		X"02",X"32",X"10",X"85",X"DD",X"7E",X"03",X"32",X"11",X"85",X"DD",X"E1",X"C9",X"F5",X"3A",X"8F",
		X"80",X"FE",X"00",X"28",X"52",X"7B",X"FE",X"00",X"28",X"4D",X"FE",X"FF",X"28",X"49",X"C5",X"E5",
		X"DD",X"E5",X"3A",X"A0",X"81",X"3D",X"26",X"00",X"6F",X"29",X"44",X"4D",X"29",X"09",X"DD",X"21",
		X"38",X"DE",X"44",X"4D",X"DD",X"09",X"DD",X"7E",X"02",X"DD",X"E1",X"E1",X"01",X"00",X"00",X"FE",
		X"04",X"38",X"06",X"06",X"10",X"3D",X"3D",X"3D",X"3D",X"FE",X"00",X"28",X"12",X"FE",X"01",X"20",
		X"04",X"0E",X"10",X"18",X"0A",X"FE",X"02",X"20",X"04",X"0E",X"40",X"18",X"02",X"0E",X"50",X"7A",
		X"B7",X"B0",X"57",X"7B",X"81",X"5F",X"C1",X"F1",X"C9",X"F5",X"C5",X"D5",X"E5",X"3A",X"94",X"80",
		X"FE",X"FF",X"CA",X"0B",X"5C",X"3A",X"91",X"80",X"3C",X"32",X"91",X"80",X"FE",X"03",X"DA",X"0B",
		X"5C",X"3E",X"00",X"32",X"91",X"80",X"21",X"0A",X"0F",X"11",X"B2",X"8C",X"01",X"0E",X"00",X"ED",
		X"B0",X"3A",X"92",X"80",X"3C",X"FE",X"07",X"38",X"02",X"3E",X"00",X"32",X"92",X"80",X"87",X"16",
		X"00",X"5F",X"21",X"B2",X"8C",X"19",X"36",X"FF",X"23",X"36",X"0F",X"E1",X"D1",X"C1",X"F1",X"C9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C3",X"E7",X"5A",X"C3",X"6D",X"5B",X"C3",X"FC",X"56",X"C3",X"C9",X"5B",X"00",X"C3",X"07",X"5A",
		X"C3",X"00",X"51",X"C3",X"3E",X"53",X"C3",X"E9",X"54",X"C3",X"EA",X"54",X"C3",X"AD",X"55",X"C3",
		X"EF",X"55",X"C3",X"31",X"56",X"C3",X"0F",X"57",X"C3",X"09",X"50",X"C3",X"15",X"58",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
