library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity galaga_cpu1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of galaga_cpu1 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"3E",X"10",X"32",X"00",X"71",X"C3",X"C4",X"02",X"87",X"30",X"05",X"24",X"C3",X"10",X"00",X"FF",
		X"85",X"6F",X"D0",X"24",X"C9",X"FF",X"FF",X"FF",X"77",X"23",X"10",X"FC",X"C9",X"FF",X"FF",X"FF",
		X"7B",X"D6",X"20",X"5F",X"D0",X"15",X"C9",X"FF",X"21",X"00",X"91",X"06",X"F0",X"AF",X"DF",X"C9",
		X"37",X"08",X"C3",X"B5",X"13",X"FF",X"FF",X"FF",X"C3",X"37",X"02",X"E9",X"21",X"00",X"93",X"06",
		X"80",X"AF",X"DF",X"21",X"00",X"9B",X"06",X"80",X"DF",X"21",X"00",X"88",X"3E",X"80",X"06",X"80",
		X"DF",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"D9",X"ED",X"A0",X"EA",X"8F",X"00",X"F5",X"21",X"00",X"71",
		X"36",X"10",X"3A",X"B9",X"9A",X"A7",X"28",X"16",X"AF",X"32",X"B9",X"9A",X"21",X"92",X"00",X"11",
		X"00",X"70",X"01",X"04",X"00",X"D9",X"3E",X"A8",X"32",X"00",X"71",X"F1",X"ED",X"45",X"F1",X"D9",
		X"ED",X"45",X"10",X"10",X"20",X"20",X"3A",X"08",X"3B",X"08",X"B2",X"17",X"00",X"17",X"86",X"1A",
		X"6A",X"08",X"3A",X"08",X"3A",X"08",X"24",X"29",X"EC",X"1D",X"9E",X"2A",X"B9",X"1D",X"EB",X"23",
		X"AA",X"1E",X"38",X"1D",X"48",X"09",X"6B",X"1B",X"B2",X"19",X"7C",X"1D",X"3A",X"08",X"8B",X"1F",
		X"0A",X"1F",X"3A",X"08",X"D8",X"1D",X"30",X"22",X"D9",X"21",X"3A",X"08",X"3A",X"08",X"F2",X"20",
		X"00",X"20",X"3A",X"08",X"8A",X"09",X"11",X"ED",X"83",X"21",X"B9",X"02",X"01",X"05",X"00",X"ED",
		X"B0",X"1E",X"CB",X"21",X"EB",X"00",X"0E",X"11",X"ED",X"B0",X"C9",X"0E",X"1B",X"18",X"0C",X"1C",
		X"24",X"11",X"10",X"12",X"11",X"24",X"24",X"24",X"24",X"19",X"1E",X"01",X"FF",X"FF",X"FF",X"FF",
		X"14",X"06",X"14",X"0C",X"14",X"08",X"14",X"0A",X"1C",X"00",X"1C",X"12",X"1E",X"00",X"1E",X"12",
		X"1C",X"02",X"1C",X"10",X"1E",X"02",X"1E",X"10",X"1C",X"04",X"1C",X"0E",X"1E",X"04",X"1E",X"0E",
		X"1C",X"06",X"1C",X"0C",X"1E",X"06",X"1E",X"0C",X"1C",X"08",X"1C",X"0A",X"1E",X"08",X"1E",X"0A",
		X"16",X"06",X"16",X"0C",X"16",X"08",X"16",X"0A",X"18",X"00",X"18",X"12",X"1A",X"00",X"1A",X"12",
		X"18",X"02",X"18",X"10",X"1A",X"02",X"1A",X"10",X"18",X"04",X"18",X"0E",X"1A",X"04",X"1A",X"0E",
		X"18",X"06",X"18",X"0C",X"1A",X"06",X"1A",X"0C",X"18",X"08",X"18",X"0A",X"1A",X"08",X"1A",X"0A",
		X"21",X"40",X"80",X"11",X"41",X"80",X"01",X"7F",X"03",X"36",X"24",X"ED",X"B0",X"21",X"40",X"84",
		X"11",X"41",X"84",X"01",X"7F",X"03",X"36",X"00",X"ED",X"B0",X"3E",X"04",X"06",X"20",X"DF",X"3E",
		X"4E",X"06",X"20",X"DF",X"C9",X"21",X"21",X"98",X"34",X"7E",X"3C",X"E6",X"03",X"32",X"25",X"98",
		X"28",X"10",X"0E",X"06",X"F7",X"EB",X"3A",X"21",X"98",X"6F",X"26",X"00",X"CD",X"66",X"0A",X"AF",
		X"18",X"0A",X"0E",X"07",X"F7",X"3E",X"01",X"32",X"AD",X"9A",X"3E",X"08",X"32",X"A8",X"92",X"3E",
		X"03",X"32",X"AE",X"92",X"32",X"0B",X"92",X"3A",X"25",X"98",X"A7",X"08",X"CD",X"7F",X"11",X"3A",
		X"AE",X"92",X"A7",X"20",X"FA",X"3E",X"78",X"32",X"AE",X"92",X"CD",X"A4",X"28",X"CD",X"B0",X"25",
		X"3E",X"02",X"32",X"AC",X"92",X"AF",X"CD",X"D5",X"12",X"AF",X"06",X"30",X"21",X"00",X"92",X"77",
		X"2C",X"2C",X"10",X"FB",X"32",X"09",X"90",X"32",X"10",X"90",X"32",X"04",X"90",X"32",X"88",X"92",
		X"32",X"2C",X"98",X"32",X"41",X"98",X"32",X"42",X"98",X"32",X"26",X"98",X"32",X"B0",X"99",X"32",
		X"24",X"98",X"3C",X"32",X"2D",X"98",X"32",X"6D",X"98",X"32",X"28",X"98",X"32",X"0B",X"90",X"32",
		X"08",X"90",X"32",X"0A",X"90",X"CD",X"00",X"2C",X"21",X"30",X"98",X"11",X"B5",X"01",X"06",X"04",
		X"72",X"2C",X"73",X"2C",X"10",X"FA",X"3A",X"05",X"68",X"CB",X"4F",X"C0",X"0E",X"0B",X"21",X"B0",
		X"83",X"CD",X"B3",X"13",X"C3",X"85",X"01",X"F5",X"08",X"F5",X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",
		X"E5",X"3A",X"04",X"68",X"57",X"3A",X"A0",X"92",X"E6",X"1C",X"4F",X"0F",X"A9",X"E6",X"18",X"4F",
		X"3A",X"BE",X"99",X"CB",X"4A",X"20",X"02",X"3E",X"07",X"E6",X"07",X"B1",X"06",X"05",X"21",X"00",
		X"A0",X"77",X"2C",X"0F",X"10",X"FB",X"32",X"30",X"68",X"AF",X"32",X"20",X"68",X"CB",X"4A",X"CA",
		X"A8",X"02",X"4F",X"21",X"00",X"90",X"79",X"85",X"6F",X"7E",X"A7",X"20",X"03",X"0C",X"18",X"F3",
		X"47",X"21",X"96",X"00",X"79",X"CB",X"27",X"85",X"6F",X"5E",X"23",X"56",X"EB",X"C5",X"CD",X"3B",
		X"00",X"C1",X"78",X"81",X"4F",X"E6",X"E0",X"28",X"DA",X"21",X"00",X"70",X"11",X"B5",X"99",X"01",
		X"03",X"00",X"D9",X"3E",X"71",X"32",X"00",X"71",X"3E",X"01",X"32",X"20",X"68",X"FD",X"E1",X"DD",
		X"E1",X"E1",X"D1",X"C1",X"F1",X"08",X"F1",X"FB",X"C9",X"00",X"00",X"00",X"00",X"02",X"24",X"17",
		X"0A",X"16",X"0C",X"18",X"ED",X"56",X"AF",X"21",X"E0",X"99",X"06",X"10",X"77",X"23",X"10",X"FC",
		X"C3",X"6C",X"33",X"31",X"A0",X"90",X"AF",X"21",X"AC",X"92",X"06",X"04",X"DF",X"21",X"A0",X"9A",
		X"06",X"20",X"DF",X"32",X"07",X"A0",X"32",X"15",X"92",X"32",X"B9",X"99",X"3D",X"21",X"CA",X"92",
		X"06",X"10",X"DF",X"3E",X"01",X"32",X"20",X"68",X"21",X"C0",X"83",X"06",X"40",X"3E",X"24",X"DF",
		X"26",X"80",X"06",X"40",X"DF",X"21",X"00",X"84",X"06",X"40",X"3E",X"03",X"DF",X"CD",X"60",X"01",
		X"11",X"20",X"8A",X"3E",X"05",X"06",X"00",X"21",X"B9",X"02",X"0E",X"06",X"ED",X"B0",X"3D",X"20",
		X"F6",X"21",X"BF",X"02",X"3E",X"2A",X"06",X"05",X"0E",X"FF",X"ED",X"A0",X"2B",X"12",X"1C",X"ED",
		X"A0",X"10",X"F7",X"3E",X"01",X"32",X"01",X"92",X"21",X"05",X"A0",X"36",X"00",X"77",X"CD",X"3C",
		X"00",X"CD",X"D6",X"00",X"CD",X"42",X"12",X"EF",X"3E",X"20",X"32",X"1E",X"90",X"3A",X"B5",X"99",
		X"32",X"B8",X"99",X"AF",X"32",X"1E",X"90",X"32",X"20",X"90",X"AF",X"32",X"07",X"A0",X"32",X"15",
		X"92",X"32",X"12",X"90",X"06",X"80",X"21",X"00",X"92",X"DF",X"3E",X"06",X"32",X"BE",X"99",X"EF",
		X"CD",X"3C",X"00",X"CD",X"42",X"12",X"3A",X"B8",X"99",X"A7",X"3E",X"01",X"28",X"02",X"3E",X"02",
		X"32",X"01",X"92",X"20",X"18",X"AF",X"32",X"03",X"92",X"3C",X"32",X"02",X"90",X"3A",X"01",X"92",
		X"3D",X"28",X"FA",X"CD",X"42",X"12",X"CD",X"60",X"01",X"EF",X"CD",X"3C",X"00",X"AF",X"32",X"0B",
		X"92",X"0E",X"13",X"F7",X"0E",X"01",X"F7",X"21",X"52",X"04",X"22",X"80",X"92",X"3A",X"80",X"99",
		X"FE",X"FF",X"28",X"24",X"5F",X"0E",X"1B",X"CD",X"3D",X"04",X"3A",X"81",X"99",X"FE",X"FF",X"28",
		X"17",X"E6",X"7F",X"5F",X"0E",X"1C",X"CD",X"3D",X"04",X"3A",X"81",X"99",X"CB",X"7F",X"20",X"08",
		X"E6",X"7F",X"5F",X"0E",X"1D",X"CD",X"3D",X"04",X"3A",X"01",X"92",X"FE",X"02",X"28",X"F9",X"32",
		X"B7",X"9A",X"CD",X"60",X"01",X"CD",X"3C",X"00",X"21",X"05",X"A0",X"36",X"00",X"36",X"01",X"21",
		X"20",X"98",X"AF",X"06",X"A0",X"DF",X"32",X"B7",X"9A",X"32",X"B9",X"99",X"3C",X"32",X"AB",X"9A",
		X"32",X"12",X"90",X"32",X"F2",X"98",X"CD",X"66",X"04",X"CD",X"7B",X"12",X"0E",X"04",X"F7",X"21",
		X"AF",X"92",X"36",X"08",X"7E",X"A7",X"20",X"FC",X"21",X"90",X"92",X"06",X"10",X"DF",X"06",X"30",
		X"21",X"B0",X"98",X"DF",X"21",X"B0",X"83",X"0E",X"0B",X"CD",X"B3",X"13",X"3E",X"01",X"32",X"80",
		X"98",X"3A",X"80",X"99",X"32",X"3E",X"98",X"32",X"7E",X"98",X"C3",X"22",X"06",X"F7",X"EB",X"7B",
		X"C6",X"40",X"5F",X"26",X"00",X"CD",X"66",X"0A",X"EB",X"0E",X"1E",X"CD",X"B3",X"13",X"CD",X"9E",
		X"12",X"C9",X"00",X"81",X"19",X"56",X"02",X"81",X"19",X"62",X"04",X"81",X"19",X"6E",X"CD",X"3B",
		X"07",X"CD",X"1E",X"08",X"18",X"F8",X"3A",X"00",X"68",X"4F",X"21",X"B3",X"99",X"3A",X"82",X"99",
		X"CB",X"46",X"28",X"08",X"CB",X"49",X"20",X"04",X"3C",X"87",X"36",X"00",X"32",X"20",X"98",X"32",
		X"60",X"98",X"11",X"F8",X"83",X"21",X"A8",X"04",X"CD",X"99",X"04",X"11",X"E3",X"83",X"21",X"A8",
		X"04",X"3A",X"B3",X"99",X"A7",X"20",X"02",X"23",X"23",X"0E",X"07",X"ED",X"B0",X"21",X"AA",X"04",
		X"11",X"C3",X"83",X"0E",X"04",X"ED",X"B0",X"C9",X"00",X"00",X"24",X"24",X"24",X"24",X"24",X"24",
		X"24",X"E1",X"21",X"AF",X"92",X"36",X"04",X"3A",X"1D",X"90",X"A7",X"28",X"17",X"AF",X"32",X"13",
		X"92",X"3C",X"32",X"25",X"90",X"3A",X"A7",X"92",X"A7",X"C2",X"5E",X"04",X"3A",X"1D",X"90",X"A7",
		X"20",X"FA",X"18",X"1B",X"7E",X"A7",X"20",X"DF",X"CD",X"3B",X"07",X"3A",X"A7",X"92",X"32",X"43",
		X"98",X"4F",X"3A",X"13",X"92",X"B1",X"20",X"0D",X"3A",X"25",X"98",X"A7",X"CA",X"63",X"06",X"CD",
		X"85",X"01",X"C3",X"45",X"06",X"21",X"20",X"98",X"7E",X"35",X"A7",X"C2",X"8C",X"05",X"3A",X"B3",
		X"99",X"A7",X"28",X"0C",X"21",X"4E",X"82",X"3A",X"40",X"98",X"C6",X"04",X"4F",X"CD",X"B3",X"13",
		X"0E",X"02",X"F7",X"CD",X"31",X"13",X"CD",X"31",X"13",X"21",X"18",X"90",X"7E",X"A7",X"20",X"FC",
		X"EF",X"CD",X"3C",X"00",X"CD",X"60",X"01",X"0E",X"15",X"F7",X"0E",X"16",X"F7",X"11",X"32",X"81",
		X"2A",X"46",X"98",X"CD",X"66",X"0A",X"0E",X"18",X"F7",X"11",X"35",X"81",X"2A",X"44",X"98",X"CD",
		X"66",X"0A",X"0E",X"19",X"F7",X"CD",X"85",X"0A",X"EB",X"0E",X"1A",X"CD",X"B3",X"13",X"21",X"AE",
		X"92",X"36",X"0E",X"7E",X"A7",X"20",X"FC",X"CD",X"60",X"01",X"CD",X"00",X"30",X"AF",X"32",X"B0",
		X"9A",X"21",X"AC",X"9A",X"11",X"B6",X"9A",X"1A",X"46",X"B0",X"28",X"09",X"04",X"05",X"28",X"02",
		X"36",X"01",X"76",X"18",X"F2",X"CD",X"60",X"01",X"3A",X"B3",X"99",X"A7",X"CA",X"F1",X"06",X"3A",
		X"60",X"98",X"3C",X"CA",X"F1",X"06",X"3A",X"13",X"92",X"3D",X"20",X"15",X"3A",X"B3",X"99",X"A7",
		X"CA",X"17",X"06",X"3A",X"60",X"98",X"3C",X"CA",X"25",X"06",X"3A",X"13",X"92",X"3D",X"C2",X"25",
		X"06",X"3A",X"A7",X"92",X"A7",X"28",X"06",X"3A",X"87",X"92",X"A7",X"20",X"FA",X"AF",X"32",X"B4",
		X"99",X"3C",X"21",X"0E",X"90",X"77",X"7E",X"A7",X"20",X"FC",X"3A",X"A0",X"9A",X"32",X"48",X"98",
		X"3A",X"AE",X"92",X"32",X"3F",X"98",X"CD",X"0C",X"11",X"CD",X"00",X"2C",X"3A",X"3F",X"98",X"32",
		X"AE",X"92",X"3A",X"48",X"98",X"32",X"A0",X"9A",X"CD",X"7E",X"13",X"3A",X"43",X"98",X"A7",X"28",
		X"03",X"CD",X"B0",X"25",X"3A",X"40",X"98",X"4F",X"3A",X"83",X"99",X"A1",X"32",X"07",X"A0",X"32",
		X"15",X"92",X"3E",X"3F",X"CD",X"D5",X"12",X"37",X"08",X"CD",X"7F",X"11",X"3A",X"43",X"98",X"A7",
		X"28",X"20",X"0E",X"03",X"F7",X"3E",X"80",X"32",X"B4",X"99",X"21",X"0E",X"90",X"3E",X"01",X"77",
		X"7E",X"A7",X"20",X"FC",X"C3",X"25",X"06",X"3A",X"43",X"98",X"A7",X"20",X"14",X"CD",X"85",X"01",
		X"18",X"0F",X"CD",X"85",X"01",X"3A",X"40",X"98",X"C6",X"04",X"4F",X"21",X"6E",X"82",X"CD",X"B3",
		X"13",X"CD",X"3D",X"13",X"3A",X"AE",X"92",X"C6",X"1E",X"FE",X"78",X"38",X"02",X"3E",X"78",X"32",
		X"AE",X"92",X"CD",X"31",X"13",X"3E",X"01",X"32",X"15",X"90",X"32",X"25",X"90",X"32",X"42",X"98",
		X"0E",X"0B",X"21",X"B0",X"83",X"CD",X"B3",X"13",X"0E",X"0B",X"21",X"AE",X"83",X"CD",X"B3",X"13",
		X"C3",X"5E",X"04",X"3A",X"88",X"92",X"5F",X"21",X"AE",X"9A",X"FE",X"28",X"20",X"03",X"21",X"B4",
		X"9A",X"36",X"01",X"CD",X"31",X"13",X"0E",X"08",X"F7",X"CD",X"31",X"13",X"6B",X"26",X"00",X"11",
		X"10",X"81",X"CD",X"66",X"0A",X"CD",X"31",X"13",X"3A",X"88",X"92",X"FE",X"28",X"28",X"1D",X"0E",
		X"09",X"F7",X"CD",X"31",X"13",X"EB",X"3A",X"88",X"92",X"A7",X"28",X"0A",X"6F",X"26",X"00",X"CD",
		X"66",X"0A",X"AF",X"12",X"E7",X"AF",X"12",X"3A",X"88",X"92",X"18",X"21",X"06",X"07",X"3A",X"A0",
		X"92",X"E6",X"0F",X"20",X"F9",X"0E",X"0B",X"CB",X"40",X"28",X"01",X"0C",X"C5",X"F7",X"C1",X"3A",
		X"A0",X"92",X"E6",X"0F",X"28",X"F9",X"10",X"E6",X"0E",X"0D",X"F7",X"3E",X"64",X"21",X"9F",X"92",
		X"86",X"77",X"CD",X"3B",X"07",X"CD",X"31",X"13",X"CD",X"31",X"13",X"21",X"B0",X"83",X"0E",X"0B",
		X"CD",X"B3",X"13",X"21",X"B3",X"83",X"0E",X"0B",X"CD",X"B3",X"13",X"0E",X"0B",X"F7",X"C3",X"EF",
		X"04",X"76",X"F3",X"3A",X"00",X"71",X"FE",X"10",X"20",X"F9",X"21",X"38",X"07",X"11",X"00",X"70",
		X"01",X"03",X"00",X"D9",X"3E",X"61",X"32",X"00",X"71",X"76",X"AF",X"CD",X"4F",X"09",X"FB",X"AF",
		X"06",X"20",X"21",X"A0",X"9A",X"DF",X"11",X"F9",X"83",X"CD",X"3A",X"0A",X"11",X"E4",X"83",X"CD",
		X"3A",X"0A",X"3A",X"B3",X"99",X"3C",X"21",X"E1",X"99",X"86",X"27",X"77",X"D2",X"5A",X"03",X"2B",
		X"7E",X"C6",X"01",X"27",X"77",X"C3",X"5A",X"03",X"02",X"02",X"02",X"3A",X"40",X"98",X"A7",X"3E",
		X"F9",X"28",X"02",X"3E",X"E4",X"DD",X"6F",X"06",X"10",X"21",X"90",X"92",X"EB",X"21",X"0D",X"08",
		X"78",X"D7",X"4E",X"EB",X"7E",X"A7",X"28",X"1D",X"35",X"EB",X"26",X"83",X"DD",X"7D",X"6F",X"79",
		X"E6",X"0F",X"CD",X"EB",X"07",X"DD",X"7D",X"3C",X"6F",X"79",X"07",X"07",X"07",X"07",X"E6",X"0F",
		X"CD",X"EB",X"07",X"18",X"DE",X"2C",X"10",X"D4",X"DD",X"7D",X"C6",X"04",X"5F",X"21",X"F2",X"83",
		X"16",X"83",X"06",X"06",X"1A",X"96",X"C6",X"09",X"FE",X"E5",X"30",X"0F",X"D6",X"0A",X"FE",X"09",
		X"38",X"09",X"3C",X"20",X"0C",X"2D",X"1D",X"10",X"EB",X"18",X"06",X"1A",X"77",X"2D",X"1D",X"10",
		X"FA",X"DD",X"7D",X"C6",X"04",X"6F",X"7E",X"FE",X"24",X"20",X"01",X"AF",X"E6",X"3F",X"07",X"4F",
		X"07",X"07",X"81",X"4F",X"2D",X"7E",X"FE",X"24",X"20",X"01",X"AF",X"81",X"21",X"3E",X"98",X"BE",
		X"C0",X"3A",X"81",X"99",X"47",X"E6",X"7F",X"4F",X"7E",X"B9",X"30",X"03",X"79",X"18",X"01",X"80",
		X"77",X"32",X"AA",X"9A",X"21",X"20",X"98",X"34",X"CD",X"7E",X"13",X"21",X"EB",X"99",X"7E",X"C6",
		X"01",X"27",X"77",X"D0",X"2D",X"7E",X"C6",X"01",X"27",X"77",X"C9",X"A7",X"C8",X"86",X"FE",X"24",
		X"38",X"02",X"D6",X"24",X"FE",X"0A",X"30",X"02",X"77",X"C9",X"D6",X"0A",X"77",X"2C",X"7E",X"FE",
		X"24",X"20",X"01",X"AF",X"FE",X"09",X"28",X"03",X"3C",X"77",X"C9",X"AF",X"18",X"EE",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"08",X"08",X"08",X"05",X"08",X"15",X"00",X"3A",X"08",
		X"90",X"47",X"3A",X"A7",X"92",X"B0",X"20",X"06",X"32",X"A0",X"9A",X"C3",X"B1",X"04",X"3A",X"13",
		X"92",X"A7",X"C8",X"AF",X"32",X"42",X"98",X"C3",X"B1",X"04",X"C9",X"3E",X"01",X"32",X"D6",X"92",
		X"21",X"40",X"8B",X"11",X"C0",X"8B",X"01",X"40",X"00",X"ED",X"B0",X"21",X"40",X"93",X"11",X"C0",
		X"93",X"0E",X"40",X"ED",X"B0",X"21",X"40",X"9B",X"11",X"C0",X"9B",X"0E",X"40",X"ED",X"B0",X"AF",
		X"32",X"D6",X"92",X"3A",X"D7",X"92",X"3D",X"28",X"FA",X"C9",X"3A",X"AE",X"92",X"47",X"FE",X"3C",
		X"30",X"06",X"3A",X"C5",X"99",X"32",X"C4",X"99",X"3A",X"A7",X"92",X"4F",X"3A",X"C0",X"99",X"21",
		X"1C",X"09",X"CD",X"D1",X"08",X"32",X"C8",X"92",X"3A",X"AA",X"92",X"A7",X"28",X"0D",X"21",X"C4",
		X"92",X"3E",X"02",X"06",X"03",X"DF",X"AF",X"32",X"A0",X"9A",X"C9",X"3A",X"C1",X"99",X"21",X"3C",
		X"09",X"CD",X"D1",X"08",X"32",X"C4",X"92",X"3A",X"C2",X"99",X"21",X"E0",X"08",X"CD",X"C0",X"08",
		X"32",X"C5",X"92",X"3A",X"C3",X"99",X"21",X"FE",X"08",X"CD",X"C0",X"08",X"32",X"C6",X"92",X"C9",
		X"5F",X"CB",X"27",X"83",X"D7",X"78",X"FE",X"28",X"30",X"01",X"23",X"A7",X"20",X"01",X"23",X"7E",
		X"C9",X"CB",X"27",X"CF",X"EB",X"61",X"3E",X"0A",X"CD",X"61",X"10",X"EB",X"7A",X"D7",X"7E",X"C9",
		X"09",X"07",X"05",X"08",X"06",X"04",X"07",X"05",X"04",X"06",X"04",X"03",X"05",X"03",X"03",X"04",
		X"03",X"03",X"04",X"02",X"02",X"03",X"03",X"02",X"03",X"02",X"02",X"02",X"02",X"02",X"06",X"05",
		X"04",X"05",X"04",X"03",X"05",X"03",X"03",X"04",X"03",X"02",X"04",X"02",X"02",X"03",X"03",X"02",
		X"03",X"02",X"01",X"02",X"02",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"03",X"03",X"01",X"01",
		X"03",X"03",X"03",X"01",X"07",X"03",X"03",X"01",X"07",X"03",X"03",X"03",X"07",X"07",X"03",X"03",
		X"0F",X"07",X"03",X"03",X"0F",X"07",X"07",X"03",X"0F",X"07",X"07",X"07",X"06",X"0A",X"0F",X"0F",
		X"04",X"08",X"0D",X"0D",X"04",X"06",X"0A",X"0A",X"3A",X"A0",X"92",X"07",X"07",X"07",X"07",X"4F",
		X"3A",X"01",X"92",X"FE",X"03",X"C0",X"3A",X"40",X"98",X"47",X"2F",X"A1",X"21",X"81",X"09",X"11",
		X"D9",X"83",X"CD",X"72",X"09",X"3A",X"B3",X"99",X"A7",X"C8",X"78",X"A1",X"21",X"84",X"09",X"11",
		X"C4",X"83",X"C5",X"E6",X"01",X"28",X"03",X"21",X"87",X"09",X"01",X"03",X"00",X"ED",X"B0",X"C1",
		X"C9",X"19",X"1E",X"01",X"19",X"1E",X"02",X"24",X"24",X"24",X"3A",X"B5",X"99",X"FE",X"BB",X"CA",
		X"6C",X"33",X"3A",X"01",X"92",X"FE",X"03",X"20",X"19",X"21",X"E9",X"99",X"7E",X"C6",X"01",X"27",
		X"FE",X"60",X"20",X"01",X"AF",X"06",X"04",X"3F",X"77",X"2D",X"7E",X"CE",X"00",X"27",X"10",X"F8",
		X"18",X"42",X"3A",X"B8",X"99",X"FE",X"A0",X"11",X"3C",X"80",X"28",X"30",X"3A",X"B5",X"99",X"21",
		X"E2",X"09",X"01",X"06",X"00",X"ED",X"B8",X"1D",X"4F",X"07",X"07",X"07",X"07",X"E6",X"0F",X"28",
		X"02",X"12",X"1D",X"79",X"E6",X"0F",X"12",X"1D",X"3E",X"24",X"12",X"18",X"17",X"1D",X"12",X"0D",
		X"0E",X"1B",X"0C",X"22",X"0A",X"15",X"19",X"24",X"0E",X"0E",X"1B",X"0F",X"21",X"EB",X"09",X"01",
		X"09",X"00",X"ED",X"B8",X"3A",X"01",X"92",X"A7",X"C8",X"3D",X"20",X"16",X"3A",X"B5",X"99",X"A7",
		X"28",X"10",X"3E",X"02",X"32",X"01",X"92",X"AF",X"21",X"A0",X"9A",X"06",X"08",X"DF",X"2C",X"06",
		X"0F",X"DF",X"3A",X"B5",X"99",X"4F",X"3A",X"B8",X"99",X"47",X"91",X"C8",X"38",X"0F",X"27",X"3D",
		X"32",X"B3",X"99",X"79",X"32",X"B8",X"99",X"3E",X"03",X"32",X"01",X"92",X"C9",X"79",X"32",X"B8",
		X"99",X"FE",X"A0",X"C8",X"90",X"27",X"32",X"79",X"9A",X"C9",X"21",X"03",X"91",X"06",X"05",X"1A",
		X"1C",X"FE",X"24",X"20",X"01",X"AF",X"ED",X"67",X"CB",X"40",X"20",X"01",X"2D",X"10",X"F0",X"AF",
		X"ED",X"67",X"2D",X"36",X"00",X"2E",X"03",X"11",X"E5",X"99",X"06",X"04",X"A7",X"1A",X"8E",X"27",
		X"12",X"1D",X"2D",X"10",X"F8",X"C9",X"06",X"01",X"25",X"24",X"20",X"05",X"7D",X"FE",X"0A",X"38",
		X"0A",X"3E",X"0A",X"CD",X"61",X"10",X"F5",X"04",X"18",X"EE",X"F1",X"CD",X"81",X"0A",X"10",X"FA",
		X"C9",X"12",X"C3",X"20",X"00",X"2A",X"44",X"98",X"ED",X"5B",X"46",X"98",X"7A",X"B3",X"20",X"05",
		X"11",X"00",X"00",X"18",X"51",X"CB",X"7A",X"20",X"0A",X"CB",X"7C",X"20",X"06",X"29",X"EB",X"29",
		X"EB",X"18",X"F2",X"7A",X"CD",X"61",X"10",X"E5",X"67",X"2E",X"00",X"7A",X"CD",X"61",X"10",X"E3",
		X"11",X"B0",X"99",X"06",X"04",X"7C",X"26",X"00",X"EB",X"ED",X"6F",X"CB",X"40",X"28",X"01",X"2C",
		X"EB",X"CD",X"19",X"0B",X"08",X"E3",X"CD",X"19",X"0B",X"E3",X"D7",X"08",X"84",X"26",X"00",X"10",
		X"E7",X"D1",X"FE",X"05",X"38",X"14",X"ED",X"5B",X"B0",X"99",X"7A",X"C6",X"01",X"27",X"57",X"30",
		X"05",X"7B",X"C6",X"01",X"27",X"5F",X"ED",X"53",X"B0",X"99",X"06",X"04",X"0E",X"00",X"21",X"B0",
		X"99",X"11",X"38",X"81",X"05",X"20",X"04",X"3E",X"2A",X"12",X"E7",X"04",X"AF",X"ED",X"6F",X"CB",
		X"40",X"28",X"01",X"2C",X"A7",X"20",X"04",X"CB",X"41",X"28",X"04",X"CB",X"C1",X"12",X"E7",X"78",
		X"FE",X"03",X"20",X"02",X"CB",X"C1",X"10",X"DC",X"C9",X"3E",X"0A",X"CD",X"4E",X"10",X"7C",X"26",
		X"00",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C4",
		X"E5",X"ED",X"5F",X"67",X"3A",X"A0",X"92",X"84",X"6F",X"26",X"01",X"7E",X"67",X"ED",X"5F",X"84",
		X"E1",X"C9",X"C5",X"D5",X"7B",X"95",X"06",X"00",X"30",X"04",X"CB",X"C0",X"ED",X"44",X"4F",X"7A",
		X"94",X"30",X"0A",X"57",X"78",X"EE",X"01",X"F6",X"02",X"47",X"7A",X"ED",X"44",X"B9",X"F5",X"17",
		X"A8",X"1F",X"3F",X"CB",X"10",X"F1",X"30",X"03",X"51",X"4F",X"7A",X"61",X"2E",X"00",X"CD",X"61",
		X"10",X"7C",X"A8",X"E6",X"01",X"28",X"03",X"7D",X"2F",X"6F",X"60",X"D1",X"C1",X"C9",X"D5",X"EB",
		X"21",X"00",X"00",X"CB",X"3F",X"30",X"01",X"19",X"CB",X"23",X"CB",X"12",X"A7",X"20",X"F4",X"D1",
		X"C9",X"C5",X"4F",X"AF",X"06",X"11",X"8F",X"38",X"0B",X"B9",X"38",X"01",X"91",X"3F",X"ED",X"6A",
		X"10",X"F4",X"C1",X"C9",X"91",X"37",X"C3",X"6E",X"10",X"7D",X"E6",X"80",X"3C",X"08",X"CB",X"BD",
		X"C3",X"8A",X"10",X"7D",X"0F",X"0F",X"E6",X"80",X"3C",X"08",X"D5",X"11",X"14",X"00",X"06",X"0C",
		X"DD",X"21",X"00",X"91",X"DD",X"CB",X"13",X"46",X"28",X"06",X"DD",X"19",X"10",X"F6",X"D1",X"C9",
		X"D1",X"DD",X"73",X"08",X"DD",X"72",X"09",X"DD",X"36",X"0D",X"01",X"DD",X"36",X"04",X"00",X"DD",
		X"36",X"05",X"01",X"4D",X"DD",X"71",X"10",X"08",X"57",X"36",X"09",X"DD",X"7D",X"2C",X"77",X"3A",
		X"15",X"92",X"5F",X"69",X"26",X"93",X"4E",X"2C",X"46",X"26",X"9B",X"7E",X"0F",X"CB",X"18",X"CB",
		X"43",X"20",X"09",X"08",X"78",X"C6",X"50",X"ED",X"44",X"47",X"08",X"3F",X"DD",X"70",X"01",X"1F",
		X"E6",X"80",X"DD",X"77",X"00",X"79",X"CB",X"43",X"28",X"03",X"C6",X"0D",X"2F",X"CB",X"3F",X"DD",
		X"77",X"03",X"1F",X"E6",X"80",X"DD",X"77",X"02",X"DD",X"72",X"13",X"DD",X"36",X"0E",X"1E",X"3A",
		X"0B",X"92",X"A7",X"28",X"03",X"3A",X"C8",X"92",X"DD",X"77",X"0F",X"C9",X"3E",X"1F",X"32",X"00",
		X"90",X"32",X"E0",X"98",X"21",X"20",X"98",X"11",X"60",X"98",X"06",X"40",X"4E",X"1A",X"77",X"79",
		X"12",X"2C",X"1C",X"10",X"F7",X"21",X"00",X"88",X"11",X"B0",X"98",X"06",X"30",X"7E",X"4F",X"26",
		X"8B",X"7E",X"E6",X"7F",X"0D",X"20",X"0B",X"E6",X"78",X"4F",X"2C",X"7E",X"2D",X"E6",X"07",X"B1",
		X"F6",X"80",X"EB",X"4E",X"77",X"EB",X"CB",X"79",X"28",X"10",X"79",X"E6",X"78",X"C6",X"06",X"77",
		X"2C",X"79",X"E6",X"07",X"77",X"2D",X"3E",X"01",X"18",X"07",X"71",X"26",X"93",X"36",X"00",X"3E",
		X"80",X"26",X"88",X"77",X"13",X"2C",X"2C",X"10",X"C4",X"21",X"00",X"90",X"11",X"E0",X"98",X"06",
		X"20",X"4E",X"1A",X"77",X"79",X"12",X"2C",X"1C",X"10",X"F7",X"AF",X"32",X"00",X"90",X"C9",X"21",
		X"02",X"80",X"06",X"12",X"7E",X"FE",X"4A",X"30",X"02",X"36",X"24",X"2C",X"10",X"F6",X"2E",X"22",
		X"06",X"12",X"7E",X"FE",X"4A",X"30",X"02",X"36",X"24",X"2C",X"10",X"F6",X"3A",X"21",X"98",X"06",
		X"00",X"21",X"01",X"80",X"FE",X"32",X"38",X"07",X"D6",X"32",X"04",X"2C",X"2C",X"18",X"F5",X"EB",
		X"6F",X"26",X"00",X"3E",X"0A",X"CD",X"61",X"10",X"67",X"E5",X"EB",X"FE",X"05",X"38",X"02",X"D6",
		X"04",X"4F",X"7B",X"CB",X"47",X"28",X"02",X"3E",X"02",X"81",X"D7",X"04",X"10",X"20",X"C1",X"79",
		X"CD",X"F5",X"11",X"78",X"FE",X"05",X"38",X"08",X"16",X"38",X"CD",X"13",X"12",X"78",X"D6",X"05",
		X"47",X"04",X"10",X"03",X"C3",X"7E",X"13",X"16",X"36",X"CD",X"13",X"12",X"18",X"F4",X"3E",X"04",
		X"CD",X"FB",X"11",X"18",X"D7",X"A7",X"C8",X"FE",X"04",X"28",X"07",X"07",X"07",X"C6",X"36",X"57",
		X"18",X"0A",X"16",X"42",X"CD",X"13",X"12",X"CD",X"28",X"12",X"16",X"3A",X"CD",X"13",X"12",X"CD",
		X"28",X"12",X"C9",X"08",X"38",X"11",X"08",X"3A",X"A0",X"92",X"C6",X"08",X"5F",X"3A",X"A0",X"92",
		X"93",X"20",X"FA",X"08",X"32",X"B5",X"9A",X"08",X"72",X"14",X"CB",X"ED",X"72",X"14",X"CB",X"D4",
		X"7A",X"E6",X"0C",X"FE",X"08",X"3E",X"01",X"28",X"01",X"3C",X"77",X"CB",X"AD",X"77",X"CB",X"94",
		X"2D",X"C9",X"21",X"5B",X"12",X"11",X"00",X"90",X"01",X"20",X"00",X"C5",X"E5",X"ED",X"B0",X"E1",
		X"C1",X"11",X"E0",X"98",X"ED",X"B0",X"AF",X"32",X"00",X"90",X"C9",X"1F",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"21",X"64",X"8B",X"11",X"30",
		X"09",X"0E",X"00",X"06",X"0A",X"73",X"26",X"93",X"36",X"00",X"26",X"9B",X"71",X"26",X"8B",X"2C",
		X"72",X"2C",X"78",X"FE",X"09",X"20",X"04",X"0E",X"01",X"16",X"0B",X"10",X"E8",X"C9",X"26",X"8B",
		X"ED",X"5B",X"80",X"92",X"1A",X"6F",X"13",X"1A",X"4F",X"E6",X"78",X"C6",X"06",X"77",X"2C",X"79",
		X"E6",X"07",X"CB",X"79",X"28",X"02",X"F6",X"08",X"77",X"13",X"2D",X"26",X"88",X"36",X"01",X"26",
		X"93",X"1A",X"77",X"13",X"2C",X"1A",X"CB",X"27",X"77",X"3E",X"00",X"17",X"26",X"9B",X"77",X"13",
		X"ED",X"53",X"80",X"92",X"C9",X"DD",X"6F",X"3A",X"15",X"92",X"4F",X"21",X"00",X"99",X"11",X"21",
		X"13",X"06",X"10",X"36",X"00",X"2C",X"1A",X"13",X"77",X"2C",X"10",X"F7",X"21",X"00",X"98",X"11",
		X"21",X"13",X"06",X"0A",X"1A",X"13",X"CB",X"41",X"28",X"03",X"C6",X"0D",X"2F",X"77",X"2C",X"2C",
		X"10",X"F2",X"06",X"06",X"1A",X"DD",X"85",X"13",X"CB",X"41",X"20",X"03",X"C6",X"4F",X"2F",X"CB",
		X"27",X"77",X"2C",X"3E",X"00",X"17",X"77",X"2C",X"10",X"EA",X"3A",X"15",X"92",X"32",X"0F",X"92",
		X"C9",X"31",X"41",X"51",X"61",X"71",X"81",X"91",X"A1",X"B1",X"C1",X"92",X"8A",X"82",X"7C",X"76",
		X"70",X"E5",X"21",X"AF",X"92",X"36",X"03",X"7E",X"A7",X"20",X"FC",X"E1",X"C9",X"3E",X"01",X"32",
		X"14",X"90",X"3A",X"70",X"82",X"FE",X"24",X"20",X"03",X"0E",X"03",X"F7",X"3A",X"87",X"92",X"A7",
		X"20",X"FA",X"CD",X"7E",X"13",X"21",X"06",X"09",X"22",X"62",X"8B",X"21",X"62",X"93",X"3A",X"15",
		X"92",X"E6",X"01",X"3E",X"29",X"0E",X"01",X"28",X"03",X"C6",X"0E",X"0D",X"36",X"7A",X"2C",X"77",
		X"26",X"9B",X"71",X"2D",X"AF",X"77",X"32",X"13",X"92",X"3C",X"32",X"B9",X"99",X"C9",X"3A",X"20",
		X"98",X"2F",X"C6",X"09",X"5F",X"16",X"49",X"21",X"1D",X"80",X"CD",X"98",X"13",X"2D",X"CD",X"98",
		X"13",X"CB",X"ED",X"2C",X"CD",X"98",X"13",X"2D",X"E5",X"14",X"4A",X"06",X"08",X"78",X"BB",X"20",
		X"02",X"0E",X"24",X"7E",X"FE",X"36",X"38",X"04",X"FE",X"4A",X"38",X"01",X"71",X"2D",X"2D",X"10",
		X"EC",X"E1",X"C9",X"A7",X"08",X"D5",X"EB",X"79",X"21",X"EF",X"13",X"CF",X"7E",X"23",X"66",X"6F",
		X"08",X"30",X"06",X"2B",X"2B",X"5E",X"23",X"56",X"23",X"4E",X"23",X"EB",X"1A",X"FE",X"2F",X"28",
		X"1E",X"D6",X"30",X"30",X"04",X"3E",X"24",X"18",X"06",X"FE",X"11",X"38",X"02",X"D6",X"07",X"77",
		X"CB",X"D4",X"71",X"CB",X"94",X"13",X"7D",X"D6",X"20",X"6F",X"30",X"E0",X"25",X"18",X"DD",X"D1",
		X"C9",X"2F",X"14",X"44",X"14",X"51",X"14",X"5C",X"14",X"66",X"14",X"72",X"14",X"7C",X"14",X"91",
		X"14",X"A3",X"14",X"AE",X"14",X"C2",X"14",X"E1",X"14",X"EE",X"14",X"09",X"15",X"13",X"15",X"22",
		X"15",X"2F",X"15",X"3C",X"15",X"40",X"15",X"59",X"15",X"5D",X"15",X"6A",X"15",X"81",X"15",X"8F",
		X"15",X"A8",X"15",X"BF",X"15",X"C5",X"15",X"D9",X"15",X"ED",X"15",X"FF",X"15",X"EB",X"82",X"00",
		X"50",X"55",X"53",X"48",X"20",X"53",X"54",X"41",X"52",X"54",X"20",X"42",X"55",X"54",X"54",X"4F",
		X"4E",X"2F",X"70",X"82",X"00",X"47",X"41",X"4D",X"45",X"20",X"4F",X"56",X"45",X"52",X"2F",X"70",
		X"82",X"00",X"52",X"45",X"41",X"44",X"59",X"20",X"21",X"2F",X"50",X"82",X"00",X"50",X"4C",X"41",
		X"59",X"45",X"52",X"20",X"31",X"2F",X"00",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"32",X"2F",
		X"70",X"82",X"00",X"53",X"54",X"41",X"47",X"45",X"20",X"2F",X"10",X"83",X"00",X"43",X"48",X"41",
		X"4C",X"4C",X"45",X"4E",X"47",X"49",X"4E",X"47",X"20",X"53",X"54",X"41",X"47",X"45",X"2F",X"10",
		X"83",X"00",X"4E",X"55",X"4D",X"42",X"45",X"52",X"20",X"4F",X"46",X"20",X"48",X"49",X"54",X"53",
		X"2F",X"B3",X"82",X"00",X"42",X"4F",X"4E",X"55",X"53",X"20",X"20",X"2F",X"F1",X"82",X"04",X"46",
		X"49",X"47",X"48",X"54",X"45",X"52",X"20",X"43",X"41",X"50",X"54",X"55",X"52",X"45",X"44",X"2F",
		X"AD",X"83",X"00",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"2F",X"6D",
		X"82",X"04",X"50",X"45",X"52",X"46",X"45",X"43",X"54",X"20",X"63",X"2F",X"73",X"83",X"05",X"53",
		X"50",X"45",X"43",X"49",X"41",X"4C",X"20",X"42",X"4F",X"4E",X"55",X"53",X"20",X"31",X"30",X"30",
		X"30",X"30",X"20",X"50",X"54",X"53",X"2F",X"42",X"82",X"00",X"47",X"41",X"4C",X"41",X"47",X"41",
		X"2F",X"A5",X"82",X"00",X"5D",X"5D",X"20",X"53",X"43",X"4F",X"52",X"45",X"20",X"5D",X"5D",X"2F",
		X"28",X"82",X"00",X"35",X"30",X"20",X"20",X"20",X"20",X"31",X"30",X"30",X"2F",X"2A",X"82",X"00",
		X"38",X"30",X"20",X"20",X"20",X"20",X"31",X"36",X"30",X"2F",X"2B",X"82",X"00",X"2F",X"3B",X"83",
		X"03",X"65",X"20",X"31",X"39",X"38",X"31",X"20",X"4D",X"49",X"44",X"57",X"41",X"59",X"20",X"4D",
		X"46",X"47",X"61",X"43",X"4F",X"61",X"2F",X"5E",X"82",X"04",X"2F",X"8F",X"82",X"04",X"5D",X"52",
		X"45",X"53",X"55",X"4C",X"54",X"53",X"5D",X"2F",X"32",X"83",X"05",X"53",X"48",X"4F",X"54",X"53",
		X"20",X"46",X"49",X"52",X"45",X"44",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"2F",X"05",X"20",X"20",X"4D",X"49",X"53",X"53",X"49",X"4C",X"45",X"53",X"2F",X"35",X"83",X"05",
		X"4E",X"55",X"4D",X"42",X"45",X"52",X"20",X"4F",X"46",X"20",X"48",X"49",X"54",X"53",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"2F",X"38",X"83",X"03",X"48",X"49",X"54",X"5D",X"4D",X"49",X"53",
		X"53",X"20",X"52",X"41",X"54",X"49",X"4F",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"2F",X"03",
		X"24",X"60",X"2F",X"2F",X"83",X"05",X"31",X"53",X"54",X"20",X"42",X"4F",X"4E",X"55",X"53",X"20",
		X"46",X"4F",X"52",X"20",X"20",X"20",X"2F",X"32",X"83",X"05",X"32",X"4E",X"44",X"20",X"42",X"4F",
		X"4E",X"55",X"53",X"20",X"46",X"4F",X"52",X"20",X"20",X"20",X"2F",X"35",X"83",X"05",X"41",X"4E",
		X"44",X"20",X"46",X"4F",X"52",X"20",X"45",X"56",X"45",X"52",X"59",X"20",X"20",X"20",X"2F",X"05",
		X"30",X"30",X"30",X"30",X"20",X"50",X"54",X"53",X"2F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"ED",X"5B",X"82",X"92",X"1A",X"07",X"07",X"07",X"E6",X"07",X"21",X"13",X"17",X"CF",X"7E",X"23",
		X"66",X"6F",X"E9",X"66",X"17",X"66",X"17",X"1F",X"17",X"66",X"17",X"34",X"17",X"2D",X"17",X"3A",
		X"A0",X"92",X"E6",X"0F",X"C0",X"21",X"07",X"92",X"35",X"C0",X"C3",X"66",X"17",X"CD",X"15",X"1F",
		X"ED",X"5B",X"82",X"92",X"1A",X"21",X"27",X"98",X"5E",X"CB",X"47",X"20",X"04",X"E6",X"0A",X"18",
		X"14",X"3A",X"09",X"92",X"6F",X"26",X"93",X"3A",X"62",X"93",X"96",X"3E",X"0A",X"28",X"06",X"3E",
		X"08",X"38",X"02",X"3E",X"02",X"CD",X"98",X"1F",X"3A",X"A0",X"92",X"E6",X"03",X"C0",X"21",X"07",
		X"92",X"35",X"C0",X"CD",X"15",X"1F",X"ED",X"5B",X"82",X"92",X"1A",X"E6",X"C0",X"FE",X"80",X"20",
		X"01",X"13",X"13",X"1A",X"ED",X"53",X"82",X"92",X"07",X"07",X"07",X"E6",X"07",X"21",X"86",X"17",
		X"CF",X"7E",X"23",X"66",X"6F",X"E9",X"94",X"17",X"94",X"17",X"A1",X"17",X"A8",X"17",X"AE",X"17",
		X"AE",X"17",X"9C",X"17",X"1A",X"07",X"E6",X"7E",X"32",X"09",X"92",X"C9",X"AF",X"32",X"03",X"90",
		X"C9",X"1A",X"E6",X"1F",X"32",X"07",X"92",X"C9",X"1A",X"E6",X"1F",X"4F",X"F7",X"C9",X"13",X"1A",
		X"18",X"F2",X"3A",X"01",X"92",X"3D",X"C0",X"3A",X"03",X"92",X"21",X"C3",X"17",X"CF",X"5E",X"23",
		X"56",X"EB",X"E9",X"40",X"19",X"48",X"19",X"84",X"19",X"D9",X"18",X"D1",X"18",X"AC",X"18",X"40",
		X"19",X"F5",X"17",X"52",X"18",X"D1",X"18",X"08",X"18",X"D1",X"18",X"40",X"18",X"40",X"19",X"E1",
		X"17",X"3A",X"AF",X"92",X"A7",X"28",X"05",X"3D",X"CA",X"A7",X"19",X"C9",X"CD",X"14",X"32",X"3E",
		X"0A",X"32",X"AF",X"92",X"C9",X"3A",X"A0",X"92",X"E6",X"1F",X"FE",X"1F",X"C0",X"3E",X"01",X"32",
		X"05",X"90",X"0E",X"02",X"F7",X"C3",X"A7",X"19",X"CD",X"4C",X"13",X"21",X"1F",X"18",X"22",X"82",
		X"92",X"3E",X"01",X"32",X"03",X"90",X"32",X"15",X"90",X"32",X"25",X"90",X"C3",X"A7",X"19",X"08",
		X"18",X"8A",X"08",X"88",X"06",X"81",X"28",X"81",X"05",X"54",X"1A",X"88",X"12",X"81",X"0F",X"A2",
		X"16",X"AA",X"14",X"88",X"18",X"88",X"10",X"43",X"82",X"10",X"88",X"06",X"A2",X"20",X"56",X"C0",
		X"EF",X"CD",X"42",X"12",X"AF",X"32",X"10",X"90",X"32",X"0B",X"92",X"3C",X"32",X"02",X"90",X"C3",
		X"A7",X"19",X"AF",X"32",X"2B",X"98",X"3C",X"32",X"B7",X"9A",X"32",X"21",X"98",X"32",X"03",X"90",
		X"32",X"15",X"90",X"32",X"25",X"98",X"21",X"87",X"18",X"22",X"82",X"92",X"CD",X"C5",X"01",X"CD",
		X"4C",X"13",X"3E",X"01",X"32",X"0B",X"92",X"32",X"42",X"98",X"32",X"2C",X"98",X"3C",X"32",X"C4",
		X"99",X"32",X"C5",X"99",X"C3",X"A7",X"19",X"02",X"8A",X"04",X"82",X"07",X"AA",X"28",X"88",X"10",
		X"AA",X"38",X"82",X"12",X"AA",X"20",X"88",X"14",X"AA",X"20",X"82",X"06",X"A8",X"0E",X"A2",X"17",
		X"88",X"12",X"A2",X"14",X"18",X"88",X"1B",X"81",X"2A",X"5F",X"4C",X"C0",X"3A",X"AE",X"92",X"A7",
		X"28",X"09",X"3D",X"CA",X"A7",X"19",X"FE",X"05",X"28",X"0C",X"C9",X"3E",X"34",X"32",X"34",X"92",
		X"3E",X"09",X"32",X"AE",X"92",X"C9",X"AF",X"32",X"62",X"93",X"0E",X"13",X"F7",X"0E",X"14",X"F7",
		X"C9",X"3A",X"03",X"90",X"A7",X"CA",X"A7",X"19",X"C9",X"06",X"07",X"CD",X"9E",X"12",X"10",X"FB",
		X"AF",X"32",X"20",X"98",X"32",X"05",X"90",X"CD",X"4C",X"13",X"21",X"0D",X"FF",X"22",X"C5",X"92",
		X"22",X"C4",X"92",X"22",X"C1",X"92",X"22",X"C0",X"92",X"21",X"28",X"19",X"22",X"82",X"92",X"AF",
		X"06",X"10",X"21",X"CA",X"92",X"DF",X"32",X"27",X"98",X"32",X"0B",X"92",X"3C",X"32",X"2B",X"98",
		X"32",X"10",X"90",X"32",X"0B",X"90",X"32",X"03",X"90",X"3A",X"03",X"68",X"0F",X"E6",X"01",X"32",
		X"B7",X"9A",X"CD",X"7B",X"12",X"C3",X"A7",X"19",X"08",X"1B",X"81",X"3D",X"81",X"0A",X"42",X"19",
		X"81",X"28",X"81",X"08",X"18",X"81",X"2E",X"81",X"03",X"1A",X"81",X"11",X"81",X"05",X"42",X"C0",
		X"CD",X"60",X"01",X"CD",X"3C",X"00",X"18",X"5F",X"21",X"5C",X"19",X"22",X"80",X"92",X"AF",X"32",
		X"05",X"92",X"32",X"A8",X"92",X"3E",X"02",X"32",X"AE",X"92",X"18",X"4B",X"08",X"1B",X"44",X"3A",
		X"0A",X"12",X"44",X"42",X"0C",X"08",X"7C",X"50",X"34",X"08",X"34",X"5C",X"30",X"08",X"64",X"5C",
		X"32",X"08",X"94",X"5C",X"4A",X"12",X"A4",X"64",X"36",X"08",X"C4",X"5C",X"58",X"12",X"B4",X"64",
		X"52",X"12",X"D4",X"64",X"3A",X"AE",X"92",X"A7",X"C0",X"3E",X"02",X"32",X"AE",X"92",X"3A",X"05",
		X"92",X"FE",X"05",X"28",X"12",X"3C",X"32",X"05",X"92",X"C6",X"0D",X"4F",X"F7",X"3A",X"05",X"92",
		X"FE",X"03",X"D8",X"CD",X"9E",X"12",X"C9",X"21",X"03",X"92",X"34",X"7E",X"FE",X"0F",X"C0",X"36",
		X"00",X"C9",X"3A",X"8E",X"92",X"A7",X"20",X"1A",X"21",X"AD",X"92",X"B6",X"28",X"28",X"FE",X"04",
		X"20",X"05",X"3D",X"77",X"32",X"A9",X"9A",X"3A",X"29",X"98",X"C6",X"0D",X"6F",X"26",X"91",X"36",
		X"04",X"C9",X"0E",X"0A",X"F7",X"3E",X"06",X"32",X"AD",X"92",X"3C",X"32",X"63",X"8B",X"AF",X"32",
		X"8B",X"92",X"32",X"8E",X"92",X"C9",X"3A",X"D1",X"82",X"FE",X"24",X"28",X"29",X"21",X"62",X"93",
		X"3A",X"28",X"98",X"E6",X"07",X"5F",X"54",X"7E",X"12",X"36",X"00",X"2C",X"1C",X"7E",X"12",X"26",
		X"9B",X"54",X"ED",X"A8",X"ED",X"A0",X"26",X"8B",X"6B",X"36",X"07",X"2D",X"36",X"07",X"0E",X"0B",
		X"21",X"B1",X"83",X"CD",X"B3",X"13",X"3A",X"28",X"98",X"6F",X"E6",X"07",X"5F",X"26",X"88",X"3A",
		X"15",X"92",X"4F",X"7E",X"FE",X"09",X"20",X"1D",X"26",X"93",X"54",X"7E",X"12",X"2C",X"1C",X"3E",
		X"10",X"CB",X"41",X"28",X"02",X"ED",X"44",X"47",X"86",X"12",X"1F",X"A8",X"07",X"E6",X"01",X"26",
		X"9B",X"54",X"AE",X"12",X"C9",X"21",X"8B",X"92",X"7E",X"A7",X"20",X"05",X"16",X"8B",X"3E",X"06",
		X"12",X"34",X"FE",X"24",X"28",X"1A",X"06",X"01",X"CB",X"41",X"20",X"02",X"05",X"05",X"6B",X"2C",
		X"26",X"93",X"78",X"86",X"77",X"1F",X"A8",X"07",X"D0",X"26",X"9B",X"7E",X"EE",X"01",X"77",X"C9",
		X"AF",X"32",X"11",X"90",X"32",X"A9",X"9A",X"16",X"88",X"3C",X"12",X"32",X"28",X"98",X"32",X"B9",
		X"99",X"3C",X"32",X"13",X"92",X"C9",X"3A",X"CA",X"99",X"4F",X"3A",X"A7",X"92",X"B9",X"D0",X"3A",
		X"41",X"98",X"A7",X"20",X"46",X"21",X"07",X"88",X"01",X"FF",X"14",X"3E",X"01",X"2C",X"ED",X"A1",
		X"28",X"0F",X"10",X"F9",X"21",X"3F",X"88",X"06",X"10",X"2C",X"ED",X"A1",X"28",X"03",X"10",X"F9",
		X"C9",X"3E",X"C0",X"32",X"41",X"98",X"2D",X"5D",X"16",X"8B",X"1C",X"1A",X"1D",X"4F",X"3A",X"21",
		X"98",X"CB",X"3F",X"CB",X"3F",X"6F",X"26",X"00",X"3E",X"03",X"CD",X"61",X"10",X"C6",X"04",X"21",
		X"2D",X"98",X"73",X"2C",X"71",X"2C",X"77",X"32",X"B2",X"9A",X"C9",X"3C",X"28",X"1C",X"32",X"41",
		X"98",X"08",X"21",X"2D",X"98",X"5E",X"16",X"88",X"1A",X"3D",X"C2",X"5A",X"1B",X"16",X"8B",X"2C",
		X"08",X"CB",X"67",X"28",X"01",X"2C",X"7E",X"1C",X"12",X"C9",X"3A",X"15",X"90",X"A7",X"20",X"06",
		X"3E",X"E0",X"32",X"41",X"98",X"C9",X"3A",X"2D",X"98",X"6F",X"26",X"88",X"7E",X"3D",X"20",X"4A",
		X"26",X"92",X"7E",X"CB",X"7F",X"20",X"43",X"3A",X"2F",X"98",X"D6",X"04",X"21",X"5F",X"1B",X"CF",
		X"11",X"B0",X"99",X"3E",X"03",X"12",X"1C",X"ED",X"A0",X"ED",X"A0",X"3A",X"2F",X"98",X"D6",X"04",
		X"E6",X"0F",X"4F",X"21",X"65",X"1B",X"CF",X"5E",X"23",X"56",X"26",X"8B",X"3A",X"2D",X"98",X"6F",
		X"79",X"07",X"07",X"07",X"C6",X"56",X"4E",X"77",X"79",X"E6",X"F8",X"4F",X"3A",X"2E",X"98",X"E6",
		X"07",X"B1",X"32",X"2E",X"98",X"26",X"88",X"CD",X"83",X"10",X"AF",X"32",X"04",X"90",X"C9",X"1E",
		X"BD",X"0A",X"B8",X"14",X"BC",X"EA",X"04",X"73",X"04",X"AB",X"04",X"3A",X"0B",X"92",X"A7",X"28",
		X"0A",X"3A",X"15",X"90",X"4F",X"3A",X"1D",X"90",X"2F",X"A1",X"C8",X"06",X"04",X"21",X"CA",X"92",
		X"7E",X"3C",X"20",X"0D",X"2C",X"2C",X"2C",X"10",X"F7",X"3A",X"A0",X"92",X"E6",X"0F",X"28",X"1E",
		X"C9",X"36",X"FF",X"3D",X"16",X"88",X"5F",X"CB",X"BB",X"08",X"1A",X"3D",X"C0",X"2C",X"5E",X"2C",
		X"56",X"08",X"6F",X"26",X"88",X"CD",X"79",X"10",X"3E",X"01",X"32",X"B3",X"9A",X"C9",X"21",X"C0",
		X"92",X"06",X"03",X"35",X"28",X"04",X"2C",X"10",X"FA",X"C9",X"3A",X"C4",X"99",X"4F",X"3A",X"87",
		X"92",X"B9",X"38",X"02",X"34",X"C9",X"CB",X"D5",X"7E",X"CB",X"95",X"77",X"78",X"3D",X"21",X"D7",
		X"1B",X"CF",X"7E",X"23",X"66",X"6F",X"E9",X"DD",X"1B",X"FD",X"1B",X"07",X"1C",X"06",X"14",X"21",
		X"08",X"88",X"11",X"4F",X"03",X"3A",X"2D",X"98",X"4F",X"7E",X"3D",X"20",X"04",X"79",X"BD",X"20",
		X"05",X"2C",X"2C",X"10",X"F4",X"C9",X"32",X"B3",X"9A",X"CD",X"83",X"10",X"C9",X"06",X"10",X"21",
		X"40",X"88",X"11",X"A9",X"03",X"18",X"DE",X"3A",X"2B",X"98",X"A7",X"20",X"29",X"21",X"2C",X"98",
		X"34",X"CB",X"46",X"20",X"21",X"DD",X"2E",X"02",X"FD",X"21",X"54",X"04",X"11",X"30",X"88",X"06",
		X"04",X"1A",X"3D",X"28",X"05",X"1C",X"1C",X"10",X"F8",X"C9",X"3E",X"01",X"32",X"2B",X"98",X"7B",
		X"32",X"28",X"98",X"C3",X"B4",X"1C",X"21",X"32",X"1D",X"16",X"88",X"01",X"00",X"06",X"5E",X"23",
		X"3A",X"2D",X"98",X"BB",X"28",X"04",X"1A",X"3D",X"D6",X"01",X"CB",X"11",X"10",X"F0",X"DD",X"2E",
		X"00",X"06",X"04",X"DD",X"61",X"79",X"E6",X"07",X"FE",X"04",X"28",X"05",X"FE",X"03",X"D4",X"93",
		X"1C",X"CB",X"19",X"10",X"F0",X"DD",X"2C",X"DD",X"4C",X"06",X"04",X"79",X"E6",X"07",X"C4",X"93",
		X"1C",X"CB",X"19",X"10",X"F6",X"DD",X"2C",X"11",X"30",X"88",X"06",X"04",X"1A",X"3D",X"28",X"26",
		X"1C",X"1C",X"10",X"F8",X"21",X"00",X"88",X"06",X"04",X"7E",X"3D",X"CA",X"2B",X"1D",X"2C",X"2C",
		X"10",X"F7",X"C9",X"78",X"CB",X"4F",X"28",X"02",X"EE",X"01",X"E6",X"03",X"CB",X"27",X"C6",X"30",
		X"5F",X"1A",X"FE",X"01",X"C0",X"E1",X"FD",X"21",X"11",X"04",X"3A",X"0B",X"92",X"A7",X"20",X"04",
		X"FD",X"21",X"F1",X"00",X"7B",X"0F",X"0F",X"7B",X"17",X"0F",X"32",X"CA",X"92",X"08",X"FD",X"22",
		X"CB",X"92",X"04",X"7B",X"E6",X"07",X"21",X"30",X"98",X"D7",X"DD",X"7D",X"EB",X"21",X"03",X"1D",
		X"CF",X"7E",X"12",X"23",X"1C",X"7E",X"12",X"DD",X"7D",X"FE",X"02",X"28",X"0C",X"11",X"CD",X"92",
		X"3D",X"28",X"03",X"CD",X"09",X"1D",X"CD",X"09",X"1D",X"3A",X"CA",X"92",X"E6",X"07",X"6F",X"26",
		X"88",X"7E",X"3D",X"C0",X"4D",X"21",X"CA",X"92",X"2C",X"2C",X"2C",X"7E",X"3C",X"20",X"F9",X"08",
		X"79",X"18",X"19",X"0D",X"BA",X"05",X"B7",X"01",X"B5",X"CB",X"09",X"38",X"06",X"05",X"CB",X"09",
		X"38",X"01",X"05",X"78",X"05",X"21",X"32",X"1D",X"D7",X"08",X"7E",X"EB",X"17",X"0F",X"77",X"08",
		X"2C",X"FD",X"7D",X"77",X"2C",X"FD",X"7C",X"77",X"2C",X"EB",X"C9",X"11",X"44",X"04",X"CD",X"83",
		X"10",X"C9",X"4A",X"52",X"5A",X"58",X"50",X"48",X"21",X"B4",X"99",X"7E",X"E6",X"7F",X"D6",X"7E",
		X"28",X"36",X"4E",X"34",X"3A",X"15",X"92",X"CB",X"01",X"A9",X"0F",X"3E",X"01",X"38",X"02",X"ED",
		X"44",X"4F",X"21",X"14",X"98",X"06",X"06",X"7E",X"81",X"77",X"1F",X"A9",X"2C",X"07",X"30",X"04",
		X"7E",X"EE",X"01",X"77",X"2C",X"10",X"F0",X"3A",X"A0",X"92",X"E6",X"FC",X"3C",X"F5",X"CD",X"EE",
		X"23",X"F1",X"C6",X"02",X"CD",X"EE",X"23",X"C9",X"32",X"0E",X"90",X"C9",X"3A",X"15",X"92",X"47",
		X"21",X"B9",X"99",X"7E",X"2C",X"A7",X"28",X"26",X"7E",X"A7",X"3E",X"FD",X"20",X"13",X"2C",X"7E",
		X"2C",X"BE",X"28",X"01",X"34",X"7E",X"2C",X"86",X"4F",X"E6",X"3F",X"77",X"79",X"07",X"07",X"E6",
		X"03",X"CB",X"40",X"20",X"02",X"ED",X"44",X"3D",X"E6",X"07",X"32",X"BE",X"99",X"C9",X"AF",X"77",
		X"2C",X"2C",X"77",X"2C",X"77",X"3E",X"07",X"18",X"F1",X"21",X"00",X"92",X"06",X"30",X"CB",X"7E",
		X"20",X"05",X"2C",X"2C",X"10",X"F8",X"C9",X"CB",X"BE",X"26",X"88",X"36",X"04",X"2C",X"36",X"40",
		X"26",X"8B",X"36",X"0A",X"26",X"92",X"18",X"EB",X"3A",X"A2",X"92",X"E6",X"01",X"C0",X"21",X"AC",
		X"92",X"06",X"04",X"7E",X"A7",X"28",X"01",X"35",X"2C",X"10",X"F8",X"C9",X"3A",X"A0",X"92",X"E6",
		X"03",X"C0",X"21",X"0F",X"92",X"7E",X"5F",X"16",X"FF",X"CB",X"7F",X"20",X"05",X"14",X"14",X"34",
		X"18",X"01",X"35",X"FE",X"1F",X"20",X"02",X"CB",X"FE",X"FE",X"81",X"20",X"02",X"CB",X"BE",X"4E",
		X"E6",X"07",X"7A",X"32",X"11",X"92",X"7B",X"20",X"10",X"21",X"6A",X"1E",X"79",X"E6",X"18",X"CF",
		X"7B",X"11",X"20",X"99",X"01",X"10",X"00",X"ED",X"B0",X"21",X"15",X"92",X"07",X"AE",X"0F",X"21",
		X"20",X"99",X"11",X"00",X"99",X"30",X"05",X"01",X"FF",X"01",X"18",X"03",X"01",X"01",X"FF",X"DD",
		X"2E",X"05",X"CD",X"49",X"1E",X"41",X"DD",X"2E",X"0B",X"CB",X"0E",X"30",X"15",X"1A",X"80",X"12",
		X"16",X"98",X"1A",X"80",X"12",X"1F",X"A8",X"07",X"30",X"06",X"1C",X"1A",X"EE",X"01",X"12",X"1D",
		X"16",X"99",X"1C",X"1C",X"2C",X"DD",X"2D",X"20",X"E0",X"C9",X"FF",X"77",X"55",X"14",X"10",X"10",
		X"14",X"55",X"77",X"FF",X"00",X"10",X"14",X"55",X"77",X"FF",X"FF",X"77",X"55",X"51",X"10",X"10",
		X"51",X"55",X"77",X"FF",X"00",X"10",X"51",X"55",X"77",X"FF",X"FF",X"77",X"57",X"15",X"10",X"10",
		X"15",X"57",X"77",X"FF",X"00",X"10",X"15",X"57",X"77",X"FF",X"FF",X"F7",X"D5",X"91",X"10",X"10",
		X"91",X"D5",X"F7",X"FF",X"00",X"10",X"91",X"D5",X"F7",X"FF",X"3A",X"A0",X"92",X"E6",X"01",X"C6",
		X"02",X"47",X"3A",X"15",X"92",X"A7",X"78",X"28",X"02",X"ED",X"44",X"DD",X"67",X"2E",X"68",X"11",
		X"B0",X"92",X"DD",X"2E",X"08",X"26",X"8B",X"7E",X"FE",X"30",X"20",X"39",X"26",X"93",X"7E",X"A7",
		X"28",X"33",X"EB",X"46",X"78",X"E6",X"7E",X"2C",X"86",X"4F",X"E6",X"1F",X"77",X"2C",X"79",X"07",
		X"07",X"07",X"E6",X"07",X"CB",X"78",X"28",X"02",X"ED",X"44",X"EB",X"86",X"77",X"2C",X"7E",X"DD",
		X"84",X"77",X"1F",X"DD",X"AC",X"07",X"30",X"07",X"26",X"9B",X"CB",X"0E",X"3F",X"CB",X"16",X"2C",
		X"DD",X"2D",X"20",X"C1",X"C9",X"2C",X"1C",X"1C",X"18",X"F5",X"3A",X"15",X"92",X"C6",X"B6",X"6F",
		X"26",X"99",X"CB",X"66",X"C0",X"21",X"64",X"93",X"11",X"A4",X"92",X"AF",X"BE",X"28",X"05",X"2E",
		X"66",X"1C",X"BE",X"C0",X"D5",X"EB",X"21",X"63",X"9B",X"54",X"1C",X"CB",X"56",X"28",X"02",X"D1",
		X"C9",X"ED",X"A8",X"26",X"93",X"54",X"ED",X"A0",X"ED",X"A8",X"26",X"9B",X"54",X"46",X"EB",X"3A",
		X"27",X"98",X"E6",X"01",X"07",X"07",X"07",X"B0",X"77",X"16",X"8B",X"1A",X"62",X"E6",X"07",X"0E",
		X"30",X"FE",X"05",X"30",X"07",X"0C",X"FE",X"02",X"30",X"02",X"0C",X"0C",X"71",X"FE",X"04",X"38",
		X"03",X"2F",X"C6",X"47",X"CB",X"27",X"4F",X"78",X"0F",X"0F",X"0F",X"E6",X"60",X"47",X"3A",X"15",
		X"92",X"A7",X"78",X"20",X"02",X"EE",X"60",X"B1",X"D1",X"12",X"26",X"88",X"36",X"06",X"3E",X"01",
		X"32",X"AF",X"9A",X"2A",X"46",X"98",X"23",X"22",X"46",X"98",X"C9",X"3A",X"27",X"98",X"5F",X"3A",
		X"15",X"92",X"C6",X"B6",X"6F",X"26",X"99",X"7E",X"E6",X"0A",X"FE",X"0A",X"28",X"37",X"21",X"15",
		X"92",X"CB",X"46",X"28",X"02",X"EE",X"0A",X"21",X"A3",X"92",X"47",X"0E",X"01",X"7E",X"EE",X"01",
		X"77",X"20",X"01",X"0C",X"21",X"62",X"93",X"7E",X"A7",X"C8",X"CB",X"48",X"20",X"0F",X"7E",X"FE",
		X"D1",X"38",X"03",X"CB",X"43",X"C0",X"FE",X"E1",X"D0",X"81",X"77",X"18",X"0D",X"7E",X"FE",X"12",
		X"D8",X"91",X"77",X"18",X"05",X"AF",X"32",X"A3",X"92",X"C9",X"CB",X"43",X"C8",X"C6",X"0F",X"32",
		X"60",X"93",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",
		X"3A",X"28",X"98",X"6F",X"26",X"88",X"7E",X"A7",X"C2",X"BF",X"20",X"3A",X"8B",X"92",X"A7",X"CA",
		X"C7",X"20",X"3D",X"CA",X"D1",X"20",X"26",X"93",X"7E",X"FE",X"80",X"28",X"09",X"F2",X"23",X"20",
		X"34",X"18",X"3B",X"35",X"18",X"38",X"2C",X"3A",X"15",X"92",X"A7",X"20",X"1F",X"7E",X"FE",X"29",
		X"20",X"0F",X"26",X"9B",X"7E",X"26",X"93",X"3D",X"20",X"07",X"3E",X"03",X"32",X"8B",X"92",X"18",
		X"1D",X"34",X"20",X"1A",X"26",X"9B",X"7E",X"EE",X"01",X"77",X"18",X"12",X"7E",X"FE",X"37",X"20",
		X"08",X"26",X"9B",X"7E",X"26",X"93",X"A7",X"28",X"E1",X"35",X"7E",X"3C",X"28",X"E6",X"21",X"62",
		X"8B",X"7E",X"D6",X"06",X"4F",X"26",X"93",X"20",X"0C",X"7E",X"FE",X"71",X"28",X"07",X"F2",X"73",
		X"20",X"34",X"C9",X"35",X"C9",X"3A",X"8B",X"92",X"FE",X"03",X"C0",X"3A",X"28",X"98",X"6F",X"36",
		X"00",X"2C",X"0D",X"0C",X"28",X"09",X"11",X"63",X"93",X"AF",X"32",X"2B",X"98",X"18",X"08",X"3E",
		X"01",X"32",X"27",X"98",X"11",X"61",X"93",X"7E",X"12",X"26",X"9B",X"54",X"7E",X"12",X"2D",X"26",
		X"88",X"36",X"80",X"26",X"8B",X"6B",X"2D",X"36",X"06",X"2C",X"36",X"09",X"2D",X"26",X"93",X"36",
		X"80",X"3E",X"01",X"32",X"14",X"90",X"32",X"15",X"90",X"32",X"25",X"90",X"32",X"B9",X"99",X"AF",
		X"32",X"1D",X"90",X"32",X"B1",X"9A",X"C9",X"3C",X"32",X"8B",X"92",X"3E",X"02",X"32",X"AD",X"92",
		X"C9",X"26",X"9B",X"3A",X"AD",X"92",X"5F",X"3A",X"87",X"92",X"B3",X"32",X"8D",X"92",X"CD",X"96",
		X"21",X"05",X"C0",X"32",X"14",X"90",X"32",X"15",X"90",X"32",X"25",X"90",X"3E",X"02",X"32",X"8B",
		X"92",X"C9",X"21",X"62",X"8B",X"7E",X"FE",X"40",X"38",X"08",X"AF",X"32",X"1C",X"90",X"32",X"BA",
		X"99",X"C9",X"26",X"9B",X"CD",X"96",X"21",X"CB",X"40",X"20",X"54",X"3A",X"8B",X"92",X"CB",X"7F",
		X"20",X"59",X"3A",X"8D",X"92",X"A7",X"C8",X"26",X"93",X"3A",X"28",X"98",X"5F",X"54",X"1A",X"BE",
		X"28",X"07",X"F2",X"28",X"21",X"35",X"18",X"01",X"34",X"2C",X"3A",X"15",X"92",X"A7",X"28",X"0B",
		X"34",X"7E",X"FE",X"7A",X"28",X"24",X"FE",X"80",X"28",X"16",X"C9",X"35",X"7E",X"3C",X"20",X"08",
		X"26",X"9B",X"7E",X"EE",X"01",X"77",X"26",X"93",X"7E",X"FE",X"E6",X"28",X"0D",X"FE",X"E0",X"C0",
		X"AF",X"32",X"8D",X"92",X"3E",X"07",X"32",X"63",X"8B",X"C9",X"AF",X"32",X"15",X"90",X"C9",X"3A",
		X"15",X"90",X"A7",X"20",X"06",X"3C",X"32",X"0D",X"92",X"18",X"22",X"26",X"93",X"2C",X"3A",X"15",
		X"92",X"A7",X"28",X"07",X"7E",X"FE",X"37",X"28",X"12",X"35",X"C9",X"7E",X"FE",X"29",X"28",X"0B",
		X"34",X"C0",X"26",X"9B",X"7E",X"EE",X"01",X"77",X"26",X"93",X"C9",X"05",X"C0",X"AF",X"32",X"1C",
		X"90",X"3C",X"32",X"25",X"90",X"C9",X"7E",X"4F",X"CB",X"3F",X"A9",X"4F",X"26",X"8B",X"06",X"00",
		X"7E",X"E6",X"07",X"FE",X"06",X"20",X"0E",X"0D",X"0C",X"20",X"0A",X"08",X"3A",X"8D",X"92",X"A7",
		X"20",X"02",X"04",X"C9",X"08",X"CB",X"41",X"20",X"07",X"FE",X"06",X"28",X"09",X"34",X"18",X"0E",
		X"A7",X"28",X"03",X"35",X"18",X"08",X"0D",X"F2",X"B5",X"21",X"0E",X"03",X"18",X"E7",X"79",X"CB",
		X"4F",X"28",X"02",X"EE",X"01",X"26",X"9B",X"77",X"C9",X"21",X"28",X"98",X"5E",X"16",X"88",X"1A",
		X"FE",X"09",X"20",X"44",X"2C",X"7E",X"DD",X"6F",X"DD",X"26",X"91",X"DD",X"7E",X"0A",X"A7",X"C0",
		X"3E",X"0C",X"DD",X"CB",X"05",X"46",X"28",X"02",X"ED",X"44",X"DD",X"77",X"0C",X"DD",X"7E",X"05",
		X"0F",X"DD",X"7E",X"04",X"1F",X"D6",X"78",X"FE",X"10",X"D0",X"3A",X"C6",X"99",X"32",X"2A",X"98",
		X"AF",X"DD",X"77",X"0C",X"32",X"19",X"90",X"32",X"8B",X"92",X"32",X"0D",X"92",X"3C",X"32",X"18",
		X"90",X"32",X"8C",X"92",X"32",X"8D",X"92",X"C9",X"AF",X"32",X"19",X"90",X"32",X"2B",X"98",X"C9",
		X"3A",X"A0",X"92",X"4F",X"E6",X"03",X"20",X"2D",X"3A",X"8A",X"92",X"ED",X"44",X"D6",X"18",X"26",
		X"21",X"07",X"CB",X"14",X"07",X"CB",X"14",X"E6",X"E0",X"C6",X"15",X"6F",X"79",X"0F",X"0F",X"E6",
		X"03",X"20",X"01",X"3C",X"C6",X"17",X"11",X"16",X"00",X"0E",X"06",X"06",X"0A",X"77",X"2C",X"10",
		X"FC",X"19",X"0D",X"20",X"F6",X"21",X"8B",X"92",X"CB",X"7E",X"20",X"0C",X"3A",X"28",X"98",X"5F",
		X"16",X"88",X"1A",X"FE",X"09",X"C2",X"35",X"23",X"21",X"8C",X"92",X"35",X"C2",X"4B",X"23",X"3A",
		X"2A",X"98",X"77",X"21",X"8B",X"92",X"CB",X"7E",X"20",X"2F",X"32",X"A5",X"9A",X"3A",X"29",X"98",
		X"C6",X"0D",X"5F",X"16",X"91",X"3E",X"FF",X"12",X"34",X"7E",X"E6",X"0F",X"FE",X"0B",X"28",X"40",
		X"CB",X"76",X"20",X"2B",X"F5",X"4F",X"07",X"81",X"21",X"A9",X"23",X"CF",X"F1",X"CD",X"98",X"23",
		X"06",X"06",X"7E",X"12",X"23",X"E7",X"10",X"FA",X"C9",X"34",X"7E",X"E6",X"0F",X"FE",X"0B",X"20",
		X"12",X"AF",X"32",X"18",X"90",X"32",X"A5",X"9A",X"32",X"A6",X"9A",X"32",X"2B",X"98",X"C9",X"ED",
		X"44",X"C6",X"0B",X"CD",X"98",X"23",X"06",X"06",X"0E",X"24",X"79",X"12",X"E7",X"10",X"FB",X"C9",
		X"CB",X"76",X"28",X"46",X"3A",X"0D",X"92",X"A7",X"28",X"07",X"CB",X"6E",X"20",X"03",X"36",X"68",
		X"C9",X"AF",X"32",X"18",X"90",X"32",X"A5",X"9A",X"32",X"A6",X"9A",X"3A",X"0D",X"92",X"A7",X"3A",
		X"29",X"98",X"20",X"0F",X"C6",X"0D",X"5F",X"16",X"91",X"AF",X"32",X"2B",X"98",X"3C",X"32",X"28",
		X"98",X"12",X"C9",X"C6",X"08",X"6F",X"26",X"91",X"11",X"6B",X"04",X"73",X"2C",X"72",X"AF",X"32",
		X"BA",X"99",X"3C",X"32",X"11",X"90",X"32",X"8E",X"92",X"C9",X"3E",X"40",X"32",X"8C",X"92",X"3E",
		X"40",X"32",X"8B",X"92",X"C9",X"3E",X"03",X"32",X"2A",X"98",X"36",X"80",X"AF",X"32",X"8D",X"92",
		X"32",X"BA",X"99",X"3C",X"32",X"8C",X"92",X"32",X"14",X"90",X"C9",X"3A",X"8B",X"92",X"FE",X"40",
		X"C0",X"3A",X"15",X"92",X"4F",X"3A",X"62",X"93",X"CB",X"41",X"28",X"04",X"C6",X"0E",X"ED",X"44",
		X"47",X"3A",X"8A",X"92",X"90",X"C6",X"1B",X"FE",X"36",X"D0",X"3A",X"01",X"92",X"3D",X"28",X"0B",
		X"3A",X"14",X"90",X"4F",X"3A",X"13",X"92",X"EE",X"01",X"A1",X"C8",X"AF",X"32",X"14",X"90",X"32",
		X"A5",X"9A",X"32",X"25",X"90",X"32",X"13",X"92",X"3C",X"32",X"1C",X"90",X"32",X"A6",X"9A",X"32",
		X"BA",X"99",X"3E",X"0A",X"32",X"2A",X"98",X"C9",X"4F",X"3A",X"8A",X"92",X"ED",X"44",X"C6",X"10",
		X"16",X"20",X"07",X"CB",X"12",X"07",X"CB",X"12",X"E6",X"E0",X"C6",X"14",X"81",X"5F",X"C9",X"24",
		X"4E",X"4F",X"50",X"51",X"24",X"24",X"52",X"53",X"54",X"55",X"24",X"24",X"56",X"57",X"58",X"59",
		X"24",X"24",X"5A",X"5B",X"5C",X"5D",X"24",X"24",X"5E",X"5F",X"60",X"61",X"24",X"62",X"63",X"64",
		X"65",X"66",X"67",X"68",X"69",X"6A",X"6B",X"6C",X"6D",X"6E",X"6F",X"70",X"71",X"72",X"73",X"74",
		X"75",X"76",X"77",X"78",X"79",X"7A",X"7B",X"7C",X"7D",X"7E",X"7F",X"3A",X"A0",X"92",X"CB",X"47",
		X"CA",X"A4",X"25",X"E6",X"02",X"5F",X"3A",X"A6",X"92",X"DD",X"6F",X"06",X"20",X"16",X"88",X"1A",
		X"CB",X"27",X"38",X"20",X"21",X"0D",X"24",X"D7",X"7E",X"23",X"66",X"6F",X"E9",X"24",X"24",X"96",
		X"24",X"6D",X"24",X"5B",X"25",X"C0",X"24",X"43",X"25",X"5B",X"25",X"9E",X"25",X"4A",X"24",X"30",
		X"24",X"1D",X"DD",X"2C",X"3E",X"04",X"83",X"5F",X"10",X"D3",X"DD",X"7D",X"32",X"A6",X"92",X"C9",
		X"6B",X"26",X"01",X"4E",X"2C",X"6E",X"26",X"99",X"7E",X"08",X"69",X"4E",X"1C",X"1A",X"C6",X"11",
		X"6F",X"26",X"91",X"08",X"77",X"2C",X"71",X"C3",X"21",X"24",X"26",X"8B",X"6B",X"1C",X"1A",X"3D",
		X"28",X"0D",X"12",X"1D",X"E6",X"03",X"20",X"CC",X"7E",X"C6",X"04",X"77",X"C3",X"24",X"24",X"26",
		X"93",X"AF",X"77",X"26",X"9B",X"77",X"1D",X"3E",X"80",X"12",X"C3",X"24",X"24",X"26",X"9B",X"6B",
		X"7E",X"E6",X"01",X"26",X"8B",X"20",X"0A",X"7E",X"E6",X"07",X"FE",X"06",X"28",X"13",X"34",X"18",
		X"28",X"7E",X"E6",X"07",X"20",X"08",X"26",X"9B",X"CB",X"86",X"26",X"8B",X"18",X"1B",X"35",X"18",
		X"18",X"3E",X"01",X"12",X"18",X"13",X"26",X"8B",X"6B",X"3A",X"A2",X"92",X"CB",X"0E",X"0F",X"0F",
		X"CB",X"16",X"3A",X"0B",X"92",X"A7",X"CA",X"22",X"24",X"26",X"01",X"4E",X"2C",X"6E",X"26",X"98",
		X"7E",X"16",X"93",X"12",X"1C",X"69",X"7E",X"12",X"16",X"9B",X"2C",X"7E",X"12",X"C3",X"21",X"24",
		X"6B",X"1C",X"1A",X"FE",X"45",X"28",X"2D",X"3C",X"12",X"1D",X"FE",X"45",X"20",X"02",X"C6",X"03",
		X"FE",X"44",X"20",X"1A",X"26",X"93",X"08",X"7E",X"D6",X"08",X"77",X"2C",X"7E",X"D6",X"08",X"77",
		X"30",X"06",X"26",X"9B",X"7E",X"EE",X"01",X"77",X"2D",X"26",X"9B",X"36",X"0C",X"08",X"26",X"8B",
		X"77",X"C3",X"24",X"24",X"1D",X"26",X"92",X"7E",X"FE",X"01",X"20",X"0F",X"26",X"93",X"36",X"00",
		X"26",X"9B",X"36",X"00",X"26",X"88",X"36",X"80",X"C3",X"24",X"24",X"26",X"8B",X"77",X"FE",X"37",
		X"38",X"0A",X"0E",X"0D",X"2C",X"FE",X"3A",X"38",X"01",X"0C",X"71",X"2D",X"26",X"93",X"0E",X"08",
		X"FE",X"3B",X"30",X"06",X"0E",X"00",X"7E",X"C6",X"08",X"77",X"2C",X"7E",X"C6",X"08",X"77",X"26",
		X"9B",X"30",X"04",X"7E",X"EE",X"01",X"77",X"2D",X"71",X"26",X"88",X"36",X"05",X"2C",X"36",X"13",
		X"C3",X"24",X"24",X"6B",X"2C",X"62",X"35",X"C2",X"24",X"24",X"2D",X"36",X"80",X"26",X"93",X"36",
		X"00",X"26",X"9B",X"36",X"00",X"3E",X"80",X"12",X"C3",X"24",X"24",X"26",X"93",X"6B",X"CB",X"FD",
		X"7E",X"FE",X"F4",X"30",X"1A",X"2C",X"4E",X"26",X"9B",X"7E",X"2D",X"0F",X"79",X"1F",X"FE",X"0B",
		X"38",X"0D",X"FE",X"A5",X"30",X"09",X"1A",X"FE",X"06",X"C2",X"22",X"24",X"C3",X"24",X"24",X"CB",
		X"BD",X"1A",X"FE",X"03",X"28",X"0A",X"3E",X"80",X"12",X"26",X"93",X"36",X"00",X"C3",X"24",X"24",
		X"1C",X"1A",X"1D",X"C6",X"13",X"6F",X"26",X"91",X"36",X"00",X"6B",X"C3",X"86",X"25",X"3E",X"03",
		X"12",X"C3",X"22",X"24",X"CB",X"4F",X"C8",X"21",X"A6",X"92",X"7E",X"36",X"00",X"2C",X"77",X"C9",
		X"21",X"7C",X"28",X"22",X"E0",X"92",X"3A",X"21",X"98",X"4F",X"FE",X"17",X"38",X"04",X"D6",X"04",
		X"18",X"F8",X"47",X"3C",X"E6",X"03",X"28",X"19",X"3A",X"84",X"99",X"2E",X"11",X"CD",X"4E",X"10",
		X"7D",X"21",X"B6",X"26",X"D7",X"11",X"02",X"27",X"78",X"CB",X"38",X"CB",X"38",X"90",X"3D",X"18",
		X"0D",X"21",X"FA",X"26",X"79",X"CB",X"3F",X"CB",X"3F",X"E6",X"07",X"11",X"EC",X"27",X"D7",X"7E",
		X"EB",X"D7",X"7E",X"23",X"32",X"E2",X"92",X"7E",X"23",X"32",X"E3",X"92",X"11",X"20",X"89",X"3E",
		X"7E",X"12",X"1C",X"7E",X"23",X"FE",X"FF",X"CA",X"8F",X"26",X"4F",X"D5",X"E5",X"21",X"00",X"91",
		X"3E",X"FF",X"06",X"10",X"DF",X"79",X"E6",X"0F",X"28",X"2A",X"47",X"CB",X"3F",X"C6",X"04",X"5F",
		X"CD",X"00",X"10",X"6F",X"26",X"00",X"7B",X"CD",X"61",X"10",X"CB",X"40",X"28",X"02",X"CB",X"DF",
		X"26",X"91",X"6F",X"7E",X"3C",X"20",X"E9",X"78",X"07",X"CB",X"01",X"30",X"02",X"F6",X"40",X"F6",
		X"38",X"77",X"10",X"DC",X"21",X"00",X"91",X"ED",X"5B",X"E0",X"92",X"06",X"08",X"7E",X"FE",X"FF",
		X"28",X"03",X"23",X"18",X"F8",X"1A",X"77",X"13",X"23",X"78",X"FE",X"05",X"20",X"02",X"2E",X"08",
		X"10",X"EB",X"ED",X"53",X"E0",X"92",X"E1",X"D1",X"46",X"23",X"4E",X"23",X"E5",X"21",X"00",X"91",
		X"78",X"12",X"7E",X"FE",X"FF",X"28",X"10",X"1C",X"12",X"1C",X"79",X"12",X"1C",X"CB",X"DD",X"7E",
		X"12",X"1C",X"CB",X"9D",X"23",X"18",X"E9",X"3E",X"7E",X"12",X"1C",X"E1",X"C3",X"03",X"26",X"1D",
		X"3A",X"2B",X"98",X"47",X"3A",X"27",X"98",X"3D",X"A0",X"28",X"17",X"3A",X"25",X"98",X"A7",X"28",
		X"11",X"62",X"7B",X"D6",X"04",X"6F",X"7E",X"12",X"1C",X"3E",X"04",X"12",X"1C",X"3E",X"87",X"32",
		X"04",X"8B",X"3E",X"7F",X"12",X"C9",X"00",X"12",X"24",X"36",X"00",X"48",X"6C",X"5A",X"48",X"6C",
		X"00",X"7E",X"A2",X"90",X"B4",X"D8",X"C6",X"00",X"12",X"48",X"6C",X"5A",X"7E",X"A2",X"00",X"7E",
		X"D8",X"C6",X"B4",X"D8",X"C6",X"B4",X"D8",X"C6",X"00",X"12",X"7E",X"A2",X"90",X"7E",X"D8",X"C6",
		X"B4",X"D8",X"C6",X"B4",X"D8",X"C6",X"B4",X"D8",X"C6",X"00",X"12",X"48",X"36",X"24",X"48",X"6C",
		X"00",X"7E",X"A2",X"90",X"B4",X"D8",X"00",X"B4",X"D8",X"C6",X"00",X"12",X"24",X"36",X"48",X"5A",
		X"6C",X"7E",X"14",X"00",X"00",X"00",X"C0",X"00",X"01",X"01",X"00",X"41",X"41",X"00",X"40",X"40",
		X"00",X"00",X"00",X"FF",X"14",X"01",X"00",X"42",X"82",X"00",X"03",X"85",X"00",X"43",X"C5",X"00",
		X"42",X"C4",X"00",X"02",X"84",X"FF",X"14",X"01",X"82",X"00",X"C0",X"00",X"01",X"01",X"00",X"41",
		X"41",X"02",X"40",X"40",X"02",X"00",X"00",X"FF",X"14",X"01",X"82",X"02",X"C2",X"00",X"03",X"85",
		X"00",X"43",X"C5",X"02",X"42",X"C4",X"02",X"02",X"84",X"FF",X"14",X"01",X"82",X"00",X"C0",X"00",
		X"01",X"C1",X"00",X"41",X"81",X"02",X"40",X"80",X"02",X"40",X"80",X"FF",X"14",X"01",X"82",X"00",
		X"C0",X"42",X"01",X"01",X"F2",X"41",X"41",X"02",X"40",X"40",X"02",X"00",X"00",X"FF",X"14",X"01",
		X"A4",X"02",X"C2",X"52",X"03",X"85",X"F2",X"43",X"C5",X"02",X"42",X"C4",X"02",X"02",X"84",X"FF",
		X"14",X"01",X"82",X"00",X"C0",X"52",X"01",X"C1",X"F2",X"41",X"81",X"02",X"40",X"80",X"02",X"40",
		X"80",X"FF",X"14",X"01",X"A4",X"00",X"C0",X"42",X"01",X"01",X"F4",X"41",X"41",X"04",X"40",X"40",
		X"04",X"00",X"00",X"FF",X"14",X"01",X"A4",X"02",X"C2",X"52",X"03",X"85",X"F4",X"43",X"C5",X"04",
		X"42",X"C4",X"04",X"02",X"84",X"FF",X"14",X"03",X"A4",X"00",X"C0",X"54",X"01",X"C1",X"F4",X"41",
		X"81",X"04",X"40",X"80",X"04",X"40",X"80",X"FF",X"14",X"03",X"A4",X"00",X"C0",X"54",X"01",X"01",
		X"F4",X"41",X"41",X"04",X"40",X"40",X"04",X"00",X"00",X"FF",X"14",X"03",X"A4",X"02",X"C2",X"54",
		X"03",X"85",X"F4",X"43",X"C5",X"04",X"42",X"C4",X"04",X"02",X"84",X"FF",X"FF",X"00",X"00",X"06",
		X"C6",X"00",X"07",X"07",X"00",X"47",X"47",X"00",X"46",X"46",X"00",X"06",X"06",X"FF",X"FF",X"00",
		X"00",X"08",X"C8",X"00",X"09",X"C9",X"00",X"09",X"C9",X"00",X"48",X"48",X"00",X"08",X"08",X"FF",
		X"FF",X"00",X"00",X"0A",X"4A",X"00",X"0B",X"CB",X"00",X"0B",X"CB",X"00",X"0A",X"4A",X"00",X"16",
		X"56",X"FF",X"FF",X"00",X"00",X"0C",X"CC",X"00",X"0D",X"0D",X"00",X"4D",X"4D",X"00",X"0C",X"CC",
		X"00",X"17",X"D7",X"FF",X"FF",X"00",X"00",X"0E",X"0E",X"00",X"0F",X"0F",X"00",X"4F",X"4F",X"00",
		X"0E",X"0E",X"00",X"4E",X"4E",X"FF",X"FF",X"00",X"00",X"10",X"10",X"00",X"11",X"D1",X"00",X"11",
		X"D1",X"00",X"50",X"50",X"00",X"10",X"10",X"FF",X"FF",X"00",X"00",X"12",X"12",X"00",X"13",X"13",
		X"00",X"53",X"53",X"00",X"52",X"52",X"00",X"12",X"12",X"FF",X"FF",X"00",X"00",X"14",X"D4",X"00",
		X"15",X"15",X"00",X"55",X"55",X"00",X"14",X"D4",X"00",X"14",X"D4",X"FF",X"58",X"5A",X"5C",X"5E",
		X"28",X"2A",X"2C",X"2E",X"30",X"34",X"36",X"32",X"50",X"52",X"54",X"56",X"42",X"46",X"40",X"44",
		X"4A",X"4E",X"48",X"4C",X"1A",X"1E",X"20",X"24",X"22",X"26",X"18",X"1C",X"08",X"0C",X"12",X"16",
		X"10",X"14",X"0A",X"0E",X"21",X"20",X"89",X"22",X"22",X"98",X"FD",X"21",X"16",X"29",X"3A",X"25",
		X"98",X"A7",X"20",X"27",X"3A",X"21",X"98",X"0F",X"0F",X"4F",X"0F",X"47",X"E6",X"1C",X"78",X"28",
		X"02",X"3E",X"03",X"E6",X"03",X"21",X"0E",X"29",X"CF",X"11",X"84",X"92",X"79",X"ED",X"A0",X"ED",
		X"A0",X"21",X"1C",X"29",X"E6",X"07",X"D7",X"56",X"5A",X"18",X"03",X"11",X"24",X"36",X"21",X"08",
		X"8B",X"DD",X"2E",X"01",X"06",X"14",X"DD",X"62",X"CD",X"F7",X"28",X"06",X"08",X"DD",X"26",X"10",
		X"CD",X"F7",X"28",X"06",X"10",X"DD",X"63",X"DD",X"2D",X"20",X"08",X"FD",X"4E",X"00",X"FD",X"23",
		X"DD",X"2E",X"08",X"CB",X"01",X"DD",X"7C",X"1F",X"77",X"2C",X"2C",X"10",X"EA",X"C9",X"0A",X"B8",
		X"0F",X"B9",X"14",X"BC",X"1E",X"BD",X"A5",X"5A",X"A9",X"0F",X"0A",X"50",X"36",X"24",X"D4",X"BA",
		X"E4",X"CC",X"A8",X"F4",X"2A",X"22",X"98",X"7E",X"FE",X"7F",X"CA",X"37",X"2A",X"FE",X"7E",X"20",
		X"30",X"3A",X"42",X"98",X"A7",X"C8",X"3A",X"87",X"92",X"A7",X"20",X"1F",X"3A",X"25",X"98",X"47",
		X"A7",X"20",X"0F",X"3A",X"AC",X"92",X"FE",X"01",X"20",X"06",X"3E",X"08",X"32",X"A8",X"92",X"C9",
		X"A7",X"C0",X"23",X"22",X"22",X"98",X"21",X"26",X"98",X"34",X"C9",X"3E",X"02",X"32",X"AC",X"92",
		X"C9",X"4F",X"CB",X"7F",X"20",X"06",X"3A",X"A0",X"92",X"E6",X"07",X"C0",X"CB",X"21",X"06",X"0C",
		X"11",X"14",X"00",X"DD",X"21",X"00",X"91",X"DD",X"CB",X"13",X"46",X"28",X"05",X"DD",X"19",X"10",
		X"F6",X"C9",X"23",X"7E",X"47",X"E6",X"78",X"FE",X"78",X"78",X"20",X"02",X"CB",X"B7",X"DD",X"77",
		X"10",X"23",X"22",X"22",X"98",X"26",X"88",X"6F",X"36",X"07",X"2C",X"DD",X"5D",X"73",X"26",X"93",
		X"E6",X"38",X"FE",X"38",X"28",X"1B",X"2D",X"26",X"8B",X"7E",X"57",X"E6",X"78",X"77",X"2C",X"7A",
		X"E6",X"07",X"CB",X"7A",X"77",X"3E",X"00",X"28",X"03",X"3A",X"E3",X"92",X"DD",X"77",X"0F",X"18",
		X"1E",X"11",X"10",X"02",X"CB",X"70",X"20",X"0D",X"11",X"18",X"03",X"3A",X"26",X"98",X"FE",X"02",
		X"20",X"03",X"11",X"08",X"00",X"26",X"8B",X"72",X"2D",X"73",X"2C",X"DD",X"36",X"0F",X"00",X"51",
		X"CB",X"B9",X"06",X"08",X"CB",X"49",X"28",X"02",X"06",X"44",X"DD",X"70",X"0E",X"06",X"00",X"21",
		X"4A",X"2A",X"09",X"7E",X"23",X"DD",X"77",X"08",X"AF",X"ED",X"6F",X"47",X"7E",X"E6",X"1F",X"DD",
		X"77",X"09",X"78",X"E6",X"0E",X"47",X"07",X"80",X"21",X"7A",X"2A",X"D7",X"CB",X"7A",X"28",X"03",
		X"23",X"23",X"23",X"7E",X"23",X"DD",X"77",X"01",X"7E",X"23",X"DD",X"77",X"03",X"7E",X"23",X"DD",
		X"77",X"05",X"AF",X"DD",X"77",X"00",X"DD",X"77",X"02",X"DD",X"77",X"04",X"3C",X"DD",X"77",X"0D",
		X"B2",X"E6",X"81",X"DD",X"77",X"13",X"C9",X"3A",X"87",X"92",X"A7",X"C0",X"32",X"08",X"90",X"3C",
		X"32",X"04",X"90",X"32",X"10",X"90",X"32",X"24",X"98",X"C9",X"1D",X"00",X"67",X"20",X"9F",X"40",
		X"D4",X"20",X"7B",X"01",X"B0",X"61",X"E8",X"01",X"F5",X"21",X"0B",X"02",X"1B",X"22",X"2B",X"82",
		X"41",X"22",X"5D",X"82",X"79",X"22",X"9E",X"02",X"BA",X"22",X"D9",X"02",X"FB",X"22",X"1D",X"03",
		X"33",X"23",X"DA",X"0F",X"F0",X"2F",X"2B",X"A2",X"5D",X"A2",X"9B",X"34",X"03",X"9B",X"44",X"03",
		X"23",X"00",X"00",X"23",X"78",X"02",X"9B",X"2C",X"03",X"9B",X"4C",X"03",X"2B",X"00",X"00",X"2B",
		X"78",X"02",X"9B",X"34",X"03",X"9B",X"34",X"03",X"9B",X"44",X"03",X"9B",X"44",X"03",X"3A",X"A0",
		X"92",X"3D",X"E6",X"03",X"C0",X"3A",X"A7",X"92",X"47",X"3A",X"08",X"90",X"B0",X"28",X"48",X"3A",
		X"0F",X"92",X"A7",X"0E",X"01",X"28",X"02",X"0D",X"0D",X"2E",X"00",X"06",X"0A",X"26",X"99",X"7E",
		X"81",X"77",X"26",X"98",X"7E",X"81",X"77",X"2C",X"2C",X"10",X"F2",X"3A",X"24",X"98",X"A7",X"3A",
		X"00",X"99",X"28",X"03",X"A7",X"28",X"11",X"FE",X"20",X"20",X"06",X"3E",X"01",X"32",X"0F",X"92",
		X"C9",X"D6",X"E0",X"C0",X"32",X"0F",X"92",X"C9",X"AF",X"32",X"0F",X"92",X"32",X"0A",X"90",X"3C",
		X"32",X"A0",X"9A",X"32",X"09",X"90",X"C9",X"32",X"0A",X"90",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3A",X"21",X"98",X"FE",X"1B",X"38",X"04",X"D6",X"04",X"18",X"F8",X"3D",X"6F",X"07",X"07",X"85",
		X"5F",X"3A",X"84",X"99",X"21",X"65",X"2C",X"CF",X"7E",X"23",X"66",X"6F",X"7B",X"D7",X"11",X"C0",
		X"99",X"06",X"05",X"7E",X"4F",X"07",X"07",X"07",X"07",X"E6",X"0F",X"12",X"1C",X"79",X"E6",X"0F",
		X"12",X"1C",X"23",X"10",X"EE",X"3A",X"21",X"98",X"FE",X"03",X"30",X"03",X"AF",X"18",X"07",X"F6",
		X"FC",X"3C",X"28",X"02",X"3E",X"0A",X"12",X"01",X"16",X"02",X"ED",X"43",X"C1",X"92",X"ED",X"43",
		X"C0",X"92",X"3A",X"21",X"98",X"FE",X"10",X"38",X"02",X"3E",X"10",X"07",X"07",X"E6",X"70",X"C6",
		X"40",X"32",X"BB",X"99",X"C9",X"EF",X"2C",X"71",X"2D",X"F3",X"2D",X"6D",X"2C",X"00",X"00",X"22",
		X"C6",X"00",X"00",X"11",X"23",X"C7",X"00",X"00",X"00",X"00",X"C0",X"00",X"11",X"12",X"23",X"97",
		X"00",X"11",X"23",X"23",X"98",X"00",X"21",X"24",X"33",X"98",X"00",X"00",X"00",X"00",X"90",X"00",
		X"22",X"25",X"33",X"99",X"10",X"22",X"36",X"34",X"69",X"10",X"10",X"11",X"23",X"97",X"00",X"00",
		X"00",X"00",X"60",X"00",X"32",X"46",X"34",X"67",X"11",X"32",X"67",X"44",X"68",X"11",X"32",X"67",
		X"45",X"68",X"11",X"00",X"00",X"00",X"60",X"00",X"42",X"78",X"45",X"69",X"11",X"42",X"78",X"45",
		X"69",X"11",X"11",X"22",X"23",X"97",X"11",X"00",X"00",X"00",X"60",X"00",X"52",X"88",X"46",X"3A",
		X"11",X"52",X"88",X"56",X"3A",X"11",X"52",X"88",X"56",X"3C",X"11",X"00",X"00",X"00",X"30",X"00",
		X"62",X"89",X"57",X"3C",X"11",X"62",X"99",X"57",X"3C",X"11",X"62",X"99",X"57",X"3C",X"11",X"00",
		X"00",X"12",X"C6",X"00",X"00",X"11",X"22",X"C6",X"00",X"00",X"00",X"00",X"C0",X"00",X"11",X"12",
		X"23",X"97",X"00",X"11",X"12",X"23",X"97",X"00",X"00",X"11",X"23",X"C7",X"00",X"00",X"00",X"00",
		X"90",X"00",X"21",X"23",X"33",X"98",X"10",X"21",X"24",X"33",X"98",X"10",X"21",X"25",X"34",X"98",
		X"10",X"00",X"00",X"00",X"60",X"00",X"22",X"25",X"34",X"68",X"11",X"32",X"36",X"44",X"68",X"11",
		X"11",X"11",X"23",X"67",X"01",X"00",X"00",X"00",X"60",X"00",X"32",X"36",X"45",X"68",X"11",X"32",
		X"46",X"45",X"69",X"11",X"32",X"67",X"45",X"69",X"11",X"00",X"00",X"00",X"60",X"00",X"42",X"67",
		X"46",X"3A",X"11",X"42",X"78",X"56",X"3A",X"11",X"52",X"78",X"56",X"3A",X"11",X"00",X"00",X"00",
		X"30",X"00",X"52",X"88",X"56",X"3C",X"11",X"62",X"99",X"57",X"3C",X"11",X"62",X"99",X"57",X"3C",
		X"11",X"00",X"00",X"23",X"C6",X"00",X"10",X"11",X"23",X"97",X"00",X"00",X"00",X"00",X"C0",X"00",
		X"11",X"12",X"33",X"98",X"00",X"21",X"23",X"34",X"68",X"00",X"21",X"24",X"34",X"68",X"00",X"00",
		X"00",X"00",X"90",X"00",X"32",X"36",X"34",X"67",X"10",X"32",X"46",X"44",X"68",X"10",X"11",X"11",
		X"23",X"97",X"10",X"00",X"00",X"00",X"60",X"00",X"42",X"67",X"45",X"68",X"11",X"42",X"67",X"45",
		X"69",X"11",X"42",X"78",X"46",X"69",X"11",X"00",X"00",X"00",X"60",X"00",X"52",X"78",X"46",X"3A",
		X"11",X"52",X"88",X"56",X"3A",X"11",X"52",X"88",X"56",X"3A",X"11",X"00",X"00",X"00",X"60",X"00",
		X"62",X"88",X"56",X"3C",X"11",X"62",X"89",X"57",X"3C",X"11",X"62",X"89",X"57",X"3E",X"11",X"00",
		X"00",X"00",X"30",X"00",X"72",X"99",X"57",X"3E",X"11",X"72",X"99",X"68",X"3E",X"11",X"72",X"99",
		X"68",X"3E",X"11",X"00",X"00",X"23",X"C6",X"00",X"10",X"11",X"23",X"97",X"00",X"00",X"00",X"00",
		X"C0",X"00",X"11",X"12",X"34",X"98",X"00",X"21",X"23",X"34",X"68",X"00",X"21",X"24",X"34",X"68",
		X"00",X"00",X"00",X"00",X"90",X"00",X"32",X"36",X"45",X"67",X"11",X"32",X"46",X"46",X"68",X"11",
		X"32",X"56",X"46",X"69",X"11",X"00",X"00",X"00",X"60",X"00",X"42",X"67",X"56",X"6A",X"11",X"42",
		X"67",X"56",X"6A",X"11",X"42",X"78",X"57",X"6A",X"11",X"00",X"00",X"00",X"60",X"00",X"52",X"78",
		X"57",X"3A",X"11",X"52",X"88",X"57",X"3A",X"11",X"52",X"88",X"68",X"3C",X"11",X"00",X"00",X"00",
		X"60",X"00",X"62",X"88",X"68",X"3C",X"11",X"62",X"89",X"68",X"3C",X"11",X"62",X"89",X"68",X"3E",
		X"11",X"00",X"00",X"00",X"30",X"00",X"72",X"99",X"68",X"3E",X"11",X"72",X"99",X"68",X"3E",X"11",
		X"72",X"99",X"68",X"3E",X"11",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"50",
		X"21",X"FD",X"83",X"3A",X"40",X"98",X"A7",X"28",X"03",X"21",X"E8",X"83",X"22",X"00",X"8A",X"11",
		X"3D",X"8A",X"CD",X"F7",X"31",X"D0",X"11",X"37",X"8A",X"CD",X"F7",X"31",X"3E",X"05",X"30",X"27",
		X"11",X"31",X"8A",X"CD",X"F7",X"31",X"3E",X"04",X"30",X"1D",X"11",X"2B",X"8A",X"CD",X"F7",X"31",
		X"3E",X"03",X"30",X"13",X"11",X"25",X"8A",X"CD",X"F7",X"31",X"3E",X"02",X"30",X"09",X"3E",X"FF",
		X"32",X"AC",X"9A",X"3E",X"01",X"18",X"03",X"32",X"B0",X"9A",X"32",X"11",X"8A",X"21",X"A6",X"31",
		X"3D",X"CF",X"CD",X"18",X"31",X"3A",X"11",X"8A",X"21",X"A1",X"31",X"3D",X"D7",X"7E",X"21",X"49",
		X"8A",X"11",X"4C",X"8A",X"A7",X"28",X"05",X"4F",X"06",X"00",X"ED",X"B8",X"06",X"03",X"3E",X"24",
		X"22",X"04",X"8A",X"2C",X"77",X"10",X"FC",X"3E",X"49",X"32",X"10",X"8A",X"21",X"7F",X"32",X"CD",
		X"28",X"33",X"CD",X"1B",X"33",X"CD",X"28",X"33",X"11",X"09",X"83",X"2A",X"00",X"8A",X"CD",X"75",
		X"32",X"21",X"49",X"81",X"11",X"E0",X"FF",X"36",X"0A",X"19",X"36",X"0A",X"19",X"36",X"0A",X"CD",
		X"1D",X"32",X"CD",X"80",X"31",X"3E",X"04",X"32",X"AE",X"92",X"3A",X"AE",X"92",X"A7",X"20",X"FA",
		X"3E",X"28",X"32",X"AE",X"92",X"CD",X"1D",X"32",X"CD",X"80",X"31",X"3A",X"A0",X"92",X"4F",X"CD",
		X"ED",X"32",X"3A",X"A0",X"92",X"B9",X"28",X"F7",X"4F",X"E6",X"0F",X"CC",X"41",X"31",X"21",X"B6",
		X"99",X"3A",X"15",X"92",X"A7",X"28",X"01",X"23",X"CB",X"66",X"CA",X"4C",X"31",X"7E",X"E6",X"0A",
		X"21",X"02",X"8A",X"11",X"03",X"8A",X"BE",X"28",X"04",X"77",X"3E",X"FD",X"12",X"1A",X"3C",X"12",
		X"E6",X"0F",X"20",X"CB",X"7E",X"FE",X"08",X"28",X"24",X"FE",X"02",X"20",X"C2",X"3E",X"28",X"32",
		X"AE",X"92",X"3A",X"10",X"8A",X"6F",X"26",X"81",X"7E",X"3D",X"FE",X"09",X"CC",X"38",X"31",X"FE",
		X"29",X"CC",X"3B",X"31",X"77",X"C3",X"BF",X"30",X"7E",X"23",X"66",X"6F",X"E9",X"3A",X"10",X"8A",
		X"6F",X"26",X"81",X"3E",X"28",X"32",X"AE",X"92",X"7E",X"3C",X"FE",X"2B",X"CC",X"3E",X"31",X"FE",
		X"25",X"CC",X"38",X"31",X"77",X"C3",X"BF",X"30",X"3E",X"2A",X"C9",X"3E",X"24",X"C9",X"3E",X"0A",
		X"C9",X"3A",X"10",X"8A",X"6F",X"26",X"85",X"7E",X"EE",X"05",X"77",X"C9",X"3A",X"10",X"8A",X"6F",
		X"26",X"85",X"36",X"00",X"26",X"81",X"4E",X"3E",X"28",X"32",X"AE",X"92",X"2A",X"04",X"8A",X"23",
		X"71",X"22",X"04",X"8A",X"21",X"10",X"8A",X"7E",X"D6",X"20",X"77",X"D2",X"B5",X"30",X"CD",X"1D",
		X"32",X"CD",X"80",X"31",X"3E",X"4C",X"32",X"A0",X"92",X"3A",X"A0",X"92",X"A7",X"20",X"FA",X"C9",
		X"3A",X"11",X"8A",X"21",X"97",X"31",X"3D",X"CF",X"7E",X"23",X"66",X"6F",X"06",X"16",X"11",X"E0",
		X"FF",X"36",X"05",X"19",X"10",X"FB",X"C9",X"74",X"87",X"76",X"87",X"78",X"87",X"7A",X"87",X"7C",
		X"87",X"0C",X"09",X"06",X"03",X"00",X"B0",X"31",X"B4",X"31",X"B8",X"31",X"CE",X"31",X"D9",X"31",
		X"3E",X"12",X"18",X"06",X"3E",X"0C",X"18",X"02",X"3E",X"06",X"21",X"37",X"8A",X"11",X"3D",X"8A",
		X"01",X"06",X"00",X"ED",X"B8",X"11",X"37",X"8A",X"4F",X"ED",X"B8",X"C3",X"D9",X"31",X"11",X"3D",
		X"8A",X"21",X"37",X"8A",X"01",X"06",X"00",X"ED",X"B8",X"3A",X"11",X"8A",X"3D",X"21",X"ED",X"31",
		X"CF",X"5E",X"23",X"56",X"2A",X"00",X"8A",X"01",X"06",X"00",X"ED",X"B8",X"C9",X"25",X"8A",X"2B",
		X"8A",X"31",X"8A",X"37",X"8A",X"3D",X"8A",X"2A",X"00",X"8A",X"06",X"06",X"1A",X"FE",X"24",X"28",
		X"0D",X"7E",X"FE",X"24",X"C8",X"1A",X"BE",X"C0",X"2D",X"1D",X"10",X"F0",X"AF",X"C9",X"BE",X"28",
		X"F7",X"AF",X"18",X"F2",X"21",X"45",X"33",X"CD",X"28",X"33",X"CD",X"28",X"33",X"21",X"B4",X"32",
		X"CD",X"1B",X"33",X"06",X"01",X"CD",X"31",X"32",X"CD",X"31",X"32",X"CD",X"31",X"32",X"CD",X"31",
		X"32",X"78",X"3D",X"87",X"87",X"87",X"21",X"C5",X"32",X"D7",X"5E",X"23",X"56",X"23",X"78",X"12",
		X"CD",X"73",X"32",X"CD",X"70",X"32",X"CD",X"70",X"32",X"CD",X"73",X"32",X"CD",X"73",X"32",X"7E",
		X"23",X"4E",X"23",X"E5",X"61",X"6F",X"CD",X"75",X"32",X"7B",X"D6",X"C0",X"5F",X"30",X"01",X"15",
		X"E1",X"7E",X"23",X"66",X"6F",X"CD",X"70",X"32",X"CD",X"70",X"32",X"CD",X"70",X"32",X"04",X"C9",
		X"7E",X"12",X"23",X"E7",X"C9",X"0E",X"06",X"7E",X"12",X"2B",X"E7",X"0D",X"20",X"F9",X"C9",X"24",
		X"83",X"15",X"04",X"0E",X"17",X"1D",X"0E",X"1B",X"24",X"22",X"18",X"1E",X"1B",X"24",X"12",X"17",
		X"12",X"1D",X"12",X"0A",X"15",X"1C",X"24",X"2C",X"E7",X"82",X"10",X"1C",X"0C",X"18",X"1B",X"0E",
		X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"17",X"0A",X"16",X"0E",X"50",X"82",X"05",X"04",X"1D",
		X"18",X"19",X"24",X"05",X"92",X"82",X"0E",X"1C",X"0C",X"18",X"1B",X"0E",X"24",X"24",X"24",X"24",
		X"24",X"17",X"0A",X"16",X"0E",X"54",X"83",X"1C",X"1D",X"25",X"8A",X"3E",X"8A",X"56",X"83",X"17",
		X"0D",X"2B",X"8A",X"41",X"8A",X"58",X"83",X"1B",X"0D",X"31",X"8A",X"44",X"8A",X"5A",X"83",X"1D",
		X"11",X"37",X"8A",X"47",X"8A",X"5C",X"83",X"1D",X"11",X"3D",X"8A",X"4A",X"8A",X"3A",X"B5",X"99",
		X"FE",X"A0",X"28",X"07",X"47",X"3A",X"B8",X"99",X"B8",X"38",X"05",X"3A",X"AE",X"92",X"A7",X"C0",
		X"E1",X"26",X"81",X"3A",X"10",X"8A",X"6F",X"ED",X"5B",X"04",X"8A",X"13",X"ED",X"A0",X"3E",X"DF",
		X"25",X"85",X"30",X"01",X"24",X"6F",X"CB",X"44",X"20",X"F2",X"C9",X"5E",X"23",X"56",X"23",X"46",
		X"23",X"7E",X"12",X"23",X"E7",X"10",X"FA",X"C9",X"5E",X"23",X"56",X"23",X"46",X"23",X"4E",X"23",
		X"EB",X"1A",X"77",X"CB",X"D4",X"71",X"CB",X"94",X"13",X"3E",X"E0",X"25",X"85",X"30",X"01",X"24",
		X"6F",X"10",X"EE",X"EB",X"C9",X"25",X"83",X"13",X"02",X"1D",X"11",X"0E",X"24",X"10",X"0A",X"15",
		X"0A",X"0C",X"1D",X"12",X"0C",X"24",X"11",X"0E",X"1B",X"18",X"0E",X"1C",X"CC",X"82",X"0C",X"04",
		X"26",X"26",X"24",X"0B",X"0E",X"1C",X"1D",X"24",X"05",X"24",X"26",X"26",X"AF",X"32",X"23",X"68",
		X"3C",X"32",X"22",X"68",X"F3",X"32",X"30",X"68",X"06",X"0A",X"D9",X"11",X"00",X"80",X"21",X"00",
		X"00",X"01",X"00",X"04",X"7D",X"AC",X"2F",X"87",X"87",X"ED",X"6A",X"7D",X"32",X"30",X"68",X"12",
		X"13",X"0B",X"78",X"B1",X"20",X"EE",X"11",X"00",X"80",X"21",X"00",X"00",X"01",X"00",X"04",X"7D",
		X"AC",X"2F",X"87",X"87",X"ED",X"6A",X"1A",X"AD",X"C2",X"C0",X"34",X"13",X"32",X"30",X"68",X"0B",
		X"78",X"B1",X"20",X"EB",X"11",X"00",X"80",X"21",X"55",X"55",X"01",X"00",X"04",X"7D",X"AC",X"2F",
		X"87",X"87",X"ED",X"6A",X"7D",X"32",X"30",X"68",X"12",X"13",X"0B",X"78",X"B1",X"20",X"EE",X"11",
		X"00",X"80",X"21",X"55",X"55",X"01",X"00",X"04",X"7D",X"AC",X"2F",X"87",X"87",X"ED",X"6A",X"1A",
		X"AD",X"C2",X"C0",X"34",X"13",X"32",X"30",X"68",X"0B",X"78",X"B1",X"20",X"EB",X"11",X"00",X"80",
		X"21",X"AA",X"AA",X"01",X"00",X"04",X"7D",X"AC",X"2F",X"87",X"87",X"ED",X"6A",X"7D",X"32",X"30",
		X"68",X"12",X"13",X"0B",X"78",X"B1",X"20",X"EE",X"11",X"00",X"80",X"21",X"AA",X"AA",X"01",X"00",
		X"04",X"7D",X"AC",X"2F",X"87",X"87",X"ED",X"6A",X"1A",X"AD",X"C2",X"C0",X"34",X"13",X"32",X"30",
		X"68",X"0B",X"78",X"B1",X"20",X"EB",X"D9",X"05",X"C2",X"7A",X"33",X"31",X"00",X"84",X"11",X"00",
		X"84",X"CD",X"7F",X"34",X"11",X"00",X"88",X"CD",X"7F",X"34",X"11",X"00",X"90",X"CD",X"7F",X"34",
		X"21",X"E0",X"99",X"11",X"00",X"90",X"01",X"20",X"00",X"ED",X"B0",X"11",X"00",X"98",X"CD",X"7F",
		X"34",X"21",X"00",X"90",X"11",X"E0",X"99",X"01",X"20",X"00",X"ED",X"B0",X"31",X"00",X"8B",X"11",
		X"00",X"80",X"CD",X"7F",X"34",X"CD",X"58",X"39",X"21",X"81",X"3B",X"CD",X"1B",X"33",X"32",X"30",
		X"68",X"CD",X"3C",X"3A",X"3E",X"07",X"32",X"20",X"90",X"CD",X"72",X"39",X"C3",X"50",X"35",X"06",
		X"1E",X"21",X"00",X"00",X"C5",X"CD",X"8C",X"34",X"C1",X"10",X"F9",X"C9",X"D5",X"E5",X"01",X"00",
		X"04",X"7D",X"AC",X"2F",X"87",X"87",X"ED",X"6A",X"7D",X"32",X"30",X"68",X"12",X"13",X"0B",X"78",
		X"B1",X"20",X"EE",X"E1",X"D1",X"D5",X"01",X"00",X"04",X"7D",X"AC",X"2F",X"87",X"87",X"ED",X"6A",
		X"1A",X"AD",X"C2",X"C0",X"34",X"13",X"32",X"30",X"68",X"0B",X"78",X"B1",X"20",X"EB",X"D1",X"C9",
		X"47",X"7A",X"1F",X"1F",X"E6",X"07",X"FE",X"04",X"38",X"01",X"3D",X"FE",X"05",X"38",X"01",X"3D",
		X"5F",X"78",X"16",X"15",X"E6",X"0F",X"20",X"02",X"16",X"11",X"32",X"30",X"68",X"D9",X"21",X"00",
		X"80",X"11",X"01",X"80",X"01",X"00",X"04",X"36",X"24",X"ED",X"B0",X"36",X"00",X"01",X"FF",X"03",
		X"ED",X"B0",X"32",X"30",X"68",X"D9",X"21",X"E2",X"82",X"36",X"1B",X"3E",X"E0",X"25",X"D7",X"36",
		X"0A",X"3E",X"E0",X"25",X"D7",X"36",X"16",X"3E",X"A0",X"25",X"D7",X"73",X"3E",X"E0",X"25",X"D7",
		X"72",X"21",X"80",X"93",X"06",X"80",X"36",X"F1",X"23",X"10",X"FB",X"32",X"30",X"68",X"C3",X"1B",
		X"35",X"E5",X"EB",X"16",X"10",X"AF",X"47",X"86",X"32",X"30",X"68",X"23",X"10",X"F9",X"15",X"20",
		X"F6",X"EB",X"E1",X"B9",X"C8",X"21",X"8B",X"3B",X"CD",X"1B",X"33",X"11",X"44",X"82",X"21",X"02",
		X"91",X"AF",X"ED",X"6F",X"12",X"E7",X"AF",X"ED",X"6F",X"12",X"32",X"30",X"68",X"C3",X"4A",X"35",
		X"21",X"00",X"91",X"36",X"00",X"23",X"36",X"00",X"23",X"36",X"01",X"AF",X"32",X"70",X"92",X"3C",
		X"32",X"23",X"68",X"11",X"00",X"00",X"0E",X"00",X"CD",X"21",X"35",X"34",X"0E",X"00",X"CD",X"21",
		X"35",X"34",X"0E",X"00",X"CD",X"21",X"35",X"34",X"0E",X"00",X"CD",X"21",X"35",X"36",X"FF",X"3A",
		X"00",X"91",X"32",X"30",X"68",X"A7",X"28",X"F7",X"3C",X"28",X"07",X"3D",X"32",X"02",X"91",X"C3",
		X"35",X"35",X"3A",X"01",X"91",X"32",X"30",X"68",X"A7",X"28",X"F7",X"3C",X"28",X"17",X"3D",X"32",
		X"02",X"91",X"C3",X"35",X"35",X"05",X"05",X"05",X"05",X"30",X"40",X"00",X"02",X"DF",X"40",X"30",
		X"30",X"03",X"DF",X"10",X"20",X"21",X"8B",X"3B",X"CD",X"1B",X"33",X"CD",X"F4",X"37",X"21",X"00",
		X"91",X"06",X"03",X"36",X"00",X"23",X"10",X"FB",X"3E",X"20",X"32",X"00",X"90",X"21",X"A5",X"35",
		X"11",X"00",X"70",X"01",X"04",X"00",X"D9",X"3E",X"A1",X"32",X"00",X"71",X"32",X"30",X"68",X"CD",
		X"EC",X"37",X"AF",X"32",X"30",X"68",X"32",X"A0",X"92",X"3A",X"A0",X"92",X"FE",X"02",X"20",X"F9",
		X"21",X"A9",X"35",X"11",X"00",X"70",X"01",X"0C",X"00",X"D9",X"3E",X"A8",X"32",X"00",X"71",X"32",
		X"30",X"68",X"CD",X"EC",X"37",X"32",X"30",X"68",X"ED",X"56",X"21",X"20",X"68",X"36",X"00",X"36",
		X"01",X"FB",X"CD",X"F2",X"39",X"AF",X"32",X"A0",X"92",X"3A",X"A0",X"92",X"E6",X"08",X"28",X"F9",
		X"3A",X"A0",X"92",X"4F",X"3A",X"A0",X"92",X"B9",X"28",X"FA",X"21",X"16",X"91",X"11",X"17",X"91",
		X"01",X"07",X"00",X"ED",X"B8",X"EB",X"11",X"B5",X"99",X"1A",X"CB",X"7F",X"C2",X"BA",X"36",X"77",
		X"23",X"B6",X"23",X"2F",X"A6",X"23",X"A6",X"77",X"47",X"23",X"13",X"1A",X"77",X"23",X"B6",X"23",
		X"2F",X"A6",X"23",X"A6",X"77",X"6F",X"60",X"06",X"10",X"29",X"DC",X"D6",X"39",X"10",X"FA",X"CD",
		X"F4",X"37",X"2A",X"72",X"92",X"7C",X"B5",X"28",X"09",X"2B",X"22",X"72",X"92",X"7C",X"B5",X"CC",
		X"BB",X"39",X"3A",X"10",X"91",X"1F",X"30",X"07",X"AF",X"32",X"71",X"92",X"C3",X"20",X"36",X"3A",
		X"17",X"91",X"E6",X"0F",X"CA",X"20",X"36",X"4F",X"21",X"82",X"37",X"11",X"71",X"92",X"1A",X"D7",
		X"7E",X"B9",X"28",X"05",X"AF",X"12",X"C3",X"20",X"36",X"EB",X"34",X"13",X"1A",X"3C",X"C2",X"20",
		X"36",X"CD",X"58",X"39",X"CD",X"72",X"39",X"11",X"98",X"37",X"21",X"42",X"80",X"06",X"1C",X"CD",
		X"66",X"37",X"10",X"FB",X"3A",X"B5",X"99",X"87",X"30",X"FA",X"AF",X"32",X"A0",X"92",X"3A",X"A0",
		X"92",X"FE",X"08",X"38",X"F9",X"3A",X"B5",X"99",X"87",X"D2",X"20",X"36",X"CD",X"72",X"39",X"21",
		X"00",X"80",X"06",X"10",X"36",X"28",X"23",X"36",X"27",X"23",X"10",X"F8",X"06",X"10",X"36",X"2D",
		X"23",X"36",X"2B",X"23",X"10",X"F8",X"06",X"10",X"36",X"28",X"23",X"36",X"2D",X"23",X"10",X"F8",
		X"06",X"10",X"36",X"27",X"23",X"36",X"2B",X"23",X"10",X"F8",X"EB",X"21",X"40",X"80",X"01",X"40",
		X"03",X"ED",X"B0",X"21",X"00",X"80",X"01",X"40",X"00",X"ED",X"B0",X"AF",X"32",X"A0",X"92",X"3A",
		X"A0",X"92",X"87",X"30",X"FA",X"3A",X"B5",X"99",X"87",X"30",X"FA",X"F3",X"CD",X"EC",X"37",X"3E",
		X"FE",X"32",X"A0",X"92",X"3A",X"A0",X"92",X"A7",X"20",X"FA",X"32",X"30",X"68",X"21",X"80",X"92",
		X"11",X"00",X"70",X"01",X"08",X"00",X"D9",X"3E",X"E1",X"32",X"00",X"71",X"CD",X"EC",X"37",X"21",
		X"00",X"70",X"11",X"88",X"92",X"01",X"03",X"00",X"D9",X"3E",X"B1",X"32",X"00",X"71",X"CD",X"EC",
		X"37",X"3A",X"88",X"92",X"FE",X"A1",X"30",X"D5",X"E6",X"0F",X"FE",X"0A",X"30",X"CF",X"FB",X"AF",
		X"32",X"10",X"82",X"C3",X"D3",X"02",X"CD",X"74",X"37",X"CD",X"74",X"37",X"CD",X"74",X"37",X"3E",
		X"05",X"C3",X"10",X"00",X"1A",X"0E",X"08",X"87",X"30",X"01",X"34",X"23",X"0D",X"20",X"F8",X"13",
		X"23",X"C9",X"02",X"02",X"02",X"02",X"02",X"08",X"08",X"08",X"08",X"08",X"08",X"02",X"02",X"02",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"FF",X"01",X"3E",X"00",X"7F",X"41",X"00",X"21",X"41",
		X"00",X"00",X"41",X"00",X"36",X"3E",X"00",X"49",X"00",X"03",X"49",X"22",X"03",X"49",X"41",X"00",
		X"36",X"41",X"3E",X"00",X"3E",X"41",X"3E",X"00",X"41",X"49",X"7F",X"41",X"49",X"20",X"7F",X"49",
		X"18",X"00",X"32",X"20",X"40",X"00",X"7F",X"40",X"01",X"00",X"7F",X"7F",X"3F",X"40",X"21",X"44",
		X"40",X"00",X"44",X"00",X"3C",X"44",X"01",X"42",X"3F",X"01",X"81",X"00",X"01",X"A5",X"7F",X"01",
		X"A5",X"04",X"7F",X"99",X"08",X"00",X"42",X"10",X"00",X"3C",X"7F",X"00",X"3A",X"00",X"71",X"FE",
		X"10",X"C8",X"18",X"F8",X"3A",X"07",X"68",X"1F",X"3C",X"E6",X"01",X"32",X"83",X"99",X"21",X"CC",
		X"3A",X"CF",X"CD",X"61",X"3A",X"3A",X"B5",X"99",X"0E",X"00",X"E6",X"0C",X"20",X"01",X"0C",X"79",
		X"32",X"07",X"A0",X"21",X"01",X"68",X"7E",X"1F",X"E6",X"01",X"4F",X"23",X"7E",X"E6",X"02",X"B1",
		X"32",X"84",X"99",X"21",X"68",X"3A",X"D7",X"11",X"2C",X"82",X"ED",X"A0",X"21",X"E4",X"3A",X"CD",
		X"1B",X"33",X"21",X"06",X"68",X"7E",X"23",X"4E",X"CB",X"19",X"8F",X"E6",X"03",X"3C",X"32",X"82",
		X"99",X"3C",X"32",X"EA",X"82",X"21",X"EB",X"3A",X"CD",X"1B",X"33",X"21",X"C4",X"3A",X"11",X"80",
		X"92",X"01",X"08",X"00",X"ED",X"B0",X"21",X"00",X"68",X"06",X"03",X"AF",X"4E",X"CB",X"19",X"8F",
		X"23",X"10",X"F9",X"E6",X"07",X"28",X"34",X"3D",X"87",X"87",X"87",X"21",X"6C",X"3A",X"D7",X"11",
		X"81",X"92",X"01",X"04",X"00",X"ED",X"B0",X"11",X"E8",X"82",X"ED",X"A0",X"11",X"28",X"82",X"ED",
		X"A0",X"11",X"E8",X"81",X"ED",X"A0",X"11",X"E8",X"80",X"ED",X"A0",X"3E",X"24",X"32",X"08",X"82",
		X"21",X"F6",X"3A",X"CD",X"1B",X"33",X"CD",X"1B",X"33",X"18",X"10",X"21",X"81",X"92",X"06",X"04",
		X"36",X"00",X"23",X"10",X"FB",X"21",X"07",X"3B",X"CD",X"1B",X"33",X"21",X"03",X"68",X"06",X"03",
		X"AF",X"4E",X"CB",X"19",X"8F",X"23",X"10",X"F9",X"E6",X"07",X"CA",X"2D",X"39",X"4F",X"3A",X"82",
		X"99",X"E6",X"04",X"87",X"81",X"87",X"21",X"A4",X"3A",X"D7",X"11",X"80",X"99",X"ED",X"A0",X"ED",
		X"A0",X"2B",X"0E",X"01",X"CD",X"DA",X"38",X"2B",X"0E",X"00",X"7E",X"3C",X"CA",X"3B",X"39",X"79",
		X"87",X"E5",X"21",X"1D",X"3B",X"D7",X"7E",X"23",X"66",X"6F",X"C5",X"CD",X"1B",X"33",X"CD",X"1B",
		X"33",X"C1",X"E1",X"7E",X"E6",X"7F",X"EB",X"21",X"F0",X"81",X"41",X"10",X"02",X"23",X"23",X"CD",
		X"1E",X"39",X"EB",X"0D",X"C0",X"EB",X"1A",X"CB",X"7F",X"C2",X"49",X"39",X"21",X"F4",X"81",X"CD",
		X"1E",X"39",X"D5",X"21",X"50",X"3B",X"CD",X"1B",X"33",X"CD",X"1B",X"33",X"E1",X"C9",X"FE",X"0A",
		X"06",X"24",X"38",X"04",X"06",X"01",X"D6",X"0A",X"70",X"CB",X"AD",X"77",X"C9",X"21",X"67",X"3B",
		X"CD",X"1B",X"33",X"21",X"80",X"99",X"36",X"FF",X"23",X"36",X"FF",X"EB",X"21",X"32",X"83",X"06",
		X"16",X"36",X"24",X"3E",X"E0",X"25",X"D7",X"10",X"F8",X"21",X"34",X"83",X"06",X"16",X"36",X"24",
		X"3E",X"E0",X"25",X"D7",X"10",X"F8",X"EB",X"C9",X"21",X"00",X"80",X"11",X"01",X"80",X"01",X"00",
		X"04",X"36",X"24",X"ED",X"B0",X"36",X"03",X"01",X"FF",X"03",X"ED",X"B0",X"3E",X"07",X"32",X"BE",
		X"99",X"C9",X"21",X"80",X"93",X"06",X"80",X"36",X"F1",X"23",X"10",X"FB",X"C9",X"21",X"E0",X"99",
		X"11",X"5E",X"83",X"0E",X"02",X"06",X"01",X"CD",X"97",X"39",X"06",X"03",X"CD",X"97",X"39",X"06",
		X"02",X"CD",X"97",X"39",X"23",X"06",X"01",X"CD",X"AA",X"39",X"CD",X"A0",X"39",X"10",X"FB",X"C9",
		X"3E",X"99",X"96",X"1F",X"1F",X"1F",X"1F",X"CD",X"AE",X"39",X"3E",X"99",X"96",X"23",X"E6",X"0F",
		X"12",X"E7",X"0D",X"C0",X"3E",X"2A",X"0E",X"04",X"12",X"E7",X"C9",X"21",X"5E",X"83",X"06",X"17",
		X"11",X"E0",X"FF",X"36",X"24",X"19",X"10",X"FB",X"C9",X"E5",X"CD",X"7D",X"39",X"21",X"84",X"03",
		X"22",X"72",X"92",X"E1",X"C1",X"C9",X"C5",X"78",X"FE",X"0F",X"28",X"ED",X"FE",X"02",X"28",X"15",
		X"FE",X"04",X"20",X"3D",X"3A",X"70",X"92",X"D6",X"01",X"30",X"02",X"3E",X"11",X"32",X"70",X"92",
		X"18",X"0A",X"C5",X"18",X"07",X"3A",X"70",X"92",X"3C",X"32",X"70",X"92",X"3A",X"70",X"92",X"FE",
		X"12",X"38",X"01",X"AF",X"32",X"70",X"92",X"E5",X"0E",X"00",X"FE",X"0A",X"38",X"03",X"0C",X"D6",
		X"0A",X"21",X"2E",X"82",X"71",X"2E",X"0E",X"77",X"21",X"47",X"3A",X"CD",X"1B",X"33",X"E1",X"C1",
		X"C9",X"3A",X"70",X"92",X"FE",X"12",X"38",X"01",X"AF",X"32",X"70",X"92",X"EB",X"CD",X"3C",X"3A",
		X"21",X"4F",X"3A",X"D7",X"6E",X"26",X"9A",X"36",X"01",X"EB",X"C1",X"C9",X"21",X"A0",X"9A",X"06",
		X"40",X"36",X"00",X"23",X"10",X"FB",X"C9",X"EE",X"82",X"05",X"1C",X"18",X"1E",X"17",X"0D",X"A1",
		X"A2",X"A3",X"A4",X"A7",X"AA",X"AB",X"AC",X"AD",X"AE",X"AF",X"B0",X"B2",X"B3",X"B4",X"B5",X"B6",
		X"B9",X"7E",X"23",X"66",X"6F",X"C3",X"1B",X"33",X"0B",X"0C",X"0D",X"0A",X"04",X"01",X"04",X"01",
		X"04",X"1C",X"01",X"24",X"03",X"01",X"03",X"01",X"03",X"1C",X"01",X"24",X"02",X"01",X"02",X"01",
		X"02",X"1C",X"01",X"24",X"02",X"03",X"02",X"03",X"02",X"1C",X"03",X"1C",X"01",X"03",X"01",X"03",
		X"01",X"24",X"03",X"1C",X"01",X"02",X"01",X"02",X"01",X"24",X"02",X"1C",X"01",X"01",X"01",X"01",
		X"01",X"24",X"01",X"24",X"FF",X"FF",X"02",X"06",X"02",X"07",X"02",X"08",X"03",X"0A",X"03",X"0C",
		X"02",X"86",X"03",X"88",X"FF",X"FF",X"03",X"0A",X"03",X"0C",X"03",X"0F",X"03",X"8A",X"03",X"8C",
		X"03",X"8F",X"03",X"FF",X"01",X"01",X"01",X"01",X"01",X"02",X"03",X"00",X"D0",X"3A",X"DA",X"3A",
		X"E6",X"82",X"07",X"1E",X"19",X"1B",X"12",X"10",X"11",X"1D",X"E6",X"82",X"07",X"1D",X"0A",X"0B",
		X"15",X"0E",X"24",X"24",X"EC",X"82",X"04",X"1B",X"0A",X"17",X"14",X"AA",X"82",X"08",X"0F",X"12",
		X"10",X"11",X"1D",X"0E",X"1B",X"1C",X"C8",X"82",X"05",X"24",X"0C",X"18",X"12",X"17",X"A8",X"81",
		X"06",X"0C",X"1B",X"0E",X"0D",X"12",X"1D",X"E8",X"82",X"12",X"0F",X"1B",X"0E",X"0E",X"24",X"19",
		X"15",X"0A",X"22",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"21",X"3B",X"39",
		X"3B",X"30",X"83",X"0A",X"01",X"1C",X"1D",X"24",X"0B",X"18",X"17",X"1E",X"1C",X"24",X"B0",X"81",
		X"08",X"00",X"00",X"00",X"00",X"24",X"19",X"1D",X"1C",X"32",X"83",X"09",X"02",X"17",X"0D",X"24",
		X"0B",X"18",X"17",X"1E",X"1C",X"B2",X"81",X"08",X"00",X"00",X"00",X"00",X"24",X"19",X"1D",X"1C",
		X"34",X"83",X"09",X"0A",X"17",X"0D",X"24",X"0E",X"1F",X"0E",X"1B",X"22",X"B4",X"81",X"08",X"00",
		X"00",X"00",X"00",X"24",X"19",X"1D",X"1C",X"30",X"83",X"16",X"0B",X"18",X"17",X"1E",X"1C",X"24",
		X"17",X"18",X"1D",X"11",X"12",X"17",X"10",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",
		X"24",X"E2",X"82",X"07",X"1B",X"0A",X"16",X"24",X"24",X"18",X"14",X"E4",X"82",X"07",X"1B",X"18",
		X"16",X"24",X"24",X"18",X"14",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"D9");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
