library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity gfx1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of gfx1 is
	type rom is array(0 to  6143) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"14",X"1C",X"7A",X"FA",X"FC",X"FC",X"FC",X"FC",X"FC",X"7A",X"7A",X"3C",X"1C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"6C",X"7C",X"7C",X"7C",X"38",X"38",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"44",X"28",X"10",X"44",X"28",X"10",
		X"02",X"22",X"31",X"1A",X"05",X"83",X"53",X"15",X"1C",X"28",X"08",X"20",X"00",X"82",X"40",X"00",
		X"04",X"70",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"08",X"68",X"80",X"90",X"30",X"18",
		X"00",X"00",X"03",X"05",X"0A",X"0D",X"17",X"0F",X"00",X"00",X"C0",X"A0",X"50",X"B0",X"E8",X"F8",
		X"15",X"13",X"0D",X"0A",X"05",X"03",X"00",X"00",X"D8",X"88",X"B0",X"50",X"A0",X"C0",X"00",X"00",
		X"82",X"C6",X"3E",X"3C",X"18",X"FE",X"FE",X"00",X"FC",X"FE",X"02",X"02",X"02",X"06",X"04",X"00",
		X"FC",X"FE",X"02",X"02",X"02",X"FE",X"FC",X"00",X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"18",X"00",X"00",X"00",
		X"00",X"00",X"00",X"5E",X"4E",X"0E",X"04",X"00",X"04",X"4E",X"1E",X"5E",X"4E",X"0E",X"04",X"00",
		X"80",X"0E",X"0E",X"1F",X"3F",X"3F",X"7F",X"7F",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"7F",X"3F",X"3F",X"1F",X"0E",X"0E",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",
		X"10",X"01",X"01",X"03",X"07",X"07",X"0F",X"0F",X"01",X"C1",X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",
		X"0F",X"0F",X"07",X"07",X"03",X"01",X"01",X"10",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",X"C1",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"2E",X"28",X"28",X"28",X"28",X"38",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"28",X"28",X"28",X"28",X"2E",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"20",X"20",X"20",X"2E",X"28",X"38",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"28",X"2E",X"20",X"20",X"20",X"38",X"00",
		X"00",X"3C",X"44",X"5A",X"BC",X"BD",X"98",X"81",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",
		X"81",X"98",X"BD",X"BC",X"5A",X"44",X"3C",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"18",X"24",X"42",X"58",X"98",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"80",
		X"80",X"80",X"98",X"58",X"42",X"24",X"18",X"00",X"80",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"43",X"07",X"3C",X"5C",X"58",X"70",X"72",X"72",X"F2",X"F2",
		X"8C",X"80",X"10",X"20",X"20",X"B0",X"94",X"00",X"72",X"70",X"78",X"7C",X"7C",X"7C",X"78",X"70",
		X"07",X"47",X"07",X"23",X"03",X"01",X"00",X"00",X"F2",X"F2",X"F2",X"F2",X"F2",X"F0",X"F8",X"3C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"0F",X"3C",X"4C",X"4C",X"FC",X"F0",X"E0",X"E6",X"E6",
		X"18",X"10",X"38",X"38",X"38",X"38",X"28",X"20",X"E0",X"E0",X"F0",X"FC",X"FC",X"FC",X"FC",X"F0",
		X"3F",X"1F",X"1F",X"0F",X"0F",X"07",X"01",X"00",X"E0",X"E6",X"E6",X"E0",X"E0",X"F0",X"FC",X"7C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"01",X"03",X"03",X"03",X"1F",X"3F",X"E4",X"24",X"24",X"CC",X"80",X"80",X"98",X"98",
		X"63",X"43",X"E3",X"E3",X"E3",X"E3",X"A3",X"83",X"80",X"C0",X"FC",X"E4",X"E4",X"E4",X"CC",X"80",
		X"FF",X"7F",X"7F",X"3F",X"3F",X"1F",X"07",X"01",X"80",X"98",X"98",X"80",X"80",X"CC",X"E4",X"E4",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"28",X"04",X"40",X"54",X"2C",X"18",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"20",X"44",X"96",X"5A",X"A6",X"BE",X"5C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"20",X"44",X"96",X"5A",X"A6",X"BE",X"5C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"04",X"56",X"A4",X"8A",X"5E",X"64",X"38",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",X"44",X"C6",X"82",X"82",X"C6",X"7C",X"38",X"00",
		X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",X"82",X"92",X"92",X"92",X"92",X"FE",X"FE",X"00",
		X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",X"00",X"82",X"82",X"FE",X"FE",X"82",X"82",X"00",
		X"00",X"02",X"02",X"02",X"02",X"FE",X"FE",X"00",X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",X"00",
		X"70",X"F8",X"88",X"88",X"88",X"FE",X"FE",X"00",X"72",X"F6",X"9E",X"8C",X"88",X"FE",X"FE",X"00",
		X"0C",X"5E",X"D2",X"92",X"92",X"F6",X"64",X"00",X"00",X"80",X"80",X"FE",X"FE",X"80",X"80",X"00",
		X"00",X"C0",X"F0",X"1E",X"1E",X"F0",X"C0",X"00",X"9E",X"9E",X"92",X"82",X"C6",X"7C",X"38",X"00",
		X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",X"80",X"90",X"90",X"90",X"90",X"FE",X"FE",X"00",
		X"00",X"42",X"22",X"36",X"1F",X"08",X"1A",X"0F",X"00",X"22",X"06",X"8C",X"28",X"80",X"D0",X"A4",
		X"3F",X"1F",X"18",X"1D",X"2D",X"33",X"01",X"00",X"F0",X"90",X"C8",X"A8",X"B8",X"44",X"C4",X"80",
		X"04",X"12",X"08",X"42",X"28",X"80",X"51",X"03",X"20",X"48",X"10",X"42",X"14",X"00",X"08",X"80",
		X"07",X"03",X"51",X"80",X"28",X"42",X"08",X"10",X"C0",X"88",X"00",X"14",X"42",X"10",X"48",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"48",X"45",X"25",X"27",X"DF",X"7E",X"7F",X"78",X"FC",X"FC",X"EE",X"46",X"56",X"02",X"56",
		X"FF",X"7E",X"F3",X"E3",X"01",X"01",X"00",X"00",X"56",X"02",X"56",X"16",X"BE",X"FC",X"FC",X"78",
		X"00",X"7E",X"42",X"42",X"42",X"42",X"7E",X"00",X"00",X"06",X"3C",X"3C",X"3C",X"3C",X"06",X"00",
		X"00",X"40",X"18",X"38",X"38",X"18",X"40",X"00",X"FF",X"FF",X"FF",X"80",X"80",X"FF",X"FF",X"FF",
		X"00",X"3F",X"7F",X"7F",X"7F",X"7F",X"3F",X"1F",X"FF",X"BE",X"BE",X"80",X"80",X"BE",X"BE",X"FF",
		X"3F",X"00",X"00",X"0C",X"0C",X"00",X"00",X"3F",X"00",X"F0",X"00",X"C6",X"C6",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"38",X"70",X"F0",X"E9",X"E1",X"E1",X"D5",X"87",
		X"87",X"D5",X"E1",X"E1",X"E9",X"F0",X"70",X"38",X"00",X"00",X"00",X"C0",X"F0",X"EB",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"38",X"78",X"41",X"63",X"F3",X"FF",X"FF",X"FF",X"40",X"E8",X"DC",X"B6",X"A0",X"C0",X"E0",X"C0",
		X"F7",X"DB",X"AB",X"AB",X"DB",X"71",X"30",X"1C",X"80",X"80",X"C0",X"E0",X"D6",X"9C",X"88",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"FC",X"1E",X"0E",X"07",X"C7",X"E7",
		X"E7",X"C7",X"07",X"0E",X"1E",X"FC",X"F8",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"18",X"3C",X"3C",X"18",X"00",X"00",X"01",X"FF",X"FF",X"01",X"01",X"FF",X"FF",X"01",
		X"0C",X"1E",X"36",X"6F",X"6B",X"23",X"27",X"4F",X"96",X"AC",X"DC",X"56",X"57",X"23",X"6B",X"5D",
		X"8F",X"87",X"CE",X"6C",X"3E",X"1E",X"16",X"0C",X"1C",X"36",X"6F",X"4B",X"47",X"AF",X"EE",X"BE",
		X"D6",X"47",X"63",X"2B",X"17",X"37",X"2E",X"2E",X"26",X"13",X"09",X"19",X"19",X"16",X"0E",X"04",
		X"7C",X"44",X"44",X"7C",X"00",X"7C",X"54",X"54",X"7C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7C",X"44",X"44",X"7C",X"00",X"7C",X"44",X"44",X"7C",X"00",X"7C",X"00",X"00",X"00",X"00",X"00",
		X"7C",X"44",X"44",X"7C",X"00",X"5C",X"54",X"54",X"74",X"00",X"7C",X"00",X"00",X"00",X"00",X"00",
		X"7C",X"44",X"44",X"7C",X"00",X"7C",X"44",X"44",X"7C",X"00",X"74",X"54",X"54",X"5C",X"00",X"00",
		X"7C",X"44",X"44",X"7C",X"00",X"5C",X"54",X"54",X"74",X"00",X"74",X"54",X"54",X"5C",X"00",X"00",
		X"7C",X"44",X"44",X"7C",X"00",X"7C",X"44",X"44",X"7C",X"00",X"7C",X"54",X"54",X"44",X"00",X"00",
		X"7C",X"44",X"44",X"7C",X"00",X"7C",X"44",X"44",X"7C",X"00",X"08",X"7C",X"08",X"78",X"00",X"00",
		X"7C",X"44",X"44",X"7C",X"00",X"7C",X"44",X"44",X"7C",X"00",X"5C",X"54",X"54",X"74",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"50",X"5A",X"40",X"60",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"01",X"04",X"04",X"04",X"0C",X"18",X"70",X"96",X"16",
		X"00",X"00",X"00",X"10",X"30",X"30",X"30",X"10",X"90",X"18",X"0C",X"3C",X"3C",X"24",X"2C",X"38",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"16",X"16",X"10",X"18",X"0C",X"04",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FE",X"BF",X"FE",X"F7",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"3E",X"3F",X"57",X"57",X"57",
		X"F7",X"57",X"46",X"06",X"06",X"06",X"06",X"00",X"00",X"06",X"06",X"06",X"06",X"46",X"57",X"F7",
		X"D7",X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"F7",X"F7",X"D6",X"D6",X"D6",X"06",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"D7",X"00",X"06",X"06",X"D6",X"D6",X"D6",X"F7",X"F7",
		X"00",X"10",X"08",X"00",X"00",X"00",X"04",X"0C",X"00",X"47",X"07",X"06",X"0F",X"17",X"13",X"09",
		X"0F",X"0C",X"04",X"00",X"00",X"00",X"04",X"00",X"AC",X"7D",X"50",X"54",X"4E",X"85",X"4A",X"47",
		X"00",X"00",X"08",X"10",X"00",X"00",X"02",X"00",X"45",X"CA",X"87",X"C3",X"76",X"7E",X"7E",X"79",
		X"00",X"00",X"00",X"00",X"20",X"10",X"00",X"00",X"35",X"34",X"0C",X"0A",X"26",X"4F",X"07",X"02",
		X"3C",X"32",X"32",X"3F",X"0F",X"07",X"67",X"67",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"F0",
		X"07",X"07",X"0F",X"3F",X"3F",X"3F",X"3F",X"0F",X"18",X"08",X"0C",X"04",X"04",X"04",X"04",X"04",
		X"07",X"67",X"67",X"07",X"07",X"0F",X"3F",X"3E",X"FC",X"18",X"18",X"30",X"F0",X"E0",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"40",X"24",X"1C",X"18",X"60",X"18",X"10",X"30",X"18",X"18",X"0C",X"0E",X"03",X"07",X"08",
		X"10",X"28",X"E8",X"54",X"54",X"28",X"88",X"CC",X"37",X"36",X"16",X"78",X"3E",X"3C",X"1C",X"14",
		X"FC",X"38",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"12",X"0C",X"00",X"00",X"00",X"00",X"00",
		X"54",X"00",X"AA",X"00",X"54",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F1",X"00",X"00",X"1F",X"1F",X"00",X"00",X"F1",X"03",X"0F",X"03",X"01",X"01",X"03",X"07",X"01",
		X"7F",X"FF",X"9F",X"FF",X"FF",X"9F",X"5F",X"FF",X"0F",X"11",X"07",X"01",X"00",X"03",X"0D",X"00",
		X"00",X"00",X"00",X"16",X"72",X"46",X"44",X"60",X"30",X"40",X"02",X"10",X"38",X"3C",X"6E",X"46",
		X"44",X"68",X"20",X"10",X"1C",X"00",X"18",X"0E",X"18",X"36",X"36",X"16",X"20",X"18",X"14",X"04",
		X"01",X"01",X"83",X"43",X"72",X"38",X"2E",X"22",X"01",X"06",X"8C",X"58",X"34",X"64",X"E8",X"E8",
		X"11",X"1D",X"3D",X"71",X"43",X"D3",X"BB",X"BD",X"F8",X"E6",X"CF",X"D9",X"D9",X"CF",X"E6",X"F2",
		X"3B",X"F1",X"19",X"8D",X"85",X"81",X"FD",X"F1",X"F3",X"F6",X"F4",X"FC",X"E6",X"CF",X"C9",X"C9",
		X"71",X"71",X"2D",X"3D",X"7E",X"C7",X"00",X"00",X"CF",X"E2",X"F2",X"FA",X"FE",X"76",X"C2",X"81",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"10",X"00",X"00",X"00",X"01",X"03",X"07",X"00",X"80",X"C0",X"E0",X"F0",X"B8",X"8C",X"80",
		X"67",X"03",X"01",X"00",X"00",X"00",X"10",X"20",X"80",X"8C",X"B8",X"F0",X"E0",X"C0",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"39",X"1D",X"1D",X"0F",X"07",X"03",X"01",X"00",X"E0",X"E0",X"E0",X"E0",X"F0",X"F8",X"F8",X"78",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",
		X"44",X"C6",X"82",X"82",X"C6",X"7C",X"38",X"00",X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",
		X"82",X"92",X"92",X"92",X"92",X"FE",X"FE",X"00",X"80",X"90",X"90",X"90",X"90",X"FE",X"FE",X"00",
		X"9E",X"9E",X"92",X"82",X"C6",X"7C",X"38",X"00",X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",
		X"00",X"82",X"82",X"FE",X"FE",X"82",X"82",X"00",X"FC",X"FE",X"02",X"02",X"02",X"06",X"04",X"00",
		X"82",X"C6",X"3E",X"3C",X"18",X"FE",X"FE",X"00",X"00",X"02",X"02",X"02",X"02",X"FE",X"FE",X"00",
		X"FE",X"FE",X"70",X"38",X"70",X"FE",X"FE",X"00",X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",
		X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",X"00",X"70",X"F8",X"88",X"88",X"88",X"FE",X"FE",X"00",
		X"7A",X"FC",X"8E",X"8A",X"82",X"FE",X"7C",X"00",X"72",X"F6",X"9E",X"8C",X"88",X"FE",X"FE",X"00",
		X"0C",X"5E",X"D2",X"92",X"92",X"F6",X"64",X"00",X"00",X"80",X"80",X"FE",X"FE",X"80",X"80",X"00",
		X"FC",X"FE",X"02",X"02",X"02",X"FE",X"FC",X"00",X"F0",X"F8",X"1C",X"0E",X"1C",X"F8",X"F0",X"00",
		X"F8",X"FE",X"1C",X"38",X"1C",X"FE",X"F8",X"00",X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",
		X"00",X"C0",X"F0",X"1E",X"1E",X"F0",X"C0",X"00",X"C2",X"E2",X"F2",X"BA",X"9E",X"8E",X"86",X"00",
		X"00",X"00",X"00",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"18",X"00",X"00",X"00",
		X"00",X"00",X"00",X"06",X"0D",X"0C",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"06",X"00",X"00",
		X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"00",X"81",X"81",X"42",X"3C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"3C",X"42",X"81",X"81",X"00",X"00",X"08",X"10",X"34",X"38",X"30",X"10",X"40",
		X"7C",X"7C",X"5C",X"7C",X"08",X"5C",X"54",X"54",X"7C",X"0C",X"06",X"04",X"04",X"08",X"00",X"00",
		X"38",X"78",X"41",X"63",X"F3",X"FF",X"FF",X"FF",X"40",X"E8",X"CC",X"B6",X"A0",X"C0",X"E0",X"C0",
		X"F7",X"DB",X"AB",X"AB",X"DB",X"71",X"30",X"1C",X"80",X"80",X"C0",X"E0",X"D6",X"9C",X"88",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"10",X"18",X"00",X"00",X"F1",X"F1",X"00",X"00",X"1F",X"0F",X"00",X"00",X"01",
		X"01",X"00",X"00",X"0F",X"1F",X"00",X"00",X"F1",X"F1",X"00",X"00",X"18",X"10",X"00",X"00",X"80",
		X"44",X"11",X"00",X"44",X"11",X"00",X"44",X"11",X"00",X"01",X"00",X"04",X"11",X"00",X"44",X"11",
		X"44",X"11",X"00",X"44",X"10",X"00",X"40",X"00",X"07",X"7F",X"0F",X"03",X"07",X"FF",X"1F",X"03",
		X"C0",X"F8",X"FF",X"E0",X"C0",X"F0",X"FE",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"7F",X"7F",X"01",X"01",X"01",X"00",X"40",X"60",X"60",X"60",X"60",X"40",X"00",
		X"11",X"86",X"1C",X"29",X"90",X"2C",X"C2",X"14",X"20",X"C6",X"88",X"32",X"64",X"11",X"14",X"CB",
		X"48",X"02",X"A8",X"18",X"B6",X"1B",X"04",X"33",X"22",X"4C",X"91",X"7A",X"B2",X"C8",X"64",X"32",
		X"58",X"2E",X"5D",X"B2",X"EC",X"E2",X"D2",X"9C",X"50",X"4D",X"49",X"26",X"60",X"74",X"D0",X"BA",
		X"B5",X"EC",X"E2",X"A0",X"53",X"44",X"20",X"08",X"00",X"82",X"00",X"81",X"30",X"0C",X"01",X"C1",
		X"11",X"B6",X"3C",X"79",X"90",X"6D",X"F6",X"1E",X"28",X"F6",X"CA",X"B2",X"74",X"71",X"34",X"CB",
		X"3A",X"6C",X"D7",X"B1",X"EC",X"E2",X"D3",X"5C",X"5A",X"4D",X"49",X"26",X"10",X"70",X"70",X"FD",
		X"F8",X"C2",X"DA",X"44",X"50",X"23",X"10",X"04",X"00",X"04",X"50",X"01",X"44",X"01",X"20",X"04",
		X"9C",X"D2",X"E2",X"EC",X"B2",X"5D",X"2E",X"58",X"BA",X"D0",X"74",X"60",X"26",X"49",X"4D",X"50",
		X"08",X"20",X"44",X"53",X"A0",X"E2",X"EC",X"B5",X"C1",X"01",X"0C",X"30",X"81",X"00",X"82",X"00",
		X"5C",X"D3",X"E2",X"EC",X"B1",X"D7",X"6C",X"3A",X"FD",X"70",X"70",X"10",X"26",X"49",X"4D",X"5A",
		X"04",X"10",X"23",X"50",X"44",X"DA",X"C2",X"F8",X"04",X"20",X"01",X"44",X"01",X"50",X"04",X"00",
		X"B2",X"57",X"AD",X"42",X"D2",X"6A",X"D4",X"33",X"3B",X"6D",X"D6",X"34",X"50",X"A2",X"6D",X"1B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"01",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"FC",X"00",X"00",X"FC",X"00",X"8C",
		X"00",X"00",X"00",X"01",X"00",X"01",X"01",X"01",X"50",X"20",X"50",X"8C",X"00",X"24",X"24",X"FC",
		X"00",X"78",X"63",X"6C",X"08",X"45",X"35",X"3A",X"00",X"DA",X"22",X"40",X"24",X"18",X"24",X"80",
		X"3A",X"35",X"45",X"08",X"6C",X"63",X"78",X"00",X"80",X"24",X"18",X"24",X"40",X"22",X"DA",X"00",
		X"00",X"00",X"00",X"30",X"78",X"F8",X"FD",X"FC",X"00",X"00",X"00",X"01",X"07",X"01",X"80",X"80",
		X"FC",X"FD",X"F8",X"78",X"30",X"00",X"00",X"00",X"80",X"80",X"01",X"07",X"01",X"00",X"00",X"00",
		X"78",X"1E",X"0F",X"1F",X"0F",X"07",X"27",X"03",X"00",X"00",X"80",X"E0",X"F9",X"FE",X"F9",X"E0",
		X"03",X"27",X"07",X"0F",X"1F",X"0F",X"1E",X"78",X"E0",X"F9",X"FE",X"F9",X"E0",X"80",X"00",X"00",
		X"0E",X"1F",X"30",X"30",X"60",X"6D",X"63",X"7C",X"09",X"1F",X"8F",X"86",X"C2",X"E2",X"52",X"62",
		X"7C",X"63",X"6D",X"60",X"30",X"30",X"1F",X"0E",X"62",X"52",X"E2",X"C2",X"86",X"8F",X"1F",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"16",X"16",X"10",X"18",X"0C",X"04",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7E",X"3C",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3C",X"7E",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"1F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"3F",X"0F",X"0F",X"0F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",X"1F",X"07",
		X"FF",X"FF",X"FE",X"FE",X"FC",X"F8",X"F0",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E0",X"F8",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"F0",X"F0",X"E0",X"E0",X"C0",X"C0",X"80",X"80",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"80",X"80",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",
		X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"07",X"03",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"07",X"03",X"01",X"01",X"03",X"07",X"0F",X"00",X"00",X"00",X"00",X"03",X"07",X"0F",X"0F",
		X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"F8",X"FC",X"FC",X"FC",X"F8",X"F0",X"C0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"C0",X"FF",X"7F",X"3F",X"1F",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"7E",X"3C",X"87",X"C7",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"CF",X"87",X"87",X"07",X"1F",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",
		X"FF",X"7F",X"00",X"00",X"00",X"7E",X"FF",X"FF",X"FF",X"FC",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"03",X"0F",X"07",X"07",X"07",X"03",X"03",X"01",X"01",
		X"03",X"07",X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FC",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FE",X"FF",X"80",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",
		X"FC",X"F8",X"F8",X"F0",X"E0",X"80",X"00",X"00",X"3F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"20",X"12",X"19",X"09",X"09",X"19",X"12",X"20",X"10",X"10",X"18",X"08",X"4C",X"46",X"23",X"10",
		X"10",X"23",X"46",X"4C",X"08",X"18",X"10",X"10",X"00",X"18",X"18",X"18",X"18",X"18",X"18",X"00",
		X"3C",X"42",X"81",X"A5",X"A5",X"99",X"42",X"3C",X"F0",X"F8",X"1C",X"0E",X"1C",X"F8",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F8",X"1C",X"0E",X"1C",X"F8",X"F0",X"00",X"FE",X"FE",X"70",X"38",X"70",X"FE",X"FE",X"00",
		X"FF",X"99",X"99",X"FF",X"FF",X"99",X"99",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"FF",X"38",X"F8",X"38",X"F8",X"3F",X"FF",X"82",X"18",X"3C",X"3C",X"3C",X"3C",X"18",X"82",
		X"54",X"DC",X"AA",X"AA",X"76",X"DC",X"AA",X"AA",X"20",X"70",X"50",X"60",X"30",X"70",X"50",X"20",
		X"22",X"88",X"00",X"22",X"88",X"00",X"22",X"88",X"07",X"1F",X"39",X"51",X"58",X"46",X"30",X"0E",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"0F",X"03",X"03",X"0F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"0F",X"03",X"FF",X"3F",X"0F",X"03",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"60",X"38",X"E0",X"30",X"8C",X"30",X"E0",X"3C",X"68",X"BD",X"B0",X"69",X"5C",X"B0",X"95",X"78",
		X"00",X"00",X"77",X"CA",X"AC",X"77",X"00",X"00",X"08",X"0E",X"7E",X"CE",X"AE",X"7E",X"0E",X"08",
		X"39",X"64",X"40",X"2D",X"2D",X"40",X"64",X"39",X"50",X"8C",X"00",X"00",X"A4",X"A4",X"A4",X"FC",
		X"00",X"00",X"FC",X"00",X"00",X"8C",X"50",X"20",X"00",X"00",X"00",X"80",X"80",X"FC",X"80",X"80",
		X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",
		X"00",X"40",X"00",X"10",X"00",X"04",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",
		X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"01",X"00",X"01",X"00",X"01",
		X"01",X"00",X"04",X"00",X"10",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"04",X"00",X"00",X"20",X"70",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"E0",X"40",
		X"10",X"38",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0E",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"70",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"70",X"20",X"00",X"00",X"00",X"00",X"00",
		X"EF",X"3F",X"0E",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0E",X"3F",X"F7",
		X"FF",X"EF",X"FD",X"BF",X"FF",X"FB",X"DF",X"FF",X"0D",X"0F",X"0F",X"0B",X"0F",X"0F",X"0D",X"0F",
		X"24",X"6A",X"D1",X"E8",X"E2",X"D4",X"68",X"24",X"04",X"14",X"1E",X"04",X"06",X"0C",X"04",X"04",
		X"00",X"60",X"F0",X"F0",X"F0",X"F0",X"60",X"00",X"04",X"08",X"04",X"04",X"00",X"04",X"04",X"02",
		X"00",X"01",X"02",X"05",X"FC",X"05",X"04",X"05",X"04",X"05",X"02",X"01",X"00",X"01",X"06",X"01",
		X"00",X"01",X"06",X"01",X"00",X"01",X"06",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"C0",X"90",X"30",X"20",
		X"00",X"00",X"26",X"7F",X"26",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"24",X"2D",X"1E",X"1C",X"1C",X"1E",X"2D",X"24",X"06",X"1F",X"1F",X"3F",X"07",X"07",X"06",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"10",X"14",X"1C",X"18",X"30",
		X"68",X"70",X"70",X"7A",X"68",X"7C",X"14",X"22",X"70",X"78",X"30",X"10",X"00",X"00",X"08",X"00",
		X"38",X"78",X"41",X"63",X"F3",X"FF",X"FF",X"FF",X"40",X"E8",X"DC",X"B6",X"A0",X"C0",X"E0",X"C0",
		X"F7",X"DB",X"AB",X"AB",X"DB",X"71",X"30",X"1C",X"80",X"80",X"C0",X"E0",X"D6",X"9C",X"88",X"40",
		X"FF",X"FF",X"3F",X"3F",X"FF",X"FF",X"FF",X"FF",X"3F",X"0F",X"80",X"80",X"F8",X"7F",X"1F",X"03",
		X"3F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"07",X"1F",X"FF",X"03",X"03",
		X"0C",X"38",X"62",X"E2",X"C3",X"00",X"20",X"30",X"80",X"80",X"80",X"84",X"CF",X"7F",X"7F",X"3F",
		X"3F",X"0F",X"8F",X"FF",X"FC",X"FC",X"F1",X"C1",X"B6",X"96",X"C7",X"63",X"79",X"E1",X"FC",X"E3",
		X"03",X"04",X"04",X"0E",X"0E",X"07",X"83",X"80",X"81",X"81",X"03",X"03",X"03",X"73",X"0F",X"FF",
		X"00",X"00",X"01",X"82",X"04",X"04",X"04",X"65",X"00",X"00",X"00",X"01",X"03",X"03",X"03",X"03",
		X"00",X"08",X"10",X"34",X"38",X"30",X"10",X"40",X"7C",X"7C",X"5C",X"7C",X"08",X"5C",X"54",X"54",
		X"7C",X"0C",X"06",X"04",X"04",X"08",X"00",X"00",X"00",X"08",X"10",X"34",X"38",X"50",X"10",X"40",
		X"7C",X"7C",X"5C",X"7C",X"08",X"7C",X"54",X"54",X"7C",X"0C",X"06",X"04",X"04",X"08",X"00",X"00",
		X"7C",X"44",X"44",X"7C",X"00",X"7C",X"54",X"54",X"7C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7C",X"44",X"44",X"7C",X"00",X"7C",X"44",X"44",X"7C",X"00",X"7C",X"00",X"00",X"00",X"00",X"00",
		X"7C",X"44",X"44",X"7C",X"00",X"5C",X"54",X"54",X"74",X"00",X"74",X"00",X"00",X"00",X"00",X"00",
		X"7C",X"44",X"44",X"7C",X"00",X"7C",X"44",X"44",X"7C",X"00",X"74",X"54",X"54",X"5C",X"00",X"00",
		X"7C",X"44",X"44",X"7C",X"00",X"5C",X"54",X"54",X"74",X"00",X"74",X"54",X"54",X"5C",X"00",X"00",
		X"7C",X"44",X"44",X"7C",X"00",X"7C",X"44",X"44",X"7C",X"00",X"7C",X"54",X"54",X"44",X"00",X"00",
		X"7C",X"44",X"44",X"7C",X"00",X"7C",X"44",X"44",X"7C",X"00",X"08",X"7C",X"08",X"78",X"00",X"00",
		X"7C",X"44",X"44",X"7C",X"00",X"7C",X"44",X"44",X"7C",X"00",X"5C",X"54",X"54",X"74",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"50",X"5A",X"40",X"60",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"01",X"04",X"04",X"04",X"0C",X"18",X"70",X"96",X"16",
		X"00",X"00",X"00",X"10",X"30",X"30",X"30",X"10",X"90",X"18",X"0C",X"3C",X"3C",X"24",X"2C",X"38",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"16",X"16",X"10",X"18",X"0C",X"04",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"10",X"18",X"00",X"00",X"F1",X"F1",X"00",X"00",X"1F",X"0F",X"00",X"00",X"01",
		X"01",X"00",X"00",X"0F",X"1F",X"00",X"00",X"F1",X"F1",X"00",X"00",X"18",X"10",X"00",X"00",X"80",
		X"44",X"11",X"00",X"44",X"11",X"00",X"44",X"11",X"00",X"01",X"00",X"04",X"11",X"00",X"44",X"11",
		X"44",X"11",X"00",X"44",X"10",X"00",X"40",X"00",X"07",X"7F",X"0F",X"03",X"07",X"FF",X"1F",X"03",
		X"C0",X"F8",X"FF",X"E0",X"C0",X"F0",X"FE",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"7F",X"7F",X"01",X"01",X"01",X"00",X"40",X"60",X"60",X"60",X"60",X"40",X"00",
		X"11",X"86",X"1C",X"29",X"90",X"2C",X"C2",X"14",X"20",X"C6",X"88",X"32",X"64",X"11",X"14",X"CB",
		X"48",X"02",X"A8",X"18",X"B6",X"1B",X"04",X"33",X"22",X"4C",X"91",X"7A",X"B2",X"C8",X"64",X"32",
		X"58",X"2E",X"5D",X"B2",X"EC",X"E2",X"D2",X"9C",X"50",X"4D",X"49",X"26",X"60",X"74",X"D0",X"BA",
		X"B5",X"EC",X"E2",X"A0",X"53",X"44",X"20",X"08",X"00",X"82",X"00",X"81",X"30",X"0C",X"01",X"C1",
		X"11",X"B6",X"3C",X"79",X"90",X"6D",X"F6",X"1E",X"28",X"F6",X"CA",X"B2",X"74",X"71",X"34",X"CB",
		X"3A",X"6C",X"D7",X"B1",X"EC",X"E2",X"D3",X"5C",X"5A",X"4D",X"49",X"26",X"10",X"70",X"70",X"FD",
		X"F8",X"C2",X"DA",X"44",X"50",X"23",X"10",X"04",X"00",X"04",X"50",X"01",X"44",X"01",X"20",X"04",
		X"9C",X"D2",X"E2",X"EC",X"B2",X"5D",X"2E",X"58",X"BA",X"D0",X"74",X"60",X"26",X"49",X"4D",X"50",
		X"08",X"20",X"44",X"53",X"A0",X"E2",X"EC",X"B5",X"C1",X"01",X"0C",X"30",X"81",X"00",X"82",X"00",
		X"5C",X"D3",X"E2",X"EC",X"B1",X"D7",X"6C",X"3A",X"FD",X"70",X"70",X"10",X"26",X"49",X"4D",X"5A",
		X"04",X"10",X"23",X"50",X"44",X"DA",X"C2",X"F8",X"04",X"20",X"01",X"44",X"01",X"50",X"04",X"00",
		X"B2",X"57",X"AD",X"42",X"D2",X"6A",X"D4",X"33",X"3B",X"6D",X"D6",X"34",X"50",X"A2",X"6D",X"1B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"01",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"FC",X"00",X"00",X"FC",X"00",X"8C",
		X"00",X"00",X"00",X"01",X"00",X"01",X"01",X"01",X"50",X"20",X"50",X"8C",X"00",X"24",X"24",X"FC",
		X"00",X"78",X"63",X"6C",X"08",X"45",X"35",X"3A",X"00",X"DA",X"22",X"40",X"24",X"18",X"24",X"80",
		X"3A",X"35",X"45",X"08",X"6C",X"63",X"78",X"00",X"80",X"24",X"18",X"24",X"40",X"22",X"DA",X"00",
		X"00",X"00",X"01",X"32",X"7A",X"F8",X"FE",X"FE",X"01",X"23",X"C5",X"24",X"04",X"A8",X"AC",X"54",
		X"FE",X"FE",X"F8",X"7A",X"32",X"01",X"00",X"00",X"54",X"AC",X"A8",X"04",X"24",X"C5",X"23",X"01",
		X"00",X"00",X"03",X"0F",X"1F",X"07",X"27",X"03",X"00",X"F8",X"E0",X"C0",X"E4",X"F8",X"E4",X"C0",
		X"03",X"27",X"07",X"1F",X"0F",X"03",X"00",X"00",X"C0",X"E4",X"F8",X"E4",X"C0",X"E0",X"F8",X"00",
		X"DC",X"66",X"33",X"6F",X"C5",X"75",X"7B",X"7C",X"19",X"6F",X"1F",X"06",X"82",X"82",X"46",X"02",
		X"7C",X"67",X"75",X"D1",X"6B",X"EB",X"76",X"BC",X"02",X"46",X"82",X"82",X"06",X"1F",X"6F",X"19",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"16",X"16",X"10",X"18",X"0C",X"04",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7C",X"7E",X"75",X"2D",X"2D",X"11",X"0D",X"02",X"FC",X"FA",X"F5",X"ED",X"ED",X"F5",X"FA",X"FC",
		X"02",X"0D",X"11",X"2D",X"2D",X"75",X"7A",X"7C",X"13",X"4F",X"3C",X"F2",X"C8",X"20",X"00",X"00",
		X"00",X"00",X"20",X"C8",X"F2",X"3C",X"4F",X"13",X"BB",X"EE",X"44",X"00",X"00",X"44",X"EE",X"BB",
		X"01",X"05",X"02",X"0A",X"15",X"4C",X"38",X"E4",X"E4",X"38",X"4C",X"15",X"0A",X"02",X"05",X"01",
		X"00",X"00",X"01",X"00",X"00",X"01",X"02",X"07",X"04",X"88",X"B0",X"00",X"00",X"68",X"94",X"80",
		X"07",X"02",X"01",X"00",X"00",X"01",X"00",X"00",X"80",X"94",X"68",X"00",X"00",X"B0",X"88",X"04",
		X"40",X"11",X"04",X"10",X"00",X"40",X"00",X"00",X"01",X"03",X"47",X"1F",X"07",X"03",X"27",X"09",
		X"E0",X"A0",X"50",X"50",X"48",X"24",X"1A",X"07",X"E0",X"B8",X"CC",X"F3",X"E6",X"CF",X"9B",X"F3",
		X"07",X"1E",X"24",X"48",X"48",X"5C",X"BC",X"EC",X"00",X"00",X"00",X"00",X"00",X"7F",X"04",X"7F",
		X"E7",X"77",X"36",X"1A",X"0A",X"06",X"02",X"01",X"FF",X"BE",X"BE",X"FE",X"FF",X"BF",X"BE",X"FE",
		X"01",X"02",X"06",X"0A",X"1A",X"36",X"77",X"E7",X"FF",X"5F",X"4E",X"0E",X"0C",X"06",X"06",X"01",
		X"FF",X"FF",X"FE",X"FE",X"FC",X"FE",X"FE",X"FF",X"01",X"05",X"06",X"0E",X"0C",X"4E",X"5E",X"FF",
		X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"01",X"01",X"01",X"00",X"00",X"41",X"01",X"00",X"E0",X"A0",X"B0",X"F0",X"60",X"60",X"20",X"00",
		X"00",X"00",X"00",X"06",X"00",X"03",X"00",X"01",X"00",X"00",X"00",X"60",X"00",X"C0",X"00",X"80",
		X"00",X"03",X"00",X"07",X"00",X"07",X"00",X"01",X"00",X"C0",X"00",X"E0",X"00",X"E0",X"00",X"80",
		X"FF",X"FF",X"7E",X"5C",X"7E",X"5C",X"5C",X"5C",X"03",X"FD",X"13",X"E0",X"C0",X"40",X"80",X"80",
		X"7F",X"7F",X"5D",X"5E",X"5E",X"5E",X"5E",X"7E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"02",X"02",X"04",X"02",X"02",X"01",X"01",X"01",X"02",X"04",X"18",X"04",X"02",X"01",
		X"7C",X"44",X"44",X"7C",X"00",X"7C",X"54",X"54",X"7C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7C",X"44",X"44",X"7C",X"00",X"7C",X"44",X"44",X"7C",X"00",X"7C",X"00",X"00",X"00",X"00",X"00",
		X"7C",X"44",X"44",X"7C",X"00",X"5C",X"54",X"54",X"74",X"00",X"7C",X"00",X"00",X"00",X"00",X"00",
		X"7C",X"44",X"44",X"7C",X"00",X"7C",X"44",X"44",X"7C",X"00",X"74",X"54",X"54",X"5C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"81",X"42",X"24",X"00",X"00",X"24",X"42",X"81",
		X"18",X"18",X"04",X"03",X"00",X"0C",X"0E",X"0F",X"30",X"70",X"78",X"78",X"3C",X"0E",X"00",X"00",
		X"07",X"41",X"60",X"14",X"00",X"00",X"0E",X"1C",X"00",X"80",X"30",X"00",X"00",X"C0",X"00",X"00",
		X"38",X"38",X"31",X"02",X"00",X"0C",X"18",X"18",X"00",X"00",X"0F",X"3C",X"78",X"78",X"70",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"18",X"18",X"04",X"03",X"00",X"0C",X"0E",X"0F",X"30",X"70",X"78",X"78",X"3C",X"0E",X"00",X"00",
		X"07",X"41",X"60",X"14",X"00",X"00",X"0E",X"1C",X"00",X"80",X"30",X"00",X"00",X"C0",X"00",X"00",
		X"38",X"38",X"31",X"02",X"00",X"0C",X"18",X"18",X"00",X"00",X"0F",X"3C",X"78",X"78",X"70",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"64",X"D0",X"00",X"2F",X"CF",X"8F",X"63",X"42",X"5A",X"5A",X"5A",X"EA",X"E8",X"F0",X"F0",
		X"00",X"00",X"10",X"40",X"00",X"00",X"00",X"00",X"E0",X"00",X"0C",X"12",X"02",X"10",X"05",X"10",
		X"0C",X"04",X"40",X"40",X"8F",X"2F",X"0F",X"83",X"42",X"5A",X"5A",X"5A",X"EA",X"E8",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"08",X"10",X"10",X"02",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"06",X"06",X"05",X"06",X"06",X"0F",X"37",
		X"BF",X"7E",X"7E",X"9D",X"06",X"06",X"07",X"07",X"0F",X"0E",X"0E",X"0D",X"0E",X"0C",X"08",X"08",
		X"24",X"00",X"24",X"18",X"00",X"3C",X"C3",X"7E",X"00",X"00",X"00",X"00",X"24",X"00",X"24",X"18",
		X"3C",X"3C",X"3C",X"18",X"00",X"00",X"00",X"00",X"00",X"3C",X"C3",X"7E",X"3C",X"3C",X"3C",X"18",
		X"01",X"08",X"84",X"B2",X"58",X"6C",X"F4",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"08",
		X"F6",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"84",X"B2",X"58",X"6C",X"F4",X"F8",X"F6",X"60",
		X"00",X"00",X"02",X"01",X"00",X"00",X"01",X"01",X"00",X"08",X"38",X"79",X"FF",X"BC",X"9C",X"DC",
		X"01",X"01",X"00",X"00",X"01",X"02",X"00",X"00",X"DC",X"9C",X"BC",X"FF",X"79",X"38",X"08",X"00",
		X"09",X"A0",X"02",X"50",X"04",X"21",X"88",X"22",X"00",X"20",X"04",X"10",X"02",X"40",X"08",X"00",
		X"00",X"00",X"08",X"00",X"00",X"20",X"02",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",
		X"01",X"01",X"02",X"02",X"04",X"02",X"02",X"01",X"01",X"01",X"02",X"04",X"18",X"04",X"02",X"01",
		X"0C",X"1E",X"36",X"6F",X"6B",X"23",X"27",X"4F",X"96",X"AC",X"DC",X"56",X"57",X"23",X"6B",X"5D",
		X"8F",X"87",X"CE",X"6C",X"3E",X"1E",X"16",X"0C",X"1C",X"36",X"6F",X"4B",X"47",X"AF",X"EE",X"BE",
		X"D6",X"47",X"63",X"2B",X"17",X"37",X"2E",X"2E",X"26",X"13",X"09",X"19",X"19",X"16",X"0E",X"04",
		X"00",X"08",X"0C",X"FE",X"FF",X"FE",X"0C",X"08",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"F0",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"FE",X"FF",X"7F",X"3F",X"1F",X"0E",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C6",X"44",X"44",X"28",X"28",X"44",X"44",X"28",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"28",X"44",X"44",X"44",X"00",X"0C",X"00",X"00",
		X"00",X"00",X"20",X"7F",X"C7",X"7F",X"20",X"00",X"00",X"00",X"00",X"82",X"C4",X"82",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"38",X"00",X"00",X"00",X"00",X"00",X"CA",X"10",X"15",X"10",X"CA",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
