library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity snd_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of snd_rom is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"F3",X"ED",X"56",X"31",X"00",X"84",X"C3",X"7E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"38",X"30",X"48",
		X"2C",X"31",X"33",X"48",X"2C",X"30",X"2C",X"30",X"F5",X"3E",X"01",X"32",X"10",X"80",X"F1",X"FB",
		X"C9",X"44",X"45",X"46",X"57",X"09",X"54",X"41",X"42",X"30",X"30",X"0D",X"0A",X"09",X"44",X"45",
		X"46",X"42",X"09",X"30",X"2C",X"46",X"4C",X"47",X"56",X"4F",X"4C",X"2C",X"30",X"2C",X"30",X"0D",
		X"0A",X"0D",X"0A",X"0D",X"0A",X"54",X"F5",X"E5",X"3A",X"00",X"E0",X"2A",X"11",X"80",X"77",X"23",
		X"CB",X"65",X"28",X"03",X"21",X"00",X"80",X"22",X"11",X"80",X"E1",X"F1",X"ED",X"45",X"CD",X"98",
		X"04",X"21",X"00",X"80",X"11",X"01",X"80",X"01",X"FF",X"07",X"36",X"00",X"ED",X"B0",X"21",X"12",
		X"80",X"36",X"80",X"21",X"00",X"80",X"11",X"01",X"80",X"01",X"0F",X"00",X"36",X"80",X"ED",X"B0",
		X"FB",X"CD",X"B3",X"04",X"3A",X"10",X"80",X"A7",X"28",X"F7",X"AF",X"32",X"10",X"80",X"DD",X"21",
		X"30",X"80",X"06",X"10",X"C5",X"DD",X"CB",X"00",X"7E",X"C4",X"C7",X"00",X"11",X"20",X"00",X"DD",
		X"19",X"C1",X"10",X"F0",X"C3",X"A1",X"00",X"DD",X"5E",X"03",X"DD",X"56",X"04",X"13",X"DD",X"73",
		X"03",X"DD",X"72",X"04",X"DD",X"6E",X"05",X"DD",X"66",X"06",X"B7",X"ED",X"52",X"CC",X"4D",X"02",
		X"DD",X"CB",X"03",X"46",X"C0",X"DD",X"5E",X"11",X"DD",X"56",X"12",X"7B",X"B2",X"20",X"07",X"DD",
		X"36",X"17",X"0F",X"C3",X"C2",X"01",X"DD",X"CB",X"00",X"6E",X"20",X"33",X"DD",X"7E",X"0B",X"B7",
		X"20",X"08",X"DD",X"73",X"13",X"DD",X"72",X"14",X"18",X"59",X"3D",X"21",X"79",X"07",X"23",X"DD",
		X"4E",X"0E",X"06",X"00",X"09",X"09",X"4E",X"23",X"66",X"69",X"0E",X"04",X"09",X"4E",X"23",X"66",
		X"69",X"4F",X"06",X"00",X"09",X"09",X"7E",X"23",X"66",X"6F",X"CD",X"1A",X"02",X"18",X"34",X"D5",
		X"DD",X"6E",X"15",X"DD",X"66",X"16",X"B7",X"ED",X"52",X"F5",X"7D",X"F2",X"40",X"01",X"ED",X"44",
		X"67",X"DD",X"5E",X"03",X"CD",X"5A",X"07",X"DD",X"5E",X"05",X"CD",X"66",X"07",X"5F",X"16",X"00",
		X"F1",X"7B",X"F2",X"5B",X"01",X"ED",X"44",X"28",X"02",X"15",X"5F",X"E1",X"19",X"DD",X"75",X"13",
		X"DD",X"74",X"14",X"DD",X"7E",X"0C",X"B7",X"20",X"0B",X"DD",X"7E",X"0D",X"2F",X"E6",X"0F",X"DD",
		X"77",X"17",X"18",X"23",X"3D",X"21",X"79",X"07",X"23",X"DD",X"4E",X"0E",X"06",X"00",X"09",X"09",
		X"4E",X"23",X"66",X"69",X"0E",X"02",X"09",X"4E",X"23",X"66",X"69",X"4F",X"06",X"00",X"09",X"09",
		X"7E",X"23",X"66",X"6F",X"CD",X"E0",X"01",X"DD",X"CB",X"00",X"76",X"20",X"25",X"DD",X"7E",X"01",
		X"E6",X"0F",X"4F",X"06",X"00",X"21",X"D5",X"01",X"09",X"4E",X"DD",X"7E",X"13",X"E6",X"0F",X"B1",
		X"CD",X"5C",X"04",X"DD",X"7E",X"13",X"E6",X"F0",X"DD",X"B6",X"14",X"0F",X"0F",X"0F",X"0F",X"CD",
		X"5C",X"04",X"DD",X"7E",X"01",X"E6",X"0F",X"4F",X"06",X"00",X"21",X"D9",X"01",X"09",X"7E",X"DD",
		X"B6",X"17",X"C3",X"5C",X"04",X"80",X"A0",X"C0",X"C0",X"90",X"B0",X"D0",X"F0",X"DD",X"77",X"0F",
		X"E5",X"DD",X"7E",X"0F",X"CB",X"3F",X"F5",X"4F",X"06",X"00",X"09",X"F1",X"7E",X"E1",X"38",X"14",
		X"0F",X"0F",X"0F",X"0F",X"B7",X"28",X"E6",X"FE",X"10",X"20",X"05",X"DD",X"35",X"0F",X"18",X"E0",
		X"FE",X"20",X"28",X"0B",X"DD",X"34",X"0F",X"F6",X"F0",X"DD",X"86",X"0D",X"3C",X"38",X"01",X"AF",
		X"2F",X"E6",X"0F",X"DD",X"77",X"17",X"C9",X"DD",X"77",X"10",X"E5",X"DD",X"7E",X"10",X"CB",X"3F",
		X"F5",X"4F",X"06",X"00",X"09",X"F1",X"7E",X"E1",X"38",X"11",X"0F",X"0F",X"0F",X"0F",X"B7",X"CA",
		X"17",X"02",X"FE",X"10",X"20",X"05",X"DD",X"35",X"10",X"18",X"DF",X"DD",X"34",X"10",X"2F",X"E6",
		X"0F",X"6F",X"26",X"00",X"EB",X"19",X"DD",X"75",X"13",X"DD",X"74",X"14",X"C9",X"DD",X"5E",X"07",
		X"DD",X"56",X"08",X"1A",X"13",X"B7",X"FA",X"D2",X"02",X"DD",X"CB",X"00",X"5E",X"20",X"59",X"B7",
		X"28",X"03",X"DD",X"86",X"09",X"21",X"C6",X"06",X"4F",X"06",X"00",X"09",X"09",X"7E",X"DD",X"77",
		X"11",X"23",X"7E",X"DD",X"77",X"12",X"DD",X"CB",X"00",X"6E",X"28",X"16",X"1A",X"13",X"DD",X"86",
		X"09",X"21",X"C6",X"06",X"4F",X"06",X"00",X"09",X"09",X"7E",X"DD",X"77",X"15",X"23",X"7E",X"DD",
		X"77",X"16",X"D5",X"1A",X"67",X"DD",X"5E",X"02",X"CD",X"5A",X"07",X"D1",X"DD",X"75",X"05",X"DD",
		X"74",X"06",X"AF",X"DD",X"77",X"0F",X"DD",X"77",X"10",X"13",X"DD",X"73",X"07",X"DD",X"72",X"08",
		X"AF",X"DD",X"77",X"03",X"DD",X"77",X"04",X"C9",X"DD",X"77",X"12",X"1A",X"13",X"DD",X"77",X"11",
		X"DD",X"CB",X"00",X"6E",X"28",X"CC",X"1A",X"13",X"DD",X"77",X"16",X"1A",X"13",X"DD",X"77",X"15",
		X"18",X"C0",X"21",X"E5",X"02",X"E5",X"E6",X"3F",X"21",X"E9",X"02",X"4F",X"06",X"00",X"09",X"09",
		X"7E",X"23",X"66",X"6F",X"E9",X"13",X"C3",X"53",X"02",X"C4",X"03",X"1D",X"03",X"22",X"03",X"37",
		X"03",X"E9",X"03",X"4B",X"03",X"62",X"03",X"67",X"03",X"72",X"03",X"8D",X"03",X"6C",X"03",X"A0",
		X"03",X"A8",X"03",X"C0",X"03",X"C6",X"03",X"CC",X"03",X"D2",X"03",X"D8",X"03",X"E0",X"03",X"F3",
		X"03",X"00",X"04",X"15",X"04",X"1D",X"04",X"25",X"04",X"34",X"04",X"45",X"04",X"1A",X"DD",X"77",
		X"02",X"C9",X"1A",X"DD",X"77",X"0D",X"C9",X"0F",X"0E",X"0D",X"0C",X"0B",X"0A",X"09",X"07",X"08",
		X"06",X"05",X"04",X"03",X"02",X"01",X"00",X"1A",X"D5",X"5F",X"DD",X"66",X"02",X"CD",X"5A",X"07",
		X"DD",X"75",X"03",X"DD",X"74",X"04",X"D1",X"E1",X"C3",X"A9",X"02",X"1A",X"F6",X"E0",X"F5",X"CD",
		X"5C",X"04",X"F1",X"F6",X"FC",X"3C",X"20",X"05",X"DD",X"CB",X"00",X"B6",X"C9",X"DD",X"CB",X"00",
		X"F6",X"C9",X"1A",X"DD",X"77",X"0C",X"C9",X"1A",X"DD",X"77",X"0B",X"C9",X"EB",X"5E",X"23",X"56",
		X"1B",X"C9",X"1A",X"4F",X"13",X"1A",X"47",X"C5",X"DD",X"E5",X"E1",X"DD",X"35",X"0A",X"DD",X"4E",
		X"0A",X"DD",X"35",X"0A",X"06",X"00",X"09",X"72",X"2B",X"73",X"D1",X"1B",X"C9",X"DD",X"E5",X"E1",
		X"DD",X"4E",X"0A",X"06",X"00",X"09",X"5E",X"23",X"56",X"DD",X"34",X"0A",X"DD",X"34",X"0A",X"C9",
		X"1A",X"DD",X"86",X"09",X"DD",X"77",X"09",X"C9",X"1A",X"13",X"C6",X"18",X"4F",X"06",X"00",X"DD",
		X"E5",X"E1",X"09",X"7E",X"B7",X"20",X"02",X"1A",X"77",X"13",X"35",X"C2",X"6C",X"03",X"13",X"C9",
		X"DD",X"CB",X"00",X"EE",X"1B",X"C9",X"DD",X"CB",X"00",X"AE",X"1B",X"C9",X"DD",X"CB",X"00",X"DE",
		X"1B",X"C9",X"DD",X"CB",X"00",X"9E",X"1B",X"C9",X"1A",X"DD",X"B6",X"00",X"DD",X"77",X"00",X"C9",
		X"1A",X"2F",X"DD",X"A6",X"00",X"DD",X"77",X"00",X"C9",X"CD",X"4D",X"04",X"DD",X"36",X"00",X"00",
		X"E1",X"E1",X"C9",X"21",X"20",X"80",X"CB",X"96",X"21",X"90",X"80",X"CB",X"96",X"C3",X"E9",X"03",
		X"21",X"20",X"80",X"36",X"00",X"06",X"04",X"11",X"20",X"00",X"21",X"30",X"80",X"CB",X"96",X"19",
		X"10",X"FB",X"C3",X"E9",X"03",X"21",X"90",X"80",X"CB",X"96",X"C3",X"E9",X"03",X"21",X"30",X"80",
		X"CB",X"96",X"C3",X"E9",X"03",X"21",X"20",X"80",X"CB",X"9E",X"CB",X"96",X"21",X"90",X"80",X"CB",
		X"96",X"C3",X"E9",X"03",X"21",X"20",X"80",X"CB",X"A6",X"CB",X"9E",X"CB",X"96",X"21",X"90",X"80",
		X"CB",X"96",X"C3",X"E9",X"03",X"21",X"70",X"80",X"CB",X"96",X"C3",X"E9",X"03",X"DD",X"7E",X"01",
		X"E6",X"0F",X"4F",X"06",X"00",X"21",X"D9",X"01",X"09",X"7E",X"F6",X"0F",X"DD",X"CB",X"00",X"56",
		X"C0",X"ED",X"47",X"DD",X"7E",X"01",X"E6",X"F0",X"FE",X"10",X"28",X"06",X"ED",X"57",X"32",X"00",
		X"C0",X"C9",X"ED",X"57",X"32",X"00",X"A0",X"C9",X"E5",X"21",X"00",X"80",X"11",X"01",X"80",X"01",
		X"0F",X"00",X"36",X"80",X"ED",X"B0",X"CD",X"8B",X"04",X"E1",X"C9",X"21",X"30",X"80",X"11",X"31",
		X"80",X"01",X"FF",X"01",X"36",X"00",X"ED",X"B0",X"21",X"AF",X"04",X"11",X"00",X"A0",X"01",X"04",
		X"00",X"ED",X"B0",X"21",X"AF",X"04",X"11",X"00",X"C0",X"01",X"04",X"00",X"ED",X"B0",X"C9",X"9F",
		X"BF",X"DF",X"FF",X"06",X"10",X"21",X"00",X"80",X"7E",X"A7",X"28",X"BC",X"FE",X"80",X"28",X"09",
		X"36",X"80",X"C5",X"E5",X"CD",X"CD",X"04",X"E1",X"C1",X"23",X"10",X"EC",X"C9",X"21",X"F4",X"04",
		X"01",X"13",X"00",X"ED",X"B9",X"C0",X"21",X"F5",X"04",X"09",X"09",X"7E",X"23",X"66",X"6F",X"79",
		X"08",X"E9",X"81",X"82",X"83",X"84",X"85",X"86",X"87",X"88",X"89",X"8A",X"8B",X"8C",X"8D",X"8E",
		X"8F",X"90",X"91",X"92",X"93",X"1B",X"05",X"2F",X"05",X"43",X"05",X"6E",X"05",X"57",X"05",X"8F",
		X"05",X"A3",X"05",X"B7",X"05",X"D0",X"05",X"E4",X"05",X"0B",X"06",X"24",X"06",X"25",X"06",X"26",
		X"06",X"37",X"06",X"48",X"06",X"5F",X"06",X"78",X"06",X"79",X"06",X"CD",X"8B",X"04",X"21",X"20",
		X"80",X"36",X"00",X"23",X"36",X"00",X"21",X"A1",X"07",X"11",X"30",X"80",X"C3",X"A4",X"06",X"CD",
		X"8B",X"04",X"21",X"20",X"80",X"36",X"00",X"23",X"36",X"00",X"21",X"D9",X"08",X"11",X"30",X"80",
		X"C3",X"A4",X"06",X"CD",X"8B",X"04",X"21",X"20",X"80",X"36",X"00",X"23",X"36",X"00",X"21",X"95",
		X"0C",X"11",X"30",X"80",X"C3",X"A4",X"06",X"21",X"20",X"80",X"3A",X"20",X"80",X"E6",X"C0",X"C0",
		X"CB",X"EE",X"CD",X"94",X"06",X"21",X"A7",X"10",X"11",X"30",X"81",X"C3",X"A4",X"06",X"3A",X"21",
		X"80",X"CB",X"7F",X"C2",X"EA",X"05",X"21",X"20",X"80",X"3A",X"20",X"80",X"E6",X"F8",X"C0",X"CB",
		X"D6",X"21",X"90",X"80",X"CB",X"D6",X"21",X"EB",X"0F",X"11",X"30",X"81",X"C3",X"A4",X"06",X"CD",
		X"8B",X"04",X"21",X"20",X"80",X"36",X"00",X"23",X"36",X"00",X"21",X"F2",X"10",X"11",X"30",X"80",
		X"C3",X"A4",X"06",X"CD",X"8B",X"04",X"21",X"20",X"80",X"36",X"00",X"23",X"36",X"00",X"21",X"10",
		X"12",X"11",X"30",X"80",X"C3",X"A4",X"06",X"21",X"21",X"80",X"CB",X"FE",X"3A",X"20",X"80",X"E6",
		X"FC",X"C0",X"21",X"90",X"80",X"CB",X"D6",X"21",X"2C",X"13",X"11",X"30",X"81",X"C3",X"A4",X"06",
		X"3A",X"20",X"80",X"E6",X"E0",X"C0",X"21",X"30",X"80",X"CB",X"D6",X"21",X"A1",X"13",X"11",X"B0",
		X"81",X"C3",X"A4",X"06",X"21",X"21",X"80",X"CB",X"7E",X"C8",X"21",X"21",X"80",X"CB",X"BE",X"21",
		X"20",X"80",X"3A",X"20",X"80",X"E6",X"F8",X"C0",X"CB",X"D6",X"21",X"90",X"80",X"CB",X"D6",X"21",
		X"25",X"14",X"11",X"30",X"81",X"3E",X"09",X"08",X"C3",X"A4",X"06",X"21",X"20",X"80",X"3A",X"20",
		X"80",X"E6",X"F0",X"C0",X"CB",X"DE",X"21",X"90",X"80",X"CB",X"D6",X"21",X"39",X"15",X"11",X"30",
		X"81",X"C3",X"A4",X"06",X"C9",X"C9",X"CD",X"8B",X"04",X"21",X"20",X"80",X"36",X"00",X"21",X"1F",
		X"16",X"11",X"30",X"80",X"C3",X"A4",X"06",X"21",X"20",X"80",X"CB",X"FE",X"CD",X"94",X"06",X"21",
		X"AE",X"16",X"11",X"30",X"81",X"C3",X"A4",X"06",X"21",X"20",X"80",X"3A",X"20",X"80",X"E6",X"80",
		X"C0",X"CB",X"F6",X"CD",X"94",X"06",X"21",X"29",X"17",X"11",X"30",X"81",X"C3",X"A4",X"06",X"21",
		X"20",X"80",X"3A",X"20",X"80",X"E6",X"E0",X"C0",X"CB",X"CE",X"21",X"90",X"80",X"CB",X"D6",X"21",
		X"D2",X"17",X"11",X"30",X"81",X"C3",X"A4",X"06",X"C9",X"21",X"20",X"80",X"3A",X"20",X"80",X"E6",
		X"E0",X"C0",X"21",X"70",X"80",X"CB",X"D6",X"21",X"A3",X"18",X"11",X"F0",X"81",X"C3",X"A4",X"06",
		X"06",X"04",X"18",X"02",X"06",X"10",X"11",X"20",X"00",X"21",X"30",X"80",X"CB",X"D6",X"19",X"10",
		X"FB",X"C3",X"98",X"04",X"7E",X"23",X"66",X"6F",X"46",X"23",X"C5",X"7E",X"23",X"E5",X"66",X"6F",
		X"01",X"0E",X"00",X"ED",X"B0",X"08",X"12",X"08",X"13",X"AF",X"06",X"11",X"12",X"13",X"10",X"FC",
		X"E1",X"23",X"C1",X"10",X"E5",X"C9",X"00",X"00",X"FF",X"03",X"C7",X"03",X"90",X"03",X"5D",X"03",
		X"2D",X"03",X"FF",X"02",X"D4",X"02",X"AB",X"02",X"85",X"02",X"61",X"02",X"3F",X"02",X"1E",X"02",
		X"00",X"02",X"E3",X"01",X"C8",X"01",X"AF",X"01",X"96",X"01",X"80",X"01",X"6A",X"01",X"56",X"01",
		X"43",X"01",X"30",X"01",X"1F",X"01",X"0F",X"01",X"00",X"01",X"F2",X"00",X"E4",X"00",X"D7",X"00",
		X"CB",X"00",X"C0",X"00",X"B5",X"00",X"AB",X"00",X"A1",X"00",X"98",X"00",X"90",X"00",X"88",X"00",
		X"80",X"00",X"79",X"00",X"72",X"00",X"6C",X"00",X"66",X"00",X"60",X"00",X"5B",X"00",X"55",X"00",
		X"51",X"00",X"4C",X"00",X"48",X"00",X"44",X"00",X"40",X"00",X"3C",X"00",X"39",X"00",X"36",X"00",
		X"33",X"00",X"30",X"00",X"2D",X"00",X"2B",X"00",X"28",X"00",X"26",X"00",X"24",X"00",X"22",X"00",
		X"20",X"00",X"1E",X"00",X"1C",X"00",X"1B",X"00",X"19",X"00",X"18",X"00",X"16",X"00",X"15",X"00",
		X"13",X"00",X"12",X"00",X"11",X"00",X"10",X"00",X"0F",X"00",X"16",X"00",X"6A",X"06",X"08",X"29",
		X"30",X"01",X"19",X"10",X"FA",X"C9",X"06",X"08",X"ED",X"6A",X"7C",X"38",X"03",X"BB",X"38",X"03",
		X"93",X"67",X"B7",X"10",X"F3",X"7D",X"17",X"2F",X"C9",X"13",X"A1",X"07",X"D9",X"08",X"95",X"0C",
		X"EB",X"0F",X"A7",X"10",X"F2",X"10",X"10",X"12",X"2C",X"13",X"A1",X"13",X"25",X"14",X"39",X"15",
		X"C1",X"15",X"DB",X"15",X"1F",X"16",X"AE",X"16",X"29",X"17",X"D2",X"17",X"36",X"18",X"A3",X"18",
		X"FF",X"A5",X"07",X"CA",X"08",X"04",X"AE",X"07",X"BB",X"07",X"C8",X"07",X"D5",X"07",X"80",X"10",
		X"00",X"00",X"00",X"01",X"00",X"E2",X"07",X"07",X"20",X"00",X"00",X"80",X"11",X"00",X"00",X"00",
		X"01",X"00",X"F7",X"07",X"07",X"20",X"00",X"00",X"80",X"12",X"00",X"00",X"00",X"01",X"00",X"21",
		X"08",X"07",X"20",X"00",X"00",X"80",X"22",X"00",X"00",X"00",X"01",X"00",X"0C",X"08",X"EF",X"20",
		X"00",X"00",X"82",X"0D",X"81",X"14",X"86",X"01",X"88",X"36",X"08",X"88",X"45",X"08",X"88",X"52",
		X"08",X"88",X"5D",X"08",X"8A",X"E2",X"07",X"82",X"0E",X"81",X"14",X"86",X"02",X"88",X"62",X"08",
		X"88",X"6A",X"08",X"88",X"72",X"08",X"88",X"7A",X"08",X"8A",X"F7",X"07",X"82",X"0D",X"81",X"14",
		X"86",X"01",X"88",X"82",X"08",X"88",X"8C",X"08",X"88",X"82",X"08",X"88",X"96",X"08",X"8A",X"0C",
		X"08",X"82",X"0D",X"81",X"14",X"86",X"01",X"88",X"A0",X"08",X"88",X"AE",X"08",X"88",X"A0",X"08",
		X"88",X"BC",X"08",X"8A",X"21",X"08",X"19",X"02",X"1D",X"02",X"20",X"02",X"19",X"02",X"1D",X"02",
		X"20",X"02",X"25",X"04",X"89",X"22",X"04",X"1E",X"04",X"22",X"02",X"1E",X"02",X"22",X"02",X"25",
		X"02",X"89",X"25",X"02",X"25",X"02",X"29",X"04",X"2C",X"02",X"29",X"06",X"89",X"27",X"06",X"20",
		X"0A",X"89",X"2C",X"01",X"8C",X"00",X"10",X"62",X"08",X"89",X"2A",X"01",X"8C",X"00",X"10",X"6A",
		X"08",X"89",X"29",X"01",X"8C",X"00",X"10",X"72",X"08",X"89",X"27",X"01",X"8C",X"00",X"10",X"7A",
		X"08",X"89",X"20",X"02",X"1D",X"02",X"8C",X"01",X"04",X"82",X"08",X"89",X"22",X"02",X"1E",X"02",
		X"8C",X"01",X"04",X"8C",X"08",X"89",X"24",X"02",X"20",X"02",X"8C",X"01",X"04",X"96",X"08",X"89",
		X"1D",X"02",X"19",X"02",X"20",X"02",X"19",X"02",X"8C",X"02",X"02",X"A0",X"08",X"89",X"1E",X"02",
		X"19",X"02",X"22",X"02",X"19",X"02",X"8C",X"02",X"02",X"AE",X"08",X"89",X"20",X"02",X"1B",X"02",
		X"20",X"02",X"18",X"02",X"8C",X"02",X"02",X"A0",X"08",X"89",X"CE",X"08",X"D4",X"08",X"CE",X"FE",
		X"DC",X"BA",X"A9",X"01",X"EF",X"EC",X"BA",X"01",X"FF",X"DD",X"08",X"0C",X"0C",X"03",X"E4",X"08",
		X"F1",X"08",X"FE",X"08",X"80",X"10",X"00",X"00",X"00",X"01",X"00",X"33",X"09",X"0C",X"20",X"00",
		X"00",X"80",X"11",X"00",X"00",X"00",X"01",X"00",X"0E",X"09",X"0C",X"20",X"00",X"00",X"80",X"12",
		X"00",X"00",X"00",X"01",X"00",X"52",X"09",X"18",X"20",X"00",X"00",X"81",X"1A",X"89",X"88",X"0B",
		X"09",X"82",X"0E",X"88",X"6D",X"09",X"82",X"0D",X"88",X"F2",X"09",X"88",X"17",X"0A",X"88",X"3C",
		X"0A",X"88",X"61",X"0A",X"88",X"86",X"0A",X"88",X"AB",X"0A",X"88",X"CA",X"0A",X"88",X"E5",X"0A",
		X"8A",X"16",X"09",X"88",X"0B",X"09",X"82",X"0E",X"88",X"9E",X"09",X"82",X"0C",X"88",X"0E",X"0B",
		X"88",X"1F",X"0B",X"88",X"2C",X"0B",X"88",X"45",X"0B",X"88",X"5A",X"0B",X"88",X"75",X"0B",X"8A",
		X"3B",X"09",X"88",X"0B",X"09",X"82",X"0E",X"88",X"CF",X"09",X"82",X"0D",X"86",X"0C",X"88",X"84",
		X"0B",X"88",X"A5",X"0B",X"88",X"C6",X"0B",X"88",X"E7",X"0B",X"8A",X"5A",X"09",X"86",X"01",X"2C",
		X"01",X"2E",X"01",X"2C",X"01",X"2B",X"01",X"86",X"02",X"2C",X"02",X"20",X"02",X"86",X"07",X"2C",
		X"02",X"2A",X"02",X"29",X"02",X"27",X"02",X"86",X"03",X"25",X"03",X"86",X"02",X"27",X"01",X"86",
		X"0B",X"29",X"02",X"2A",X"02",X"2C",X"02",X"00",X"02",X"20",X"02",X"00",X"02",X"89",X"86",X"01",
		X"29",X"01",X"2A",X"01",X"29",X"01",X"28",X"01",X"86",X"02",X"29",X"02",X"00",X"02",X"86",X"07",
		X"29",X"02",X"27",X"02",X"25",X"02",X"24",X"02",X"86",X"03",X"20",X"03",X"86",X"02",X"1E",X"01",
		X"86",X"0B",X"1D",X"02",X"1B",X"02",X"1D",X"02",X"00",X"02",X"1D",X"02",X"00",X"02",X"89",X"86",
		X"0C",X"01",X"06",X"86",X"0B",X"01",X"02",X"86",X"07",X"01",X"02",X"08",X"02",X"0D",X"02",X"08",
		X"02",X"86",X"0C",X"01",X"04",X"05",X"04",X"86",X"0B",X"01",X"02",X"00",X"02",X"01",X"02",X"00",
		X"02",X"89",X"86",X"01",X"29",X"01",X"2A",X"01",X"29",X"01",X"2A",X"01",X"2C",X"01",X"2A",X"01",
		X"2C",X"01",X"2A",X"01",X"29",X"01",X"2A",X"01",X"29",X"01",X"2A",X"01",X"2C",X"01",X"2A",X"01",
		X"2C",X"01",X"86",X"02",X"2A",X"01",X"89",X"86",X"01",X"29",X"01",X"2A",X"01",X"2C",X"01",X"2E",
		X"01",X"30",X"01",X"31",X"01",X"30",X"01",X"29",X"01",X"2A",X"01",X"2C",X"01",X"2A",X"01",X"86",
		X"02",X"29",X"01",X"86",X"03",X"2A",X"02",X"86",X"04",X"27",X"02",X"89",X"86",X"01",X"27",X"01",
		X"29",X"01",X"27",X"01",X"29",X"01",X"2A",X"01",X"29",X"01",X"2A",X"01",X"29",X"01",X"27",X"01",
		X"29",X"01",X"27",X"01",X"29",X"01",X"2A",X"01",X"29",X"01",X"2A",X"01",X"86",X"02",X"29",X"01",
		X"89",X"86",X"01",X"27",X"01",X"29",X"01",X"2A",X"01",X"2C",X"01",X"2E",X"01",X"30",X"01",X"2E",
		X"01",X"2C",X"01",X"2A",X"01",X"2E",X"01",X"2C",X"01",X"86",X"02",X"2B",X"01",X"86",X"03",X"2C",
		X"02",X"86",X"04",X"29",X"02",X"89",X"86",X"01",X"29",X"01",X"2A",X"01",X"29",X"01",X"2A",X"01",
		X"2C",X"01",X"2B",X"01",X"2C",X"01",X"2A",X"01",X"29",X"01",X"2A",X"01",X"29",X"01",X"2A",X"01",
		X"2C",X"01",X"2B",X"01",X"2C",X"01",X"86",X"02",X"2A",X"01",X"89",X"86",X"01",X"29",X"01",X"2A",
		X"01",X"2C",X"01",X"2E",X"01",X"30",X"01",X"31",X"01",X"30",X"01",X"2E",X"01",X"2C",X"01",X"30",
		X"01",X"2E",X"01",X"2D",X"01",X"86",X"05",X"2E",X"04",X"89",X"86",X"06",X"31",X"01",X"30",X"01",
		X"31",X"02",X"25",X"01",X"24",X"01",X"25",X"02",X"2E",X"01",X"2D",X"01",X"2E",X"02",X"22",X"01",
		X"21",X"01",X"22",X"02",X"89",X"86",X"01",X"2C",X"01",X"2E",X"01",X"2C",X"01",X"86",X"02",X"20",
		X"01",X"86",X"01",X"2A",X"01",X"2C",X"01",X"2A",X"01",X"86",X"02",X"20",X"01",X"86",X"01",X"27",
		X"01",X"26",X"01",X"27",X"01",X"86",X"02",X"20",X"01",X"2C",X"02",X"20",X"02",X"89",X"86",X"08",
		X"20",X"0A",X"86",X"09",X"1D",X"02",X"1E",X"02",X"1F",X"02",X"86",X"08",X"20",X"0A",X"89",X"86",
		X"09",X"25",X"02",X"24",X"02",X"22",X"02",X"86",X"08",X"20",X"0A",X"89",X"86",X"09",X"1E",X"02",
		X"1D",X"02",X"1B",X"02",X"86",X"08",X"1E",X"0A",X"86",X"09",X"1D",X"02",X"1B",X"02",X"19",X"02",
		X"86",X"08",X"20",X"0A",X"89",X"86",X"09",X"1D",X"02",X"1E",X"02",X"1F",X"02",X"86",X"08",X"20",
		X"0A",X"86",X"09",X"1E",X"02",X"1D",X"02",X"1E",X"02",X"89",X"86",X"06",X"29",X"01",X"28",X"01",
		X"29",X"02",X"1D",X"01",X"1C",X"01",X"1D",X"02",X"2A",X"01",X"29",X"01",X"2A",X"02",X"1E",X"01",
		X"1D",X"01",X"1E",X"02",X"89",X"86",X"08",X"1B",X"09",X"00",X"01",X"86",X"09",X"1B",X"02",X"1D",
		X"02",X"1E",X"02",X"89",X"01",X"02",X"0D",X"02",X"08",X"02",X"0D",X"02",X"01",X"02",X"0D",X"02",
		X"08",X"02",X"0D",X"02",X"01",X"02",X"0D",X"02",X"08",X"02",X"0D",X"02",X"0A",X"02",X"08",X"02",
		X"06",X"02",X"05",X"02",X"89",X"03",X"02",X"0C",X"02",X"0F",X"02",X"0C",X"02",X"08",X"02",X"0C",
		X"02",X"08",X"02",X"0C",X"02",X"08",X"02",X"0C",X"02",X"0F",X"02",X"0C",X"02",X"0D",X"02",X"08",
		X"02",X"05",X"02",X"01",X"02",X"89",X"01",X"02",X"0D",X"02",X"08",X"02",X"0D",X"02",X"01",X"02",
		X"0D",X"02",X"08",X"02",X"0D",X"02",X"01",X"02",X"0D",X"02",X"08",X"02",X"0D",X"02",X"0A",X"02",
		X"06",X"02",X"0D",X"02",X"06",X"02",X"89",X"86",X"0C",X"01",X"04",X"86",X"0B",X"08",X"02",X"0D",
		X"02",X"86",X"0C",X"01",X"04",X"86",X"0B",X"06",X"02",X"0D",X"02",X"86",X"0C",X"0C",X"04",X"08",
		X"04",X"86",X"0B",X"08",X"02",X"06",X"02",X"05",X"02",X"03",X"02",X"89",X"24",X"0C",X"2C",X"0C",
		X"24",X"0C",X"2C",X"0C",X"33",X"0C",X"43",X"0C",X"4F",X"0C",X"5C",X"0C",X"5C",X"0C",X"65",X"0C",
		X"7D",X"0C",X"86",X"0C",X"DE",X"FF",X"FF",X"EE",X"DC",X"BA",X"99",X"01",X"DE",X"FF",X"ED",X"B9",
		X"75",X"32",X"01",X"CD",X"EF",X"FF",X"FE",X"ED",X"DC",X"CB",X"BB",X"AA",X"AA",X"99",X"99",X"98",
		X"88",X"77",X"01",X"CD",X"ED",X"FF",X"FE",X"EE",X"DD",X"DC",X"CB",X"97",X"53",X"21",X"01",X"DE",
		X"FF",X"FE",X"ED",X"DC",X"CC",X"BB",X"AA",X"99",X"88",X"76",X"65",X"01",X"DD",X"DD",X"EE",X"EE",
		X"FF",X"FF",X"EE",X"EE",X"00",X"AB",X"CD",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",
		X"EE",X"ED",X"DD",X"DD",X"CC",X"CC",X"CB",X"BB",X"BB",X"AA",X"AA",X"A9",X"01",X"DE",X"FF",X"FF",
		X"FF",X"ED",X"DA",X"87",X"43",X"01",X"EF",X"FF",X"FE",X"EE",X"EE",X"DD",X"DD",X"DC",X"CC",X"BB",
		X"BA",X"A9",X"98",X"01",X"FF",X"99",X"0C",X"BE",X"0F",X"05",X"A4",X"0C",X"B2",X"0C",X"C0",X"0C",
		X"CE",X"0C",X"DC",X"0C",X"80",X"20",X"00",X"00",X"00",X"01",X"00",X"EA",X"0C",X"0C",X"20",X"00",
		X"00",X"0F",X"80",X"21",X"00",X"00",X"00",X"01",X"00",X"17",X"0D",X"0C",X"20",X"00",X"00",X"0E",
		X"80",X"10",X"00",X"00",X"00",X"01",X"00",X"40",X"0D",X"00",X"20",X"00",X"00",X"0F",X"80",X"11",
		X"00",X"00",X"00",X"05",X"00",X"EA",X"0C",X"0C",X"20",X"00",X"00",X"0E",X"80",X"12",X"00",X"00",
		X"00",X"01",X"00",X"70",X"0D",X"00",X"20",X"00",X"00",X"0E",X"81",X"18",X"86",X"01",X"20",X"02",
		X"88",X"9D",X"0D",X"88",X"A8",X"0D",X"88",X"B7",X"0D",X"88",X"C2",X"0D",X"88",X"9D",X"0D",X"88",
		X"A8",X"0D",X"88",X"B7",X"0D",X"88",X"CD",X"0D",X"88",X"DA",X"0D",X"88",X"EB",X"0D",X"88",X"FC",
		X"0D",X"88",X"0D",X"0E",X"8A",X"F0",X"0C",X"81",X"18",X"86",X"03",X"1D",X"02",X"88",X"18",X"0E",
		X"88",X"2D",X"0E",X"88",X"42",X"0E",X"88",X"57",X"0E",X"8C",X"00",X"02",X"1D",X"0D",X"88",X"57",
		X"0E",X"88",X"57",X"0E",X"88",X"6E",X"0E",X"88",X"8F",X"0E",X"88",X"8F",X"0E",X"8A",X"1D",X"0D",
		X"81",X"18",X"86",X"04",X"0D",X"02",X"88",X"A4",X"0E",X"88",X"B9",X"0E",X"88",X"CE",X"0E",X"88",
		X"E3",X"0E",X"88",X"A4",X"0E",X"88",X"B9",X"0E",X"88",X"CE",X"0E",X"88",X"F8",X"0E",X"88",X"0D",
		X"0F",X"88",X"0D",X"0F",X"88",X"1E",X"0F",X"88",X"2F",X"0F",X"88",X"3C",X"0F",X"8A",X"46",X"0D",
		X"81",X"18",X"00",X"02",X"86",X"02",X"88",X"51",X"0F",X"88",X"60",X"0F",X"88",X"6D",X"0F",X"88",
		X"7A",X"0F",X"88",X"51",X"0F",X"88",X"60",X"0F",X"88",X"6D",X"0F",X"88",X"85",X"0F",X"88",X"92",
		X"0F",X"88",X"A3",X"0F",X"88",X"B4",X"0F",X"88",X"BB",X"0F",X"8A",X"74",X"0D",X"25",X"04",X"25",
		X"02",X"29",X"02",X"2C",X"06",X"2C",X"02",X"89",X"2E",X"02",X"2C",X"02",X"2A",X"02",X"29",X"02",
		X"2A",X"04",X"27",X"02",X"20",X"02",X"89",X"24",X"04",X"24",X"02",X"25",X"02",X"27",X"06",X"20",
		X"02",X"89",X"2C",X"04",X"2A",X"02",X"27",X"02",X"29",X"06",X"20",X"02",X"89",X"2C",X"02",X"2A",
		X"02",X"29",X"02",X"27",X"02",X"25",X"06",X"20",X"02",X"89",X"27",X"02",X"27",X"02",X"27",X"02",
		X"20",X"02",X"29",X"02",X"29",X"02",X"29",X"02",X"20",X"02",X"89",X"27",X"02",X"27",X"02",X"27",
		X"02",X"20",X"02",X"29",X"02",X"2C",X"02",X"2E",X"02",X"30",X"02",X"89",X"31",X"02",X"2C",X"02",
		X"2C",X"02",X"29",X"02",X"2A",X"02",X"25",X"02",X"25",X"02",X"22",X"02",X"89",X"25",X"0F",X"86",
		X"03",X"25",X"0F",X"86",X"01",X"20",X"02",X"89",X"25",X"02",X"1D",X"01",X"20",X"02",X"25",X"01",
		X"1D",X"02",X"25",X"02",X"1D",X"01",X"20",X"02",X"25",X"01",X"1D",X"02",X"89",X"25",X"02",X"1D",
		X"01",X"20",X"02",X"25",X"01",X"1D",X"02",X"25",X"02",X"1E",X"01",X"20",X"02",X"27",X"01",X"18",
		X"02",X"89",X"20",X"02",X"18",X"01",X"1B",X"02",X"20",X"01",X"18",X"02",X"20",X"02",X"18",X"01",
		X"1B",X"02",X"20",X"01",X"18",X"02",X"89",X"20",X"02",X"18",X"01",X"1B",X"01",X"1E",X"01",X"20",
		X"01",X"18",X"02",X"25",X"02",X"1D",X"01",X"20",X"02",X"25",X"01",X"1D",X"02",X"89",X"25",X"01",
		X"2C",X"01",X"2C",X"01",X"29",X"01",X"2C",X"01",X"29",X"01",X"29",X"01",X"25",X"01",X"2A",X"01",
		X"19",X"01",X"19",X"01",X"16",X"01",X"19",X"01",X"16",X"01",X"16",X"01",X"12",X"01",X"89",X"19",
		X"02",X"1D",X"01",X"20",X"02",X"1D",X"01",X"19",X"02",X"19",X"02",X"1D",X"01",X"20",X"02",X"1D",
		X"01",X"19",X"02",X"89",X"11",X"02",X"0D",X"02",X"14",X"02",X"0D",X"02",X"11",X"01",X"11",X"01",
		X"0D",X"02",X"14",X"01",X"14",X"01",X"0D",X"02",X"89",X"11",X"02",X"0D",X"02",X"14",X"02",X"0D",
		X"02",X"12",X"01",X"12",X"01",X"0D",X"02",X"0F",X"01",X"0F",X"01",X"08",X"02",X"89",X"0C",X"02",
		X"08",X"02",X"0F",X"02",X"08",X"02",X"0C",X"01",X"0C",X"01",X"08",X"02",X"0F",X"01",X"0F",X"01",
		X"08",X"02",X"89",X"0C",X"02",X"08",X"02",X"0F",X"02",X"08",X"02",X"11",X"01",X"11",X"01",X"0D",
		X"02",X"14",X"01",X"14",X"01",X"14",X"02",X"89",X"0C",X"02",X"08",X"02",X"0F",X"02",X"08",X"02",
		X"11",X"01",X"11",X"01",X"0D",X"02",X"0D",X"01",X"0D",X"01",X"0D",X"02",X"89",X"0C",X"02",X"08",
		X"02",X"0F",X"02",X"08",X"02",X"11",X"02",X"0D",X"02",X"14",X"02",X"0D",X"02",X"89",X"0D",X"02",
		X"01",X"02",X"0D",X"02",X"01",X"02",X"12",X"02",X"06",X"02",X"12",X"02",X"06",X"02",X"89",X"0D",
		X"02",X"0D",X"01",X"0D",X"05",X"0D",X"02",X"0D",X"01",X"0D",X"05",X"89",X"0D",X"02",X"11",X"01",
		X"14",X"02",X"11",X"01",X"0D",X"02",X"0D",X"02",X"11",X"01",X"14",X"02",X"11",X"01",X"0D",X"02",
		X"89",X"00",X"02",X"2C",X"02",X"2C",X"02",X"2C",X"02",X"29",X"06",X"25",X"01",X"25",X"01",X"89",
		X"25",X"02",X"24",X"02",X"20",X"02",X"20",X"02",X"1E",X"04",X"1B",X"04",X"89",X"00",X"02",X"27",
		X"02",X"27",X"02",X"27",X"02",X"24",X"06",X"20",X"02",X"89",X"1B",X"02",X"1B",X"02",X"20",X"02",
		X"20",X"02",X"20",X"08",X"89",X"1B",X"02",X"1B",X"02",X"20",X"04",X"20",X"02",X"1D",X"02",X"19",
		X"04",X"89",X"20",X"02",X"20",X"02",X"20",X"02",X"20",X"02",X"20",X"02",X"20",X"02",X"20",X"02",
		X"20",X"02",X"89",X"20",X"02",X"20",X"02",X"20",X"02",X"20",X"02",X"20",X"02",X"20",X"02",X"22",
		X"02",X"24",X"02",X"89",X"86",X"04",X"25",X"08",X"25",X"08",X"89",X"25",X"20",X"89",X"C6",X"0F",
		X"D0",X"0F",X"D9",X"0F",X"DF",X"0F",X"CE",X"FF",X"FE",X"DC",X"BB",X"BB",X"AA",X"AA",X"98",X"01",
		X"BC",X"DE",X"FD",X"CB",X"BB",X"BB",X"BB",X"AA",X"01",X"CD",X"EF",X"FF",X"ED",X"CB",X"01",X"EF",
		X"ED",X"CB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BA",X"98",X"01",X"FF",X"EF",X"0F",X"9B",X"10",X"03",
		X"F6",X"0F",X"03",X"10",X"10",X"10",X"80",X"20",X"00",X"00",X"00",X"01",X"00",X"1D",X"10",X"00",
		X"20",X"00",X"00",X"80",X"21",X"00",X"00",X"00",X"01",X"00",X"47",X"10",X"00",X"20",X"00",X"00",
		X"80",X"22",X"00",X"00",X"00",X"01",X"00",X"71",X"10",X"00",X"20",X"00",X"00",X"81",X"01",X"86",
		X"01",X"82",X"0E",X"31",X"02",X"36",X"03",X"3A",X"03",X"82",X"0F",X"8C",X"00",X"03",X"23",X"10",
		X"3A",X"03",X"3D",X"03",X"42",X"03",X"82",X"0E",X"86",X"02",X"8D",X"31",X"3D",X"0A",X"8E",X"82",
		X"0F",X"8C",X"00",X"03",X"3A",X"10",X"93",X"81",X"01",X"86",X"01",X"82",X"0E",X"3D",X"02",X"3A",
		X"03",X"36",X"03",X"82",X"0F",X"8C",X"01",X"03",X"23",X"10",X"36",X"03",X"3A",X"03",X"3D",X"05",
		X"82",X"0E",X"86",X"02",X"8D",X"38",X"44",X"0A",X"8E",X"82",X"0F",X"8C",X"01",X"03",X"64",X"10",
		X"84",X"81",X"01",X"86",X"01",X"82",X"0E",X"36",X"02",X"31",X"03",X"36",X"03",X"82",X"0F",X"8C",
		X"02",X"03",X"23",X"10",X"31",X"04",X"36",X"03",X"3A",X"03",X"86",X"02",X"82",X"0E",X"8D",X"29",
		X"35",X"0A",X"8E",X"82",X"0F",X"8C",X"02",X"03",X"8E",X"10",X"84",X"9F",X"10",X"A2",X"10",X"FE",
		X"DD",X"01",X"FE",X"DC",X"A9",X"01",X"FF",X"AB",X"10",X"E6",X"10",X"03",X"B2",X"10",X"BF",X"10",
		X"CC",X"10",X"80",X"20",X"00",X"00",X"00",X"01",X"00",X"D9",X"10",X"02",X"20",X"00",X"00",X"80",
		X"21",X"00",X"00",X"00",X"01",X"00",X"D9",X"10",X"0A",X"20",X"00",X"00",X"80",X"22",X"00",X"00",
		X"00",X"01",X"00",X"D9",X"10",X"0E",X"20",X"00",X"00",X"82",X"0F",X"81",X"01",X"86",X"01",X"28",
		X"01",X"29",X"1E",X"00",X"32",X"94",X"E8",X"10",X"EF",X"FE",X"DD",X"CC",X"BA",X"99",X"88",X"77",
		X"01",X"FF",X"F6",X"10",X"A0",X"11",X"05",X"01",X"11",X"0E",X"11",X"1B",X"11",X"28",X"11",X"35",
		X"11",X"80",X"20",X"00",X"00",X"00",X"01",X"00",X"42",X"11",X"11",X"20",X"00",X"00",X"80",X"21",
		X"00",X"00",X"00",X"01",X"00",X"42",X"11",X"05",X"20",X"00",X"00",X"80",X"22",X"00",X"00",X"00",
		X"01",X"00",X"62",X"11",X"05",X"20",X"00",X"00",X"80",X"10",X"00",X"00",X"00",X"01",X"00",X"62",
		X"11",X"05",X"20",X"00",X"00",X"80",X"11",X"00",X"00",X"00",X"01",X"00",X"86",X"11",X"05",X"20",
		X"00",X"00",X"81",X"14",X"82",X"0F",X"86",X"01",X"25",X"01",X"26",X"01",X"25",X"01",X"26",X"01",
		X"86",X"02",X"25",X"02",X"1D",X"02",X"86",X"03",X"20",X"04",X"8D",X"86",X"04",X"25",X"19",X"08",
		X"8E",X"84",X"81",X"14",X"82",X"0F",X"86",X"05",X"00",X"04",X"29",X"02",X"25",X"02",X"86",X"01",
		X"25",X"01",X"26",X"01",X"25",X"01",X"26",X"01",X"86",X"02",X"25",X"02",X"1D",X"02",X"8D",X"86",
		X"04",X"20",X"19",X"04",X"8E",X"84",X"81",X"14",X"82",X"0F",X"86",X"05",X"31",X"02",X"2C",X"02",
		X"25",X"02",X"20",X"02",X"19",X"02",X"14",X"02",X"8D",X"86",X"04",X"0D",X"19",X"08",X"8E",X"84",
		X"AA",X"11",X"B0",X"11",X"BB",X"11",X"D0",X"11",X"FA",X"11",X"BC",X"EF",X"FF",X"FE",X"DC",X"01",
		X"DF",X"FE",X"DC",X"CC",X"CC",X"CC",X"CC",X"CB",X"A9",X"75",X"01",X"67",X"89",X"AB",X"CD",X"ED",
		X"DF",X"DF",X"DF",X"CF",X"CF",X"CF",X"CF",X"BF",X"BF",X"BF",X"AF",X"AF",X"AE",X"DC",X"85",X"01",
		X"EF",X"EF",X"EF",X"EF",X"EF",X"DE",X"DE",X"DE",X"DE",X"DE",X"CD",X"CD",X"CD",X"CD",X"CD",X"BC",
		X"BC",X"BC",X"BC",X"BC",X"AB",X"AB",X"AB",X"AB",X"AB",X"9A",X"9A",X"9A",X"9A",X"9A",X"89",X"89",
		X"89",X"78",X"78",X"67",X"67",X"67",X"56",X"56",X"42",X"01",X"EF",X"FF",X"FE",X"DC",X"BA",X"99",
		X"88",X"77",X"66",X"55",X"44",X"77",X"66",X"55",X"44",X"33",X"55",X"44",X"33",X"22",X"01",X"FF",
		X"14",X"12",X"FD",X"12",X"06",X"21",X"12",X"2E",X"12",X"3B",X"12",X"48",X"12",X"55",X"12",X"62",
		X"12",X"80",X"20",X"00",X"00",X"00",X"01",X"00",X"6F",X"12",X"00",X"20",X"00",X"00",X"80",X"21",
		X"00",X"00",X"00",X"01",X"00",X"6F",X"12",X"F4",X"20",X"00",X"00",X"80",X"22",X"00",X"00",X"00",
		X"01",X"00",X"99",X"12",X"00",X"20",X"00",X"00",X"80",X"10",X"00",X"00",X"00",X"01",X"00",X"99",
		X"12",X"00",X"20",X"00",X"00",X"80",X"11",X"00",X"00",X"00",X"01",X"00",X"D0",X"12",X"0C",X"20",
		X"00",X"00",X"80",X"12",X"00",X"00",X"00",X"01",X"00",X"D0",X"12",X"00",X"20",X"00",X"00",X"82",
		X"0F",X"81",X"14",X"86",X"01",X"3D",X"01",X"38",X"01",X"35",X"01",X"31",X"01",X"2C",X"01",X"29",
		X"01",X"25",X"01",X"20",X"01",X"86",X"04",X"1D",X"01",X"19",X"01",X"14",X"01",X"11",X"01",X"8C",
		X"00",X"02",X"6F",X"12",X"86",X"02",X"3D",X"04",X"84",X"82",X"0F",X"81",X"14",X"86",X"02",X"00",
		X"04",X"3D",X"01",X"38",X"01",X"35",X"01",X"31",X"01",X"86",X"04",X"2C",X"01",X"29",X"01",X"25",
		X"01",X"20",X"01",X"1D",X"01",X"19",X"01",X"14",X"01",X"11",X"01",X"0D",X"01",X"11",X"01",X"14",
		X"01",X"19",X"01",X"1D",X"01",X"20",X"01",X"25",X"01",X"29",X"01",X"86",X"02",X"25",X"04",X"84",
		X"82",X"0F",X"81",X"14",X"86",X"03",X"00",X"08",X"01",X"01",X"05",X"01",X"08",X"01",X"0D",X"01",
		X"11",X"01",X"14",X"01",X"19",X"01",X"1D",X"01",X"20",X"01",X"25",X"01",X"29",X"01",X"2C",X"01",
		X"25",X"01",X"20",X"01",X"1D",X"01",X"19",X"01",X"86",X"02",X"01",X"04",X"84",X"05",X"13",X"11",
		X"13",X"26",X"13",X"0B",X"13",X"FE",X"DD",X"DC",X"BB",X"BA",X"01",X"DE",X"FF",X"FE",X"DC",X"BA",
		X"01",X"CD",X"FF",X"FE",X"EE",X"DD",X"CC",X"CC",X"CC",X"CC",X"CC",X"BB",X"BA",X"AA",X"A9",X"99",
		X"99",X"99",X"88",X"88",X"87",X"01",X"DE",X"FF",X"DC",X"BB",X"01",X"FF",X"30",X"13",X"8C",X"13",
		X"03",X"37",X"13",X"44",X"13",X"51",X"13",X"80",X"20",X"00",X"00",X"00",X"01",X"00",X"5E",X"13",
		X"0B",X"20",X"00",X"00",X"80",X"21",X"00",X"00",X"00",X"01",X"00",X"75",X"13",X"F7",X"20",X"00",
		X"00",X"80",X"22",X"00",X"00",X"00",X"01",X"00",X"75",X"13",X"FD",X"20",X"00",X"00",X"82",X"0F",
		X"81",X"01",X"86",X"01",X"2B",X"01",X"2C",X"09",X"86",X"00",X"2F",X"01",X"30",X"09",X"86",X"02",
		X"30",X"01",X"31",X"10",X"95",X"82",X"0F",X"81",X"01",X"86",X"02",X"2B",X"01",X"2C",X"09",X"86",
		X"01",X"2F",X"01",X"30",X"09",X"86",X"03",X"30",X"01",X"31",X"10",X"84",X"92",X"13",X"96",X"13",
		X"9B",X"13",X"DF",X"ED",X"CC",X"01",X"DF",X"EE",X"DC",X"B7",X"01",X"EF",X"FF",X"EC",X"A8",X"01",
		X"FF",X"A5",X"13",X"1C",X"14",X"01",X"A8",X"13",X"80",X"10",X"00",X"00",X"00",X"01",X"00",X"B5",
		X"13",X"FF",X"20",X"00",X"00",X"81",X"01",X"82",X"0F",X"86",X"01",X"1B",X"02",X"1D",X"0D",X"1D",
		X"02",X"1E",X"0D",X"1D",X"02",X"1F",X"0D",X"22",X"02",X"24",X"0D",X"18",X"02",X"19",X"0D",X"1B",
		X"02",X"1D",X"0D",X"1D",X"02",X"1F",X"0D",X"24",X"02",X"25",X"0D",X"22",X"02",X"24",X"0D",X"24",
		X"02",X"25",X"0D",X"1B",X"02",X"1D",X"0D",X"29",X"02",X"2A",X"0D",X"29",X"02",X"2A",X"0D",X"1E",
		X"02",X"20",X"0D",X"16",X"02",X"18",X"0D",X"24",X"02",X"25",X"0D",X"25",X"02",X"27",X"0D",X"2A",
		X"02",X"2C",X"0D",X"25",X"02",X"28",X"0D",X"22",X"02",X"24",X"0D",X"24",X"02",X"25",X"0D",X"25",
		X"02",X"27",X"0D",X"2A",X"02",X"2D",X"0D",X"22",X"02",X"30",X"0D",X"96",X"1E",X"14",X"FF",X"FF",
		X"EC",X"A8",X"77",X"01",X"FF",X"27",X"14",X"03",X"2E",X"14",X"3B",X"14",X"48",X"14",X"80",X"20",
		X"00",X"00",X"00",X"01",X"00",X"55",X"14",X"00",X"20",X"00",X"00",X"80",X"21",X"00",X"00",X"00",
		X"09",X"00",X"C5",X"14",X"F4",X"20",X"00",X"00",X"80",X"22",X"00",X"00",X"00",X"0C",X"00",X"C5",
		X"14",X"F4",X"20",X"00",X"00",X"81",X"01",X"8F",X"82",X"0F",X"00",X"14",X"01",X"00",X"17",X"01",
		X"00",X"1C",X"01",X"00",X"1E",X"01",X"00",X"20",X"01",X"00",X"24",X"01",X"00",X"28",X"01",X"00",
		X"2C",X"01",X"00",X"30",X"01",X"00",X"37",X"01",X"00",X"41",X"01",X"00",X"4B",X"01",X"00",X"55",
		X"01",X"00",X"64",X"01",X"00",X"78",X"01",X"00",X"82",X"01",X"00",X"8C",X"01",X"00",X"96",X"01",
		X"00",X"A0",X"01",X"82",X"0E",X"00",X"AA",X"01",X"00",X"B4",X"01",X"00",X"BE",X"01",X"00",X"C8",
		X"01",X"00",X"DC",X"01",X"00",X"F0",X"01",X"01",X"05",X"01",X"01",X"19",X"01",X"01",X"2D",X"01",
		X"01",X"41",X"01",X"82",X"0D",X"01",X"55",X"01",X"01",X"69",X"01",X"01",X"7D",X"01",X"01",X"91",
		X"01",X"01",X"A5",X"01",X"93",X"81",X"01",X"8F",X"82",X"0F",X"00",X"23",X"01",X"00",X"28",X"01",
		X"00",X"2D",X"01",X"00",X"32",X"01",X"00",X"37",X"01",X"00",X"3C",X"01",X"00",X"41",X"01",X"00",
		X"46",X"01",X"00",X"4B",X"01",X"00",X"50",X"01",X"00",X"55",X"01",X"00",X"5A",X"01",X"00",X"64",
		X"01",X"00",X"6E",X"01",X"00",X"78",X"01",X"00",X"82",X"01",X"00",X"8C",X"01",X"00",X"96",X"01",
		X"00",X"A0",X"01",X"00",X"AA",X"01",X"82",X"0E",X"00",X"B4",X"01",X"00",X"BE",X"01",X"00",X"C8",
		X"01",X"00",X"D2",X"01",X"00",X"DC",X"01",X"00",X"E6",X"01",X"00",X"F0",X"01",X"00",X"FA",X"01",
		X"01",X"05",X"01",X"01",X"0F",X"01",X"82",X"0D",X"01",X"19",X"01",X"01",X"23",X"01",X"01",X"2D",
		X"01",X"01",X"41",X"01",X"01",X"55",X"01",X"84",X"FF",X"3D",X"15",X"B6",X"15",X"03",X"44",X"15",
		X"51",X"15",X"5E",X"15",X"80",X"20",X"00",X"00",X"00",X"01",X"00",X"6B",X"15",X"00",X"20",X"00",
		X"00",X"80",X"21",X"00",X"00",X"00",X"02",X"00",X"6B",X"15",X"00",X"20",X"00",X"00",X"80",X"22",
		X"00",X"00",X"00",X"01",X"00",X"6B",X"15",X"00",X"20",X"00",X"00",X"81",X"01",X"86",X"02",X"82",
		X"0C",X"36",X"01",X"82",X"0C",X"3A",X"01",X"82",X"0C",X"3A",X"01",X"82",X"0D",X"3B",X"01",X"82",
		X"0D",X"3B",X"01",X"82",X"0E",X"3C",X"01",X"82",X"0F",X"3C",X"02",X"3D",X"02",X"82",X"0E",X"86",
		X"01",X"3E",X"03",X"86",X"02",X"82",X"0D",X"30",X"02",X"82",X"0D",X"35",X"02",X"82",X"0C",X"33",
		X"01",X"82",X"0E",X"31",X"01",X"82",X"0D",X"2F",X"02",X"82",X"0D",X"2F",X"02",X"2E",X"02",X"82",
		X"0C",X"86",X"01",X"2D",X"09",X"97",X"BA",X"15",X"BE",X"15",X"FC",X"A7",X"51",X"01",X"FE",X"01",
		X"FF",X"C3",X"15",X"01",X"C6",X"15",X"80",X"21",X"00",X"00",X"00",X"01",X"00",X"D3",X"15",X"00",
		X"20",X"00",X"00",X"81",X"32",X"82",X"0F",X"00",X"0A",X"96",X"FF",X"DF",X"15",X"15",X"16",X"02",
		X"E4",X"15",X"F1",X"15",X"80",X"23",X"00",X"00",X"00",X"01",X"00",X"FE",X"15",X"00",X"20",X"00",
		X"00",X"80",X"13",X"00",X"00",X"00",X"01",X"00",X"06",X"16",X"00",X"20",X"00",X"00",X"88",X"0E",
		X"16",X"85",X"04",X"0D",X"04",X"84",X"88",X"0E",X"16",X"85",X"00",X"3D",X"04",X"84",X"81",X"16",
		X"82",X"0F",X"86",X"01",X"89",X"17",X"16",X"13",X"46",X"79",X"AB",X"AD",X"EF",X"00",X"FF",X"23",
		X"16",X"9E",X"16",X"03",X"2A",X"16",X"37",X"16",X"44",X"16",X"80",X"20",X"00",X"00",X"00",X"01",
		X"00",X"51",X"16",X"07",X"20",X"00",X"00",X"80",X"21",X"00",X"00",X"00",X"08",X"00",X"51",X"16",
		X"FB",X"20",X"00",X"00",X"80",X"22",X"00",X"00",X"00",X"01",X"00",X"7E",X"16",X"FB",X"20",X"00",
		X"00",X"81",X"15",X"82",X"0F",X"86",X"01",X"2E",X"01",X"2C",X"01",X"2A",X"02",X"2A",X"02",X"2A",
		X"02",X"2E",X"01",X"2C",X"01",X"2A",X"02",X"2A",X"02",X"2A",X"02",X"2E",X"01",X"2C",X"01",X"2A",
		X"02",X"35",X"01",X"33",X"01",X"31",X"02",X"38",X"01",X"35",X"01",X"36",X"02",X"84",X"81",X"15",
		X"82",X"0F",X"86",X"02",X"00",X"02",X"22",X"01",X"1E",X"01",X"25",X"01",X"1E",X"01",X"8C",X"01",
		X"05",X"86",X"16",X"19",X"01",X"19",X"01",X"19",X"01",X"19",X"01",X"1E",X"02",X"84",X"A2",X"16",
		X"A8",X"16",X"AC",X"EF",X"FF",X"EC",X"BA",X"01",X"EF",X"FE",X"DC",X"BA",X"01",X"FF",X"B2",X"16",
		X"21",X"17",X"03",X"B9",X"16",X"C6",X"16",X"D3",X"16",X"80",X"20",X"00",X"00",X"00",X"01",X"00",
		X"E0",X"16",X"00",X"20",X"00",X"00",X"80",X"21",X"00",X"00",X"00",X"01",X"00",X"FB",X"16",X"00",
		X"20",X"00",X"00",X"80",X"13",X"00",X"00",X"00",X"01",X"00",X"0A",X"17",X"00",X"20",X"00",X"00",
		X"82",X"0F",X"81",X"01",X"86",X"01",X"2C",X"08",X"25",X"08",X"29",X"08",X"2C",X"07",X"31",X"07",
		X"35",X"07",X"38",X"06",X"3D",X"06",X"41",X"06",X"41",X"03",X"94",X"82",X"0F",X"81",X"01",X"86",
		X"01",X"19",X"10",X"25",X"0F",X"20",X"14",X"01",X"0C",X"84",X"82",X"0F",X"81",X"01",X"86",X"01",
		X"85",X"07",X"8F",X"00",X"03",X"10",X"00",X"05",X"0F",X"00",X"07",X"14",X"00",X"14",X"0C",X"90",
		X"84",X"23",X"17",X"EF",X"EF",X"CB",X"AA",X"01",X"FF",X"2D",X"17",X"C4",X"17",X"06",X"3A",X"17",
		X"47",X"17",X"54",X"17",X"61",X"17",X"6E",X"17",X"7B",X"17",X"80",X"20",X"00",X"00",X"00",X"01",
		X"00",X"88",X"17",X"00",X"20",X"00",X"00",X"80",X"21",X"00",X"00",X"00",X"0A",X"00",X"9B",X"17",
		X"00",X"20",X"00",X"00",X"80",X"22",X"00",X"00",X"00",X"14",X"00",X"AE",X"17",X"00",X"20",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"01",X"00",X"C1",X"17",X"00",X"20",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"01",X"00",X"C1",X"17",X"00",X"20",X"00",X"00",X"00",X"12",X"00",X"00",X"00",
		X"01",X"00",X"C1",X"17",X"00",X"20",X"00",X"00",X"81",X"08",X"82",X"0F",X"86",X"01",X"25",X"02",
		X"31",X"02",X"3D",X"02",X"25",X"02",X"31",X"02",X"3D",X"06",X"94",X"81",X"08",X"82",X"0F",X"86",
		X"01",X"2C",X"02",X"38",X"02",X"44",X"02",X"2C",X"02",X"38",X"02",X"44",X"06",X"94",X"81",X"08",
		X"82",X"0F",X"86",X"01",X"29",X"02",X"35",X"02",X"41",X"02",X"29",X"02",X"35",X"02",X"41",X"05",
		X"94",X"00",X"01",X"84",X"C6",X"17",X"CD",X"EF",X"FF",X"ED",X"DC",X"CB",X"BA",X"A9",X"98",X"87",
		X"01",X"FF",X"D6",X"17",X"31",X"18",X"03",X"DD",X"17",X"EA",X"17",X"F7",X"17",X"80",X"20",X"00",
		X"00",X"00",X"01",X"00",X"04",X"18",X"00",X"20",X"00",X"00",X"80",X"21",X"00",X"00",X"00",X"01",
		X"00",X"04",X"18",X"00",X"20",X"00",X"00",X"80",X"22",X"00",X"00",X"00",X"01",X"00",X"04",X"18",
		X"00",X"20",X"00",X"00",X"81",X"04",X"86",X"01",X"82",X"0B",X"20",X"01",X"82",X"0D",X"2C",X"01",
		X"82",X"0C",X"25",X"01",X"82",X"0E",X"31",X"01",X"82",X"0D",X"29",X"01",X"82",X"0F",X"35",X"01",
		X"82",X"0E",X"2C",X"01",X"82",X"0E",X"38",X"01",X"82",X"0D",X"31",X"01",X"82",X"0C",X"3D",X"01",
		X"98",X"33",X"18",X"EF",X"01",X"FF",X"38",X"18",X"03",X"3F",X"18",X"4C",X"18",X"59",X"18",X"80",
		X"10",X"00",X"00",X"00",X"01",X"00",X"66",X"18",X"00",X"20",X"00",X"00",X"80",X"11",X"00",X"00",
		X"00",X"01",X"00",X"7A",X"18",X"00",X"20",X"00",X"00",X"80",X"12",X"00",X"00",X"00",X"01",X"00",
		X"8E",X"18",X"00",X"20",X"00",X"00",X"81",X"0D",X"82",X"0F",X"0D",X"01",X"01",X"01",X"05",X"01",
		X"08",X"01",X"0D",X"01",X"8C",X"00",X"02",X"66",X"18",X"99",X"81",X"0D",X"82",X"0F",X"01",X"01",
		X"0D",X"01",X"08",X"01",X"05",X"01",X"01",X"01",X"8C",X"00",X"02",X"7A",X"18",X"99",X"81",X"0D",
		X"82",X"0F",X"05",X"01",X"11",X"01",X"01",X"01",X"01",X"01",X"05",X"01",X"8C",X"00",X"02",X"8E",
		X"18",X"99",X"FF",X"A5",X"18",X"01",X"A8",X"18",X"80",X"13",X"00",X"00",X"00",X"01",X"00",X"B5",
		X"18",X"00",X"20",X"00",X"00",X"82",X"0F",X"81",X"05",X"85",X"07",X"8F",X"8D",X"00",X"01",X"00",
		X"05",X"01",X"00",X"05",X"00",X"0A",X"01",X"00",X"0A",X"00",X"0F",X"01",X"00",X"0F",X"00",X"14",
		X"01",X"00",X"14",X"00",X"1E",X"01",X"00",X"1E",X"00",X"28",X"01",X"00",X"28",X"00",X"3C",X"01",
		X"00",X"3C",X"00",X"37",X"01",X"00",X"37",X"00",X"32",X"01",X"8C",X"00",X"0A",X"DB",X"18",X"82",
		X"0E",X"00",X"37",X"00",X"32",X"01",X"82",X"0D",X"00",X"36",X"00",X"31",X"01",X"82",X"0C",X"00",
		X"35",X"00",X"30",X"01",X"82",X"0B",X"00",X"34",X"00",X"2F",X"01",X"82",X"0A",X"00",X"33",X"00",
		X"2E",X"01",X"82",X"09",X"00",X"32",X"00",X"2D",X"01",X"99",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
