library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity kick_sound_cpu is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of kick_sound_cpu is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"F3",X"31",X"FF",X"83",X"ED",X"56",X"18",X"58",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F5",X"3A",X"00",X"E0",X"3A",X"75",X"83",X"3D",
		X"28",X"06",X"32",X"75",X"83",X"F1",X"FB",X"C9",X"3C",X"32",X"74",X"83",X"3E",X"06",X"32",X"75",
		X"83",X"F1",X"FB",X"C9",X"74",X"72",X"6F",X"6E",X"69",X"78",X"20",X"20",X"20",X"20",X"20",X"20",
		X"21",X"00",X"B0",X"36",X"0F",X"21",X"02",X"B0",X"36",X"F0",X"3A",X"00",X"F0",X"CB",X"47",X"20",
		X"4F",X"CB",X"4F",X"20",X"2E",X"AF",X"32",X"77",X"83",X"CD",X"15",X"05",X"CD",X"CD",X"05",X"3A",
		X"77",X"83",X"FE",X"00",X"28",X"1D",X"CB",X"67",X"20",X"05",X"01",X"00",X"10",X"18",X"03",X"01",
		X"00",X"80",X"11",X"01",X"00",X"60",X"69",X"32",X"00",X"D0",X"37",X"3F",X"ED",X"52",X"20",X"FC",
		X"2F",X"18",X"F2",X"3E",X"FF",X"32",X"00",X"D0",X"3A",X"00",X"F0",X"CB",X"57",X"20",X"08",X"CD",
		X"41",X"06",X"18",X"EF",X"3A",X"00",X"F0",X"CB",X"5F",X"20",X"F9",X"CD",X"68",X"06",X"18",X"F4",
		X"06",X"00",X"CD",X"24",X"06",X"06",X"FF",X"CD",X"24",X"06",X"06",X"55",X"CD",X"24",X"06",X"06",
		X"AA",X"CD",X"24",X"06",X"AF",X"32",X"77",X"83",X"CD",X"15",X"05",X"CD",X"CD",X"05",X"3A",X"77",
		X"83",X"32",X"00",X"C0",X"CD",X"E7",X"00",X"31",X"FF",X"83",X"F3",X"ED",X"56",X"CD",X"09",X"01",
		X"CD",X"18",X"39",X"FB",X"AF",X"32",X"74",X"83",X"CD",X"78",X"01",X"CD",X"D4",X"34",X"CD",X"18",
		X"39",X"3A",X"74",X"83",X"B7",X"28",X"FA",X"18",X"EB",X"21",X"B7",X"3C",X"06",X"20",X"11",X"20",
		X"80",X"DD",X"21",X"00",X"80",X"7E",X"DD",X"77",X"00",X"2F",X"12",X"13",X"23",X"DD",X"23",X"10",
		X"F4",X"06",X"06",X"11",X"09",X"00",X"DD",X"21",X"BC",X"82",X"DD",X"36",X"00",X"FF",X"DD",X"36",
		X"01",X"FF",X"DD",X"36",X"02",X"00",X"DD",X"36",X"03",X"00",X"DD",X"36",X"04",X"00",X"DD",X"36",
		X"05",X"00",X"DD",X"36",X"06",X"00",X"DD",X"19",X"10",X"E0",X"06",X"03",X"21",X"6B",X"83",X"36",
		X"00",X"23",X"10",X"FB",X"3E",X"01",X"32",X"0C",X"83",X"32",X"20",X"83",X"3D",X"32",X"1F",X"83",
		X"3A",X"00",X"90",X"E6",X"80",X"32",X"6E",X"83",X"3E",X"55",X"32",X"71",X"83",X"3E",X"06",X"32",
		X"75",X"83",X"3E",X"31",X"32",X"76",X"83",X"C9",X"3A",X"6E",X"83",X"47",X"3A",X"00",X"90",X"A8",
		X"CB",X"7F",X"20",X"31",X"CB",X"40",X"28",X"1E",X"CB",X"80",X"78",X"32",X"6E",X"83",X"CD",X"D6",
		X"01",X"3A",X"70",X"83",X"CB",X"47",X"28",X"0E",X"CD",X"81",X"02",X"CD",X"8F",X"03",X"CD",X"F2",
		X"03",X"CD",X"53",X"39",X"18",X"23",X"CD",X"8F",X"03",X"3A",X"6F",X"83",X"CB",X"47",X"28",X"19",
		X"CD",X"53",X"39",X"18",X"14",X"78",X"2F",X"CB",X"C7",X"32",X"6E",X"83",X"CD",X"8F",X"03",X"3A",
		X"6F",X"83",X"CB",X"47",X"28",X"03",X"CD",X"53",X"39",X"3E",X"01",X"32",X"20",X"83",X"32",X"0C",
		X"83",X"3D",X"32",X"1F",X"83",X"C9",X"3E",X"01",X"32",X"70",X"83",X"DD",X"21",X"00",X"90",X"DD",
		X"46",X"00",X"CB",X"70",X"28",X"23",X"FD",X"21",X"00",X"80",X"FD",X"7E",X"0F",X"E6",X"8F",X"4F",
		X"78",X"17",X"E6",X"70",X"B1",X"FD",X"77",X"0F",X"FD",X"7E",X"1F",X"E6",X"8F",X"4F",X"78",X"17",
		X"17",X"17",X"17",X"E6",X"70",X"B1",X"FD",X"77",X"1F",X"DD",X"7E",X"01",X"4F",X"FE",X"00",X"28",
		X"22",X"CB",X"7F",X"28",X"64",X"DD",X"7E",X"02",X"CB",X"7F",X"20",X"5D",X"79",X"E6",X"7F",X"4F",
		X"06",X"06",X"FD",X"21",X"BC",X"82",X"11",X"09",X"00",X"FD",X"7E",X"06",X"B9",X"28",X"23",X"FD",
		X"19",X"10",X"F6",X"FD",X"21",X"6B",X"83",X"DD",X"46",X"02",X"78",X"E6",X"7F",X"28",X"1B",X"FD",
		X"77",X"01",X"DD",X"7E",X"01",X"CB",X"7F",X"C0",X"DD",X"7E",X"03",X"FE",X"00",X"C8",X"FD",X"77",
		X"02",X"C9",X"DD",X"7E",X"03",X"FD",X"77",X"07",X"18",X"D9",X"DD",X"4E",X"01",X"79",X"FE",X"00",
		X"20",X"09",X"DD",X"7E",X"03",X"FE",X"00",X"20",X"D9",X"18",X"09",X"CB",X"79",X"28",X"D3",X"CB",
		X"78",X"20",X"CF",X"AF",X"32",X"70",X"83",X"18",X"C9",X"79",X"E6",X"7F",X"32",X"6B",X"83",X"18",
		X"B2",X"06",X"03",X"21",X"6B",X"83",X"C5",X"7E",X"4F",X"FE",X"00",X"CA",X"52",X"03",X"3A",X"76",
		X"83",X"91",X"DA",X"52",X"03",X"79",X"FE",X"31",X"20",X"04",X"F3",X"C3",X"00",X"00",X"79",X"FE",
		X"01",X"20",X"0C",X"DD",X"21",X"00",X"80",X"DD",X"7E",X"1F",X"F6",X"80",X"DD",X"77",X"1F",X"79",
		X"FE",X"02",X"20",X"0F",X"DD",X"21",X"00",X"80",X"DD",X"7E",X"1F",X"E6",X"7F",X"DD",X"77",X"1F",
		X"CD",X"59",X"03",X"79",X"FE",X"03",X"20",X"03",X"CD",X"59",X"03",X"79",X"FE",X"0A",X"20",X"07",
		X"3E",X"31",X"32",X"76",X"83",X"18",X"0A",X"79",X"FE",X"0C",X"20",X"05",X"3E",X"1E",X"32",X"76",
		X"83",X"79",X"D9",X"6F",X"26",X"00",X"54",X"5D",X"29",X"29",X"19",X"19",X"19",X"11",X"8F",X"08",
		X"19",X"EB",X"1A",X"FE",X"00",X"20",X"1F",X"01",X"0C",X"83",X"60",X"69",X"3E",X"06",X"08",X"13",
		X"1A",X"FE",X"00",X"28",X"4A",X"7E",X"CD",X"51",X"3B",X"1A",X"77",X"60",X"69",X"34",X"08",X"3D",
		X"FE",X"00",X"20",X"EA",X"18",X"39",X"3E",X"06",X"21",X"20",X"83",X"08",X"13",X"1A",X"FE",X"00",
		X"28",X"2D",X"7E",X"CD",X"51",X"3B",X"1A",X"77",X"26",X"00",X"6F",X"29",X"01",X"E6",X"09",X"09",
		X"01",X"20",X"83",X"0A",X"CB",X"27",X"E5",X"21",X"33",X"83",X"CD",X"51",X"3B",X"EB",X"E3",X"7E",
		X"12",X"23",X"13",X"7E",X"12",X"0A",X"3C",X"02",X"D1",X"60",X"69",X"08",X"3D",X"20",X"CC",X"D9",
		X"AF",X"77",X"23",X"C1",X"05",X"C2",X"86",X"02",X"C9",X"D9",X"DD",X"21",X"BC",X"82",X"01",X"09",
		X"00",X"11",X"0C",X"83",X"3E",X"01",X"12",X"62",X"6B",X"3E",X"06",X"08",X"DD",X"7E",X"03",X"FE",
		X"00",X"28",X"0B",X"1A",X"CD",X"51",X"3B",X"DD",X"7E",X"03",X"77",X"62",X"6B",X"34",X"DD",X"09",
		X"08",X"3D",X"20",X"E7",X"3E",X"00",X"32",X"1F",X"83",X"3C",X"32",X"20",X"83",X"D9",X"C9",X"AF",
		X"32",X"6F",X"83",X"21",X"0C",X"83",X"7E",X"D6",X"01",X"28",X"2A",X"11",X"09",X"00",X"4F",X"DD",
		X"21",X"BC",X"82",X"06",X"06",X"23",X"7E",X"DD",X"BE",X"04",X"20",X"13",X"AF",X"DD",X"77",X"06",
		X"DD",X"77",X"04",X"DD",X"77",X"05",X"3C",X"32",X"6F",X"83",X"0D",X"20",X"E2",X"18",X"06",X"DD",
		X"19",X"10",X"E4",X"18",X"F5",X"21",X"1F",X"83",X"7E",X"4F",X"FE",X"00",X"C8",X"3E",X"01",X"32",
		X"6F",X"83",X"06",X"06",X"21",X"E0",X"3C",X"DD",X"21",X"BC",X"82",X"11",X"09",X"00",X"79",X"A6",
		X"28",X"0A",X"AF",X"DD",X"77",X"06",X"DD",X"77",X"04",X"DD",X"77",X"05",X"DD",X"19",X"23",X"10",
		X"ED",X"C9",X"3A",X"20",X"83",X"D6",X"01",X"C8",X"08",X"CD",X"24",X"04",X"CD",X"40",X"04",X"79",
		X"CB",X"27",X"21",X"33",X"83",X"CD",X"51",X"3B",X"7A",X"FE",X"00",X"20",X"11",X"CB",X"7E",X"20",
		X"0A",X"E5",X"CD",X"81",X"04",X"E1",X"7A",X"FE",X"00",X"20",X"03",X"CD",X"BA",X"04",X"23",X"36",
		X"00",X"08",X"18",X"D1",X"06",X"00",X"0E",X"01",X"16",X"01",X"3A",X"20",X"83",X"5F",X"21",X"33",
		X"83",X"23",X"7A",X"BB",X"C8",X"23",X"23",X"78",X"BE",X"30",X"02",X"46",X"4A",X"14",X"18",X"F2",
		X"79",X"CB",X"27",X"21",X"33",X"83",X"CD",X"51",X"3B",X"C5",X"06",X"06",X"4E",X"11",X"09",X"00",
		X"21",X"E0",X"3C",X"DD",X"21",X"BC",X"82",X"7E",X"A1",X"28",X"1D",X"DD",X"7E",X"04",X"FE",X"00",
		X"20",X"16",X"21",X"20",X"83",X"C1",X"79",X"CD",X"51",X"3B",X"7E",X"DD",X"77",X"04",X"DD",X"70",
		X"05",X"AF",X"DD",X"77",X"03",X"16",X"01",X"C9",X"DD",X"19",X"23",X"10",X"DA",X"16",X"00",X"C1",
		X"C9",X"26",X"06",X"11",X"09",X"00",X"DD",X"21",X"BC",X"82",X"DD",X"7E",X"04",X"FE",X"00",X"20",
		X"15",X"79",X"21",X"20",X"83",X"CD",X"51",X"3B",X"7E",X"DD",X"77",X"04",X"DD",X"70",X"05",X"AF",
		X"DD",X"77",X"03",X"16",X"01",X"C9",X"DD",X"19",X"25",X"20",X"DF",X"16",X"00",X"21",X"33",X"83",
		X"79",X"CB",X"27",X"CD",X"51",X"3B",X"F6",X"3F",X"77",X"C9",X"16",X"FF",X"1E",X"00",X"E5",X"C5",
		X"4E",X"06",X"00",X"DD",X"21",X"BC",X"82",X"21",X"E0",X"3C",X"7E",X"A1",X"28",X"08",X"DD",X"7E",
		X"05",X"BA",X"30",X"02",X"57",X"58",X"D5",X"11",X"09",X"00",X"DD",X"19",X"D1",X"23",X"04",X"78",
		X"FE",X"06",X"20",X"E6",X"C1",X"7A",X"B8",X"30",X"24",X"21",X"20",X"83",X"79",X"CD",X"51",X"3B",
		X"4E",X"6B",X"26",X"00",X"54",X"5D",X"29",X"29",X"29",X"19",X"EB",X"DD",X"21",X"BC",X"82",X"DD",
		X"19",X"DD",X"71",X"04",X"DD",X"70",X"05",X"AF",X"DD",X"77",X"03",X"E1",X"C9",X"E1",X"C0",X"CB",
		X"76",X"C8",X"E5",X"18",X"D4",X"DD",X"21",X"BD",X"05",X"AF",X"F5",X"DD",X"6E",X"00",X"DD",X"66",
		X"01",X"7C",X"B5",X"20",X"0A",X"F1",X"47",X"3A",X"77",X"83",X"B0",X"32",X"77",X"83",X"C9",X"DD",
		X"5E",X"04",X"DD",X"56",X"05",X"DD",X"4E",X"02",X"DD",X"46",X"03",X"ED",X"B0",X"DD",X"6E",X"00",
		X"DD",X"66",X"01",X"DD",X"5E",X"02",X"DD",X"56",X"03",X"7A",X"B3",X"28",X"11",X"06",X"02",X"3E",
		X"00",X"77",X"BE",X"C2",X"B8",X"05",X"F6",X"FF",X"10",X"F7",X"23",X"1B",X"18",X"EB",X"DD",X"66",
		X"01",X"DD",X"6E",X"00",X"DD",X"5E",X"02",X"DD",X"56",X"03",X"7A",X"B3",X"28",X"06",X"36",X"00",
		X"23",X"1B",X"18",X"F6",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"DD",X"5E",X"02",X"DD",X"56",X"03",
		X"7A",X"B3",X"28",X"14",X"7E",X"FE",X"00",X"20",X"2F",X"3E",X"01",X"77",X"BE",X"C2",X"B8",X"05",
		X"CB",X"27",X"30",X"F7",X"23",X"1B",X"18",X"E8",X"AF",X"DD",X"66",X"05",X"DD",X"6E",X"04",X"DD",
		X"56",X"01",X"DD",X"5E",X"00",X"DD",X"4E",X"02",X"DD",X"46",X"03",X"ED",X"B0",X"47",X"F1",X"B0",
		X"11",X"07",X"00",X"DD",X"19",X"C3",X"1A",X"05",X"DD",X"7E",X"06",X"18",X"DC",X"00",X"80",X"00",
		X"02",X"00",X"80",X"10",X"00",X"82",X"00",X"02",X"00",X"80",X"10",X"00",X"00",X"DD",X"21",X"09",
		X"06",X"16",X"00",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"DD",X"4E",X"00",X"DD",X"46",X"01",X"78",
		X"B1",X"28",X"1A",X"AF",X"86",X"23",X"0D",X"20",X"FB",X"05",X"20",X"F8",X"DD",X"BE",X"04",X"28",
		X"05",X"7A",X"DD",X"B6",X"05",X"57",X"01",X"06",X"00",X"DD",X"09",X"18",X"D6",X"7A",X"B7",X"C8",
		X"47",X"3A",X"77",X"83",X"B0",X"32",X"77",X"83",X"C9",X"00",X"10",X"00",X"00",X"86",X"01",X"00",
		X"10",X"00",X"10",X"EC",X"02",X"00",X"10",X"00",X"20",X"41",X"04",X"00",X"10",X"00",X"30",X"F7",
		X"08",X"00",X"00",X"7A",X"3A",X"00",X"90",X"B8",X"20",X"FA",X"3A",X"01",X"90",X"B8",X"20",X"F4",
		X"3A",X"02",X"90",X"B8",X"20",X"EE",X"3A",X"03",X"90",X"B8",X"20",X"E8",X"78",X"32",X"00",X"C0",
		X"C9",X"06",X"00",X"CD",X"A1",X"06",X"0E",X"00",X"3E",X"AD",X"CD",X"E1",X"06",X"0E",X"01",X"3E",
		X"07",X"CD",X"E1",X"06",X"06",X"01",X"CD",X"A1",X"06",X"0E",X"00",X"3E",X"AD",X"CD",X"E1",X"06",
		X"0E",X"01",X"3E",X"77",X"CD",X"E1",X"06",X"C9",X"CD",X"41",X"06",X"16",X"10",X"3E",X"00",X"1E",
		X"FF",X"06",X"00",X"0E",X"00",X"CD",X"E1",X"06",X"2F",X"0E",X"01",X"CD",X"E1",X"06",X"06",X"01",
		X"32",X"78",X"83",X"E6",X"7F",X"CD",X"E1",X"06",X"3A",X"78",X"83",X"2F",X"0E",X"00",X"CD",X"E1",
		X"06",X"3C",X"E6",X"0F",X"47",X"07",X"07",X"07",X"07",X"B0",X"1D",X"20",X"FD",X"15",X"20",X"CF",
		X"C9",X"CD",X"F8",X"06",X"36",X"00",X"DD",X"36",X"00",X"F4",X"36",X"01",X"DD",X"36",X"00",X"01",
		X"36",X"02",X"DD",X"36",X"00",X"FA",X"36",X"03",X"DD",X"36",X"00",X"00",X"36",X"04",X"DD",X"36",
		X"00",X"7D",X"36",X"05",X"DD",X"36",X"00",X"00",X"36",X"08",X"DD",X"36",X"00",X"0B",X"36",X"09",
		X"DD",X"36",X"00",X"0B",X"36",X"0A",X"DD",X"36",X"00",X"0B",X"36",X"07",X"DD",X"36",X"00",X"F8",
		X"C9",X"CD",X"F8",X"06",X"32",X"72",X"83",X"AF",X"A9",X"28",X"09",X"36",X"0F",X"3A",X"72",X"83",
		X"DD",X"77",X"00",X"C9",X"36",X"0E",X"18",X"F5",X"32",X"72",X"83",X"AF",X"A8",X"3A",X"72",X"83",
		X"20",X"08",X"21",X"00",X"A0",X"DD",X"21",X"02",X"A0",X"C9",X"21",X"00",X"B0",X"DD",X"21",X"02",
		X"B0",X"C9",X"11",X"94",X"00",X"CD",X"B9",X"06",X"0E",X"05",X"C5",X"1E",X"4A",X"01",X"50",X"00",
		X"CD",X"DF",X"04",X"0E",X"05",X"C5",X"1E",X"02",X"01",X"F3",X"02",X"CD",X"DF",X"04",X"0E",X"05",
		X"C5",X"1E",X"02",X"01",X"F3",X"02",X"CD",X"DF",X"04",X"21",X"50",X"00",X"36",X"0C",X"21",X"94",
		X"16",X"36",X"04",X"C9",X"21",X"73",X"17",X"73",X"2B",X"70",X"2B",X"71",X"3A",X"73",X"17",X"32",
		X"74",X"17",X"4F",X"3E",X"50",X"B9",X"D2",X"5E",X"07",X"21",X"74",X"17",X"36",X"50",X"01",X"01",
		X"00",X"C5",X"3A",X"74",X"17",X"11",X"71",X"17",X"CD",X"1B",X"13",X"2B",X"EB",X"01",X"5B",X"03",
		X"CD",X"0F",X"13",X"3A",X"C7",X"13",X"1F",X"D2",X"99",X"07",X"3E",X"37",X"21",X"94",X"16",X"BE",
		X"D2",X"86",X"07",X"CD",X"06",X"07",X"0E",X"05",X"C5",X"2A",X"71",X"17",X"44",X"4D",X"2A",X"74",
		X"17",X"EB",X"CD",X"DF",X"04",X"21",X"94",X"16",X"34",X"3A",X"CA",X"13",X"1F",X"D2",X"AF",X"07",
		X"0E",X"01",X"C5",X"2A",X"71",X"17",X"44",X"4D",X"2A",X"74",X"17",X"EB",X"CD",X"DF",X"04",X"C9",
		X"2A",X"25",X"14",X"26",X"00",X"01",X"CB",X"13",X"09",X"7E",X"FE",X"20",X"C2",X"C6",X"07",X"21",
		X"25",X"14",X"35",X"C3",X"B0",X"07",X"21",X"25",X"14",X"34",X"C9",X"01",X"0B",X"00",X"C5",X"2A",
		X"25",X"14",X"26",X"00",X"01",X"CB",X"13",X"09",X"EB",X"01",X"F4",X"02",X"CD",X"0F",X"13",X"01",
		X"08",X"00",X"C5",X"01",X"05",X"00",X"2A",X"68",X"16",X"09",X"E5",X"2A",X"25",X"14",X"26",X"00",
		X"01",X"D6",X"13",X"09",X"EB",X"C1",X"CD",X"0F",X"13",X"3A",X"25",X"14",X"C6",X"12",X"32",X"25",
		X"00",X"8B",X"32",X"93",X"32",X"9B",X"32",X"A6",X"32",X"B1",X"32",X"BC",X"32",X"C7",X"32",X"D2",
		X"32",X"DD",X"32",X"E8",X"32",X"F3",X"32",X"FE",X"32",X"09",X"33",X"14",X"33",X"1F",X"33",X"2A",
		X"33",X"35",X"33",X"3A",X"33",X"3F",X"33",X"44",X"33",X"49",X"33",X"4E",X"33",X"59",X"33",X"64",
		X"33",X"6F",X"33",X"7A",X"33",X"85",X"33",X"90",X"33",X"95",X"33",X"9A",X"33",X"9F",X"33",X"1C",
		X"34",X"32",X"34",X"48",X"34",X"5E",X"34",X"74",X"34",X"7F",X"34",X"A4",X"33",X"95",X"34",X"AB",
		X"34",X"B0",X"34",X"AF",X"33",X"B5",X"34",X"BA",X"34",X"27",X"34",X"3D",X"34",X"53",X"34",X"69",
		X"34",X"B4",X"33",X"A0",X"34",X"BF",X"33",X"CA",X"33",X"D5",X"33",X"E0",X"33",X"EB",X"33",X"F6",
		X"33",X"BF",X"33",X"CA",X"33",X"D5",X"33",X"E0",X"33",X"FB",X"33",X"06",X"34",X"11",X"34",X"14",
		X"33",X"E8",X"32",X"DD",X"32",X"C7",X"32",X"9B",X"32",X"49",X"33",X"44",X"33",X"3A",X"33",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"00",X"00",X"00",
		X"00",X"00",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"01",X"04",X"00",X"00",X"00",X"00",X"00",
		X"01",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"01",X"06",
		X"06",X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1E",X"1E",X"1E",
		X"1E",X"1E",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"10",X"00",X"00",X"00",X"00",
		X"00",X"01",X"11",X"12",X"00",X"00",X"00",X"00",X"01",X"1F",X"20",X"21",X"00",X"00",X"00",X"01",
		X"15",X"16",X"17",X"18",X"19",X"00",X"01",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"1A",X"1B",
		X"1C",X"1D",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"2B",X"00",X"00",X"00",X"00",X"00",X"01",X"1E",X"1E",X"00",X"00",X"00",X"00",
		X"01",X"2C",X"00",X"00",X"00",X"00",X"00",X"01",X"43",X"44",X"45",X"46",X"47",X"48",X"01",X"2D",
		X"00",X"00",X"00",X"00",X"00",X"01",X"2E",X"00",X"00",X"00",X"00",X"00",X"01",X"30",X"00",X"00",
		X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"01",X"31",X"42",X"00",X"00",X"00",
		X"00",X"00",X"31",X"42",X"00",X"00",X"00",X"00",X"01",X"13",X"14",X"13",X"14",X"00",X"00",X"01",
		X"1A",X"1B",X"1C",X"1D",X"00",X"00",X"01",X"23",X"24",X"25",X"26",X"00",X"00",X"01",X"08",X"09",
		X"29",X"2A",X"00",X"00",X"00",X"0A",X"0B",X"0C",X"49",X"00",X"00",X"00",X"23",X"24",X"25",X"26",
		X"00",X"00",X"00",X"08",X"09",X"29",X"2A",X"00",X"00",X"01",X"0A",X"0B",X"0C",X"49",X"00",X"00",
		X"01",X"0D",X"0E",X"0F",X"00",X"00",X"00",X"01",X"32",X"33",X"34",X"35",X"00",X"00",X"00",X"32",
		X"33",X"34",X"35",X"00",X"00",X"01",X"36",X"37",X"38",X"39",X"00",X"00",X"00",X"36",X"37",X"38",
		X"39",X"00",X"00",X"01",X"3A",X"3B",X"3C",X"3D",X"00",X"00",X"00",X"3A",X"3B",X"3C",X"3D",X"00",
		X"00",X"01",X"3E",X"3F",X"40",X"41",X"00",X"00",X"00",X"3E",X"3F",X"40",X"41",X"00",X"00",X"01",
		X"4A",X"4B",X"00",X"00",X"00",X"00",X"00",X"00",X"81",X"0F",X"81",X"05",X"81",X"14",X"81",X"0A",
		X"E0",X"1E",X"1E",X"19",X"BC",X"23",X"86",X"55",X"86",X"55",X"88",X"5A",X"82",X"5A",X"84",X"5A",
		X"9E",X"2D",X"9E",X"2D",X"9E",X"2D",X"9E",X"32",X"9E",X"37",X"9E",X"37",X"9E",X"3C",X"9E",X"3C",
		X"BE",X"41",X"BE",X"41",X"BE",X"41",X"BE",X"41",X"BE",X"41",X"9E",X"46",X"9E",X"46",X"9E",X"46",
		X"9E",X"46",X"A1",X"64",X"E5",X"50",X"E5",X"50",X"E5",X"50",X"C1",X"16",X"86",X"55",X"86",X"55",
		X"98",X"55",X"98",X"55",X"BC",X"3C",X"BC",X"3C",X"98",X"55",X"98",X"55",X"81",X"15",X"C1",X"18",
		X"81",X"18",X"81",X"18",X"81",X"18",X"A0",X"23",X"8A",X"4B",X"82",X"5A",X"88",X"5A",X"84",X"5A",
		X"90",X"5A",X"82",X"5A",X"88",X"5A",X"84",X"5A",X"90",X"5A",X"82",X"5A",X"84",X"5A",X"88",X"5A",
		X"90",X"5A",X"82",X"5A",X"88",X"5A",X"84",X"5A",X"90",X"5A",X"8A",X"4B",X"81",X"43",X"82",X"44",
		X"84",X"45",X"88",X"46",X"90",X"47",X"A0",X"48",X"90",X"4B",X"8A",X"50",X"8A",X"50",X"46",X"0C",
		X"FF",X"FF",X"FF",X"FF",X"50",X"0C",X"69",X"0C",X"5C",X"0C",X"81",X"0C",X"96",X"0C",X"8F",X"0C",
		X"A5",X"0C",X"B8",X"0C",X"B1",X"0C",X"C4",X"0C",X"DF",X"0C",X"D2",X"0C",X"FF",X"0C",X"1A",X"0D",
		X"0D",X"0D",X"3A",X"0D",X"4D",X"0D",X"46",X"0D",X"7A",X"0D",X"FF",X"FF",X"84",X"0D",X"7A",X"0D",
		X"8A",X"0D",X"84",X"0D",X"7A",X"0D",X"9D",X"0D",X"84",X"0D",X"7A",X"0D",X"B6",X"0D",X"84",X"0D",
		X"7A",X"0D",X"D9",X"0D",X"84",X"0D",X"7A",X"0D",X"FC",X"0D",X"84",X"0D",X"7A",X"0D",X"2F",X"0E",
		X"84",X"0D",X"7A",X"0D",X"3C",X"0E",X"84",X"0D",X"7A",X"0D",X"47",X"0E",X"84",X"0D",X"52",X"0E",
		X"73",X"0E",X"60",X"0E",X"7A",X"0D",X"A6",X"0E",X"84",X"0D",X"7A",X"0D",X"B1",X"0E",X"84",X"0D",
		X"7A",X"0D",X"BC",X"0E",X"84",X"0D",X"7A",X"0D",X"CF",X"0E",X"84",X"0D",X"E0",X"0E",X"F5",X"0E",
		X"EA",X"0E",X"E0",X"0E",X"0F",X"0F",X"EA",X"0E",X"E0",X"0E",X"1A",X"0F",X"EA",X"0E",X"E0",X"0E",
		X"25",X"0F",X"EA",X"0E",X"E0",X"0E",X"30",X"0F",X"EA",X"0E",X"7A",X"0D",X"3B",X"0F",X"7A",X"0D",
		X"7A",X"0D",X"62",X"0F",X"84",X"0D",X"7A",X"0D",X"89",X"0F",X"84",X"0D",X"7A",X"0D",X"B0",X"0F",
		X"84",X"0D",X"D8",X"11",X"BB",X"0F",X"E6",X"11",X"CD",X"0F",X"E8",X"0F",X"DB",X"0F",X"03",X"10",
		X"11",X"10",X"DB",X"0F",X"20",X"10",X"2E",X"10",X"DB",X"0F",X"3D",X"10",X"52",X"10",X"4B",X"10",
		X"7A",X"0D",X"59",X"10",X"84",X"0D",X"7A",X"0D",X"99",X"10",X"84",X"0D",X"7A",X"0D",X"CC",X"10",
		X"84",X"0D",X"7A",X"0D",X"33",X"11",X"84",X"0D",X"7A",X"0D",X"FF",X"FF",X"84",X"0D",X"7A",X"0D",
		X"FF",X"FF",X"84",X"0D",X"7A",X"0D",X"82",X"11",X"84",X"0D",X"7A",X"0D",X"B7",X"11",X"84",X"0D",
		X"D8",X"11",X"ED",X"11",X"E6",X"11",X"02",X"12",X"1C",X"12",X"10",X"12",X"7C",X"12",X"97",X"12",
		X"8A",X"12",X"61",X"13",X"6F",X"13",X"10",X"12",X"46",X"0C",X"FF",X"FF",X"FF",X"FF",X"52",X"15",
		X"66",X"15",X"60",X"15",X"B7",X"15",X"D0",X"15",X"C5",X"15",X"7A",X"0D",X"14",X"16",X"84",X"0D",
		X"7A",X"0D",X"5B",X"16",X"84",X"0D",X"7A",X"0D",X"BC",X"16",X"84",X"0D",X"7A",X"0D",X"07",X"17",
		X"84",X"0D",X"7A",X"0D",X"58",X"17",X"84",X"0D",X"7A",X"0D",X"9F",X"17",X"84",X"0D",X"7A",X"0D",
		X"00",X"18",X"84",X"0D",X"7A",X"0D",X"4B",X"18",X"84",X"0D",X"7A",X"0D",X"9C",X"18",X"84",X"0D",
		X"7A",X"0D",X"BF",X"18",X"84",X"0D",X"7A",X"0D",X"E2",X"18",X"84",X"0D",X"7A",X"0D",X"FD",X"18",
		X"84",X"0D",X"7A",X"0D",X"16",X"19",X"84",X"0D",X"7A",X"0D",X"5B",X"19",X"84",X"0D",X"7A",X"0D",
		X"82",X"19",X"84",X"0D",X"7A",X"0D",X"A9",X"19",X"84",X"0D",X"B7",X"15",X"D0",X"19",X"C5",X"15",
		X"14",X"1A",X"29",X"1A",X"22",X"1A",X"3B",X"1A",X"49",X"1A",X"22",X"1A",X"5E",X"1A",X"6C",X"1A",
		X"22",X"1A",X"81",X"1A",X"8F",X"1A",X"22",X"1A",X"A4",X"1A",X"B2",X"1A",X"22",X"1A",X"C7",X"1A",
		X"D5",X"1A",X"22",X"1A",X"7A",X"0D",X"ED",X"1A",X"84",X"0D",X"7A",X"0D",X"16",X"1B",X"84",X"0D",
		X"7A",X"0D",X"23",X"1B",X"84",X"0D",X"CD",X"B6",X"39",X"00",X"00",X"FF",X"0A",X"00",X"FF",X"C9",
		X"CD",X"B6",X"39",X"10",X"01",X"FF",X"0A",X"04",X"04",X"16",X"FF",X"C9",X"CD",X"7A",X"3A",X"00",
		X"0A",X"0A",X"CD",X"7A",X"3A",X"01",X"04",X"04",X"C9",X"CD",X"FC",X"34",X"75",X"0C",X"00",X"01",
		X"00",X"0A",X"01",X"01",X"00",X"CD",X"FC",X"34",X"98",X"10",X"01",X"01",X"00",X"0A",X"01",X"FF",
		X"00",X"CD",X"B6",X"39",X"01",X"01",X"FF",X"0A",X"01",X"00",X"1E",X"02",X"00",X"FF",X"C9",X"CD",
		X"7A",X"3A",X"00",X"0A",X"0A",X"C9",X"CD",X"FC",X"34",X"98",X"10",X"00",X"01",X"00",X"01",X"01",
		X"0B",X"08",X"03",X"FF",X"00",X"CD",X"B6",X"39",X"10",X"00",X"FF",X"0A",X"0F",X"04",X"0B",X"FF",
		X"C9",X"CD",X"7A",X"3A",X"00",X"0A",X"0A",X"C9",X"CD",X"FC",X"34",X"98",X"10",X"00",X"01",X"00",
		X"0F",X"01",X"FF",X"00",X"CD",X"B6",X"39",X"01",X"03",X"FF",X"0A",X"01",X"00",X"FF",X"02",X"00",
		X"FF",X"C9",X"CD",X"7A",X"3A",X"00",X"00",X"00",X"CD",X"7A",X"3A",X"01",X"0A",X"0A",X"C9",X"CD",
		X"FC",X"34",X"F0",X"0C",X"00",X"02",X"10",X"05",X"01",X"0F",X"00",X"07",X"01",X"F3",X"FF",X"00",
		X"CD",X"FC",X"34",X"98",X"10",X"01",X"01",X"00",X"02",X"02",X"07",X"0F",X"07",X"FF",X"00",X"CD",
		X"B6",X"39",X"01",X"04",X"FF",X"0A",X"00",X"00",X"68",X"02",X"00",X"FF",X"C9",X"CD",X"7A",X"3A",
		X"00",X"00",X"00",X"CD",X"7A",X"3A",X"01",X"0A",X"0A",X"C9",X"CD",X"FC",X"34",X"2B",X"0D",X"00",
		X"02",X"00",X"90",X"03",X"02",X"00",X"FF",X"02",X"02",X"00",X"00",X"CD",X"FC",X"34",X"98",X"10",
		X"01",X"01",X"00",X"05",X"01",X"02",X"80",X"FF",X"00",X"00",X"CD",X"B6",X"39",X"10",X"07",X"FF",
		X"0A",X"01",X"04",X"1F",X"FF",X"C9",X"CD",X"7A",X"3A",X"00",X"0A",X"0A",X"C9",X"CD",X"FC",X"34",
		X"98",X"10",X"00",X"01",X"00",X"02",X"01",X"05",X"02",X"01",X"FF",X"01",X"05",X"00",X"02",X"01",
		X"FD",X"02",X"01",X"05",X"02",X"01",X"FF",X"01",X"05",X"00",X"02",X"01",X"FD",X"02",X"01",X"05",
		X"02",X"01",X"FF",X"01",X"05",X"00",X"0D",X"05",X"FF",X"00",X"CD",X"B6",X"39",X"01",X"03",X"FF",
		X"0A",X"00",X"FF",X"C9",X"CD",X"D9",X"3A",X"00",X"C9",X"C9",X"CD",X"E9",X"36",X"89",X"0D",X"00",
		X"18",X"3E",X"25",X"CC",X"23",X"6A",X"24",X"CC",X"23",X"E7",X"24",X"00",X"00",X"CD",X"E9",X"36",
		X"89",X"0D",X"00",X"18",X"4E",X"25",X"EB",X"23",X"5D",X"24",X"86",X"24",X"EB",X"23",X"5D",X"24",
		X"D1",X"24",X"EB",X"23",X"00",X"00",X"CD",X"E9",X"36",X"98",X"10",X"00",X"FF",X"38",X"30",X"3F",
		X"30",X"6D",X"30",X"3F",X"30",X"77",X"30",X"3F",X"30",X"6D",X"30",X"3F",X"30",X"77",X"30",X"3F",
		X"30",X"6D",X"30",X"3F",X"30",X"77",X"30",X"00",X"00",X"CD",X"E9",X"36",X"98",X"10",X"00",X"FF",
		X"EA",X"30",X"EE",X"30",X"04",X"31",X"EE",X"30",X"14",X"31",X"EE",X"30",X"04",X"31",X"EE",X"30",
		X"14",X"31",X"EE",X"30",X"04",X"31",X"EE",X"30",X"14",X"31",X"00",X"00",X"CD",X"E9",X"36",X"98",
		X"10",X"00",X"FF",X"8A",X"31",X"8E",X"31",X"8E",X"31",X"8E",X"31",X"95",X"31",X"8E",X"31",X"A8",
		X"31",X"EA",X"30",X"8E",X"31",X"8E",X"31",X"8E",X"31",X"95",X"31",X"8E",X"31",X"A8",X"31",X"EA",
		X"30",X"8E",X"31",X"8E",X"31",X"8E",X"31",X"95",X"31",X"8E",X"31",X"A8",X"31",X"00",X"00",X"CD",
		X"E9",X"36",X"89",X"0D",X"00",X"00",X"81",X"1B",X"A0",X"1F",X"00",X"00",X"CD",X"E9",X"36",X"89",
		X"0D",X"00",X"00",X"F5",X"1F",X"00",X"00",X"CD",X"E9",X"36",X"89",X"0D",X"00",X"00",X"3E",X"20",
		X"00",X"00",X"CD",X"B6",X"39",X"01",X"05",X"FF",X"0A",X"02",X"00",X"88",X"02",X"00",X"FF",X"C9",
		X"CD",X"7A",X"3A",X"00",X"0A",X"0A",X"CD",X"7A",X"3A",X"01",X"00",X"00",X"CD",X"7A",X"3A",X"02",
		X"00",X"00",X"C9",X"CD",X"FC",X"34",X"85",X"0E",X"00",X"01",X"00",X"04",X"01",X"03",X"01",X"6E",
		X"00",X"0B",X"02",X"FF",X"00",X"CD",X"FC",X"34",X"97",X"0E",X"01",X"01",X"00",X"04",X"01",X"F8",
		X"01",X"6E",X"00",X"0B",X"02",X"04",X"00",X"CD",X"FC",X"34",X"98",X"10",X"02",X"01",X"FF",X"02",
		X"01",X"FA",X"02",X"01",X"06",X"00",X"CD",X"E9",X"36",X"89",X"0D",X"00",X"00",X"91",X"20",X"00",
		X"00",X"CD",X"E9",X"36",X"89",X"0D",X"00",X"00",X"A1",X"20",X"00",X"00",X"CD",X"E9",X"36",X"89",
		X"0D",X"00",X"00",X"30",X"1B",X"88",X"1E",X"A7",X"1E",X"62",X"1B",X"87",X"20",X"00",X"00",X"CD",
		X"E9",X"36",X"89",X"0D",X"00",X"00",X"49",X"1B",X"C3",X"1E",X"E2",X"1E",X"62",X"1B",X"00",X"00",
		X"CD",X"B6",X"39",X"01",X"01",X"FF",X"0A",X"00",X"FF",X"C9",X"CD",X"D9",X"3A",X"00",X"CD",X"7A",
		X"3A",X"01",X"0A",X"0A",X"C9",X"CD",X"E9",X"36",X"00",X"0F",X"00",X"00",X"B1",X"20",X"00",X"00",
		X"CD",X"FC",X"34",X"98",X"10",X"01",X"01",X"FF",X"01",X"06",X"01",X"01",X"06",X"FF",X"00",X"CD",
		X"E9",X"36",X"00",X"0F",X"00",X"00",X"CD",X"20",X"00",X"00",X"CD",X"E9",X"36",X"00",X"0F",X"00",
		X"00",X"B8",X"20",X"00",X"00",X"CD",X"E9",X"36",X"00",X"0F",X"00",X"00",X"BF",X"20",X"00",X"00",
		X"CD",X"E9",X"36",X"00",X"0F",X"00",X"00",X"C6",X"20",X"00",X"00",X"CD",X"E9",X"36",X"89",X"0D",
		X"00",X"18",X"94",X"1B",X"C4",X"1B",X"EB",X"1B",X"EB",X"1B",X"EB",X"1B",X"0B",X"1C",X"94",X"1B",
		X"94",X"1B",X"94",X"1B",X"C4",X"1B",X"94",X"1B",X"94",X"1B",X"C4",X"1B",X"0B",X"1C",X"EB",X"1C",
		X"00",X"00",X"CD",X"E9",X"36",X"89",X"0D",X"00",X"18",X"A4",X"1B",X"D1",X"1B",X"A4",X"1B",X"A4",
		X"1B",X"A4",X"1B",X"D1",X"1B",X"A4",X"1B",X"A4",X"1B",X"A4",X"1B",X"D1",X"1B",X"25",X"1C",X"25",
		X"1C",X"D1",X"1B",X"D1",X"1B",X"07",X"1D",X"00",X"00",X"CD",X"E9",X"36",X"89",X"0D",X"00",X"18",
		X"B4",X"1B",X"DE",X"1B",X"FB",X"1B",X"FB",X"1B",X"FB",X"1B",X"18",X"1C",X"B4",X"1B",X"B4",X"1B",
		X"B4",X"1B",X"DE",X"1B",X"35",X"1C",X"35",X"1C",X"DE",X"1B",X"18",X"1C",X"14",X"1D",X"00",X"00",
		X"CD",X"E9",X"36",X"89",X"0D",X"00",X"18",X"45",X"1C",X"00",X"00",X"CD",X"FC",X"34",X"98",X"10",
		X"00",X"01",X"FF",X"02",X"01",X"07",X"01",X"07",X"00",X"07",X"01",X"FE",X"00",X"CD",X"B6",X"39",
		X"01",X"05",X"FF",X"0A",X"0C",X"00",X"28",X"02",X"00",X"FF",X"C9",X"CD",X"7A",X"3A",X"00",X"0A",
		X"0A",X"CD",X"7A",X"3A",X"01",X"0A",X"0A",X"C9",X"CD",X"FC",X"34",X"F7",X"0F",X"00",X"01",X"FF",
		X"01",X"02",X"01",X"01",X"02",X"FF",X"00",X"CD",X"FC",X"34",X"98",X"10",X"01",X"01",X"00",X"0B",
		X"07",X"FF",X"00",X"CD",X"B6",X"39",X"01",X"05",X"FF",X"0A",X"0C",X"00",X"3C",X"02",X"00",X"FF",
		X"C9",X"CD",X"FC",X"34",X"F7",X"0F",X"00",X"01",X"FF",X"01",X"01",X"01",X"01",X"01",X"FF",X"00",
		X"CD",X"B6",X"39",X"01",X"05",X"FF",X"0A",X"0C",X"00",X"50",X"02",X"00",X"FF",X"C9",X"CD",X"FC",
		X"34",X"F7",X"0F",X"00",X"01",X"FF",X"01",X"03",X"01",X"01",X"03",X"FF",X"00",X"CD",X"B6",X"39",
		X"10",X"00",X"FF",X"16",X"03",X"0A",X"0D",X"04",X"00",X"FF",X"C9",X"CD",X"02",X"3B",X"00",X"16",
		X"04",X"C9",X"CD",X"6E",X"38",X"98",X"10",X"00",X"01",X"CD",X"E9",X"36",X"89",X"0D",X"00",X"18",
		X"D4",X"20",X"E7",X"20",X"0F",X"21",X"2B",X"21",X"0F",X"21",X"32",X"21",X"E7",X"20",X"39",X"21",
		X"6A",X"21",X"E7",X"20",X"0F",X"21",X"2B",X"21",X"0F",X"21",X"32",X"21",X"E7",X"20",X"39",X"21",
		X"7A",X"21",X"CC",X"23",X"6A",X"24",X"CC",X"23",X"E7",X"24",X"3E",X"25",X"CC",X"23",X"6A",X"24",
		X"CC",X"23",X"E7",X"24",X"6C",X"25",X"00",X"00",X"C9",X"CD",X"E9",X"36",X"89",X"0D",X"00",X"18",
		X"87",X"21",X"B3",X"21",X"62",X"22",X"B3",X"21",X"62",X"22",X"EB",X"23",X"5D",X"24",X"86",X"24",
		X"EB",X"23",X"5D",X"24",X"D1",X"24",X"EB",X"23",X"4E",X"25",X"EB",X"23",X"5D",X"24",X"86",X"24",
		X"EB",X"23",X"5D",X"24",X"D1",X"24",X"EB",X"23",X"7C",X"25",X"00",X"00",X"CD",X"E9",X"36",X"89",
		X"0D",X"00",X"18",X"69",X"22",X"7C",X"22",X"7C",X"22",X"DE",X"22",X"DE",X"22",X"8E",X"21",X"8E",
		X"21",X"F1",X"22",X"8F",X"22",X"8F",X"22",X"A2",X"22",X"7C",X"22",X"C7",X"22",X"7C",X"22",X"7C",
		X"22",X"DE",X"22",X"DE",X"22",X"8E",X"21",X"8E",X"21",X"F1",X"22",X"8F",X"22",X"8F",X"22",X"A2",
		X"22",X"7C",X"22",X"D7",X"22",X"FE",X"23",X"FE",X"23",X"2A",X"24",X"A5",X"24",X"2A",X"24",X"CA",
		X"24",X"FE",X"23",X"FE",X"23",X"2A",X"24",X"FA",X"24",X"5E",X"25",X"FE",X"23",X"FE",X"23",X"2A",
		X"24",X"A5",X"24",X"2A",X"24",X"CA",X"24",X"FE",X"23",X"FE",X"23",X"2A",X"24",X"FA",X"24",X"83",
		X"25",X"00",X"00",X"CD",X"E9",X"36",X"89",X"0D",X"00",X"18",X"16",X"23",X"1D",X"23",X"54",X"23",
		X"54",X"23",X"67",X"23",X"C5",X"23",X"1D",X"23",X"54",X"23",X"54",X"23",X"67",X"23",X"C5",X"23",
		X"11",X"24",X"43",X"24",X"43",X"24",X"50",X"24",X"50",X"24",X"43",X"24",X"43",X"24",X"11",X"24",
		X"43",X"24",X"43",X"24",X"2E",X"25",X"65",X"25",X"11",X"24",X"43",X"24",X"43",X"24",X"50",X"24",
		X"50",X"24",X"43",X"24",X"43",X"24",X"11",X"24",X"43",X"24",X"43",X"24",X"2E",X"25",X"65",X"25",
		X"00",X"00",X"CD",X"E9",X"36",X"89",X"0D",X"00",X"18",X"93",X"25",X"FE",X"23",X"FE",X"23",X"2A",
		X"24",X"A5",X"24",X"2A",X"24",X"CA",X"24",X"FE",X"23",X"FE",X"23",X"2A",X"24",X"FA",X"24",X"5E",
		X"25",X"FE",X"23",X"FE",X"23",X"2A",X"24",X"A5",X"24",X"2A",X"24",X"CA",X"24",X"FE",X"23",X"FE",
		X"23",X"2A",X"24",X"FA",X"24",X"00",X"00",X"CD",X"E9",X"36",X"89",X"0D",X"00",X"18",X"65",X"25",
		X"11",X"24",X"43",X"24",X"43",X"24",X"50",X"24",X"50",X"24",X"43",X"24",X"43",X"24",X"11",X"24",
		X"43",X"24",X"43",X"24",X"2E",X"25",X"00",X"00",X"CD",X"B6",X"39",X"01",X"01",X"FF",X"0A",X"02",
		X"00",X"A9",X"02",X"00",X"FF",X"C9",X"CD",X"7A",X"3A",X"00",X"0A",X"0A",X"C9",X"CD",X"FC",X"34",
		X"98",X"10",X"00",X"01",X"04",X"04",X"01",X"03",X"02",X"02",X"FF",X"01",X"03",X"00",X"05",X"01",
		X"FE",X"00",X"CD",X"B6",X"39",X"01",X"03",X"FF",X"0A",X"08",X"00",X"FA",X"02",X"00",X"FF",X"C9",
		X"CD",X"B1",X"3A",X"00",X"00",X"CD",X"7A",X"3A",X"01",X"0A",X"0A",X"C9",X"CD",X"0D",X"36",X"5B",
		X"12",X"00",X"02",X"FF",X"02",X"FA",X"00",X"02",X"13",X"01",X"02",X"31",X"01",X"02",X"57",X"01",
		X"02",X"88",X"01",X"02",X"CA",X"01",X"02",X"25",X"02",X"02",X"AF",X"02",X"0A",X"94",X"03",X"02",
		X"AF",X"02",X"02",X"25",X"02",X"02",X"CA",X"01",X"02",X"88",X"01",X"02",X"57",X"01",X"02",X"31",
		X"01",X"02",X"13",X"01",X"02",X"FA",X"00",X"02",X"00",X"00",X"00",X"CD",X"FC",X"34",X"98",X"10",
		X"01",X"01",X"00",X"01",X"01",X"04",X"01",X"11",X"FC",X"01",X"01",X"FC",X"01",X"05",X"04",X"01",
		X"01",X"04",X"01",X"11",X"FC",X"01",X"01",X"FC",X"01",X"01",X"04",X"00",X"CD",X"B6",X"39",X"01",
		X"03",X"FF",X"0A",X"0A",X"00",X"C3",X"02",X"01",X"FF",X"C9",X"CD",X"7A",X"3A",X"00",X"0A",X"0A",
		X"CD",X"7A",X"3A",X"01",X"00",X"00",X"C9",X"CD",X"FC",X"34",X"54",X"13",X"00",X"01",X"00",X"01",
		X"03",X"01",X"01",X"02",X"FF",X"01",X"02",X"01",X"01",X"02",X"FF",X"01",X"02",X"01",X"01",X"02",
		X"FF",X"01",X"02",X"01",X"01",X"01",X"FF",X"01",X"02",X"01",X"01",X"01",X"FF",X"01",X"01",X"01",
		X"01",X"01",X"FF",X"01",X"01",X"01",X"01",X"01",X"FF",X"01",X"01",X"01",X"01",X"01",X"FF",X"01",
		X"01",X"01",X"01",X"01",X"FF",X"01",X"01",X"01",X"01",X"01",X"FF",X"01",X"01",X"01",X"01",X"01",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"FF",X"01",X"01",X"01",X"01",X"01",X"FF",X"01",X"01",X"01",
		X"01",X"01",X"FF",X"01",X"01",X"01",X"01",X"01",X"FF",X"01",X"01",X"01",X"01",X"01",X"FF",X"01",
		X"01",X"01",X"01",X"01",X"FF",X"01",X"01",X"01",X"01",X"01",X"FF",X"01",X"01",X"01",X"01",X"01",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"FF",X"01",X"01",X"01",X"01",X"01",X"FF",X"01",X"01",X"01",
		X"01",X"01",X"FF",X"01",X"01",X"01",X"01",X"01",X"FF",X"01",X"01",X"01",X"01",X"01",X"FF",X"01",
		X"01",X"01",X"01",X"01",X"FF",X"01",X"01",X"01",X"01",X"01",X"FF",X"01",X"01",X"01",X"01",X"01",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"FF",X"01",X"01",X"01",X"01",X"01",X"FF",X"01",X"01",X"01",
		X"01",X"01",X"FF",X"00",X"CD",X"FC",X"34",X"98",X"10",X"01",X"02",X"00",X"16",X"03",X"EF",X"FF",
		X"00",X"CD",X"B6",X"39",X"01",X"03",X"FF",X"0A",X"03",X"00",X"CC",X"02",X"00",X"FF",X"C9",X"CD",
		X"0D",X"36",X"37",X"15",X"00",X"02",X"00",X"02",X"CC",X"00",X"02",X"C4",X"00",X"02",X"BD",X"00",
		X"02",X"B7",X"00",X"02",X"B1",X"00",X"02",X"AC",X"00",X"02",X"A7",X"00",X"02",X"BD",X"00",X"02",
		X"C4",X"00",X"02",X"CC",X"00",X"02",X"D3",X"00",X"02",X"DC",X"00",X"02",X"E5",X"00",X"02",X"DC",
		X"00",X"02",X"D3",X"00",X"02",X"CC",X"00",X"02",X"C4",X"00",X"02",X"BD",X"00",X"02",X"B7",X"00",
		X"02",X"CC",X"00",X"02",X"D3",X"00",X"02",X"DC",X"00",X"02",X"E5",X"00",X"02",X"EF",X"00",X"02",
		X"FA",X"00",X"02",X"EF",X"00",X"02",X"E5",X"00",X"02",X"DC",X"00",X"02",X"D3",X"00",X"02",X"CC",
		X"00",X"02",X"C4",X"00",X"02",X"DC",X"00",X"02",X"E5",X"00",X"02",X"EF",X"00",X"02",X"FA",X"00",
		X"02",X"06",X"01",X"02",X"13",X"01",X"02",X"06",X"01",X"02",X"FA",X"00",X"02",X"EF",X"00",X"02",
		X"E5",X"00",X"02",X"DC",X"00",X"02",X"D3",X"00",X"02",X"EF",X"00",X"02",X"FA",X"00",X"02",X"06",
		X"01",X"02",X"13",X"01",X"02",X"21",X"01",X"02",X"31",X"01",X"02",X"21",X"01",X"02",X"13",X"01",
		X"02",X"06",X"01",X"02",X"FA",X"00",X"02",X"EF",X"00",X"02",X"E5",X"00",X"02",X"06",X"01",X"02",
		X"13",X"01",X"02",X"21",X"01",X"02",X"31",X"01",X"02",X"43",X"01",X"02",X"57",X"01",X"02",X"43",
		X"01",X"02",X"31",X"01",X"02",X"21",X"01",X"02",X"13",X"01",X"02",X"06",X"01",X"02",X"FA",X"00",
		X"02",X"21",X"01",X"02",X"31",X"01",X"02",X"43",X"01",X"02",X"57",X"01",X"02",X"6E",X"01",X"02",
		X"88",X"01",X"02",X"6E",X"01",X"02",X"57",X"01",X"02",X"43",X"01",X"02",X"31",X"01",X"02",X"21",
		X"01",X"02",X"13",X"01",X"02",X"43",X"01",X"02",X"57",X"01",X"02",X"6E",X"01",X"02",X"88",X"01",
		X"02",X"A7",X"01",X"02",X"CA",X"01",X"02",X"A7",X"01",X"02",X"88",X"01",X"02",X"6E",X"01",X"02",
		X"57",X"01",X"02",X"43",X"01",X"02",X"31",X"01",X"02",X"6E",X"01",X"02",X"88",X"01",X"02",X"A7",
		X"01",X"02",X"CA",X"01",X"02",X"F4",X"01",X"02",X"25",X"02",X"02",X"F4",X"01",X"02",X"CA",X"01",
		X"02",X"A7",X"01",X"02",X"88",X"01",X"02",X"6E",X"01",X"02",X"57",X"01",X"02",X"A7",X"01",X"02",
		X"CA",X"01",X"02",X"F4",X"01",X"02",X"25",X"02",X"02",X"63",X"02",X"02",X"AF",X"02",X"02",X"63",
		X"02",X"02",X"25",X"02",X"02",X"F4",X"01",X"02",X"CA",X"01",X"02",X"A7",X"01",X"02",X"88",X"01",
		X"02",X"F4",X"01",X"02",X"25",X"02",X"02",X"63",X"02",X"02",X"AF",X"02",X"02",X"11",X"03",X"02",
		X"94",X"03",X"02",X"11",X"03",X"02",X"AF",X"02",X"02",X"63",X"02",X"02",X"25",X"02",X"02",X"F4",
		X"01",X"02",X"CA",X"01",X"02",X"AF",X"02",X"02",X"57",X"01",X"02",X"E5",X"00",X"02",X"AC",X"00",
		X"02",X"89",X"00",X"02",X"72",X"00",X"02",X"62",X"00",X"02",X"56",X"00",X"02",X"4C",X"00",X"02",
		X"45",X"00",X"02",X"3E",X"00",X"02",X"AF",X"02",X"02",X"57",X"01",X"02",X"E5",X"00",X"02",X"AC",
		X"00",X"02",X"89",X"00",X"02",X"72",X"00",X"02",X"62",X"00",X"02",X"56",X"00",X"02",X"4C",X"00",
		X"02",X"45",X"00",X"02",X"3E",X"00",X"00",X"CD",X"FC",X"34",X"98",X"10",X"01",X"01",X"00",X"02",
		X"01",X"04",X"02",X"7E",X"FF",X"02",X"01",X"01",X"01",X"14",X"FE",X"02",X"01",X"01",X"01",X"14",
		X"FA",X"00",X"CD",X"B6",X"39",X"01",X"03",X"FF",X"0A",X"0A",X"00",X"7D",X"02",X"00",X"FF",X"C9",
		X"CD",X"B1",X"3A",X"00",X"00",X"C9",X"CD",X"0D",X"36",X"98",X"10",X"00",X"02",X"FF",X"02",X"57",
		X"01",X"02",X"31",X"01",X"02",X"13",X"01",X"02",X"FA",X"00",X"02",X"E5",X"00",X"02",X"D3",X"00",
		X"02",X"C4",X"00",X"02",X"B7",X"00",X"02",X"AC",X"00",X"02",X"A2",X"00",X"02",X"99",X"00",X"02",
		X"91",X"00",X"02",X"89",X"00",X"02",X"91",X"00",X"02",X"99",X"00",X"02",X"A2",X"00",X"02",X"AC",
		X"00",X"02",X"B7",X"00",X"02",X"C4",X"00",X"02",X"D3",X"00",X"02",X"E5",X"00",X"02",X"FA",X"00",
		X"02",X"13",X"01",X"02",X"31",X"01",X"00",X"CD",X"B6",X"39",X"01",X"03",X"FF",X"0A",X"03",X"00",
		X"00",X"02",X"00",X"FF",X"C9",X"CD",X"B1",X"3A",X"00",X"00",X"CD",X"B1",X"3A",X"01",X"0A",X"C9",
		X"CD",X"0D",X"36",X"03",X"16",X"00",X"02",X"FF",X"03",X"00",X"00",X"02",X"E8",X"02",X"02",X"BE",
		X"01",X"02",X"3F",X"01",X"02",X"F8",X"00",X"02",X"CB",X"00",X"02",X"AC",X"00",X"02",X"95",X"00",
		X"03",X"00",X"00",X"02",X"CB",X"00",X"02",X"F8",X"00",X"02",X"3F",X"01",X"02",X"BE",X"01",X"02",
		X"E8",X"02",X"00",X"CD",X"0D",X"36",X"98",X"10",X"01",X"01",X"FF",X"03",X"00",X"0E",X"0B",X"03",
		X"00",X"0A",X"0B",X"00",X"CD",X"E9",X"36",X"98",X"10",X"00",X"FF",X"9A",X"25",X"9E",X"25",X"9E",
		X"25",X"AE",X"25",X"D0",X"25",X"D0",X"25",X"E0",X"25",X"02",X"26",X"02",X"26",X"12",X"26",X"43",
		X"26",X"50",X"26",X"AF",X"28",X"B6",X"28",X"C6",X"28",X"B6",X"28",X"CA",X"28",X"D7",X"28",X"E4",
		X"28",X"D7",X"28",X"E4",X"28",X"D7",X"28",X"E4",X"28",X"D7",X"28",X"C6",X"28",X"AF",X"28",X"AF",
		X"28",X"B6",X"28",X"F1",X"28",X"B6",X"28",X"04",X"29",X"00",X"00",X"CD",X"E9",X"36",X"98",X"10",
		X"00",X"FF",X"A8",X"26",X"AF",X"26",X"B9",X"26",X"BD",X"26",X"CA",X"26",X"BD",X"26",X"D4",X"26",
		X"DE",X"26",X"D4",X"26",X"E2",X"26",X"AF",X"26",X"EC",X"26",X"F0",X"26",X"03",X"27",X"F0",X"26",
		X"07",X"27",X"AF",X"26",X"B9",X"26",X"BD",X"26",X"CA",X"26",X"BD",X"26",X"20",X"27",X"43",X"26",
		X"3C",X"27",X"AF",X"28",X"63",X"29",X"C6",X"28",X"63",X"29",X"73",X"29",X"80",X"29",X"8D",X"29",
		X"80",X"29",X"8D",X"29",X"80",X"29",X"8D",X"29",X"80",X"29",X"91",X"29",X"AF",X"28",X"63",X"29",
		X"A4",X"29",X"E7",X"29",X"FD",X"29",X"E7",X"29",X"16",X"2A",X"00",X"00",X"CD",X"E9",X"36",X"98",
		X"10",X"00",X"FF",X"79",X"27",X"80",X"27",X"8D",X"27",X"80",X"27",X"97",X"27",X"A1",X"27",X"97",
		X"27",X"A5",X"27",X"B2",X"27",X"C5",X"27",X"B2",X"27",X"C9",X"27",X"79",X"27",X"80",X"27",X"8D",
		X"27",X"80",X"27",X"DF",X"27",X"32",X"2A",X"32",X"2A",X"32",X"2A",X"4B",X"2A",X"4B",X"2A",X"4B",
		X"2A",X"4B",X"2A",X"32",X"2A",X"32",X"2A",X"32",X"2A",X"32",X"2A",X"64",X"2A",X"7D",X"2A",X"96",
		X"2A",X"7D",X"2A",X"64",X"2A",X"00",X"00",X"CD",X"E9",X"36",X"98",X"10",X"00",X"FF",X"34",X"28",
		X"3E",X"28",X"3E",X"28",X"4E",X"28",X"4E",X"28",X"5B",X"28",X"5B",X"28",X"5B",X"28",X"6B",X"28",
		X"6B",X"28",X"3E",X"28",X"3E",X"28",X"3E",X"28",X"4E",X"28",X"4E",X"28",X"78",X"28",X"AF",X"2A",
		X"CB",X"2A",X"D2",X"2A",X"D2",X"2A",X"DF",X"2A",X"EC",X"2A",X"DF",X"2A",X"76",X"2B",X"AF",X"2A",
		X"F0",X"2A",X"03",X"2B",X"16",X"2B",X"03",X"2B",X"20",X"2B",X"2A",X"2B",X"3D",X"2B",X"56",X"2B",
		X"3D",X"2B",X"6C",X"2B",X"2A",X"2B",X"00",X"00",X"CD",X"E9",X"36",X"98",X"10",X"00",X"FF",X"AF",
		X"28",X"B6",X"28",X"C6",X"28",X"B6",X"28",X"CA",X"28",X"D7",X"28",X"E4",X"28",X"D7",X"28",X"E4",
		X"28",X"D7",X"28",X"E4",X"28",X"D7",X"28",X"C6",X"28",X"AF",X"28",X"AF",X"28",X"B6",X"28",X"F1",
		X"28",X"B6",X"28",X"04",X"29",X"9A",X"25",X"9E",X"25",X"9E",X"25",X"AE",X"25",X"D0",X"25",X"D0",
		X"25",X"E0",X"25",X"02",X"26",X"02",X"26",X"12",X"26",X"43",X"26",X"50",X"26",X"00",X"00",X"CD",
		X"E9",X"36",X"98",X"10",X"00",X"FF",X"56",X"29",X"63",X"29",X"C6",X"28",X"63",X"29",X"73",X"29",
		X"80",X"29",X"8D",X"29",X"80",X"29",X"8D",X"29",X"80",X"29",X"8D",X"29",X"80",X"29",X"91",X"29",
		X"AF",X"28",X"63",X"29",X"A4",X"29",X"E7",X"29",X"FD",X"29",X"E7",X"29",X"16",X"2A",X"EC",X"2A",
		X"AF",X"26",X"B9",X"26",X"BD",X"26",X"CA",X"26",X"BD",X"26",X"D4",X"26",X"DE",X"26",X"D4",X"26",
		X"E2",X"26",X"AF",X"26",X"EC",X"26",X"F0",X"26",X"03",X"27",X"F0",X"26",X"07",X"27",X"AF",X"26",
		X"B9",X"26",X"BD",X"26",X"CA",X"26",X"BD",X"26",X"20",X"27",X"43",X"26",X"3C",X"27",X"00",X"00",
		X"CD",X"E9",X"36",X"98",X"10",X"00",X"FF",X"32",X"2A",X"32",X"2A",X"32",X"2A",X"4B",X"2A",X"4B",
		X"2A",X"4B",X"2A",X"4B",X"2A",X"32",X"2A",X"32",X"2A",X"32",X"2A",X"32",X"2A",X"64",X"2A",X"7D",
		X"2A",X"96",X"2A",X"7D",X"2A",X"64",X"2A",X"79",X"27",X"80",X"27",X"8D",X"27",X"80",X"27",X"97",
		X"27",X"A1",X"27",X"97",X"27",X"A5",X"27",X"B2",X"27",X"C5",X"27",X"B2",X"27",X"C9",X"27",X"79",
		X"27",X"80",X"27",X"8D",X"27",X"80",X"27",X"DF",X"27",X"00",X"00",X"CD",X"E9",X"36",X"98",X"10",
		X"00",X"FF",X"AF",X"2A",X"CB",X"2A",X"D2",X"2A",X"D2",X"2A",X"DF",X"2A",X"EC",X"2A",X"DF",X"2A",
		X"76",X"2B",X"AF",X"2A",X"F0",X"2A",X"03",X"2B",X"16",X"2B",X"03",X"2B",X"20",X"2B",X"2A",X"2B",
		X"3D",X"2B",X"56",X"2B",X"3D",X"2B",X"6C",X"2B",X"2A",X"2B",X"9A",X"25",X"3E",X"28",X"3E",X"28",
		X"4E",X"28",X"4E",X"28",X"5B",X"28",X"5B",X"28",X"5B",X"28",X"6B",X"28",X"6B",X"28",X"3E",X"28",
		X"3E",X"28",X"3E",X"28",X"4E",X"28",X"4E",X"28",X"78",X"28",X"00",X"00",X"CD",X"E9",X"36",X"98",
		X"10",X"00",X"FF",X"F4",X"2B",X"FE",X"2B",X"05",X"2C",X"0F",X"2C",X"1C",X"2C",X"23",X"2C",X"2D",
		X"2C",X"37",X"2C",X"41",X"2C",X"4B",X"2C",X"52",X"2C",X"5F",X"2C",X"69",X"2C",X"00",X"00",X"CD",
		X"E9",X"36",X"98",X"10",X"00",X"FF",X"37",X"2C",X"6D",X"2C",X"41",X"2C",X"52",X"2C",X"74",X"2C",
		X"5F",X"2C",X"7B",X"2C",X"F4",X"2B",X"05",X"2C",X"85",X"2C",X"0F",X"2C",X"23",X"2C",X"8C",X"2C",
		X"00",X"00",X"CD",X"E9",X"36",X"98",X"10",X"00",X"FF",X"90",X"2C",X"12",X"2D",X"1C",X"2D",X"12",
		X"2D",X"20",X"2D",X"12",X"2D",X"24",X"2D",X"12",X"2D",X"28",X"2D",X"00",X"00",X"CD",X"E9",X"36",
		X"98",X"10",X"00",X"FF",X"59",X"2D",X"69",X"2D",X"70",X"2D",X"7D",X"2D",X"59",X"2D",X"81",X"2D",
		X"70",X"2D",X"88",X"2D",X"00",X"00",X"CD",X"E9",X"36",X"98",X"10",X"00",X"FF",X"E6",X"2D",X"ED",
		X"2D",X"0C",X"2E",X"1C",X"2E",X"ED",X"2D",X"2C",X"2E",X"1C",X"2E",X"ED",X"2D",X"0C",X"2E",X"39",
		X"2E",X"79",X"2E",X"ED",X"2D",X"0C",X"2E",X"1C",X"2E",X"ED",X"2D",X"2C",X"2E",X"1C",X"2E",X"ED",
		X"2D",X"0C",X"2E",X"39",X"2E",X"79",X"2E",X"ED",X"2D",X"0C",X"2E",X"1C",X"2E",X"ED",X"2D",X"2C",
		X"2E",X"1C",X"2E",X"ED",X"2D",X"0C",X"2E",X"39",X"2E",X"00",X"00",X"CD",X"E9",X"36",X"98",X"10",
		X"00",X"FF",X"80",X"2E",X"84",X"2E",X"A9",X"2E",X"84",X"2E",X"CB",X"2E",X"F0",X"2E",X"84",X"2E",
		X"A9",X"2E",X"84",X"2E",X"CB",X"2E",X"F0",X"2E",X"84",X"2E",X"A9",X"2E",X"84",X"2E",X"CB",X"2E",
		X"00",X"00",X"CD",X"E9",X"36",X"98",X"10",X"00",X"FF",X"80",X"2E",X"95",X"2F",X"CC",X"2F",X"95",
		X"2F",X"03",X"30",X"31",X"30",X"95",X"2F",X"CC",X"2F",X"95",X"2F",X"03",X"30",X"31",X"30",X"95",
		X"2F",X"CC",X"2F",X"95",X"2F",X"03",X"30",X"00",X"00",X"CD",X"E9",X"36",X"98",X"10",X"00",X"FF",
		X"F7",X"2E",X"FB",X"2E",X"2C",X"2F",X"FB",X"2E",X"5D",X"2F",X"91",X"2F",X"FB",X"2E",X"2C",X"2F",
		X"FB",X"2E",X"5D",X"2F",X"91",X"2F",X"FB",X"2E",X"2C",X"2F",X"FB",X"2E",X"5D",X"2F",X"00",X"00",
		X"CD",X"0D",X"36",X"03",X"1A",X"00",X"02",X"FF",X"03",X"00",X"00",X"02",X"D0",X"05",X"02",X"7D",
		X"03",X"02",X"7E",X"02",X"02",X"F0",X"01",X"02",X"96",X"01",X"02",X"57",X"01",X"02",X"2A",X"01",
		X"03",X"00",X"00",X"02",X"96",X"01",X"02",X"F0",X"01",X"02",X"7E",X"02",X"02",X"7D",X"03",X"02",
		X"D0",X"05",X"00",X"CD",X"0D",X"36",X"98",X"10",X"01",X"01",X"FF",X"03",X"00",X"0E",X"08",X"03",
		X"00",X"0A",X"08",X"00",X"CD",X"B6",X"39",X"01",X"02",X"FF",X"0A",X"01",X"00",X"DE",X"02",X"01",
		X"FF",X"C9",X"CD",X"7A",X"3A",X"00",X"0A",X"0A",X"C9",X"CD",X"FC",X"34",X"98",X"10",X"00",X"01",
		X"00",X"04",X"01",X"03",X"01",X"34",X"00",X"04",X"01",X"FD",X"00",X"CD",X"B6",X"39",X"01",X"02",
		X"FF",X"0A",X"01",X"00",X"AA",X"02",X"01",X"FF",X"C9",X"CD",X"FC",X"34",X"98",X"10",X"00",X"01",
		X"00",X"01",X"3C",X"00",X"04",X"01",X"03",X"01",X"34",X"00",X"04",X"01",X"FD",X"00",X"CD",X"B6",
		X"39",X"01",X"02",X"FF",X"0A",X"01",X"00",X"7B",X"02",X"01",X"FF",X"C9",X"CD",X"FC",X"34",X"98",
		X"10",X"00",X"01",X"00",X"01",X"78",X"00",X"04",X"01",X"03",X"01",X"34",X"00",X"04",X"01",X"FD",
		X"00",X"CD",X"B6",X"39",X"01",X"02",X"FF",X"0A",X"01",X"00",X"52",X"02",X"01",X"FF",X"C9",X"CD",
		X"FC",X"34",X"98",X"10",X"00",X"01",X"00",X"01",X"B4",X"00",X"04",X"01",X"03",X"01",X"34",X"00",
		X"04",X"01",X"FD",X"00",X"CD",X"B6",X"39",X"01",X"02",X"FF",X"0A",X"01",X"00",X"2D",X"02",X"01",
		X"FF",X"C9",X"CD",X"FC",X"34",X"98",X"10",X"00",X"01",X"00",X"01",X"F0",X"00",X"04",X"01",X"03",
		X"01",X"34",X"00",X"04",X"01",X"FD",X"00",X"CD",X"B6",X"39",X"01",X"02",X"FF",X"0A",X"01",X"00",
		X"0C",X"02",X"01",X"FF",X"C9",X"CD",X"FC",X"34",X"98",X"10",X"00",X"01",X"00",X"01",X"C8",X"00",
		X"01",X"64",X"00",X"04",X"01",X"03",X"01",X"34",X"00",X"04",X"01",X"FD",X"00",X"CD",X"E9",X"36",
		X"98",X"10",X"00",X"FF",X"E8",X"31",X"EA",X"30",X"EF",X"31",X"08",X"32",X"EF",X"31",X"21",X"32",
		X"EA",X"30",X"EF",X"31",X"08",X"32",X"EF",X"31",X"21",X"32",X"EA",X"30",X"EF",X"31",X"08",X"32",
		X"EF",X"31",X"21",X"32",X"00",X"00",X"CD",X"E9",X"36",X"98",X"10",X"00",X"00",X"AF",X"2A",X"C2",
		X"2B",X"00",X"00",X"CD",X"E9",X"36",X"98",X"10",X"00",X"00",X"32",X"2A",X"DB",X"2B",X"00",X"00",
		X"0D",X"77",X"00",X"0D",X"7F",X"00",X"05",X"86",X"00",X"05",X"7F",X"00",X"05",X"86",X"00",X"05",
		X"8E",X"00",X"0D",X"96",X"00",X"0D",X"9F",X"00",X"00",X"0D",X"8E",X"00",X"0D",X"96",X"00",X"05",
		X"9F",X"00",X"05",X"96",X"00",X"05",X"9F",X"00",X"05",X"A9",X"00",X"0D",X"B3",X"00",X"0D",X"BE",
		X"00",X"00",X"05",X"FD",X"00",X"05",X"EF",X"00",X"05",X"E1",X"00",X"05",X"D5",X"00",X"05",X"C9",
		X"00",X"05",X"BE",X"00",X"05",X"B3",X"00",X"05",X"A9",X"00",X"05",X"9F",X"00",X"05",X"96",X"00",
		X"00",X"05",X"9F",X"00",X"21",X"00",X"00",X"05",X"D5",X"00",X"05",X"D5",X"00",X"0D",X"E1",X"00",
		X"0D",X"D5",X"00",X"00",X"23",X"00",X"00",X"05",X"77",X"00",X"05",X"77",X"00",X"0D",X"77",X"00",
		X"0D",X"77",X"00",X"00",X"23",X"00",X"00",X"05",X"9F",X"00",X"05",X"9F",X"00",X"0D",X"9F",X"00",
		X"0D",X"9F",X"00",X"00",X"23",X"00",X"00",X"05",X"BE",X"00",X"05",X"BE",X"00",X"0D",X"BE",X"00",
		X"0D",X"BE",X"00",X"00",X"23",X"00",X"00",X"0D",X"77",X"00",X"23",X"00",X"00",X"0D",X"77",X"00",
		X"00",X"23",X"00",X"00",X"0D",X"9F",X"00",X"23",X"00",X"00",X"0D",X"9F",X"00",X"00",X"23",X"00",
		X"00",X"0D",X"BE",X"00",X"23",X"00",X"00",X"0D",X"BE",X"00",X"00",X"23",X"00",X"00",X"05",X"7F",
		X"00",X"05",X"7F",X"00",X"0D",X"7F",X"00",X"0D",X"7F",X"00",X"00",X"23",X"00",X"00",X"05",X"B3",
		X"00",X"05",X"B3",X"00",X"0D",X"B3",X"00",X"0D",X"B3",X"00",X"00",X"23",X"00",X"00",X"0D",X"7F",
		X"00",X"23",X"00",X"00",X"0D",X"7F",X"00",X"00",X"23",X"00",X"00",X"0D",X"B3",X"00",X"23",X"00",
		X"00",X"0D",X"B3",X"00",X"00",X"23",X"00",X"00",X"05",X"A9",X"00",X"05",X"A9",X"00",X"0D",X"A9",
		X"00",X"0D",X"A9",X"00",X"00",X"23",X"00",X"00",X"05",X"C9",X"00",X"05",X"C9",X"00",X"0D",X"C9",
		X"00",X"0D",X"C9",X"00",X"00",X"19",X"BC",X"03",X"0F",X"FB",X"04",X"0F",X"BC",X"03",X"07",X"F4",
		X"03",X"07",X"BC",X"03",X"07",X"86",X"03",X"07",X"53",X"03",X"07",X"24",X"03",X"07",X"F6",X"02",
		X"19",X"CC",X"02",X"0F",X"F6",X"02",X"19",X"53",X"03",X"23",X"00",X"00",X"19",X"38",X"02",X"0F",
		X"7F",X"02",X"07",X"CC",X"02",X"07",X"7F",X"02",X"07",X"CC",X"02",X"07",X"F6",X"02",X"07",X"53",
		X"03",X"07",X"F6",X"02",X"07",X"CC",X"02",X"07",X"53",X"03",X"19",X"BC",X"03",X"0F",X"F6",X"02",
		X"19",X"FB",X"04",X"23",X"00",X"00",X"19",X"BC",X"03",X"0F",X"FB",X"04",X"0F",X"BC",X"03",X"07",
		X"F4",X"03",X"07",X"BC",X"03",X"07",X"53",X"03",X"07",X"F6",X"02",X"07",X"CC",X"02",X"07",X"7F",
		X"02",X"19",X"A4",X"02",X"0F",X"38",X"02",X"15",X"DE",X"01",X"0F",X"FA",X"01",X"0F",X"DE",X"01",
		X"15",X"7B",X"01",X"15",X"DE",X"01",X"15",X"AA",X"01",X"15",X"7F",X"02",X"0F",X"DE",X"01",X"07",
		X"FA",X"01",X"07",X"38",X"02",X"07",X"7F",X"02",X"07",X"CC",X"02",X"07",X"F6",X"02",X"07",X"53",
		X"03",X"0F",X"BC",X"03",X"23",X"00",X"00",X"15",X"FB",X"04",X"00",X"0D",X"77",X"00",X"05",X"7F",
		X"00",X"05",X"8E",X"00",X"05",X"9F",X"00",X"05",X"B3",X"00",X"05",X"BE",X"00",X"05",X"D5",X"00",
		X"0D",X"EF",X"00",X"27",X"00",X"00",X"00",X"0D",X"9F",X"00",X"27",X"00",X"00",X"25",X"00",X"00",
		X"15",X"3F",X"01",X"00",X"0D",X"BE",X"00",X"27",X"00",X"00",X"29",X"00",X"00",X"00",X"0D",X"C9",
		X"00",X"0D",X"BE",X"00",X"00",X"0D",X"A9",X"00",X"0D",X"9F",X"00",X"00",X"0D",X"B3",X"00",X"0D",
		X"BE",X"00",X"05",X"BE",X"00",X"05",X"B3",X"00",X"05",X"BE",X"00",X"05",X"C9",X"00",X"0D",X"D5",
		X"00",X"0D",X"EF",X"00",X"0D",X"FD",X"00",X"0D",X"EF",X"00",X"00",X"0D",X"77",X"07",X"0D",X"BE",
		X"00",X"0D",X"FB",X"04",X"0D",X"BE",X"00",X"0D",X"BC",X"03",X"0D",X"BE",X"00",X"0D",X"FB",X"04",
		X"0D",X"BE",X"00",X"0D",X"77",X"07",X"0D",X"BE",X"00",X"0D",X"FB",X"04",X"0D",X"BE",X"00",X"0D",
		X"BC",X"03",X"0D",X"BE",X"00",X"0D",X"FB",X"04",X"0D",X"BE",X"00",X"00",X"05",X"8E",X"00",X"05",
		X"7F",X"00",X"0D",X"8E",X"00",X"0D",X"9F",X"00",X"00",X"05",X"D5",X"00",X"21",X"00",X"00",X"05",
		X"FD",X"00",X"05",X"FD",X"00",X"0D",X"0C",X"01",X"0D",X"FD",X"00",X"00",X"23",X"00",X"00",X"0D",
		X"AA",X"01",X"23",X"00",X"00",X"0D",X"AA",X"01",X"23",X"00",X"00",X"0D",X"AA",X"01",X"23",X"00",
		X"00",X"0D",X"AA",X"01",X"00",X"0D",X"FB",X"04",X"0D",X"66",X"01",X"0D",X"53",X"03",X"0D",X"66",
		X"01",X"0D",X"7F",X"02",X"0D",X"66",X"01",X"0D",X"53",X"03",X"0D",X"66",X"01",X"00",X"0D",X"FD",
		X"00",X"05",X"C9",X"00",X"05",X"C9",X"00",X"0D",X"A9",X"00",X"0D",X"FD",X"00",X"05",X"9F",X"00",
		X"05",X"8E",X"00",X"05",X"9F",X"00",X"05",X"A9",X"00",X"0D",X"BE",X"00",X"0D",X"FD",X"00",X"0D",
		X"7F",X"00",X"05",X"7F",X"00",X"05",X"7F",X"00",X"0D",X"7F",X"00",X"0D",X"7F",X"00",X"0D",X"7F",
		X"00",X"0D",X"7F",X"00",X"0D",X"7F",X"00",X"0D",X"7F",X"00",X"00",X"0D",X"92",X"01",X"0D",X"52",
		X"01",X"0D",X"FD",X"00",X"0D",X"92",X"01",X"0D",X"FD",X"00",X"05",X"FD",X"00",X"05",X"FD",X"00",
		X"0D",X"FD",X"00",X"0D",X"3F",X"01",X"0D",X"92",X"01",X"05",X"92",X"01",X"05",X"92",X"01",X"0D",
		X"92",X"01",X"0D",X"92",X"01",X"0D",X"FD",X"00",X"0D",X"FD",X"00",X"0D",X"FD",X"00",X"0D",X"FD",
		X"00",X"00",X"0D",X"F4",X"03",X"05",X"FA",X"01",X"05",X"FA",X"01",X"0D",X"F4",X"03",X"0D",X"FA",
		X"01",X"0D",X"ED",X"05",X"05",X"F6",X"02",X"05",X"F6",X"02",X"0D",X"F6",X"02",X"0D",X"F6",X"02",
		X"0D",X"F4",X"03",X"05",X"FA",X"01",X"05",X"FA",X"01",X"0D",X"F4",X"03",X"0D",X"FA",X"01",X"05",
		X"FA",X"01",X"05",X"18",X"02",X"05",X"38",X"02",X"05",X"5A",X"02",X"05",X"7F",X"02",X"05",X"A4",
		X"02",X"05",X"CC",X"02",X"05",X"53",X"03",X"00",X"05",X"A9",X"00",X"05",X"9F",X"00",X"05",X"A9",
		X"00",X"05",X"B3",X"00",X"0D",X"BE",X"00",X"0D",X"C9",X"00",X"05",X"D5",X"00",X"05",X"C9",X"00",
		X"05",X"D5",X"00",X"05",X"E1",X"00",X"00",X"0D",X"EF",X"00",X"0D",X"FD",X"00",X"05",X"0C",X"01",
		X"05",X"FD",X"00",X"05",X"0C",X"01",X"05",X"1C",X"01",X"05",X"2D",X"01",X"05",X"1C",X"01",X"05",
		X"0C",X"01",X"00",X"05",X"C9",X"00",X"05",X"BE",X"00",X"05",X"C9",X"00",X"05",X"D5",X"00",X"0D",
		X"E1",X"00",X"0D",X"EF",X"00",X"05",X"FD",X"00",X"05",X"EF",X"00",X"05",X"FD",X"00",X"05",X"0C",
		X"01",X"00",X"0D",X"1C",X"01",X"0D",X"2D",X"01",X"05",X"3F",X"01",X"05",X"2D",X"01",X"05",X"3F",
		X"01",X"05",X"52",X"01",X"05",X"66",X"01",X"05",X"52",X"01",X"05",X"3F",X"01",X"05",X"2D",X"01",
		X"05",X"1C",X"01",X"05",X"0C",X"01",X"00",X"0D",X"D5",X"00",X"05",X"D5",X"00",X"05",X"D5",X"00",
		X"0D",X"8E",X"00",X"0D",X"D5",X"00",X"0D",X"C9",X"00",X"05",X"C9",X"00",X"05",X"C9",X"00",X"13",
		X"86",X"00",X"05",X"7F",X"00",X"05",X"6A",X"00",X"05",X"71",X"00",X"05",X"77",X"00",X"0D",X"7F",
		X"00",X"0D",X"8E",X"00",X"0D",X"9F",X"00",X"27",X"00",X"00",X"00",X"23",X"00",X"00",X"0D",X"52",
		X"01",X"23",X"00",X"00",X"0D",X"52",X"01",X"23",X"00",X"00",X"0D",X"3F",X"01",X"23",X"00",X"00",
		X"0D",X"3F",X"01",X"23",X"00",X"00",X"0D",X"3F",X"01",X"23",X"00",X"00",X"0D",X"52",X"01",X"0D",
		X"3F",X"01",X"27",X"00",X"00",X"00",X"0D",X"53",X"03",X"0D",X"DE",X"01",X"0D",X"53",X"03",X"0D",
		X"DE",X"01",X"0D",X"86",X"03",X"0D",X"18",X"02",X"0D",X"86",X"03",X"0D",X"92",X"01",X"0D",X"53",
		X"03",X"23",X"00",X"00",X"0D",X"A7",X"06",X"0D",X"A7",X"06",X"0F",X"FB",X"04",X"0B",X"FB",X"04",
		X"03",X"70",X"04",X"07",X"FB",X"04",X"07",X"98",X"05",X"07",X"ED",X"05",X"07",X"A7",X"06",X"00",
		X"0D",X"96",X"00",X"05",X"C9",X"00",X"05",X"C9",X"00",X"0D",X"D5",X"00",X"0D",X"C9",X"00",X"0D",
		X"8E",X"00",X"05",X"BE",X"00",X"05",X"BE",X"00",X"0D",X"C9",X"00",X"0D",X"BE",X"00",X"0D",X"86",
		X"00",X"05",X"B3",X"00",X"05",X"B3",X"00",X"0D",X"BE",X"00",X"0D",X"B3",X"00",X"0D",X"7F",X"00",
		X"05",X"9F",X"00",X"05",X"9F",X"00",X"0D",X"A9",X"00",X"0D",X"9F",X"00",X"05",X"9F",X"00",X"05",
		X"A9",X"00",X"05",X"9F",X"00",X"05",X"96",X"00",X"05",X"8E",X"00",X"05",X"96",X"00",X"05",X"8E",
		X"00",X"05",X"7F",X"00",X"00",X"23",X"00",X"00",X"0D",X"FD",X"00",X"23",X"00",X"00",X"0D",X"FD",
		X"00",X"23",X"00",X"00",X"0D",X"EF",X"00",X"23",X"00",X"00",X"0D",X"EF",X"00",X"23",X"00",X"00",
		X"0D",X"E1",X"00",X"23",X"00",X"00",X"0D",X"E1",X"00",X"23",X"00",X"00",X"0D",X"D5",X"00",X"23",
		X"00",X"00",X"0D",X"D5",X"00",X"23",X"00",X"00",X"0D",X"B3",X"00",X"23",X"00",X"00",X"0D",X"B3",
		X"00",X"23",X"00",X"00",X"0D",X"B3",X"00",X"23",X"00",X"00",X"0D",X"B3",X"00",X"00",X"0D",X"FB",
		X"04",X"0D",X"3F",X"01",X"0D",X"FB",X"04",X"0D",X"3F",X"01",X"0D",X"B4",X"04",X"0D",X"2D",X"01",
		X"0D",X"B4",X"04",X"0D",X"2D",X"01",X"0D",X"70",X"04",X"0D",X"1C",X"01",X"0D",X"70",X"04",X"0D",
		X"1C",X"01",X"0D",X"31",X"04",X"0D",X"0C",X"01",X"0D",X"31",X"04",X"0D",X"0C",X"01",X"0D",X"FB",
		X"04",X"0D",X"D5",X"00",X"0D",X"FB",X"04",X"0D",X"D5",X"00",X"0D",X"FB",X"04",X"0D",X"98",X"05",
		X"0D",X"ED",X"05",X"0D",X"A7",X"06",X"00",X"05",X"8E",X"00",X"05",X"86",X"00",X"05",X"7F",X"00",
		X"00",X"11",X"9F",X"00",X"01",X"B3",X"00",X"01",X"BE",X"00",X"01",X"D5",X"00",X"07",X"EF",X"00",
		X"00",X"11",X"7F",X"02",X"01",X"CC",X"02",X"01",X"F6",X"02",X"01",X"53",X"03",X"07",X"BC",X"03",
		X"00",X"1F",X"EF",X"00",X"1F",X"EF",X"00",X"00",X"1F",X"1C",X"01",X"1F",X"3F",X"01",X"00",X"1F",
		X"66",X"01",X"1F",X"7B",X"01",X"00",X"1F",X"CC",X"02",X"1F",X"BC",X"03",X"00",X"1F",X"EE",X"00",
		X"1F",X"EE",X"00",X"00",X"2B",X"77",X"00",X"3B",X"00",X"00",X"2B",X"9F",X"00",X"2B",X"9F",X"00",
		X"2B",X"A9",X"00",X"2B",X"9F",X"00",X"00",X"2B",X"8E",X"00",X"39",X"00",X"00",X"2F",X"8E",X"00",
		X"2B",X"7F",X"00",X"39",X"00",X"00",X"2F",X"7F",X"00",X"2B",X"6A",X"00",X"39",X"00",X"00",X"31",
		X"77",X"00",X"2B",X"77",X"00",X"2B",X"77",X"00",X"2B",X"7F",X"00",X"2B",X"8E",X"00",X"00",X"2B",
		X"9F",X"00",X"37",X"00",X"00",X"2B",X"96",X"00",X"2B",X"8E",X"00",X"37",X"00",X"00",X"2B",X"96",
		X"00",X"2D",X"9F",X"00",X"2B",X"9F",X"00",X"2B",X"9F",X"00",X"00",X"2B",X"9F",X"00",X"2B",X"9F",
		X"00",X"00",X"2B",X"A9",X"00",X"2B",X"9F",X"00",X"00",X"2D",X"7F",X"00",X"2B",X"7F",X"00",X"2B",
		X"7F",X"00",X"2B",X"77",X"00",X"2B",X"71",X"00",X"2D",X"6A",X"00",X"2B",X"D5",X"00",X"2B",X"D5",
		X"00",X"2B",X"BE",X"00",X"2B",X"A9",X"00",X"2B",X"9F",X"00",X"37",X"00",X"00",X"2B",X"A9",X"00",
		X"2B",X"9F",X"00",X"37",X"00",X"00",X"2B",X"A9",X"00",X"00",X"2D",X"9F",X"00",X"2B",X"9F",X"00",
		X"2B",X"9F",X"00",X"2B",X"A9",X"00",X"2B",X"9F",X"00",X"00",X"2D",X"9F",X"00",X"2B",X"3F",X"01",
		X"2D",X"3F",X"01",X"2B",X"3F",X"01",X"00",X"2B",X"BE",X"00",X"3D",X"00",X"00",X"00",X"2B",X"3F",
		X"01",X"37",X"00",X"00",X"2B",X"2D",X"01",X"2B",X"1C",X"01",X"37",X"00",X"00",X"2B",X"2D",X"01",
		X"2B",X"3F",X"01",X"37",X"00",X"00",X"2B",X"3F",X"01",X"2B",X"3F",X"01",X"37",X"00",X"00",X"2B",
		X"3F",X"01",X"00",X"2B",X"B3",X"00",X"39",X"00",X"00",X"2F",X"B3",X"00",X"2B",X"B3",X"00",X"39",
		X"00",X"00",X"2F",X"B3",X"00",X"2B",X"BE",X"00",X"39",X"00",X"00",X"31",X"BE",X"00",X"3B",X"00",
		X"00",X"2B",X"B3",X"00",X"37",X"00",X"00",X"2B",X"B3",X"00",X"2B",X"B3",X"00",X"37",X"00",X"00",
		X"2B",X"B3",X"00",X"2D",X"B3",X"00",X"2B",X"B3",X"00",X"2B",X"B3",X"00",X"2B",X"B3",X"00",X"2B",
		X"B3",X"00",X"2B",X"BE",X"00",X"37",X"00",X"00",X"2B",X"BE",X"00",X"2B",X"BE",X"00",X"37",X"00",
		X"00",X"2B",X"BE",X"00",X"2D",X"BE",X"00",X"3B",X"00",X"00",X"2B",X"D5",X"00",X"39",X"00",X"00",
		X"2F",X"D5",X"00",X"2B",X"D5",X"00",X"39",X"00",X"00",X"2F",X"D5",X"00",X"2B",X"9F",X"00",X"39",
		X"00",X"00",X"31",X"9F",X"00",X"2B",X"9F",X"00",X"2B",X"9F",X"00",X"2B",X"9F",X"00",X"2B",X"9F",
		X"00",X"2D",X"9F",X"00",X"2B",X"9F",X"00",X"2B",X"9F",X"00",X"2B",X"9F",X"00",X"2B",X"9F",X"00",
		X"2D",X"A9",X"00",X"2B",X"EF",X"00",X"2B",X"EF",X"00",X"2B",X"EF",X"00",X"2B",X"EF",X"00",X"2B",
		X"FD",X"00",X"37",X"00",X"00",X"2B",X"EF",X"00",X"2B",X"FD",X"00",X"37",X"00",X"00",X"2B",X"EF",
		X"00",X"00",X"2D",X"FD",X"00",X"3B",X"00",X"00",X"00",X"2B",X"BC",X"03",X"3B",X"00",X"00",X"2B",
		X"3F",X"01",X"2B",X"3F",X"01",X"2B",X"52",X"01",X"2B",X"3F",X"01",X"00",X"2B",X"AA",X"01",X"37",
		X"00",X"00",X"2B",X"AA",X"01",X"2B",X"AA",X"01",X"37",X"00",X"00",X"2B",X"AA",X"01",X"00",X"2B",
		X"EF",X"00",X"37",X"00",X"00",X"2B",X"EF",X"00",X"2B",X"EF",X"00",X"37",X"00",X"00",X"2B",X"EF",
		X"00",X"00",X"2B",X"FD",X"00",X"37",X"00",X"00",X"2B",X"FD",X"00",X"2B",X"FD",X"00",X"37",X"00",
		X"00",X"2B",X"FD",X"00",X"2B",X"EF",X"00",X"37",X"00",X"00",X"2B",X"52",X"01",X"2B",X"52",X"01",
		X"37",X"00",X"00",X"2B",X"52",X"01",X"00",X"2D",X"AA",X"01",X"2B",X"3F",X"01",X"2B",X"3F",X"01",
		X"2B",X"52",X"01",X"2B",X"3F",X"01",X"00",X"2D",X"AA",X"01",X"3B",X"00",X"00",X"00",X"2B",X"DE",
		X"01",X"37",X"00",X"00",X"2B",X"DE",X"01",X"2B",X"DE",X"01",X"37",X"00",X"00",X"2B",X"DE",X"01",
		X"00",X"2B",X"DE",X"01",X"37",X"00",X"00",X"2B",X"DE",X"01",X"2B",X"DE",X"01",X"37",X"00",X"00",
		X"2B",X"52",X"01",X"2B",X"3F",X"01",X"37",X"00",X"00",X"2B",X"3F",X"01",X"2B",X"3F",X"01",X"37",
		X"00",X"00",X"2B",X"FD",X"00",X"00",X"2B",X"77",X"07",X"3D",X"00",X"00",X"00",X"2B",X"98",X"05",
		X"37",X"00",X"00",X"2B",X"66",X"01",X"2B",X"98",X"05",X"37",X"00",X"00",X"2B",X"66",X"01",X"2B",
		X"FB",X"04",X"37",X"00",X"00",X"2B",X"66",X"01",X"2B",X"FB",X"04",X"37",X"00",X"00",X"2B",X"66",
		X"01",X"2B",X"BC",X"03",X"39",X"00",X"00",X"31",X"BC",X"03",X"2B",X"7F",X"02",X"2D",X"F6",X"02",
		X"2B",X"BC",X"03",X"00",X"2B",X"F4",X"03",X"37",X"00",X"00",X"2B",X"66",X"01",X"2B",X"FB",X"04",
		X"37",X"00",X"00",X"2B",X"66",X"01",X"00",X"2B",X"BC",X"03",X"37",X"00",X"00",X"2B",X"7B",X"01",
		X"2B",X"FB",X"04",X"37",X"00",X"00",X"2B",X"7B",X"01",X"2B",X"BC",X"03",X"37",X"00",X"00",X"2B",
		X"7B",X"01",X"2F",X"FB",X"04",X"2B",X"47",X"05",X"37",X"00",X"00",X"2B",X"AA",X"01",X"2F",X"47",
		X"05",X"2B",X"98",X"05",X"37",X"00",X"00",X"2B",X"AA",X"01",X"2F",X"98",X"05",X"2B",X"ED",X"05",
		X"37",X"00",X"00",X"2B",X"3F",X"01",X"2F",X"ED",X"05",X"33",X"47",X"06",X"2F",X"A7",X"06",X"2F",
		X"A7",X"06",X"2F",X"A7",X"06",X"2F",X"A7",X"06",X"2D",X"FB",X"04",X"2B",X"A7",X"06",X"2D",X"FB",
		X"04",X"2B",X"A7",X"06",X"00",X"2D",X"FB",X"04",X"3B",X"00",X"00",X"00",X"2F",X"3F",X"01",X"2D",
		X"FD",X"00",X"2B",X"D5",X"00",X"2F",X"8E",X"00",X"2F",X"8E",X"00",X"35",X"8E",X"00",X"2B",X"9F",
		X"00",X"2B",X"9F",X"00",X"2B",X"BE",X"00",X"2B",X"9F",X"00",X"00",X"2B",X"66",X"01",X"37",X"00",
		X"00",X"2B",X"66",X"01",X"2B",X"66",X"01",X"37",X"00",X"00",X"2B",X"66",X"01",X"00",X"2B",X"FA",
		X"01",X"37",X"00",X"00",X"2B",X"FA",X"01",X"2B",X"FA",X"01",X"37",X"00",X"00",X"2B",X"FA",X"01",
		X"00",X"2D",X"F4",X"03",X"37",X"00",X"00",X"2D",X"FB",X"04",X"37",X"00",X"00",X"2D",X"F4",X"03",
		X"2B",X"66",X"01",X"2D",X"FB",X"04",X"2B",X"66",X"01",X"00",X"37",X"00",X"00",X"2B",X"EF",X"00",
		X"2B",X"D5",X"00",X"2B",X"BE",X"00",X"2B",X"B3",X"00",X"2B",X"9F",X"00",X"2D",X"8E",X"00",X"2B",
		X"EF",X"00",X"00",X"2D",X"BC",X"03",X"2B",X"DE",X"01",X"2D",X"FB",X"04",X"2B",X"DE",X"01",X"00",
		X"2D",X"F4",X"03",X"2B",X"3F",X"01",X"2D",X"FB",X"04",X"2B",X"3F",X"01",X"00",X"2F",X"B3",X"00",
		X"2F",X"B3",X"00",X"35",X"BE",X"00",X"2B",X"BE",X"00",X"00",X"35",X"8E",X"00",X"2B",X"B3",X"00",
		X"2B",X"B3",X"00",X"2B",X"D5",X"00",X"2B",X"B3",X"00",X"35",X"8E",X"00",X"2B",X"9F",X"00",X"2D",
		X"BE",X"00",X"2B",X"EF",X"00",X"00",X"2D",X"BE",X"00",X"2B",X"BE",X"00",X"35",X"B3",X"00",X"2B",
		X"B3",X"00",X"2D",X"B3",X"00",X"2B",X"B3",X"00",X"35",X"BE",X"00",X"2B",X"BE",X"00",X"2D",X"EF",
		X"00",X"2B",X"3F",X"01",X"00",X"2D",X"EF",X"00",X"2B",X"EF",X"00",X"2B",X"3F",X"01",X"2B",X"D5",
		X"00",X"2B",X"BE",X"00",X"2B",X"B3",X"00",X"2B",X"9F",X"00",X"2B",X"96",X"00",X"2D",X"8E",X"00",
		X"2B",X"FD",X"00",X"2D",X"FD",X"00",X"2B",X"FD",X"00",X"00",X"2D",X"3F",X"01",X"2B",X"7B",X"01",
		X"00",X"2B",X"BE",X"00",X"2B",X"EF",X"00",X"2B",X"BE",X"00",X"2F",X"A9",X"00",X"2F",X"52",X"01",
		X"2F",X"EF",X"00",X"2F",X"3F",X"01",X"00",X"2F",X"77",X"00",X"2D",X"EF",X"00",X"2B",X"D5",X"00",
		X"2F",X"BE",X"00",X"2F",X"EF",X"00",X"33",X"D5",X"00",X"00",X"2B",X"EF",X"00",X"2B",X"3F",X"01",
		X"2B",X"EF",X"00",X"2F",X"C9",X"00",X"2F",X"92",X"01",X"37",X"00",X"00",X"2B",X"DE",X"01",X"2B",
		X"AA",X"01",X"2B",X"7B",X"01",X"2B",X"66",X"01",X"2B",X"52",X"01",X"2B",X"3F",X"01",X"2B",X"52",
		X"01",X"2B",X"3F",X"01",X"2B",X"2D",X"01",X"2B",X"1C",X"01",X"2B",X"FD",X"00",X"00",X"33",X"B4",
		X"04",X"2F",X"FB",X"04",X"2F",X"FB",X"04",X"2F",X"FB",X"04",X"2F",X"FB",X"04",X"00",X"2D",X"EF",
		X"00",X"2B",X"EF",X"00",X"2B",X"EF",X"00",X"2B",X"FD",X"00",X"2B",X"1C",X"01",X"00",X"2D",X"7B",
		X"01",X"2B",X"DE",X"01",X"2B",X"DE",X"01",X"2B",X"AA",X"01",X"2B",X"7B",X"01",X"00",X"2D",X"EF",
		X"00",X"3B",X"00",X"00",X"00",X"2D",X"BC",X"03",X"3B",X"00",X"00",X"00",X"2D",X"EF",X"00",X"2B",
		X"9F",X"00",X"2B",X"9F",X"00",X"2B",X"8E",X"00",X"2B",X"7F",X"00",X"00",X"2D",X"7B",X"01",X"3B",
		X"00",X"00",X"00",X"2D",X"EF",X"00",X"2B",X"7F",X"02",X"2B",X"CC",X"02",X"2B",X"F6",X"02",X"2B",
		X"53",X"03",X"00",X"2D",X"77",X"00",X"3B",X"00",X"00",X"00",X"57",X"00",X"00",X"00",X"51",X"00",
		X"00",X"41",X"52",X"01",X"45",X"3F",X"01",X"41",X"EF",X"00",X"4D",X"BE",X"00",X"00",X"51",X"00",
		X"00",X"41",X"52",X"01",X"45",X"3F",X"01",X"47",X"EF",X"00",X"41",X"52",X"01",X"45",X"3F",X"01",
		X"47",X"EF",X"00",X"41",X"52",X"01",X"45",X"3F",X"01",X"41",X"D5",X"00",X"4D",X"B3",X"00",X"00",
		X"51",X"00",X"00",X"41",X"2D",X"01",X"45",X"1C",X"01",X"41",X"D5",X"00",X"4D",X"B3",X"00",X"00",
		X"51",X"00",X"00",X"41",X"2D",X"01",X"45",X"1C",X"01",X"47",X"D5",X"00",X"41",X"2D",X"01",X"45",
		X"1C",X"01",X"47",X"C9",X"00",X"41",X"FD",X"00",X"45",X"EF",X"00",X"41",X"BE",X"00",X"4D",X"9F",
		X"00",X"00",X"51",X"00",X"00",X"41",X"C9",X"00",X"45",X"BE",X"00",X"41",X"9F",X"00",X"4D",X"77",
		X"00",X"00",X"51",X"00",X"00",X"41",X"C9",X"00",X"45",X"BE",X"00",X"41",X"9F",X"00",X"45",X"96",
		X"00",X"41",X"BE",X"00",X"45",X"D5",X"00",X"41",X"BE",X"00",X"45",X"B3",X"00",X"41",X"96",X"00",
		X"45",X"8E",X"00",X"41",X"77",X"00",X"45",X"71",X"00",X"41",X"8E",X"00",X"45",X"96",X"00",X"41",
		X"8E",X"00",X"00",X"51",X"00",X"00",X"41",X"1C",X"01",X"45",X"2D",X"01",X"41",X"1C",X"01",X"00",
		X"47",X"EF",X"00",X"45",X"D5",X"00",X"41",X"C9",X"00",X"45",X"BE",X"00",X"41",X"A9",X"00",X"45",
		X"9F",X"00",X"41",X"96",X"00",X"3F",X"8E",X"00",X"3F",X"7F",X"00",X"3F",X"8E",X"00",X"3F",X"7F",
		X"00",X"3F",X"8E",X"00",X"3F",X"7F",X"00",X"45",X"96",X"00",X"41",X"8E",X"00",X"45",X"77",X"00",
		X"41",X"8E",X"00",X"45",X"A9",X"00",X"41",X"C9",X"00",X"45",X"7F",X"00",X"41",X"9F",X"00",X"45",
		X"B3",X"00",X"41",X"D5",X"00",X"45",X"EF",X"00",X"41",X"1C",X"01",X"45",X"3F",X"01",X"41",X"7B",
		X"01",X"45",X"DE",X"01",X"55",X"00",X"00",X"00",X"41",X"77",X"00",X"4F",X"00",X"00",X"00",X"41",
		X"3F",X"01",X"45",X"EF",X"00",X"41",X"FD",X"00",X"00",X"4D",X"7B",X"01",X"00",X"51",X"00",X"00",
		X"41",X"7B",X"01",X"45",X"92",X"01",X"41",X"7B",X"01",X"00",X"45",X"1C",X"01",X"41",X"52",X"01",
		X"47",X"3F",X"01",X"00",X"45",X"1C",X"01",X"41",X"52",X"01",X"45",X"3F",X"01",X"00",X"41",X"EF",
		X"00",X"00",X"41",X"1C",X"01",X"4D",X"FD",X"00",X"51",X"00",X"00",X"00",X"4D",X"66",X"01",X"00",
		X"51",X"00",X"00",X"41",X"66",X"01",X"45",X"7B",X"01",X"41",X"66",X"01",X"45",X"FD",X"00",X"41",
		X"2D",X"01",X"00",X"47",X"1C",X"01",X"00",X"45",X"1C",X"01",X"41",X"52",X"01",X"45",X"3F",X"01",
		X"41",X"7B",X"01",X"45",X"66",X"01",X"41",X"92",X"01",X"4D",X"7B",X"01",X"51",X"00",X"00",X"00",
		X"45",X"3F",X"01",X"41",X"EF",X"00",X"45",X"3F",X"01",X"41",X"EF",X"00",X"45",X"2D",X"01",X"41",
		X"EF",X"00",X"45",X"2D",X"01",X"41",X"EF",X"00",X"4D",X"1C",X"01",X"00",X"4D",X"D5",X"00",X"47",
		X"EF",X"00",X"45",X"FD",X"00",X"41",X"1C",X"01",X"45",X"3F",X"01",X"41",X"52",X"01",X"45",X"3F",
		X"01",X"41",X"FD",X"00",X"45",X"1C",X"01",X"41",X"1C",X"01",X"45",X"2D",X"01",X"41",X"1C",X"01",
		X"45",X"EF",X"00",X"41",X"1C",X"01",X"45",X"EF",X"00",X"41",X"1C",X"01",X"47",X"BE",X"00",X"47",
		X"D5",X"00",X"4D",X"EF",X"00",X"57",X"00",X"00",X"00",X"57",X"00",X"00",X"4D",X"DE",X"01",X"00",
		X"51",X"00",X"00",X"41",X"DE",X"01",X"45",X"FA",X"01",X"41",X"DE",X"01",X"00",X"45",X"66",X"01",
		X"41",X"92",X"01",X"47",X"7B",X"01",X"00",X"45",X"66",X"01",X"41",X"92",X"01",X"45",X"7B",X"01",
		X"00",X"41",X"3F",X"01",X"00",X"41",X"66",X"01",X"4D",X"3F",X"01",X"57",X"00",X"00",X"4D",X"AA",
		X"01",X"00",X"51",X"00",X"00",X"41",X"AA",X"01",X"45",X"C3",X"01",X"41",X"AA",X"01",X"45",X"3F",
		X"01",X"41",X"7B",X"01",X"00",X"47",X"66",X"01",X"00",X"45",X"66",X"01",X"41",X"92",X"01",X"45",
		X"7B",X"01",X"41",X"DE",X"01",X"45",X"AA",X"01",X"41",X"FA",X"01",X"4D",X"DE",X"01",X"00",X"45",
		X"3F",X"01",X"41",X"7B",X"01",X"45",X"3F",X"01",X"41",X"7B",X"01",X"45",X"2D",X"01",X"41",X"7B",
		X"01",X"45",X"2D",X"01",X"41",X"7B",X"01",X"4D",X"66",X"01",X"57",X"00",X"00",X"4D",X"66",X"01",
		X"4D",X"52",X"01",X"45",X"7B",X"01",X"41",X"92",X"01",X"45",X"7B",X"01",X"41",X"AA",X"01",X"45",
		X"C3",X"01",X"41",X"7B",X"01",X"45",X"38",X"02",X"41",X"C3",X"01",X"45",X"AA",X"01",X"41",X"66",
		X"01",X"45",X"92",X"01",X"41",X"52",X"01",X"47",X"3F",X"01",X"47",X"66",X"01",X"4D",X"7B",X"01",
		X"57",X"00",X"00",X"00",X"41",X"77",X"07",X"4F",X"00",X"00",X"55",X"00",X"00",X"00",X"51",X"00",
		X"00",X"41",X"BC",X"03",X"45",X"BC",X"03",X"41",X"BC",X"03",X"4D",X"BC",X"03",X"00",X"51",X"00",
		X"00",X"41",X"BC",X"03",X"51",X"00",X"00",X"41",X"BC",X"03",X"00",X"51",X"00",X"00",X"41",X"FB",
		X"04",X"45",X"FB",X"04",X"41",X"FB",X"04",X"4D",X"FB",X"04",X"00",X"51",X"00",X"00",X"41",X"FB",
		X"04",X"51",X"00",X"00",X"41",X"FB",X"04",X"00",X"47",X"BC",X"03",X"47",X"BC",X"03",X"47",X"86",
		X"03",X"47",X"86",X"03",X"47",X"53",X"03",X"47",X"53",X"03",X"47",X"24",X"03",X"47",X"24",X"03",
		X"4B",X"BC",X"03",X"41",X"F4",X"03",X"4B",X"70",X"04",X"41",X"FB",X"04",X"47",X"98",X"05",X"47",
		X"47",X"05",X"47",X"FB",X"04",X"47",X"FB",X"04",X"4D",X"77",X"07",X"57",X"00",X"00",X"00",X"57",
		X"00",X"00",X"57",X"00",X"00",X"00",X"51",X"00",X"00",X"41",X"3F",X"01",X"45",X"52",X"01",X"41",
		X"66",X"01",X"45",X"7B",X"01",X"00",X"55",X"00",X"00",X"00",X"41",X"AA",X"01",X"45",X"92",X"01",
		X"41",X"7B",X"01",X"45",X"66",X"01",X"00",X"41",X"AA",X"01",X"45",X"7B",X"01",X"41",X"DE",X"01",
		X"45",X"AA",X"01",X"00",X"53",X"00",X"00",X"3F",X"9F",X"00",X"3F",X"A9",X"00",X"45",X"9F",X"00",
		X"00",X"41",X"FA",X"01",X"45",X"DE",X"01",X"41",X"AA",X"01",X"45",X"7B",X"01",X"55",X"00",X"00",
		X"57",X"00",X"00",X"00",X"55",X"00",X"00",X"45",X"52",X"01",X"55",X"00",X"00",X"45",X"3F",X"01",
		X"55",X"00",X"00",X"47",X"3F",X"01",X"41",X"3F",X"01",X"41",X"52",X"01",X"41",X"66",X"01",X"45",
		X"7B",X"01",X"41",X"C3",X"01",X"45",X"DE",X"01",X"41",X"C3",X"01",X"45",X"AA",X"01",X"53",X"00",
		X"00",X"41",X"52",X"01",X"45",X"3F",X"01",X"41",X"3F",X"01",X"45",X"66",X"01",X"41",X"AA",X"01",
		X"47",X"DE",X"01",X"45",X"3F",X"01",X"3F",X"1C",X"01",X"3F",X"FD",X"00",X"41",X"EF",X"00",X"4F",
		X"00",X"00",X"55",X"00",X"00",X"00",X"41",X"77",X"00",X"4F",X"00",X"00",X"55",X"00",X"00",X"57",
		X"00",X"00",X"00",X"51",X"00",X"00",X"41",X"BE",X"00",X"45",X"C9",X"00",X"41",X"D5",X"00",X"45",
		X"EF",X"00",X"00",X"41",X"FD",X"00",X"45",X"EF",X"00",X"41",X"E1",X"00",X"45",X"D5",X"00",X"00",
		X"41",X"FD",X"00",X"45",X"EF",X"00",X"41",X"1C",X"01",X"45",X"FD",X"00",X"00",X"57",X"00",X"00",
		X"00",X"41",X"FD",X"00",X"45",X"1C",X"01",X"41",X"FD",X"00",X"45",X"3F",X"01",X"55",X"00",X"00",
		X"57",X"00",X"00",X"00",X"41",X"3F",X"01",X"45",X"1C",X"01",X"41",X"FD",X"00",X"41",X"EF",X"00",
		X"41",X"FD",X"00",X"41",X"EF",X"00",X"45",X"3F",X"01",X"41",X"7B",X"01",X"45",X"1C",X"01",X"41",
		X"7B",X"01",X"45",X"3F",X"01",X"41",X"1C",X"01",X"45",X"EF",X"00",X"41",X"BE",X"00",X"45",X"C9",
		X"00",X"41",X"D5",X"00",X"45",X"EF",X"00",X"4F",X"00",X"00",X"41",X"EF",X"00",X"41",X"FD",X"00",
		X"41",X"EF",X"00",X"45",X"1C",X"01",X"00",X"47",X"D5",X"00",X"41",X"EF",X"00",X"45",X"FD",X"00",
		X"41",X"FD",X"00",X"45",X"EF",X"00",X"41",X"D5",X"00",X"47",X"BE",X"00",X"00",X"41",X"BE",X"00",
		X"41",X"C9",X"00",X"41",X"D5",X"00",X"45",X"E1",X"00",X"41",X"1C",X"01",X"45",X"2D",X"01",X"41",
		X"3F",X"01",X"45",X"52",X"01",X"00",X"45",X"BE",X"00",X"3F",X"C9",X"00",X"3F",X"D5",X"00",X"43",
		X"EF",X"00",X"3F",X"3F",X"01",X"3F",X"1C",X"01",X"3F",X"FD",X"00",X"41",X"EF",X"00",X"51",X"00",
		X"00",X"00",X"41",X"BC",X"03",X"51",X"00",X"00",X"41",X"FB",X"04",X"51",X"00",X"00",X"41",X"BC",
		X"03",X"51",X"00",X"00",X"41",X"FB",X"04",X"51",X"00",X"00",X"00",X"41",X"FB",X"04",X"51",X"00",
		X"00",X"41",X"A7",X"06",X"51",X"00",X"00",X"41",X"FB",X"04",X"51",X"00",X"00",X"41",X"A7",X"06",
		X"51",X"00",X"00",X"00",X"41",X"BC",X"03",X"51",X"00",X"00",X"41",X"FB",X"04",X"51",X"00",X"00",
		X"41",X"BC",X"03",X"51",X"00",X"00",X"41",X"BC",X"03",X"51",X"00",X"00",X"00",X"41",X"A7",X"06",
		X"51",X"00",X"00",X"41",X"53",X"03",X"51",X"00",X"00",X"41",X"FB",X"04",X"51",X"00",X"00",X"41",
		X"53",X"03",X"51",X"00",X"00",X"00",X"41",X"77",X"07",X"51",X"00",X"00",X"41",X"BC",X"03",X"51",
		X"00",X"00",X"41",X"70",X"04",X"51",X"00",X"00",X"41",X"F6",X"02",X"51",X"00",X"00",X"00",X"5B",
		X"F6",X"02",X"5B",X"24",X"03",X"5B",X"F6",X"02",X"5F",X"7F",X"02",X"5B",X"F6",X"02",X"5F",X"38",
		X"02",X"5B",X"F6",X"02",X"5F",X"7F",X"02",X"5B",X"38",X"02",X"00",X"63",X"DE",X"01",X"51",X"00",
		X"00",X"00",X"5B",X"7F",X"02",X"5F",X"38",X"02",X"5B",X"FA",X"01",X"5F",X"DE",X"01",X"00",X"5B",
		X"7F",X"02",X"5F",X"38",X"02",X"5B",X"18",X"02",X"63",X"FA",X"01",X"00",X"51",X"00",X"00",X"00",
		X"5F",X"DE",X"01",X"5B",X"38",X"02",X"5F",X"7F",X"02",X"5B",X"F6",X"02",X"5F",X"BC",X"03",X"55",
		X"00",X"00",X"00",X"5B",X"F6",X"02",X"5B",X"24",X"03",X"5B",X"F6",X"02",X"5B",X"7F",X"02",X"5B",
		X"A4",X"02",X"5B",X"7F",X"02",X"00",X"5B",X"BC",X"03",X"5B",X"F4",X"03",X"5B",X"BC",X"03",X"00",
		X"5B",X"5A",X"02",X"5B",X"38",X"02",X"5B",X"FA",X"01",X"00",X"5D",X"DE",X"01",X"59",X"7F",X"02",
		X"59",X"38",X"02",X"59",X"FA",X"01",X"5B",X"DE",X"01",X"51",X"00",X"00",X"00",X"51",X"00",X"00",
		X"61",X"AA",X"01",X"5B",X"DE",X"01",X"5F",X"FA",X"01",X"5B",X"7F",X"02",X"5F",X"38",X"02",X"5B",
		X"FA",X"01",X"61",X"DE",X"01",X"00",X"5B",X"DE",X"01",X"5B",X"FA",X"01",X"5B",X"18",X"02",X"5F",
		X"38",X"02",X"5B",X"38",X"02",X"5F",X"5A",X"02",X"5B",X"38",X"02",X"00",X"5F",X"7F",X"02",X"59",
		X"38",X"02",X"59",X"FA",X"01",X"00",X"51",X"00",X"00",X"5B",X"FA",X"01",X"5F",X"DE",X"01",X"5B",
		X"C3",X"01",X"63",X"AA",X"01",X"51",X"00",X"00",X"5B",X"AA",X"01",X"5F",X"7B",X"01",X"5B",X"66",
		X"01",X"5F",X"3F",X"01",X"5B",X"3F",X"01",X"5F",X"1C",X"01",X"5B",X"66",X"01",X"5F",X"3F",X"01",
		X"5B",X"3F",X"01",X"5F",X"66",X"01",X"5B",X"3F",X"01",X"5F",X"7B",X"01",X"5B",X"DE",X"01",X"5F",
		X"38",X"02",X"5B",X"DE",X"01",X"5F",X"7F",X"02",X"5B",X"7F",X"02",X"5F",X"38",X"02",X"5B",X"CC",
		X"02",X"00",X"5F",X"DE",X"01",X"4F",X"00",X"00",X"5F",X"3F",X"01",X"4F",X"00",X"00",X"5F",X"EF",
		X"00",X"59",X"EF",X"00",X"59",X"EF",X"00",X"61",X"EF",X"00",X"00",X"41",X"BC",X"03",X"51",X"00",
		X"00",X"41",X"FB",X"04",X"51",X"00",X"00",X"45",X"BC",X"03",X"3F",X"BC",X"03",X"3F",X"BC",X"03",
		X"47",X"BC",X"03",X"00",X"7D",X"77",X"00",X"7D",X"7F",X"00",X"7D",X"8E",X"00",X"00",X"7B",X"8E",
		X"00",X"79",X"96",X"00",X"00",X"7D",X"9F",X"00",X"7D",X"B3",X"00",X"7D",X"BE",X"00",X"00",X"7D",
		X"D5",X"00",X"7D",X"EF",X"00",X"7D",X"FD",X"00",X"7D",X"1C",X"01",X"00",X"7B",X"1C",X"01",X"79",
		X"2D",X"01",X"00",X"7D",X"3F",X"01",X"7D",X"66",X"01",X"7D",X"7B",X"01",X"00",X"7B",X"7B",X"01",
		X"79",X"92",X"01",X"7D",X"AA",X"01",X"00",X"7D",X"DE",X"01",X"7D",X"FA",X"01",X"7D",X"38",X"02",
		X"00",X"7D",X"7F",X"02",X"7D",X"CC",X"02",X"7D",X"F6",X"02",X"00",X"7B",X"F6",X"02",X"79",X"24",
		X"03",X"00",X"7D",X"53",X"03",X"7D",X"BC",X"03",X"7D",X"F4",X"03",X"7D",X"70",X"04",X"00",X"7D",
		X"FB",X"04",X"7D",X"98",X"05",X"7D",X"ED",X"05",X"00",X"7D",X"A7",X"06",X"00",X"7B",X"38",X"02",
		X"79",X"5A",X"02",X"00",X"7B",X"70",X"04",X"79",X"B4",X"04",X"00",X"7B",X"ED",X"05",X"79",X"47",
		X"06",X"7D",X"6A",X"00",X"00",X"7B",X"BE",X"00",X"79",X"C9",X"00",X"00",X"7D",X"AA",X"01",X"00",
		X"73",X"7B",X"01",X"77",X"EF",X"00",X"73",X"3F",X"01",X"75",X"BE",X"00",X"71",X"EF",X"00",X"75",
		X"D5",X"00",X"71",X"EF",X"00",X"71",X"FD",X"00",X"71",X"EF",X"00",X"71",X"E1",X"00",X"71",X"D5",
		X"00",X"71",X"C9",X"00",X"71",X"BE",X"00",X"71",X"B3",X"00",X"71",X"A9",X"00",X"73",X"9F",X"00",
		X"73",X"9F",X"00",X"73",X"8E",X"00",X"73",X"B3",X"00",X"73",X"BE",X"00",X"77",X"77",X"00",X"73",
		X"9F",X"00",X"75",X"5F",X"00",X"71",X"77",X"00",X"75",X"6A",X"00",X"71",X"77",X"00",X"71",X"7F",
		X"00",X"71",X"77",X"00",X"71",X"71",X"00",X"71",X"6A",X"00",X"71",X"64",X"00",X"71",X"5F",X"00",
		X"71",X"59",X"00",X"71",X"54",X"00",X"71",X"50",X"00",X"71",X"9F",X"00",X"71",X"50",X"00",X"71",
		X"9F",X"00",X"71",X"8E",X"00",X"71",X"9F",X"00",X"71",X"50",X"00",X"71",X"9F",X"00",X"73",X"7F",
		X"00",X"00",X"73",X"9F",X"00",X"73",X"8E",X"00",X"73",X"9F",X"00",X"00",X"73",X"B3",X"00",X"00",
		X"73",X"77",X"00",X"00",X"73",X"BE",X"00",X"00",X"73",X"A9",X"00",X"73",X"8E",X"00",X"73",X"BE",
		X"00",X"73",X"8E",X"00",X"73",X"D5",X"00",X"73",X"8E",X"00",X"73",X"EF",X"00",X"73",X"8E",X"00",
		X"73",X"FD",X"00",X"73",X"D5",X"00",X"73",X"1C",X"01",X"73",X"D5",X"00",X"73",X"3F",X"01",X"73",
		X"3F",X"01",X"73",X"1C",X"01",X"73",X"66",X"01",X"00",X"6B",X"DE",X"01",X"69",X"AA",X"01",X"65",
		X"92",X"01",X"67",X"7B",X"01",X"67",X"DE",X"01",X"00",X"69",X"38",X"02",X"65",X"5A",X"02",X"00",
		X"6D",X"7F",X"02",X"6F",X"00",X"00",X"67",X"7F",X"02",X"67",X"38",X"02",X"00",X"67",X"FA",X"01",
		X"00",X"69",X"CC",X"02",X"65",X"A4",X"02",X"00",X"67",X"18",X"02",X"6B",X"FA",X"01",X"69",X"DE",
		X"01",X"65",X"C3",X"01",X"67",X"AA",X"01",X"67",X"7F",X"02",X"67",X"38",X"02",X"67",X"FA",X"01",
		X"6B",X"DE",X"01",X"69",X"AA",X"01",X"65",X"92",X"01",X"67",X"7B",X"01",X"67",X"DE",X"01",X"67",
		X"AA",X"01",X"67",X"7B",X"01",X"6B",X"52",X"01",X"69",X"3F",X"01",X"65",X"2D",X"01",X"67",X"1C",
		X"01",X"67",X"AA",X"01",X"67",X"7B",X"01",X"67",X"52",X"01",X"65",X"3F",X"01",X"65",X"52",X"01",
		X"67",X"3F",X"01",X"67",X"AA",X"01",X"67",X"FA",X"01",X"67",X"7F",X"02",X"67",X"7F",X"02",X"67",
		X"38",X"02",X"67",X"FA",X"01",X"00",X"85",X"77",X"00",X"8B",X"00",X"00",X"00",X"83",X"66",X"01",
		X"87",X"7B",X"01",X"83",X"66",X"01",X"87",X"7B",X"01",X"85",X"66",X"01",X"85",X"3F",X"01",X"87",
		X"FD",X"00",X"87",X"1C",X"01",X"87",X"3F",X"01",X"87",X"66",X"01",X"00",X"83",X"7B",X"01",X"87",
		X"92",X"01",X"83",X"7B",X"01",X"87",X"92",X"01",X"85",X"7B",X"01",X"00",X"85",X"3F",X"01",X"87",
		X"1C",X"01",X"87",X"3F",X"01",X"87",X"66",X"01",X"87",X"7B",X"01",X"00",X"85",X"EF",X"00",X"81",
		X"1C",X"01",X"85",X"EF",X"00",X"85",X"FD",X"00",X"00",X"85",X"3F",X"01",X"87",X"EF",X"00",X"87",
		X"FD",X"00",X"87",X"1C",X"01",X"87",X"3F",X"01",X"87",X"1C",X"01",X"87",X"2D",X"01",X"85",X"1C",
		X"01",X"85",X"EF",X"00",X"85",X"D5",X"00",X"87",X"BE",X"00",X"87",X"C9",X"00",X"85",X"BE",X"00",
		X"85",X"B3",X"00",X"85",X"BE",X"00",X"87",X"BE",X"00",X"87",X"D5",X"00",X"87",X"EF",X"00",X"87",
		X"1C",X"01",X"85",X"BE",X"00",X"85",X"D5",X"00",X"00",X"85",X"EF",X"00",X"8B",X"00",X"00",X"00",
		X"89",X"00",X"00",X"00",X"83",X"FA",X"01",X"87",X"18",X"02",X"83",X"FA",X"01",X"87",X"18",X"02",
		X"85",X"FA",X"01",X"8B",X"00",X"00",X"83",X"DE",X"01",X"87",X"FA",X"01",X"83",X"DE",X"01",X"87",
		X"FA",X"01",X"85",X"DE",X"01",X"8B",X"00",X"00",X"00",X"83",X"AA",X"01",X"87",X"C3",X"01",X"83",
		X"AA",X"01",X"87",X"C3",X"01",X"85",X"AA",X"01",X"8B",X"00",X"00",X"85",X"7B",X"01",X"81",X"92",
		X"01",X"85",X"7B",X"01",X"85",X"66",X"01",X"8B",X"00",X"00",X"00",X"87",X"66",X"01",X"87",X"7B",
		X"01",X"85",X"66",X"01",X"81",X"2D",X"01",X"87",X"3F",X"01",X"87",X"52",X"01",X"85",X"3F",X"01",
		X"85",X"1C",X"01",X"85",X"3F",X"01",X"81",X"52",X"01",X"85",X"3F",X"01",X"85",X"66",X"01",X"00",
		X"85",X"7B",X"01",X"8B",X"00",X"00",X"00",X"85",X"BC",X"03",X"00",X"85",X"FB",X"04",X"85",X"70",
		X"04",X"85",X"31",X"04",X"85",X"F4",X"03",X"8D",X"00",X"00",X"85",X"FB",X"04",X"8D",X"00",X"00",
		X"85",X"F4",X"03",X"85",X"FB",X"04",X"85",X"70",X"04",X"85",X"F4",X"03",X"85",X"BC",X"03",X"8D",
		X"00",X"00",X"85",X"FB",X"04",X"8D",X"00",X"00",X"85",X"BC",X"03",X"00",X"85",X"F6",X"02",X"85",
		X"CC",X"02",X"85",X"A4",X"02",X"85",X"7F",X"02",X"8D",X"00",X"00",X"85",X"53",X"03",X"8D",X"00",
		X"00",X"85",X"7F",X"02",X"85",X"7F",X"02",X"85",X"38",X"02",X"85",X"FA",X"01",X"85",X"DE",X"01",
		X"85",X"38",X"02",X"85",X"7F",X"02",X"85",X"F6",X"02",X"85",X"53",X"03",X"00",X"85",X"BC",X"03",
		X"85",X"53",X"03",X"85",X"F6",X"02",X"85",X"CC",X"02",X"87",X"F6",X"02",X"87",X"24",X"03",X"85",
		X"53",X"03",X"85",X"CC",X"02",X"85",X"BC",X"03",X"87",X"F4",X"03",X"87",X"31",X"04",X"85",X"70",
		X"04",X"85",X"86",X"03",X"85",X"53",X"03",X"85",X"A4",X"02",X"85",X"7F",X"02",X"85",X"FA",X"01",
		X"00",X"85",X"DE",X"01",X"00",X"7F",X"B3",X"00",X"87",X"B3",X"00",X"87",X"9F",X"00",X"87",X"B3",
		X"00",X"87",X"9F",X"00",X"87",X"B3",X"00",X"87",X"9F",X"00",X"87",X"B3",X"00",X"87",X"9F",X"00",
		X"7F",X"BE",X"00",X"87",X"BE",X"00",X"87",X"9F",X"00",X"87",X"BE",X"00",X"87",X"9F",X"00",X"87",
		X"BE",X"00",X"87",X"9F",X"00",X"87",X"BE",X"00",X"87",X"9F",X"00",X"00",X"7F",X"D5",X"00",X"87",
		X"D5",X"00",X"87",X"7F",X"00",X"87",X"D5",X"00",X"87",X"7F",X"00",X"87",X"D5",X"00",X"87",X"7F",
		X"00",X"87",X"D5",X"00",X"87",X"7F",X"00",X"87",X"BE",X"00",X"87",X"77",X"00",X"87",X"C9",X"00",
		X"87",X"8E",X"00",X"87",X"C9",X"00",X"87",X"8E",X"00",X"87",X"BE",X"00",X"87",X"77",X"00",X"7F",
		X"B3",X"00",X"00",X"81",X"8E",X"00",X"87",X"96",X"00",X"87",X"77",X"00",X"87",X"96",X"00",X"87",
		X"6A",X"00",X"81",X"9F",X"00",X"87",X"8E",X"00",X"87",X"59",X"00",X"87",X"9F",X"00",X"87",X"5F",
		X"00",X"81",X"A9",X"00",X"87",X"9F",X"00",X"87",X"5F",X"00",X"87",X"B3",X"00",X"87",X"6A",X"00",
		X"00",X"85",X"BE",X"00",X"8B",X"00",X"00",X"00",X"41",X"77",X"00",X"51",X"00",X"00",X"00",X"41",
		X"3F",X"01",X"41",X"1C",X"01",X"41",X"FD",X"00",X"41",X"EF",X"00",X"41",X"FD",X"00",X"41",X"EF",
		X"00",X"45",X"3F",X"01",X"41",X"7B",X"01",X"41",X"1C",X"01",X"41",X"3F",X"01",X"41",X"1C",X"01",
		X"45",X"66",X"01",X"41",X"AA",X"01",X"45",X"3F",X"01",X"41",X"3F",X"01",X"00",X"45",X"52",X"01",
		X"41",X"52",X"01",X"47",X"66",X"01",X"00",X"45",X"3F",X"01",X"41",X"3F",X"01",X"47",X"3F",X"01",
		X"41",X"7B",X"01",X"41",X"66",X"01",X"41",X"3F",X"01",X"41",X"1C",X"01",X"41",X"2D",X"01",X"41",
		X"1C",X"01",X"45",X"EF",X"00",X"41",X"E1",X"00",X"41",X"D5",X"00",X"41",X"D5",X"00",X"55",X"00",
		X"00",X"41",X"D5",X"00",X"41",X"EF",X"00",X"41",X"D5",X"00",X"45",X"FD",X"00",X"41",X"D5",X"00",
		X"41",X"BE",X"00",X"41",X"BE",X"00",X"55",X"00",X"00",X"41",X"BE",X"00",X"41",X"D5",X"00",X"41",
		X"BE",X"00",X"45",X"E1",X"00",X"41",X"BE",X"00",X"41",X"B3",X"00",X"41",X"BE",X"00",X"41",X"B3",
		X"00",X"41",X"D5",X"00",X"41",X"BE",X"00",X"41",X"A9",X"00",X"45",X"9F",X"00",X"41",X"9F",X"00",
		X"45",X"9F",X"00",X"41",X"9F",X"00",X"47",X"9F",X"00",X"00",X"53",X"00",X"00",X"00",X"41",X"FA",
		X"01",X"41",X"DE",X"01",X"41",X"AA",X"01",X"47",X"7B",X"01",X"47",X"DE",X"01",X"47",X"AA",X"01",
		X"47",X"FA",X"01",X"00",X"45",X"7B",X"01",X"41",X"7B",X"01",X"45",X"92",X"01",X"41",X"92",X"01",
		X"47",X"AA",X"01",X"00",X"47",X"DE",X"01",X"47",X"FA",X"01",X"47",X"18",X"02",X"41",X"DE",X"01",
		X"41",X"AA",X"01",X"41",X"7B",X"01",X"47",X"66",X"01",X"47",X"1C",X"01",X"41",X"2D",X"01",X"41",
		X"3F",X"01",X"41",X"2D",X"01",X"45",X"66",X"01",X"41",X"2D",X"01",X"41",X"FD",X"00",X"41",X"1C",
		X"01",X"41",X"FD",X"00",X"45",X"2D",X"01",X"41",X"FD",X"00",X"41",X"EF",X"00",X"41",X"FD",X"00",
		X"41",X"EF",X"00",X"45",X"1C",X"01",X"41",X"EF",X"00",X"41",X"E1",X"00",X"41",X"FD",X"00",X"41",
		X"E1",X"00",X"45",X"1C",X"01",X"41",X"E1",X"00",X"41",X"D5",X"00",X"41",X"E1",X"00",X"41",X"D5",
		X"00",X"41",X"52",X"01",X"41",X"3F",X"01",X"41",X"1C",X"01",X"45",X"FD",X"00",X"41",X"FD",X"00",
		X"45",X"EF",X"00",X"41",X"EF",X"00",X"47",X"D5",X"00",X"00",X"57",X"00",X"00",X"00",X"57",X"00",
		X"00",X"57",X"00",X"00",X"00",X"45",X"7B",X"01",X"41",X"7B",X"01",X"45",X"7B",X"01",X"41",X"7B",
		X"01",X"47",X"7B",X"01",X"53",X"00",X"00",X"00",X"45",X"5A",X"02",X"41",X"38",X"02",X"45",X"FA",
		X"01",X"41",X"AA",X"01",X"45",X"38",X"02",X"41",X"FA",X"01",X"45",X"DE",X"01",X"41",X"7B",X"01",
		X"45",X"C3",X"01",X"41",X"AA",X"01",X"45",X"7B",X"01",X"41",X"3F",X"01",X"45",X"AA",X"01",X"41",
		X"7B",X"01",X"45",X"DE",X"01",X"41",X"AA",X"01",X"45",X"AA",X"01",X"41",X"AA",X"01",X"45",X"7B",
		X"01",X"41",X"7B",X"01",X"47",X"66",X"01",X"00",X"41",X"77",X"07",X"51",X"00",X"00",X"00",X"45",
		X"BC",X"03",X"4F",X"00",X"00",X"45",X"7F",X"02",X"4F",X"00",X"00",X"45",X"53",X"03",X"4F",X"00",
		X"00",X"45",X"7F",X"02",X"4F",X"00",X"00",X"00",X"45",X"BC",X"03",X"4F",X"00",X"00",X"45",X"24",
		X"03",X"4F",X"00",X"00",X"45",X"53",X"03",X"4F",X"00",X"00",X"45",X"FB",X"04",X"4F",X"00",X"00",
		X"00",X"45",X"F6",X"02",X"4F",X"00",X"00",X"45",X"7F",X"02",X"4F",X"00",X"00",X"45",X"18",X"02",
		X"41",X"DE",X"01",X"45",X"38",X"02",X"41",X"7F",X"02",X"45",X"CC",X"02",X"4F",X"00",X"00",X"45",
		X"38",X"02",X"4F",X"00",X"00",X"45",X"5A",X"02",X"4F",X"00",X"00",X"45",X"FA",X"01",X"4F",X"00",
		X"00",X"45",X"F6",X"02",X"4F",X"00",X"00",X"45",X"5A",X"02",X"4F",X"00",X"00",X"45",X"38",X"02",
		X"4F",X"00",X"00",X"45",X"DE",X"01",X"4F",X"00",X"00",X"45",X"38",X"02",X"4F",X"00",X"00",X"45",
		X"C3",X"01",X"4F",X"00",X"00",X"45",X"AA",X"01",X"4F",X"00",X"00",X"45",X"38",X"02",X"4F",X"00",
		X"00",X"47",X"7F",X"02",X"47",X"38",X"02",X"47",X"FA",X"01",X"00",X"05",X"05",X"01",X"01",X"01",
		X"02",X"FC",X"00",X"06",X"05",X"01",X"01",X"01",X"02",X"FC",X"00",X"06",X"04",X"02",X"01",X"01",
		X"02",X"00",X"04",X"01",X"FF",X"00",X"03",X"08",X"01",X"01",X"01",X"04",X"00",X"02",X"01",X"FC",
		X"00",X"02",X"08",X"01",X"01",X"01",X"0B",X"00",X"02",X"01",X"FC",X"00",X"03",X"08",X"01",X"01",
		X"01",X"0B",X"00",X"02",X"01",X"FC",X"00",X"02",X"08",X"01",X"01",X"01",X"12",X"00",X"02",X"01",
		X"FC",X"00",X"03",X"08",X"01",X"01",X"01",X"12",X"00",X"02",X"01",X"FC",X"00",X"02",X"08",X"01",
		X"01",X"01",X"20",X"00",X"02",X"01",X"FC",X"00",X"02",X"08",X"01",X"01",X"01",X"2E",X"00",X"02",
		X"01",X"FC",X"00",X"03",X"08",X"01",X"01",X"01",X"2E",X"00",X"02",X"01",X"FC",X"00",X"02",X"08",
		X"01",X"01",X"01",X"4A",X"00",X"02",X"01",X"FC",X"00",X"03",X"08",X"01",X"01",X"01",X"4A",X"00",
		X"02",X"01",X"FC",X"00",X"02",X"08",X"01",X"01",X"01",X"66",X"00",X"02",X"01",X"FC",X"00",X"02",
		X"08",X"01",X"01",X"01",X"D6",X"00",X"02",X"01",X"FC",X"00",X"04",X"02",X"01",X"03",X"01",X"DC",
		X"00",X"02",X"01",X"FC",X"00",X"00",X"01",X"0E",X"00",X"00",X"00",X"01",X"1C",X"00",X"00",X"00",
		X"01",X"38",X"00",X"00",X"00",X"01",X"54",X"00",X"00",X"00",X"01",X"70",X"00",X"00",X"02",X"08",
		X"01",X"01",X"01",X"0A",X"00",X"02",X"01",X"FC",X"00",X"02",X"08",X"01",X"01",X"01",X"1E",X"00",
		X"02",X"01",X"FC",X"00",X"02",X"08",X"01",X"01",X"01",X"32",X"00",X"02",X"01",X"FC",X"00",X"02",
		X"08",X"01",X"01",X"01",X"5A",X"00",X"02",X"01",X"FC",X"00",X"02",X"08",X"01",X"01",X"01",X"6E",
		X"00",X"02",X"01",X"FC",X"00",X"02",X"08",X"01",X"01",X"01",X"96",X"00",X"02",X"01",X"FC",X"00",
		X"00",X"01",X"14",X"00",X"00",X"00",X"01",X"28",X"00",X"00",X"00",X"01",X"50",X"00",X"00",X"00",
		X"01",X"A0",X"00",X"00",X"01",X"03",X"01",X"03",X"01",X"46",X"00",X"07",X"01",X"FF",X"00",X"00",
		X"01",X"30",X"00",X"00",X"02",X"03",X"01",X"03",X"01",X"26",X"00",X"07",X"01",X"FF",X"00",X"06",
		X"05",X"01",X"01",X"01",X"06",X"00",X"02",X"01",X"FD",X"00",X"03",X"08",X"01",X"01",X"01",X"10",
		X"00",X"02",X"01",X"FC",X"00",X"03",X"08",X"01",X"01",X"01",X"1D",X"00",X"02",X"01",X"FC",X"00",
		X"03",X"08",X"01",X"01",X"01",X"2A",X"00",X"02",X"01",X"FC",X"00",X"03",X"08",X"01",X"01",X"01",
		X"5E",X"00",X"02",X"01",X"FC",X"00",X"00",X"01",X"1A",X"00",X"00",X"05",X"05",X"01",X"01",X"01",
		X"06",X"00",X"02",X"01",X"FD",X"00",X"02",X"08",X"01",X"01",X"01",X"1D",X"00",X"02",X"01",X"FC",
		X"00",X"02",X"08",X"01",X"01",X"01",X"2A",X"00",X"02",X"01",X"FC",X"00",X"07",X"03",X"01",X"01",
		X"01",X"02",X"00",X"03",X"01",X"FF",X"00",X"08",X"03",X"01",X"01",X"01",X"02",X"00",X"03",X"01",
		X"FF",X"00",X"07",X"03",X"01",X"01",X"01",X"06",X"00",X"07",X"01",X"FF",X"00",X"08",X"03",X"01",
		X"01",X"01",X"06",X"00",X"07",X"01",X"FF",X"00",X"01",X"03",X"01",X"03",X"01",X"0E",X"00",X"07",
		X"01",X"FF",X"00",X"02",X"03",X"01",X"03",X"01",X"0E",X"00",X"07",X"01",X"FF",X"00",X"01",X"03",
		X"01",X"03",X"01",X"16",X"00",X"07",X"01",X"FF",X"00",X"02",X"03",X"01",X"03",X"01",X"16",X"00",
		X"07",X"01",X"FF",X"00",X"01",X"03",X"01",X"03",X"01",X"26",X"00",X"07",X"01",X"FF",X"00",X"01",
		X"03",X"01",X"03",X"01",X"36",X"00",X"07",X"01",X"FF",X"00",X"02",X"03",X"01",X"03",X"01",X"36",
		X"00",X"07",X"01",X"FF",X"00",X"01",X"03",X"01",X"03",X"01",X"56",X"00",X"07",X"01",X"FF",X"00",
		X"02",X"03",X"01",X"03",X"01",X"56",X"00",X"07",X"01",X"FF",X"00",X"00",X"01",X"10",X"00",X"00",
		X"00",X"01",X"20",X"00",X"00",X"00",X"01",X"40",X"00",X"00",X"00",X"01",X"60",X"00",X"00",X"00",
		X"00",X"00",X"00",X"45",X"61",X"72",X"6C",X"43",X"6F",X"72",X"62",X"61",X"6E",X"56",X"69",X"63",
		X"6B",X"65",X"72",X"73",X"06",X"06",X"11",X"09",X"00",X"DD",X"21",X"BC",X"82",X"DD",X"7E",X"01",
		X"FE",X"FF",X"28",X"13",X"DD",X"4E",X"02",X"21",X"F0",X"34",X"E5",X"DD",X"6E",X"00",X"67",X"E9",
		X"11",X"09",X"00",X"DD",X"36",X"02",X"00",X"DD",X"19",X"10",X"E2",X"C9",X"FD",X"E1",X"C5",X"3E",
		X"06",X"90",X"4F",X"FD",X"5E",X"02",X"CD",X"65",X"3B",X"C1",X"C5",X"E5",X"DD",X"E3",X"79",X"FE",
		X"00",X"28",X"33",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"DD",X"5E",X"02",X"DD",X"56",X"03",X"7E",
		X"12",X"FD",X"CB",X"03",X"4E",X"28",X"04",X"23",X"13",X"7E",X"12",X"FD",X"7E",X"06",X"DD",X"77",
		X"04",X"FD",X"7E",X"05",X"DD",X"77",X"05",X"AF",X"DD",X"77",X"06",X"FD",X"7E",X"04",X"DD",X"77",
		X"07",X"DD",X"E1",X"C3",X"04",X"36",X"DD",X"35",X"04",X"28",X"05",X"DD",X"E1",X"C3",X"04",X"36",
		X"FD",X"46",X"03",X"CB",X"48",X"26",X"00",X"DD",X"6E",X"06",X"54",X"5D",X"20",X"04",X"0E",X"03",
		X"18",X"03",X"0E",X"04",X"29",X"19",X"19",X"16",X"00",X"1E",X"05",X"19",X"EB",X"FD",X"E5",X"FD",
		X"19",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"DD",X"5E",X"02",X"DD",X"56",X"03",X"CB",X"48",X"20",
		X"07",X"FD",X"7E",X"02",X"86",X"12",X"18",X"10",X"C5",X"4E",X"23",X"46",X"FD",X"6E",X"02",X"FD",
		X"66",X"03",X"09",X"C1",X"EB",X"73",X"23",X"72",X"DD",X"35",X"05",X"20",X"5D",X"DD",X"34",X"06",
		X"16",X"00",X"59",X"FD",X"19",X"FD",X"7E",X"00",X"FE",X"00",X"20",X"3C",X"DD",X"7E",X"07",X"FE",
		X"00",X"28",X"1D",X"FE",X"FF",X"28",X"03",X"DD",X"35",X"07",X"AF",X"DD",X"77",X"06",X"FD",X"E1",
		X"FD",X"7E",X"05",X"DD",X"77",X"05",X"FD",X"7E",X"06",X"DD",X"77",X"04",X"DD",X"E1",X"18",X"34",
		X"FD",X"E1",X"DD",X"E1",X"C1",X"3E",X"06",X"90",X"21",X"E0",X"3C",X"16",X"00",X"5F",X"19",X"3A",
		X"1F",X"83",X"B6",X"32",X"1F",X"83",X"18",X"1D",X"FD",X"7E",X"01",X"DD",X"77",X"04",X"FD",X"7E",
		X"00",X"DD",X"77",X"05",X"FD",X"E1",X"DD",X"E1",X"18",X"0A",X"FD",X"7E",X"01",X"DD",X"77",X"04",
		X"FD",X"E1",X"DD",X"E1",X"C1",X"FD",X"6E",X"00",X"FD",X"66",X"01",X"E5",X"C9",X"FD",X"E1",X"C5",
		X"3E",X"06",X"90",X"4F",X"FD",X"5E",X"02",X"CD",X"65",X"3B",X"C1",X"E5",X"DD",X"E3",X"79",X"FE",
		X"00",X"28",X"2A",X"FD",X"7E",X"06",X"DD",X"5E",X"02",X"DD",X"56",X"03",X"12",X"FD",X"CB",X"03",
		X"4E",X"28",X"05",X"13",X"FD",X"7E",X"07",X"12",X"FD",X"7E",X"05",X"DD",X"77",X"04",X"AF",X"DD",
		X"77",X"06",X"FD",X"7E",X"04",X"DD",X"77",X"07",X"DD",X"E1",X"C3",X"E1",X"36",X"DD",X"35",X"04",
		X"28",X"05",X"DD",X"E1",X"C3",X"E1",X"36",X"DD",X"34",X"06",X"C5",X"FD",X"46",X"03",X"CB",X"48",
		X"26",X"00",X"DD",X"6E",X"06",X"54",X"5D",X"29",X"28",X"01",X"19",X"FD",X"E5",X"16",X"00",X"1E",
		X"05",X"19",X"EB",X"FD",X"19",X"FD",X"7E",X"00",X"FE",X"00",X"28",X"1D",X"DD",X"77",X"04",X"FD",
		X"7E",X"01",X"DD",X"5E",X"02",X"DD",X"56",X"03",X"12",X"CB",X"48",X"28",X"05",X"FD",X"7E",X"02",
		X"13",X"12",X"FD",X"E1",X"C1",X"DD",X"E1",X"18",X"48",X"DD",X"7E",X"07",X"FE",X"00",X"28",X"2B",
		X"FE",X"FF",X"28",X"03",X"DD",X"35",X"07",X"AF",X"DD",X"77",X"06",X"FD",X"E1",X"FD",X"7E",X"05",
		X"DD",X"77",X"04",X"FD",X"7E",X"06",X"DD",X"5E",X"02",X"DD",X"56",X"03",X"12",X"CB",X"48",X"28",
		X"05",X"FD",X"7E",X"07",X"13",X"12",X"C1",X"DD",X"E1",X"18",X"16",X"FD",X"E1",X"C1",X"DD",X"E1",
		X"3E",X"06",X"90",X"21",X"E0",X"3C",X"16",X"00",X"5F",X"19",X"3A",X"1F",X"83",X"B6",X"32",X"1F",
		X"83",X"FD",X"6E",X"00",X"FD",X"66",X"01",X"E5",X"C9",X"FD",X"E1",X"C5",X"3E",X"06",X"90",X"4F",
		X"FD",X"5E",X"02",X"CD",X"65",X"3B",X"C1",X"E5",X"DD",X"E3",X"79",X"FE",X"00",X"28",X"0C",X"FD",
		X"7E",X"03",X"DD",X"77",X"00",X"CD",X"C8",X"37",X"C3",X"BE",X"37",X"DD",X"35",X"0C",X"C2",X"BE",
		X"37",X"DD",X"5E",X"09",X"DD",X"56",X"0A",X"21",X"02",X"00",X"19",X"7E",X"DD",X"6E",X"0F",X"DD",
		X"66",X"10",X"86",X"77",X"DD",X"35",X"0B",X"C2",X"B6",X"37",X"21",X"03",X"00",X"19",X"DD",X"75",
		X"09",X"DD",X"74",X"0A",X"7E",X"FE",X"00",X"20",X"70",X"DD",X"5E",X"05",X"DD",X"56",X"06",X"21",
		X"03",X"00",X"19",X"DD",X"75",X"05",X"DD",X"74",X"06",X"7E",X"FE",X"00",X"20",X"54",X"DD",X"6E",
		X"01",X"DD",X"66",X"02",X"23",X"23",X"DD",X"75",X"01",X"DD",X"74",X"02",X"23",X"7E",X"FE",X"00",
		X"20",X"26",X"DD",X"7E",X"00",X"FE",X"00",X"20",X"13",X"3E",X"06",X"90",X"21",X"E0",X"3C",X"16",
		X"00",X"5F",X"19",X"3A",X"1F",X"83",X"B6",X"32",X"1F",X"83",X"18",X"42",X"FE",X"FF",X"28",X"03",
		X"DD",X"35",X"00",X"CD",X"C8",X"37",X"18",X"36",X"DD",X"6E",X"01",X"DD",X"66",X"02",X"5E",X"23",
		X"56",X"DD",X"73",X"03",X"DD",X"72",X"04",X"DD",X"73",X"05",X"DD",X"72",X"06",X"CD",X"2B",X"38",
		X"18",X"1C",X"54",X"5D",X"CD",X"2B",X"38",X"18",X"15",X"DD",X"77",X"0B",X"11",X"01",X"00",X"19",
		X"7E",X"DD",X"77",X"0C",X"18",X"08",X"21",X"01",X"00",X"19",X"7E",X"DD",X"77",X"0C",X"DD",X"E1",
		X"FD",X"6E",X"00",X"FD",X"66",X"01",X"E5",X"C9",X"FD",X"E5",X"E1",X"11",X"04",X"00",X"19",X"DD",
		X"75",X"01",X"DD",X"74",X"02",X"FD",X"7E",X"04",X"DD",X"77",X"03",X"DD",X"77",X"05",X"6F",X"FD",
		X"7E",X"05",X"DD",X"77",X"04",X"DD",X"77",X"06",X"67",X"23",X"DD",X"5E",X"0D",X"DD",X"56",X"0E",
		X"7E",X"12",X"23",X"13",X"7E",X"12",X"2B",X"2B",X"16",X"00",X"5E",X"21",X"00",X"08",X"19",X"5E",
		X"DD",X"73",X"07",X"23",X"56",X"DD",X"72",X"08",X"21",X"00",X"00",X"19",X"7E",X"DD",X"6E",X"0F",
		X"DD",X"66",X"10",X"77",X"21",X"01",X"00",X"19",X"DD",X"75",X"09",X"DD",X"74",X"0A",X"7E",X"DD",
		X"77",X"0B",X"11",X"01",X"00",X"19",X"7E",X"DD",X"77",X"0C",X"C9",X"13",X"DD",X"6E",X"0D",X"DD",
		X"66",X"0E",X"1A",X"77",X"13",X"23",X"1A",X"77",X"1B",X"1B",X"26",X"00",X"1A",X"6F",X"11",X"00",
		X"08",X"19",X"5E",X"23",X"56",X"DD",X"73",X"07",X"DD",X"72",X"08",X"21",X"00",X"00",X"19",X"7E",
		X"DD",X"6E",X"0F",X"DD",X"66",X"10",X"77",X"21",X"01",X"00",X"19",X"DD",X"75",X"09",X"DD",X"74",
		X"0A",X"7E",X"DD",X"77",X"0B",X"11",X"01",X"00",X"19",X"7E",X"DD",X"77",X"0C",X"C9",X"3E",X"06",
		X"90",X"6F",X"26",X"00",X"29",X"54",X"5D",X"29",X"29",X"19",X"11",X"44",X"82",X"19",X"FD",X"E1",
		X"E5",X"26",X"00",X"FD",X"6E",X"02",X"54",X"5D",X"29",X"29",X"19",X"DD",X"E3",X"EB",X"DD",X"19",
		X"DD",X"7E",X"04",X"FE",X"00",X"28",X"05",X"DD",X"35",X"04",X"18",X"35",X"3A",X"71",X"83",X"C5",
		X"4F",X"E6",X"33",X"EA",X"A7",X"38",X"37",X"79",X"1F",X"32",X"71",X"83",X"47",X"FD",X"7E",X"03",
		X"DD",X"77",X"04",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"5E",X"16",X"00",X"21",X"D7",X"3C",X"19",
		X"4E",X"79",X"A0",X"47",X"79",X"2F",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"4E",X"A1",X"B0",X"77",
		X"C1",X"DD",X"E1",X"FD",X"6E",X"00",X"FD",X"66",X"01",X"E5",X"C9",X"C5",X"3E",X"06",X"90",X"47",
		X"57",X"1E",X"2E",X"CD",X"56",X"3B",X"EB",X"FD",X"21",X"83",X"3B",X"FD",X"19",X"16",X"00",X"58",
		X"21",X"3E",X"82",X"19",X"FD",X"7E",X"14",X"4F",X"FE",X"0F",X"7E",X"20",X"17",X"CB",X"27",X"CB",
		X"27",X"CB",X"27",X"CB",X"27",X"E6",X"F0",X"47",X"FD",X"6E",X"12",X"FD",X"66",X"13",X"7E",X"A1",
		X"B0",X"77",X"C1",X"C9",X"E6",X"0F",X"18",X"EF",X"01",X"1F",X"00",X"21",X"00",X"80",X"11",X"20",
		X"80",X"09",X"EB",X"09",X"06",X"0F",X"DD",X"21",X"00",X"B0",X"1A",X"BE",X"28",X"07",X"77",X"DD",
		X"70",X"00",X"32",X"02",X"B0",X"1B",X"2B",X"05",X"F2",X"2A",X"39",X"06",X"0F",X"DD",X"21",X"00",
		X"A0",X"1A",X"BE",X"28",X"07",X"77",X"DD",X"70",X"00",X"32",X"02",X"A0",X"1B",X"2B",X"05",X"F2",
		X"41",X"39",X"C9",X"DD",X"21",X"BC",X"82",X"06",X"00",X"DD",X"7E",X"04",X"DD",X"BE",X"03",X"28",
		X"49",X"DD",X"77",X"03",X"DD",X"36",X"02",X"01",X"26",X"00",X"DD",X"6E",X"04",X"29",X"54",X"5D",
		X"19",X"19",X"11",X"7E",X"0A",X"19",X"5E",X"23",X"56",X"DD",X"E5",X"E5",X"EB",X"11",X"82",X"39",
		X"D5",X"E9",X"E1",X"DD",X"E1",X"23",X"7E",X"DD",X"77",X"00",X"23",X"7E",X"DD",X"77",X"01",X"DD",
		X"7E",X"04",X"FE",X"00",X"28",X"14",X"23",X"23",X"7E",X"FE",X"FF",X"28",X"0D",X"DD",X"E5",X"57",
		X"2B",X"5E",X"EB",X"11",X"A8",X"39",X"D5",X"E9",X"DD",X"E1",X"11",X"09",X"00",X"DD",X"19",X"04",
		X"78",X"FE",X"06",X"20",X"A4",X"C9",X"50",X"1E",X"2E",X"CD",X"56",X"3B",X"11",X"83",X"3B",X"19",
		X"E5",X"FD",X"E1",X"DD",X"E3",X"DD",X"CB",X"00",X"46",X"20",X"10",X"FD",X"7E",X"09",X"2F",X"4F",
		X"FD",X"5E",X"06",X"FD",X"56",X"07",X"1A",X"B1",X"12",X"18",X"0B",X"FD",X"5E",X"06",X"FD",X"56",
		X"07",X"1A",X"FD",X"A6",X"09",X"12",X"DD",X"CB",X"00",X"66",X"20",X"0A",X"FD",X"7E",X"08",X"2F",
		X"4F",X"1A",X"B1",X"12",X"18",X"05",X"1A",X"FD",X"A6",X"08",X"12",X"DD",X"4E",X"01",X"FD",X"7E",
		X"14",X"FE",X"0F",X"20",X"0A",X"79",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"4F",X"FD",
		X"5E",X"12",X"FD",X"56",X"13",X"1A",X"FD",X"A6",X"14",X"B1",X"12",X"DD",X"7E",X"02",X"4F",X"FE",
		X"FF",X"28",X"2F",X"26",X"00",X"68",X"5D",X"54",X"29",X"29",X"29",X"19",X"11",X"BC",X"82",X"19",
		X"11",X"01",X"90",X"3E",X"06",X"CD",X"51",X"3B",X"1A",X"E6",X"7F",X"77",X"23",X"FD",X"E5",X"D1",
		X"EB",X"79",X"CD",X"51",X"3B",X"7E",X"12",X"23",X"13",X"66",X"6F",X"EB",X"72",X"21",X"03",X"90",
		X"7E",X"12",X"DD",X"E5",X"E1",X"1E",X"03",X"16",X"00",X"19",X"D9",X"FD",X"E5",X"D1",X"D9",X"7E",
		X"FE",X"FF",X"28",X"12",X"D9",X"62",X"6B",X"CD",X"51",X"3B",X"4E",X"23",X"46",X"D9",X"23",X"7E",
		X"D9",X"02",X"D9",X"23",X"18",X"E9",X"23",X"D1",X"E5",X"C9",X"DD",X"E1",X"48",X"DD",X"5E",X"00",
		X"CD",X"65",X"3B",X"DD",X"5E",X"01",X"FD",X"E5",X"16",X"00",X"FD",X"19",X"FD",X"7E",X"00",X"77",
		X"23",X"FD",X"7E",X"01",X"77",X"FD",X"E1",X"DD",X"5E",X"02",X"FD",X"E5",X"FD",X"19",X"FD",X"7E",
		X"00",X"23",X"77",X"23",X"FD",X"7E",X"01",X"77",X"1E",X"03",X"DD",X"19",X"FD",X"E1",X"DD",X"E5",
		X"C9",X"DD",X"E1",X"FD",X"E5",X"E1",X"16",X"00",X"DD",X"5E",X"01",X"19",X"E5",X"48",X"DD",X"5E",
		X"00",X"CD",X"65",X"3B",X"16",X"00",X"1E",X"02",X"19",X"D1",X"1A",X"77",X"13",X"23",X"1A",X"77",
		X"16",X"00",X"1E",X"02",X"DD",X"19",X"DD",X"E5",X"C9",X"DD",X"E1",X"DD",X"5E",X"00",X"48",X"CD",
		X"65",X"3B",X"EB",X"21",X"0D",X"00",X"19",X"FD",X"7E",X"00",X"77",X"FD",X"7E",X"01",X"23",X"77",
		X"21",X"0F",X"00",X"19",X"FD",X"7E",X"0A",X"77",X"FD",X"7E",X"0B",X"23",X"77",X"DD",X"23",X"DD",
		X"E5",X"C9",X"DD",X"E1",X"26",X"00",X"68",X"29",X"54",X"5D",X"29",X"29",X"19",X"E5",X"DD",X"6E",
		X"00",X"26",X"00",X"54",X"5D",X"29",X"29",X"19",X"D1",X"19",X"11",X"44",X"82",X"19",X"DD",X"5E",
		X"01",X"16",X"00",X"FD",X"E5",X"FD",X"19",X"FD",X"7E",X"00",X"77",X"23",X"FD",X"7E",X"01",X"77",
		X"1E",X"02",X"19",X"FD",X"E1",X"FD",X"E5",X"DD",X"5E",X"02",X"FD",X"19",X"FD",X"7E",X"01",X"77",
		X"2B",X"FD",X"7E",X"00",X"77",X"23",X"23",X"72",X"1E",X"03",X"DD",X"19",X"FD",X"E1",X"DD",X"E5",
		X"C9",X"85",X"6F",X"D0",X"24",X"C9",X"C5",X"42",X"21",X"00",X"00",X"54",X"78",X"B7",X"28",X"03",
		X"19",X"10",X"FD",X"C1",X"C9",X"21",X"F2",X"3C",X"16",X"00",X"19",X"56",X"21",X"E6",X"3C",X"79",
		X"CB",X"27",X"5F",X"7A",X"16",X"00",X"19",X"5E",X"23",X"56",X"6F",X"26",X"00",X"19",X"11",X"40",
		X"80",X"19",X"C9",X"00",X"80",X"01",X"80",X"06",X"80",X"07",X"80",X"F7",X"FE",X"08",X"80",X"0B",
		X"80",X"0C",X"80",X"0D",X"80",X"0E",X"80",X"F0",X"00",X"48",X"80",X"59",X"80",X"6A",X"80",X"7B",
		X"80",X"8C",X"80",X"44",X"80",X"55",X"80",X"66",X"80",X"77",X"80",X"88",X"80",X"3E",X"82",X"F4",
		X"82",X"02",X"80",X"03",X"80",X"06",X"80",X"07",X"80",X"EF",X"FD",X"09",X"80",X"0B",X"80",X"0C",
		X"80",X"0D",X"80",X"0E",X"80",X"0F",X"00",X"9D",X"80",X"AE",X"80",X"BF",X"80",X"D0",X"80",X"E1",
		X"80",X"99",X"80",X"AA",X"80",X"BB",X"80",X"CC",X"80",X"DD",X"80",X"3F",X"82",X"F7",X"82",X"04",
		X"80",X"05",X"80",X"06",X"80",X"07",X"80",X"DF",X"FB",X"0A",X"80",X"0B",X"80",X"0C",X"80",X"0D",
		X"80",X"0F",X"80",X"F0",X"00",X"F2",X"80",X"03",X"81",X"14",X"81",X"25",X"81",X"36",X"81",X"EE",
		X"80",X"FF",X"80",X"10",X"81",X"21",X"81",X"32",X"81",X"40",X"82",X"FA",X"82",X"10",X"80",X"11",
		X"80",X"16",X"80",X"17",X"80",X"F7",X"FE",X"18",X"80",X"1B",X"80",X"1C",X"80",X"1D",X"80",X"1E",
		X"80",X"F0",X"00",X"47",X"81",X"58",X"81",X"69",X"81",X"7A",X"81",X"8B",X"81",X"43",X"81",X"54",
		X"81",X"65",X"81",X"76",X"81",X"87",X"81",X"41",X"82",X"FD",X"82",X"12",X"80",X"13",X"80",X"16",
		X"80",X"17",X"80",X"EF",X"FD",X"19",X"80",X"1B",X"80",X"1C",X"80",X"1D",X"80",X"1E",X"80",X"0F",
		X"00",X"9C",X"81",X"AD",X"81",X"BE",X"81",X"CF",X"81",X"E0",X"81",X"98",X"81",X"A9",X"81",X"BA",
		X"81",X"CB",X"81",X"DC",X"81",X"42",X"82",X"00",X"83",X"14",X"80",X"15",X"80",X"16",X"80",X"17",
		X"80",X"DF",X"FB",X"1A",X"80",X"1B",X"80",X"1C",X"80",X"1D",X"80",X"1F",X"80",X"F0",X"00",X"F1",
		X"81",X"02",X"82",X"13",X"82",X"24",X"82",X"35",X"82",X"ED",X"81",X"FE",X"81",X"0F",X"82",X"20",
		X"82",X"31",X"82",X"43",X"82",X"03",X"83",X"80",X"00",X"00",X"01",X"00",X"02",X"00",X"03",X"00",
		X"04",X"00",X"05",X"00",X"06",X"00",X"07",X"00",X"08",X"00",X"09",X"00",X"0A",X"00",X"0B",X"00",
		X"0C",X"00",X"0D",X"00",X"0E",X"FF",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"01",X"03",X"07",X"0F",X"1F",X"3F",X"7F",X"FF",
		X"01",X"02",X"04",X"08",X"10",X"20",X"00",X"00",X"55",X"00",X"AA",X"00",X"FF",X"00",X"54",X"01",
		X"A9",X"01",X"00",X"11",X"22",X"33",X"44",X"2C",X"85",X"01",X"86",X"01",X"03",X"05",X"0D",X"86",
		X"08",X"0E",X"07",X"07",X"03",X"07",X"06",X"07",X"07",X"02",X"8C",X"4A",X"08",X"0F",X"03",X"0A",
		X"F6",X"84",X"0B",X"F5",X"41",X"03",X"0D",X"08",X"0B",X"FD",X"84",X"07",X"01",X"03",X"0B",X"FC",
		X"35",X"07",X"02",X"03",X"0B",X"2B",X"87",X"02",X"F3",X"92",X"3D",X"01",X"8A",X"0B",X"2D",X"8C",
		X"02",X"EA",X"89",X"3D",X"13",X"00",X"07",X"04",X"07",X"08",X"03",X"09",X"FC",X"04",X"0B",X"DE",
		X"92",X"21",X"0B",X"20",X"81",X"0B",X"F9",X"86",X"08",X"07",X"06",X"0A",X"03",X"02",X"08",X"2C",
		X"01",X"79",X"0B",X"DF",X"89",X"02",X"C5",X"24",X"06",X"0B",X"03",X"01",X"33",X"0B",X"E0",X"C4",
		X"21",X"0B",X"20",X"81",X"0B",X"F7",X"9F",X"0B",X"2C",X"12",X"0B",X"28",X"0F",X"0B",X"F6",X"87",
		X"1F",X"07",X"01",X"A0",X"01",X"06",X"1F",X"DB",X"02",X"A2",X"7A",X"0B",X"29",X"77",X"07",X"04",
		X"06",X"01",X"03",X"01",X"14",X"0B",X"F9",X"96",X"1F",X"06",X"0B",X"2C",X"68",X"0B",X"28",X"65",
		X"0B",X"F6",X"62",X"0B",X"29",X"5F",X"07",X"03",X"06",X"0C",X"03",X"0D",X"08",X"02",X"3D",X"55",
		X"21",X"01",X"68",X"0B",X"E1",X"A9",X"21",X"0B",X"28",X"4B",X"0A",X"F6",X"91",X"1F",X"D3",X"02",
		X"6B",X"43",X"0B",X"29",X"40",X"0B",X"2C",X"3D",X"0B",X"F7",X"3A",X"01",X"42",X"0B",X"29",X"35",
		X"0B",X"2C",X"32",X"0A",X"F7",X"84",X"02",X"14",X"2C",X"21",X"01",X"4B",X"01",X"27",X"0B",X"E2",
		X"B2",X"0B",X"20",X"81",X"0B",X"FA",X"8C",X"0B",X"2C",X"73",X"1F",X"EB",X"0B",X"FE",X"6E",X"06",
		X"01",X"03",X"0B",X"F9",X"8B",X"0B",X"2C",X"65",X"0B",X"F9",X"62",X"1F",X"08",X"01",X"71",X"0B",
		X"28",X"5B",X"0B",X"F8",X"58",X"0B",X"29",X"55",X"0B",X"2C",X"52",X"1F",X"E3",X"02",X"05",X"5D",
		X"01",X"5E",X"0B",X"E3",X"8A",X"02",X"15",X"45",X"3D",X"07",X"03",X"06",X"0D",X"03",X"04",X"04",
		X"00",X"00",X"00",X"00",X"69",X"60",X"4E",X"23",X"46",X"1A",X"81",X"6F",X"13",X"1A",X"88",X"67",
		X"C9",X"EB",X"5F",X"16",X"00",X"EB",X"1A",X"85",X"6F",X"13",X"1A",X"8C",X"67",X"C9",X"EB",X"5F",
		X"16",X"00",X"EB",X"1A",X"A5",X"6F",X"13",X"1A",X"A4",X"67",X"C9",X"44",X"4D",X"21",X"00",X"00",
		X"3E",X"10",X"F5",X"29",X"EB",X"97",X"29",X"EB",X"8D",X"91",X"6F",X"7C",X"98",X"67",X"13",X"D2",
		X"54",X"3E",X"09",X"1B",X"F1",X"3D",X"C2",X"42",X"3E",X"C9",X"5E",X"23",X"56",X"EB",X"29",X"E5",
		X"29",X"29",X"C1",X"09",X"C9",X"44",X"4D",X"21",X"00",X"00",X"3E",X"10",X"29",X"EB",X"29",X"EB",
		X"D2",X"74",X"3E",X"09",X"3D",X"C2",X"6C",X"3E",X"C9",X"59",X"50",X"EB",X"97",X"95",X"6F",X"3E",
		X"00",X"9C",X"67",X"C9",X"EB",X"5F",X"16",X"00",X"EB",X"1A",X"B5",X"6F",X"13",X"1A",X"B4",X"67",
		X"C9",X"5F",X"16",X"00",X"7B",X"95",X"6F",X"7A",X"9C",X"67",X"C9",X"4F",X"06",X"00",X"7B",X"91",
		X"6F",X"7A",X"98",X"67",X"C9",X"69",X"60",X"4E",X"23",X"46",X"1A",X"91",X"6F",X"13",X"1A",X"98",
		X"67",X"C9",X"6F",X"26",X"00",X"1A",X"95",X"6F",X"13",X"1A",X"9C",X"67",X"C9",X"5F",X"16",X"00",
		X"7B",X"96",X"5F",X"7A",X"23",X"9E",X"57",X"EB",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"2D",X"99",X"2D",X"99",
		X"2D",X"99",X"2D",X"26",X"1E",X"99",X"2D",X"94",X"2B",X"F2",X"28",X"F2",X"28",X"00",X"00",X"C9",
		X"2E",X"26",X"1E",X"BE",X"1F",X"FF",X"FF",X"70",X"03",X"01",X"07",X"00",X"04",X"23",X"00",X"6D",
		X"36",X"BE",X"39",X"B7",X"0F",X"5B",X"3E",X"17",X"35",X"24",X"35",X"4F",X"37",X"5C",X"40",X"E4",
		X"3E",X"62",X"3F",X"C2",X"3A",X"BC",X"3B",X"3E",X"00",X"C8",X"39",X"B8",X"3A",X"C1",X"FC",X"35",
		X"F7",X"07",X"C5",X"54",X"55",X"4C",X"4F",X"53",X"42",X"41",X"A2",X"3C",X"A9",X"00",X"C3",X"44",
		X"41",X"82",X"35",X"DC",X"88",X"4A",X"C4",X"44",X"41",X"34",X"11",X"DB",X"80",X"09",X"C6",X"41",
		X"64",X"36",X"F9",X"30",X"C4",X"4E",X"41",X"60",X"00",X"DA",X"A0",X"C9",X"49",X"43",X"53",X"41",
		X"F6",X"22",X"82",X"D4",X"45",X"53",X"41",X"C0",X"23",X"94",X"C2",X"EC",X"22",X"F5",X"00",X"C5",
		X"53",X"41",X"42",X"77",X"36",X"A6",X"C3",X"42",X"D8",X"3A",X"FB",X"00",X"D4",X"49",X"42",X"36",
		X"35",X"D8",X"40",X"CB",X"43",X"4F",X"4C",X"42",X"88",X"00",X"83",X"C5",X"54",X"59",X"42",X"F4",
		X"3D",X"84",X"C3",X"A7",X"35",X"F6",X"01",X"CC",X"4C",X"41",X"43",X"AF",X"00",X"D6",X"CD",X"C6",
		X"43",X"43",X"A8",X"00",X"D1",X"3F",X"C4",X"4E",X"43",X"40",X"35",X"96",X"08",X"CE",X"4F",X"4D",
		X"4D",X"4F",X"43",X"75",X"37",X"A2",X"02",X"CE",X"4F",X"43",X"11",X"3A",X"96",X"20",X"D0",X"43",
		X"D3",X"00",X"DA",X"B8",X"C4",X"50",X"43",X"0B",X"3B",X"D2",X"A9",X"D2",X"44",X"50",X"43",X"22",
		X"39",X"D2",X"B9",X"C9",X"50",X"43",X"57",X"38",X"D2",X"A1",X"D2",X"49",X"50",X"43",X"B1",X"35");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
