library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity dderby_sp_bits_4 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of dderby_sp_bits_4 is
	type rom is array(0 to  32767) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"99",X"99",X"99",X"00",X"77",X"77",X"22",X"00",X"26",X"22",X"99",
		X"00",X"22",X"22",X"99",X"00",X"77",X"97",X"22",X"00",X"02",X"97",X"66",X"00",X"02",X"27",X"66",
		X"00",X"77",X"26",X"66",X"00",X"77",X"22",X"66",X"00",X"22",X"26",X"66",X"00",X"62",X"92",X"66",
		X"00",X"26",X"92",X"66",X"00",X"22",X"26",X"66",X"00",X"77",X"22",X"66",X"00",X"77",X"26",X"66",
		X"00",X"02",X"27",X"66",X"00",X"02",X"97",X"66",X"00",X"77",X"97",X"22",X"00",X"22",X"22",X"99",
		X"00",X"26",X"22",X"99",X"00",X"77",X"77",X"22",X"00",X"99",X"99",X"99",X"00",X"00",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"90",X"00",X"00",X"77",X"97",X"00",X"00",X"27",X"77",X"00",X"00",X"67",X"66",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",
		X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"62",X"00",X"00",
		X"99",X"26",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",
		X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"99",X"00",X"00",
		X"67",X"66",X"00",X"00",X"27",X"77",X"00",X"00",X"77",X"97",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"79",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"62",X"00",
		X"00",X"00",X"26",X"00",X"00",X"00",X"22",X"00",X"00",X"09",X"99",X"97",X"00",X"09",X"22",X"27",
		X"00",X"77",X"22",X"79",X"00",X"77",X"72",X"97",X"00",X"97",X"77",X"99",X"00",X"97",X"29",X"22",
		X"00",X"97",X"29",X"66",X"00",X"90",X"99",X"66",X"00",X"00",X"99",X"66",X"00",X"02",X"99",X"66",
		X"00",X"22",X"27",X"66",X"00",X"29",X"29",X"66",X"00",X"66",X"29",X"66",X"00",X"72",X"22",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"29",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"62",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"66",X"99",X"00",X"00",
		X"27",X"99",X"00",X"00",X"29",X"66",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"99",X"00",X"00",
		X"00",X"07",X"27",X"66",X"00",X"00",X"22",X"66",X"00",X"00",X"22",X"66",X"00",X"00",X"27",X"66",
		X"00",X"00",X"72",X"22",X"00",X"00",X"79",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"76",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"22",X"90",X"00",X"99",X"22",X"90",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",
		X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"97",X"67",X"00",X"00",X"92",X"26",X"00",X"00",
		X"72",X"62",X"00",X"00",X"22",X"27",X"00",X"00",X"22",X"27",X"00",X"00",X"29",X"27",X"00",X"00",
		X"22",X"70",X"00",X"00",X"76",X"70",X"00",X"00",X"99",X"70",X"00",X"00",X"99",X"00",X"00",X"00",
		X"09",X"69",X"00",X"00",X"00",X"79",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"07",X"00",X"00",X"00",X"02",X"90",X"00",X"00",X"72",X"97",X"00",X"00",X"27",X"99",
		X"00",X"00",X"77",X"29",X"00",X"00",X"22",X"22",X"00",X"EE",X"22",X"22",X"00",X"EE",X"66",X"22",
		X"00",X"E3",X"69",X"99",X"00",X"37",X"29",X"67",X"00",X"26",X"22",X"99",X"00",X"22",X"29",X"92",
		X"00",X"92",X"29",X"96",X"00",X"09",X"92",X"66",X"00",X"09",X"22",X"66",X"00",X"07",X"29",X"66",
		X"00",X"00",X"27",X"66",X"00",X"00",X"26",X"66",X"00",X"00",X"29",X"66",X"00",X"00",X"27",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"79",X"00",X"00",X"00",X"27",X"00",X"00",X"00",
		X"62",X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"66",X"00",X"00",X"00",
		X"00",X"00",X"27",X"66",X"00",X"00",X"22",X"66",X"00",X"00",X"92",X"66",X"00",X"00",X"92",X"66",
		X"00",X"00",X"09",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"72",
		X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"79",X"00",X"00",X"97",X"67",X"00",X"00",X"92",X"67",X"00",X"00",
		X"22",X"26",X"00",X"00",X"22",X"92",X"00",X"00",X"22",X"29",X"00",X"00",X"29",X"29",X"00",X"00",
		X"92",X"97",X"00",X"00",X"22",X"70",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"09",X"00",X"00",
		X"22",X"09",X"00",X"00",X"92",X"99",X"00",X"00",X"92",X"90",X"00",X"00",X"29",X"00",X"00",X"00",
		X"62",X"00",X"00",X"00",X"76",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",
		X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"07",X"00",X"00",X"09",X"02",X"00",X"00",X"97",X"02",X"00",X"00",X"97",X"29",
		X"00",X"00",X"09",X"29",X"00",X"00",X"92",X"72",X"00",X"00",X"92",X"72",X"00",X"00",X"92",X"72",
		X"00",X"00",X"29",X"22",X"00",X"00",X"29",X"29",X"00",X"00",X"29",X"92",X"00",X"00",X"22",X"22",
		X"00",X"00",X"62",X"99",X"00",X"00",X"29",X"62",X"00",X"00",X"29",X"99",X"00",X"00",X"22",X"99",
		X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"66",X"00",X"00",X"22",X"66",
		X"00",X"00",X"22",X"66",X"00",X"00",X"92",X"66",X"00",X"00",X"92",X"66",X"00",X"00",X"97",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",X"00",X"00",X"00",
		X"70",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"27",X"00",X"00",X"00",X"27",X"00",X"00",X"00",
		X"27",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"96",X"00",X"00",X"00",
		X"00",X"00",X"09",X"66",X"00",X"00",X"09",X"66",X"00",X"00",X"09",X"66",X"00",X"00",X"00",X"66",
		X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"27",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"96",
		X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"96",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"26",X"00",X"00",X"00",
		X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"97",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"27",X"00",X"00",X"00",X"79",X"00",X"00",X"00",X"92",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"22",X"90",X"00",X"00",X"22",X"90",X"00",X"00",X"22",X"90",X"00",X"00",
		X"22",X"00",X"00",X"00",X"62",X"00",X"00",X"00",X"22",X"70",X"00",X"00",X"77",X"70",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"E0",X"00",X"00",X"77",X"E3",X"00",
		X"09",X"76",X"99",X"00",X"09",X"22",X"62",X"00",X"09",X"26",X"62",X"00",X"09",X"22",X"22",X"00",
		X"09",X"26",X"62",X"00",X"09",X"22",X"22",X"00",X"77",X"26",X"67",X"00",X"99",X"22",X"27",X"00",
		X"99",X"29",X"67",X"00",X"99",X"29",X"27",X"00",X"99",X"99",X"67",X"00",X"99",X"29",X"27",X"00",
		X"99",X"77",X"27",X"00",X"97",X"62",X"22",X"00",X"97",X"99",X"22",X"00",X"07",X"99",X"92",X"00",
		X"07",X"99",X"27",X"00",X"07",X"77",X"79",X"00",X"07",X"66",X"97",X"00",X"09",X"66",X"62",X"00",
		X"09",X"66",X"22",X"00",X"09",X"66",X"22",X"00",X"09",X"66",X"92",X"00",X"09",X"66",X"92",X"00",
		X"09",X"66",X"92",X"00",X"09",X"66",X"96",X"00",X"09",X"66",X"96",X"00",X"09",X"66",X"96",X"00",
		X"09",X"66",X"96",X"00",X"09",X"22",X"96",X"00",X"09",X"99",X"97",X"00",X"09",X"99",X"27",X"00",
		X"09",X"99",X"27",X"00",X"09",X"99",X"27",X"00",X"09",X"99",X"77",X"00",X"99",X"77",X"67",X"00",
		X"99",X"22",X"67",X"00",X"99",X"22",X"67",X"00",X"99",X"79",X"67",X"00",X"99",X"26",X"67",X"00",
		X"99",X"22",X"67",X"00",X"99",X"26",X"67",X"00",X"97",X"22",X"67",X"00",X"97",X"26",X"67",X"00",
		X"07",X"22",X"67",X"00",X"07",X"99",X"67",X"00",X"09",X"77",X"67",X"00",X"00",X"00",X"69",X"00",
		X"00",X"99",X"69",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"9A",X"00",X"00",X"00",X"AC",X"00",X"00",X"00",X"BA",X"00",
		X"00",X"00",X"AD",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",
		X"00",X"09",X"00",X"00",X"00",X"9A",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"15",X"00",X"00",
		X"00",X"11",X"00",X"00",X"09",X"51",X"00",X"00",X"91",X"51",X"00",X"00",X"11",X"09",X"00",X"00",
		X"14",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"90",X"00",X"00",X"11",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"19",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"9D",X"00",
		X"00",X"00",X"DA",X"00",X"00",X"00",X"AD",X"00",X"00",X"00",X"D9",X"00",X"00",X"09",X"99",X"00",
		X"00",X"9A",X"99",X"00",X"00",X"AD",X"90",X"00",X"00",X"AD",X"00",X"00",X"99",X"A9",X"00",X"00",
		X"DD",X"D9",X"00",X"00",X"DA",X"DD",X"00",X"00",X"AA",X"DD",X"00",X"00",X"AA",X"DD",X"00",X"00",
		X"A9",X"DD",X"00",X"00",X"A9",X"D9",X"00",X"00",X"DA",X"D9",X"00",X"00",X"DA",X"99",X"00",X"00",
		X"DD",X"90",X"00",X"00",X"9D",X"90",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"90",X"00",X"00",X"77",X"97",X"00",X"00",X"27",X"72",X"00",X"00",X"67",X"62",X"00",X"00",
		X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",
		X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"69",X"00",X"00",
		X"99",X"29",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"67",X"99",X"00",X"00",X"27",X"66",X"00",X"00",X"77",X"97",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"29",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"62",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"66",X"99",X"00",X"00",
		X"27",X"99",X"00",X"00",X"29",X"66",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",
		X"99",X"22",X"90",X"00",X"99",X"22",X"90",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"97",X"97",X"00",X"00",X"92",X"99",X"00",X"00",
		X"72",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"97",X"00",X"00",X"29",X"97",X"00",X"00",
		X"22",X"70",X"00",X"00",X"76",X"70",X"00",X"00",X"99",X"70",X"00",X"00",X"99",X"00",X"00",X"00",
		X"09",X"69",X"00",X"00",X"00",X"79",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"79",X"00",X"00",X"97",X"67",X"00",X"00",X"92",X"67",X"00",X"00",
		X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"29",X"22",X"00",X"00",
		X"92",X"97",X"00",X"00",X"22",X"90",X"00",X"00",X"29",X"99",X"00",X"00",X"99",X"09",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",
		X"69",X"00",X"00",X"00",X"76",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",
		X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"96",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"26",X"00",X"00",X"00",
		X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"27",X"00",X"00",X"00",X"79",X"00",X"00",X"00",X"92",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"22",X"90",X"00",X"00",X"22",X"90",X"00",X"00",X"22",X"20",X"00",X"00",
		X"99",X"20",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"70",X"00",X"00",X"77",X"70",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"66",X"00",X"00",X"09",X"66",X"00",X"00",X"09",X"66",X"00",X"00",X"00",X"66",
		X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"27",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"66",
		X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"66",X"92",X"00",X"09",X"66",X"96",X"00",X"09",X"66",X"96",X"00",X"09",X"66",X"96",X"00",
		X"09",X"66",X"96",X"00",X"09",X"22",X"96",X"00",X"09",X"99",X"97",X"00",X"09",X"99",X"27",X"00",
		X"09",X"99",X"27",X"00",X"09",X"99",X"27",X"00",X"09",X"99",X"77",X"00",X"99",X"77",X"67",X"00",
		X"99",X"22",X"67",X"00",X"99",X"22",X"67",X"00",X"99",X"79",X"67",X"00",X"99",X"26",X"97",X"00",
		X"99",X"22",X"97",X"00",X"99",X"99",X"29",X"00",X"96",X"99",X"27",X"00",X"96",X"99",X"27",X"00",
		X"07",X"99",X"22",X"00",X"07",X"99",X"22",X"00",X"09",X"77",X"97",X"00",X"00",X"09",X"69",X"00",
		X"00",X"99",X"69",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"99",X"99",X"99",X"00",X"E9",X"77",X"22",X"00",X"EE",X"22",X"99",
		X"00",X"E3",X"22",X"99",X"00",X"32",X"97",X"22",X"00",X"09",X"27",X"66",X"00",X"09",X"27",X"66",
		X"00",X"77",X"22",X"66",X"00",X"9D",X"22",X"66",X"00",X"9D",X"92",X"66",X"00",X"99",X"92",X"66",
		X"00",X"99",X"92",X"66",X"00",X"99",X"92",X"66",X"00",X"9D",X"92",X"66",X"00",X"7D",X"22",X"66",
		X"00",X"09",X"97",X"66",X"00",X"09",X"97",X"66",X"00",X"22",X"97",X"22",X"00",X"22",X"22",X"99",
		X"00",X"26",X"22",X"99",X"00",X"77",X"77",X"22",X"00",X"99",X"99",X"99",X"00",X"00",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"79",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"09",X"99",X"00",X"00",X"09",X"22",X"00",X"00",X"09",X"62",X"97",X"00",X"09",X"99",X"27",
		X"00",X"07",X"99",X"79",X"00",X"09",X"99",X"97",X"00",X"07",X"DD",X"99",X"00",X"07",X"DD",X"22",
		X"00",X"97",X"92",X"66",X"00",X"90",X"92",X"66",X"00",X"30",X"22",X"66",X"00",X"32",X"29",X"66",
		X"00",X"32",X"27",X"66",X"00",X"22",X"29",X"66",X"00",X"66",X"29",X"66",X"00",X"72",X"22",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"00",
		X"00",X"00",X"07",X"00",X"00",X"00",X"09",X"90",X"00",X"00",X"D9",X"97",X"00",X"00",X"D9",X"99",
		X"00",X"00",X"DD",X"29",X"00",X"09",X"9D",X"22",X"00",X"09",X"DD",X"22",X"00",X"EE",X"D9",X"22",
		X"00",X"EE",X"9D",X"99",X"00",X"E3",X"DD",X"67",X"00",X"33",X"D2",X"99",X"00",X"22",X"22",X"92",
		X"00",X"92",X"99",X"96",X"00",X"09",X"92",X"66",X"00",X"09",X"22",X"66",X"00",X"07",X"29",X"66",
		X"00",X"00",X"27",X"66",X"00",X"00",X"26",X"66",X"00",X"00",X"29",X"66",X"00",X"00",X"27",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",X"00",X"00",X"00",
		X"70",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"27",X"00",X"00",X"00",X"27",X"00",X"00",X"00",
		X"27",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"96",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"03",X"00",X"00",X"90",X"02",X"00",X"00",X"90",X"92",
		X"00",X"00",X"09",X"96",X"00",X"00",X"99",X"92",X"00",X"00",X"9D",X"96",X"00",X"00",X"99",X"99",
		X"00",X"00",X"29",X"99",X"00",X"00",X"29",X"29",X"00",X"00",X"29",X"22",X"00",X"00",X"22",X"99",
		X"00",X"00",X"62",X"99",X"00",X"00",X"22",X"62",X"00",X"00",X"29",X"99",X"00",X"00",X"22",X"99",
		X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"66",X"00",X"00",X"22",X"66",
		X"00",X"00",X"22",X"66",X"00",X"00",X"92",X"66",X"00",X"00",X"92",X"66",X"00",X"00",X"97",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"99",X"00",
		X"09",X"09",X"99",X"00",X"09",X"99",X"33",X"00",X"09",X"99",X"92",X"00",X"09",X"D9",X"26",X"00",
		X"09",X"DD",X"62",X"00",X"09",X"D9",X"29",X"00",X"77",X"DD",X"29",X"00",X"99",X"D9",X"99",X"00",
		X"99",X"2D",X"99",X"00",X"99",X"29",X"97",X"00",X"99",X"29",X"67",X"00",X"99",X"92",X"27",X"00",
		X"99",X"77",X"27",X"00",X"97",X"62",X"22",X"00",X"97",X"99",X"22",X"00",X"07",X"99",X"92",X"00",
		X"07",X"99",X"27",X"00",X"07",X"77",X"79",X"00",X"07",X"66",X"97",X"00",X"09",X"66",X"62",X"00",
		X"09",X"66",X"22",X"00",X"09",X"66",X"22",X"00",X"09",X"66",X"92",X"00",X"09",X"66",X"92",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E9",X"09",X"99",X"00",X"EE",X"77",X"22",X"00",X"E3",X"22",X"99",
		X"00",X"32",X"22",X"99",X"00",X"22",X"97",X"22",X"00",X"09",X"27",X"66",X"00",X"09",X"27",X"66",
		X"00",X"77",X"22",X"66",X"00",X"9D",X"22",X"66",X"00",X"9D",X"92",X"66",X"00",X"99",X"92",X"66",
		X"00",X"99",X"92",X"66",X"00",X"99",X"92",X"66",X"00",X"9D",X"92",X"66",X"00",X"7D",X"22",X"66",
		X"00",X"09",X"97",X"66",X"00",X"09",X"97",X"66",X"00",X"32",X"97",X"22",X"00",X"32",X"22",X"99",
		X"00",X"36",X"22",X"99",X"00",X"77",X"77",X"22",X"00",X"99",X"99",X"99",X"00",X"00",X"90",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"29",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"62",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"66",X"99",X"00",X"00",
		X"27",X"99",X"00",X"00",X"29",X"66",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",
		X"00",X"09",X"99",X"00",X"00",X"09",X"22",X"00",X"00",X"09",X"62",X"97",X"00",X"09",X"99",X"27",
		X"00",X"07",X"99",X"79",X"00",X"09",X"99",X"97",X"00",X"07",X"DD",X"99",X"00",X"07",X"DD",X"22",
		X"00",X"97",X"92",X"66",X"00",X"30",X"92",X"66",X"00",X"30",X"22",X"66",X"00",X"32",X"29",X"66",
		X"00",X"32",X"27",X"66",X"00",X"32",X"29",X"66",X"00",X"66",X"29",X"66",X"00",X"72",X"22",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"00",
		X"00",X"00",X"07",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"D9",X"99",
		X"00",X"00",X"DD",X"29",X"00",X"09",X"9D",X"22",X"00",X"09",X"DD",X"22",X"00",X"EE",X"D9",X"22",
		X"00",X"EE",X"9D",X"99",X"00",X"EE",X"DD",X"67",X"00",X"26",X"D2",X"99",X"00",X"22",X"22",X"92",
		X"00",X"92",X"99",X"96",X"00",X"99",X"92",X"66",X"00",X"99",X"22",X"66",X"00",X"99",X"29",X"66",
		X"00",X"09",X"27",X"66",X"00",X"09",X"26",X"66",X"00",X"00",X"29",X"66",X"00",X"00",X"27",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",X"00",X"00",X"00",
		X"70",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"27",X"00",X"00",X"00",X"27",X"00",X"00",X"00",
		X"27",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"96",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",
		X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"03",X"00",X"00",X"90",X"02",X"00",X"00",X"90",X"92",
		X"00",X"00",X"09",X"96",X"00",X"00",X"99",X"92",X"00",X"00",X"9D",X"96",X"00",X"00",X"99",X"99",
		X"00",X"00",X"29",X"99",X"00",X"00",X"29",X"29",X"00",X"00",X"29",X"22",X"00",X"00",X"22",X"99",
		X"00",X"00",X"62",X"99",X"00",X"00",X"22",X"62",X"00",X"00",X"29",X"99",X"00",X"00",X"22",X"99",
		X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"66",X"00",X"00",X"22",X"66",
		X"00",X"00",X"22",X"66",X"00",X"00",X"92",X"66",X"00",X"00",X"92",X"66",X"00",X"00",X"97",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"99",X"00",
		X"09",X"09",X"99",X"00",X"09",X"99",X"62",X"00",X"09",X"99",X"92",X"00",X"09",X"D9",X"26",X"00",
		X"09",X"DD",X"62",X"00",X"09",X"D9",X"29",X"00",X"77",X"DD",X"29",X"00",X"99",X"D9",X"99",X"00",
		X"99",X"2D",X"99",X"00",X"99",X"29",X"97",X"00",X"99",X"29",X"67",X"00",X"99",X"92",X"27",X"00",
		X"99",X"77",X"27",X"00",X"97",X"62",X"22",X"00",X"97",X"99",X"22",X"00",X"07",X"99",X"92",X"00",
		X"07",X"99",X"27",X"00",X"07",X"77",X"79",X"00",X"07",X"66",X"97",X"00",X"09",X"66",X"62",X"00",
		X"09",X"66",X"22",X"00",X"09",X"66",X"22",X"00",X"09",X"66",X"92",X"00",X"09",X"66",X"92",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"90",X"00",X"00",X"77",X"97",X"00",X"00",X"27",X"77",X"00",X"00",X"67",X"77",X"00",X"00",
		X"99",X"92",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",
		X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"62",X"00",X"00",X"99",X"22",X"00",X"00",
		X"99",X"29",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"67",X"99",X"00",X"00",X"27",X"66",X"00",X"00",X"77",X"07",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"22",X"90",X"00",X"99",X"22",X"90",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",
		X"99",X"22",X"00",X"00",X"99",X"29",X"00",X"00",X"97",X"99",X"00",X"00",X"92",X"99",X"00",X"00",
		X"72",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"97",X"00",X"00",X"29",X"97",X"00",X"00",
		X"22",X"70",X"00",X"00",X"76",X"70",X"00",X"00",X"09",X"70",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"69",X"00",X"00",X"00",X"79",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"27",X"66",X"00",X"99",X"22",X"66",X"00",X"09",X"22",X"66",X"00",X"00",X"27",X"66",
		X"00",X"00",X"72",X"22",X"00",X"00",X"79",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"76",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"97",X"69",X"00",X"00",X"92",X"69",X"00",X"00",X"22",X"22",X"00",X"00",
		X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"29",X"99",X"00",X"00",X"92",X"97",X"00",X"00",
		X"22",X"90",X"00",X"00",X"22",X"99",X"00",X"00",X"99",X"09",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"69",X"00",X"00",X"00",
		X"76",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"07",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"96",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"26",X"00",X"00",X"00",
		X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"27",X"00",X"00",X"00",X"79",X"90",X"00",X"00",X"92",X"90",X"00",X"00",
		X"22",X"90",X"00",X"00",X"22",X"90",X"00",X"00",X"22",X"90",X"00",X"00",X"22",X"00",X"00",X"00",
		X"22",X"20",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"70",X"00",X"00",X"77",X"70",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"66",X"00",X"00",X"09",X"66",X"00",X"00",X"09",X"66",X"00",X"00",X"00",X"66",
		X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"27",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"66",
		X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"66",X"92",X"00",X"09",X"66",X"96",X"00",X"09",X"66",X"96",X"00",X"09",X"66",X"96",X"00",
		X"09",X"66",X"96",X"00",X"09",X"22",X"96",X"00",X"09",X"99",X"97",X"00",X"09",X"99",X"27",X"00",
		X"09",X"99",X"27",X"00",X"09",X"99",X"27",X"00",X"09",X"99",X"77",X"00",X"09",X"77",X"67",X"00",
		X"09",X"22",X"67",X"00",X"09",X"22",X"67",X"00",X"09",X"79",X"67",X"00",X"09",X"22",X"97",X"00",
		X"09",X"22",X"27",X"00",X"09",X"22",X"29",X"00",X"06",X"99",X"27",X"00",X"06",X"99",X"22",X"00",
		X"09",X"99",X"92",X"00",X"09",X"99",X"99",X"00",X"09",X"77",X"97",X"00",X"00",X"09",X"69",X"00",
		X"00",X"99",X"69",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"91",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"10",X"00",
		X"00",X"00",X"10",X"00",X"00",X"01",X"21",X"00",X"00",X"10",X"29",X"00",X"00",X"10",X"11",X"00",
		X"01",X"91",X"11",X"00",X"00",X"12",X"02",X"00",X"00",X"12",X"0F",X"00",X"00",X"21",X"09",X"00",
		X"00",X"11",X"F1",X"10",X"09",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"0F",X"90",X"00",X"01",X"21",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"10",X"00",X"00",
		X"10",X"11",X"00",X"11",X"11",X"02",X"10",X"11",X"92",X"90",X"10",X"00",X"92",X"00",X"01",X"00",
		X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"01",X"00",X"10",X"99",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"91",X"00",X"00",X"00",
		X"01",X"09",X"10",X"00",X"22",X"20",X"11",X"00",X"11",X"11",X"00",X"00",X"10",X"01",X"90",X"00",
		X"00",X"00",X"99",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"11",X"00",X"10",X"00",X"11",X"00",X"11",X"00",X"01",X"00",X"11",X"00",X"02",
		X"00",X"11",X"01",X"10",X"00",X"19",X"10",X"11",X"00",X"91",X"00",X"11",X"00",X"11",X"10",X"10",
		X"00",X"90",X"00",X"10",X"00",X"09",X"00",X"10",X"00",X"01",X"99",X"91",X"00",X"01",X"19",X"90",
		X"00",X"11",X"00",X"00",X"00",X"10",X"99",X"99",X"99",X"01",X"99",X"99",X"09",X"10",X"09",X"99",
		X"10",X"11",X"99",X"99",X"11",X"11",X"99",X"90",X"00",X"00",X"99",X"00",X"10",X"00",X"99",X"00",
		X"11",X"09",X"00",X"09",X"11",X"09",X"00",X"00",X"11",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"01",X"00",X"10",X"90",X"11",X"00",
		X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"10",X"00",X"11",X"00",X"09",X"00",
		X"00",X"00",X"00",X"00",X"01",X"09",X"90",X"00",X"01",X"99",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"90",X"00",X"01",X"00",X"99",X"00",X"11",X"99",X"99",X"00",X"10",X"99",X"99",X"20",X"00",
		X"99",X"90",X"10",X"00",X"99",X"91",X"00",X"11",X"90",X"99",X"11",X"10",X"00",X"10",X"00",X"00",
		X"00",X"10",X"19",X"90",X"00",X"20",X"99",X"90",X"00",X"01",X"00",X"00",X"00",X"01",X"99",X"00",
		X"19",X"09",X"00",X"00",X"00",X"91",X"00",X"00",X"11",X"99",X"00",X"00",X"01",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"11",X"99",X"00",X"00",X"01",X"90",X"00",X"00",
		X"11",X"00",X"10",X"00",X"01",X"01",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"10",X"00",X"00",X"99",X"12",X"00",X"99",X"99",X"10",X"11",X"00",X"99",X"00",X"00",X"10",
		X"00",X"01",X"10",X"00",X"00",X"00",X"11",X"00",X"00",X"09",X"19",X"09",X"09",X"19",X"00",X"99",
		X"00",X"11",X"99",X"09",X"11",X"11",X"90",X"09",X"00",X"01",X"99",X"09",X"00",X"09",X"99",X"99",
		X"11",X"99",X"00",X"99",X"00",X"91",X"90",X"09",X"99",X"91",X"11",X"11",X"99",X"00",X"11",X"00",
		X"00",X"99",X"90",X"99",X"99",X"90",X"90",X"99",X"99",X"00",X"90",X"09",X"99",X"99",X"99",X"00",
		X"09",X"10",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",
		X"09",X"10",X"00",X"00",X"90",X"10",X"10",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"11",X"00",
		X"00",X"00",X"11",X"00",X"00",X"90",X"01",X"00",X"99",X"90",X"01",X"10",X"11",X"00",X"99",X"99",
		X"10",X"00",X"99",X"00",X"11",X"10",X"99",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",
		X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"99",X"00",X"00",X"11",X"99",X"00",X"00",
		X"01",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"14",X"00",X"00",X"00",
		X"14",X"99",X"00",X"00",X"14",X"99",X"00",X"00",X"14",X"00",X"00",X"00",X"14",X"00",X"00",X"00",
		X"14",X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"19",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"14",X"14",X"00",X"00",X"41",X"11",X"00",
		X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"10",X"00",X"00",X"11",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"11",X"09",X"00",X"00",X"14",X"99",X"00",X"00",X"11",X"90",X"00",
		X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"11",X"11",X"00",
		X"11",X"11",X"00",X"00",X"11",X"11",X"99",X"00",X"91",X"11",X"99",X"00",X"09",X"11",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"10",X"00",X"00",
		X"00",X"10",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"1F",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"01",X"10",X"00",X"00",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"20",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"1F",X"00",X"00",
		X"00",X"21",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"90",X"00",X"00",X"99",X"FF",X"00",X"0F",X"99",X"09",X"00",
		X"9F",X"FF",X"F0",X"00",X"F0",X"0F",X"F0",X"00",X"FF",X"0F",X"F0",X"00",X"9F",X"F0",X"FF",X"00",
		X"99",X"09",X"09",X"00",X"09",X"00",X"9F",X"00",X"09",X"FF",X"9F",X"00",X"00",X"FF",X"9F",X"00",
		X"09",X"FF",X"90",X"00",X"00",X"FF",X"99",X"90",X"00",X"FF",X"09",X"90",X"09",X"99",X"FF",X"00",
		X"09",X"F9",X"FF",X"00",X"90",X"F9",X"F9",X"00",X"90",X"FF",X"00",X"00",X"F9",X"F0",X"FF",X"00",
		X"00",X"FF",X"FF",X"00",X"09",X"F9",X"F9",X"00",X"09",X"0F",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"F9",X"00",X"00",X"99",X"00",X"00",X"00",
		X"9F",X"0F",X"00",X"00",X"F9",X"FF",X"00",X"00",X"09",X"F9",X"00",X"00",X"F9",X"99",X"00",X"00",
		X"F0",X"90",X"00",X"00",X"9F",X"F9",X"00",X"00",X"90",X"FF",X"00",X"00",X"99",X"9F",X"90",X"00",
		X"9F",X"99",X"00",X"00",X"FF",X"F0",X"00",X"00",X"F0",X"FF",X"00",X"00",X"FF",X"F0",X"00",X"00",
		X"FF",X"F9",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"9F",X"F0",X"00",X"F9",X"99",X"90",X"00",
		X"F9",X"F0",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"F0",X"00",
		X"90",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"90",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"0F",X"00",X"F0",X"00",X"99",X"00",X"0F",X"00",X"99",X"F0",X"00",X"00",X"00",X"09",X"99",X"00",
		X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"A9",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"A9",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"DA",X"00",
		X"00",X"00",X"99",X"00",X"00",X"09",X"00",X"00",X"00",X"9A",X"00",X"00",X"00",X"AB",X"00",X"00",
		X"00",X"BD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"D9",X"00",X"00",
		X"00",X"99",X"00",X"00",X"AD",X"90",X"00",X"00",X"AA",X"00",X"00",X"00",X"9A",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",
		X"AA",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"90",X"99",X"00",X"00",X"39",X"99",X"99",X"00",X"32",X"99",X"22",X"00",X"32",X"22",X"99",
		X"00",X"32",X"62",X"99",X"00",X"92",X"22",X"99",X"00",X"92",X"22",X"66",X"00",X"22",X"29",X"66",
		X"00",X"27",X"29",X"66",X"00",X"26",X"92",X"66",X"00",X"22",X"92",X"66",X"00",X"22",X"96",X"66",
		X"00",X"22",X"96",X"66",X"00",X"22",X"92",X"66",X"00",X"26",X"92",X"66",X"00",X"27",X"29",X"66",
		X"00",X"22",X"29",X"66",X"00",X"92",X"22",X"66",X"00",X"92",X"22",X"99",X"00",X"32",X"62",X"99",
		X"00",X"32",X"22",X"99",X"00",X"32",X"99",X"22",X"00",X"99",X"99",X"99",X"00",X"90",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"99",X"72",X"00",X"00",
		X"92",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"29",X"77",X"00",X"00",X"99",X"22",X"00",X"00",
		X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"29",X"00",X"00",
		X"99",X"29",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",
		X"99",X"22",X"00",X"00",X"29",X"77",X"00",X"00",X"22",X"22",X"00",X"00",X"92",X"22",X"00",X"00",
		X"99",X"72",X"00",X"00",X"22",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"29",X"00",
		X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"62",X"90",X"00",X"92",X"26",X"99",
		X"00",X"22",X"22",X"29",X"00",X"22",X"92",X"92",X"00",X"22",X"92",X"99",X"00",X"72",X"29",X"99",
		X"00",X"22",X"29",X"29",X"00",X"92",X"99",X"66",X"00",X"29",X"96",X"66",X"00",X"22",X"96",X"66",
		X"00",X"22",X"96",X"66",X"00",X"22",X"96",X"66",X"00",X"22",X"92",X"66",X"00",X"22",X"92",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"90",X"00",X"00",X"62",X"99",X"00",X"00",X"69",X"99",X"00",X"00",X"99",X"22",X"00",X"00",
		X"00",X"99",X"92",X"66",X"00",X"99",X"99",X"66",X"00",X"09",X"29",X"66",X"00",X"00",X"22",X"66",
		X"00",X"00",X"92",X"66",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"92",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"26",X"00",X"00",X"99",X"22",X"90",X"00",
		X"99",X"22",X"00",X"00",X"99",X"22",X"90",X"00",X"99",X"22",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"92",X"96",X"00",X"00",X"22",X"96",X"00",X"00",X"22",X"99",X"00",X"00",
		X"22",X"69",X"00",X"00",X"77",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"09",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"9E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"99",X"00",
		X"00",X"99",X"77",X"99",X"00",X"99",X"27",X"99",X"00",X"99",X"77",X"99",X"00",X"99",X"27",X"99",
		X"00",X"99",X"26",X"22",X"00",X"99",X"22",X"22",X"00",X"99",X"26",X"22",X"00",X"99",X"22",X"22",
		X"00",X"E9",X"26",X"92",X"00",X"92",X"72",X"99",X"00",X"E9",X"26",X"92",X"00",X"92",X"72",X"99",
		X"00",X"99",X"29",X"96",X"00",X"09",X"29",X"66",X"00",X"99",X"29",X"96",X"00",X"09",X"29",X"66",
		X"00",X"00",X"29",X"66",X"00",X"00",X"29",X"66",X"00",X"00",X"29",X"66",X"00",X"00",X"29",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"29",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"00",X"00",X"92",X"66",X"00",X"00",X"99",X"66",X"00",X"00",X"92",X"66",X"00",X"00",X"99",X"66",
		X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"96",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"29",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"22",X"00",X"00",X"99",X"92",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"92",X"00",X"00",
		X"92",X"29",X"00",X"00",X"22",X"92",X"00",X"00",X"92",X"29",X"00",X"00",X"22",X"92",X"00",X"00",
		X"22",X"99",X"00",X"00",X"62",X"00",X"00",X"00",X"22",X"99",X"00",X"00",X"62",X"00",X"00",X"00",
		X"22",X"99",X"00",X"00",X"72",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"72",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"E9",X"00",X"00",X"99",X"E9",X"00",X"00",X"09",X"E9",X"00",X"00",X"99",X"E9",
		X"00",X"00",X"22",X"29",X"00",X"00",X"22",X"62",X"00",X"00",X"22",X"29",X"00",X"00",X"22",X"62",
		X"00",X"09",X"22",X"26",X"00",X"99",X"62",X"26",X"00",X"09",X"22",X"26",X"00",X"99",X"62",X"26",
		X"00",X"00",X"27",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"27",X"22",X"00",X"00",X"22",X"22",
		X"00",X"00",X"22",X"92",X"00",X"00",X"62",X"00",X"00",X"00",X"22",X"92",X"00",X"00",X"62",X"99",
		X"00",X"00",X"29",X"99",X"00",X"00",X"92",X"99",X"00",X"00",X"29",X"99",X"00",X"00",X"92",X"99",
		X"00",X"00",X"29",X"66",X"00",X"00",X"29",X"66",X"00",X"00",X"29",X"66",X"00",X"00",X"29",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",
		X"00",X"00",X"92",X"66",X"00",X"00",X"92",X"66",X"00",X"00",X"92",X"66",X"00",X"00",X"09",X"66",
		X"00",X"00",X"09",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"72",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"29",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"92",X"00",X"00",X"00",
		X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",
		X"92",X"00",X"00",X"00",X"22",X"09",X"00",X"00",X"92",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"66",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"39",X"00",X"00",X"99",X"00",X"00",X"99",X"92",X"39",X"00",
		X"9E",X"22",X"EE",X"00",X"09",X"22",X"97",X"00",X"99",X"22",X"93",X"00",X"09",X"22",X"97",X"00",
		X"09",X"22",X"27",X"00",X"09",X"62",X"62",X"00",X"09",X"62",X"62",X"00",X"09",X"62",X"62",X"00",
		X"97",X"62",X"67",X"00",X"99",X"62",X"69",X"00",X"99",X"62",X"67",X"00",X"99",X"22",X"67",X"00",
		X"99",X"99",X"67",X"00",X"99",X"66",X"67",X"00",X"99",X"99",X"67",X"00",X"99",X"99",X"27",X"00",
		X"07",X"99",X"77",X"00",X"07",X"99",X"92",X"00",X"07",X"99",X"72",X"00",X"09",X"66",X"92",X"00",
		X"09",X"66",X"92",X"00",X"09",X"66",X"92",X"00",X"09",X"66",X"92",X"00",X"09",X"66",X"92",X"00",
		X"09",X"66",X"92",X"00",X"09",X"66",X"92",X"00",X"09",X"66",X"92",X"00",X"09",X"66",X"92",X"00",
		X"09",X"66",X"92",X"00",X"09",X"66",X"92",X"00",X"09",X"99",X"92",X"00",X"07",X"99",X"92",X"00",
		X"07",X"99",X"97",X"00",X"07",X"99",X"92",X"00",X"07",X"99",X"97",X"00",X"97",X"99",X"27",X"00",
		X"97",X"99",X"27",X"00",X"97",X"22",X"27",X"00",X"97",X"99",X"27",X"00",X"97",X"22",X"27",X"00",
		X"97",X"22",X"27",X"00",X"97",X"29",X"27",X"00",X"99",X"22",X"27",X"00",X"99",X"29",X"27",X"00",
		X"09",X"99",X"27",X"00",X"09",X"77",X"90",X"00",X"09",X"77",X"00",X"00",X"09",X"77",X"99",X"00",
		X"09",X"00",X"00",X"00",X"09",X"99",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"50",X"00",X"00",X"D9",X"00",X"00",X"00",X"99",X"50",X"00",
		X"00",X"99",X"55",X"00",X"00",X"95",X"90",X"00",X"00",X"50",X"95",X"00",X"00",X"05",X"90",X"00",
		X"00",X"90",X"95",X"00",X"00",X"00",X"90",X"00",X"00",X"90",X"95",X"00",X"00",X"99",X"50",X"00",
		X"00",X"99",X"05",X"00",X"00",X"99",X"50",X"00",X"00",X"99",X"05",X"00",X"00",X"99",X"50",X"00",
		X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0B",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"0B",X"00",X"00",
		X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"B0",X"99",X"B0",X"00",X"00",X"99",X"00",X"00",X"0B",X"9D",X"00",X"00",
		X"B0",X"99",X"00",X"00",X"00",X"99",X"B0",X"00",X"B0",X"95",X"00",X"00",X"00",X"59",X"B0",X"00",
		X"00",X"59",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"BB",X"00",X"09",X"99",X"00",X"00",
		X"09",X"99",X"55",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"B0",X"00",X"00",X"00",
		X"00",X"B0",X"00",X"00",X"00",X"BB",X"50",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"B0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"99",X"72",X"00",X"00",
		X"92",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"29",X"22",X"00",X"00",X"99",X"22",X"00",X"00",
		X"99",X"29",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"29",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"29",X"00",X"00",X"92",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"92",X"22",X"00",X"00",
		X"29",X"72",X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"69",X"90",X"00",X"00",X"62",X"99",X"00",X"00",X"69",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"92",X"00",X"00",X"99",X"22",X"99",X"00",X"99",X"22",X"90",X"00",X"99",X"22",X"99",X"00",
		X"99",X"22",X"90",X"00",X"99",X"22",X"90",X"00",X"99",X"22",X"90",X"00",X"99",X"77",X"00",X"00",
		X"99",X"99",X"00",X"00",X"92",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"99",X"00",X"00",
		X"99",X"09",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"09",X"00",X"00",X"99",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"90",X"00",X"00",X"69",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"29",X"00",X"00",X"99",X"92",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"92",X"00",X"00",
		X"99",X"69",X"00",X"00",X"22",X"72",X"00",X"00",X"92",X"29",X"00",X"00",X"22",X"72",X"00",X"00",
		X"29",X"77",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"99",X"00",X"00",
		X"29",X"00",X"00",X"00",X"97",X"99",X"00",X"00",X"92",X"00",X"00",X"00",X"72",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"29",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"92",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"92",X"66",X"00",X"00",X"09",X"66",X"00",X"00",X"92",X"66",X"00",X"00",X"09",X"66",
		X"00",X"00",X"09",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"29",
		X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"66",X"92",X"00",X"09",X"66",X"92",X"00",X"09",X"66",X"92",X"00",X"09",X"66",X"92",X"00",
		X"09",X"99",X"72",X"00",X"09",X"66",X"92",X"00",X"09",X"99",X"92",X"00",X"07",X"99",X"92",X"00",
		X"09",X"99",X"92",X"00",X"09",X"99",X"92",X"00",X"09",X"99",X"97",X"00",X"99",X"99",X"27",X"00",
		X"97",X"99",X"29",X"00",X"99",X"22",X"97",X"00",X"97",X"99",X"97",X"00",X"97",X"22",X"97",X"00",
		X"92",X"22",X"97",X"00",X"92",X"77",X"77",X"00",X"92",X"77",X"77",X"00",X"92",X"77",X"77",X"00",
		X"02",X"99",X"00",X"00",X"09",X"99",X"90",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"99",X"00",
		X"09",X"00",X"00",X"00",X"09",X"00",X"99",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"E2",X"99",X"00",X"00",X"99",X"22",X"99",X"00",X"E2",X"99",X"22",X"00",X"E2",X"22",X"99",
		X"00",X"E2",X"62",X"66",X"00",X"22",X"22",X"99",X"00",X"92",X"22",X"66",X"00",X"22",X"29",X"66",
		X"00",X"27",X"92",X"66",X"00",X"26",X"92",X"66",X"00",X"22",X"92",X"66",X"00",X"22",X"96",X"66",
		X"00",X"26",X"92",X"66",X"00",X"22",X"29",X"66",X"00",X"26",X"92",X"66",X"00",X"27",X"29",X"66",
		X"00",X"99",X"29",X"66",X"00",X"99",X"62",X"99",X"00",X"99",X"22",X"99",X"00",X"E9",X"62",X"99",
		X"00",X"EE",X"99",X"99",X"00",X"00",X"99",X"00",X"00",X"99",X"99",X"99",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"26",X"99",X"00",X"99",X"99",X"90",X"00",X"92",X"26",X"99",
		X"00",X"22",X"92",X"99",X"00",X"22",X"92",X"99",X"00",X"22",X"92",X"99",X"00",X"72",X"29",X"99",
		X"00",X"22",X"29",X"29",X"00",X"92",X"96",X"66",X"00",X"99",X"96",X"66",X"00",X"92",X"96",X"66",
		X"00",X"99",X"96",X"66",X"00",X"99",X"92",X"66",X"00",X"99",X"92",X"66",X"00",X"99",X"92",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"E9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"99",X"00",
		X"00",X"99",X"92",X"00",X"00",X"09",X"27",X"99",X"00",X"99",X"77",X"99",X"00",X"09",X"27",X"99",
		X"00",X"99",X"26",X"99",X"00",X"9E",X"22",X"92",X"00",X"99",X"26",X"99",X"00",X"9E",X"22",X"92",
		X"00",X"EE",X"22",X"92",X"00",X"EE",X"22",X"22",X"00",X"EE",X"26",X"92",X"00",X"EE",X"72",X"99",
		X"00",X"99",X"29",X"96",X"00",X"99",X"29",X"99",X"00",X"99",X"29",X"96",X"00",X"09",X"29",X"66",
		X"00",X"00",X"29",X"66",X"00",X"00",X"29",X"66",X"00",X"00",X"29",X"66",X"00",X"00",X"29",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"E9",X"00",X"00",X"99",X"E9",
		X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"69",X"00",X"00",X"22",X"29",X"00",X"00",X"22",X"69",
		X"00",X"00",X"22",X"99",X"00",X"03",X"62",X"29",X"00",X"00",X"22",X"99",X"00",X"03",X"62",X"29",
		X"00",X"03",X"62",X"29",X"00",X"03",X"22",X"22",X"00",X"03",X"27",X"29",X"00",X"03",X"22",X"22",
		X"00",X"00",X"22",X"92",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"92",X"00",X"00",X"62",X"99",
		X"00",X"00",X"29",X"99",X"00",X"00",X"92",X"99",X"00",X"00",X"29",X"99",X"00",X"00",X"92",X"99",
		X"00",X"00",X"29",X"66",X"00",X"00",X"29",X"66",X"00",X"00",X"29",X"66",X"00",X"00",X"29",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"92",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"92",X"99",X"00",
		X"00",X"22",X"EE",X"00",X"00",X"22",X"EE",X"00",X"99",X"22",X"99",X"00",X"09",X"22",X"22",X"00",
		X"09",X"22",X"22",X"00",X"09",X"62",X"99",X"00",X"09",X"62",X"99",X"00",X"09",X"62",X"99",X"00",
		X"97",X"62",X"99",X"00",X"99",X"62",X"99",X"00",X"99",X"62",X"99",X"00",X"99",X"22",X"99",X"00",
		X"99",X"99",X"69",X"00",X"99",X"99",X"27",X"00",X"99",X"99",X"69",X"00",X"99",X"99",X"27",X"00",
		X"99",X"99",X"77",X"00",X"07",X"66",X"72",X"00",X"07",X"99",X"72",X"00",X"09",X"66",X"92",X"00",
		X"09",X"66",X"92",X"00",X"09",X"66",X"92",X"00",X"09",X"66",X"92",X"00",X"09",X"66",X"92",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"32",X"99",X"22",X"00",X"32",X"22",X"99",X"00",X"32",X"99",X"22",X"00",X"32",X"22",X"99",
		X"00",X"92",X"22",X"66",X"00",X"22",X"29",X"66",X"00",X"92",X"22",X"66",X"00",X"22",X"29",X"66",
		X"00",X"22",X"92",X"66",X"00",X"22",X"96",X"66",X"00",X"22",X"92",X"66",X"00",X"22",X"96",X"66",
		X"00",X"26",X"92",X"66",X"00",X"27",X"29",X"66",X"00",X"26",X"92",X"66",X"00",X"27",X"29",X"66",
		X"00",X"99",X"22",X"99",X"00",X"E9",X"62",X"99",X"00",X"99",X"22",X"99",X"00",X"E9",X"62",X"99",
		X"00",X"99",X"99",X"99",X"00",X"00",X"99",X"00",X"00",X"99",X"99",X"99",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"92",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"90",X"00",X"00",
		X"69",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"69",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"90",X"00",X"92",X"26",X"99",X"00",X"99",X"99",X"90",X"00",X"92",X"26",X"99",
		X"00",X"22",X"92",X"99",X"00",X"72",X"29",X"99",X"00",X"22",X"92",X"99",X"00",X"72",X"29",X"99",
		X"00",X"99",X"96",X"66",X"00",X"92",X"96",X"66",X"00",X"99",X"96",X"66",X"00",X"92",X"96",X"66",
		X"00",X"99",X"96",X"66",X"00",X"99",X"96",X"66",X"00",X"99",X"92",X"66",X"00",X"99",X"92",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"9E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"92",X"00",X"00",X"09",X"22",X"00",X"00",X"99",X"77",X"00",X"00",X"09",X"27",X"90",
		X"00",X"99",X"67",X"99",X"00",X"99",X"22",X"99",X"00",X"99",X"26",X"99",X"00",X"9E",X"22",X"92",
		X"00",X"EE",X"22",X"99",X"00",X"EE",X"22",X"22",X"00",X"EE",X"26",X"92",X"00",X"9E",X"72",X"99",
		X"00",X"9E",X"72",X"99",X"00",X"99",X"29",X"99",X"00",X"99",X"29",X"96",X"00",X"09",X"29",X"66",
		X"00",X"09",X"29",X"66",X"00",X"00",X"29",X"66",X"00",X"00",X"29",X"66",X"00",X"00",X"29",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"E9",X"00",X"00",X"99",X"E9",
		X"00",X"00",X"99",X"99",X"00",X"00",X"22",X"29",X"00",X"00",X"22",X"29",X"00",X"00",X"22",X"69",
		X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"62",X"29",
		X"00",X"00",X"62",X"26",X"00",X"00",X"72",X"22",X"00",X"00",X"27",X"29",X"00",X"00",X"22",X"22",
		X"00",X"00",X"22",X"99",X"00",X"09",X"22",X"22",X"00",X"09",X"22",X"92",X"00",X"09",X"62",X"99",
		X"00",X"00",X"69",X"99",X"00",X"00",X"69",X"99",X"00",X"00",X"29",X"99",X"00",X"00",X"92",X"99",
		X"00",X"00",X"92",X"66",X"00",X"00",X"92",X"66",X"00",X"00",X"29",X"66",X"00",X"00",X"29",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"92",X"99",X"00",
		X"00",X"22",X"EE",X"00",X"03",X"22",X"EE",X"00",X"99",X"22",X"99",X"00",X"09",X"22",X"22",X"00",
		X"09",X"22",X"22",X"00",X"09",X"62",X"99",X"00",X"09",X"62",X"99",X"00",X"09",X"62",X"99",X"00",
		X"97",X"62",X"99",X"00",X"99",X"62",X"99",X"00",X"99",X"62",X"99",X"00",X"99",X"22",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"66",X"99",X"00",X"99",X"99",X"69",X"00",X"99",X"99",X"27",X"00",
		X"99",X"99",X"77",X"00",X"07",X"99",X"72",X"00",X"07",X"99",X"72",X"00",X"09",X"66",X"92",X"00",
		X"09",X"66",X"92",X"00",X"09",X"66",X"92",X"00",X"09",X"66",X"92",X"00",X"09",X"66",X"92",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"99",X"72",X"00",X"00",
		X"92",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"29",X"22",X"00",X"00",X"99",X"22",X"00",X"00",
		X"99",X"22",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"29",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"29",X"00",X"00",X"29",X"27",X"00",X"00",X"22",X"22",X"00",X"00",X"92",X"22",X"00",X"00",
		X"29",X"72",X"00",X"00",X"99",X"92",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"92",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"22",X"90",X"00",X"99",X"22",X"99",X"00",
		X"99",X"22",X"90",X"00",X"99",X"22",X"90",X"00",X"99",X"22",X"90",X"00",X"99",X"77",X"00",X"00",
		X"99",X"99",X"00",X"00",X"92",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"99",X"00",X"00",
		X"92",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"09",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"92",X"66",X"00",X"99",X"99",X"66",X"00",X"09",X"29",X"66",X"00",X"09",X"22",X"66",
		X"00",X"00",X"92",X"96",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"69",X"00",X"00",X"00",X"69",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"92",X"00",X"00",
		X"99",X"69",X"00",X"00",X"99",X"22",X"00",X"00",X"92",X"29",X"00",X"00",X"22",X"72",X"00",X"00",
		X"29",X"77",X"00",X"00",X"92",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"99",X"00",X"00",
		X"29",X"99",X"00",X"00",X"97",X"99",X"00",X"00",X"92",X"00",X"00",X"00",X"72",X"00",X"00",X"00",
		X"79",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"29",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"92",X"00",X"00",X"00",
		X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",
		X"29",X"90",X"00",X"00",X"92",X"90",X"00",X"00",X"22",X"90",X"00",X"00",X"22",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"92",X"66",X"00",X"00",X"92",X"66",X"00",X"00",X"92",X"66",X"00",X"00",X"09",X"66",
		X"00",X"00",X"09",X"66",X"00",X"00",X"09",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",
		X"00",X"00",X"00",X"67",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"29",
		X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"66",X"92",X"00",X"09",X"66",X"92",X"00",X"09",X"66",X"92",X"00",X"09",X"66",X"92",X"00",
		X"09",X"66",X"72",X"00",X"09",X"66",X"92",X"00",X"09",X"99",X"92",X"00",X"07",X"99",X"92",X"00",
		X"09",X"99",X"92",X"00",X"09",X"99",X"92",X"00",X"09",X"99",X"97",X"00",X"09",X"99",X"27",X"00",
		X"09",X"99",X"29",X"00",X"09",X"22",X"99",X"00",X"07",X"99",X"97",X"00",X"07",X"22",X"97",X"00",
		X"02",X"22",X"97",X"00",X"02",X"22",X"97",X"00",X"02",X"77",X"77",X"00",X"02",X"77",X"77",X"00",
		X"02",X"99",X"27",X"00",X"00",X"99",X"90",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"99",X"00",
		X"09",X"99",X"99",X"00",X"00",X"00",X"99",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"26",X"00",X"00",X"00",
		X"26",X"99",X"00",X"00",X"26",X"99",X"00",X"00",X"26",X"00",X"00",X"00",X"26",X"00",X"00",X"00",
		X"26",X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"22",X"00",X"00",X"00",
		X"29",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"90",X"00",X"02",X"00",X"90",X"00",X"26",X"26",X"00",X"00",X"62",X"22",X"00",
		X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"20",X"00",X"00",X"22",X"00",X"00",
		X"00",X"22",X"00",X"00",X"00",X"22",X"09",X"00",X"00",X"26",X"99",X"00",X"00",X"22",X"90",X"00",
		X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"00",X"00",X"22",X"22",X"00",
		X"22",X"22",X"00",X"00",X"22",X"22",X"99",X"00",X"92",X"22",X"99",X"00",X"09",X"22",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"99",X"00",X"00",X"99",X"99",X"99",X"00",X"EE",X"11",X"55",X"00",X"EE",X"44",X"55",
		X"00",X"EE",X"44",X"59",X"00",X"55",X"59",X"59",X"00",X"55",X"11",X"55",X"00",X"55",X"44",X"14",
		X"00",X"51",X"44",X"14",X"00",X"51",X"44",X"44",X"00",X"51",X"44",X"44",X"00",X"51",X"11",X"44",
		X"00",X"91",X"59",X"14",X"00",X"51",X"44",X"44",X"00",X"91",X"41",X"14",X"00",X"55",X"44",X"44",
		X"00",X"55",X"11",X"14",X"00",X"59",X"11",X"14",X"00",X"EE",X"55",X"59",X"00",X"EE",X"99",X"59",
		X"00",X"EE",X"11",X"59",X"00",X"95",X"11",X"55",X"00",X"99",X"99",X"99",X"00",X"09",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"55",X"11",X"00",X"00",X"15",X"59",X"00",X"00",
		X"91",X"99",X"00",X"00",X"55",X"99",X"00",X"00",X"49",X"59",X"00",X"00",X"11",X"44",X"00",X"00",
		X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",
		X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",
		X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"49",X"99",X"00",X"00",X"55",X"99",X"00",X"00",
		X"94",X"99",X"00",X"00",X"59",X"55",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"11",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"54",X"90",X"00",X"00",X"59",X"19",X"00",X"09",X"11",X"11",
		X"00",X"09",X"44",X"55",X"00",X"09",X"44",X"99",X"00",X"95",X"14",X"19",X"00",X"91",X"44",X"59",
		X"00",X"94",X"51",X"91",X"00",X"94",X"59",X"54",X"00",X"95",X"45",X"44",X"00",X"55",X"44",X"14",
		X"00",X"E3",X"44",X"44",X"00",X"E3",X"44",X"44",X"00",X"E3",X"44",X"44",X"00",X"95",X"51",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"51",X"00",X"00",X"00",
		X"91",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"55",X"00",X"00",X"11",X"54",X"00",X"00",
		X"44",X"15",X"90",X"00",X"44",X"94",X"90",X"00",X"44",X"99",X"90",X"00",X"44",X"41",X"00",X"00",
		X"00",X"95",X"95",X"44",X"00",X"99",X"19",X"44",X"00",X"00",X"14",X"44",X"00",X"00",X"51",X"54",
		X"00",X"00",X"95",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"55",
		X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"49",X"00",X"00",X"44",X"49",X"00",X"00",
		X"44",X"45",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"54",X"59",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"95",X"00",X"00",X"59",X"99",X"00",X"00",X"55",X"59",X"00",X"00",
		X"51",X"95",X"00",X"00",X"59",X"95",X"00",X"00",X"99",X"55",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"59",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E3",X"00",
		X"00",X"00",X"33",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"55",X"90",X"00",X"00",X"11",X"99",
		X"00",X"00",X"14",X"59",X"00",X"09",X"94",X"15",X"00",X"99",X"11",X"41",X"00",X"99",X"44",X"41",
		X"00",X"9E",X"94",X"91",X"00",X"EE",X"55",X"95",X"00",X"E3",X"49",X"91",X"00",X"33",X"41",X"91",
		X"00",X"51",X"44",X"91",X"00",X"91",X"44",X"91",X"00",X"95",X"44",X"51",X"00",X"09",X"44",X"14",
		X"00",X"09",X"15",X"14",X"00",X"00",X"59",X"14",X"00",X"00",X"99",X"44",X"00",X"00",X"55",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"19",X"00",X"00",X"00",
		X"51",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"14",X"00",X"00",X"00",
		X"00",X"00",X"54",X"44",X"00",X"00",X"55",X"44",X"00",X"00",X"51",X"44",X"00",X"00",X"55",X"44",
		X"00",X"00",X"91",X"44",X"00",X"00",X"09",X"44",X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"94",
		X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"45",
		X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"59",X"00",X"00",X"00",X"45",X"90",X"00",X"00",X"14",X"90",X"00",X"00",X"44",X"99",X"00",X"00",
		X"44",X"59",X"00",X"00",X"44",X"15",X"00",X"00",X"44",X"54",X"00",X"00",X"44",X"95",X"00",X"00",
		X"44",X"41",X"00",X"00",X"44",X"55",X"00",X"00",X"44",X"95",X"00",X"00",X"44",X"94",X"00",X"00",
		X"44",X"15",X"00",X"00",X"44",X"55",X"00",X"00",X"44",X"55",X"00",X"00",X"44",X"99",X"00",X"00",
		X"44",X"00",X"00",X"00",X"49",X"00",X"00",X"00",X"45",X"00",X"00",X"00",X"19",X"00",X"00",X"00",
		X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"19",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"55",X"00",X"00",X"99",X"95",X"00",X"00",X"99",X"19",
		X"00",X"00",X"54",X"15",X"00",X"00",X"95",X"11",X"00",X"00",X"95",X"41",X"00",X"00",X"95",X"44",
		X"00",X"00",X"95",X"14",X"00",X"00",X"55",X"44",X"00",X"00",X"55",X"44",X"00",X"00",X"15",X"41",
		X"00",X"00",X"49",X"44",X"00",X"00",X"49",X"14",X"00",X"00",X"45",X"59",X"00",X"00",X"11",X"99",
		X"00",X"00",X"14",X"99",X"00",X"00",X"54",X"99",X"00",X"00",X"94",X"99",X"00",X"00",X"91",X"51",
		X"00",X"00",X"91",X"14",X"00",X"00",X"95",X"44",X"00",X"00",X"09",X"44",X"00",X"00",X"09",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"19",X"00",X"00",X"00",
		X"19",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"91",X"00",X"00",X"00",
		X"95",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"00",X"00",X"09",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",
		X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"14",
		X"00",X"00",X"00",X"94",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"59",
		X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"55",
		X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"95",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"41",X"00",X"00",X"00",X"45",X"00",X"00",X"00",
		X"45",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"44",X"90",X"00",X"00",X"44",X"90",X"00",X"00",X"44",X"90",X"00",X"00",
		X"44",X"90",X"00",X"00",X"44",X"90",X"00",X"00",X"44",X"19",X"00",X"00",X"49",X"45",X"00",X"00",
		X"99",X"15",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"00",X"00",X"00",X"59",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"59",X"99",X"99",X"00",X"95",X"15",X"E5",X"00",X"59",X"99",X"E9",X"00",
		X"59",X"19",X"35",X"00",X"95",X"59",X"15",X"00",X"09",X"59",X"19",X"00",X"99",X"49",X"19",X"00",
		X"99",X"49",X"49",X"00",X"99",X"49",X"49",X"00",X"99",X"49",X"49",X"00",X"99",X"49",X"19",X"00",
		X"99",X"49",X"49",X"00",X"99",X"49",X"19",X"00",X"99",X"11",X"19",X"00",X"09",X"99",X"19",X"00",
		X"09",X"99",X"49",X"00",X"09",X"99",X"59",X"00",X"09",X"99",X"19",X"00",X"09",X"99",X"59",X"00",
		X"09",X"11",X"19",X"00",X"09",X"44",X"59",X"00",X"09",X"44",X"19",X"00",X"09",X"44",X"59",X"00",
		X"09",X"44",X"19",X"00",X"09",X"44",X"59",X"00",X"09",X"44",X"19",X"00",X"09",X"44",X"59",X"00",
		X"09",X"44",X"19",X"00",X"09",X"44",X"59",X"00",X"09",X"44",X"19",X"00",X"09",X"44",X"19",X"00",
		X"09",X"44",X"59",X"00",X"99",X"44",X"19",X"00",X"99",X"44",X"19",X"00",X"99",X"44",X"59",X"00",
		X"99",X"44",X"19",X"00",X"99",X"44",X"59",X"00",X"99",X"44",X"19",X"00",X"99",X"44",X"59",X"00",
		X"99",X"44",X"19",X"00",X"99",X"11",X"59",X"00",X"99",X"99",X"19",X"00",X"09",X"99",X"59",X"00",
		X"95",X"55",X"19",X"00",X"91",X"15",X"41",X"00",X"95",X"99",X"91",X"00",X"91",X"55",X"51",X"00",
		X"99",X"99",X"99",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"9A",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"39",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"33",X"00",X"00",
		X"99",X"39",X"00",X"00",X"99",X"93",X"00",X"00",X"90",X"93",X"00",X"00",X"90",X"99",X"00",X"00",
		X"90",X"93",X"00",X"00",X"90",X"99",X"00",X"00",X"90",X"93",X"00",X"00",X"99",X"93",X"00",X"00",
		X"99",X"93",X"00",X"00",X"99",X"39",X"00",X"00",X"39",X"93",X"00",X"00",X"93",X"39",X"50",X"00",
		X"99",X"99",X"05",X"00",X"99",X"99",X"50",X"00",X"99",X"99",X"05",X"00",X"99",X"90",X"50",X"00",
		X"99",X"05",X"05",X"00",X"09",X"50",X"50",X"00",X"00",X"05",X"05",X"00",X"00",X"50",X"50",X"00",
		X"00",X"05",X"05",X"00",X"00",X"00",X"50",X"00",X"00",X"05",X"05",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"39",X"00",X"00",
		X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"93",X"99",X"00",X"00",X"93",X"99",X"00",X"00",
		X"99",X"D9",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"05",X"00",X"99",X"00",X"50",X"00",
		X"99",X"00",X"05",X"00",X"99",X"00",X"50",X"00",X"99",X"00",X"05",X"00",X"99",X"00",X"50",X"00",
		X"99",X"00",X"05",X"00",X"09",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"55",X"11",X"00",X"00",X"15",X"59",X"00",X"00",
		X"91",X"55",X"00",X"00",X"55",X"51",X"00",X"00",X"49",X"59",X"00",X"00",X"11",X"99",X"00",X"00",
		X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",
		X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",
		X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"49",X"19",X"00",X"00",X"55",X"14",X"00",X"00",
		X"94",X"54",X"00",X"00",X"51",X"51",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"51",X"90",X"00",X"00",
		X"91",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"55",X"00",X"00",X"11",X"54",X"00",X"00",
		X"44",X"15",X"90",X"00",X"44",X"94",X"90",X"00",X"44",X"14",X"90",X"00",X"44",X"59",X"00",X"00",
		X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",
		X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"54",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"59",X"95",X"00",X"00",X"55",X"59",X"00",X"00",
		X"51",X"95",X"00",X"00",X"59",X"95",X"00",X"00",X"99",X"55",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"59",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"59",X"90",X"00",X"00",X"45",X"99",X"00",X"00",X"14",X"99",X"00",X"00",X"44",X"99",X"00",X"00",
		X"44",X"59",X"00",X"00",X"44",X"15",X"00",X"00",X"44",X"54",X"00",X"00",X"54",X"15",X"00",X"00",
		X"45",X"59",X"00",X"00",X"99",X"55",X"00",X"00",X"99",X"95",X"00",X"00",X"99",X"54",X"00",X"00",
		X"99",X"15",X"00",X"00",X"95",X"55",X"00",X"00",X"55",X"55",X"00",X"00",X"55",X"99",X"00",X"00",
		X"95",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"19",X"00",X"00",X"00",
		X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"19",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"41",X"00",X"00",X"00",X"45",X"00",X"00",X"00",
		X"45",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"90",X"00",X"00",X"44",X"90",X"00",X"00",
		X"44",X"90",X"00",X"00",X"44",X"90",X"00",X"00",X"45",X"90",X"00",X"00",X"55",X"90",X"00",X"00",
		X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"19",X"00",X"00",X"99",X"45",X"00",X"00",
		X"99",X"15",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"59",X"00",X"00",X"00",
		X"91",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",
		X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"14",
		X"00",X"00",X"00",X"94",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"59",
		X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"55",
		X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"95",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"44",X"19",X"00",X"09",X"44",X"59",X"00",X"09",X"44",X"19",X"00",X"09",X"44",X"59",X"00",
		X"09",X"44",X"19",X"00",X"09",X"44",X"59",X"00",X"09",X"44",X"19",X"00",X"09",X"44",X"19",X"00",
		X"09",X"44",X"59",X"00",X"59",X"44",X"19",X"00",X"59",X"44",X"19",X"00",X"59",X"54",X"59",X"00",
		X"59",X"45",X"19",X"00",X"59",X"99",X"59",X"00",X"59",X"99",X"19",X"00",X"59",X"99",X"59",X"00",
		X"59",X"99",X"19",X"00",X"59",X"99",X"59",X"00",X"59",X"99",X"19",X"00",X"09",X"99",X"59",X"00",
		X"95",X"99",X"19",X"00",X"91",X"55",X"41",X"00",X"95",X"99",X"91",X"00",X"91",X"55",X"51",X"00",
		X"99",X"99",X"99",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"99",X"00",X"00",X"99",X"99",X"99",X"00",X"9E",X"11",X"55",X"00",X"9E",X"44",X"15",
		X"00",X"9E",X"44",X"59",X"00",X"55",X"55",X"59",X"00",X"55",X"55",X"55",X"00",X"99",X"99",X"14",
		X"00",X"99",X"D9",X"14",X"00",X"DD",X"D9",X"44",X"00",X"DD",X"9D",X"44",X"00",X"DD",X"DD",X"44",
		X"00",X"DD",X"DD",X"14",X"00",X"DD",X"9D",X"44",X"00",X"DD",X"D9",X"14",X"00",X"99",X"D9",X"44",
		X"00",X"99",X"99",X"14",X"00",X"59",X"99",X"14",X"00",X"9E",X"55",X"59",X"00",X"9E",X"99",X"59",
		X"00",X"5E",X"11",X"59",X"00",X"95",X"11",X"11",X"00",X"99",X"99",X"99",X"00",X"09",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"15",X"90",X"00",X"00",X"11",X"90",
		X"00",X"00",X"44",X"99",X"00",X"00",X"54",X"99",X"00",X"00",X"55",X"19",X"00",X"09",X"99",X"11",
		X"00",X"09",X"99",X"55",X"00",X"09",X"DD",X"99",X"00",X"95",X"9D",X"19",X"00",X"91",X"99",X"59",
		X"00",X"94",X"9D",X"91",X"00",X"94",X"D9",X"54",X"00",X"95",X"99",X"44",X"00",X"EE",X"D9",X"14",
		X"00",X"EE",X"D9",X"44",X"00",X"E3",X"95",X"44",X"00",X"E3",X"51",X"44",X"00",X"95",X"51",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"3E",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"E3",X"90",X"00",X"00",X"55",X"99",X"00",X"00",X"95",X"99",X"00",X"00",X"99",X"99",
		X"00",X"00",X"D9",X"59",X"00",X"09",X"DD",X"15",X"00",X"99",X"9D",X"41",X"00",X"99",X"D9",X"41",
		X"00",X"95",X"99",X"51",X"00",X"EE",X"99",X"95",X"00",X"E3",X"D9",X"91",X"00",X"33",X"99",X"91",
		X"00",X"51",X"D9",X"91",X"00",X"91",X"95",X"91",X"00",X"95",X"91",X"51",X"00",X"09",X"11",X"14",
		X"00",X"09",X"15",X"14",X"00",X"00",X"59",X"14",X"00",X"00",X"99",X"44",X"00",X"00",X"55",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"19",X"00",X"00",X"00",
		X"19",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"91",X"00",X"00",X"00",
		X"95",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E3",X"00",X"00",X"99",X"35",X"00",X"00",X"99",X"95",
		X"00",X"00",X"54",X"D9",X"00",X"00",X"95",X"D9",X"00",X"00",X"95",X"DD",X"00",X"00",X"95",X"9D",
		X"00",X"00",X"95",X"9D",X"00",X"00",X"55",X"99",X"00",X"00",X"55",X"D9",X"00",X"00",X"15",X"99",
		X"00",X"00",X"49",X"94",X"00",X"00",X"49",X"14",X"00",X"00",X"45",X"59",X"00",X"00",X"11",X"99",
		X"00",X"00",X"14",X"99",X"00",X"00",X"54",X"99",X"00",X"00",X"94",X"99",X"00",X"00",X"91",X"51",
		X"00",X"00",X"91",X"14",X"00",X"00",X"95",X"44",X"00",X"00",X"09",X"44",X"00",X"00",X"09",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"59",X"99",X"99",X"00",X"95",X"D5",X"E5",X"00",X"59",X"DD",X"E9",X"00",
		X"53",X"99",X"33",X"00",X"95",X"99",X"15",X"00",X"09",X"DD",X"19",X"00",X"09",X"D9",X"19",X"00",
		X"09",X"99",X"49",X"00",X"99",X"99",X"49",X"00",X"09",X"D9",X"49",X"00",X"09",X"99",X"19",X"00",
		X"99",X"99",X"49",X"00",X"09",X"99",X"19",X"00",X"09",X"11",X"19",X"00",X"09",X"99",X"19",X"00",
		X"09",X"99",X"49",X"00",X"09",X"99",X"59",X"00",X"09",X"99",X"19",X"00",X"09",X"99",X"59",X"00",
		X"09",X"11",X"19",X"00",X"09",X"44",X"59",X"00",X"09",X"44",X"19",X"00",X"09",X"44",X"59",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"99",X"00",X"00",X"99",X"99",X"99",X"00",X"EE",X"11",X"55",X"00",X"EE",X"44",X"15",
		X"00",X"EE",X"44",X"59",X"00",X"55",X"55",X"59",X"00",X"55",X"55",X"55",X"00",X"99",X"99",X"14",
		X"00",X"99",X"D9",X"14",X"00",X"DD",X"D9",X"44",X"00",X"DD",X"9D",X"44",X"00",X"DD",X"DD",X"44",
		X"00",X"DD",X"DD",X"14",X"00",X"DD",X"9D",X"44",X"00",X"DD",X"D9",X"14",X"00",X"99",X"D9",X"44",
		X"00",X"99",X"99",X"14",X"00",X"59",X"99",X"14",X"00",X"EE",X"55",X"59",X"00",X"EE",X"99",X"59",
		X"00",X"EE",X"11",X"59",X"00",X"95",X"11",X"11",X"00",X"99",X"99",X"99",X"00",X"09",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"51",X"00",X"00",X"00",
		X"91",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"55",X"00",X"00",X"11",X"54",X"00",X"00",
		X"44",X"15",X"90",X"00",X"44",X"94",X"90",X"00",X"44",X"14",X"90",X"00",X"44",X"59",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"11",X"00",
		X"00",X"00",X"44",X"90",X"00",X"00",X"54",X"99",X"00",X"00",X"55",X"19",X"00",X"09",X"99",X"11",
		X"00",X"09",X"99",X"55",X"00",X"09",X"DD",X"99",X"00",X"95",X"9D",X"19",X"00",X"91",X"99",X"59",
		X"00",X"94",X"9D",X"91",X"00",X"94",X"D9",X"54",X"00",X"95",X"99",X"44",X"00",X"5E",X"D9",X"14",
		X"00",X"EE",X"D9",X"44",X"00",X"E3",X"95",X"44",X"00",X"93",X"51",X"44",X"00",X"95",X"51",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"3E",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"E3",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"95",X"90",X"00",X"00",X"99",X"90",
		X"00",X"00",X"D9",X"59",X"00",X"09",X"DD",X"15",X"00",X"99",X"9D",X"41",X"00",X"99",X"D9",X"41",
		X"00",X"95",X"99",X"51",X"00",X"EE",X"99",X"95",X"00",X"E3",X"D9",X"91",X"00",X"33",X"99",X"91",
		X"00",X"51",X"D9",X"91",X"00",X"91",X"95",X"91",X"00",X"95",X"91",X"51",X"00",X"09",X"11",X"14",
		X"00",X"99",X"15",X"14",X"00",X"99",X"59",X"14",X"00",X"09",X"99",X"44",X"00",X"00",X"55",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"19",X"00",X"00",X"00",
		X"19",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"91",X"00",X"00",X"00",
		X"95",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"5E",
		X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E3",X"00",X"00",X"99",X"35",X"00",X"00",X"99",X"95",
		X"00",X"00",X"54",X"D9",X"00",X"00",X"95",X"D9",X"00",X"00",X"95",X"DD",X"00",X"00",X"95",X"9D",
		X"00",X"00",X"95",X"9D",X"00",X"00",X"55",X"99",X"00",X"00",X"55",X"D9",X"00",X"00",X"15",X"99",
		X"00",X"00",X"49",X"94",X"00",X"00",X"49",X"14",X"00",X"00",X"45",X"59",X"00",X"00",X"11",X"99",
		X"00",X"00",X"14",X"99",X"00",X"00",X"54",X"99",X"00",X"00",X"94",X"99",X"00",X"00",X"91",X"51",
		X"00",X"00",X"91",X"14",X"00",X"00",X"95",X"44",X"00",X"00",X"99",X"44",X"00",X"00",X"09",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"59",X"99",X"99",X"00",X"95",X"D5",X"E5",X"00",X"59",X"DD",X"E9",X"00",
		X"59",X"99",X"15",X"00",X"95",X"99",X"35",X"00",X"09",X"DD",X"19",X"00",X"99",X"D9",X"19",X"00",
		X"99",X"99",X"49",X"00",X"99",X"99",X"49",X"00",X"99",X"D9",X"49",X"00",X"99",X"99",X"19",X"00",
		X"99",X"99",X"49",X"00",X"99",X"99",X"19",X"00",X"99",X"11",X"19",X"00",X"09",X"99",X"19",X"00",
		X"09",X"99",X"49",X"00",X"09",X"99",X"59",X"00",X"09",X"99",X"19",X"00",X"09",X"99",X"59",X"00",
		X"09",X"11",X"19",X"00",X"09",X"44",X"59",X"00",X"09",X"44",X"19",X"00",X"09",X"44",X"59",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"55",X"11",X"00",X"00",X"15",X"59",X"00",X"00",
		X"91",X"55",X"00",X"00",X"55",X"51",X"00",X"00",X"49",X"59",X"00",X"00",X"11",X"99",X"00",X"00",
		X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",
		X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",
		X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"49",X"19",X"00",X"00",X"55",X"14",X"00",X"00",
		X"94",X"54",X"00",X"00",X"51",X"51",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",
		X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"54",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"59",X"95",X"00",X"00",X"55",X"59",X"00",X"00",
		X"51",X"95",X"00",X"00",X"59",X"95",X"00",X"00",X"99",X"55",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"59",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"95",X"95",X"44",X"00",X"99",X"19",X"44",X"00",X"99",X"14",X"44",X"00",X"99",X"51",X"54",
		X"00",X"00",X"95",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"55",
		X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"59",X"00",X"00",X"00",X"45",X"00",X"00",X"00",X"14",X"90",X"00",X"00",X"44",X"99",X"00",X"00",
		X"44",X"59",X"00",X"00",X"44",X"15",X"00",X"00",X"44",X"54",X"00",X"00",X"54",X"15",X"00",X"00",
		X"45",X"59",X"00",X"00",X"99",X"55",X"00",X"00",X"99",X"95",X"00",X"00",X"99",X"54",X"00",X"00",
		X"99",X"15",X"00",X"00",X"95",X"55",X"00",X"00",X"55",X"55",X"00",X"00",X"55",X"99",X"00",X"00",
		X"95",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"19",X"00",X"00",X"00",
		X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"19",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"41",X"00",X"00",X"00",X"45",X"00",X"00",X"00",
		X"45",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"45",X"90",X"00",X"00",X"55",X"90",X"00",X"00",
		X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"19",X"00",X"00",X"99",X"45",X"00",X"00",
		X"99",X"15",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"59",X"00",X"00",X"00",
		X"91",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",
		X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"14",
		X"00",X"00",X"00",X"94",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"59",
		X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"55",
		X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"95",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"44",X"19",X"00",X"09",X"44",X"59",X"00",X"09",X"44",X"19",X"00",X"09",X"44",X"59",X"00",
		X"09",X"44",X"19",X"00",X"09",X"44",X"59",X"00",X"09",X"44",X"19",X"00",X"09",X"44",X"19",X"00",
		X"09",X"44",X"59",X"00",X"59",X"44",X"19",X"00",X"99",X"44",X"19",X"00",X"99",X"54",X"59",X"00",
		X"99",X"45",X"19",X"00",X"99",X"99",X"59",X"00",X"99",X"99",X"19",X"00",X"99",X"99",X"59",X"00",
		X"99",X"99",X"19",X"00",X"99",X"99",X"59",X"00",X"99",X"99",X"19",X"00",X"09",X"99",X"59",X"00",
		X"95",X"99",X"19",X"00",X"91",X"55",X"41",X"00",X"95",X"99",X"91",X"00",X"91",X"55",X"51",X"00",
		X"99",X"99",X"99",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"99",X"99",X"00",X"22",X"92",X"92",X"00",X"29",X"29",X"29",X"00",X"29",X"29",X"29",X"00",
		X"29",X"29",X"29",X"00",X"99",X"29",X"29",X"00",X"22",X"29",X"29",X"00",X"22",X"29",X"29",X"00",
		X"99",X"29",X"29",X"00",X"00",X"29",X"29",X"00",X"00",X"29",X"29",X"00",X"99",X"29",X"29",X"00",
		X"29",X"29",X"29",X"00",X"29",X"29",X"29",X"00",X"29",X"29",X"29",X"00",X"92",X"92",X"92",X"00",
		X"99",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"09",X"09",X"09",X"00",X"99",X"99",X"99",X"90",X"92",X"92",X"92",X"90",
		X"92",X"92",X"92",X"90",X"92",X"92",X"92",X"90",X"92",X"92",X"92",X"90",X"92",X"92",X"92",X"90",
		X"92",X"92",X"92",X"90",X"92",X"92",X"92",X"90",X"92",X"92",X"92",X"90",X"92",X"92",X"92",X"90",
		X"92",X"92",X"92",X"90",X"92",X"92",X"92",X"90",X"99",X"99",X"99",X"90",X"09",X"09",X"09",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"29",X"90",X"90",X"90",X"99",X"99",X"99",X"99",X"09",X"29",X"29",X"29",
		X"09",X"29",X"29",X"29",X"99",X"29",X"29",X"29",X"99",X"29",X"29",X"29",X"29",X"29",X"29",X"29",
		X"29",X"29",X"29",X"29",X"29",X"29",X"29",X"29",X"29",X"29",X"29",X"29",X"29",X"29",X"29",X"29",
		X"29",X"29",X"29",X"29",X"29",X"29",X"29",X"29",X"29",X"99",X"99",X"99",X"99",X"90",X"90",X"90",
		X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"92",X"09",X"09",X"00",X"92",X"99",X"99",X"90",X"92",X"92",X"92",X"90",
		X"92",X"92",X"92",X"90",X"92",X"92",X"92",X"90",X"92",X"92",X"92",X"90",X"92",X"92",X"92",X"90",
		X"99",X"92",X"92",X"90",X"00",X"92",X"92",X"90",X"00",X"92",X"92",X"90",X"99",X"92",X"92",X"90",
		X"92",X"92",X"92",X"90",X"92",X"92",X"92",X"90",X"99",X"99",X"99",X"90",X"99",X"09",X"09",X"00",
		X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"09",X"00",X"99",X"90",X"99",X"00",X"99",X"90",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"90",X"00",
		X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"99",X"00",
		X"99",X"00",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"90",X"00",X"99",X"99",X"90",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"9A",X"99",X"99",X"99",X"A9",X"99",X"99",X"99",X"99",X"99",X"99",
		X"09",X"99",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"A9",X"99",
		X"00",X"00",X"9A",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"99",X"00",X"00",X"99",
		X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"90",X"00",X"99",X"99",X"90",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"90",X"00",X"99",X"99",X"90",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"90",X"00",X"99",X"99",X"90",X"00",X"99",X"99",X"99",X"00",X"09",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",
		X"93",X"90",X"00",X"00",X"93",X"90",X"00",X"00",X"93",X"00",X"00",X"00",X"39",X"00",X"00",X"00",
		X"39",X"00",X"00",X"00",X"99",X"00",X"50",X"00",X"99",X"00",X"05",X"00",X"99",X"00",X"50",X"00",
		X"99",X"00",X"05",X"00",X"99",X"00",X"50",X"00",X"99",X"00",X"05",X"00",X"99",X"00",X"50",X"00",
		X"99",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"95",X"99",X"00",X"00",X"59",X"99",X"00",X"00",X"55",X"51",X"59",X"00",X"E5",X"44",X"15",
		X"00",X"EE",X"44",X"99",X"00",X"EE",X"99",X"99",X"00",X"E9",X"55",X"59",X"00",X"99",X"11",X"44",
		X"00",X"99",X"11",X"14",X"00",X"99",X"41",X"44",X"00",X"99",X"41",X"44",X"00",X"95",X"41",X"44",
		X"00",X"95",X"55",X"44",X"00",X"95",X"41",X"44",X"00",X"99",X"11",X"44",X"00",X"99",X"41",X"44",
		X"00",X"99",X"41",X"44",X"00",X"E9",X"51",X"44",X"00",X"EE",X"95",X"99",X"00",X"EE",X"19",X"99",
		X"00",X"E5",X"11",X"99",X"00",X"55",X"44",X"51",X"00",X"99",X"55",X"99",X"00",X"99",X"99",X"00",
		X"00",X"50",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"09",X"95",X"00",X"00",X"99",X"11",X"00",X"00",X"15",X"44",X"00",X"00",
		X"59",X"14",X"00",X"00",X"99",X"99",X"00",X"00",X"95",X"99",X"00",X"00",X"14",X"19",X"00",X"00",
		X"44",X"49",X"00",X"00",X"44",X"49",X"00",X"00",X"44",X"49",X"00",X"00",X"44",X"49",X"00",X"00",
		X"44",X"49",X"00",X"00",X"44",X"49",X"00",X"00",X"44",X"49",X"00",X"00",X"44",X"49",X"00",X"00",
		X"44",X"45",X"00",X"00",X"54",X"59",X"00",X"00",X"95",X"95",X"00",X"00",X"99",X"99",X"00",X"00",
		X"19",X"44",X"00",X"00",X"51",X"44",X"00",X"00",X"99",X"11",X"00",X"00",X"05",X"95",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"50",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"14",X"00",
		X"00",X"00",X"41",X"00",X"00",X"00",X"14",X"95",X"00",X"00",X"44",X"19",X"00",X"00",X"55",X"44",
		X"00",X"09",X"99",X"59",X"00",X"09",X"11",X"99",X"00",X"05",X"14",X"99",X"00",X"95",X"44",X"99",
		X"00",X"95",X"14",X"99",X"00",X"95",X"51",X"91",X"00",X"99",X"44",X"91",X"00",X"54",X"44",X"14",
		X"00",X"9E",X"14",X"14",X"00",X"EE",X"14",X"44",X"00",X"5E",X"54",X"44",X"00",X"33",X"51",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"59",X"00",X"00",X"00",
		X"91",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"95",X"99",X"00",X"00",X"54",X"44",X"00",X"00",
		X"15",X"14",X"00",X"00",X"44",X"55",X"90",X"00",X"44",X"95",X"59",X"00",X"44",X"49",X"59",X"00",
		X"00",X"95",X"95",X"14",X"00",X"99",X"19",X"44",X"00",X"00",X"45",X"44",X"00",X"00",X"44",X"44",
		X"00",X"00",X"51",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"19",
		X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"41",X"59",X"00",X"44",X"44",X"59",X"00",X"44",X"44",X"50",X"00",X"44",X"41",X"90",X"00",
		X"44",X"45",X"90",X"00",X"44",X"49",X"00",X"00",X"44",X"49",X"00",X"00",X"44",X"55",X"00",X"00",
		X"44",X"95",X"00",X"00",X"54",X"55",X"00",X"00",X"54",X"51",X"00",X"00",X"19",X"55",X"00",X"00",
		X"14",X"55",X"00",X"00",X"51",X"95",X"00",X"00",X"99",X"49",X"00",X"00",X"05",X"49",X"00",X"00",
		X"00",X"49",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"05",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"3E",X"00",X"00",X"00",X"1E",X"00",
		X"00",X"00",X"95",X"00",X"00",X"00",X"91",X"90",X"00",X"00",X"91",X"99",X"00",X"00",X"99",X"99",
		X"00",X"00",X"45",X"45",X"00",X"99",X"54",X"44",X"00",X"55",X"44",X"44",X"00",X"95",X"54",X"95",
		X"00",X"9E",X"11",X"19",X"00",X"EE",X"45",X"99",X"00",X"EE",X"44",X"99",X"00",X"53",X"11",X"99",
		X"00",X"55",X"14",X"99",X"00",X"95",X"44",X"91",X"00",X"09",X"44",X"14",X"00",X"09",X"14",X"44",
		X"00",X"00",X"54",X"44",X"00",X"00",X"95",X"44",X"00",X"00",X"99",X"44",X"00",X"00",X"99",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"19",X"00",X"00",X"00",
		X"91",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"59",X"00",X"00",X"00",
		X"00",X"00",X"19",X"44",X"00",X"00",X"51",X"44",X"00",X"00",X"59",X"44",X"00",X"00",X"99",X"14",
		X"00",X"00",X"09",X"44",X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"94",X"00",X"00",X"00",X"94",
		X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"49",X"00",X"00",X"00",X"45",X"00",X"00",X"00",X"55",
		X"00",X"00",X"00",X"94",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"59",X"50",X"00",X"00",X"45",X"90",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"49",X"00",X"00",
		X"45",X"41",X"00",X"00",X"99",X"44",X"00",X"00",X"55",X"44",X"00",X"00",X"99",X"54",X"00",X"00",
		X"95",X"94",X"00",X"00",X"94",X"59",X"00",X"00",X"14",X"55",X"00",X"00",X"44",X"59",X"00",X"00",
		X"44",X"59",X"00",X"00",X"44",X"91",X"00",X"00",X"44",X"51",X"00",X"00",X"45",X"11",X"00",X"00",
		X"95",X"55",X"00",X"00",X"55",X"55",X"00",X"00",X"55",X"50",X"00",X"00",X"49",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"45",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"55",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"1E",X"00",X"00",X"05",X"EE",
		X"00",X"00",X"99",X"EE",X"00",X"00",X"95",X"33",X"00",X"00",X"59",X"41",X"00",X"00",X"99",X"54",
		X"00",X"00",X"99",X"91",X"00",X"00",X"49",X"59",X"00",X"00",X"49",X"19",X"00",X"00",X"49",X"41",
		X"00",X"00",X"49",X"14",X"00",X"00",X"49",X"44",X"00",X"00",X"49",X"44",X"00",X"00",X"49",X"44",
		X"00",X"00",X"49",X"15",X"00",X"00",X"49",X"99",X"00",X"00",X"49",X"99",X"00",X"00",X"49",X"99",
		X"00",X"00",X"45",X"99",X"00",X"00",X"15",X"54",X"00",X"00",X"51",X"11",X"00",X"00",X"59",X"44",
		X"00",X"00",X"99",X"44",X"00",X"00",X"99",X"44",X"00",X"00",X"99",X"44",X"00",X"00",X"09",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"95",X"00",X"00",X"00",
		X"15",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"91",X"00",X"00",X"00",
		X"95",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"00",X"00",X"05",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",
		X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"54",
		X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"41",X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"14",
		X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",
		X"00",X"00",X"00",X"49",X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"14",
		X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"59",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"59",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"95",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"44",X"50",X"00",X"00",X"44",X"50",X"00",X"00",
		X"44",X"90",X"00",X"00",X"44",X"90",X"00",X"00",X"19",X"50",X"00",X"00",X"55",X"99",X"00",X"00",
		X"55",X"95",X"00",X"00",X"51",X"55",X"00",X"00",X"55",X"59",X"00",X"00",X"55",X"50",X"00",X"00",
		X"95",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"50",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"99",X"99",X"00",X"99",X"55",X"E5",X"00",
		X"99",X"99",X"EE",X"00",X"99",X"95",X"E9",X"00",X"99",X"55",X"31",X"00",X"59",X"49",X"41",X"00",
		X"55",X"55",X"41",X"00",X"99",X"11",X"41",X"00",X"99",X"45",X"11",X"00",X"99",X"15",X"11",X"00",
		X"99",X"45",X"41",X"00",X"99",X"41",X"41",X"00",X"99",X"41",X"41",X"00",X"99",X"45",X"41",X"00",
		X"55",X"41",X"44",X"00",X"55",X"59",X"14",X"00",X"55",X"99",X"14",X"00",X"59",X"99",X"54",X"00",
		X"55",X"99",X"94",X"00",X"99",X"99",X"15",X"00",X"99",X"41",X"99",X"00",X"59",X"11",X"49",X"00",
		X"59",X"41",X"59",X"00",X"09",X"44",X"19",X"00",X"59",X"44",X"99",X"00",X"09",X"44",X"19",X"00",
		X"09",X"44",X"99",X"00",X"09",X"44",X"19",X"00",X"09",X"44",X"59",X"00",X"09",X"44",X"19",X"00",
		X"09",X"44",X"49",X"00",X"09",X"44",X"49",X"00",X"09",X"44",X"19",X"00",X"09",X"44",X"15",X"00",
		X"59",X"11",X"55",X"00",X"95",X"99",X"51",X"00",X"95",X"99",X"55",X"00",X"95",X"99",X"54",X"00",
		X"95",X"41",X"54",X"00",X"95",X"41",X"14",X"00",X"95",X"44",X"14",X"00",X"95",X"41",X"44",X"00",
		X"95",X"44",X"44",X"00",X"95",X"95",X"44",X"00",X"95",X"59",X"44",X"00",X"95",X"15",X"44",X"00",
		X"55",X"55",X"44",X"00",X"59",X"55",X"99",X"00",X"99",X"15",X"99",X"00",X"99",X"55",X"55",X"00",
		X"99",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"09",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"A9",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"33",X"99",X"00",X"00",X"39",X"99",X"00",X"00",
		X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"00",X"05",X"00",X"99",X"00",X"50",X"00",
		X"99",X"00",X"05",X"00",X"99",X"00",X"50",X"00",X"99",X"00",X"05",X"00",X"90",X"00",X"50",X"00",
		X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"39",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"39",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"50",X"00",
		X"09",X"99",X"05",X"00",X"00",X"90",X"50",X"00",X"00",X"05",X"05",X"00",X"00",X"50",X"50",X"00",
		X"00",X"05",X"05",X"00",X"00",X"50",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"09",X"95",X"00",X"00",X"99",X"11",X"00",X"00",X"15",X"45",X"00",X"00",
		X"59",X"14",X"00",X"00",X"99",X"99",X"00",X"00",X"95",X"99",X"00",X"00",X"14",X"19",X"00",X"00",
		X"44",X"59",X"00",X"00",X"44",X"59",X"00",X"00",X"44",X"59",X"00",X"00",X"44",X"59",X"00",X"00",
		X"44",X"59",X"00",X"00",X"44",X"59",X"00",X"00",X"44",X"59",X"00",X"00",X"44",X"59",X"00",X"00",
		X"44",X"49",X"00",X"00",X"54",X"59",X"00",X"00",X"95",X"95",X"00",X"00",X"99",X"99",X"00",X"00",
		X"19",X"45",X"00",X"00",X"51",X"54",X"00",X"00",X"99",X"15",X"00",X"00",X"05",X"95",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"59",X"00",X"00",X"00",
		X"91",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"95",X"99",X"00",X"00",X"54",X"44",X"00",X"00",
		X"15",X"14",X"00",X"00",X"44",X"55",X"90",X"00",X"44",X"95",X"59",X"00",X"44",X"49",X"59",X"00",
		X"44",X"41",X"59",X"00",X"44",X"45",X"59",X"00",X"44",X"54",X"50",X"00",X"44",X"49",X"90",X"00",
		X"44",X"59",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",
		X"44",X"99",X"00",X"00",X"54",X"99",X"00",X"00",X"54",X"99",X"00",X"00",X"19",X"55",X"00",X"00",
		X"14",X"55",X"00",X"00",X"51",X"95",X"00",X"00",X"99",X"59",X"00",X"00",X"05",X"59",X"00",X"00",
		X"00",X"59",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"05",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"59",X"59",X"00",X"00",X"45",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"49",X"00",X"00",
		X"45",X"41",X"00",X"00",X"99",X"44",X"00",X"00",X"55",X"44",X"00",X"00",X"99",X"54",X"00",X"00",
		X"95",X"94",X"00",X"00",X"94",X"59",X"00",X"00",X"14",X"95",X"00",X"00",X"44",X"99",X"00",X"00",
		X"45",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"45",X"59",X"00",X"00",X"45",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"59",X"90",X"00",X"00",X"55",X"90",X"00",X"00",X"49",X"00",X"00",X"00",
		X"54",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"55",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"59",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"54",X"90",X"00",X"00",X"95",X"90",X"00",X"00",
		X"99",X"99",X"00",X"00",X"54",X"99",X"00",X"00",X"44",X"59",X"00",X"00",X"44",X"50",X"00",X"00",
		X"54",X"90",X"00",X"00",X"55",X"90",X"00",X"00",X"59",X"50",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"95",X"00",X"00",X"99",X"55",X"00",X"00",X"99",X"59",X"00",X"00",X"99",X"50",X"00",X"00",
		X"99",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"05",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",
		X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"54",
		X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"41",X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"14",
		X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",
		X"00",X"00",X"00",X"49",X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"49",X"00",X"00",X"00",X"14",
		X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"59",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"44",X"99",X"00",X"09",X"44",X"19",X"00",X"09",X"44",X"59",X"00",X"09",X"44",X"19",X"00",
		X"09",X"44",X"49",X"00",X"09",X"44",X"49",X"00",X"09",X"44",X"19",X"00",X"09",X"44",X"15",X"00",
		X"59",X"11",X"55",X"00",X"95",X"99",X"51",X"00",X"95",X"99",X"55",X"00",X"95",X"99",X"54",X"00",
		X"95",X"41",X"54",X"00",X"95",X"41",X"14",X"00",X"95",X"45",X"14",X"00",X"95",X"51",X"41",X"00",
		X"95",X"15",X"41",X"00",X"95",X"99",X"41",X"00",X"99",X"99",X"19",X"00",X"95",X"99",X"91",X"00",
		X"55",X"99",X"19",X"00",X"59",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"55",X"55",X"00",
		X"99",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",
		X"00",X"95",X"99",X"00",X"00",X"59",X"99",X"00",X"00",X"55",X"51",X"59",X"00",X"EE",X"44",X"15",
		X"00",X"EE",X"44",X"99",X"00",X"EE",X"99",X"99",X"00",X"15",X"59",X"59",X"00",X"99",X"99",X"44",
		X"00",X"99",X"99",X"14",X"00",X"99",X"D9",X"44",X"00",X"99",X"99",X"44",X"00",X"95",X"99",X"44",
		X"00",X"95",X"D9",X"44",X"00",X"95",X"99",X"44",X"00",X"99",X"99",X"44",X"00",X"99",X"D9",X"44",
		X"00",X"99",X"99",X"44",X"00",X"1E",X"99",X"44",X"00",X"EE",X"95",X"99",X"00",X"EE",X"19",X"99",
		X"00",X"EE",X"11",X"99",X"00",X"55",X"44",X"51",X"00",X"99",X"55",X"99",X"00",X"99",X"99",X"00",
		X"00",X"50",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"50",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"54",X"90",
		X"00",X"00",X"41",X"99",X"00",X"00",X"14",X"95",X"00",X"00",X"44",X"19",X"00",X"05",X"55",X"44",
		X"00",X"00",X"99",X"19",X"00",X"00",X"99",X"99",X"00",X"50",X"D9",X"99",X"00",X"00",X"DD",X"99",
		X"00",X"55",X"D9",X"99",X"00",X"55",X"99",X"91",X"00",X"59",X"99",X"91",X"00",X"53",X"D9",X"14",
		X"00",X"93",X"D9",X"14",X"00",X"9E",X"9D",X"44",X"00",X"5E",X"99",X"44",X"00",X"15",X"51",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"35",X"00",X"00",X"00",X"3E",X"90",
		X"00",X"00",X"9E",X"99",X"00",X"00",X"9E",X"99",X"00",X"00",X"93",X"99",X"00",X"00",X"99",X"99",
		X"00",X"00",X"9D",X"45",X"00",X"99",X"99",X"44",X"00",X"55",X"DD",X"44",X"00",X"95",X"99",X"95",
		X"00",X"95",X"99",X"19",X"00",X"9E",X"DD",X"99",X"00",X"5E",X"D9",X"99",X"00",X"53",X"DD",X"99",
		X"00",X"55",X"99",X"99",X"00",X"95",X"99",X"91",X"00",X"09",X"94",X"14",X"00",X"09",X"94",X"44",
		X"00",X"00",X"54",X"44",X"00",X"00",X"91",X"44",X"00",X"00",X"91",X"44",X"00",X"00",X"99",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"95",X"00",X"00",X"00",
		X"15",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"91",X"00",X"00",X"00",
		X"95",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"3E",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"09",X"EE",X"00",X"00",X"95",X"E3",X"00",X"00",X"59",X"31",X"00",X"00",X"99",X"54",
		X"00",X"00",X"E9",X"91",X"00",X"00",X"E9",X"99",X"00",X"00",X"39",X"99",X"00",X"00",X"49",X"D9",
		X"00",X"00",X"49",X"D9",X"00",X"00",X"49",X"99",X"00",X"00",X"49",X"99",X"00",X"00",X"49",X"41",
		X"00",X"00",X"49",X"15",X"00",X"00",X"49",X"99",X"00",X"00",X"49",X"99",X"00",X"00",X"49",X"99",
		X"00",X"00",X"45",X"99",X"00",X"00",X"11",X"54",X"00",X"00",X"51",X"11",X"00",X"00",X"59",X"44",
		X"00",X"00",X"99",X"44",X"00",X"00",X"99",X"44",X"00",X"00",X"99",X"44",X"00",X"00",X"09",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"99",X"99",X"00",X"99",X"55",X"95",X"00",
		X"99",X"99",X"E5",X"00",X"99",X"DD",X"E5",X"00",X"95",X"59",X"33",X"00",X"59",X"D9",X"45",X"00",
		X"55",X"DD",X"51",X"00",X"99",X"DD",X"45",X"00",X"99",X"D9",X"11",X"00",X"99",X"D9",X"11",X"00",
		X"99",X"DD",X"41",X"00",X"99",X"D9",X"41",X"00",X"99",X"99",X"41",X"00",X"99",X"99",X"41",X"00",
		X"55",X"11",X"44",X"00",X"55",X"59",X"14",X"00",X"55",X"99",X"14",X"00",X"59",X"99",X"54",X"00",
		X"55",X"99",X"94",X"00",X"99",X"99",X"15",X"00",X"99",X"41",X"99",X"00",X"59",X"11",X"49",X"00",
		X"59",X"41",X"59",X"00",X"09",X"44",X"19",X"00",X"59",X"44",X"99",X"00",X"09",X"44",X"19",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"95",X"09",X"00",X"00",X"59",X"99",X"00",X"00",X"55",X"51",X"59",X"00",X"E5",X"44",X"15",
		X"00",X"EE",X"44",X"99",X"00",X"EE",X"99",X"99",X"00",X"15",X"59",X"59",X"00",X"99",X"99",X"44",
		X"00",X"99",X"99",X"14",X"00",X"99",X"D9",X"44",X"00",X"99",X"99",X"44",X"00",X"95",X"99",X"44",
		X"00",X"95",X"D9",X"44",X"00",X"95",X"99",X"44",X"00",X"99",X"99",X"44",X"00",X"99",X"D9",X"44",
		X"00",X"99",X"99",X"44",X"00",X"1E",X"99",X"44",X"00",X"EE",X"95",X"99",X"00",X"EE",X"19",X"99",
		X"00",X"35",X"11",X"99",X"00",X"55",X"44",X"51",X"00",X"99",X"55",X"99",X"00",X"99",X"99",X"00",
		X"00",X"50",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"59",X"00",X"00",X"00",
		X"91",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"95",X"99",X"00",X"00",X"54",X"44",X"00",X"00",
		X"15",X"14",X"00",X"00",X"44",X"55",X"90",X"00",X"44",X"95",X"59",X"00",X"44",X"49",X"59",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"50",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"34",X"00",
		X"00",X"00",X"31",X"90",X"00",X"00",X"14",X"95",X"00",X"00",X"44",X"19",X"00",X"05",X"55",X"44",
		X"00",X"00",X"99",X"19",X"00",X"00",X"99",X"99",X"00",X"50",X"D9",X"99",X"00",X"00",X"DD",X"99",
		X"00",X"55",X"D9",X"99",X"00",X"55",X"99",X"91",X"00",X"59",X"99",X"91",X"00",X"54",X"D9",X"14",
		X"00",X"95",X"D9",X"14",X"00",X"9E",X"9D",X"44",X"00",X"5E",X"99",X"44",X"00",X"15",X"51",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"3E",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"9E",X"90",X"00",X"00",X"91",X"99",X"00",X"00",X"99",X"99",
		X"00",X"00",X"9D",X"45",X"00",X"99",X"99",X"44",X"00",X"55",X"DD",X"44",X"00",X"95",X"99",X"95",
		X"00",X"95",X"99",X"19",X"00",X"9E",X"DD",X"99",X"00",X"5E",X"D9",X"99",X"00",X"53",X"DD",X"99",
		X"00",X"55",X"99",X"99",X"00",X"95",X"99",X"91",X"00",X"99",X"94",X"14",X"00",X"99",X"94",X"44",
		X"00",X"99",X"54",X"44",X"00",X"99",X"91",X"44",X"00",X"09",X"91",X"44",X"00",X"00",X"99",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"95",X"00",X"00",X"00",
		X"15",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"91",X"00",X"00",X"00",
		X"95",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"1E",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"09",X"EE",X"00",X"00",X"95",X"E3",X"00",X"00",X"59",X"33",X"00",X"00",X"99",X"54",
		X"00",X"00",X"E9",X"91",X"00",X"00",X"E9",X"99",X"00",X"00",X"39",X"99",X"00",X"00",X"49",X"D9",
		X"00",X"00",X"49",X"D9",X"00",X"00",X"49",X"99",X"00",X"00",X"49",X"99",X"00",X"00",X"49",X"41",
		X"00",X"00",X"49",X"15",X"00",X"00",X"49",X"99",X"00",X"00",X"49",X"99",X"00",X"00",X"49",X"99",
		X"00",X"00",X"45",X"99",X"00",X"00",X"11",X"54",X"00",X"00",X"51",X"11",X"00",X"00",X"59",X"44",
		X"00",X"00",X"99",X"44",X"00",X"00",X"99",X"44",X"00",X"00",X"99",X"44",X"00",X"00",X"09",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"99",X"99",X"00",X"99",X"55",X"95",X"00",
		X"99",X"99",X"E5",X"00",X"99",X"DD",X"E5",X"00",X"95",X"59",X"35",X"00",X"59",X"D9",X"45",X"00",
		X"55",X"DD",X"51",X"00",X"99",X"DD",X"45",X"00",X"99",X"D9",X"11",X"00",X"99",X"D9",X"11",X"00",
		X"99",X"DD",X"41",X"00",X"99",X"D9",X"41",X"00",X"99",X"99",X"41",X"00",X"99",X"99",X"41",X"00",
		X"55",X"11",X"44",X"00",X"55",X"59",X"14",X"00",X"55",X"99",X"14",X"00",X"59",X"99",X"54",X"00",
		X"55",X"99",X"94",X"00",X"99",X"99",X"15",X"00",X"99",X"41",X"99",X"00",X"59",X"11",X"49",X"00",
		X"59",X"41",X"59",X"00",X"09",X"44",X"19",X"00",X"59",X"44",X"99",X"00",X"09",X"44",X"19",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"00",X"09",X"95",X"00",X"00",X"99",X"11",X"00",X"00",X"15",X"45",X"00",X"00",
		X"59",X"14",X"00",X"00",X"99",X"99",X"00",X"00",X"95",X"99",X"00",X"00",X"14",X"19",X"00",X"00",
		X"44",X"59",X"00",X"00",X"44",X"59",X"00",X"00",X"44",X"59",X"00",X"00",X"44",X"59",X"00",X"00",
		X"44",X"59",X"00",X"00",X"44",X"59",X"00",X"00",X"44",X"59",X"00",X"00",X"44",X"59",X"00",X"00",
		X"44",X"49",X"00",X"00",X"54",X"59",X"00",X"00",X"95",X"95",X"00",X"00",X"99",X"99",X"00",X"00",
		X"19",X"45",X"00",X"00",X"51",X"54",X"00",X"00",X"99",X"15",X"00",X"00",X"05",X"95",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"41",X"59",X"00",X"44",X"45",X"59",X"00",X"44",X"54",X"50",X"00",X"44",X"49",X"90",X"00",
		X"44",X"59",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",
		X"44",X"99",X"00",X"00",X"54",X"99",X"00",X"00",X"54",X"99",X"00",X"00",X"19",X"55",X"00",X"00",
		X"14",X"55",X"00",X"00",X"51",X"95",X"00",X"00",X"99",X"59",X"00",X"00",X"99",X"59",X"00",X"00",
		X"99",X"59",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"05",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"95",X"95",X"14",X"00",X"99",X"19",X"44",X"00",X"99",X"45",X"44",X"00",X"99",X"44",X"44",
		X"00",X"99",X"51",X"99",X"00",X"09",X"99",X"99",X"00",X"00",X"90",X"99",X"00",X"00",X"00",X"19",
		X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"59",X"00",X"00",X"00",X"45",X"90",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"49",X"00",X"00",
		X"45",X"41",X"00",X"00",X"99",X"44",X"00",X"00",X"55",X"44",X"00",X"00",X"99",X"54",X"00",X"00",
		X"95",X"94",X"00",X"00",X"94",X"59",X"00",X"00",X"14",X"95",X"00",X"00",X"44",X"99",X"00",X"00",
		X"45",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"45",X"59",X"00",X"00",X"45",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"59",X"90",X"00",X"00",X"55",X"90",X"00",X"00",X"49",X"00",X"00",X"00",
		X"54",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"55",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"59",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"95",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"44",X"50",X"00",X"00",X"44",X"50",X"00",X"00",
		X"54",X"90",X"00",X"00",X"55",X"90",X"00",X"00",X"59",X"50",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"95",X"00",X"00",X"99",X"55",X"00",X"00",X"99",X"59",X"00",X"00",X"99",X"50",X"00",X"00",
		X"99",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"05",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",
		X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"54",
		X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"41",X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"14",
		X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",
		X"00",X"00",X"00",X"49",X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"49",X"00",X"00",X"00",X"14",
		X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"59",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"44",X"99",X"00",X"09",X"44",X"19",X"00",X"09",X"44",X"59",X"00",X"09",X"44",X"19",X"00",
		X"09",X"44",X"49",X"00",X"09",X"44",X"49",X"00",X"09",X"44",X"19",X"00",X"09",X"44",X"15",X"00",
		X"59",X"11",X"55",X"00",X"95",X"99",X"51",X"00",X"95",X"99",X"55",X"00",X"95",X"99",X"54",X"00",
		X"95",X"41",X"54",X"00",X"95",X"41",X"14",X"00",X"95",X"45",X"14",X"00",X"95",X"51",X"41",X"00",
		X"95",X"15",X"41",X"00",X"95",X"99",X"41",X"00",X"99",X"99",X"19",X"00",X"95",X"99",X"91",X"00",
		X"55",X"99",X"19",X"00",X"59",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"55",X"55",X"00",
		X"99",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",
		X"C0",X"99",X"CC",X"00",X"CC",X"99",X"C0",X"00",X"0C",X"D9",X"CC",X"00",X"00",X"99",X"0C",X"00",
		X"00",X"99",X"00",X"00",X"00",X"95",X"50",X"00",X"C0",X"50",X"05",X"00",X"0C",X"05",X"50",X"00",
		X"CC",X"50",X"05",X"00",X"CC",X"00",X"50",X"00",X"0C",X"90",X"0C",X"00",X"CC",X"99",X"5C",X"00",
		X"0C",X"99",X"00",X"00",X"C0",X"99",X"50",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"05",X"CC",X"00",X"00",X"50",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"0C",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"77",X"00",X"00",X"07",X"75",X"00",X"00",X"75",X"75",X"00",X"00",X"57",X"57",
		X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",
		X"00",X"00",X"77",X"11",X"00",X"00",X"74",X"32",X"00",X"00",X"74",X"33",X"00",X"00",X"41",X"33",
		X"00",X"00",X"42",X"33",X"00",X"00",X"41",X"33",X"00",X"00",X"11",X"33",X"00",X"00",X"12",X"33",
		X"00",X"00",X"41",X"33",X"00",X"00",X"42",X"32",X"00",X"00",X"44",X"33",X"00",X"00",X"44",X"23",
		X"00",X"00",X"74",X"21",X"00",X"00",X"77",X"21",X"00",X"00",X"74",X"31",X"00",X"00",X"41",X"31",
		X"00",X"00",X"42",X"24",X"00",X"00",X"12",X"24",X"00",X"00",X"12",X"24",X"00",X"00",X"42",X"24",
		X"00",X"00",X"41",X"24",X"00",X"00",X"41",X"24",X"00",X"00",X"71",X"34",X"00",X"00",X"71",X"34",
		X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",
		X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"70",X"00",X"77",X"77",X"77",X"00",
		X"77",X"77",X"70",X"00",X"77",X"77",X"07",X"00",X"77",X"77",X"70",X"00",X"77",X"77",X"77",X"00",
		X"77",X"77",X"77",X"00",X"47",X"77",X"77",X"00",X"14",X"77",X"77",X"00",X"14",X"77",X"77",X"00",
		X"14",X"77",X"77",X"00",X"14",X"77",X"77",X"00",X"77",X"77",X"77",X"00",X"77",X"77",X"77",X"00",
		X"77",X"77",X"77",X"00",X"77",X"77",X"77",X"00",X"77",X"77",X"77",X"70",X"77",X"77",X"77",X"00",
		X"41",X"77",X"77",X"00",X"22",X"77",X"77",X"04",X"22",X"77",X"77",X"70",X"32",X"77",X"77",X"74",
		X"22",X"77",X"77",X"70",X"22",X"77",X"77",X"40",X"21",X"77",X"77",X"40",X"21",X"77",X"77",X"74",
		X"00",X"00",X"74",X"17",X"00",X"00",X"77",X"11",X"00",X"00",X"77",X"22",X"00",X"00",X"77",X"22",
		X"00",X"00",X"77",X"44",X"00",X"00",X"77",X"6F",X"00",X"00",X"77",X"11",X"00",X"00",X"77",X"12",
		X"00",X"00",X"07",X"14",X"00",X"00",X"07",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"41",
		X"00",X"00",X"00",X"42",X"00",X"00",X"00",X"42",X"00",X"00",X"0B",X"42",X"00",X"00",X"BB",X"22",
		X"00",X"00",X"CB",X"22",X"00",X"9B",X"B9",X"22",X"00",X"99",X"B9",X"22",X"99",X"B9",X"99",X"22",
		X"AA",X"BB",X"99",X"22",X"AB",X"9A",X"99",X"22",X"AC",X"AA",X"79",X"22",X"CB",X"AA",X"79",X"22",
		X"BB",X"AA",X"79",X"22",X"BB",X"AA",X"77",X"22",X"BB",X"AA",X"77",X"22",X"BB",X"AA",X"99",X"22",
		X"21",X"77",X"77",X"77",X"24",X"77",X"77",X"77",X"24",X"77",X"77",X"77",X"22",X"77",X"77",X"77",
		X"22",X"77",X"77",X"77",X"21",X"77",X"77",X"77",X"21",X"77",X"77",X"77",X"14",X"77",X"77",X"77",
		X"14",X"77",X"77",X"77",X"47",X"77",X"77",X"77",X"77",X"97",X"77",X"77",X"47",X"A9",X"77",X"77",
		X"77",X"77",X"77",X"77",X"44",X"47",X"77",X"77",X"44",X"17",X"77",X"77",X"44",X"11",X"77",X"77",
		X"11",X"11",X"77",X"77",X"11",X"22",X"77",X"77",X"11",X"12",X"47",X"77",X"21",X"12",X"77",X"77",
		X"12",X"11",X"99",X"77",X"21",X"11",X"A9",X"77",X"22",X"11",X"A9",X"77",X"22",X"14",X"A9",X"99",
		X"22",X"29",X"AA",X"99",X"32",X"4A",X"AA",X"99",X"23",X"9A",X"AA",X"99",X"22",X"9A",X"BA",X"99",
		X"22",X"9C",X"AA",X"99",X"22",X"AC",X"9A",X"99",X"22",X"AB",X"9A",X"99",X"22",X"BB",X"99",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"9B",X"00",X"00",X"00",X"9B",
		X"00",X"00",X"00",X"9C",X"00",X"00",X"00",X"9C",X"00",X"00",X"00",X"BC",X"00",X"00",X"00",X"CB",
		X"00",X"00",X"00",X"CB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"AB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BA",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"7A",X"00",X"00",X"00",X"77",
		X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",
		X"00",X"00",X"02",X"21",X"00",X"00",X"02",X"11",X"00",X"00",X"23",X"21",X"00",X"00",X"23",X"14",
		X"00",X"00",X"22",X"11",X"00",X"00",X"32",X"14",X"00",X"00",X"22",X"11",X"00",X"00",X"22",X"11",
		X"BB",X"A9",X"79",X"22",X"BA",X"AA",X"99",X"22",X"BA",X"AA",X"99",X"22",X"AB",X"AA",X"99",X"22",
		X"A9",X"AA",X"A9",X"22",X"AA",X"AA",X"A9",X"12",X"AA",X"AA",X"99",X"22",X"AA",X"AA",X"99",X"12",
		X"A9",X"AA",X"99",X"11",X"A9",X"AA",X"99",X"12",X"94",X"AA",X"99",X"11",X"94",X"AA",X"99",X"12",
		X"44",X"AA",X"99",X"11",X"49",X"AA",X"99",X"11",X"4A",X"AA",X"99",X"11",X"4A",X"A9",X"A9",X"11",
		X"99",X"AA",X"99",X"11",X"99",X"A9",X"97",X"11",X"9A",X"AA",X"79",X"41",X"AA",X"AA",X"97",X"41",
		X"AB",X"AA",X"99",X"41",X"BB",X"AA",X"97",X"41",X"BA",X"BA",X"99",X"41",X"BB",X"AA",X"97",X"41",
		X"BB",X"AA",X"99",X"41",X"BB",X"AA",X"99",X"44",X"BB",X"BB",X"97",X"41",X"BC",X"BA",X"99",X"44",
		X"BD",X"BA",X"99",X"41",X"CC",X"BA",X"99",X"44",X"BB",X"BB",X"97",X"41",X"AA",X"BA",X"99",X"47",
		X"22",X"BA",X"7B",X"BA",X"12",X"BA",X"97",X"BB",X"22",X"A9",X"97",X"CB",X"22",X"99",X"99",X"CB",
		X"22",X"9A",X"99",X"BB",X"22",X"99",X"AA",X"BB",X"2A",X"99",X"BB",X"BA",X"2A",X"9A",X"AA",X"BB",
		X"49",X"AA",X"BB",X"BA",X"4B",X"AA",X"BB",X"BA",X"BB",X"AA",X"AB",X"AA",X"BB",X"AA",X"BB",X"BA",
		X"BA",X"AA",X"AA",X"7A",X"AA",X"AB",X"BA",X"AA",X"AA",X"AA",X"BA",X"AA",X"AA",X"BA",X"BB",X"AA",
		X"BA",X"BA",X"BA",X"BB",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A9",X"AA",X"AA",X"AA",X"A9",X"AA",
		X"AA",X"AA",X"A9",X"AA",X"AA",X"AA",X"99",X"AA",X"AA",X"AA",X"99",X"AA",X"BA",X"AA",X"97",X"AA",
		X"AA",X"AA",X"77",X"AA",X"BB",X"AA",X"77",X"AA",X"AB",X"AA",X"77",X"AA",X"BB",X"AA",X"77",X"AA",
		X"BB",X"AA",X"77",X"7A",X"BB",X"BB",X"77",X"77",X"BB",X"BB",X"77",X"21",X"BB",X"BB",X"77",X"11",
		X"00",X"00",X"22",X"10",X"00",X"00",X"22",X"10",X"00",X"00",X"22",X"10",X"00",X"00",X"22",X"00",
		X"00",X"00",X"22",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"21",X"00",
		X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"02",X"21",X"00",X"00",X"22",X"11",X"00",
		X"00",X"22",X"14",X"00",X"00",X"22",X"41",X"00",X"00",X"22",X"10",X"00",X"00",X"22",X"41",X"00",
		X"00",X"22",X"11",X"00",X"00",X"22",X"14",X"00",X"00",X"12",X"11",X"00",X"00",X"22",X"11",X"00",
		X"00",X"12",X"12",X"00",X"00",X"22",X"12",X"00",X"00",X"12",X"21",X"00",X"00",X"11",X"21",X"00",
		X"00",X"01",X"21",X"00",X"00",X"01",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",
		X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"32",X"00",X"00",X"00",X"32",X"00",
		X"AA",X"BA",X"99",X"9B",X"AA",X"AA",X"99",X"7A",X"AA",X"AA",X"97",X"BA",X"AA",X"AA",X"79",X"BA",
		X"AA",X"AA",X"99",X"BA",X"A9",X"AA",X"79",X"AA",X"9A",X"A9",X"99",X"AA",X"B9",X"99",X"99",X"AA",
		X"99",X"99",X"A9",X"99",X"99",X"99",X"AA",X"99",X"99",X"AA",X"AA",X"99",X"99",X"AA",X"AA",X"99",
		X"99",X"AA",X"B9",X"99",X"74",X"99",X"B9",X"99",X"77",X"B9",X"B9",X"99",X"77",X"B9",X"BB",X"99",
		X"97",X"9B",X"BB",X"A9",X"09",X"94",X"BB",X"AA",X"09",X"79",X"AB",X"DA",X"00",X"17",X"9A",X"99",
		X"00",X"11",X"9B",X"9B",X"00",X"12",X"BB",X"BA",X"00",X"21",X"AB",X"AA",X"00",X"22",X"99",X"BB",
		X"00",X"22",X"BA",X"AA",X"00",X"22",X"BB",X"AA",X"00",X"22",X"BB",X"77",X"00",X"22",X"9B",X"44",
		X"00",X"22",X"77",X"DC",X"00",X"22",X"79",X"22",X"00",X"22",X"27",X"22",X"00",X"22",X"27",X"22",
		X"BB",X"AA",X"77",X"21",X"BC",X"A7",X"77",X"21",X"CC",X"99",X"77",X"21",X"CC",X"9A",X"77",X"21",
		X"CC",X"99",X"77",X"22",X"CD",X"A9",X"77",X"22",X"CD",X"A9",X"77",X"22",X"BC",X"BA",X"77",X"22",
		X"BC",X"AA",X"77",X"22",X"BB",X"AA",X"77",X"22",X"BB",X"AA",X"77",X"22",X"AB",X"A9",X"77",X"22",
		X"AA",X"A9",X"77",X"22",X"AA",X"99",X"79",X"22",X"A9",X"99",X"97",X"22",X"A9",X"77",X"77",X"22",
		X"99",X"97",X"07",X"22",X"99",X"79",X"07",X"22",X"99",X"77",X"04",X"22",X"99",X"77",X"04",X"22",
		X"A9",X"77",X"04",X"22",X"BB",X"77",X"04",X"22",X"B9",X"77",X"04",X"22",X"99",X"77",X"00",X"22",
		X"77",X"77",X"04",X"22",X"99",X"77",X"04",X"21",X"77",X"77",X"04",X"22",X"77",X"79",X"04",X"21",
		X"21",X"77",X"04",X"22",X"11",X"94",X"04",X"21",X"11",X"20",X"04",X"12",X"11",X"40",X"04",X"21",
		X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",
		X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"20",X"00",X"00",X"22",X"20",X"00",X"00",X"12",X"20",
		X"00",X"00",X"12",X"12",X"00",X"00",X"11",X"12",X"00",X"00",X"01",X"11",X"00",X"00",X"01",X"21",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"21",
		X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"21",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"12",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"22",X"21",X"22",X"00",X"22",X"21",X"22",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",
		X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"32",X"00",X"22",X"22",X"23",
		X"00",X"22",X"22",X"32",X"00",X"22",X"22",X"23",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",
		X"00",X"22",X"22",X"23",X"00",X"12",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"41",X"22",X"22",
		X"00",X"42",X"22",X"22",X"00",X"44",X"22",X"22",X"22",X"44",X"22",X"22",X"11",X"11",X"22",X"22",
		X"22",X"C2",X"11",X"22",X"21",X"22",X"11",X"22",X"12",X"12",X"11",X"25",X"22",X"11",X"41",X"5E",
		X"22",X"22",X"44",X"EE",X"11",X"22",X"77",X"55",X"21",X"12",X"77",X"EE",X"21",X"41",X"44",X"75",
		X"22",X"41",X"55",X"57",X"12",X"74",X"EE",X"57",X"21",X"77",X"7E",X"57",X"02",X"77",X"75",X"55",
		X"21",X"27",X"04",X"22",X"22",X"27",X"00",X"12",X"22",X"42",X"00",X"22",X"22",X"44",X"00",X"22",
		X"22",X"47",X"00",X"22",X"22",X"4E",X"00",X"22",X"22",X"75",X"00",X"22",X"22",X"57",X"00",X"22",
		X"22",X"57",X"00",X"22",X"22",X"55",X"00",X"22",X"22",X"57",X"00",X"22",X"22",X"77",X"00",X"22",
		X"22",X"77",X"00",X"22",X"22",X"77",X"E0",X"12",X"22",X"75",X"50",X"12",X"27",X"75",X"7E",X"11",
		X"7E",X"57",X"55",X"41",X"EE",X"55",X"57",X"01",X"EE",X"E5",X"75",X"04",X"7E",X"75",X"57",X"00",
		X"7E",X"55",X"75",X"00",X"57",X"55",X"77",X"00",X"57",X"55",X"57",X"00",X"57",X"55",X"75",X"00",
		X"5E",X"55",X"57",X"00",X"57",X"55",X"55",X"00",X"55",X"55",X"57",X"00",X"55",X"55",X"55",X"00",
		X"75",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"41",
		X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"32",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"23",
		X"00",X"00",X"00",X"32",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",
		X"00",X"00",X"01",X"22",X"00",X"00",X"11",X"22",X"00",X"00",X"12",X"22",X"00",X"00",X"22",X"22",
		X"00",X"00",X"22",X"22",X"00",X"00",X"21",X"22",X"00",X"00",X"22",X"12",X"00",X"00",X"22",X"22",
		X"00",X"77",X"77",X"55",X"00",X"77",X"57",X"55",X"04",X"77",X"55",X"55",X"07",X"77",X"55",X"55",
		X"47",X"77",X"55",X"57",X"77",X"75",X"45",X"55",X"55",X"57",X"54",X"55",X"55",X"55",X"75",X"57",
		X"5E",X"55",X"57",X"75",X"EE",X"55",X"55",X"57",X"55",X"55",X"55",X"75",X"27",X"55",X"75",X"54",
		X"21",X"55",X"77",X"77",X"2E",X"55",X"55",X"77",X"EE",X"5E",X"E5",X"77",X"55",X"55",X"E5",X"77",
		X"22",X"55",X"E5",X"77",X"22",X"E5",X"5E",X"77",X"22",X"EE",X"55",X"77",X"22",X"5E",X"55",X"77",
		X"21",X"77",X"55",X"77",X"22",X"11",X"55",X"77",X"12",X"22",X"57",X"77",X"21",X"12",X"77",X"77",
		X"22",X"22",X"77",X"57",X"22",X"22",X"77",X"77",X"12",X"22",X"77",X"55",X"22",X"21",X"77",X"00",
		X"22",X"11",X"77",X"00",X"22",X"11",X"74",X"00",X"22",X"11",X"17",X"00",X"11",X"17",X"74",X"00",
		X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"E5",X"55",X"00",
		X"55",X"55",X"55",X"00",X"75",X"55",X"55",X"00",X"55",X"E5",X"55",X"00",X"57",X"E5",X"55",X"00",
		X"55",X"5E",X"55",X"00",X"75",X"EE",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",
		X"55",X"EE",X"55",X"00",X"55",X"E5",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"77",X"55",X"00",
		X"55",X"11",X"75",X"00",X"77",X"11",X"77",X"00",X"11",X"22",X"17",X"00",X"12",X"22",X"21",X"00",
		X"22",X"22",X"12",X"00",X"22",X"22",X"21",X"00",X"22",X"23",X"22",X"00",X"22",X"22",X"21",X"00",
		X"22",X"22",X"21",X"00",X"22",X"22",X"21",X"00",X"22",X"22",X"11",X"00",X"22",X"22",X"21",X"00",
		X"22",X"22",X"12",X"00",X"22",X"22",X"21",X"00",X"22",X"22",X"11",X"00",X"22",X"22",X"11",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"70",X"00",X"CC",X"00",X"44",X"44",X"CC",X"00",
		X"CC",X"BC",X"C9",X"00",X"CC",X"BA",X"99",X"00",X"CC",X"BD",X"49",X"00",X"CC",X"CD",X"49",X"00",
		X"CC",X"CD",X"49",X"00",X"CC",X"CD",X"4B",X"00",X"CC",X"CD",X"7D",X"00",X"CC",X"CD",X"7D",X"00",
		X"CC",X"DD",X"7D",X"00",X"CC",X"DD",X"7F",X"00",X"CC",X"DD",X"CD",X"00",X"1C",X"DD",X"DD",X"00",
		X"CC",X"DD",X"DC",X"00",X"CC",X"DD",X"D7",X"00",X"0C",X"DD",X"C7",X"00",X"7C",X"DD",X"70",X"00",
		X"0C",X"CD",X"70",X"00",X"D4",X"DD",X"00",X"00",X"D4",X"DD",X"00",X"00",X"7D",X"CD",X"00",X"00",
		X"7D",X"DD",X"00",X"00",X"77",X"D4",X"00",X"00",X"07",X"4C",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"DC",X"00",X"00",X"00",X"DC",X"00",X"00",X"00",X"DC",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"BC",X"00",X"00",X"00",X"BC",X"00",X"00",X"0C",X"DD",X"00",X"00",X"7C",X"DD",X"00",X"00",
		X"7C",X"DD",X"00",X"00",X"7C",X"CD",X"00",X"00",X"77",X"77",X"70",X"00",X"77",X"77",X"70",X"00",
		X"77",X"77",X"70",X"00",X"57",X"77",X"70",X"00",X"57",X"77",X"70",X"00",X"57",X"77",X"70",X"00",
		X"57",X"77",X"70",X"00",X"57",X"77",X"70",X"00",X"57",X"77",X"70",X"00",X"57",X"77",X"70",X"00",
		X"57",X"77",X"70",X"00",X"57",X"77",X"70",X"00",X"55",X"77",X"70",X"00",X"57",X"77",X"70",X"00",
		X"77",X"77",X"70",X"00",X"77",X"77",X"70",X"00",X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BB",X"A9",X"79",X"22",X"BA",X"AA",X"99",X"22",X"BA",X"AA",X"99",X"22",X"AB",X"AA",X"99",X"22",
		X"A9",X"AA",X"A9",X"22",X"AA",X"AA",X"A9",X"12",X"AA",X"AA",X"99",X"22",X"AA",X"AA",X"99",X"12",
		X"A9",X"AA",X"99",X"11",X"A9",X"AA",X"99",X"12",X"94",X"AA",X"99",X"11",X"94",X"AA",X"99",X"12",
		X"44",X"AA",X"99",X"11",X"49",X"AA",X"99",X"11",X"4A",X"AA",X"99",X"11",X"4A",X"A9",X"A9",X"11",
		X"99",X"AA",X"99",X"11",X"99",X"A9",X"97",X"11",X"9A",X"AA",X"79",X"41",X"AA",X"AA",X"97",X"41",
		X"AB",X"AA",X"99",X"41",X"BB",X"AA",X"97",X"41",X"BA",X"BA",X"99",X"41",X"BB",X"AA",X"97",X"41",
		X"BB",X"AA",X"99",X"41",X"BB",X"AA",X"99",X"44",X"BB",X"BB",X"97",X"41",X"BC",X"BA",X"99",X"44",
		X"BD",X"BA",X"99",X"41",X"CC",X"BA",X"99",X"44",X"BB",X"BB",X"97",X"41",X"AA",X"BA",X"99",X"47",
		X"BB",X"AA",X"77",X"21",X"BC",X"AA",X"77",X"21",X"CC",X"BA",X"77",X"21",X"CC",X"AB",X"77",X"21",
		X"CC",X"9A",X"77",X"22",X"CD",X"A9",X"77",X"22",X"CD",X"A9",X"77",X"22",X"BC",X"BA",X"77",X"22",
		X"BC",X"AA",X"77",X"22",X"BB",X"AA",X"77",X"22",X"BB",X"AA",X"77",X"22",X"AB",X"A9",X"77",X"22",
		X"AA",X"A9",X"77",X"22",X"AA",X"99",X"79",X"22",X"A9",X"99",X"97",X"22",X"A9",X"77",X"77",X"22",
		X"99",X"97",X"07",X"22",X"99",X"79",X"07",X"22",X"99",X"77",X"04",X"22",X"99",X"77",X"04",X"22",
		X"A9",X"77",X"04",X"22",X"BB",X"77",X"04",X"22",X"B9",X"77",X"04",X"22",X"99",X"77",X"00",X"22",
		X"77",X"77",X"04",X"22",X"99",X"77",X"04",X"21",X"77",X"77",X"04",X"22",X"77",X"79",X"04",X"21",
		X"21",X"77",X"04",X"22",X"11",X"94",X"04",X"21",X"11",X"20",X"04",X"12",X"11",X"40",X"04",X"21",
		X"00",X"07",X"00",X"00",X"00",X"77",X"70",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",
		X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"14",X"77",X"00",X"00",X"32",X"77",X"00",
		X"00",X"33",X"77",X"00",X"00",X"33",X"77",X"00",X"00",X"32",X"77",X"00",X"00",X"33",X"77",X"00",
		X"00",X"21",X"77",X"00",X"00",X"37",X"77",X"70",X"00",X"24",X"77",X"00",X"00",X"24",X"77",X"70",
		X"00",X"27",X"77",X"70",X"00",X"37",X"77",X"70",X"00",X"17",X"77",X"77",X"00",X"22",X"77",X"77",
		X"00",X"44",X"77",X"77",X"00",X"22",X"77",X"77",X"00",X"14",X"77",X"77",X"00",X"23",X"97",X"77",
		X"00",X"22",X"7A",X"77",X"00",X"14",X"17",X"77",X"00",X"41",X"11",X"70",X"00",X"42",X"12",X"70",
		X"00",X"12",X"11",X"70",X"99",X"22",X"14",X"77",X"BB",X"22",X"2A",X"97",X"A9",X"22",X"9A",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"9B",
		X"00",X"00",X"00",X"BC",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"00",X"AB",X"00",X"00",X"00",X"B7",X"00",X"00",X"00",X"31",X"00",X"00",X"00",X"21",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"21",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BA",X"12",X"AB",X"BB",X"BA",X"12",X"BA",X"CC",X"AA",X"12",X"A7",X"CB",X"AA",X"12",X"79",X"BB",
		X"AA",X"41",X"AA",X"BB",X"AA",X"41",X"AA",X"BA",X"9A",X"41",X"AA",X"B7",X"AA",X"41",X"BA",X"AA",
		X"AA",X"A7",X"AB",X"AB",X"AA",X"94",X"BA",X"AA",X"AA",X"94",X"AA",X"AA",X"AB",X"94",X"AA",X"BA",
		X"BA",X"94",X"AA",X"BA",X"BB",X"74",X"BA",X"BA",X"BB",X"AA",X"BA",X"77",X"AA",X"AA",X"BB",X"22",
		X"AA",X"AA",X"BA",X"22",X"AA",X"AA",X"BA",X"12",X"AA",X"99",X"BA",X"12",X"99",X"7A",X"AA",X"12",
		X"99",X"19",X"AA",X"12",X"99",X"A9",X"99",X"12",X"9A",X"99",X"99",X"12",X"AB",X"99",X"99",X"12",
		X"49",X"BA",X"77",X"12",X"17",X"91",X"97",X"22",X"11",X"99",X"77",X"22",X"22",X"9A",X"77",X"22",
		X"22",X"BA",X"77",X"22",X"22",X"77",X"77",X"22",X"22",X"2D",X"47",X"22",X"22",X"22",X"42",X"21",
		X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"12",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"21",
		X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"12",
		X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"32",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"21",
		X"22",X"92",X"42",X"22",X"22",X"72",X"14",X"22",X"12",X"22",X"14",X"22",X"12",X"23",X"47",X"22",
		X"12",X"33",X"45",X"22",X"12",X"22",X"75",X"12",X"42",X"22",X"57",X"42",X"42",X"22",X"77",X"01",
		X"74",X"22",X"E5",X"04",X"17",X"11",X"EE",X"00",X"1C",X"77",X"E5",X"00",X"21",X"55",X"E5",X"00",
		X"22",X"5E",X"75",X"00",X"11",X"5E",X"55",X"00",X"24",X"55",X"55",X"00",X"17",X"55",X"55",X"00",
		X"47",X"55",X"55",X"50",X"77",X"55",X"55",X"50",X"77",X"55",X"E5",X"50",X"45",X"55",X"5E",X"50",
		X"55",X"57",X"55",X"50",X"55",X"47",X"E5",X"50",X"55",X"77",X"EE",X"50",X"55",X"77",X"55",X"50",
		X"55",X"57",X"77",X"50",X"7E",X"77",X"22",X"50",X"27",X"57",X"22",X"50",X"22",X"77",X"22",X"00",
		X"22",X"75",X"22",X"00",X"22",X"75",X"22",X"00",X"21",X"50",X"22",X"00",X"21",X"00",X"22",X"00",
		X"06",X"00",X"D0",X"00",X"FF",X"FF",X"D0",X"00",X"00",X"66",X"D0",X"00",X"00",X"06",X"D0",X"00",
		X"0F",X"06",X"D0",X"00",X"FF",X"00",X"D0",X"00",X"F0",X"00",X"D0",X"00",X"F0",X"00",X"D0",X"00",
		X"F0",X"00",X"D0",X"00",X"F0",X"00",X"D0",X"00",X"FF",X"00",X"DD",X"00",X"6F",X"00",X"00",X"00",
		X"06",X"00",X"00",X"00",X"00",X"06",X"D0",X"00",X"00",X"6F",X"DD",X"00",X"00",X"F0",X"DD",X"00",
		X"F0",X"00",X"C0",X"00",X"6F",X"00",X"DD",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"0D",X"00",
		X"00",X"00",X"DD",X"D0",X"00",X"00",X"D0",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0D",X"00",X"00",X"00",X"0D",X"D0",X"00",X"0D",X"0D",X"D0",X"00",X"D0",X"0D",X"0D",
		X"00",X"00",X"0D",X"0D",X"00",X"00",X"0D",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"0D",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"D0",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0D",X"0D",X"00",X"00",X"D0",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"D0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"33",X"33",X"00",X"03",X"13",X"13",X"00",
		X"03",X"11",X"11",X"00",X"31",X"31",X"31",X"00",X"31",X"31",X"31",X"00",X"11",X"31",X"31",X"00",
		X"31",X"31",X"31",X"00",X"31",X"31",X"31",X"00",X"31",X"31",X"31",X"00",X"31",X"31",X"31",X"00",
		X"31",X"11",X"11",X"00",X"11",X"13",X"13",X"00",X"33",X"33",X"33",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"33",X"00",X"11",X"11",X"31",X"00",
		X"13",X"13",X"11",X"00",X"33",X"13",X"13",X"00",X"30",X"13",X"13",X"00",X"03",X"11",X"13",X"00",
		X"03",X"33",X"13",X"00",X"31",X"00",X"13",X"00",X"31",X"30",X"13",X"00",X"11",X"33",X"13",X"00",
		X"13",X"13",X"11",X"00",X"11",X"11",X"31",X"00",X"33",X"33",X"33",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"33",X"00",X"11",X"31",X"31",X"00",
		X"13",X"11",X"11",X"00",X"13",X"13",X"13",X"00",X"13",X"13",X"13",X"00",X"11",X"13",X"13",X"00",
		X"33",X"13",X"13",X"00",X"00",X"13",X"13",X"00",X"30",X"13",X"13",X"00",X"33",X"13",X"13",X"00",
		X"13",X"11",X"11",X"00",X"11",X"31",X"31",X"00",X"33",X"33",X"33",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"33",X"00",X"11",X"11",X"31",X"00",
		X"11",X"13",X"11",X"00",X"33",X"13",X"13",X"00",X"00",X"13",X"13",X"00",X"00",X"11",X"13",X"00",
		X"03",X"33",X"13",X"00",X"31",X"00",X"13",X"00",X"11",X"30",X"13",X"00",X"11",X"33",X"13",X"00",
		X"11",X"13",X"11",X"00",X"11",X"11",X"31",X"00",X"33",X"33",X"33",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"00",
		X"33",X"33",X"33",X"00",X"31",X"31",X"31",X"00",X"31",X"31",X"31",X"00",X"31",X"31",X"31",X"00",
		X"31",X"31",X"31",X"00",X"31",X"31",X"31",X"00",X"31",X"31",X"31",X"00",X"31",X"31",X"31",X"00",
		X"33",X"33",X"33",X"00",X"33",X"03",X"03",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"30",X"00",X"03",X"33",X"30",X"00",
		X"03",X"33",X"33",X"30",X"03",X"33",X"03",X"30",X"03",X"33",X"03",X"30",X"00",X"33",X"33",X"30",
		X"00",X"33",X"33",X"30",X"00",X"30",X"33",X"30",X"00",X"03",X"33",X"30",X"03",X"33",X"33",X"30",
		X"33",X"33",X"33",X"30",X"33",X"33",X"00",X"00",X"33",X"30",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"03",X"00",X"00",X"00",
		X"33",X"03",X"33",X"30",X"33",X"03",X"33",X"30",X"33",X"03",X"33",X"30",X"33",X"33",X"33",X"30",
		X"33",X"33",X"33",X"30",X"30",X"33",X"33",X"30",X"33",X"33",X"33",X"30",X"33",X"33",X"33",X"30",
		X"33",X"33",X"33",X"30",X"33",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"33",X"33",X"00",X"03",X"23",X"23",X"00",
		X"03",X"22",X"22",X"00",X"32",X"32",X"32",X"00",X"32",X"32",X"32",X"00",X"22",X"32",X"32",X"00",
		X"32",X"32",X"32",X"00",X"32",X"32",X"32",X"00",X"32",X"32",X"32",X"00",X"32",X"32",X"32",X"00",
		X"32",X"22",X"22",X"00",X"22",X"23",X"23",X"00",X"33",X"33",X"33",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"33",X"00",X"22",X"22",X"32",X"00",
		X"23",X"23",X"22",X"00",X"33",X"23",X"23",X"00",X"30",X"23",X"23",X"00",X"03",X"22",X"23",X"00",
		X"03",X"33",X"23",X"00",X"32",X"00",X"23",X"00",X"32",X"30",X"23",X"00",X"22",X"33",X"23",X"00",
		X"23",X"23",X"22",X"00",X"22",X"22",X"32",X"00",X"33",X"33",X"33",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"33",X"00",X"22",X"32",X"32",X"00",
		X"23",X"22",X"22",X"00",X"23",X"23",X"23",X"00",X"23",X"23",X"23",X"00",X"22",X"23",X"23",X"00",
		X"33",X"23",X"23",X"00",X"00",X"23",X"23",X"00",X"30",X"23",X"23",X"00",X"33",X"23",X"23",X"00",
		X"23",X"22",X"22",X"00",X"22",X"32",X"32",X"00",X"33",X"33",X"33",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"33",X"00",X"22",X"22",X"32",X"00",
		X"22",X"23",X"22",X"00",X"33",X"23",X"23",X"00",X"00",X"23",X"23",X"00",X"00",X"22",X"23",X"00",
		X"03",X"33",X"23",X"00",X"32",X"00",X"23",X"00",X"22",X"30",X"23",X"00",X"22",X"33",X"23",X"00",
		X"22",X"23",X"22",X"00",X"22",X"22",X"32",X"00",X"33",X"33",X"33",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"00",
		X"33",X"33",X"33",X"00",X"32",X"32",X"32",X"00",X"32",X"32",X"32",X"00",X"32",X"32",X"32",X"00",
		X"32",X"32",X"32",X"00",X"32",X"32",X"32",X"00",X"32",X"32",X"32",X"00",X"32",X"32",X"32",X"00",
		X"33",X"33",X"33",X"00",X"33",X"03",X"03",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"30",X"00",X"03",X"33",X"30",X"00",
		X"03",X"33",X"33",X"30",X"03",X"33",X"03",X"30",X"03",X"33",X"03",X"30",X"00",X"33",X"33",X"30",
		X"00",X"33",X"33",X"30",X"00",X"30",X"33",X"30",X"00",X"03",X"33",X"30",X"03",X"33",X"33",X"30",
		X"33",X"33",X"33",X"30",X"33",X"33",X"00",X"00",X"33",X"30",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"03",X"00",X"00",X"00",
		X"33",X"03",X"33",X"30",X"33",X"03",X"33",X"30",X"33",X"03",X"33",X"30",X"33",X"33",X"33",X"30",
		X"33",X"33",X"33",X"30",X"30",X"33",X"33",X"30",X"33",X"33",X"33",X"30",X"33",X"33",X"33",X"30",
		X"33",X"33",X"33",X"30",X"33",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
