
module TTL74_257(
	GN,
	SEL,
	B4,
	A4,
	B3,
	A3,
	B2,
	A2,
	B1,
	A1,
	Y4,
	Y3,
	Y2,
	Y1
);


input wire	GN;
input wire	SEL;
input wire	B4;
input wire	A4;
input wire	B3;
input wire	A3;
input wire	B2;
input wire	A2;
input wire	B1;
input wire	A1;
output wire	Y4;
output wire	Y3;
output wire	Y2;
output wire	Y1;

wire	SYNTHESIZED_WIRE_0;
wire	SYNTHESIZED_WIRE_1;
wire	SYNTHESIZED_WIRE_2;
wire	SYNTHESIZED_WIRE_20;
wire	SYNTHESIZED_WIRE_4;
wire	SYNTHESIZED_WIRE_5;
wire	SYNTHESIZED_WIRE_6;
wire	SYNTHESIZED_WIRE_8;
wire	SYNTHESIZED_WIRE_9;
wire	SYNTHESIZED_WIRE_10;
wire	SYNTHESIZED_WIRE_12;
wire	SYNTHESIZED_WIRE_14;
wire	SYNTHESIZED_WIRE_15;
wire	SYNTHESIZED_WIRE_21;




assign	SYNTHESIZED_WIRE_2 = SYNTHESIZED_WIRE_0 | SYNTHESIZED_WIRE_1;

assign	SYNTHESIZED_WIRE_1 = B1 & SEL;

assign	Y1 = SYNTHESIZED_WIRE_20 ? SYNTHESIZED_WIRE_2 : 1'bz;

assign	SYNTHESIZED_WIRE_6 = SYNTHESIZED_WIRE_4 | SYNTHESIZED_WIRE_5;

assign	Y2 = SYNTHESIZED_WIRE_20 ? SYNTHESIZED_WIRE_6 : 1'bz;

assign	SYNTHESIZED_WIRE_10 = SYNTHESIZED_WIRE_8 | SYNTHESIZED_WIRE_9;

assign	Y3 = SYNTHESIZED_WIRE_20 ? SYNTHESIZED_WIRE_10 : 1'bz;

assign	Y4 = SYNTHESIZED_WIRE_20 ? SYNTHESIZED_WIRE_12 : 1'bz;

assign	SYNTHESIZED_WIRE_12 = SYNTHESIZED_WIRE_14 | SYNTHESIZED_WIRE_15;

assign	SYNTHESIZED_WIRE_20 =  ~GN;

assign	SYNTHESIZED_WIRE_21 =  ~SEL;

assign	SYNTHESIZED_WIRE_0 = A1 & SYNTHESIZED_WIRE_21;

assign	SYNTHESIZED_WIRE_4 = A2 & SYNTHESIZED_WIRE_21;

assign	SYNTHESIZED_WIRE_8 = A3 & SYNTHESIZED_WIRE_21;

assign	SYNTHESIZED_WIRE_14 = A4 & SYNTHESIZED_WIRE_21;

assign	SYNTHESIZED_WIRE_5 = B2 & SEL;

assign	SYNTHESIZED_WIRE_9 = B3 & SEL;

assign	SYNTHESIZED_WIRE_15 = B4 & SEL;


endmodule
