library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity travusa_spr_bit1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of travusa_spr_bit1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"7F",X"7F",X"7F",X"7F",X"3E",X"19",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"19",X"3E",X"7F",X"7F",X"7F",X"7F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C1",X"C1",X"C1",X"C1",X"C0",X"C0",X"E0",X"E0",X"E1",X"F7",X"FF",X"FF",X"1F",X"08",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"83",X"03",X"FF",X"FF",X"FC",X"0A",X"00",X"00",
		X"00",X"00",X"08",X"1F",X"FF",X"FF",X"F7",X"E1",X"E0",X"E0",X"C0",X"C0",X"C1",X"C1",X"C1",X"C1",
		X"00",X"00",X"0A",X"FC",X"FF",X"FF",X"03",X"83",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"87",X"87",X"87",X"87",X"87",X"CF",X"FF",X"FF",X"3F",X"F9",X"F8",X"FE",X"3E",X"0C",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"07",X"03",X"03",X"00",X"00",X"00",X"00",X"00",
		X"03",X"01",X"1F",X"0C",X"6D",X"DF",X"CF",X"FF",X"F7",X"E7",X"03",X"00",X"00",X"01",X"01",X"00",
		X"FE",X"BE",X"3C",X"28",X"80",X"C0",X"80",X"03",X"03",X"27",X"7F",X"FF",X"F8",X"FF",X"87",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"FC",X"FE",X"FE",X"FE",X"BA",X"80",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"07",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"BC",X"FE",X"FE",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"07",X"03",X"03",X"00",X"00",X"00",X"00",X"00",
		X"03",X"01",X"1F",X"0C",X"6D",X"DF",X"CF",X"FF",X"F7",X"E7",X"03",X"00",X"00",X"01",X"01",X"00",
		X"FC",X"FC",X"78",X"50",X"80",X"C0",X"80",X"03",X"07",X"0F",X"7F",X"FF",X"F8",X"FF",X"87",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"FC",X"FE",X"FE",X"FE",X"BA",X"80",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"07",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"F8",X"FC",X"FC",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"07",X"07",X"03",X"01",X"03",X"06",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1B",X"3B",X"C9",X"8E",X"FE",X"FC",X"EF",X"EF",X"57",X"11",X"07",X"0F",X"0F",X"1E",X"18",X"00",
		X"A0",X"00",X"00",X"00",X"00",X"00",X"10",X"7E",X"FE",X"FF",X"BF",X"2D",X"C1",X"F0",X"3C",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"3F",X"7F",X"7F",X"7F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"07",X"07",X"03",X"01",X"03",X"06",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"3E",X"CA",X"8E",X"FE",X"FC",X"EF",X"EF",X"57",X"11",X"07",X"0F",X"0F",X"1C",X"19",X"00",
		X"40",X"00",X"00",X"00",X"00",X"00",X"30",X"7E",X"FE",X"FF",X"BF",X"2D",X"C1",X"F0",X"3C",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"3F",X"7F",X"7F",X"7F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"2D",X"7F",X"4C",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"4C",X"7F",X"2D",X"00",
		X"00",X"00",X"80",X"80",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"80",X"80",X"00",X"00",
		X"00",X"12",X"7F",X"33",X"61",X"61",X"61",X"61",X"61",X"61",X"61",X"61",X"33",X"7F",X"12",X"00",
		X"00",X"00",X"80",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"80",X"00",X"00",
		X"01",X"01",X"01",X"01",X"02",X"02",X"03",X"03",X"01",X"01",X"03",X"03",X"01",X"00",X"00",X"00",
		X"E0",X"14",X"3E",X"F6",X"E4",X"04",X"44",X"E0",X"E0",X"E0",X"E0",X"C0",X"80",X"40",X"C0",X"C0",
		X"00",X"01",X"01",X"01",X"02",X"02",X"03",X"03",X"01",X"01",X"03",X"03",X"01",X"00",X"00",X"00",
		X"F0",X"14",X"9E",X"F6",X"E4",X"04",X"44",X"E0",X"E0",X"E0",X"E0",X"C0",X"80",X"40",X"C0",X"C0",
		X"FF",X"FF",X"FF",X"7F",X"0F",X"0C",X"08",X"00",X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"07",X"07",X"03",X"81",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FE",X"FE",X"E1",X"05",X"64",X"7C",X"26",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"26",X"7C",X"64",X"05",X"E1",X"FE",X"FE",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",
		X"FE",X"FE",X"FE",X"E1",X"05",X"64",X"7C",X"26",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"26",X"7C",X"64",X"05",X"E1",X"FE",X"FE",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",
		X"0E",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"0B",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"F8",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"F0",X"F8",X"70",
		X"7F",X"FF",X"FF",X"DB",X"E1",X"30",X"82",X"67",X"7A",X"FC",X"3C",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"37",X"7F",X"7E",X"FF",X"FF",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",
		X"7F",X"FF",X"FF",X"DB",X"E1",X"30",X"82",X"67",X"7A",X"FC",X"3C",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"C0",X"C0",X"80",X"80",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"1F",X"0F",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F8",X"E0",X"80",X"00",X"00",X"60",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"33",X"3F",X"0F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"0F",X"3F",X"33",X"01",
		X"00",X"40",X"80",X"80",X"C0",X"F0",X"80",X"80",X"80",X"80",X"F0",X"C0",X"80",X"80",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"40",X"01",X"40",X"F1",X"E3",X"E3",X"E3",X"E3",X"F1",X"40",X"01",X"40",X"40",X"00",
		X"00",X"00",X"20",X"E0",X"60",X"F0",X"F8",X"E0",X"E0",X"F8",X"F0",X"60",X"E0",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"0E",X"1C",X"3C",X"3C",X"1C",X"0E",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"70",X"30",X"70",X"F0",X"F0",X"70",X"30",X"70",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"0F",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"9C",X"1C",X"38",X"1C",X"9C",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"18",X"30",X"18",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"04",X"00",X"06",X"0F",X"3F",X"7F",X"7F",X"7F",X"7F",X"3F",X"0F",X"06",X"00",X"04",X"04",
		X"00",X"0C",X"0F",X"03",X"8F",X"1E",X"1E",X"1E",X"1F",X"1F",X"0F",X"83",X"0F",X"0C",X"00",X"00",
		X"40",X"C0",X"E0",X"E0",X"F0",X"D0",X"C0",X"C0",X"C0",X"F0",X"F0",X"E0",X"E0",X"60",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"0F",X"0F",X"07",X"01",X"07",X"00",X"00",X"00",
		X"1F",X"1F",X"0F",X"1B",X"13",X"57",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"18",X"1C",X"1C",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"0F",
		X"FC",X"FC",X"FC",X"FC",X"E4",X"C1",X"C1",X"81",X"82",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"C0",X"80",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"70",X"F8",X"C8",X"01",X"01",X"01",X"01",X"F3",X"F9",X"F9",X"FC",
		X"00",X"00",X"00",X"00",X"30",X"78",X"F8",X"FC",X"F8",X"E0",X"E0",X"E0",X"E0",X"C0",X"D0",X"F0",
		X"0F",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"F0",X"F0",X"EC",X"7E",X"5F",X"73",X"7D",X"FF",X"E6",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"0F",X"0F",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"E7",X"FF",
		X"FC",X"FC",X"FE",X"FE",X"7E",X"FE",X"DE",X"8C",X"00",X"00",X"01",X"03",X"07",X"1C",X"38",X"00",
		X"00",X"00",X"00",X"00",X"1E",X"3E",X"FF",X"FF",X"FB",X"F1",X"E0",X"C0",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"E0",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"60",X"20",
		X"7F",X"FF",X"FF",X"7F",X"1F",X"0F",X"07",X"01",X"00",X"00",X"01",X"04",X"06",X"03",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"2E",X"2E",X"2E",X"3E",X"1E",X"1F",X"1F",X"1F",X"0F",X"1E",X"3E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FC",X"F8",X"70",X"06",X"8F",X"FF",X"7F",X"3F",X"1B",X"0C",X"04",X"00",X"00",X"00",X"00",
		X"18",X"30",X"00",X"00",X"00",X"C0",X"E0",X"E0",X"F0",X"F0",X"70",X"78",X"70",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"30",X"F8",X"38",X"00",X"38",X"7C",X"FC",X"FC",X"FE",X"FE",X"FE",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"38",X"38",X"18",
		X"C7",X"CF",X"6F",X"27",X"23",X"30",X"3F",X"3F",X"3F",X"2F",X"2F",X"07",X"01",X"03",X"07",X"0F",
		X"F8",X"F8",X"F0",X"E0",X"86",X"06",X"06",X"0C",X"18",X"80",X"80",X"80",X"80",X"80",X"80",X"00",
		X"00",X"00",X"19",X"3F",X"3F",X"0F",X"0F",X"0F",X"1F",X"1F",X"0F",X"0F",X"07",X"81",X"80",X"80",
		X"7C",X"F8",X"F8",X"F0",X"E0",X"E0",X"B0",X"9C",X"9E",X"8E",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"1E",X"3E",X"7E",X"7C",X"FE",X"FE",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"1B",X"3D",X"7C",X"7C",X"7C",X"7E",X"7F",X"7F",X"3F",X"03",X"01",
		X"E0",X"70",X"38",X"00",X"00",X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"3F",X"37",X"01",
		X"18",X"18",X"18",X"58",X"F8",X"F0",X"F0",X"F0",X"B0",X"B0",X"B0",X"80",X"80",X"E0",X"E0",X"E0",
		X"10",X"10",X"10",X"19",X"0F",X"03",X"87",X"C7",X"E7",X"F7",X"F3",X"FA",X"E8",X"C4",X"C8",X"C0",
		X"20",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F1",X"23",X"03",X"03",X"16",X"1C",X"18",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"41",X"E2",X"E7",X"F7",X"7C",X"08",
		X"00",X"00",X"00",X"00",X"60",X"40",X"C0",X"80",X"82",X"06",X"04",X"CC",X"E8",X"F8",X"D0",X"30",
		X"00",X"00",X"01",X"01",X"03",X"03",X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"C7",X"E3",X"F3",X"F3",X"F3",X"F3",X"F3",X"E7",X"FF",X"1F",X"0E",X"06",X"02",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"E0",X"E0",X"E0",X"31",X"1F",X"0F",X"0F",X"3F",X"7F",
		X"1C",X"0C",X"80",X"80",X"C0",X"60",X"31",X"15",X"1F",X"0E",X"06",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"FE",X"F0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"07",X"0E",X"0C",X"18",X"01",X"07",X"1C",X"70",X"E0",X"20",X"20",X"B0",X"B8",X"BC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"1F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"17",X"07",X"04",X"00",X"00",X"00",X"00",X"00",
		X"2C",X"3E",X"3E",X"3E",X"C7",X"E5",X"E5",X"C6",X"02",X"02",X"02",X"00",X"00",X"00",X"00",X"00",
		X"02",X"02",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"40",X"60",X"20",X"00",X"00",X"00",X"00",
		X"E7",X"E7",X"C7",X"C7",X"C3",X"83",X"83",X"83",X"81",X"C1",X"C1",X"01",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"C0",X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E8",X"F8",X"7C",X"7C",X"36",
		X"03",X"06",X"0C",X"18",X"18",X"11",X"11",X"10",X"18",X"78",X"70",X"18",X"08",X"08",X"6C",X"F6",
		X"00",X"00",X"00",X"00",X"00",X"80",X"A0",X"38",X"38",X"18",X"08",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E1",X"E1",X"E1",X"E0",X"F0",X"FC",X"F8",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"03",X"03",X"1F",X"3F",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"E0",X"E0",X"E0",X"E1",
		X"FF",X"FF",X"FF",X"FF",X"3E",X"CE",X"CF",X"1E",X"FC",X"FC",X"FE",X"47",X"03",X"02",X"00",X"00",
		X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"C0",X"C3",X"80",X"00",X"01",X"03",X"00",X"00",X"18",X"18",X"70",X"F9",X"FF",X"FF",
		X"00",X"00",X"00",X"FC",X"FE",X"FE",X"CE",X"3C",X"70",X"00",X"00",X"00",X"00",X"C0",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"7F",X"7F",X"7F",X"7F",X"3E",X"18",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"18",X"3E",X"7F",X"7F",X"7F",X"7F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C1",X"C1",X"C1",X"C1",X"C0",X"C0",X"E0",X"E0",X"E1",X"F7",X"FF",X"FF",X"1F",X"48",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"83",X"03",X"FF",X"FF",X"FC",X"08",X"00",X"00",
		X"00",X"00",X"48",X"1F",X"FF",X"FF",X"F7",X"E1",X"E0",X"E0",X"C0",X"C0",X"C1",X"C1",X"C1",X"C1",
		X"00",X"00",X"08",X"FC",X"FF",X"FF",X"03",X"83",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"87",X"87",X"87",X"87",X"87",X"CF",X"FF",X"FF",X"3F",X"F9",X"F8",X"FE",X"3E",X"8C",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"00",X"00",X"01",X"03",X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"40",X"00",X"00",X"00",
		X"00",X"00",X"03",X"07",X"0F",X"00",X"00",X"00",X"60",X"20",X"20",X"20",X"20",X"60",X"60",X"60",
		X"00",X"00",X"80",X"C0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FF",X"9F",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",X"F7",X"E1",X"F8",X"FE",X"3F",X"0F",X"03",X"00",X"00",
		X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",
		X"C0",X"FC",X"FF",X"FF",X"F7",X"E3",X"C3",X"C1",X"81",X"81",X"03",X"03",X"07",X"07",X"07",X"0F",
		X"FC",X"FC",X"F8",X"F8",X"F8",X"FC",X"7C",X"67",X"FF",X"FF",X"FF",X"3F",X"0F",X"07",X"03",X"00",
		X"3C",X"3C",X"3C",X"78",X"78",X"78",X"F8",X"F0",X"F8",X"F0",X"20",X"20",X"C0",X"80",X"00",X"00",
		X"C0",X"F8",X"FE",X"3F",X"0F",X"C7",X"F7",X"FE",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",
		X"00",X"00",X"00",X"80",X"F8",X"FC",X"FC",X"70",X"F2",X"FE",X"FE",X"1E",X"1E",X"1F",X"1E",X"1C",
		X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"03",X"07",X"07",X"03",X"03",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"1F",X"10",X"10",X"00",
		X"01",X"03",X"03",X"07",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"07",X"03",X"03",
		X"FF",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"7F",X"7F",X"C7",X"80",X"80",X"00",X"00",X"80",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"06",X"07",X"07",X"03",X"03",X"03",X"01",X"01",X"01",
		X"00",X"00",X"10",X"10",X"3F",X"FF",X"7F",X"7F",X"F0",X"E0",X"E0",X"E0",X"B0",X"BF",X"BF",X"FF",
		X"F8",X"F8",X"F8",X"FC",X"7F",X"79",X"60",X"30",X"18",X"0F",X"07",X"03",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"DF",X"FF",X"3F",X"1E",X"FC",X"F1",X"FB",X"7F",X"7C",X"00",X"00",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0F",X"1F",X"3F",X"7F",X"7F",X"FF",X"FE",X"F8",
		X"04",X"0E",X"00",X"02",X"07",X"3F",X"FF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"9F",X"0F",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"EF",X"66",X"F1",X"FF",X"FF",X"FE",X"60",X"00",X"00",
		X"88",X"F8",X"F8",X"F8",X"F8",X"98",X"98",X"F8",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"08",X"08",X"08",X"08",X"08",X"08",
		X"00",X"3F",X"FF",X"6F",X"EF",X"E6",X"F1",X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"FE",X"FE",X"FE",
		X"38",X"FC",X"F8",X"F8",X"98",X"98",X"F8",X"F8",X"18",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"F0",X"F8",X"CE",X"47",X"61",X"3F",X"1F",X"0F",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"03",X"0F",X"3F",X"7F",X"FF",X"FF",X"FD",X"F0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"CC",X"1E",X"3F",X"CF",X"00",
		X"87",X"80",X"80",X"80",X"C0",X"E0",X"F8",X"F8",X"F8",X"E8",X"E8",X"B0",X"70",X"E0",X"80",X"00",
		X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"A8",X"78",X"C8",X"80",X"80",X"00",X"00",X"80",X"80",X"87",X"87",X"87",X"87",X"87",X"87",X"87",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C7",X"1F",X"0D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"FC",X"F8",X"E8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0F",X"0F",X"04",X"06",X"03",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"0F",X"0F",X"0E",X"0E",X"0E",X"0E",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"DF",X"7F",X"3B",X"F7",X"E7",X"7F",X"00",X"00",
		X"C3",X"C3",X"C3",X"C0",X"C0",X"C0",X"E0",X"F8",X"F8",X"E8",X"E8",X"F8",X"F0",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"19",X"07",X"1B",X"7F",X"FF",X"FF",X"FF",X"FF",X"9F",X"1F",X"1F",X"1F",X"1F",
		X"00",X"00",X"18",X"FC",X"F8",X"E8",X"E8",X"F8",X"E0",X"C0",X"80",X"C0",X"C0",X"C3",X"C3",X"C3",
		X"33",X"73",X"73",X"73",X"73",X"73",X"73",X"73",X"7B",X"7F",X"27",X"31",X"1F",X"07",X"00",X"00",
		X"F0",X"F3",X"F3",X"F3",X"F3",X"F3",X"F0",X"FC",X"FC",X"F8",X"FC",X"FC",X"F8",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"1F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"FC",X"F8",X"FC",X"F0",
		X"00",X"00",X"01",X"03",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"03",X"01",X"00",X"00",
		X"1C",X"7E",X"FC",X"3E",X"3C",X"38",X"39",X"39",X"39",X"39",X"38",X"3C",X"3E",X"FC",X"7E",X"1C",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"1C",X"7E",X"DE",X"9C",X"98",X"99",X"99",X"98",X"9C",X"DE",X"7E",X"1C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0E",X"1E",X"36",X"34",X"34",X"34",X"34",X"36",X"1E",X"06",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"0A",X"0A",X"0A",X"0A",X"06",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"80",X"C0",X"40",X"4C",X"4F",X"6F",X"6F",X"2F",X"2F",X"07",X"03",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"0C",X"0E",X"CF",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"7F",X"E7",X"FF",X"FE",X"FC",X"00",X"00",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"CF",X"0E",X"0C",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"00",X"00",X"FC",X"FE",X"FF",X"E7",X"7F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"E0",X"E0",X"E0",X"FF",X"FF",X"FF",X"E0",X"60",X"60",X"7F",X"7F",X"7F",X"70",X"FE",X"FE",X"7F",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"80",
		X"7F",X"FF",X"FF",X"7F",X"60",X"60",X"60",X"7F",X"7F",X"FF",X"E0",X"E0",X"E0",X"FF",X"FF",X"FF",
		X"80",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"03",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FE",
		X"03",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",
		X"FE",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"1C",X"3E",X"63",X"5D",X"5D",X"5D",X"5D",X"63",X"3E",X"1C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"1C",X"3E",X"7F",X"7D",X"41",X"41",X"6D",X"7F",X"3E",X"1E",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"1C",X"3E",X"65",X"45",X"51",X"59",X"49",X"6D",X"3E",X"1C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"1C",X"3E",X"6B",X"41",X"55",X"5D",X"49",X"6B",X"3E",X"1C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"1C",X"3E",X"7B",X"41",X"41",X"4B",X"63",X"73",X"3E",X"1C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"1C",X"3E",X"73",X"51",X"55",X"45",X"45",X"7F",X"3E",X"1C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"1C",X"3E",X"7B",X"51",X"55",X"55",X"41",X"63",X"3E",X"1C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"1E",X"3E",X"4F",X"47",X"51",X"59",X"5F",X"4F",X"3E",X"1C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"1C",X"3E",X"6B",X"51",X"55",X"55",X"45",X"6B",X"3E",X"1C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"1C",X"3E",X"63",X"41",X"55",X"55",X"45",X"6F",X"3E",X"1C",X"00",X"00",X"00",
		X"07",X"0C",X"1B",X"1B",X"1B",X"0C",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"30",X"D8",X"D8",X"D8",X"30",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"0C",X"1E",X"1E",X"1E",X"0E",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"38",X"78",X"78",X"38",X"70",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"08",X"1E",X"18",X"19",X"0C",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"10",X"38",X"F8",X"98",X"30",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"0C",X"19",X"1C",X"19",X"0C",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"30",X"98",X"F8",X"98",X"30",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"0C",X"18",X"1C",X"1C",X"0C",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"F0",X"18",X"98",X"38",X"70",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"0C",X"19",X"18",X"1F",X"0C",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"30",X"F8",X"38",X"38",X"30",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"0C",X"19",X"1C",X"1F",X"0C",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"30",X"98",X"18",X"98",X"30",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"1E",X"1E",X"1C",X"19",X"08",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"70",X"78",X"F8",X"D8",X"10",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"0C",X"19",X"1C",X"1B",X"0C",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"30",X"D8",X"38",X"98",X"30",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"0C",X"19",X"18",X"19",X"0C",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"30",X"F8",X"38",X"98",X"30",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"14",X"5C",X"0F",X"1B",X"77",X"94",X"20",X"84",X"10",X"42",X"90",X"05",X"20",X"0A",X"00",
		X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"80",X"12",X"40",X"08",X"21",X"00",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"20",X"05",X"90",X"42",X"10",X"84",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"21",X"08",X"40",X"12",X"80",X"00",
		X"20",X"68",X"F0",X"90",X"18",X"98",X"F0",X"50",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"1F",X"3F",X"7F",X"7F",X"E0",X"E0",X"E0",X"F0",X"FF",X"7F",X"7F",X"3F",
		X"00",X"00",X"00",X"00",X"F0",X"F8",X"F8",X"FC",X"3C",X"1C",X"1C",X"1C",X"F8",X"F8",X"F0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"FF",X"FF",X"7F",X"30",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"FC",X"FC",X"F8",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"1E",X"3F",X"7F",X"FF",X"E7",X"E3",X"E3",X"F1",X"F9",X"F8",X"78",X"30",
		X"00",X"00",X"00",X"00",X"0C",X"1C",X"9C",X"9C",X"DC",X"DC",X"FC",X"FC",X"FC",X"FC",X"7C",X"18",
		X"00",X"00",X"00",X"00",X"1C",X"3E",X"7F",X"FF",X"EF",X"E7",X"E7",X"F6",X"F8",X"F8",X"78",X"30",
		X"00",X"00",X"00",X"00",X"70",X"F8",X"FC",X"FC",X"3C",X"1C",X"1C",X"1C",X"3C",X"78",X"70",X"60",
		X"02",X"82",X"92",X"92",X"92",X"FE",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"F8",X"88",X"88",X"88",X"FE",X"FE",X"00",X"FE",X"FE",X"70",X"38",X"70",X"FE",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"E0",X"F0",X"1E",X"1E",X"F0",X"E0",X"00",X"00",X"80",X"80",X"FE",X"FE",X"80",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"1F",X"1F",X"3F",X"3F",X"3F",X"3F",X"1F",X"3F",X"3F",X"3F",X"1F",X"07",X"07",X"03",X"01",
		X"6C",X"7E",X"FE",X"FE",X"FC",X"FC",X"FE",X"FF",X"FF",X"FF",X"FE",X"FC",X"FC",X"FC",X"F8",X"B0",
		X"E0",X"F8",X"FE",X"FF",X"FF",X"E7",X"40",X"00",X"40",X"E7",X"FF",X"FF",X"FE",X"F8",X"E0",X"40",
		X"00",X"00",X"00",X"80",X"E0",X"F8",X"FE",X"3F",X"FE",X"F8",X"E0",X"80",X"00",X"00",X"00",X"00",
		X"40",X"00",X"40",X"E7",X"FF",X"FF",X"FE",X"F8",X"E0",X"40",X"E0",X"FF",X"FF",X"FF",X"E0",X"40",
		X"FE",X"3F",X"FE",X"F8",X"E0",X"80",X"00",X"00",X"00",X"02",X"07",X"FF",X"FF",X"FF",X"07",X"02",
		X"00",X"00",X"01",X"07",X"1F",X"7F",X"FC",X"7F",X"1F",X"47",X"E1",X"F8",X"FE",X"FF",X"FF",X"E7",
		X"1F",X"7F",X"FF",X"FF",X"F7",X"72",X"70",X"72",X"F7",X"FF",X"FF",X"7F",X"1F",X"87",X"E2",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"78",X"FF",X"FF",X"FF",X"78",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"0F",X"CF",X"0F",X"06",X"00",X"02",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"1F",X"1F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"18",X"38",X"38",X"10",X"30",X"EF",X"FE",X"FE",X"FE",X"FE",X"EF",X"30",X"10",X"38",X"38",X"18",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"1F",X"3F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"18",X"38",X"38",X"10",X"30",X"EF",X"FE",X"FE",X"FE",X"FE",X"EF",X"30",X"10",X"38",X"38",X"18",
		X"00",X"00",X"00",X"18",X"3C",X"7E",X"FE",X"FE",X"FE",X"FE",X"7E",X"3C",X"18",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"7C",X"7F",X"7F",X"7F",X"7F",X"7C",X"00",X"00",X"00",X"00",X"00",
		X"0D",X"1F",X"1F",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"EE",X"FE",X"FE",X"FE",X"7E",X"7F",X"7F",X"73",X"30",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7C",X"FC",X"FE",X"FE",X"7E",X"3E",X"FC",X"FC",X"18",X"01",X"03",X"3F",X"70",X"70",X"E0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"7E",X"FF",X"FF",X"FF",X"FD",X"FC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F7",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"07",X"07",X"03",X"09",X"03",X"06",
		X"00",X"00",X"00",X"00",X"00",X"06",X"0E",X"2E",X"7C",X"78",X"F8",X"F7",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"8C",X"00",X"00",X"81",X"07",X"1F",X"3F",X"7B",X"38",X"70",X"60",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"FE",X"FE",X"FF",X"FF",X"FB",X"FD",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"7E",X"7E",X"7F",X"3F",X"9F",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"17",X"07",X"03",X"01",X"03",X"06",
		X"00",X"00",X"00",X"00",X"00",X"06",X"0E",X"2E",X"7C",X"78",X"F8",X"F7",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"1F",X"3F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"18",X"38",X"38",X"10",X"30",X"ED",X"FB",X"FB",X"FB",X"FB",X"ED",X"30",X"10",X"38",X"38",X"18",
		X"00",X"00",X"00",X"30",X"78",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"78",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"7C",X"7F",X"7F",X"7F",X"7F",X"7C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"1F",X"5F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"18",X"38",X"38",X"10",X"30",X"ED",X"FB",X"FB",X"FB",X"FB",X"ED",X"30",X"10",X"38",X"38",X"18",
		X"00",X"00",X"00",X"30",X"7C",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"7C",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"7C",X"7F",X"7F",X"7F",X"7F",X"7C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"0F",X"1F",X"1F",X"0F",X"01",X"07",X"0C",X"00",
		X"00",X"18",X"39",X"3B",X"33",X"A3",X"E1",X"EC",X"FF",X"FF",X"FF",X"FF",X"FF",X"3E",X"38",X"18",
		X"00",X"00",X"F0",X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",X"FC",X"D8",X"80",X"00",X"01",X"0F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1E",X"7F",X"7F",X"7F",X"F9",X"F0",X"FC",X"FC",
		X"38",X"70",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"13",X"06",X"0C",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"D8",X"CE",X"47",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"0D",X"1F",X"1F",X"4F",
		X"00",X"00",X"00",X"00",X"00",X"19",X"3B",X"3F",X"B3",X"E1",X"E4",X"EF",X"FF",X"FF",X"FF",X"F9",
		X"00",X"00",X"01",X"07",X"3F",X"3F",X"78",X"38",X"70",X"60",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"FB",X"F1",X"C0",X"FC",X"FC",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"F8",X"FC",X"FE",X"FE",X"FE",X"FE",X"DC",X"8C",X"88",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7E",X"7E",X"7F",
		X"03",X"26",X"0C",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"D8",X"CE",X"47",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"0D",X"1F",X"3F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"19",X"3B",X"3B",X"B3",X"E1",X"E4",X"EF",X"FF",X"FF",X"FF",X"F9",
		X"00",X"00",X"01",X"07",X"3F",X"3F",X"78",X"38",X"70",X"60",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"FB",X"F1",X"C0",X"FC",X"FC",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"DE",X"8E",X"8C",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7E",X"7E",X"7F",
		X"00",X"00",X"00",X"07",X"07",X"0F",X"1F",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"11",X"31",X"FD",X"FF",X"FF",X"FF",X"FF",X"FD",X"31",X"11",X"30",X"30",X"10",X"00",X"00",
		X"00",X"00",X"E0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FC",X"FF",X"FF",X"FF",X"FF",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"38",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"0F",X"1F",X"5F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"38",X"12",X"33",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"33",X"12",X"38",X"38",X"18",X"00",X"00",
		X"00",X"00",X"C0",X"E0",X"F0",X"F0",X"F0",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FC",X"FF",X"FF",X"FF",X"FF",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"38",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"0F",X"1F",X"1F",X"0F",X"01",X"07",X"0C",X"00",X"00",X"00",X"00",
		X"3F",X"3F",X"BF",X"FF",X"DF",X"CF",X"FF",X"FE",X"FC",X"DE",X"7E",X"38",X"18",X"00",X"00",X"00",
		X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F1",X"61",X"43",X"07",X"1F",X"3F",X"1C",X"38",X"30",X"00",
		X"00",X"00",X"00",X"00",X"3E",X"FF",X"FF",X"FF",X"F9",X"F0",X"FC",X"FC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"3B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"07",X"0F",X"0F",X"17",X"01",X"01",X"03",X"06",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"DF",X"CF",X"FF",X"F6",X"E4",X"E2",X"61",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"E0",X"70",X"61",X"01",X"03",X"04",X"1F",X"1F",X"3C",X"1C",X"38",X"30",
		X"00",X"00",X"1E",X"FE",X"FF",X"FF",X"FB",X"C1",X"40",X"7C",X"FC",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"3B",X"3F",X"BF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"F0",
		X"01",X"01",X"01",X"01",X"0F",X"1F",X"1F",X"0F",X"41",X"03",X"06",X"0C",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"DF",X"CF",X"FF",X"FF",X"FE",X"99",X"C0",X"C0",X"40",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"F8",X"F8",X"F8",X"F0",X"30",X"21",X"01",X"03",X"04",X"1F",X"1F",X"3C",X"1C",X"38",X"30",
		X"00",X"00",X"1E",X"FF",X"FF",X"FF",X"F9",X"C0",X"40",X"7C",X"FC",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"39",X"3D",X"BF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"F0",X"F8",
		X"00",X"00",X"00",X"00",X"0C",X"1F",X"1F",X"0F",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"1C",X"14",X"10",X"BB",X"FF",X"FE",X"FE",X"DE",X"CE",X"60",X"20",X"70",X"70",X"30",X"00",
		X"00",X"00",X"00",X"18",X"3C",X"7E",X"FE",X"FE",X"FE",X"FE",X"7E",X"3C",X"18",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"7C",X"7E",X"7F",X"7F",X"7F",X"7D",X"FC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"5B",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0F",X"2F",X"07",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"1C",X"3C",X"78",X"78",X"F8",X"F7",X"EF",X"3F",X"FF",X"FF",
		X"FE",X"CC",X"80",X"00",X"01",X"07",X"1F",X"1F",X"7B",X"38",X"70",X"60",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"FE",X"FE",X"FF",X"FF",X"FB",X"FD",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"7E",X"7E",X"7F",X"3F",X"9F",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1D",X"1C",X"0C",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"1F",X"07",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"18",X"1C",X"1C",X"1D",
		X"7F",X"7F",X"6F",X"6F",X"6D",X"6D",X"2F",X"4F",X"67",X"73",X"73",X"37",X"5F",X"7F",X"7F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"47",X"63",X"70",X"78",X"3C",X"1C",X"6E",X"77",X"7F",X"7F",X"1F",X"43",X"60",X"78",X"7C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"78",X"7C",X"7E",X"3F",X"1F",X"47",X"63",X"78",X"7C",X"7D",X"7D",X"6D",X"6D",X"7D",X"7D",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"6F",X"6D",X"6D",X"6F",X"6F",X"6F",X"6F",X"7D",X"7D",X"3D",X"5D",X"65",X"71",X"70",X"30",X"58",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"0C",X"0F",X"4F",X"6F",X"7F",X"7D",X"7D",X"7F",X"6F",X"6F",X"7F",X"7D",X"3F",X"1F",X"4F",
		X"F0",X"90",X"80",X"80",X"E0",X"F0",X"F0",X"F0",X"F0",X"90",X"80",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"98",X"9E",X"9F",X"9F",X"8F",X"97",X"91",X"80",X"80",X"80",X"80",X"80",X"C0",X"F0",X"F0",
		X"1F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"1F",X"07",X"03",X"00",X"00",X"00",
		X"9F",X"9F",X"8F",X"87",X"01",X"00",X"10",X"18",X"1E",X"9F",X"9F",X"8F",X"87",X"01",X"00",X"00",
		X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",X"23",X"03",X"03",X"03",X"C0",X"E0",X"F8",X"FD",X"FF",X"3F",
		X"00",X"00",X"00",X"90",X"98",X"9C",X"9C",X"9C",X"1C",X"1C",X"9C",X"9C",X"9C",X"9C",X"9C",X"9E",
		X"FF",X"7F",X"3F",X"1F",X"0F",X"07",X"03",X"C1",X"E0",X"F8",X"FC",X"FF",X"FF",X"FF",X"E7",X"E3",
		X"E0",X"F0",X"F3",X"F3",X"B3",X"BB",X"BF",X"BF",X"9F",X"9F",X"9F",X"9F",X"8F",X"87",X"03",X"01",
		X"00",X"00",X"00",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"80",X"A0",X"B0",X"B0",X"B0",X"B0",X"B0",X"F0",X"F0",X"F0",X"F0",X"90",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"90",X"80",X"80",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"A0",X"80",X"80",X"40",X"D0",X"D0",X"D0",X"D0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"B0",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"80",X"80",X"80",X"80",X"C0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"39",X"38",X"38",X"38",X"18",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E7",X"F7",X"F7",X"7F",X"3F",X"3F",X"1F",X"0F",X"0F",X"07",X"03",X"03",X"01",X"00",X"00",X"00",
		X"00",X"0C",X"0E",X"0E",X"2E",X"32",X"30",X"38",X"3C",X"3C",X"3E",X"3F",X"3F",X"3F",X"3B",X"3B",
		X"FB",X"7F",X"3F",X"8F",X"C7",X"F1",X"F8",X"7E",X"3F",X"0F",X"07",X"01",X"06",X"87",X"C7",X"C7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"CF",X"C7",X"F3",X"FB",X"7F",X"3F",X"8F",X"C7",X"F1",X"F8",X"FE",X"FF",X"CF",X"C7",X"F3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"E0",X"F0",X"78",X"38",X"1C",X"EE",X"FF",X"FF",X"FF",X"0F",X"80",X"C0",X"F0",X"F8",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E6",X"E7",X"E7",X"E3",X"E0",X"E0",X"E0",X"60",X"60",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"06",X"06",X"C6",X"E6",X"F6",X"F6",X"36",X"1E",X"0E",X"0E",X"0E",X"06",X"06",X"26",X"E6",
		X"FF",X"7F",X"3F",X"0F",X"07",X"01",X"00",X"00",X"40",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"0E",X"06",X"06",X"06",X"06",X"06",X"06",X"C6",X"E6",X"F6",X"F6",X"36",X"16",X"06",X"06",X"06",
		X"03",X"03",X"03",X"83",X"C3",X"F1",X"F8",X"FE",X"FF",X"FF",X"EF",X"E7",X"E7",X"E7",X"F7",X"FF",
		X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"86",X"C6",X"E6",X"F6",X"78",X"3C",X"1C",X"0E",
		X"C3",X"C3",X"C3",X"C3",X"43",X"03",X"03",X"03",X"03",X"01",X"00",X"02",X"03",X"03",X"03",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"06",X"06",X"06",X"06",
		X"00",X"00",X"00",X"02",X"03",X"03",X"03",X"03",X"03",X"83",X"C3",X"C3",X"C3",X"C1",X"C0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"3F",X"FF",X"FF",X"FF",X"FF",X"FC",X"3C",X"1C",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"7C",X"7C",X"6C",X"6C",X"7C",X"7C",X"3C",X"18",X"00",X"60",X"FC",X"FC",X"FC",X"FC",X"9C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"F7",X"E3",X"FB",X"FD",X"7D",X"3F",X"DF",X"EF",X"FF",X"FC",X"3C",X"1F",X"C7",X"E3",X"F8",
		X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"80",X"80",X"80",
		X"40",X"60",X"78",X"7C",X"7D",X"FD",X"ED",X"ED",X"FD",X"7D",X"7F",X"FF",X"EF",X"FF",X"FC",X"7C",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
