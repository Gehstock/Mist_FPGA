-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

entity GALAXIAN_1H is
  port (
    CLK         : in    std_logic;
    ADDR        : in    std_logic_vector(11 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of GALAXIAN_1H is


  type ROM_ARRAY is array(0 to 4095) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"38",x"7C",x"C2",x"82",x"86",x"7C",x"38",x"00", -- 0x0000
    x"02",x"02",x"FE",x"FE",x"42",x"02",x"00",x"00", -- 0x0008
    x"62",x"F2",x"BA",x"9A",x"9E",x"CE",x"46",x"00", -- 0x0010
    x"8C",x"DE",x"F2",x"B2",x"92",x"86",x"04",x"00", -- 0x0018
    x"08",x"FE",x"FE",x"C8",x"68",x"38",x"18",x"00", -- 0x0020
    x"1C",x"BE",x"A2",x"A2",x"A2",x"E6",x"E4",x"00", -- 0x0028
    x"0C",x"9E",x"92",x"92",x"D2",x"7E",x"3C",x"00", -- 0x0030
    x"C0",x"E0",x"B0",x"9E",x"8E",x"C0",x"C0",x"00", -- 0x0038
    x"0C",x"6E",x"9A",x"9A",x"B2",x"F2",x"6C",x"00", -- 0x0040
    x"78",x"FC",x"96",x"92",x"92",x"F2",x"60",x"00", -- 0x0048
    x"1C",x"02",x"3C",x"3D",x"14",x"10",x"00",x"00", -- 0x0050
    x"00",x"00",x"00",x"00",x"00",x"60",x"C0",x"00", -- 0x0058
    x"38",x"48",x"1E",x"3E",x"3E",x"1E",x"3C",x"30", -- 0x0060
    x"00",x"00",x"00",x"30",x"10",x"08",x"00",x"00", -- 0x0068
    x"02",x"06",x"04",x"00",x"00",x"00",x"00",x"00", -- 0x0070
    x"00",x"00",x"38",x"1C",x"70",x"30",x"34",x"18", -- 0x0078
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0080
    x"3E",x"7E",x"C8",x"88",x"C8",x"7E",x"3E",x"00", -- 0x0088
    x"6C",x"FE",x"92",x"92",x"92",x"FE",x"FE",x"00", -- 0x0090
    x"44",x"C6",x"82",x"82",x"C6",x"7C",x"38",x"00", -- 0x0098
    x"38",x"7C",x"C6",x"82",x"82",x"FE",x"FE",x"00", -- 0x00A0
    x"82",x"92",x"92",x"92",x"FE",x"FE",x"00",x"00", -- 0x00A8
    x"80",x"90",x"90",x"90",x"90",x"FE",x"FE",x"00", -- 0x00B0
    x"9E",x"9E",x"92",x"82",x"C6",x"7C",x"38",x"00", -- 0x00B8
    x"FE",x"FE",x"10",x"10",x"10",x"FE",x"FE",x"00", -- 0x00C0
    x"82",x"82",x"FE",x"FE",x"82",x"82",x"00",x"00", -- 0x00C8
    x"FC",x"FE",x"02",x"02",x"02",x"06",x"04",x"00", -- 0x00D0
    x"82",x"C6",x"6E",x"3C",x"18",x"FE",x"FE",x"00", -- 0x00D8
    x"02",x"02",x"02",x"02",x"FE",x"FE",x"00",x"00", -- 0x00E0
    x"FE",x"FE",x"70",x"38",x"70",x"FE",x"FE",x"00", -- 0x00E8
    x"FE",x"FE",x"1C",x"38",x"70",x"FE",x"FE",x"00", -- 0x00F0
    x"7C",x"FE",x"82",x"82",x"82",x"FE",x"7C",x"00", -- 0x00F8
    x"70",x"F8",x"88",x"88",x"88",x"FE",x"FE",x"00", -- 0x0100
    x"7A",x"FC",x"8E",x"8A",x"82",x"FE",x"7C",x"00", -- 0x0108
    x"72",x"F6",x"9E",x"8C",x"88",x"FE",x"FE",x"00", -- 0x0110
    x"0C",x"5E",x"D2",x"92",x"92",x"F6",x"64",x"00", -- 0x0118
    x"80",x"80",x"FE",x"FE",x"80",x"80",x"00",x"00", -- 0x0120
    x"FC",x"FE",x"02",x"02",x"02",x"FE",x"FC",x"00", -- 0x0128
    x"F0",x"F8",x"1C",x"0E",x"1C",x"F8",x"F0",x"00", -- 0x0130
    x"F8",x"FE",x"1C",x"38",x"1C",x"FE",x"F8",x"00", -- 0x0138
    x"C6",x"EE",x"7C",x"38",x"7C",x"EE",x"C6",x"00", -- 0x0140
    x"C0",x"F0",x"1E",x"1E",x"F0",x"C0",x"00",x"00", -- 0x0148
    x"C2",x"E2",x"F2",x"BA",x"9E",x"8E",x"86",x"00", -- 0x0150
    x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00", -- 0x0158
    x"00",x"00",x"00",x"00",x"00",x"04",x"00",x"00", -- 0x0160
    x"00",x"00",x"00",x"00",x"00",x"40",x"00",x"00", -- 0x0168
    x"00",x"01",x"00",x"01",x"00",x"00",x"00",x"00", -- 0x0170
    x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0178
    x"00",x"00",x"00",x"00",x"00",x"04",x"00",x"09", -- 0x0180
    x"00",x"00",x"00",x"00",x"00",x"40",x"00",x"00", -- 0x0188
    x"00",x"00",x"04",x"00",x"01",x"00",x"00",x"00", -- 0x0190
    x"10",x"80",x"40",x"00",x"00",x"00",x"00",x"00", -- 0x0198
    x"00",x"00",x"00",x"01",x"08",x"00",x"00",x"00", -- 0x01A0
    x"00",x"00",x"00",x"40",x"00",x"00",x"00",x"00", -- 0x01A8
    x"11",x"04",x"00",x"00",x"08",x"00",x"00",x"00", -- 0x01B0
    x"20",x"00",x"00",x"00",x"00",x"20",x"00",x"00", -- 0x01B8
    x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00", -- 0x01C0
    x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00", -- 0x01C8
    x"08",x"00",x"01",x"00",x"00",x"04",x"00",x"00", -- 0x01D0
    x"88",x"00",x"00",x"10",x"00",x"00",x"00",x"00", -- 0x01D8
    x"00",x"03",x"00",x"01",x"00",x"00",x"00",x"00", -- 0x01E0
    x"00",x"00",x"00",x"80",x"00",x"C0",x"00",x"60", -- 0x01E8
    x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"03", -- 0x01F0
    x"00",x"60",x"00",x"C0",x"00",x"80",x"00",x"00", -- 0x01F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0200
    x"00",x"00",x"00",x"00",x"00",x"60",x"00",x"60", -- 0x0208
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0210
    x"00",x"60",x"00",x"60",x"00",x"00",x"00",x"00", -- 0x0218
    x"10",x"02",x"00",x"20",x"00",x"00",x"40",x"00", -- 0x0220
    x"00",x"10",x"02",x"40",x"00",x"00",x"04",x"00", -- 0x0228
    x"00",x"40",x"10",x"04",x"00",x"80",x"02",x"20", -- 0x0230
    x"00",x"08",x"80",x"00",x"01",x"00",x"20",x"00", -- 0x0238
    x"00",x"20",x"58",x"48",x"24",x"19",x"01",x"00", -- 0x0240
    x"00",x"04",x"08",x"10",x"12",x"0C",x"A0",x"38", -- 0x0248
    x"00",x"01",x"19",x"24",x"48",x"58",x"20",x"00", -- 0x0250
    x"38",x"A0",x"0C",x"12",x"10",x"08",x"04",x"00", -- 0x0258
    x"00",x"02",x"20",x"10",x"00",x"02",x"46",x"00", -- 0x0260
    x"00",x"40",x"04",x"08",x"00",x"60",x"62",x"80", -- 0x0268
    x"00",x"46",x"02",x"00",x"10",x"20",x"02",x"00", -- 0x0270
    x"80",x"62",x"60",x"00",x"08",x"04",x"40",x"00", -- 0x0278
    x"00",x"18",x"34",x"34",x"14",x"08",x"09",x"00", -- 0x0280
    x"00",x"00",x"00",x"0E",x"10",x"08",x"26",x"30", -- 0x0288
    x"00",x"09",x"08",x"14",x"34",x"34",x"18",x"00", -- 0x0290
    x"30",x"26",x"08",x"10",x"0E",x"00",x"00",x"00", -- 0x0298
    x"00",x"08",x"1C",x"1E",x"1E",x"0E",x"06",x"00", -- 0x02A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02A8
    x"00",x"06",x"0E",x"1E",x"1E",x"1C",x"08",x"00", -- 0x02B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02B8
    x"00",x"08",x"1C",x"1E",x"1E",x"0E",x"06",x"00", -- 0x02C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02C8
    x"00",x"06",x"0E",x"1E",x"1E",x"1C",x"08",x"00", -- 0x02D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02D8
    x"00",x"08",x"1C",x"1E",x"1E",x"0E",x"06",x"00", -- 0x02E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02E8
    x"00",x"06",x"0E",x"1E",x"1E",x"1C",x"08",x"00", -- 0x02F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02F8
    x"00",x"00",x"00",x"01",x"03",x"1C",x"23",x"C0", -- 0x0300
    x"00",x"7E",x"FC",x"08",x"F1",x"13",x"FF",x"0F", -- 0x0308
    x"23",x"1C",x"03",x"01",x"00",x"00",x"00",x"00", -- 0x0310
    x"FF",x"13",x"F1",x"08",x"FC",x"7E",x"00",x"00", -- 0x0318
    x"1C",x"38",x"C2",x"06",x"C2",x"38",x"1C",x"00", -- 0x0320
    x"C3",x"C3",x"C3",x"C3",x"C3",x"C3",x"C3",x"C3", -- 0x0328
    x"C3",x"C3",x"C3",x"C3",x"C3",x"C3",x"FF",x"FF", -- 0x0330
    x"C3",x"C3",x"C3",x"C3",x"FF",x"FF",x"FF",x"FF", -- 0x0338
    x"C3",x"C3",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0340
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0348
    x"1F",x"C6",x"F2",x"1D",x"03",x"00",x"00",x"00", -- 0x0350
    x"CC",x"E0",x"80",x"40",x"98",x"F0",x"00",x"00", -- 0x0358
    x"03",x"06",x"0D",x"1E",x"F9",x"06",x"1C",x"FF", -- 0x0360
    x"60",x"FE",x"1F",x"61",x"70",x"F8",x"0C",x"E6", -- 0x0368
    x"06",x"D3",x"FC",x"3B",x"1D",x"0C",x"04",x"00", -- 0x0370
    x"0F",x"78",x"A0",x"18",x"C7",x"3E",x"0C",x"00", -- 0x0378
    x"00",x"01",x"03",x"07",x"03",x"07",x"0F",x"3F", -- 0x0380
    x"80",x"80",x"D8",x"F8",x"F8",x"F0",x"F0",x"F0", -- 0x0388
    x"1F",x"1F",x"1F",x"0F",x"03",x"07",x"07",x"01", -- 0x0390
    x"F8",x"F8",x"F0",x"E0",x"F8",x"FC",x"78",x"00", -- 0x0398
    x"00",x"00",x"00",x"00",x"00",x"04",x"01",x"03", -- 0x03A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"90", -- 0x03A8
    x"07",x"02",x"02",x"08",x"00",x"00",x"00",x"00", -- 0x03B0
    x"C0",x"80",x"A0",x"10",x"00",x"00",x"00",x"00", -- 0x03B8
    x"00",x"00",x"00",x"04",x"24",x"04",x"4E",x"27", -- 0x03C0
    x"00",x"00",x"20",x"40",x"11",x"80",x"A4",x"C8", -- 0x03C8
    x"07",x"03",x"25",x"00",x"08",x"00",x"00",x"00", -- 0x03D0
    x"C0",x"20",x"90",x"A0",x"20",x"50",x"00",x"00", -- 0x03D8
    x"00",x"00",x"42",x"20",x"04",x"0F",x"E7",x"3F", -- 0x03E0
    x"00",x"20",x"44",x"C8",x"80",x"80",x"D0",x"EC", -- 0x03E8
    x"07",x"07",x"0D",x"1D",x"29",x"42",x"01",x"00", -- 0x03F0
    x"C0",x"A0",x"B0",x"88",x"44",x"20",x"10",x"08", -- 0x03F8
    x"07",x"08",x"08",x"07",x"00",x"07",x"08",x"08", -- 0x0400
    x"C0",x"20",x"20",x"C0",x"00",x"C0",x"20",x"20", -- 0x0408
    x"07",x"00",x"06",x"09",x"09",x"09",x"06",x"00", -- 0x0410
    x"C0",x"00",x"C0",x"20",x"20",x"20",x"C0",x"00", -- 0x0418
    x"00",x"07",x"08",x"08",x"07",x"00",x"07",x"08", -- 0x0420
    x"00",x"C0",x"20",x"20",x"C0",x"00",x"C0",x"20", -- 0x0428
    x"08",x"07",x"00",x"00",x"0F",x"04",x"00",x"00", -- 0x0430
    x"20",x"C0",x"00",x"20",x"E0",x"20",x"00",x"00", -- 0x0438
    x"07",x"08",x"08",x"07",x"00",x"07",x"08",x"08", -- 0x0440
    x"C0",x"20",x"20",x"C0",x"00",x"C0",x"20",x"20", -- 0x0448
    x"07",x"00",x"06",x"09",x"08",x"08",x"04",x"00", -- 0x0450
    x"C0",x"00",x"20",x"20",x"A0",x"60",x"20",x"00", -- 0x0458
    x"07",x"08",x"08",x"07",x"00",x"07",x"08",x"08", -- 0x0460
    x"C0",x"20",x"20",x"C0",x"00",x"C0",x"20",x"20", -- 0x0468
    x"07",x"00",x"08",x"0D",x"0B",x"09",x"08",x"00", -- 0x0470
    x"C0",x"00",x"C0",x"20",x"20",x"20",x"20",x"00", -- 0x0478
    x"2F",x"2B",x"7D",x"7B",x"7E",x"FF",x"BF",x"4F", -- 0x0480
    x"E3",x"E3",x"E3",x"E3",x"E3",x"73",x"FB",x"FF", -- 0x0488
    x"7F",x"FF",x"FF",x"FF",x"7F",x"9F",x"5F",x"6F", -- 0x0490
    x"FF",x"FF",x"FF",x"FF",x"7F",x"3F",x"7B",x"77", -- 0x0498
    x"27",x"37",x"37",x"3B",x"3B",x"3D",x"7D",x"7F", -- 0x04A0
    x"FE",x"FC",x"DE",x"FF",x"FF",x"8F",x"EF",x"F7", -- 0x04A8
    x"7F",x"FF",x"FF",x"BE",x"BE",x"5F",x"5F",x"4F", -- 0x04B0
    x"EF",x"7F",x"7F",x"3F",x"37",x"77",x"7F",x"FE", -- 0x04B8
    x"FF",x"DF",x"DF",x"7F",x"7F",x"17",x"1B",x"1B", -- 0x04C0
    x"5F",x"8F",x"CF",x"E7",x"F7",x"FF",x"FF",x"DF", -- 0x04C8
    x"7E",x"3E",x"7E",x"37",x"37",x"3F",x"7F",x"FF", -- 0x04D0
    x"FF",x"FF",x"FD",x"FD",x"FB",x"FF",x"BF",x"DF", -- 0x04D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04E0
    x"FF",x"FF",x"E7",x"07",x"07",x"06",x"FE",x"FE", -- 0x04E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04F0
    x"66",x"06",x"06",x"64",x"3C",x"1C",x"08",x"00", -- 0x04F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0500
    x"00",x"08",x"1C",x"3C",x"64",x"06",x"06",x"66", -- 0x0508
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0510
    x"FE",x"FE",x"E7",x"07",x"07",x"07",x"FF",x"FF", -- 0x0518
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0520
    x"FF",x"E7",x"07",x"07",x"07",x"FE",x"66",x"06", -- 0x0528
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0530
    x"06",x"64",x"3C",x"1C",x"08",x"00",x"00",x"00", -- 0x0538
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0540
    x"00",x"00",x"00",x"08",x"1C",x"3C",x"64",x"06", -- 0x0548
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0550
    x"06",x"66",x"FE",x"E7",x"07",x"07",x"07",x"FF", -- 0x0558
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0560
    x"07",x"07",x"FF",x"FF",x"FF",x"66",x"06",x"06", -- 0x0568
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0570
    x"64",x"3C",x"1C",x"08",x"00",x"00",x"00",x"00", -- 0x0578
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0580
    x"00",x"00",x"00",x"00",x"08",x"1C",x"3C",x"64", -- 0x0588
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0590
    x"06",x"06",x"66",x"FF",x"FF",x"FF",x"E7",x"07", -- 0x0598
    x"FF",x"F9",x"F1",x"61",x"61",x"63",x"37",x"3F", -- 0x05A0
    x"F9",x"F8",x"F8",x"FE",x"FF",x"FF",x"F8",x"F0", -- 0x05A8
    x"3F",x"0F",x"0E",x"00",x"00",x"00",x"00",x"00", -- 0x05B0
    x"F0",x"7B",x"3F",x"3E",x"00",x"00",x"00",x"00", -- 0x05B8
    x"00",x"00",x"00",x"00",x"01",x"0F",x"0F",x"3F", -- 0x05C0
    x"00",x"00",x"00",x"00",x"FE",x"FF",x"FF",x"FE", -- 0x05C8
    x"3F",x"37",x"63",x"61",x"61",x"F1",x"F9",x"FF", -- 0x05D0
    x"FC",x"C6",x"87",x"CF",x"FE",x"FC",x"FE",x"FF", -- 0x05D8
    x"00",x"00",x"03",x"0F",x"F2",x"CE",x"3E",x"FF", -- 0x05E0
    x"00",x"03",x"F8",x"C0",x"80",x"C0",x"30",x"08", -- 0x05E8
    x"1F",x"C6",x"F2",x"1D",x"03",x"00",x"00",x"00", -- 0x05F0
    x"CC",x"E0",x"80",x"40",x"98",x"F0",x"00",x"00", -- 0x05F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0600
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0608
    x"3F",x"3F",x"7F",x"0B",x"0B",x"07",x"03",x"02", -- 0x0610
    x"CE",x"FE",x"FE",x"EC",x"74",x"FC",x"FC",x"4C", -- 0x0618
    x"04",x"07",x"1F",x"1F",x"3D",x"7D",x"1F",x"2F", -- 0x0620
    x"04",x"04",x"F8",x"FC",x"F4",x"FC",x"FC",x"FE", -- 0x0628
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0630
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0638
    x"2E",x"1F",x"1F",x"1F",x"27",x"42",x"04",x"00", -- 0x0640
    x"7E",x"FE",x"FE",x"BE",x"BD",x"50",x"00",x"00", -- 0x0648
    x"F7",x"EB",x"DD",x"3D",x"FD",x"7F",x"F7",x"2D", -- 0x0650
    x"F7",x"EF",x"DB",x"B7",x"AF",x"BE",x"FE",x"EA", -- 0x0658
    x"7F",x"7F",x"FF",x"7E",x"BD",x"DB",x"FB",x"F7", -- 0x0660
    x"FF",x"FE",x"6F",x"AF",x"D7",x"DD",x"ED",x"F7", -- 0x0668
    x"00",x"00",x"87",x"5F",x"3B",x"7B",x"7F",x"FF", -- 0x0670
    x"00",x"02",x"FC",x"FC",x"D4",x"BE",x"4E",x"CD", -- 0x0678
    x"60",x"74",x"D8",x"CE",x"64",x"68",x"FF",x"10", -- 0x0680
    x"0B",x"37",x"7B",x"BB",x"32",x"F0",x"24",x"02", -- 0x0688
    x"FF",x"BF",x"1F",x"3F",x"2F",x"14",x"00",x"03", -- 0x0690
    x"6F",x"EF",x"F7",x"F7",x"36",x"2E",x"5E",x"85", -- 0x0698
    x"3C",x"23",x"8E",x"CF",x"4F",x"7B",x"3D",x"FE", -- 0x06A0
    x"9E",x"12",x"3B",x"7D",x"9D",x"ED",x"FB",x"F7", -- 0x06A8
    x"00",x"00",x"20",x"6C",x"F8",x"58",x"26",x"16", -- 0x06B0
    x"80",x"80",x"80",x"98",x"8C",x"16",x"1C",x"1E", -- 0x06B8
    x"1C",x"0C",x"00",x"21",x"41",x"08",x"08",x"00", -- 0x06C0
    x"40",x"20",x"60",x"C0",x"80",x"84",x"82",x"00", -- 0x06C8
    x"38",x"3C",x"18",x"00",x"01",x"03",x"08",x"1C", -- 0x06D0
    x"00",x"08",x"0C",x"0E",x"C6",x"C4",x"86",x"42", -- 0x06D8
    x"4E",x"06",x"01",x"01",x"03",x"03",x"01",x"00", -- 0x06E0
    x"20",x"00",x"06",x"0F",x"07",x"03",x"01",x"00", -- 0x06E8
    x"00",x"00",x"10",x"10",x"00",x"00",x"04",x"8E", -- 0x06F0
    x"00",x"00",x"00",x"02",x"24",x"A0",x"60",x"30", -- 0x06F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0700
    x"00",x"01",x"21",x"13",x"0F",x"0F",x"07",x"1F", -- 0x0708
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0710
    x"3F",x"5F",x"17",x"0F",x"07",x"09",x"08",x"00", -- 0x0718
    x"00",x"00",x"04",x"88",x"B0",x"F0",x"F8",x"FE", -- 0x0720
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0728
    x"C8",x"F0",x"B8",x"D8",x"E4",x"C0",x"00",x"00", -- 0x0730
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0738
    x"02",x"01",x"00",x"00",x"00",x"00",x"00",x"03", -- 0x0740
    x"00",x"07",x"8F",x"FF",x"3F",x"7C",x"7B",x"73", -- 0x0748
    x"3F",x"0E",x"00",x"00",x"01",x"02",x"00",x"00", -- 0x0750
    x"F7",x"77",x"7B",x"FD",x"1E",x"0F",x"07",x"05", -- 0x0758
    x"00",x"30",x"F8",x"FF",x"FF",x"EF",x"EF",x"F7", -- 0x0760
    x"00",x"00",x"40",x"80",x"00",x"80",x"C0",x"C0", -- 0x0768
    x"F3",x"F7",x"EF",x"FF",x"9C",x"F8",x"E4",x"80", -- 0x0770
    x"B8",x"84",x"00",x"00",x"C0",x"20",x"00",x"00", -- 0x0778
    x"10",x"08",x"00",x"00",x"11",x"1F",x"0F",x"1F", -- 0x0780
    x"0E",x"1E",x"3E",x"BF",x"DF",x"EE",x"FF",x"FF", -- 0x0788
    x"1F",x"07",x"03",x"31",x"00",x"01",x"03",x"00", -- 0x0790
    x"FF",x"CF",x"BF",x"7F",x"FE",x"BF",x"1F",x"07", -- 0x0798
    x"00",x"F8",x"FF",x"FF",x"FF",x"FF",x"F8",x"E7", -- 0x07A0
    x"00",x"10",x"30",x"F0",x"F8",x"FC",x"0C",x"FC", -- 0x07A8
    x"EF",x"FF",x"FF",x"FF",x"EF",x"1C",x"F8",x"80", -- 0x07B0
    x"FC",x"FC",x"F8",x"F0",x"80",x"46",x"22",x"00", -- 0x07B8
    x"00",x"00",x"39",x"31",x"69",x"00",x"00",x"00", -- 0x07C0
    x"00",x"00",x"8F",x"DF",x"C6",x"07",x"01",x"00", -- 0x07C8
    x"0C",x"38",x"00",x"0C",x"1E",x"0C",x"00",x"00", -- 0x07D0
    x"01",x"39",x"38",x"18",x"00",x"00",x"00",x"00", -- 0x07D8
    x"00",x"18",x"1A",x"1A",x"03",x"02",x"44",x"C0", -- 0x07E0
    x"00",x"00",x"00",x"00",x"70",x"60",x"00",x"00", -- 0x07E8
    x"C1",x"01",x"00",x"70",x"70",x"60",x"00",x"00", -- 0x07F0
    x"80",x"80",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07F8
    x"38",x"7C",x"C2",x"82",x"86",x"7C",x"38",x"00", -- 0x0800
    x"02",x"02",x"FE",x"FE",x"42",x"02",x"00",x"00", -- 0x0808
    x"62",x"F2",x"BA",x"9A",x"9E",x"CE",x"46",x"00", -- 0x0810
    x"8C",x"DE",x"F2",x"B2",x"92",x"86",x"04",x"00", -- 0x0818
    x"08",x"FE",x"FE",x"C8",x"68",x"38",x"18",x"00", -- 0x0820
    x"1C",x"BE",x"A2",x"A2",x"A2",x"E6",x"E4",x"00", -- 0x0828
    x"0C",x"9E",x"92",x"92",x"D2",x"7E",x"3C",x"00", -- 0x0830
    x"C0",x"E0",x"B0",x"9E",x"8E",x"C0",x"C0",x"00", -- 0x0838
    x"0C",x"6E",x"9A",x"9A",x"B2",x"F2",x"6C",x"00", -- 0x0840
    x"78",x"FC",x"96",x"92",x"92",x"F2",x"60",x"00", -- 0x0848
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0850
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0858
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0860
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0868
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0870
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0878
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0880
    x"3E",x"7E",x"C8",x"88",x"C8",x"7E",x"3E",x"00", -- 0x0888
    x"6C",x"FE",x"92",x"92",x"92",x"FE",x"FE",x"00", -- 0x0890
    x"44",x"C6",x"82",x"82",x"C6",x"7C",x"38",x"00", -- 0x0898
    x"38",x"7C",x"C6",x"82",x"82",x"FE",x"FE",x"00", -- 0x08A0
    x"82",x"92",x"92",x"92",x"FE",x"FE",x"00",x"00", -- 0x08A8
    x"80",x"90",x"90",x"90",x"90",x"FE",x"FE",x"00", -- 0x08B0
    x"9E",x"9E",x"92",x"82",x"C6",x"7C",x"38",x"00", -- 0x08B8
    x"FE",x"FE",x"10",x"10",x"10",x"FE",x"FE",x"00", -- 0x08C0
    x"82",x"82",x"FE",x"FE",x"82",x"82",x"00",x"00", -- 0x08C8
    x"FC",x"FE",x"02",x"02",x"02",x"06",x"04",x"00", -- 0x08D0
    x"82",x"C6",x"6E",x"3C",x"18",x"FE",x"FE",x"00", -- 0x08D8
    x"02",x"02",x"02",x"02",x"FE",x"FE",x"00",x"00", -- 0x08E0
    x"FE",x"FE",x"70",x"38",x"70",x"FE",x"FE",x"00", -- 0x08E8
    x"FE",x"FE",x"1C",x"38",x"70",x"FE",x"FE",x"00", -- 0x08F0
    x"7C",x"FE",x"82",x"82",x"82",x"FE",x"7C",x"00", -- 0x08F8
    x"70",x"F8",x"88",x"88",x"88",x"FE",x"FE",x"00", -- 0x0900
    x"7A",x"FC",x"8E",x"8A",x"82",x"FE",x"7C",x"00", -- 0x0908
    x"72",x"F6",x"9E",x"8C",x"88",x"FE",x"FE",x"00", -- 0x0910
    x"0C",x"5E",x"D2",x"92",x"92",x"F6",x"64",x"00", -- 0x0918
    x"80",x"80",x"FE",x"FE",x"80",x"80",x"00",x"00", -- 0x0920
    x"FC",x"FE",x"02",x"02",x"02",x"FE",x"FC",x"00", -- 0x0928
    x"F0",x"F8",x"1C",x"0E",x"1C",x"F8",x"F0",x"00", -- 0x0930
    x"F8",x"FE",x"1C",x"38",x"1C",x"FE",x"F8",x"00", -- 0x0938
    x"C6",x"EE",x"7C",x"38",x"7C",x"EE",x"C6",x"00", -- 0x0940
    x"C0",x"F0",x"1E",x"1E",x"F0",x"C0",x"00",x"00", -- 0x0948
    x"C2",x"E2",x"F2",x"BA",x"9E",x"8E",x"86",x"00", -- 0x0950
    x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00", -- 0x0958
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0960
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0968
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0970
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0978
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0980
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0988
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0990
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0998
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x09A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x09A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x09B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x09B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x09C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x09C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x09D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x09D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x09E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x09E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x09F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x09F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A18
    x"00",x"00",x"00",x"01",x"01",x"01",x"1D",x"0F", -- 0x0A20
    x"00",x"40",x"C0",x"C0",x"C0",x"C0",x"C0",x"40", -- 0x0A28
    x"0F",x"1F",x"01",x"01",x"01",x"00",x"00",x"00", -- 0x0A30
    x"40",x"C0",x"C0",x"C0",x"C0",x"C0",x"40",x"00", -- 0x0A38
    x"1D",x"74",x"1F",x"33",x"23",x"03",x"01",x"01", -- 0x0A40
    x"80",x"C0",x"80",x"E0",x"80",x"80",x"C0",x"C0", -- 0x0A48
    x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A50
    x"C0",x"C0",x"C0",x"00",x"00",x"00",x"00",x"00", -- 0x0A58
    x"FB",x"4B",x"FD",x"47",x"47",x"67",x"03",x"03", -- 0x0A60
    x"80",x"00",x"80",x"C0",x"00",x"00",x"00",x"00", -- 0x0A68
    x"03",x"03",x"03",x"01",x"01",x"00",x"00",x"00", -- 0x0A70
    x"00",x"00",x"80",x"C0",x"C0",x"C0",x"C0",x"C0", -- 0x0A78
    x"10",x"AC",x"D6",x"98",x"6F",x"23",x"7B",x"03", -- 0x0A80
    x"C0",x"C0",x"C0",x"C0",x"C0",x"80",x"00",x"00", -- 0x0A88
    x"03",x"03",x"67",x"47",x"47",x"7D",x"CB",x"7B", -- 0x0A90
    x"00",x"00",x"00",x"00",x"C0",x"80",x"D0",x"80", -- 0x0A98
    x"EB",x"BD",x"8F",x"CF",x"1E",x"0E",x"0C",x"0C", -- 0x0AA0
    x"10",x"C0",x"20",x"80",x"40",x"00",x"00",x"00", -- 0x0AA8
    x"1C",x"1C",x"1C",x"1E",x"0E",x"0C",x"0C",x"04", -- 0x0AB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0AB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0AC0
    x"00",x"0C",x"0C",x"1C",x"38",x"78",x"70",x"D0", -- 0x0AC8
    x"00",x"39",x"A3",x"B3",x"5F",x"5C",x"FD",x"5B", -- 0x0AD0
    x"C0",x"C0",x"C0",x"80",x"E0",x"D0",x"E0",x"90", -- 0x0AD8
    x"00",x"00",x"00",x"00",x"01",x"01",x"13",x"1F", -- 0x0AE0
    x"00",x"00",x"00",x"00",x"40",x"40",x"E4",x"FC", -- 0x0AE8
    x"03",x"01",x"01",x"00",x"00",x"00",x"00",x"00", -- 0x0AF0
    x"E0",x"C0",x"C0",x"80",x"00",x"00",x"00",x"00", -- 0x0AF8
    x"00",x"00",x"00",x"01",x"03",x"1C",x"23",x"C0", -- 0x0B00
    x"00",x"7E",x"FC",x"08",x"F1",x"13",x"FF",x"0F", -- 0x0B08
    x"23",x"1C",x"03",x"01",x"00",x"00",x"00",x"00", -- 0x0B10
    x"FF",x"13",x"F1",x"08",x"FC",x"7E",x"00",x"00", -- 0x0B18
    x"1C",x"38",x"C2",x"06",x"C2",x"38",x"1C",x"00", -- 0x0B20
    x"00",x"00",x"00",x"18",x"08",x"1C",x"FE",x"F8", -- 0x0B28
    x"0C",x"06",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B30
    x"FE",x"1C",x"08",x"18",x"00",x"00",x"00",x"00", -- 0x0B38
    x"02",x"07",x"07",x"0F",x"0F",x"0F",x"1F",x"18", -- 0x0B40
    x"00",x"00",x"00",x"80",x"80",x"80",x"C0",x"C0", -- 0x0B48
    x"17",x"37",x"38",x"3F",x"70",x"7F",x"7F",x"00", -- 0x0B50
    x"40",x"60",x"E0",x"E0",x"70",x"F0",x"F0",x"00", -- 0x0B58
    x"02",x"02",x"07",x"07",x"0F",x"0F",x"1F",x"00", -- 0x0B60
    x"00",x"00",x"00",x"00",x"80",x"80",x"C0",x"00", -- 0x0B68
    x"7F",x"00",x"00",x"0F",x"7F",x"48",x"7F",x"00", -- 0x0B70
    x"00",x"03",x"03",x"00",x"00",x"7F",x"41",x"41", -- 0x0B78
    x"00",x"01",x"03",x"07",x"03",x"07",x"0F",x"3F", -- 0x0B80
    x"80",x"80",x"D8",x"F8",x"F8",x"F0",x"F0",x"F0", -- 0x0B88
    x"1F",x"1F",x"1F",x"0F",x"03",x"07",x"07",x"01", -- 0x0B90
    x"F8",x"F8",x"F0",x"E0",x"F8",x"FC",x"78",x"00", -- 0x0B98
    x"00",x"00",x"00",x"00",x"00",x"04",x"01",x"03", -- 0x0BA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"90", -- 0x0BA8
    x"07",x"02",x"02",x"08",x"00",x"00",x"00",x"00", -- 0x0BB0
    x"C0",x"80",x"A0",x"10",x"00",x"00",x"00",x"00", -- 0x0BB8
    x"00",x"00",x"00",x"04",x"24",x"04",x"4E",x"27", -- 0x0BC0
    x"00",x"00",x"20",x"40",x"11",x"80",x"A4",x"C8", -- 0x0BC8
    x"07",x"03",x"25",x"00",x"08",x"00",x"00",x"00", -- 0x0BD0
    x"C0",x"20",x"90",x"A0",x"20",x"50",x"00",x"00", -- 0x0BD8
    x"00",x"00",x"42",x"20",x"04",x"0F",x"E7",x"3F", -- 0x0BE0
    x"00",x"20",x"44",x"C8",x"80",x"80",x"D0",x"EC", -- 0x0BE8
    x"07",x"07",x"0D",x"1D",x"29",x"42",x"01",x"00", -- 0x0BF0
    x"C0",x"A0",x"B0",x"88",x"44",x"20",x"10",x"08", -- 0x0BF8
    x"07",x"08",x"08",x"07",x"00",x"07",x"08",x"08", -- 0x0C00
    x"C0",x"20",x"20",x"C0",x"00",x"C0",x"20",x"20", -- 0x0C08
    x"07",x"00",x"06",x"09",x"09",x"09",x"06",x"00", -- 0x0C10
    x"C0",x"00",x"C0",x"20",x"20",x"20",x"C0",x"00", -- 0x0C18
    x"00",x"07",x"08",x"08",x"07",x"00",x"07",x"08", -- 0x0C20
    x"00",x"C0",x"20",x"20",x"C0",x"00",x"C0",x"20", -- 0x0C28
    x"08",x"07",x"00",x"00",x"0F",x"04",x"00",x"00", -- 0x0C30
    x"20",x"C0",x"00",x"20",x"E0",x"20",x"00",x"00", -- 0x0C38
    x"07",x"08",x"08",x"07",x"00",x"07",x"08",x"08", -- 0x0C40
    x"C0",x"20",x"20",x"C0",x"00",x"C0",x"20",x"20", -- 0x0C48
    x"07",x"00",x"06",x"09",x"08",x"08",x"04",x"00", -- 0x0C50
    x"C0",x"00",x"20",x"20",x"A0",x"60",x"20",x"00", -- 0x0C58
    x"07",x"08",x"08",x"07",x"00",x"07",x"08",x"08", -- 0x0C60
    x"C0",x"20",x"20",x"C0",x"00",x"C0",x"20",x"20", -- 0x0C68
    x"07",x"00",x"08",x"0D",x"0B",x"09",x"08",x"00", -- 0x0C70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"23", -- 0x0DA0
    x"00",x"00",x"20",x"10",x"18",x"38",x"FC",x"78", -- 0x0DA8
    x"33",x"1F",x"1F",x"0F",x"01",x"00",x"00",x"00", -- 0x0DB0
    x"78",x"D8",x"48",x"20",x"B0",x"10",x"00",x"00", -- 0x0DB8
    x"00",x"00",x"00",x"00",x"00",x"20",x"31",x"1F", -- 0x0DC0
    x"00",x"00",x"00",x"08",x"08",x"1C",x"7C",x"7C", -- 0x0DC8
    x"1F",x"1F",x"06",x"02",x"00",x"00",x"00",x"00", -- 0x0DD0
    x"F8",x"B8",x"90",x"C0",x"40",x"40",x"00",x"00", -- 0x0DD8
    x"00",x"00",x"00",x"00",x"10",x"10",x"19",x"1F", -- 0x0DE0
    x"00",x"00",x"00",x"00",x"04",x"04",x"4C",x"7C", -- 0x0DE8
    x"1F",x"0E",x"06",x"02",x"00",x"00",x"00",x"00", -- 0x0DF0
    x"FC",x"B8",x"B0",x"A0",x"80",x"80",x"00",x"00", -- 0x0DF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E08
    x"3F",x"3F",x"7F",x"0B",x"0B",x"07",x"03",x"02", -- 0x0E10
    x"CE",x"FE",x"FE",x"EC",x"74",x"FC",x"FC",x"4C", -- 0x0E18
    x"04",x"07",x"1F",x"1F",x"3D",x"7D",x"1F",x"2F", -- 0x0E20
    x"04",x"04",x"F8",x"FC",x"F4",x"FC",x"FC",x"FE", -- 0x0E28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E38
    x"2E",x"1F",x"1F",x"1F",x"27",x"42",x"04",x"00", -- 0x0E40
    x"7E",x"FE",x"FE",x"BE",x"BD",x"50",x"00",x"00", -- 0x0E48
    x"F7",x"EB",x"DD",x"3D",x"FD",x"7F",x"F7",x"2D", -- 0x0E50
    x"F7",x"EF",x"DB",x"B7",x"AF",x"BE",x"FE",x"EA", -- 0x0E58
    x"7F",x"7F",x"FF",x"7E",x"BD",x"DB",x"FB",x"F7", -- 0x0E60
    x"FF",x"FE",x"6F",x"AF",x"D7",x"DD",x"ED",x"F7", -- 0x0E68
    x"00",x"00",x"87",x"5F",x"3B",x"7B",x"7F",x"FF", -- 0x0E70
    x"00",x"02",x"FC",x"FC",x"D4",x"BE",x"4E",x"CD", -- 0x0E78
    x"60",x"74",x"D8",x"CE",x"64",x"68",x"FF",x"10", -- 0x0E80
    x"0B",x"37",x"7B",x"BB",x"32",x"F0",x"24",x"02", -- 0x0E88
    x"FF",x"BF",x"1F",x"3F",x"2F",x"14",x"00",x"03", -- 0x0E90
    x"6F",x"EF",x"F7",x"F7",x"36",x"2E",x"5E",x"85", -- 0x0E98
    x"3C",x"23",x"8E",x"CF",x"4F",x"7B",x"3D",x"FE", -- 0x0EA0
    x"9E",x"12",x"3B",x"7D",x"9D",x"ED",x"FB",x"F7", -- 0x0EA8
    x"00",x"00",x"20",x"6C",x"F8",x"58",x"26",x"16", -- 0x0EB0
    x"80",x"80",x"80",x"98",x"8C",x"16",x"1C",x"1E", -- 0x0EB8
    x"1C",x"0C",x"00",x"21",x"41",x"08",x"08",x"00", -- 0x0EC0
    x"40",x"20",x"60",x"C0",x"80",x"84",x"82",x"00", -- 0x0EC8
    x"38",x"3C",x"18",x"00",x"01",x"03",x"08",x"1C", -- 0x0ED0
    x"00",x"08",x"0C",x"0E",x"C6",x"C4",x"86",x"42", -- 0x0ED8
    x"4E",x"06",x"01",x"01",x"03",x"03",x"01",x"00", -- 0x0EE0
    x"20",x"00",x"06",x"0F",x"07",x"03",x"01",x"00", -- 0x0EE8
    x"00",x"00",x"10",x"10",x"00",x"00",x"04",x"8E", -- 0x0EF0
    x"00",x"00",x"00",x"02",x"24",x"A0",x"60",x"30", -- 0x0EF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F00
    x"00",x"01",x"21",x"13",x"0F",x"0F",x"07",x"1F", -- 0x0F08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F10
    x"3F",x"5F",x"17",x"0F",x"07",x"09",x"08",x"00", -- 0x0F18
    x"00",x"00",x"04",x"88",x"B0",x"F0",x"F8",x"FE", -- 0x0F20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F28
    x"C8",x"F0",x"B8",x"D8",x"E4",x"C0",x"00",x"00", -- 0x0F30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F38
    x"02",x"01",x"00",x"00",x"00",x"00",x"00",x"03", -- 0x0F40
    x"00",x"07",x"8F",x"FF",x"3F",x"7C",x"7B",x"73", -- 0x0F48
    x"3F",x"0E",x"00",x"00",x"01",x"02",x"00",x"00", -- 0x0F50
    x"F7",x"77",x"7B",x"FD",x"1E",x"0F",x"07",x"05", -- 0x0F58
    x"00",x"30",x"F8",x"FF",x"FF",x"EF",x"EF",x"F7", -- 0x0F60
    x"00",x"00",x"40",x"80",x"00",x"80",x"C0",x"C0", -- 0x0F68
    x"F3",x"F7",x"EF",x"FF",x"9C",x"F8",x"E4",x"80", -- 0x0F70
    x"B8",x"84",x"00",x"00",x"C0",x"20",x"00",x"00", -- 0x0F78
    x"10",x"08",x"00",x"00",x"11",x"1F",x"0F",x"1F", -- 0x0F80
    x"0E",x"1E",x"3E",x"BF",x"DF",x"EE",x"FF",x"FF", -- 0x0F88
    x"1F",x"07",x"03",x"31",x"00",x"01",x"03",x"00", -- 0x0F90
    x"FF",x"CF",x"BF",x"7F",x"FE",x"BF",x"1F",x"07", -- 0x0F98
    x"00",x"F8",x"FF",x"FF",x"FF",x"FF",x"F8",x"E7", -- 0x0FA0
    x"00",x"10",x"30",x"F0",x"F8",x"FC",x"0C",x"FC", -- 0x0FA8
    x"EF",x"FF",x"FF",x"FF",x"EF",x"1C",x"F8",x"80", -- 0x0FB0
    x"FC",x"FC",x"F8",x"F0",x"80",x"46",x"22",x"00", -- 0x0FB8
    x"00",x"00",x"39",x"31",x"69",x"00",x"00",x"00", -- 0x0FC0
    x"00",x"00",x"8F",x"DF",x"C6",x"07",x"01",x"00", -- 0x0FC8
    x"0C",x"38",x"00",x"0C",x"1E",x"0C",x"00",x"00", -- 0x0FD0
    x"01",x"39",x"38",x"18",x"00",x"00",x"00",x"00", -- 0x0FD8
    x"00",x"18",x"1A",x"1A",x"03",x"02",x"44",x"C0", -- 0x0FE0
    x"00",x"00",x"00",x"00",x"70",x"60",x"00",x"00", -- 0x0FE8
    x"C1",x"01",x"00",x"70",x"70",x"60",x"00",x"00", -- 0x0FF0
    x"80",x"80",x"00",x"00",x"00",x"00",x"00",x"00"  -- 0x0FF8
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
       DATA <= ROM(to_integer(unsigned(ADDR)));
  end process;
end RTL;
