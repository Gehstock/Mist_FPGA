library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_H5 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_H5 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"6C",X"C6",X"C6",X"FE",X"C6",X"C6",
		X"00",X"FC",X"C6",X"C6",X"FC",X"C6",X"C6",X"FC",X"00",X"3C",X"66",X"C0",X"C0",X"C0",X"66",X"3C",
		X"00",X"F8",X"CC",X"C6",X"C6",X"C6",X"CC",X"F8",X"00",X"FC",X"C0",X"C0",X"F8",X"C0",X"C0",X"FE",
		X"00",X"FE",X"C0",X"C0",X"FC",X"C0",X"C0",X"C0",X"00",X"3E",X"60",X"C0",X"CE",X"C6",X"66",X"3E",
		X"00",X"C6",X"C6",X"C6",X"FE",X"C6",X"C6",X"C6",X"00",X"FC",X"30",X"30",X"30",X"30",X"30",X"FC",
		X"00",X"06",X"06",X"06",X"06",X"06",X"C6",X"7C",X"00",X"C6",X"CC",X"D8",X"F0",X"F8",X"DC",X"CE",
		X"00",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"FE",X"00",X"C6",X"EE",X"FE",X"FE",X"D6",X"C6",X"C6",
		X"00",X"C6",X"E6",X"F6",X"FE",X"DE",X"CE",X"C6",X"00",X"7C",X"C6",X"C6",X"C6",X"C6",X"C6",X"7C",
		X"00",X"FC",X"C6",X"C6",X"C6",X"FC",X"C0",X"C0",X"00",X"7C",X"C6",X"C6",X"C6",X"CE",X"CC",X"7A",
		X"00",X"FC",X"C6",X"C6",X"CE",X"F8",X"DC",X"CE",X"00",X"78",X"CC",X"C0",X"7C",X"06",X"C6",X"7C",
		X"00",X"FC",X"30",X"30",X"30",X"30",X"30",X"30",X"00",X"C6",X"C6",X"C6",X"C6",X"C6",X"C6",X"7C",
		X"00",X"C6",X"C6",X"C6",X"EE",X"7C",X"38",X"10",X"00",X"C6",X"C6",X"D6",X"FE",X"FE",X"EE",X"C6",
		X"00",X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",X"CC",X"CC",X"CC",X"78",X"30",X"30",X"30",
		X"00",X"FE",X"0E",X"1C",X"38",X"70",X"E0",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"EE",X"4A",X"4E",X"4C",X"4A",X"00",X"00",X"00",X"4D",X"E9",X"AD",X"E9",X"A9",X"00",X"00",
		X"00",X"D7",X"14",X"94",X"14",X"17",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"00",
		X"00",X"10",X"38",X"54",X"10",X"10",X"00",X"00",X"00",X"00",X"1C",X"0C",X"14",X"20",X"00",X"00",
		X"08",X"1C",X"36",X"77",X"77",X"77",X"36",X"1C",X"08",X"1C",X"22",X"7B",X"63",X"6F",X"22",X"1C",
		X"08",X"1C",X"22",X"7B",X"63",X"7B",X"22",X"1C",X"08",X"1C",X"2A",X"6B",X"63",X"7B",X"3A",X"1C",
		X"08",X"1C",X"22",X"6F",X"63",X"7B",X"22",X"1C",X"08",X"1C",X"2E",X"6F",X"63",X"6B",X"22",X"1C",
		X"08",X"1C",X"22",X"7B",X"7B",X"7B",X"3A",X"1C",X"08",X"1C",X"22",X"6B",X"63",X"6B",X"22",X"1C",
		X"08",X"1C",X"22",X"6B",X"63",X"7B",X"3A",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"38",X"4C",X"C6",X"C6",X"C6",X"64",X"38",X"00",X"30",X"70",X"30",X"30",X"30",X"30",X"FC",
		X"00",X"7C",X"C6",X"0E",X"3C",X"78",X"E0",X"FE",X"00",X"7E",X"0C",X"18",X"3C",X"06",X"C6",X"7C",
		X"00",X"1C",X"3C",X"6C",X"CC",X"FE",X"0C",X"0C",X"00",X"FC",X"C0",X"FC",X"06",X"06",X"C6",X"7C",
		X"00",X"3C",X"60",X"C0",X"FC",X"C6",X"C6",X"7C",X"00",X"FE",X"C6",X"0C",X"18",X"30",X"30",X"30",
		X"00",X"78",X"C4",X"E4",X"78",X"9E",X"86",X"7C",X"00",X"7C",X"C6",X"C6",X"7E",X"06",X"0C",X"78",
		X"00",X"10",X"38",X"AA",X"AA",X"28",X"AA",X"BA",X"00",X"10",X"38",X"BA",X"BA",X"38",X"BA",X"BA",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"FC",X"26",X"22",X"26",X"FC",X"F8",X"00",
		X"FE",X"FE",X"92",X"92",X"92",X"FE",X"6C",X"00",X"38",X"7C",X"C6",X"82",X"82",X"C6",X"44",X"00",
		X"FE",X"FE",X"82",X"82",X"C6",X"7C",X"38",X"00",X"FE",X"FE",X"92",X"92",X"92",X"82",X"80",X"00",
		X"FE",X"FE",X"12",X"12",X"12",X"12",X"02",X"00",X"38",X"7C",X"C6",X"82",X"92",X"F2",X"F2",X"00",
		X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",X"82",X"82",X"FE",X"FE",X"82",X"82",X"00",X"00",
		X"40",X"C0",X"80",X"80",X"80",X"FE",X"7E",X"00",X"FE",X"FE",X"30",X"78",X"EC",X"C6",X"82",X"00",
		X"FE",X"FE",X"80",X"80",X"80",X"80",X"80",X"00",X"FE",X"FE",X"1C",X"38",X"1C",X"FE",X"FE",X"00",
		X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",X"00",
		X"FE",X"FE",X"22",X"22",X"22",X"3E",X"1C",X"00",X"7C",X"FE",X"82",X"A2",X"E2",X"7E",X"BC",X"00",
		X"FE",X"FE",X"22",X"62",X"F2",X"DE",X"9C",X"00",X"4C",X"DE",X"92",X"92",X"96",X"F4",X"60",X"00",
		X"02",X"02",X"FE",X"FE",X"02",X"02",X"00",X"00",X"7E",X"FE",X"80",X"80",X"80",X"FE",X"7E",X"00",
		X"1E",X"3E",X"70",X"E0",X"70",X"3E",X"1E",X"00",X"FE",X"FE",X"70",X"38",X"70",X"FE",X"FE",X"00",
		X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",X"0E",X"1E",X"F0",X"F0",X"1E",X"0E",X"00",X"00",
		X"C2",X"E2",X"F2",X"B2",X"9E",X"8E",X"86",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"3E",X"02",X"00",X"3E",X"1A",X"2E",X"00",X"3C",X"16",X"3C",X"00",X"3E",X"0A",X"00",X"3E",
		X"0A",X"02",X"00",X"3E",X"00",X"3E",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"60",X"60",X"00",X"00",X"60",X"60",X"00",X"00",X"60",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"04",X"3E",X"04",X"08",X"00",X"00",X"00",X"00",X"20",X"14",X"0C",X"1C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",X"00",X"80",X"84",X"FE",X"FE",X"80",X"80",X"00",X"00",
		X"C4",X"E6",X"F2",X"B2",X"BA",X"9E",X"8C",X"00",X"40",X"C2",X"92",X"9A",X"9E",X"F6",X"62",X"00",
		X"30",X"38",X"2C",X"26",X"FE",X"FE",X"20",X"00",X"4E",X"CE",X"8A",X"8A",X"8A",X"FA",X"70",X"00",
		X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",X"00",X"06",X"06",X"E2",X"F2",X"1A",X"0E",X"06",X"00",
		X"6C",X"9E",X"9A",X"B2",X"B2",X"EC",X"60",X"00",X"0C",X"9E",X"92",X"92",X"D2",X"7E",X"3C",X"00",
		X"D8",X"00",X"FC",X"86",X"FC",X"00",X"D8",X"00",X"D8",X"00",X"FC",X"FE",X"FC",X"00",X"D8",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"63",X"63",X"7F",X"63",X"63",X"36",X"1C",X"0C",
		X"3F",X"63",X"63",X"3F",X"63",X"63",X"3F",X"00",X"3C",X"66",X"03",X"03",X"03",X"66",X"3C",X"00",
		X"1F",X"33",X"63",X"63",X"63",X"33",X"1F",X"00",X"7F",X"03",X"03",X"1F",X"03",X"03",X"3F",X"00",
		X"03",X"03",X"03",X"3F",X"03",X"03",X"7F",X"00",X"7C",X"66",X"63",X"73",X"03",X"06",X"7C",X"00",
		X"63",X"63",X"63",X"7F",X"63",X"63",X"63",X"00",X"3F",X"0C",X"0C",X"0C",X"0C",X"0C",X"3F",X"00",
		X"3E",X"63",X"60",X"60",X"60",X"60",X"60",X"00",X"73",X"3B",X"1F",X"0F",X"1B",X"33",X"63",X"00",
		X"7F",X"03",X"03",X"03",X"03",X"03",X"03",X"00",X"63",X"63",X"6B",X"7F",X"7F",X"77",X"63",X"00",
		X"63",X"73",X"7B",X"7F",X"6F",X"67",X"63",X"00",X"3E",X"63",X"63",X"63",X"63",X"63",X"3E",X"00",
		X"03",X"03",X"3F",X"63",X"63",X"63",X"3F",X"00",X"5E",X"33",X"7B",X"63",X"63",X"63",X"3E",X"00",
		X"73",X"3B",X"1F",X"73",X"63",X"63",X"3F",X"00",X"3E",X"63",X"60",X"3E",X"03",X"33",X"1E",X"00",
		X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"3F",X"00",X"3E",X"63",X"63",X"63",X"63",X"63",X"63",X"00",
		X"08",X"1C",X"3E",X"77",X"63",X"63",X"63",X"00",X"63",X"77",X"7F",X"7F",X"6B",X"63",X"63",X"00",
		X"63",X"77",X"3E",X"1C",X"3E",X"77",X"63",X"00",X"0C",X"0C",X"0C",X"1E",X"33",X"33",X"33",X"00",
		X"7F",X"07",X"0E",X"1C",X"38",X"70",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"52",X"32",X"72",X"52",X"77",X"00",X"00",X"00",X"95",X"97",X"B5",X"97",X"B2",X"00",
		X"00",X"00",X"E8",X"28",X"29",X"28",X"EB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"08",X"2A",X"1C",X"08",X"00",X"00",X"00",X"04",X"28",X"30",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1C",X"26",X"63",X"63",X"63",X"32",X"1C",X"00",X"3F",X"0C",X"0C",X"0C",X"0C",X"0E",X"0C",X"00",
		X"7F",X"07",X"1E",X"3C",X"70",X"63",X"3E",X"00",X"3E",X"63",X"60",X"3C",X"18",X"30",X"7E",X"00",
		X"30",X"30",X"7F",X"33",X"36",X"3C",X"38",X"00",X"3E",X"63",X"60",X"60",X"3F",X"03",X"3F",X"00",
		X"3E",X"63",X"63",X"3F",X"03",X"06",X"3C",X"00",X"0C",X"0C",X"0C",X"18",X"30",X"63",X"6F",X"00",
		X"3E",X"61",X"79",X"1E",X"27",X"23",X"1E",X"00",X"1E",X"30",X"60",X"7E",X"63",X"63",X"3E",X"00",
		X"5D",X"55",X"14",X"55",X"55",X"1C",X"08",X"00",X"5D",X"5D",X"1C",X"5D",X"5D",X"1C",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"3F",X"64",X"44",X"64",X"3F",X"1F",
		X"00",X"36",X"7F",X"49",X"49",X"49",X"7F",X"7F",X"00",X"22",X"63",X"41",X"41",X"63",X"3E",X"1C",
		X"00",X"1C",X"3E",X"63",X"41",X"41",X"7F",X"7F",X"00",X"01",X"41",X"49",X"49",X"49",X"7F",X"7F",
		X"00",X"40",X"48",X"48",X"48",X"48",X"7F",X"7F",X"00",X"4F",X"4F",X"49",X"41",X"63",X"3E",X"1C",
		X"00",X"7F",X"7F",X"08",X"08",X"08",X"7F",X"7F",X"00",X"00",X"41",X"41",X"7F",X"7F",X"41",X"41",
		X"00",X"7E",X"7F",X"01",X"01",X"01",X"03",X"02",X"00",X"41",X"63",X"37",X"1E",X"0C",X"7F",X"7F",
		X"00",X"01",X"01",X"01",X"01",X"01",X"7F",X"7F",X"00",X"7F",X"7F",X"38",X"1C",X"38",X"7F",X"7F",
		X"00",X"7F",X"7F",X"0E",X"1C",X"38",X"7F",X"7F",X"00",X"3E",X"7F",X"41",X"41",X"41",X"7F",X"3E",
		X"00",X"38",X"7C",X"44",X"44",X"44",X"7F",X"7F",X"00",X"3D",X"7E",X"47",X"45",X"41",X"7F",X"3E",
		X"00",X"39",X"7B",X"4F",X"46",X"44",X"7F",X"7F",X"00",X"06",X"2F",X"69",X"49",X"49",X"7B",X"32",
		X"00",X"00",X"40",X"40",X"7F",X"7F",X"40",X"40",X"00",X"7E",X"7F",X"01",X"01",X"01",X"7F",X"7E",
		X"00",X"78",X"7C",X"0E",X"07",X"0E",X"7C",X"78",X"00",X"7F",X"7F",X"0E",X"1C",X"0E",X"7F",X"7F",
		X"00",X"63",X"77",X"3E",X"1C",X"3E",X"77",X"63",X"00",X"00",X"70",X"78",X"0F",X"0F",X"78",X"70",
		X"00",X"61",X"71",X"79",X"5D",X"4F",X"47",X"43",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"74",X"58",X"7C",X"00",X"40",X"7C",X"40",X"7C",X"00",X"50",X"7C",X"00",X"3C",X"68",X"3C",
		X"44",X"44",X"7C",X"00",X"7C",X"00",X"40",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"06",X"06",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"00",
		X"00",X"00",X"10",X"20",X"7C",X"20",X"10",X"00",X"00",X"00",X"38",X"30",X"28",X"04",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"1C",X"3E",X"61",X"41",X"43",X"3E",X"1C",X"00",X"00",X"01",X"01",X"7F",X"7F",X"21",X"01",
		X"00",X"31",X"79",X"5D",X"4D",X"4F",X"67",X"23",X"00",X"46",X"6F",X"79",X"59",X"49",X"43",X"02",
		X"00",X"04",X"7F",X"7F",X"64",X"34",X"1C",X"0C",X"00",X"0E",X"5F",X"51",X"51",X"51",X"73",X"72",
		X"00",X"06",X"4F",X"49",X"49",X"69",X"3F",X"1E",X"00",X"60",X"70",X"58",X"4F",X"47",X"60",X"60",
		X"00",X"06",X"37",X"4D",X"4D",X"59",X"79",X"36",X"00",X"3C",X"7E",X"4B",X"49",X"49",X"79",X"30",
		X"00",X"1B",X"00",X"3F",X"61",X"3F",X"00",X"1B",X"00",X"1B",X"00",X"3F",X"7F",X"3F",X"00",X"1B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
