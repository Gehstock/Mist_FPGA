library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_PGM_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_PGM_1 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"30",X"10",X"21",X"FF",X"00",X"22",X"0A",X"4D",X"3A",X"0C",X"4D",X"3D",X"32",X"0C",X"4D",X"CA",
		X"F1",X"30",X"CD",X"2D",X"32",X"FE",X"0F",X"28",X"1F",X"21",X"0D",X"4D",X"CB",X"46",X"20",X"1D",
		X"2A",X"04",X"4D",X"36",X"40",X"FE",X"00",X"28",X"35",X"FE",X"01",X"28",X"46",X"FE",X"02",X"28",
		X"50",X"FE",X"03",X"28",X"59",X"C3",X"9C",X"30",X"21",X"0D",X"4D",X"CB",X"86",X"3A",X"2C",X"4C",
		X"CB",X"67",X"28",X"0D",X"2A",X"04",X"4D",X"36",X"81",X"2A",X"06",X"4D",X"36",X"80",X"C3",X"F0",
		X"27",X"2A",X"04",X"4D",X"36",X"40",X"2A",X"06",X"4D",X"36",X"40",X"C3",X"F0",X"27",X"7D",X"E6",
		X"1F",X"FE",X"06",X"28",X"07",X"7D",X"D6",X"03",X"6F",X"22",X"04",X"4D",X"21",X"0D",X"4D",X"CB",
		X"C6",X"18",X"CA",X"7C",X"FE",X"42",X"20",X"05",X"7D",X"FE",X"E0",X"30",X"EF",X"DF",X"DF",X"18",
		X"E8",X"7D",X"E6",X"1F",X"FE",X"12",X"28",X"E4",X"7D",X"C6",X"03",X"6F",X"18",X"DB",X"7C",X"FE",
		X"41",X"20",X"05",X"7D",X"FE",X"60",X"38",X"D4",X"E7",X"E7",X"18",X"CD",X"2A",X"04",X"4D",X"7C",
		X"FE",X"42",X"20",X"11",X"7D",X"FE",X"F2",X"28",X"2F",X"FE",X"B2",X"28",X"2B",X"FE",X"72",X"28",
		X"40",X"FE",X"32",X"28",X"3C",X"EB",X"2A",X"06",X"4D",X"7C",X"FE",X"40",X"20",X"05",X"7D",X"FE",
		X"B5",X"28",X"A9",X"EB",X"2B",X"7E",X"2A",X"08",X"4D",X"77",X"23",X"22",X"08",X"4D",X"2A",X"06",
		X"4D",X"77",X"E7",X"22",X"06",X"4D",X"18",X"94",X"2A",X"06",X"4D",X"7C",X"FE",X"42",X"28",X"8C",
		X"36",X"3B",X"DF",X"22",X"06",X"4D",X"2A",X"08",X"4D",X"36",X"40",X"2B",X"22",X"08",X"4D",X"18",
		X"E5",X"CD",X"F0",X"26",X"CD",X"02",X"31",X"3E",X"FF",X"CD",X"10",X"1D",X"CD",X"D6",X"24",X"C3",
		X"AF",X"01",X"CD",X"6B",X"31",X"DD",X"21",X"00",X"4E",X"0E",X"01",X"3E",X"07",X"06",X"05",X"FD",
		X"21",X"A7",X"43",X"FD",X"E5",X"E1",X"11",X"00",X"04",X"19",X"CD",X"9D",X"31",X"FD",X"71",X"00",
		X"F5",X"DD",X"7E",X"0C",X"CD",X"A8",X"31",X"F1",X"FD",X"E5",X"E1",X"11",X"20",X"FF",X"19",X"DD",
		X"E5",X"D1",X"E5",X"EB",X"11",X"0F",X"00",X"19",X"EB",X"E1",X"C5",X"F5",X"06",X"03",X"CD",X"CB",
		X"31",X"F1",X"C1",X"DD",X"E5",X"D1",X"FD",X"E5",X"E1",X"D5",X"11",X"00",X"FE",X"19",X"D1",X"C5",
		X"F5",X"06",X"0C",X"1A",X"77",X"E7",X"13",X"10",X"FA",X"F1",X"C1",X"FD",X"23",X"FD",X"23",X"FD",
		X"23",X"11",X"10",X"00",X"DD",X"19",X"0C",X"3D",X"10",X"A9",X"C9",X"CD",X"00",X"01",X"11",X"89",
		X"31",X"21",X"45",X"41",X"CD",X"ED",X"01",X"11",X"8F",X"31",X"21",X"65",X"43",X"CD",X"ED",X"01",
		X"11",X"96",X"31",X"21",X"A5",X"42",X"C3",X"ED",X"01",X"12",X"4E",X"41",X"4D",X"45",X"FF",X"12",
		X"52",X"4F",X"55",X"4E",X"44",X"FF",X"12",X"53",X"43",X"4F",X"52",X"45",X"FF",X"F5",X"C5",X"06",
		X"1C",X"77",X"E7",X"10",X"FC",X"C1",X"F1",X"C9",X"F5",X"E6",X"F0",X"0F",X"0F",X"0F",X"0F",X"FD",
		X"77",X"A0",X"F1",X"E6",X"0F",X"FD",X"77",X"80",X"C9",X"1A",X"E6",X"F0",X"0F",X"0F",X"0F",X"0F",
		X"77",X"E7",X"1A",X"E6",X"0F",X"77",X"E7",X"1B",X"10",X"EF",X"C9",X"CD",X"B9",X"31",X"36",X"00",
		X"C9",X"4E",X"4F",X"4E",X"50",X"45",X"40",X"3D",X"40",X"40",X"40",X"40",X"40",X"03",X"70",X"32",
		X"00",X"54",X"41",X"4B",X"41",X"53",X"48",X"49",X"40",X"48",X"41",X"52",X"41",X"03",X"57",X"10",
		X"00",X"46",X"55",X"4D",X"49",X"4B",X"4F",X"40",X"59",X"41",X"4D",X"41",X"3D",X"01",X"60",X"09",
		X"00",X"52",X"45",X"49",X"4B",X"4F",X"40",X"49",X"5A",X"55",X"4D",X"49",X"40",X"01",X"54",X"05",
		X"00",X"41",X"54",X"53",X"55",X"4B",X"4F",X"40",X"4B",X"49",X"42",X"41",X"40",X"01",X"32",X"04",
		X"00",X"21",X"D1",X"31",X"11",X"00",X"4E",X"01",X"50",X"00",X"ED",X"B0",X"C9",X"06",X"A0",X"10",
		X"FE",X"CD",X"62",X"01",X"3A",X"2E",X"4C",X"06",X"F0",X"10",X"FE",X"C9",X"E5",X"F5",X"DD",X"E5",
		X"E1",X"7D",X"C6",X"FD",X"6F",X"46",X"F1",X"E1",X"80",X"DD",X"77",X"21",X"C9",X"3A",X"9A",X"4C",
		X"CB",X"4F",X"C0",X"3A",X"88",X"4C",X"C3",X"99",X"32",X"3E",X"FD",X"21",X"9A",X"4C",X"18",X"20",
		X"32",X"FD",X"4C",X"32",X"FE",X"4C",X"C3",X"9F",X"19",X"CB",X"CE",X"21",X"9A",X"4C",X"CB",X"8E",
		X"AF",X"18",X"1D",X"3D",X"32",X"9E",X"4C",X"C0",X"21",X"BE",X"4C",X"CB",X"96",X"AF",X"18",X"10",
		X"CB",X"CE",X"CD",X"60",X"32",X"00",X"00",X"21",X"00",X"00",X"22",X"07",X"4C",X"C3",X"9F",X"19",
		X"CD",X"60",X"32",X"CD",X"01",X"07",X"C3",X"9F",X"19",X"FE",X"01",X"28",X"BC",X"FE",X"00",X"3E",
		X"FC",X"28",X"B8",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"0D",
		X"0F",X"0F",X"0F",X"BC",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",
		X"0B",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"0C",
		X"0E",X"0E",X"0E",X"AB",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0D",X"0F",X"0F",X"BB",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"08",X"00",X"00",X"00",X"0B",
		X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"09",X"00",X"60",X"00",X"00",X"09",X"00",X"00",X"00",
		X"0C",X"0E",X"0E",X"BB",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"07",X"00",X"00",X"00",X"0A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"0F",X"6F",X"00",X"00",X"0B",X"00",X"00",X"00",
		X"0A",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",X"97",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"0C",X"0E",X"7E",X"00",X"00",X"0A",X"00",X"00",X"00",
		X"00",X"00",X"00",X"B8",X"00",X"00",X"F0",X"F0",X"D0",X"F0",X"F0",X"F0",X"F0",X"F8",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"D0",X"F0",X"F0",X"F0",X"FB",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"B6",X"00",X"00",X"E0",X"E0",X"C0",X"E0",X"E0",X"E0",X"E0",X"E6",X"E0",X"E0",
		X"E0",X"E0",X"E0",X"C8",X"E0",X"E0",X"E0",X"EA",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"E0",X"E0",X"E0",X"B6",X"00",X"00",X"00",X"00",X"B0",X"00",X"08",X"00",X"00",X"07",X"00",X"00",
		X"00",X"00",X"00",X"B6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"B6",X"00",X"00",X"00",X"00",X"A0",X"00",X"06",X"00",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"A6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",
		X"00",X"00",X"00",X"B6",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"0E",X"0E",X"0E",X"0E",
		X"0E",X"0E",X"0E",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"06",X"00",X"00",X"00",
		X"00",X"00",X"00",X"B6",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"60",X"07",X"00",X"00",X"00",
		X"00",X"00",X"00",X"B6",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"80",X"00",X"00",X"00",X"00",
		X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"B6",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"60",X"00",X"00",X"09",X"00",
		X"00",X"00",X"00",X"98",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"B6",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"70",X"00",X"00",X"0B",X"90",
		X"00",X"00",X"00",X"D6",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"90",X"00",X"00",X"B7",X"1E",X"C3",X"40",X"09",X"63",X"42",X"09",X"C8",X"42",X"09",X"4A",X"42",
		X"08",X"96",X"41",X"08",X"17",X"43",X"08",X"CE",X"42",X"07",X"2E",X"41",X"07",X"52",X"43",X"07",
		X"B2",X"42",X"06",X"77",X"42",X"06",X"43",X"41",X"06",X"C3",X"41",X"05",X"8C",X"41",X"05",X"89",
		X"43",X"05",X"CE",X"40",X"04",X"52",X"42",X"04",X"7B",X"42",X"04",X"49",X"40",X"03",X"25",X"43",
		X"03",X"CE",X"41",X"03",X"4E",X"40",X"02",X"43",X"42",X"02",X"4E",X"42",X"02",X"EA",X"41",X"01",
		X"D6",X"41",X"01",X"AE",X"43",X"01",X"4E",X"41",X"40",X"23",X"41",X"00",X"E8",X"42",X"00",X"06",
		X"94",X"40",X"7E",X"41",X"72",X"43",X"AC",X"41",X"C6",X"41",X"E5",X"42",X"E5",X"21",X"00",X"25",
		X"22",X"85",X"4C",X"E1",X"C3",X"8F",X"20",X"CB",X"6F",X"C0",X"CB",X"77",X"C0",X"79",X"FE",X"01",
		X"CA",X"DC",X"25",X"A7",X"C0",X"C3",X"DE",X"1C",X"CD",X"9C",X"19",X"3E",X"10",X"CD",X"10",X"1D",
		X"C3",X"DC",X"25",X"21",X"C9",X"43",X"11",X"8F",X"31",X"CD",X"D5",X"01",X"3A",X"40",X"4C",X"2E",
		X"E6",X"47",X"E6",X"0F",X"77",X"23",X"78",X"E6",X"F0",X"0F",X"0F",X"0F",X"0F",X"77",X"11",X"EF",
		X"43",X"21",X"0F",X"4E",X"AF",X"12",X"1E",X"F5",X"CD",X"09",X"13",X"C3",X"E6",X"25",X"AF",X"32",
		X"2D",X"4C",X"3C",X"32",X"40",X"4C",X"CD",X"CF",X"9B",X"CD",X"00",X"01",X"CD",X"52",X"09",X"CD",
		X"12",X"0D",X"CD",X"5B",X"35",X"CD",X"77",X"35",X"CD",X"9F",X"36",X"CD",X"D6",X"9B",X"06",X"0E",
		X"CD",X"45",X"35",X"18",X"F0",X"3A",X"26",X"4C",X"A7",X"20",X"03",X"10",X"F8",X"C9",X"21",X"30",
		X"4C",X"06",X"0C",X"36",X"00",X"23",X"10",X"FB",X"C3",X"0D",X"90",X"CD",X"E0",X"06",X"CB",X"86",
		X"3E",X"30",X"CD",X"C1",X"01",X"AF",X"32",X"44",X"4C",X"3C",X"32",X"81",X"4C",X"32",X"42",X"4C",
		X"21",X"08",X"37",X"CD",X"99",X"37",X"C9",X"3A",X"41",X"4C",X"A7",X"28",X"05",X"3D",X"32",X"41",
		X"4C",X"C9",X"3E",X"40",X"32",X"41",X"4C",X"3A",X"43",X"4C",X"A7",X"C2",X"14",X"36",X"2A",X"45",
		X"4C",X"3A",X"42",X"4C",X"3D",X"28",X"03",X"23",X"18",X"FA",X"3A",X"42",X"4C",X"3C",X"32",X"42",
		X"4C",X"7E",X"47",X"E6",X"0F",X"32",X"47",X"4C",X"78",X"E6",X"F0",X"C2",X"F8",X"35",X"CD",X"0E",
		X"36",X"3E",X"08",X"32",X"43",X"4C",X"C9",X"AF",X"CD",X"0E",X"36",X"3A",X"47",X"4C",X"FE",X"01",
		X"28",X"0B",X"CD",X"26",X"36",X"3E",X"01",X"32",X"01",X"50",X"C9",X"AE",X"35",X"AF",X"CD",X"D6",
		X"24",X"CD",X"42",X"36",X"18",X"EF",X"AF",X"CD",X"D6",X"24",X"3A",X"47",X"4C",X"FE",X"01",X"3A",
		X"44",X"4C",X"CB",X"9F",X"20",X"02",X"CB",X"DF",X"CB",X"FF",X"CB",X"8F",X"32",X"44",X"4C",X"3E",
		X"20",X"32",X"43",X"4C",X"00",X"00",X"00",X"C9",X"CB",X"77",X"20",X"0B",X"CB",X"6F",X"20",X"B7",
		X"CB",X"67",X"20",X"D2",X"C3",X"6E",X"37",X"21",X"44",X"4C",X"CB",X"CE",X"18",X"A3",X"21",X"44",
		X"4C",X"CB",X"8E",X"C9",X"F5",X"3A",X"44",X"4C",X"CB",X"4F",X"20",X"04",X"00",X"C3",X"79",X"37",
		X"F1",X"3D",X"32",X"43",X"4C",X"C9",X"CD",X"0E",X"07",X"23",X"E7",X"E7",X"7E",X"FE",X"0A",X"CD",
		X"5B",X"36",X"22",X"51",X"4C",X"CD",X"E4",X"0A",X"CB",X"D6",X"CB",X"9E",X"3E",X"0C",X"32",X"FC",
		X"4F",X"C9",X"CD",X"0E",X"07",X"23",X"DF",X"7E",X"FE",X"0A",X"CD",X"7A",X"36",X"22",X"51",X"4C",
		X"CD",X"E4",X"0A",X"CB",X"D6",X"CB",X"DE",X"3E",X"0E",X"18",X"E3",X"30",X"19",X"E5",X"E7",X"7E",
		X"FE",X"0A",X"E1",X"38",X"02",X"2B",X"C9",X"C1",X"2B",X"22",X"51",X"4C",X"CD",X"B0",X"0A",X"CB",
		X"EE",X"CB",X"96",X"C3",X"3A",X"36",X"E1",X"C3",X"3C",X"36",X"30",X"19",X"E5",X"DF",X"7E",X"FE",
		X"0A",X"E1",X"38",X"02",X"2B",X"C9",X"C1",X"2B",X"22",X"51",X"4C",X"CD",X"B0",X"0A",X"CB",X"EE",
		X"CB",X"96",X"C3",X"55",X"36",X"E1",X"C3",X"57",X"36",X"CD",X"0C",X"0A",X"C3",X"14",X"10",X"3A",
		X"44",X"4C",X"CB",X"67",X"C8",X"21",X"30",X"4C",X"06",X"08",X"36",X"00",X"23",X"10",X"FB",X"3E",
		X"20",X"CD",X"C1",X"01",X"3A",X"FD",X"4F",X"32",X"7E",X"4F",X"3E",X"11",X"32",X"FD",X"4F",X"06",
		X"10",X"3E",X"80",X"32",X"FC",X"4F",X"3E",X"05",X"CD",X"C1",X"01",X"3E",X"84",X"32",X"FC",X"4F",
		X"3E",X"05",X"CD",X"C1",X"01",X"10",X"EA",X"3E",X"80",X"CD",X"C1",X"01",X"C1",X"C9",X"F5",X"3A",
		X"44",X"4C",X"CB",X"E7",X"32",X"44",X"4C",X"F1",X"C9",X"DD",X"5E",X"00",X"DD",X"56",X"01",X"2A",
		X"3A",X"4C",X"7C",X"92",X"F2",X"F9",X"36",X"ED",X"44",X"FE",X"09",X"D0",X"7D",X"93",X"F2",X"03",
		X"37",X"ED",X"44",X"FE",X"09",X"38",X"D7",X"C9",X"01",X"01",X"00",X"00",X"00",X"01",X"01",X"21",
		X"40",X"01",X"21",X"40",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"40",X"40",
		X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"01",X"21",X"40",X"40",X"01",X"03",X"03",X"00",X"00",
		X"00",X"00",X"00",X"40",X"02",X"02",X"02",X"02",X"02",X"01",X"01",X"01",X"11",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"13",X"01",X"00",X"00",X"00",X"00",
		X"23",X"40",X"03",X"03",X"23",X"40",X"03",X"03",X"03",X"13",X"03",X"03",X"23",X"03",X"02",X"02",
		X"02",X"02",X"03",X"13",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"80",X"21",X"44",
		X"4C",X"CB",X"C6",X"3E",X"F0",X"32",X"43",X"4C",X"C9",X"CB",X"47",X"20",X"04",X"F1",X"C3",X"99",
		X"08",X"F1",X"3D",X"32",X"43",X"4C",X"3A",X"3B",X"4C",X"3D",X"32",X"3B",X"4C",X"CD",X"0E",X"07",
		X"23",X"23",X"7E",X"FE",X"F6",X"D8",X"C3",X"DE",X"36",X"ED",X"5F",X"CB",X"4F",X"28",X"03",X"21",
		X"A6",X"37",X"22",X"45",X"4C",X"C9",X"03",X"03",X"03",X"00",X"00",X"00",X"03",X"21",X"01",X"01",
		X"11",X"01",X"01",X"23",X"03",X"03",X"00",X"00",X"00",X"00",X"40",X"40",X"40",X"40",X"40",X"40",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"23",X"03",
		X"03",X"03",X"03",X"23",X"01",X"11",X"03",X"23",X"40",X"03",X"40",X"40",X"40",X"40",X"40",X"40",
		X"40",X"40",X"40",X"40",X"03",X"23",X"03",X"03",X"23",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"11",X"01",X"01",X"01",X"11",X"01",X"01",X"11",X"80",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
