library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity obj2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of obj2 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"E3",X"F3",X"FB",X"B9",X"10",X"43",X"83",X"83",X"01",X"00",X"00",X"00",X"00",
		X"E0",X"E6",X"C7",X"87",X"C1",X"C0",X"00",X"40",X"00",X"80",X"80",X"C0",X"DC",X"FC",X"C0",X"00",
		X"1E",X"1C",X"20",X"60",X"C0",X"C0",X"E0",X"E3",X"E3",X"63",X"61",X"E0",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"07",X"07",X"87",X"83",X"0B",X"08",X"08",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"0F",X"0F",X"0F",X"37",X"33",X"30",X"20",X"00",X"00",X"00",X"00",
		X"C0",X"C0",X"00",X"00",X"0C",X"0E",X"0E",X"06",X"44",X"40",X"40",X"40",X"40",X"40",X"40",X"00",
		X"60",X"E0",X"E0",X"81",X"01",X"01",X"81",X"C1",X"C1",X"81",X"01",X"01",X"81",X"E0",X"E0",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"C3",X"C3",X"C1",X"80",X"43",X"03",X"83",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"C3",X"E3",X"E3",X"C1",X"C0",X"C3",X"C3",X"C3",X"C1",X"E0",X"E0",X"E0",X"C0",
		X"00",X"06",X"07",X"03",X"C1",X"C0",X"C0",X"00",X"40",X"00",X"00",X"00",X"1C",X"3C",X"00",X"00",
		X"00",X"06",X"07",X"03",X"C1",X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",X"C0",X"FC",X"FC",X"E0",X"C0",
		X"1E",X"1C",X"00",X"00",X"C0",X"C0",X"E0",X"E3",X"C3",X"A3",X"81",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"1C",X"00",X"00",X"C0",X"C0",X"E0",X"E3",X"E3",X"63",X"E1",X"60",X"60",X"E0",X"E0",X"C0",
		X"84",X"8C",X"D8",X"9C",X"C8",X"E0",X"E0",X"00",X"20",X"80",X"C0",X"40",X"40",X"C0",X"CC",X"9C",
		X"C1",X"E5",X"42",X"82",X"C1",X"C0",X"80",X"41",X"03",X"87",X"8E",X"8D",X"83",X"C6",X"CC",X"C0",
		X"00",X"20",X"70",X"58",X"7B",X"7F",X"1F",X"2F",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"A8",X"B8",X"B0",X"38",X"60",X"40",X"C0",X"80",X"D0",X"F0",X"E0",X"40",X"00",
		X"80",X"40",X"E0",X"F0",X"E0",X"C0",X"40",X"40",X"40",X"68",X"78",X"F8",X"D0",X"40",X"00",X"00",
		X"00",X"40",X"40",X"68",X"38",X"20",X"B8",X"A0",X"A0",X"B8",X"B0",X"38",X"68",X"40",X"40",X"00",
		X"40",X"C0",X"DC",X"FF",X"FF",X"C7",X"02",X"00",X"00",X"00",X"00",X"E0",X"F0",X"F0",X"60",X"00",
		X"00",X"00",X"C0",X"20",X"10",X"10",X"08",X"88",X"48",X"08",X"10",X"10",X"20",X"C0",X"00",X"00",
		X"40",X"F0",X"20",X"20",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"20",X"20",X"F0",X"40",
		X"A0",X"F0",X"D0",X"D8",X"C8",X"C8",X"C8",X"C8",X"C8",X"C8",X"C8",X"C8",X"D8",X"D0",X"F0",X"A0",
		X"00",X"00",X"00",X"00",X"F2",X"FE",X"03",X"02",X"02",X"03",X"FF",X"F2",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"C0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"C0",X"00",X"00",X"00",
		X"A0",X"F0",X"D0",X"D8",X"C8",X"C8",X"C8",X"C8",X"C8",X"C8",X"C8",X"C8",X"D8",X"D0",X"F0",X"A0",
		X"40",X"F0",X"20",X"20",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"20",X"20",X"F0",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"02",X"08",X"04",X"02",X"F8",X"FC",X"FC",X"FC",X"FC",X"FC",X"FA",X"02",X"0A",X"14",X"02",
		X"33",X"39",X"78",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7C",X"3D",X"19",X"03",
		X"33",X"39",X"78",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7C",X"3D",X"19",X"03",
		X"33",X"39",X"78",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7C",X"3D",X"19",X"03",
		X"1F",X"27",X"47",X"43",X"43",X"43",X"43",X"43",X"43",X"43",X"43",X"43",X"47",X"27",X"1F",X"1F",
		X"6F",X"F7",X"F7",X"73",X"7B",X"7B",X"7B",X"73",X"7B",X"7B",X"7B",X"73",X"F7",X"F7",X"67",X"0F",
		X"00",X"00",X"C0",X"C0",X"40",X"C0",X"C0",X"40",X"C0",X"40",X"C0",X"40",X"C0",X"C0",X"00",X"00",
		X"E0",X"E0",X"E0",X"E0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F4",X"F0",X"F0",X"28",X"00",X"00",X"00",
		X"00",X"01",X"02",X"E4",X"F8",X"FA",X"FC",X"FC",X"FC",X"F8",X"FA",X"FC",X"F8",X"F8",X"30",X"20",
		X"C0",X"E0",X"F0",X"F0",X"F8",X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",
		X"00",X"05",X"02",X"07",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FC",X"F8",X"F0",
		X"00",X"00",X"00",X"00",X"03",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"60",X"B0",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"78",X"00",X"CC",X"F8",X"FE",X"FD",X"FC",X"F9",X"F8",X"F8",X"F8",
		X"FC",X"F8",X"FC",X"FC",X"32",X"84",X"C3",X"F0",X"F8",X"F0",X"F0",X"A0",X"04",X"02",X"00",X"00",
		X"F8",X"F8",X"F8",X"F0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E6",X"FC",X"78",X"F8",X"FC",
		X"00",X"01",X"07",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"3F",X"9F",X"CF",X"E3",X"C1",X"80",X"08",X"10",X"20",X"20",X"20",X"20",X"20",X"00",
		X"60",X"F0",X"F8",X"FC",X"FC",X"FE",X"FC",X"EC",X"CE",X"CE",X"C0",X"C0",X"E0",X"E0",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0B",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0B",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"FF",X"FE",X"FC",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F8",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"18",X"30",X"F6",X"F7",X"F7",X"F3",X"FB",X"F9",X"FC",X"E4",X"C2",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"30",X"70",X"F0",X"F0",X"E0",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"49",X"2A",X"08",X"7E",X"08",X"2A",X"49",X"80",X"00",X"02",X"09",X"80",X"08",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"81",X"C3",X"E3",X"33",X"1B",X"AF",X"AF",X"1B",X"33",X"E3",X"C3",X"81",X"00",X"00",
		X"20",X"70",X"71",X"53",X"DB",X"8B",X"8B",X"FF",X"FF",X"8B",X"8B",X"DB",X"53",X"71",X"70",X"20",
		X"00",X"00",X"00",X"00",X"00",X"78",X"FC",X"CC",X"FC",X"FC",X"CC",X"78",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"78",X"FC",X"FE",X"CE",X"FE",X"FE",X"CC",X"FC",X"78",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"18",X"38",X"9F",X"37",X"25",X"09",X"5E",X"17",X"0E",X"10",X"21",X"0F",X"13",X"04",X"00",
		X"00",X"00",X"00",X"07",X"13",X"03",X"38",X"7F",X"07",X"00",X"02",X"43",X"07",X"06",X"10",X"00",
		X"20",X"04",X"02",X"0B",X"37",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F9",X"13",X"21",X"42",X"00",
		X"00",X"00",X"03",X"03",X"7F",X"FF",X"7F",X"7F",X"FF",X"FF",X"7F",X"7F",X"8D",X"00",X"22",X"00",
		X"60",X"E0",X"A0",X"20",X"20",X"20",X"A0",X"E0",X"60",X"E0",X"A0",X"20",X"20",X"20",X"A0",X"E0",
		X"FE",X"FF",X"FF",X"83",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"83",X"FF",X"FF",X"FE",
		X"00",X"00",X"00",X"FF",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"DF",X"5F",X"5F",X"5F",X"DF",X"5F",X"5F",X"DF",X"5F",X"5F",X"5F",X"DF",X"FF",X"DF",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"70",X"70",X"70",X"70",X"F0",X"70",X"70",X"70",X"F0",X"70",X"70",X"F0",X"70",X"70",X"E0",
		X"00",X"00",X"20",X"70",X"10",X"00",X"00",X"20",X"70",X"A8",X"F4",X"52",X"7A",X"34",X"00",X"00",
		X"00",X"20",X"10",X"08",X"0C",X"DE",X"FE",X"FE",X"FE",X"7C",X"F8",X"78",X"F0",X"80",X"00",X"00",
		X"00",X"00",X"10",X"08",X"08",X"FC",X"FC",X"FE",X"FE",X"7E",X"FE",X"7E",X"FC",X"98",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F8",X"F8",X"F8",X"F8",X"78",X"38",X"38",X"F0",X"F0",X"E0",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"F8",X"F8",X"78",X"78",X"78",X"78",X"78",X"70",X"70",X"E0",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"F8",X"F8",X"F8",X"38",X"38",X"78",X"F8",X"F0",X"F0",X"E0",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"20",X"10",X"08",X"04",X"04",X"04",X"04",X"04",X"04",X"08",X"10",X"20",X"C0",X"00",
		X"00",X"00",X"00",X"80",X"40",X"A0",X"50",X"50",X"50",X"50",X"A0",X"40",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"A0",X"A0",X"40",X"80",X"00",X"00",X"00",X"00",X"00",
		X"82",X"84",X"00",X"00",X"00",X"00",X"00",X"00",X"9A",X"00",X"00",X"00",X"00",X"00",X"84",X"82",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",
		X"04",X"02",X"84",X"54",X"12",X"12",X"12",X"12",X"14",X"14",X"14",X"12",X"02",X"02",X"04",X"00",
		X"00",X"00",X"00",X"00",X"DE",X"2E",X"76",X"6A",X"6A",X"6A",X"76",X"2E",X"DE",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"C0",X"E0",X"F0",X"F0",X"F8",X"FC",X"FE",X"FC",X"F8",X"F0",X"F0",X"E0",X"C0",X"00",X"00",
		X"00",X"C0",X"E0",X"F0",X"F0",X"F8",X"F4",X"E0",X"4A",X"1C",X"B8",X"F0",X"F0",X"E0",X"C0",X"00",
		X"38",X"BC",X"9C",X"CC",X"80",X"40",X"00",X"80",X"80",X"00",X"46",X"86",X"CE",X"8C",X"8C",X"00",
		X"00",X"00",X"F0",X"F8",X"FC",X"FE",X"33",X"DF",X"DE",X"88",X"20",X"03",X"07",X"0F",X"0E",X"0C",
		X"00",X"00",X"1F",X"7F",X"FF",X"7F",X"3F",X"2F",X"5E",X"0F",X"47",X"07",X"07",X"0F",X"07",X"03",
		X"C0",X"20",X"20",X"20",X"C0",X"00",X"C0",X"20",X"20",X"20",X"C0",X"00",X"20",X"E0",X"20",X"00",
		X"C0",X"20",X"20",X"C0",X"00",X"C0",X"20",X"20",X"C0",X"00",X"20",X"20",X"A0",X"60",X"20",X"00",
		X"C0",X"20",X"20",X"C0",X"00",X"C0",X"20",X"20",X"C0",X"00",X"C0",X"20",X"20",X"20",X"20",X"00",
		X"C0",X"20",X"20",X"C0",X"00",X"C0",X"20",X"20",X"C0",X"00",X"C0",X"20",X"20",X"20",X"40",X"00",
		X"C0",X"20",X"20",X"C0",X"00",X"C0",X"20",X"20",X"C0",X"00",X"C0",X"20",X"20",X"20",X"C0",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
