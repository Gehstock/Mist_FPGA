library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity kick_sp_bits_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of kick_sp_bits_1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"E0",X"00",X"EE",X"00",X"0E",X"00",X"EE",X"00",X"00",X"00",
		X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"0E",X"00",X"00",X"0E",X"E0",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"E0",X"00",X"00",X"00",X"0E",X"10",X"00",X"00",X"00",
		X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"11",X"00",X"00",X"0E",X"11",X"00",X"00",X"EE",
		X"11",X"00",X"00",X"E0",X"11",X"E0",X"00",X"00",X"11",X"EE",X"00",X"00",X"11",X"0E",X"EE",X"00",
		X"10",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",
		X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",
		X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",
		X"70",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",X"00",X"EE",X"00",
		X"00",X"0E",X"EE",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"E0",
		X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"0E",X"00",X"00",X"E0",X"0E",X"00",X"00",X"00",
		X"0E",X"E0",X"00",X"00",X"EE",X"0E",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",
		X"EE",X"00",X"00",X"00",X"EE",X"00",X"0E",X"00",X"EE",X"EE",X"E0",X"00",X"EE",X"EE",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"0E",X"EE",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"E0",
		X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"7E",X"00",X"00",X"E0",X"77",X"D0",X"88",X"00",
		X"77",X"D0",X"88",X"00",X"77",X"DE",X"88",X"00",X"77",X"D0",X"88",X"00",X"77",X"00",X"88",X"00",
		X"77",X"00",X"88",X"00",X"75",X"00",X"8E",X"00",X"77",X"2E",X"E8",X"00",X"77",X"2E",X"EE",X"EE",
		X"FF",X"33",X"77",X"77",X"FF",X"43",X"77",X"77",X"55",X"44",X"77",X"77",X"55",X"44",X"77",X"77",
		X"05",X"44",X"77",X"77",X"00",X"44",X"77",X"77",X"00",X"44",X"77",X"77",X"00",X"44",X"07",X"77",
		X"00",X"04",X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"33",X"77",X"77",X"55",X"33",X"77",X"77",X"55",X"33",X"77",X"72",X"FF",X"33",X"77",X"72",
		X"55",X"33",X"77",X"72",X"55",X"33",X"77",X"22",X"05",X"00",X"77",X"22",X"00",X"00",X"07",X"22",
		X"00",X"40",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"55",X"00",X"00",X"44",X"FF",X"00",
		X"00",X"44",X"55",X"00",X"00",X"44",X"55",X"B0",X"00",X"44",X"FF",X"00",X"00",X"44",X"55",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"33",X"77",X"77",X"55",X"33",X"77",X"77",X"FF",X"33",X"B7",X"77",X"55",X"33",X"BB",X"77",
		X"55",X"33",X"BB",X"77",X"05",X"43",X"BB",X"22",X"00",X"43",X"BB",X"22",X"00",X"44",X"07",X"22",
		X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"44",X"BB",X"00",X"00",X"44",X"BB",
		X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AB",X"00",X"00",X"00",X"AB",X"00",X"00",X"00",X"AA",
		X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"B7",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"B6",X"00",X"00",X"44",X"66",X"00",X"00",X"44",X"BB",
		X"00",X"00",X"00",X"BA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",
		X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"00",X"B6",X"00",X"00",X"00",X"B6",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"00",X"AA",X"00",X"00",X"44",X"AB",X"00",X"00",X"44",X"AB",X"00",X"00",X"00",X"AA",
		X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",
		X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"40",X"00",X"01",X"11",
		X"40",X"00",X"07",X"11",X"44",X"00",X"77",X"77",X"44",X"00",X"77",X"77",X"44",X"05",X"77",X"77",
		X"44",X"33",X"77",X"77",X"44",X"33",X"77",X"77",X"44",X"33",X"77",X"77",X"05",X"33",X"77",X"77",
		X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",
		X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"77",X"00",X"00",X"DD",X"77",X"00",X"00",X"DD",X"77",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",
		X"00",X"B0",X"00",X"77",X"00",X"B0",X"00",X"77",X"00",X"B0",X"00",X"77",X"00",X"B0",X"00",X"77",
		X"00",X"B0",X"00",X"77",X"00",X"BB",X"00",X"77",X"00",X"0B",X"00",X"77",X"00",X"0B",X"00",X"77",
		X"00",X"BB",X"00",X"77",X"00",X"BB",X"00",X"77",X"00",X"BB",X"00",X"77",X"00",X"BB",X"00",X"77",
		X"00",X"BB",X"00",X"77",X"00",X"FF",X"00",X"77",X"00",X"FF",X"00",X"77",X"00",X"FF",X"00",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"E0",X"00",X"EE",X"00",X"0E",X"00",X"EE",X"00",X"00",X"00",
		X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"0E",X"00",X"00",X"0E",X"E0",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"E0",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"E0",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"EE",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"5F",X"22",X"E0",X"00",X"5F",X"22",X"0E",X"00",X"05",X"77",X"00",X"00",X"EE",X"77",X"00",X"00",
		X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"0E",X"00",X"00",X"0E",X"E0",X"00",X"00",
		X"0E",X"00",X"00",X"E0",X"0E",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"EE",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"EE",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"EE",X"EE",X"EE",X"77",X"EE",X"0E",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",
		X"77",X"0E",X"00",X"00",X"EE",X"E0",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"EE",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"EE",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",
		X"00",X"0B",X"00",X"77",X"00",X"BB",X"00",X"77",X"00",X"BB",X"00",X"77",X"00",X"BB",X"00",X"77",
		X"00",X"BB",X"00",X"77",X"00",X"05",X"00",X"77",X"00",X"0F",X"00",X"77",X"00",X"04",X"00",X"70",
		X"00",X"04",X"00",X"70",X"05",X"34",X"00",X"70",X"05",X"33",X"77",X"77",X"55",X"33",X"77",X"77",
		X"FF",X"33",X"77",X"77",X"55",X"33",X"77",X"77",X"55",X"34",X"77",X"77",X"FF",X"44",X"77",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"B5",X"00",X"00",X"00",X"5F",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"F5",X"00",
		X"00",X"00",X"45",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"40",X"01",X"00",X"00",X"07",X"71",
		X"00",X"00",X"77",X"71",X"05",X"00",X"77",X"71",X"05",X"33",X"77",X"77",X"55",X"33",X"77",X"77",
		X"FF",X"33",X"77",X"77",X"55",X"33",X"77",X"77",X"55",X"33",X"77",X"77",X"CF",X"33",X"77",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"11",
		X"00",X"0B",X"00",X"11",X"00",X"BB",X"00",X"11",X"00",X"BB",X"00",X"11",X"00",X"BB",X"00",X"11",
		X"00",X"BF",X"00",X"11",X"00",X"5F",X"00",X"11",X"00",X"F5",X"00",X"11",X"00",X"54",X"00",X"11",
		X"00",X"04",X"00",X"11",X"00",X"04",X"00",X"11",X"00",X"00",X"07",X"11",X"00",X"00",X"07",X"71",
		X"00",X"00",X"77",X"77",X"05",X"03",X"77",X"77",X"05",X"33",X"77",X"77",X"55",X"33",X"77",X"77",
		X"FF",X"33",X"77",X"77",X"55",X"33",X"77",X"77",X"55",X"33",X"77",X"77",X"CF",X"33",X"77",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"0B",X"00",X"00",
		X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"07",X"00",X"04",X"00",X"07",X"00",X"04",X"00",X"77",X"00",X"44",X"07",X"77",
		X"00",X"33",X"77",X"77",X"05",X"33",X"77",X"77",X"05",X"33",X"77",X"77",X"55",X"33",X"77",X"77",
		X"FF",X"33",X"77",X"77",X"FF",X"33",X"77",X"77",X"55",X"33",X"77",X"77",X"55",X"33",X"77",X"77",
		X"00",X"00",X"00",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",
		X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"D0",
		X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"5B",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"F5",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"4F",X"00",X"00",X"00",X"4F",X"00",
		X"00",X"00",X"40",X"00",X"00",X"44",X"00",X"07",X"00",X"44",X"00",X"77",X"00",X"44",X"00",X"77",
		X"00",X"44",X"00",X"77",X"05",X"44",X"00",X"77",X"55",X"44",X"00",X"77",X"FF",X"44",X"00",X"77",
		X"55",X"40",X"07",X"77",X"55",X"33",X"F7",X"77",X"FF",X"33",X"F7",X"77",X"55",X"33",X"F7",X"77",
		X"55",X"33",X"F7",X"77",X"FF",X"33",X"F7",X"77",X"55",X"33",X"F7",X"77",X"55",X"40",X"07",X"77",
		X"FF",X"44",X"00",X"11",X"55",X"44",X"00",X"11",X"05",X"44",X"00",X"11",X"00",X"44",X"00",X"11",
		X"00",X"44",X"00",X"11",X"00",X"44",X"00",X"01",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",
		X"BB",X"FF",X"00",X"00",X"00",X"55",X"00",X"11",X"00",X"FF",X"00",X"11",X"00",X"55",X"00",X"11",
		X"00",X"55",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"05",X"00",X"00",X"00",X"55",X"DD",X"00",X"00",X"DB",X"DD",X"00",X"00",X"DB",X"DD",
		X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",
		X"77",X"77",X"5B",X"00",X"77",X"77",X"FB",X"00",X"77",X"77",X"50",X"00",X"77",X"EE",X"E0",X"EE",
		X"7E",X"E0",X"0E",X"00",X"EE",X"00",X"0E",X"00",X"EE",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"0E",X"00",X"00",X"0E",X"0E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"EE",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"EE",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"FB",X"D0",X"00",X"EE",X"FB",X"E0",X"00",X"EE",X"00",X"0E",X"00",X"EE",X"0D",X"00",X"00",
		X"EE",X"0D",X"00",X"00",X"EE",X"0D",X"00",X"00",X"EE",X"0E",X"E0",X"E0",X"0E",X"E0",X"E0",X"0E",
		X"0E",X"00",X"E0",X"00",X"0E",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"EE",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"EE",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"0E",X"EE",X"00",X"70",X"EE",X"00",X"00",X"70",X"E0",X"00",X"00",X"77",X"00",X"00",X"EE",
		X"77",X"00",X"00",X"EE",X"77",X"00",X"00",X"EE",X"77",X"00",X"00",X"00",X"77",X"00",X"8E",X"00",
		X"77",X"00",X"8E",X"00",X"77",X"00",X"8E",X"00",X"77",X"00",X"8E",X"00",X"77",X"00",X"E8",X"00",
		X"77",X"E0",X"E8",X"0E",X"77",X"7E",X"E8",X"E0",X"77",X"70",X"F5",X"00",X"EE",X"70",X"5F",X"00",
		X"EE",X"7F",X"DD",X"00",X"EE",X"5F",X"DD",X"00",X"EE",X"55",X"DD",X"00",X"EE",X"F5",X"DD",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"0E",X"EE",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"EE",X"30",X"00",X"00",X"EE",X"33",X"00",X"00",X"E0",X"33",X"00",X"00",X"00",
		X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"3E",X"00",X"DD",X"00",X"3E",X"00",X"DD",X"00",
		X"3E",X"00",X"DD",X"00",X"EE",X"00",X"DD",X"00",X"7E",X"E0",X"DD",X"00",X"77",X"7E",X"BB",X"00",
		X"77",X"77",X"FB",X"00",X"77",X"77",X"5F",X"00",X"77",X"77",X"FE",X"00",X"77",X"77",X"E8",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"0E",X"EE",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"E0",X"00",X"00",X"30",X"EE",X"00",X"00",X"3E",X"8E",X"00",X"00",X"3E",X"8E",X"00",X"00",
		X"3E",X"88",X"00",X"00",X"EE",X"88",X"00",X"00",X"EE",X"88",X"0E",X"00",X"7E",X"E8",X"0E",X"00",
		X"77",X"EE",X"E0",X"EE",X"77",X"77",X"50",X"00",X"77",X"77",X"FB",X"00",X"77",X"77",X"5B",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"BB",X"04",X"00",X"00",X"BB",X"44",X"00",X"00",X"BB",X"44",X"00",X"00",X"00",X"44",
		X"00",X"00",X"0B",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"44",X"BB",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"A0",
		X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",
		X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"44",X"BB",
		X"55",X"53",X"77",X"77",X"FF",X"33",X"77",X"77",X"55",X"33",X"77",X"77",X"55",X"33",X"77",X"77",
		X"FF",X"33",X"77",X"77",X"55",X"00",X"77",X"22",X"05",X"00",X"07",X"22",X"00",X"40",X"07",X"22",
		X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"40",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",
		X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",
		X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"40",X"00",X"00",
		X"00",X"40",X"07",X"22",X"05",X"00",X"07",X"22",X"55",X"00",X"77",X"22",X"FF",X"33",X"77",X"77",
		X"55",X"33",X"77",X"77",X"55",X"33",X"77",X"77",X"FF",X"33",X"77",X"77",X"55",X"53",X"77",X"77",
		X"55",X"44",X"77",X"77",X"55",X"44",X"77",X"77",X"FF",X"44",X"77",X"72",X"55",X"44",X"77",X"72",
		X"55",X"44",X"77",X"72",X"05",X"44",X"77",X"22",X"05",X"43",X"77",X"22",X"00",X"33",X"07",X"22",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"40",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",
		X"00",X"04",X"44",X"44",X"00",X"04",X"44",X"44",X"00",X"04",X"44",X"44",X"00",X"04",X"44",X"44",
		X"00",X"04",X"44",X"44",X"00",X"04",X"44",X"44",X"00",X"04",X"44",X"44",X"00",X"00",X"44",X"44",
		X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"40",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"00",X"77",X"00",X"44",X"00",X"77",X"00",X"44",X"00",X"77",X"00",X"44",X"00",X"77",
		X"00",X"44",X"03",X"77",X"00",X"44",X"33",X"77",X"00",X"44",X"33",X"77",X"00",X"44",X"33",X"77",
		X"00",X"44",X"33",X"77",X"00",X"44",X"33",X"77",X"00",X"44",X"53",X"70",X"00",X"44",X"35",X"00",
		X"00",X"44",X"53",X"00",X"00",X"44",X"33",X"00",X"00",X"43",X"33",X"00",X"00",X"33",X"33",X"00",
		X"00",X"33",X"33",X"00",X"00",X"33",X"33",X"00",X"00",X"33",X"33",X"00",X"00",X"3B",X"33",X"00",
		X"00",X"3A",X"34",X"00",X"00",X"33",X"34",X"44",X"00",X"BB",X"44",X"44",X"00",X"BB",X"44",X"44",
		X"04",X"BB",X"44",X"44",X"04",X"BB",X"44",X"44",X"04",X"AB",X"44",X"00",X"04",X"BB",X"44",X"00",
		X"04",X"AA",X"40",X"00",X"04",X"AA",X"00",X"00",X"04",X"4A",X"00",X"00",X"44",X"00",X"00",X"00",
		X"77",X"77",X"DD",X"00",X"77",X"77",X"DD",X"00",X"77",X"70",X"DD",X"00",X"77",X"00",X"DD",X"00",
		X"77",X"00",X"0D",X"0E",X"77",X"00",X"E0",X"EE",X"77",X"00",X"00",X"EE",X"77",X"00",X"00",X"E0",
		X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",
		X"00",X"EE",X"EE",X"00",X"00",X"EE",X"E0",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",
		X"55",X"B0",X"00",X"00",X"FF",X"00",X"00",X"00",X"55",X"BB",X"00",X"00",X"55",X"00",X"00",X"00",
		X"FF",X"BB",X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"E0",
		X"00",X"00",X"0E",X"EE",X"00",X"00",X"0E",X"EE",X"00",X"00",X"0E",X"EE",X"00",X"0E",X"0E",X"0E",
		X"00",X"EE",X"0E",X"0E",X"00",X"EE",X"0E",X"00",X"00",X"E0",X"0E",X"00",X"00",X"00",X"0E",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"0E",X"00",X"00",X"0E",X"E0",
		X"00",X"00",X"0E",X"E0",X"00",X"00",X"0E",X"00",X"00",X"E0",X"0E",X"00",X"00",X"0E",X"0E",X"00",
		X"00",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"EE",X"00",X"0E",X"00",
		X"EE",X"00",X"DE",X"00",X"EE",X"05",X"DD",X"00",X"EE",X"55",X"DD",X"00",X"77",X"5F",X"DD",X"EE",
		X"33",X"33",X"00",X"05",X"33",X"44",X"40",X"55",X"03",X"44",X"44",X"5F",X"03",X"44",X"44",X"F5",
		X"00",X"44",X"44",X"55",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"00",X"00",
		X"00",X"45",X"00",X"00",X"00",X"5F",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"5F",X"00",X"00",
		X"AA",X"BB",X"00",X"00",X"AA",X"BB",X"00",X"E0",X"AA",X"BB",X"00",X"0E",X"00",X"BB",X"00",X"0E",
		X"00",X"BB",X"44",X"EE",X"00",X"BA",X"44",X"EE",X"00",X"BA",X"44",X"E0",X"00",X"B6",X"44",X"00",
		X"00",X"B6",X"44",X"50",X"00",X"BB",X"44",X"0B",X"00",X"B0",X"04",X"BB",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"D0",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",
		X"00",X"B0",X"D0",X"00",X"00",X"55",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"F5",X"00",X"00",
		X"00",X"57",X"00",X"00",X"00",X"57",X"00",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",
		X"00",X"0E",X"EE",X"00",X"00",X"EE",X"EE",X"70",X"00",X"EE",X"0E",X"77",X"00",X"E0",X"07",X"77",
		X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"07",X"77",X"77",X"00",X"77",X"7E",X"70",
		X"00",X"77",X"7E",X"00",X"00",X"77",X"E7",X"E0",X"00",X"77",X"E7",X"EE",X"07",X"77",X"77",X"EE",
		X"77",X"77",X"70",X"EE",X"77",X"77",X"00",X"0E",X"77",X"77",X"00",X"00",X"77",X"37",X"00",X"EE",
		X"77",X"33",X"00",X"00",X"73",X"33",X"00",X"00",X"73",X"33",X"0E",X"00",X"73",X"33",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"40",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",
		X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",
		X"00",X"00",X"00",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",
		X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"40",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",
		X"00",X"04",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"FF",X"00",
		X"00",X"44",X"44",X"00",X"00",X"FF",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"05",
		X"00",X"44",X"44",X"55",X"00",X"44",X"44",X"05",X"00",X"44",X"44",X"00",X"00",X"44",X"45",X"00",
		X"00",X"44",X"55",X"00",X"00",X"44",X"55",X"00",X"00",X"44",X"55",X"00",X"00",X"55",X"55",X"00",
		X"00",X"05",X"55",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",
		X"00",X"06",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"6F",X"66",X"00",X"00",X"6F",X"66",X"00",
		X"00",X"FF",X"66",X"00",X"00",X"FF",X"66",X"00",X"00",X"F6",X"66",X"00",X"00",X"F6",X"66",X"06",
		X"00",X"66",X"66",X"66",X"00",X"66",X"66",X"0D",X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"00",
		X"00",X"66",X"66",X"00",X"00",X"66",X"DD",X"00",X"00",X"66",X"DD",X"00",X"00",X"86",X"DD",X"00",
		X"00",X"06",X"DD",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"C0",X"00",X"CC",X"AA",X"CC",X"00",X"CA",X"AA",X"AC",
		X"00",X"AA",X"CA",X"CC",X"00",X"AA",X"CC",X"C0",X"00",X"AA",X"FC",X"C0",X"00",X"AA",X"CC",X"CC",
		X"00",X"AA",X"CC",X"AC",X"00",X"AA",X"CC",X"AC",X"00",X"AA",X"CC",X"CC",X"00",X"AA",X"CA",X"C0",
		X"00",X"AA",X"CC",X"C0",X"00",X"AA",X"FC",X"CC",X"00",X"AA",X"CC",X"AC",X"00",X"AA",X"CC",X"AC",
		X"00",X"AA",X"CC",X"CC",X"00",X"AA",X"CC",X"C0",X"00",X"AA",X"CA",X"CC",X"00",X"AA",X"AA",X"AC",
		X"00",X"CA",X"AA",X"AC",X"00",X"CC",X"AA",X"CC",X"00",X"00",X"CC",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"C0",X"00",X"CC",X"66",X"CC",X"00",X"C6",X"66",X"6C",
		X"00",X"66",X"C6",X"CC",X"00",X"66",X"CC",X"C0",X"00",X"66",X"FC",X"C0",X"00",X"66",X"CC",X"CC",
		X"00",X"66",X"CC",X"6C",X"00",X"66",X"CC",X"6C",X"00",X"66",X"CC",X"CC",X"00",X"66",X"C6",X"C0",
		X"00",X"66",X"CC",X"C0",X"00",X"66",X"FC",X"CC",X"00",X"66",X"CC",X"6C",X"00",X"66",X"CC",X"6C",
		X"00",X"66",X"CC",X"CC",X"00",X"66",X"CC",X"C0",X"00",X"66",X"C6",X"CC",X"00",X"66",X"66",X"6C",
		X"00",X"C6",X"66",X"6C",X"00",X"CC",X"66",X"CC",X"00",X"00",X"CC",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"C0",X"00",X"CC",X"BB",X"CC",X"00",X"CB",X"BB",X"BC",
		X"00",X"BB",X"CB",X"CC",X"00",X"BB",X"CC",X"C0",X"00",X"BB",X"FC",X"C0",X"00",X"BB",X"CC",X"CC",
		X"00",X"BB",X"CC",X"BC",X"00",X"BB",X"CC",X"BC",X"00",X"BB",X"CC",X"CC",X"00",X"BB",X"CB",X"C0",
		X"00",X"BB",X"CC",X"C0",X"00",X"BB",X"FC",X"CC",X"00",X"BB",X"CC",X"BC",X"00",X"BB",X"CC",X"BC",
		X"00",X"BB",X"CC",X"CC",X"00",X"BB",X"CC",X"C0",X"00",X"BB",X"CB",X"CC",X"00",X"BB",X"BB",X"BC",
		X"00",X"CB",X"BB",X"BC",X"00",X"CC",X"BB",X"CC",X"00",X"00",X"CC",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"0A",X"AA",X"00",X"00",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"00",X"00",X"AA",X"FF",X"00",
		X"00",X"AA",X"AA",X"00",X"00",X"FF",X"AA",X"00",X"00",X"FF",X"AA",X"00",X"00",X"AA",X"AA",X"0A",
		X"00",X"AA",X"AA",X"AA",X"00",X"AA",X"AA",X"0A",X"00",X"AA",X"AA",X"00",X"00",X"AA",X"A9",X"00",
		X"00",X"AA",X"99",X"00",X"00",X"AA",X"99",X"00",X"00",X"9A",X"99",X"00",X"00",X"A9",X"99",X"00",
		X"00",X"0A",X"99",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"7F",X"00",
		X"00",X"00",X"66",X"00",X"00",X"FF",X"66",X"00",X"00",X"00",X"64",X"00",X"00",X"00",X"04",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"05",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"0A",X"00",X"00",X"00",X"A4",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"45",X"00",X"00",X"FF",X"40",X"00",X"00",X"00",X"04",X"00",
		X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"40",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"65",X"00",
		X"00",X"04",X"64",X"00",X"00",X"0A",X"54",X"00",X"00",X"0A",X"04",X"00",X"00",X"00",X"05",X"00",
		X"00",X"05",X"05",X"00",X"00",X"05",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"AA",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"40",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",
		X"00",X"00",X"44",X"44",X"00",X"00",X"04",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",
		X"00",X"00",X"00",X"44",X"00",X"00",X"04",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",
		X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"40",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"00",X"00",X"00",X"44",X"00",X"40",X"00",X"44",X"00",X"40",X"00",X"44",X"00",X"44",
		X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",
		X"00",X"44",X"04",X"44",X"00",X"44",X"04",X"44",X"00",X"44",X"04",X"40",X"00",X"04",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"04",X"00",X"99",X"90",X"00",X"00",X"A9",X"99",X"00",X"00",X"9A",X"99",
		X"0A",X"09",X"9A",X"99",X"00",X"09",X"A9",X"99",X"00",X"09",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"09",X"99",X"99",X"00",X"09",X"A9",X"99",X"00",X"09",X"9A",X"99",X"00",X"00",X"9A",X"99",
		X"00",X"00",X"A9",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",
		X"00",X"04",X"00",X"00",X"00",X"44",X"00",X"40",X"00",X"44",X"00",X"40",X"00",X"44",X"00",X"44",
		X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"04",X"44",X"00",X"44",X"04",X"44",
		X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"40",X"00",X"04",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"60",
		X"00",X"06",X"AA",X"66",X"00",X"06",X"AA",X"A6",X"00",X"06",X"A6",X"A6",X"00",X"06",X"A6",X"A6",
		X"00",X"06",X"A6",X"A6",X"00",X"06",X"A6",X"A6",X"00",X"06",X"A6",X"A6",X"00",X"06",X"A6",X"66",
		X"00",X"00",X"66",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",X"06",X"AA",X"A6",
		X"00",X"06",X"AA",X"A6",X"00",X"06",X"AA",X"A6",X"00",X"06",X"6A",X"A6",X"00",X"06",X"66",X"A6",
		X"00",X"06",X"06",X"A6",X"00",X"00",X"00",X"A6",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"60",
		X"00",X"06",X"AA",X"66",X"00",X"06",X"AA",X"A6",X"00",X"06",X"A6",X"A6",X"00",X"06",X"A6",X"A6",
		X"00",X"06",X"A6",X"A6",X"00",X"06",X"A6",X"A6",X"00",X"06",X"A6",X"A6",X"00",X"06",X"A6",X"66",
		X"00",X"00",X"66",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"60",X"00",X"06",X"AA",X"66",
		X"00",X"06",X"AA",X"A6",X"00",X"06",X"00",X"A6",X"00",X"06",X"00",X"A6",X"00",X"06",X"00",X"A6",
		X"00",X"06",X"00",X"A6",X"00",X"06",X"AA",X"A6",X"00",X"06",X"AA",X"66",X"00",X"00",X"66",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"A6",X"00",X"06",X"66",X"A6",X"00",X"06",X"AA",X"A6",
		X"00",X"06",X"AA",X"A6",X"00",X"06",X"66",X"A6",X"00",X"00",X"00",X"A6",X"00",X"00",X"00",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"60",X"00",X"06",X"AA",X"66",
		X"00",X"06",X"AA",X"A6",X"00",X"06",X"A6",X"A6",X"00",X"06",X"A6",X"A6",X"00",X"06",X"A6",X"A6",
		X"00",X"06",X"A6",X"A6",X"00",X"06",X"A6",X"A6",X"00",X"06",X"A6",X"66",X"00",X"06",X"66",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"A6",X"00",X"06",X"66",X"A6",X"00",X"06",X"AA",X"A6",
		X"00",X"06",X"AA",X"A6",X"00",X"06",X"66",X"A6",X"00",X"00",X"00",X"A6",X"00",X"00",X"00",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",
		X"00",X"06",X"A6",X"A6",X"00",X"06",X"AA",X"A6",X"00",X"06",X"AA",X"A6",X"00",X"06",X"6A",X"A6",
		X"00",X"06",X"66",X"A6",X"00",X"06",X"06",X"A6",X"00",X"06",X"00",X"A6",X"00",X"06",X"00",X"A6",
		X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"A6",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"6A",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"A6",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"60",
		X"00",X"06",X"AA",X"66",X"00",X"06",X"AA",X"A6",X"00",X"06",X"AA",X"A6",X"00",X"06",X"AA",X"A6",
		X"00",X"06",X"AA",X"A6",X"00",X"06",X"AA",X"A6",X"00",X"06",X"66",X"A6",X"00",X"06",X"00",X"66",
		X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"A6",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"6A",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"A6",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"6A",X"00",
		X"00",X"00",X"6A",X"00",X"00",X"66",X"6A",X"66",X"00",X"AA",X"AA",X"A6",X"00",X"6A",X"AA",X"A6",
		X"00",X"66",X"0A",X"66",X"00",X"06",X"0A",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"0A",X"00",
		X"00",X"00",X"0A",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"6A",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"A6",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"6A",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"A6",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"60",
		X"00",X"06",X"AA",X"66",X"00",X"06",X"AA",X"A6",X"00",X"06",X"A6",X"A6",X"00",X"06",X"A6",X"A6",
		X"00",X"06",X"A6",X"A6",X"00",X"06",X"A6",X"A6",X"00",X"06",X"A6",X"A6",X"00",X"06",X"A6",X"66",
		X"00",X"00",X"66",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"A6",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"6A",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"A6",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"C0",X"00",X"CC",X"55",X"CC",X"00",X"C5",X"55",X"5C",
		X"00",X"55",X"C5",X"CC",X"00",X"55",X"CC",X"C0",X"00",X"55",X"FC",X"C0",X"00",X"55",X"CC",X"CC",
		X"00",X"55",X"CC",X"5C",X"00",X"55",X"CC",X"5C",X"00",X"55",X"CC",X"CC",X"00",X"55",X"C5",X"C0",
		X"00",X"55",X"CC",X"C0",X"00",X"55",X"FC",X"CC",X"00",X"55",X"CC",X"5C",X"00",X"55",X"CC",X"5C",
		X"00",X"55",X"CC",X"CC",X"00",X"55",X"CC",X"C0",X"00",X"55",X"C5",X"CC",X"00",X"55",X"55",X"5C",
		X"00",X"C5",X"55",X"5C",X"00",X"CC",X"55",X"CC",X"00",X"00",X"CC",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
