library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity wacko_bg_bits_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of wacko_bg_bits_1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"5A",X"5A",X"A5",X"A5",X"5A",X"5A",X"A5",X"A5",X"5A",X"5A",X"A5",X"A5",X"5A",X"5A",X"A5",X"A5",
		X"A5",X"A5",X"5A",X"5A",X"55",X"55",X"A5",X"A5",X"5A",X"5A",X"55",X"55",X"A5",X"A5",X"5A",X"5A",
		X"55",X"55",X"A5",X"A5",X"5A",X"5A",X"55",X"55",X"A5",X"A5",X"5A",X"5A",X"55",X"55",X"55",X"55",
		X"A5",X"A5",X"5A",X"5A",X"55",X"55",X"55",X"55",X"A5",X"A5",X"5A",X"5A",X"55",X"55",X"55",X"55",
		X"A9",X"A5",X"5A",X"5A",X"55",X"55",X"55",X"55",X"55",X"55",X"A5",X"A5",X"5A",X"5A",X"55",X"55",
		X"55",X"55",X"55",X"55",X"A5",X"A5",X"5A",X"5A",X"55",X"55",X"55",X"55",X"55",X"55",X"A5",X"A5",
		X"5A",X"5A",X"55",X"55",X"55",X"55",X"55",X"55",X"A5",X"A5",X"5A",X"5A",X"55",X"55",X"55",X"55",
		X"55",X"55",X"A5",X"A5",X"5A",X"5A",X"55",X"55",X"55",X"55",X"55",X"55",X"A5",X"A5",X"5A",X"5A",
		X"55",X"55",X"55",X"55",X"55",X"55",X"A5",X"A5",X"5A",X"5A",X"55",X"55",X"55",X"55",X"55",X"55",
		X"A5",X"A5",X"5A",X"5A",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"A5",X"A5",X"5A",X"5A",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"A5",X"A5",X"5A",X"5A",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"A5",X"A5",X"5A",X"5A",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"A5",X"A5",X"5A",X"5A",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"A5",X"A5",X"5A",X"5A",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"A5",X"A5",X"5A",X"5A",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"6A",X"56",X"AB",
		X"5A",X"AF",X"5A",X"AF",X"AA",X"BF",X"AA",X"BF",X"AA",X"BF",X"AA",X"BF",X"AA",X"BF",X"AA",X"AF",
		X"AA",X"AF",X"AA",X"AA",X"AA",X"AE",X"AA",X"BE",X"AA",X"FA",X"AB",X"FA",X"AF",X"EA",X"BF",X"EA",
		X"FF",X"EA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"EA",X"FF",X"EA",
		X"FF",X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F5",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"6B",X"55",X"AB",X"56",X"AF",X"56",X"AF",X"5E",X"AF",X"FE",X"AB",X"FE",X"AB",X"FF",X"AA",
		X"FF",X"AA",X"FF",X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"FF",X"AE",X"FF",X"BE",
		X"FE",X"BE",X"FA",X"BE",X"BA",X"FE",X"AA",X"FE",X"AA",X"FF",X"AA",X"FF",X"AB",X"FF",X"AB",X"FF",
		X"AB",X"FF",X"AB",X"FF",X"AB",X"FF",X"AB",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"BF",X"AA",X"AB",
		X"AA",X"AA",X"AA",X"AA",X"FA",X"AA",X"FF",X"FE",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"A9",X"55",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"55",X"5B",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"F5",X"55",X"FD",X"55",
		X"FD",X"55",X"FD",X"55",X"FF",X"56",X"FF",X"F6",X"FF",X"FA",X"FF",X"EA",X"FF",X"AA",X"FF",X"AA",
		X"BE",X"AB",X"AA",X"AB",X"EA",X"AB",X"EA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"AA",X"FA",X"AA",X"FA",X"AA",
		X"FF",X"EA",X"FF",X"EA",X"FF",X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"BF",X"FF",X"AA",X"BF",X"AA",X"AA",X"AA",X"A5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"57",X"55",X"57",X"55",X"5F",X"55",X"7E",X"55",X"FE",X"57",X"FE",
		X"5F",X"FE",X"7F",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"FF",X"BF",X"FF",X"AF",X"FF",
		X"AF",X"FF",X"AB",X"FF",X"AA",X"FF",X"AA",X"BF",X"FA",X"AF",X"FF",X"EF",X"FF",X"FF",X"FF",X"F5",
		X"FF",X"D5",X"FD",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"A5",X"55",X"55",X"56",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"7E",X"55",X"FA",X"95",X"EA",X"A5",X"EA",X"A9",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"EA",X"AA",X"EA",X"AA",X"FA",X"AA",X"FA",X"AA",X"FE",X"AA",X"FE",X"AA",X"FF",X"AA",
		X"FF",X"EA",X"FF",X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FC",X"FF",X"F4",X"FF",X"D4",X"FF",X"54",X"FD",X"54",X"F5",X"54",X"55",X"54",X"55",X"54",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"6A",X"A9",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"0A",X"A0",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"0A",X"A0",
		X"00",X"00",X"0A",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"0A",X"A0",
		X"00",X"00",X"2A",X"A0",X"20",X"A0",X"00",X"A0",X"2A",X"A0",X"28",X"00",X"28",X"20",X"2A",X"A0",
		X"00",X"00",X"2A",X"A0",X"20",X"A0",X"00",X"A0",X"0A",X"80",X"00",X"A0",X"20",X"A0",X"2A",X"A0",
		X"00",X"00",X"00",X"A0",X"28",X"A0",X"28",X"A0",X"2A",X"A8",X"00",X"A0",X"00",X"A0",X"00",X"A0",
		X"00",X"00",X"2A",X"A0",X"28",X"20",X"28",X"00",X"2A",X"A0",X"00",X"A0",X"20",X"A0",X"2A",X"A0",
		X"00",X"00",X"2A",X"A8",X"28",X"28",X"28",X"00",X"2A",X"A8",X"28",X"28",X"28",X"28",X"2A",X"A8",
		X"00",X"00",X"2A",X"A0",X"28",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",
		X"00",X"00",X"2A",X"A8",X"28",X"28",X"28",X"28",X"0A",X"A0",X"28",X"28",X"28",X"28",X"2A",X"A8",
		X"00",X"00",X"2A",X"A8",X"28",X"28",X"28",X"28",X"2A",X"A8",X"00",X"28",X"28",X"28",X"2A",X"A8",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"A5",X"55",
		X"A9",X"55",X"A9",X"55",X"AA",X"55",X"AA",X"56",X"AA",X"5A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"05",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"AA",X"FE",X"AA",X"FF",X"FA",X"C0",X"FC",X"00",X"00",
		X"01",X"50",X"01",X"50",X"05",X"50",X"15",X"50",X"55",X"50",X"55",X"40",X"55",X"40",X"55",X"00",
		X"00",X"01",X"00",X"01",X"00",X"01",X"40",X"01",X"40",X"00",X"50",X"00",X"54",X"00",X"55",X"00",
		X"55",X"40",X"55",X"55",X"A5",X"5A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"0A",X"A0",X"28",X"28",X"28",X"28",X"28",X"28",X"2A",X"A8",X"28",X"28",X"28",X"28",
		X"00",X"00",X"2A",X"A8",X"28",X"28",X"28",X"28",X"2A",X"A0",X"28",X"28",X"28",X"28",X"2A",X"A8",
		X"00",X"00",X"2A",X"A8",X"28",X"28",X"28",X"00",X"28",X"00",X"28",X"28",X"28",X"28",X"2A",X"A8",
		X"00",X"00",X"2A",X"A0",X"28",X"A8",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"A8",X"2A",X"A0",
		X"00",X"00",X"2A",X"A8",X"28",X"28",X"28",X"00",X"2A",X"80",X"28",X"00",X"28",X"28",X"2A",X"A8",
		X"00",X"00",X"2A",X"A8",X"28",X"28",X"28",X"00",X"2A",X"80",X"28",X"00",X"28",X"00",X"28",X"00",
		X"00",X"00",X"2A",X"A8",X"28",X"28",X"28",X"00",X"28",X"A8",X"28",X"28",X"28",X"28",X"2A",X"A8",
		X"00",X"00",X"28",X"28",X"28",X"28",X"28",X"28",X"2A",X"A8",X"28",X"28",X"28",X"28",X"28",X"28",
		X"00",X"00",X"0A",X"A0",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"0A",X"A0",
		X"00",X"00",X"02",X"A8",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"28",X"A0",X"28",X"A0",X"2A",X"A0",
		X"00",X"00",X"28",X"20",X"28",X"A0",X"2A",X"A0",X"2A",X"00",X"2A",X"A0",X"28",X"A0",X"28",X"A0",
		X"00",X"00",X"28",X"00",X"28",X"00",X"28",X"00",X"28",X"00",X"28",X"28",X"28",X"28",X"2A",X"A8",
		X"00",X"00",X"A8",X"A8",X"AA",X"A8",X"A2",X"28",X"A2",X"28",X"A0",X"28",X"A0",X"28",X"A0",X"28",
		X"00",X"00",X"A0",X"28",X"A8",X"28",X"AA",X"28",X"AA",X"A8",X"A2",X"A8",X"A0",X"A8",X"A0",X"28",
		X"00",X"00",X"2A",X"A8",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"2A",X"A8",
		X"00",X"00",X"2A",X"A8",X"28",X"28",X"28",X"28",X"2A",X"A8",X"28",X"00",X"28",X"00",X"28",X"00",
		X"00",X"00",X"AA",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A2",X"A0",X"A2",X"A8",X"AA",X"A8",
		X"00",X"00",X"2A",X"A8",X"28",X"28",X"28",X"28",X"2A",X"A0",X"28",X"28",X"28",X"28",X"28",X"28",
		X"00",X"00",X"2A",X"A8",X"28",X"28",X"28",X"00",X"2A",X"A8",X"00",X"28",X"28",X"28",X"2A",X"A8",
		X"00",X"00",X"2A",X"A8",X"2A",X"A8",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",
		X"00",X"00",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"2A",X"A8",
		X"00",X"00",X"28",X"08",X"28",X"08",X"28",X"08",X"28",X"28",X"28",X"A0",X"2A",X"80",X"2A",X"00",
		X"00",X"00",X"A0",X"28",X"A0",X"28",X"A0",X"28",X"A2",X"28",X"A2",X"28",X"AA",X"A8",X"A8",X"A8",
		X"00",X"00",X"A0",X"28",X"A8",X"A8",X"2A",X"A0",X"0A",X"80",X"2A",X"A0",X"A8",X"A8",X"A0",X"28",
		X"00",X"00",X"28",X"28",X"28",X"28",X"2A",X"A8",X"0A",X"A0",X"02",X"80",X"02",X"80",X"02",X"80",
		X"00",X"00",X"2A",X"A8",X"28",X"28",X"00",X"A0",X"02",X"80",X"0A",X"00",X"28",X"28",X"2A",X"A8",
		X"55",X"56",X"55",X"5A",X"55",X"6B",X"55",X"AB",X"55",X"AF",X"56",X"AF",X"5A",X"BF",X"5A",X"BF",
		X"6A",X"BF",X"AA",X"BF",X"AA",X"BF",X"AA",X"BF",X"AA",X"AF",X"AA",X"AF",X"AA",X"AB",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A9",X"AA",X"A5",X"AA",X"95",
		X"AA",X"55",X"A9",X"55",X"A1",X"55",X"A1",X"55",X"81",X"55",X"05",X"55",X"05",X"55",X"05",X"55",
		X"05",X"55",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"A5",X"55",X"A9",X"55",X"AA",X"95",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"D5",X"55",X"F5",X"55",X"F5",X"55",X"FD",X"55",X"FD",X"55",X"FD",X"55",X"FD",X"5F",X"FF",X"7F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"A0",X"0F",X"A0",X"03",X"90",X"00",X"50",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"40",X"00",X"50",X"00",
		X"50",X"00",X"50",X"00",X"50",X"00",X"54",X"00",X"54",X"00",X"54",X"00",X"55",X"00",X"55",X"00",
		X"55",X"40",X"55",X"40",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"54",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"A5",X"55",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"D5",X"55",X"F5",X"55",
		X"F5",X"55",X"F5",X"55",X"FD",X"55",X"FF",X"D5",X"FF",X"55",X"FF",X"55",X"FD",X"55",X"FD",X"55",
		X"F5",X"55",X"C5",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"01",X"55",X"01",X"55",X"00",X"55",
		X"00",X"55",X"00",X"15",X"00",X"15",X"00",X"05",X"00",X"05",X"00",X"01",X"00",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"00",X"14",X"00",X"14",X"00",X"54",X"00",X"54",X"00",X"54",X"00",X"54",X"00",X"50",X"00",
		X"54",X"00",X"54",X"00",X"6A",X"00",X"5A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"51",X"55",X"41",X"55",X"41",X"55",
		X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",
		X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"05",X"40",X"05",X"40",X"05",X"40",X"05",X"40",X"05",
		X"40",X"01",X"40",X"01",X"50",X"01",X"50",X"00",X"50",X"00",X"50",X"00",X"54",X"00",X"55",X"00",
		X"55",X"00",X"15",X"40",X"05",X"40",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"AA",X"02",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"55",X"55",X"55",X"51",X"55",X"40",X"55",X"40",X"55",X"00",X"55",X"00",X"54",X"00",X"54",X"00",
		X"54",X"00",X"54",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",
		X"54",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"15",X"40",X"15",X"40",X"05",X"40",
		X"05",X"50",X"01",X"50",X"00",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"05",X"05",
		X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"AA",X"A0",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"56",X"1F",X"5A",X"0F",X"9A",X"0F",X"AA",
		X"03",X"EA",X"00",X"FA",X"00",X"2A",X"00",X"0A",X"00",X"02",X"00",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"A7",X"56",X"BF",X"5A",X"BF",
		X"6A",X"FF",X"6A",X"FF",X"AA",X"FF",X"AA",X"FF",X"AB",X"FF",X"AB",X"FF",X"AB",X"FF",X"AB",X"FF",
		X"AA",X"FF",X"AA",X"FF",X"AA",X"BF",X"AA",X"BF",X"AA",X"BF",X"AA",X"AF",X"AA",X"AF",X"AA",X"AB",
		X"AA",X"AA",X"2A",X"AA",X"2A",X"AA",X"0A",X"AA",X"00",X"AA",X"00",X"2A",X"00",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",X"AA",X"AA",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"F5",X"55",X"FD",X"55",X"FD",X"55",X"FF",X"55",
		X"FF",X"55",X"FF",X"D6",X"FF",X"FA",X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",
		X"FF",X"EA",X"FF",X"FA",X"FF",X"FA",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"BF",X"FF",X"AF",X"FF",X"AB",X"FF",X"AA",X"BF",X"AA",X"AA",X"AA",X"AA",X"02",X"AB",
		X"00",X"AF",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",X"02",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"F5",X"F5",X"F7",X"FD",X"FF",X"FD",X"FF",X"EE",X"FF",X"EA",X"BF",X"EA",X"BF",X"AA",X"AF",X"AA",
		X"AF",X"AA",X"AB",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"AA",X"FE",X"FA",
		X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"0F",X"FF",X"03",X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"55",X"5F",X"55",X"7F",X"55",X"7F",X"55",X"7F",X"55",X"FF",X"55",X"FF",X"56",X"FF",X"AA",X"FF",
		X"AA",X"FF",X"AB",X"FF",X"AB",X"FF",X"AB",X"FF",X"AB",X"FF",X"AB",X"FF",X"AB",X"FF",X"AB",X"FF",
		X"AB",X"FF",X"AB",X"FF",X"AB",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"BF",X"AA",X"AF",
		X"AA",X"BF",X"EA",X"FF",X"EB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"FF",X"00",X"03",
		X"00",X"00",X"00",X"AA",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"54",X"00",X"50",X"00",X"50",X"00",X"A8",X"00",X"A0",X"00",X"A0",X"00",X"A8",X"00",X"AA",X"A8",
		X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"95",X"6A",X"A5",X"EA",X"A5",X"EA",X"AD",X"EA",X"AD",
		X"EA",X"AE",X"EA",X"AE",X"EA",X"AE",X"EA",X"BE",X"AA",X"BF",X"AA",X"BF",X"AA",X"BF",X"AA",X"AF",
		X"AA",X"AF",X"AA",X"AF",X"AA",X"AF",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"EA",X"AA",X"FA",X"AA",
		X"FA",X"AA",X"FA",X"AA",X"FE",X"AA",X"FE",X"AA",X"FF",X"AA",X"FF",X"FA",X"C0",X"3F",X"C0",X"03",
		X"00",X"03",X"00",X"03",X"00",X"00",X"F0",X"00",X"FC",X"00",X"FC",X"00",X"FF",X"00",X"FF",X"00",
		X"3F",X"C0",X"00",X"FC",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"6B",X"55",
		X"AB",X"C0",X"AB",X"E4",X"AB",X"E5",X"AF",X"E5",X"AF",X"E5",X"AF",X"E9",X"AF",X"E9",X"AF",X"EA",
		X"00",X"05",X"00",X"15",X"00",X"15",X"00",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FC",X"BF",X"FC",X"BF",X"FC",X"BF",X"F0",X"AF",X"F0",X"AB",X"F0",X"EF",X"F0",X"FF",X"F0",
		X"FF",X"FC",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"FD",X"00",X"FD",X"00",X"01",
		X"00",X"02",X"00",X"2A",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"55",X"5F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"05",X"40",X"15",X"40",X"55",X"50",X"55",X"50",X"55",X"54",X"55",X"54",X"55",X"54",
		X"AA",X"80",X"AA",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"55",X"40",X"55",X"00",X"55",X"00",X"95",X"00",X"A9",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"05",X"00",X"05",X"00",X"15",X"00",X"54",X"01",X"54",X"05",X"54",X"15",X"50",X"15",X"50",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"02",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"04",X"00",X"00",X"00",X"00",X"0A",X"00",X"AA",X"A0",X"AA",X"A8",X"AA",X"AA",X"AA",X"AA",
		X"A0",X"00",X"A0",X"00",X"A8",X"00",X"AA",X"A8",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"95",X"A9",X"54",X"A9",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"01",X"55",X"01",X"55",
		X"00",X"05",X"00",X"15",X"00",X"55",X"00",X"55",X"15",X"54",X"55",X"50",X"55",X"40",X"55",X"00",
		X"00",X"15",X"00",X"55",X"01",X"55",X"15",X"55",X"55",X"54",X"55",X"50",X"55",X"40",X"55",X"00",
		X"55",X"40",X"54",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C0",X"FF",X"00",X"FC",X"00",X"F0",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"D5",X"55",X"FD",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FE",X"A8",X"FF",X"A0",X"FF",X"C0",
		X"AA",X"80",X"AA",X"00",X"AA",X"00",X"A8",X"00",X"A0",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"F0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"01",X"00",X"01",X"00",X"05",X"00",X"05",X"00",X"14",X"00",X"14",X"00",X"50",X"00",X"50",X"00",
		X"95",X"55",X"A9",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"95",X"AA",X"A9",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",X"FF",X"AA",
		X"FE",X"AA",X"FA",X"AA",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"AF",X"FF",X"AA",X"FF",X"AA",X"AA",X"EA",X"AA",X"FA",X"AA",X"FA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FF",X"FC",X"FF",X"F0",X"FF",X"C0",
		X"A5",X"55",X"A9",X"55",X"A9",X"55",X"AA",X"57",X"AA",X"5F",X"AA",X"7F",X"AA",X"FF",X"AA",X"BF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"AA",X"FA",X"AA",
		X"FA",X"AA",X"FF",X"AA",X"FF",X"FA",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"7D",X"55",X"FE",X"57",X"FA",X"5F",X"FA",X"5F",X"FA",X"5F",X"FA",X"7F",X"FA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"FF",X"0F",X"FF",X"03",X"FF",
		X"03",X"FF",X"03",X"FF",X"03",X"FF",X"03",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",X"FF",X"03",X"FF",
		X"0F",X"FF",X"03",X"FF",X"00",X"FF",X"00",X"3F",X"00",X"3F",X"00",X"0F",X"00",X"0F",X"00",X"0F",
		X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",X"00",X"03",X"40",X"00",X"50",X"00",X"50",X"00",
		X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"40",X"55",X"40",X"55",X"00",
		X"55",X"00",X"94",X"00",X"A4",X"00",X"A0",X"00",X"A0",X"00",X"A8",X"20",X"AA",X"AA",X"AA",X"AA",
		X"55",X"57",X"95",X"FF",X"BF",X"FF",X"BF",X"FF",X"AF",X"FF",X"AA",X"FF",X"AA",X"BF",X"AA",X"AF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"51",X"01",X"55",X"41",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"F5",X"55",X"E5",X"55",X"A9",X"55",X"A9",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"95",X"AA",X"95",
		X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"A8",X"FA",X"A0",X"FF",X"A0",X"FF",X"C0",X"FF",X"00",X"FC",X"00",X"F0",X"00",
		X"00",X"55",X"00",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"15",X"55",X"15",X"55",X"15",X"55",
		X"FA",X"A5",X"FA",X"9A",X"FA",X"A5",X"FA",X"AA",X"FA",X"A5",X"FA",X"AA",X"FA",X"A9",X"FA",X"AA",
		X"FA",X"A9",X"FA",X"AA",X"FA",X"AA",X"FE",X"AA",X"FE",X"AA",X"FE",X"AA",X"FE",X"AA",X"FE",X"AA",
		X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"EA",X"FF",X"EA",X"FF",X"FA",X"FF",X"FA",
		X"55",X"55",X"55",X"6A",X"56",X"AA",X"2A",X"AA",X"0A",X"AA",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"A5",X"A5",X"AA",X"5A",X"AA",X"A5",X"AA",X"BA",X"AA",X"B5",X"AA",X"BE",X"AA",X"FD",X"AA",X"FE",
		X"AA",X"FD",X"AA",X"FE",X"AB",X"FA",X"AB",X"FA",X"AF",X"FA",X"AF",X"FA",X"AF",X"FA",X"AF",X"FA",
		X"AF",X"FA",X"AF",X"FA",X"EF",X"FA",X"FF",X"FE",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"A5",X"A5",X"5A",X"5A",X"A6",X"A5",X"AA",X"5B",X"A9",X"AF",X"AA",X"7F",X"AA",X"FE",X"AB",X"FE",
		X"AB",X"FE",X"AB",X"FE",X"AB",X"FE",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"EA",X"BF",X"FA",X"BF",
		X"A5",X"A5",X"5A",X"5A",X"EA",X"A5",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"AA",X"EA",X"AA",X"FF",X"AA",X"FF",X"FF",
		X"A5",X"A5",X"5A",X"5A",X"A5",X"A5",X"5A",X"5A",X"A5",X"A5",X"AA",X"5A",X"A5",X"A5",X"AA",X"5A",
		X"AA",X"A5",X"AA",X"DA",X"AA",X"A5",X"AA",X"5A",X"AA",X"A5",X"AA",X"5A",X"FD",X"A5",X"FE",X"5A",
		X"FF",X"E5",X"FF",X"FA",X"FF",X"FD",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"A5",X"A5",X"5A",X"AA",X"A5",X"AA",X"5A",X"AA",X"AA",X"AA",X"5A",X"AA",X"AA",X"AA",X"5A",X"AA",
		X"BA",X"AA",X"FE",X"AA",X"FE",X"AA",X"FE",X"AA",X"FF",X"AA",X"FF",X"AA",X"7F",X"AA",X"BF",X"EA",
		X"3F",X"FA",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",X"AF",X"FF",X"AB",X"FF",X"AB",X"FF",
		X"AA",X"FF",X"AA",X"BF",X"AA",X"AF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"A5",X"A5",X"5A",X"5A",X"A5",X"AA",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"57",X"AA",X"5F",X"AA",X"7F",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"EA",X"FF",X"FA",X"FF",X"FA",
		X"A5",X"A5",X"5A",X"5A",X"A5",X"A5",X"5A",X"5A",X"A5",X"A5",X"5A",X"5A",X"AA",X"AA",X"6A",X"AA",
		X"FA",X"AA",X"EA",X"AA",X"FA",X"AA",X"FE",X"AA",X"FF",X"EA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"A5",X"A5",X"5A",X"5A",X"A5",X"A7",X"5A",X"5B",X"A5",X"AF",X"5A",X"5F",X"A5",X"AF",X"5A",X"9F",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"AA",X"FA",X"AA",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"AA",X"FF",X"AA",X"FF",X"EA",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"5F",X"55",X"5F",X"55",X"57",X"F5",X"55",X"D5",X"57",X"F5",X"5F",X"F6",X"57",X"59",X"57",X"E9",
		X"AA",X"AF",X"AA",X"AF",X"AA",X"AF",X"AA",X"AB",X"AA",X"AA",X"EA",X"AA",X"EA",X"AA",X"FA",X"AA",
		X"A5",X"A7",X"5A",X"5F",X"A5",X"AF",X"5A",X"5F",X"A5",X"BF",X"5A",X"7F",X"A5",X"FF",X"5A",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A9",X"AA",X"95",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A5",X"AA",X"5A",X"A5",X"A5",X"5A",X"5A",X"A5",X"A5",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"0A",X"A0",X"28",X"28",X"22",X"88",X"22",X"08",X"22",X"08",X"22",X"88",X"28",X"28",X"0A",X"A0",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",X"FC",
		X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",X"FF",
		X"00",X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"F0",
		X"FF",X"F0",X"FF",X"F0",X"03",X"F0",X"03",X"F0",X"03",X"F0",X"03",X"F0",X"03",X"F0",X"03",X"F0",
		X"03",X"F0",X"03",X"F0",X"03",X"F0",X"03",X"F0",X"03",X"F0",X"03",X"F0",X"03",X"F0",X"03",X"F0",
		X"03",X"F0",X"03",X"F0",X"03",X"FF",X"03",X"FF",X"03",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",
		X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"AA",X"80",X"AA",X"00",X"AC",X"00",X"FC",X"00",X"FC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"03",X"C0",X"03",X"C0",X"0F",X"C0",X"0F",
		X"C0",X"3F",X"C0",X"3F",X"C0",X"FF",X"C0",X"FC",X"C3",X"FC",X"C3",X"F0",X"CF",X"F0",X"CF",X"C0",
		X"FF",X"C0",X"FF",X"00",X"FF",X"00",X"FC",X"00",X"FC",X"00",X"F0",X"00",X"F0",X"00",X"C0",X"00",
		X"FC",X"00",X"FC",X"00",X"FC",X"00",X"3C",X"00",X"3C",X"00",X"3C",X"00",X"FC",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"03",X"00",X"03",X"00",X"0F",X"00",X"0F",X"00",X"3F",X"00",X"3F",X"00",X"FF",
		X"00",X"FF",X"03",X"FC",X"03",X"FC",X"0F",X"F0",X"0F",X"F0",X"3F",X"C0",X"3F",X"C0",X"FF",X"00",
		X"FF",X"00",X"FC",X"00",X"FC",X"00",X"F0",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"30",X"00",X"FC",X"00",X"FC",X"03",X"FC",X"03",X"FC",X"0F",X"FC",X"0F",X"FC",
		X"3F",X"FC",X"3F",X"3F",X"FF",X"3F",X"FC",X"3F",X"FC",X"3F",X"F0",X"3F",X"F0",X"3F",X"C0",X"3F",
		X"0C",X"00",X"0C",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"C0",X"0A",X"C0",X"0A",X"AA",X"02",X"AA",
		X"00",X"0F",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"00",X"C0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",
		X"F0",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",X"3C",X"00",X"3F",X"00",
		X"3F",X"00",X"3F",X"00",X"3F",X"C0",X"3F",X"FF",X"0F",X"FF",X"0F",X"FF",X"00",X"00",X"00",X"00",
		X"A9",X"55",X"AA",X"55",X"AA",X"95",X"AA",X"A5",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",
		X"C0",X"03",X"C0",X"03",X"C0",X"0F",X"F0",X"0F",X"F0",X"3F",X"F0",X"3F",X"F0",X"FF",X"F0",X"FF",
		X"F3",X"FC",X"F3",X"FC",X"F3",X"F0",X"FF",X"F0",X"FF",X"C0",X"FF",X"C0",X"FF",X"00",X"FF",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FA",X"AA",X"00",X"0A",X"00",X"0F",X"00",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",X"00",X"0F",
		X"00",X"0F",X"00",X"3F",X"00",X"3F",X"00",X"FF",X"00",X"FC",X"03",X"FC",X"03",X"F0",X"0F",X"F0",
		X"0F",X"C0",X"3F",X"C0",X"3F",X"00",X"FF",X"00",X"FC",X"00",X"F0",X"00",X"00",X"03",X"00",X"03",
		X"00",X"FF",X"03",X"FF",X"0F",X"FF",X"0F",X"FF",X"3F",X"C0",X"3F",X"C0",X"FF",X"00",X"FF",X"00",
		X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"FA",X"AA",X"FA",X"AA",X"FA",X"AA",X"FE",X"AA",X"FE",X"AA",
		X"0F",X"C0",X"3F",X"C0",X"3F",X"C0",X"FF",X"00",X"FC",X"00",X"FC",X"00",X"F0",X"03",X"F0",X"03",
		X"FF",X"AA",X"FF",X"EA",X"FF",X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"FF",X"00",
		X"FC",X"00",X"F0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"AA",X"FF",X"EA",X"3F",X"FA",X"0F",X"FE",X"00",X"FF",X"00",X"3F",X"00",X"0F",X"00",X"03",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5A",X"55",X"6A",X"97",
		X"03",X"C0",X"0F",X"F0",X"0F",X"F0",X"03",X"C0",X"3F",X"FC",X"03",X"C0",X"0C",X"30",X"3C",X"3C",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"BF",X"AA",X"BF",X"AA",X"FF",
		X"AA",X"BF",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"BF",
		X"AA",X"BF",X"AA",X"BF",X"EA",X"AF",X"FA",X"AB",X"FF",X"EA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FA",X"0F",X"FA",X"3F",X"EA",X"3F",X"EA",X"FF",X"AA",X"FF",X"AA",X"FE",X"AA",X"FE",X"AA",
		X"AA",X"AA",X"AA",X"AB",X"AA",X"AF",X"AA",X"AF",X"AA",X"BF",X"AA",X"BC",X"AA",X"FC",X"AA",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"AA",X"EA",X"AB",X"EA",X"AB",X"EA",X"AF",X"EA",X"AF",X"EA",X"BF",X"EA",X"BF",X"EA",X"FF",X"EA",
		X"FF",X"EA",X"FF",X"EA",X"F3",X"EA",X"C3",X"EA",X"03",X"EA",X"03",X"EA",X"03",X"EA",X"03",X"EA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",
		X"FF",X"00",X"FF",X"00",X"3F",X"00",X"3C",X"00",X"3C",X"00",X"3C",X"00",X"30",X"00",X"00",X"00",
		X"00",X"03",X"00",X"0F",X"00",X"3F",X"00",X"FF",X"00",X"FC",X"00",X"FC",X"0F",X"F0",X"0A",X"A0",
		X"FF",X"FF",X"FF",X"FE",X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",X"AF",X"FA",X"AF",X"FA",X"AF",X"FA",
		X"AB",X"FF",X"AB",X"FF",X"AB",X"FF",X"AB",X"FF",X"AA",X"FF",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"BF",X"AA",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"F0",X"0F",X"F0",X"0F",X"C0",X"0F",X"C0",X"3F",X"C0",X"3F",X"00",X"3F",X"00",X"3F",X"00",
		X"57",X"D5",X"57",X"55",X"57",X"55",X"5F",X"D5",X"5D",X"D5",X"55",X"D5",X"57",X"E5",X"57",X"55",
		X"3F",X"00",X"3F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"C0",X"0F",X"C0",X"0F",X"C0",
		X"0F",X"C0",X"03",X"F0",X"03",X"F0",X"03",X"FC",X"00",X"FC",X"00",X"FF",X"00",X"3F",X"00",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"F0",X"00",
		X"00",X"03",X"00",X"3F",X"03",X"FF",X"0F",X"FF",X"3F",X"FC",X"FF",X"C0",X"FF",X"00",X"FC",X"00",
		X"FF",X"C0",X"FC",X"00",X"F0",X"00",X"F0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FA",X"FF",X"EA",
		X"C0",X"00",X"F0",X"00",X"FC",X"00",X"FF",X"00",X"3F",X"C0",X"0F",X"F0",X"03",X"FF",X"00",X"FF",
		X"FF",X"EA",X"FF",X"EA",X"AF",X"EA",X"AF",X"EA",X"BF",X"FA",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"FF",X"03",X"FF",X"00",X"FF",X"00",X"3F",X"00",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"00",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AB",X"FF",X"AA",X"FF",X"AA",X"BF",X"AA",X"BF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"FF",X"03",X"FF",
		X"3F",X"C0",X"0F",X"C0",X"0F",X"C0",X"0F",X"F0",X"03",X"FF",X"00",X"FF",X"00",X"3F",X"00",X"03",
		X"AA",X"AF",X"AA",X"AB",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"0F",X"00",X"3F",
		X"AA",X"AB",X"AA",X"AF",X"AA",X"BF",X"AA",X"FF",X"3F",X"FF",X"3F",X"FF",X"0F",X"FF",X"03",X"FF",
		X"AA",X"AF",X"AA",X"AF",X"AA",X"AB",X"AA",X"AB",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"C0",X"00",X"C0",X"00",X"F0",X"00",X"F0",X"00",X"FC",X"00",X"FC",X"00",X"3F",X"00",X"3F",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"00",X"FC",X"03",X"FF",
		X"01",X"55",X"00",X"55",X"00",X"16",X"00",X"0A",X"00",X"02",X"00",X"02",X"00",X"00",X"00",X"00",
		X"C3",X"FF",X"F3",X"CF",X"FF",X"03",X"FF",X"00",X"3C",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"5A",X"55",X"5A",X"55",X"6A",X"5A",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",X"C0",X"0F",X"F0",X"0F",X"FC",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"0F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FC",X"3F",X"FC",X"0F",X"F0",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"03",X"F0",X"03",X"FC",X"0F",X"FF",X"3F",X"FF",X"FF",X"3F",X"FC",X"0F",X"F0",X"03",X"C0",X"00",
		X"01",X"00",X"01",X"00",X"00",X"40",X"00",X"40",X"00",X"40",X"40",X"40",X"50",X"10",X"15",X"50",
		X"05",X"54",X"05",X"41",X"01",X"41",X"01",X"41",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"00",
		X"00",X"3F",X"00",X"FF",X"00",X"FF",X"03",X"FF",X"03",X"FF",X"0F",X"FF",X"0F",X"FF",X"3F",X"3F",
		X"FF",X"3F",X"FC",X"3F",X"FC",X"3F",X"F0",X"3F",X"F0",X"3F",X"C0",X"3F",X"00",X"3F",X"00",X"3F",
		X"3F",X"FF",X"FF",X"3F",X"FC",X"3F",X"FC",X"3F",X"30",X"3F",X"00",X"3F",X"00",X"3F",X"00",X"3F",
		X"3F",X"3F",X"3F",X"FF",X"0F",X"FF",X"03",X"FF",X"03",X"FF",X"03",X"FF",X"0F",X"FF",X"0F",X"FF",
		X"FC",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",
		X"FC",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"03",X"FC",X"0F",X"FC",X"3F",
		X"FC",X"3F",X"FC",X"FF",X"FC",X"FE",X"FF",X"FA",X"FF",X"FA",X"FF",X"EA",X"FF",X"AA",X"FE",X"AA",
		X"AA",X"AA",X"EA",X"AA",X"FA",X"AA",X"FA",X"AA",X"FE",X"AA",X"FF",X"AA",X"FF",X"EA",X"FF",X"FA",
		X"FC",X"FA",X"FC",X"FE",X"FC",X"FF",X"FC",X"3F",X"FC",X"0F",X"FC",X"03",X"FC",X"00",X"FC",X"00",
		X"01",X"00",X"01",X"00",X"05",X"00",X"05",X"40",X"05",X"40",X"05",X"40",X"05",X"40",X"05",X"50",
		X"05",X"50",X"05",X"14",X"04",X"15",X"04",X"15",X"04",X"15",X"04",X"14",X"04",X"14",X"04",X"14",
		X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"05",X"04",X"01",X"04",X"01",X"05",X"01",
		X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"40",X"05",X"40",X"05",X"40",X"05",X"40",
		X"05",X"40",X"05",X"40",X"05",X"50",X"05",X"50",X"05",X"50",X"05",X"50",X"05",X"50",X"05",X"50",
		X"F0",X"00",X"FC",X"00",X"FF",X"00",X"BF",X"C0",X"AF",X"F0",X"AB",X"FC",X"AA",X"FC",X"AA",X"BF",
		X"85",X"55",X"A5",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"F0",X"00",X"C0",X"03",X"00",X"03",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"3F",X"00",X"3F",
		X"00",X"3F",X"00",X"3C",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",X"FC",
		X"C0",X"FC",X"F0",X"FC",X"F0",X"F0",X"FC",X"F0",X"FC",X"F0",X"BF",X"F0",X"AF",X"F0",X"AB",X"F0",
		X"AB",X"FC",X"AA",X"FF",X"AA",X"BF",X"AA",X"AF",X"AA",X"AF",X"AA",X"AB",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"AA",X"FA",X"AA",X"FA",X"AB",
		X"FE",X"AF",X"FF",X"BF",X"3F",X"FF",X"0F",X"FC",X"03",X"F0",X"00",X"F0",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"FF",X"00",X"3F",X"00",X"0F",X"00",X"03",
		X"FC",X"00",X"FC",X"00",X"F0",X"00",X"F0",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"F0",X"00",X"F0",X"00",X"FC",X"00",X"BF",X"00",
		X"AF",X"C0",X"AB",X"F0",X"AB",X"FC",X"AF",X"F0",X"BF",X"C0",X"FF",X"C0",X"FF",X"F0",X"F0",X"FC",
		X"C0",X"3F",X"C0",X"3F",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"FF",X"0F",X"FF",X"FF",X"F0",X"FF",X"00",
		X"00",X"05",X"15",X"55",X"55",X"55",X"55",X"00",X"54",X"00",X"10",X"00",X"10",X"00",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"FF",X"00",X"FF",X"03",X"FC",X"03",X"F0",X"0F",X"C0",
		X"0F",X"00",X"3F",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",
		X"10",X"00",X"14",X"00",X"14",X"00",X"04",X"00",X"05",X"00",X"01",X"00",X"01",X"40",X"01",X"54",
		X"05",X"55",X"05",X"55",X"15",X"54",X"55",X"50",X"05",X"40",X"01",X"40",X"01",X"40",X"01",X"40",
		X"00",X"03",X"00",X"3F",X"00",X"FF",X"FF",X"FF",X"FF",X"F0",X"FF",X"00",X"C0",X"00",X"00",X"00",
		X"00",X"3F",X"00",X"FF",X"00",X"FC",X"03",X"FC",X"0F",X"F0",X"0F",X"F0",X"3F",X"C0",X"3F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"03",X"FF",X"FF",
		X"01",X"40",X"01",X"40",X"01",X"40",X"00",X"50",X"00",X"50",X"00",X"54",X"00",X"14",X"40",X"14",
		X"50",X"04",X"50",X"05",X"50",X"01",X"54",X"01",X"55",X"01",X"15",X"41",X"15",X"45",X"15",X"55",
		X"05",X"00",X"05",X"00",X"01",X"00",X"01",X"40",X"01",X"50",X"00",X"50",X"00",X"54",X"00",X"54",
		X"00",X"15",X"00",X"15",X"40",X"15",X"50",X"05",X"54",X"01",X"95",X"00",X"A5",X"50",X"A5",X"50",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"FF",X"03",X"FF",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"54",X"3F",X"50",X"3F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"07",X"00",X"05",
		X"00",X"05",X"00",X"05",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"40",X"14",
		X"55",X"54",X"15",X"50",X"04",X"14",X"00",X"05",X"00",X"05",X"00",X"01",X"00",X"01",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"50",X"00",X"50",X"00",X"54",X"00",
		X"05",X"00",X"05",X"40",X"01",X"50",X"00",X"54",X"00",X"54",X"00",X"15",X"00",X"15",X"00",X"05",
		X"00",X"05",X"00",X"05",X"40",X"00",X"50",X"00",X"54",X"00",X"58",X"00",X"1A",X"82",X"16",X"AA",
		X"FF",X"FF",X"0C",X"FF",X"04",X"3F",X"05",X"03",X"01",X"40",X"00",X"50",X"00",X"14",X"00",X"04",
		X"00",X"05",X"00",X"01",X"00",X"01",X"00",X"01",X"40",X"05",X"40",X"05",X"50",X"15",X"54",X"15",
		X"14",X"00",X"14",X"00",X"14",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"40",X"05",X"40",
		X"01",X"50",X"01",X"55",X"01",X"55",X"00",X"55",X"00",X"55",X"00",X"15",X"00",X"15",X"00",X"05",
		X"50",X"01",X"54",X"0A",X"A8",X"2A",X"0A",X"AA",X"0A",X"AA",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"FF",X"0F",X"FF",X"03",X"FF",
		X"03",X"FC",X"03",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"50",X"01",X"55",X"00",X"54",X"00",X"14",X"00",X"14",X"00",X"14",X"00",X"05",X"00",X"05",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"AA",X"FE",X"AA",X"FF",X"EA",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FF",X"F0",X"FF",X"C0",X"FC",X"00",
		X"14",X"00",X"05",X"00",X"01",X"00",X"01",X"00",X"05",X"40",X"05",X"50",X"14",X"50",X"10",X"10",
		X"10",X"10",X"54",X"14",X"05",X"55",X"01",X"45",X"05",X"01",X"14",X"00",X"10",X"00",X"50",X"00",
		X"50",X"00",X"54",X"00",X"05",X"00",X"05",X"50",X"01",X"54",X"00",X"15",X"00",X"06",X"00",X"0A",
		X"55",X"55",X"55",X"55",X"55",X"55",X"A5",X"55",X"A5",X"55",X"AA",X"55",X"AA",X"95",X"AA",X"A5",
		X"FF",X"FF",X"FF",X"FF",X"FC",X"3F",X"C0",X"0F",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"45",X"40",X"55",X"40",X"05",X"40",X"05",X"40",X"01",X"50",
		X"00",X"50",X"00",X"50",X"00",X"15",X"00",X"05",X"00",X"00",X"00",X"00",X"A8",X"00",X"AA",X"80",
		X"55",X"5F",X"55",X"7F",X"55",X"FF",X"57",X"FF",X"5F",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"AA",X"00",X"A8",X"00",X"A0",X"00",X"80",X"00",X"00",X"00",
		X"FC",X"00",X"F0",X"00",X"F0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"F0",X"00",X"F0",X"00",
		X"F0",X"00",X"F0",X"00",X"FC",X"00",X"FC",X"00",X"3C",X"00",X"3C",X"00",X"3C",X"00",X"3F",X"00",
		X"0F",X"00",X"0F",X"00",X"0C",X"00",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"05",X"00",X"54",X"00",X"04",X"00",X"05",X"00",X"01",X"54",X"01",X"55",X"15",X"50",
		X"FF",X"C0",X"03",X"F0",X"00",X"3C",X"00",X"0C",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"55",X"00",X"15",X"00",X"05",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"50",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"0F",X"00",X"03",X"00",X"00",
		X"00",X"0F",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",X"00",X"0F",
		X"00",X"0F",X"00",X"3C",X"00",X"F0",X"03",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",
		X"3C",X"00",X"3C",X"00",X"3C",X"00",X"FC",X"00",X"FC",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"C0",
		X"FF",X"0F",X"FC",X"03",X"FC",X"03",X"F0",X"03",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"C0",X"00",
		X"00",X"0F",X"00",X"3F",X"00",X"3F",X"00",X"FF",X"00",X"FF",X"0F",X"FC",X"3F",X"F0",X"FF",X"00",
		X"FF",X"00",X"F0",X"00",X"C0",X"00",X"00",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FF",X"FC",X"FF",X"F0",X"FF",X"F0",X"FF",X"F0",X"FF",X"C0",
		X"FF",X"F0",X"FF",X"F0",X"FF",X"F0",X"FF",X"F0",X"03",X"F0",X"00",X"F0",X"00",X"FC",X"00",X"3C",
		X"00",X"00",X"00",X"02",X"00",X"0A",X"00",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"7A",X"95",X"EA",X"A5",X"E5",X"65",X"E5",X"65",X"E5",X"65",X"F5",X"D5",X"76",X"D5",X"55",X"D5",
		X"3F",X"00",X"0F",X"00",X"2A",X"00",X"AA",X"00",X"A8",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"03",X"FF",X"00",X"FF",X"00",X"3F",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"F0",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",X"FF",X"00",X"3F",X"00",
		X"3F",X"C0",X"0F",X"F0",X"00",X"FF",X"00",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"FE",X"AA",X"FC",X"2A",X"F0",X"02",X"C0",X"02",
		X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"0F",X"80",X"0E",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",
		X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"B0",X"00",X"AA",X"A0",X"AA",X"A8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"0F",X"00",X"3F",
		X"00",X"FF",X"00",X"FE",X"00",X"FD",X"00",X"75",X"01",X"55",X"01",X"55",X"01",X"55",X"01",X"55",
		X"01",X"55",X"01",X"55",X"01",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",
		X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"01",X"56",X"01",X"5A",X"01",X"6A",
		X"02",X"AA",X"00",X"AA",X"00",X"2A",X"00",X"2A",X"00",X"0A",X"00",X"02",X"00",X"00",X"00",X"00",
		X"03",X"F0",X"0F",X"FC",X"3F",X"F8",X"2F",X"FB",X"EF",X"FA",X"EF",X"F6",X"EF",X"F6",X"AF",X"D7",
		X"A7",X"D7",X"A7",X"D7",X"A5",X"D5",X"95",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"5A",X"55",X"AA",X"5A",X"AA",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"03",X"C0",X"0F",X"F0",X"0F",X"F0",X"3F",X"F0",X"AF",X"FC",X"AF",
		X"FF",X"AF",X"F5",X"9F",X"F5",X"5F",X"F5",X"5F",X"D5",X"5D",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"56",X"AA",
		X"00",X"00",X"C0",X"03",X"F0",X"0F",X"FC",X"3F",X"F8",X"FF",X"EA",X"FF",X"EA",X"BF",X"EA",X"BF",
		X"EA",X"5F",X"E9",X"5F",X"69",X"5F",X"59",X"57",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"A5",X"5A",X"A8",X"0A",X"A0",X"4A",X"56",X"95",X"5A",X"A5",X"AA",X"AA",X"AA",X"AA",
		X"55",X"56",X"55",X"5A",X"55",X"6A",X"55",X"AA",X"56",X"AA",X"5A",X"AA",X"6A",X"AA",X"6A",X"AA",
		X"55",X"56",X"55",X"59",X"55",X"6A",X"55",X"A5",X"56",X"5A",X"59",X"A5",X"6A",X"5A",X"A5",X"A5",
		X"0F",X"F0",X"3A",X"E8",X"E5",X"96",X"FA",X"EB",X"FF",X"FF",X"F7",X"FF",X"35",X"7C",X"0F",X"F0",
		X"03",X"C0",X"0F",X"B0",X"0F",X"B0",X"0F",X"F0",X"3F",X"FC",X"2A",X"A8",X"FF",X"FF",X"37",X"1C",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"5A",X"A9",X"6A",X"6A",X"A9",X"AA",X"AA",X"AA",X"AA",X"A5",X"6A",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"59",X"55",X"DF",X"55",X"77",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"7F",X"FD",X"FD",X"7F",X"DD",X"D5",X"75",X"5F",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"D7",X"FA",X"FD",X"55",X"97",X"D5",X"D5",X"FD",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"D6",X"95",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"AA",X"56",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"56",X"AA",X"55",X"55",X"55",X"55",
		X"A5",X"55",X"A5",X"55",X"A5",X"55",X"A5",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"4A",X"55",X"02",X"55",X"00",X"54",X"00",X"54",X"00",X"54",X"00",X"50",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"69",X"55",X"AA",X"55",X"AA",X"95",X"AA",X"AF",X"0A",X"BF",X"00",X"FF",X"00",X"0F",
		X"55",X"55",X"55",X"55",X"55",X"50",X"55",X"59",X"55",X"64",X"55",X"59",X"55",X"04",X"55",X"99",
		X"54",X"41",X"56",X"59",X"59",X"04",X"59",X"65",X"44",X"11",X"66",X"65",X"11",X"04",X"55",X"55",
		X"55",X"55",X"55",X"56",X"7F",X"5A",X"FF",X"EA",X"FF",X"F8",X"F5",X"FC",X"D5",X"F0",X"D5",X"C0",
		X"05",X"55",X"95",X"55",X"45",X"55",X"99",X"55",X"49",X"55",X"99",X"55",X"44",X"55",X"99",X"55",
		X"04",X"15",X"99",X"95",X"44",X"65",X"96",X"55",X"10",X"41",X"65",X"95",X"11",X"04",X"55",X"55",
		X"55",X"55",X"57",X"FF",X"5F",X"FF",X"7F",X"7F",X"FF",X"5F",X"FF",X"57",X"FF",X"57",X"FB",X"FD",
		X"FA",X"FD",X"FA",X"FF",X"FA",X"DD",X"FE",X"D5",X"7F",X"DD",X"55",X"FF",X"55",X"7F",X"55",X"55",
		X"55",X"55",X"5A",X"95",X"EA",X"AF",X"DA",X"AB",X"5A",X"AA",X"59",X"A9",X"F9",X"65",X"79",X"65",
		X"7A",X"5A",X"FE",X"5A",X"DE",X"AA",X"5D",X"9A",X"DD",X"56",X"FD",X"9A",X"FA",X"AB",X"56",X"A5",
		X"55",X"55",X"55",X"55",X"F5",X"55",X"FD",X"55",X"FD",X"55",X"F5",X"D5",X"F5",X"D5",X"75",X"D5",
		X"7F",X"D5",X"75",X"D5",X"F5",X"F5",X"FF",X"75",X"F5",X"75",X"B5",X"F5",X"F7",X"D5",X"FF",X"55",
		X"FF",X"FF",X"CF",X"FF",X"8F",X"FF",X"8F",X"FE",X"83",X"FE",X"A3",X"FF",X"53",X"FF",X"53",X"FF",
		X"60",X"FF",X"64",X"FF",X"64",X"FF",X"54",X"FF",X"50",X"FF",X"53",X"FF",X"53",X"FF",X"53",X"FD",
		X"53",X"FD",X"53",X"FD",X"43",X"FD",X"4F",X"FD",X"4F",X"FD",X"43",X"F5",X"53",X"F5",X"53",X"F5",
		X"53",X"F5",X"53",X"F5",X"50",X"F5",X"54",X"D5",X"54",X"D5",X"54",X"D5",X"57",X"55",X"57",X"55",
		X"FF",X"FF",X"8F",X"FF",X"83",X"FF",X"A3",X"FF",X"A3",X"FF",X"A0",X"FF",X"64",X"FF",X"64",X"FE",
		X"94",X"FE",X"54",X"FE",X"50",X"FE",X"53",X"FE",X"53",X"FD",X"53",X"FD",X"50",X"FD",X"54",X"FD",
		X"54",X"FD",X"54",X"F5",X"54",X"F5",X"50",X"F5",X"53",X"F5",X"53",X"F5",X"53",X"F5",X"53",X"F5",
		X"54",X"F5",X"54",X"F5",X"54",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"0F",X"FF",X"83",X"FE",X"A3",X"FE",X"A3",X"FD",
		X"A0",X"FD",X"58",X"FD",X"58",X"FD",X"54",X"F5",X"54",X"F5",X"53",X"F5",X"53",X"F5",X"53",X"F5",
		X"53",X"F5",X"53",X"F5",X"53",X"D5",X"57",X"D5",X"57",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"3F",X"FF",X"0F",X"FF",X"8F",X"FE",X"83",X"FE",X"A3",X"F6",X"A0",X"FA",X"A8",X"F6",
		X"A8",X"D6",X"64",X"D5",X"67",X"D5",X"97",X"55",X"57",X"55",X"57",X"55",X"55",X"55",X"55",X"55",
		X"55",X"50",X"55",X"00",X"54",X"00",X"50",X"00",X"50",X"00",X"40",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
