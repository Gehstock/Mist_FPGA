library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity spr_rom1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of spr_rom1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"20",X"42",X"26",X"6A",X"7E",X"F8",X"44",X"55",
		X"40",X"24",X"46",X"65",X"6F",X"F1",X"E6",X"66",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"08",
		X"02",X"02",X"02",X"11",X"00",X"00",X"00",X"00",X"A8",X"64",X"34",X"22",X"BA",X"42",X"40",X"00",
		X"77",X"66",X"C6",X"44",X"D5",X"24",X"20",X"00",X"04",X"04",X"04",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"31",X"14",X"04",X"4C",X"08",X"FB",X"9A",X"66",X"11",
		X"88",X"8C",X"42",X"C6",X"ED",X"F3",X"37",X"FD",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"8C",
		X"02",X"22",X"02",X"11",X"00",X"00",X"00",X"00",X"35",X"64",X"FE",X"10",X"BC",X"70",X"20",X"00",
		X"FD",X"46",X"E6",X"33",X"F0",X"80",X"00",X"00",X"CC",X"CC",X"C8",X"88",X"00",X"00",X"00",X"00",
		X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"16",X"11",X"91",X"89",X"33",X"E4",X"88",X"D9",
		X"00",X"08",X"86",X"E7",X"F3",X"71",X"20",X"20",X"00",X"00",X"00",X"00",X"08",X"C8",X"8C",X"44",
		X"11",X"11",X"01",X"10",X"00",X"00",X"00",X"00",X"FE",X"BB",X"99",X"DC",X"E6",X"22",X"10",X"00",
		X"F7",X"BD",X"F1",X"A0",X"F0",X"C0",X"80",X"80",X"44",X"C4",X"C0",X"88",X"00",X"80",X"00",X"00",
		X"00",X"00",X"12",X"02",X"13",X"13",X"02",X"13",X"0E",X"67",X"11",X"11",X"33",X"C8",X"AE",X"BB",
		X"00",X"08",X"8C",X"C6",X"F7",X"EA",X"75",X"57",X"00",X"00",X"00",X"00",X"08",X"8C",X"04",X"8C",
		X"02",X"13",X"01",X"11",X"00",X"00",X"00",X"00",X"64",X"56",X"BA",X"DD",X"EE",X"73",X"00",X"00",
		X"74",X"60",X"D0",X"B8",X"E0",X"C0",X"88",X"44",X"C0",X"48",X"C0",X"8C",X"44",X"00",X"00",X"00",
		X"00",X"01",X"00",X"04",X"26",X"26",X"13",X"02",X"00",X"0C",X"CF",X"31",X"52",X"40",X"CC",X"BB",
		X"00",X"00",X"08",X"8E",X"4D",X"E2",X"75",X"56",X"00",X"00",X"00",X"00",X"08",X"8C",X"04",X"8C",
		X"13",X"01",X"11",X"00",X"00",X"00",X"00",X"00",X"E8",X"74",X"76",X"88",X"89",X"77",X"00",X"00",
		X"31",X"50",X"B0",X"F8",X"30",X"C8",X"32",X"00",X"C8",X"44",X"6A",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"22",X"00",X"4C",X"14",X"04",X"00",X"00",X"0F",X"EA",X"FC",X"77",X"00",X"E6",
		X"00",X"00",X"08",X"07",X"99",X"E6",X"F9",X"76",X"00",X"00",X"00",X"80",X"08",X"8C",X"8C",X"04",
		X"13",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"39",X"14",X"31",X"88",X"55",X"33",X"00",X"00",
		X"20",X"70",X"74",X"B8",X"54",X"1C",X"00",X"00",X"F2",X"E0",X"80",X"80",X"00",X"88",X"00",X"00",
		X"00",X"00",X"00",X"07",X"22",X"00",X"CC",X"19",X"00",X"00",X"87",X"6E",X"F7",X"74",X"88",X"D4",
		X"00",X"00",X"2C",X"23",X"11",X"CC",X"F3",X"74",X"00",X"00",X"00",X"00",X"08",X"C0",X"C8",X"88",
		X"14",X"12",X"11",X"00",X"00",X"00",X"00",X"00",X"37",X"B8",X"02",X"99",X"66",X"31",X"00",X"00",
		X"20",X"B0",X"38",X"54",X"67",X"EC",X"00",X"00",X"84",X"80",X"C0",X"80",X"44",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"1E",X"44",X"00",X"CC",X"00",X"00",X"01",X"0E",X"D5",X"DA",X"88",X"C4",
		X"00",X"00",X"0E",X"01",X"5D",X"F3",X"9E",X"64",X"00",X"00",X"00",X"00",X"08",X"C0",X"A2",X"80",
		X"08",X"34",X"13",X"00",X"00",X"00",X"00",X"00",X"73",X"B0",X"8A",X"99",X"66",X"11",X"00",X"00",
		X"74",X"B2",X"DC",X"76",X"47",X"8C",X"00",X"00",X"80",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"16",X"18",X"00",X"00",X"00",X"00",X"07",X"19",X"FA",X"9F",X"98",
		X"00",X"00",X"0E",X"EF",X"AF",X"F1",X"FC",X"64",X"00",X"00",X"00",X"00",X"08",X"00",X"8C",X"80",
		X"00",X"98",X"66",X"11",X"00",X"00",X"00",X"00",X"6E",X"94",X"DD",X"88",X"77",X"00",X"00",X"00",
		X"30",X"92",X"EE",X"33",X"67",X"EE",X"00",X"00",X"C0",X"C0",X"C0",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"21",X"52",X"9D",X"00",X"00",X"21",X"06",X"19",X"BC",X"D9",X"90",
		X"00",X"C0",X"2C",X"47",X"F1",X"D5",X"FA",X"EE",X"00",X"00",X"00",X"40",X"44",X"08",X"80",X"C0",
		X"4C",X"00",X"44",X"DC",X"11",X"00",X"00",X"00",X"EE",X"B8",X"8C",X"08",X"FF",X"00",X"00",X"00",
		X"74",X"77",X"FE",X"33",X"FE",X"00",X"00",X"00",X"A4",X"62",X"C8",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"13",X"35",X"00",X"00",X"21",X"53",X"2E",X"B8",X"FB",X"7C",
		X"00",X"80",X"2C",X"DE",X"8C",X"F0",X"E8",X"FC",X"00",X"00",X"00",X"00",X"80",X"00",X"C0",X"F6",
		X"4D",X"CC",X"00",X"22",X"44",X"00",X"00",X"00",X"88",X"AA",X"64",X"F7",X"22",X"00",X"00",X"00",
		X"31",X"66",X"DD",X"99",X"02",X"00",X"00",X"00",X"60",X"C0",X"88",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"13",X"00",X"00",X"03",X"26",X"19",X"54",X"75",X"FE",
		X"00",X"00",X"48",X"9F",X"DA",X"F0",X"DC",X"DE",X"00",X"00",X"88",X"00",X"00",X"C0",X"C0",X"C0",
		X"26",X"15",X"4C",X"00",X"02",X"26",X"00",X"00",X"A2",X"EE",X"60",X"19",X"C4",X"AA",X"00",X"00",
		X"FE",X"22",X"88",X"00",X"23",X"44",X"00",X"00",X"84",X"CC",X"8C",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"02",X"00",X"00",X"43",X"84",X"3B",X"74",X"FB",X"C4",
		X"00",X"22",X"A2",X"64",X"78",X"50",X"7C",X"DC",X"00",X"00",X"00",X"00",X"80",X"E2",X"80",X"C4",
		X"13",X"00",X"36",X"44",X"44",X"00",X"11",X"00",X"00",X"66",X"76",X"11",X"64",X"73",X"CC",X"00",
		X"65",X"73",X"77",X"99",X"EE",X"88",X"00",X"00",X"C8",X"88",X"88",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"43",X"95",X"19",X"76",X"75",X"44",
		X"00",X"C4",X"C8",X"D0",X"F0",X"D8",X"FC",X"67",X"00",X"00",X"00",X"40",X"C4",X"00",X"C0",X"CC",
		X"13",X"13",X"12",X"22",X"22",X"32",X"00",X"00",X"C8",X"A2",X"B3",X"9A",X"11",X"21",X"64",X"A0",
		X"B3",X"66",X"04",X"99",X"AA",X"44",X"00",X"00",X"8C",X"8C",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"01",X"01",X"01",X"00",X"00",X"43",X"BF",X"19",X"BA",X"31",X"77",
		X"04",X"00",X"A0",X"F0",X"E9",X"B6",X"FA",X"FE",X"00",X"00",X"84",X"00",X"00",X"C0",X"8C",X"8C",
		X"01",X"01",X"01",X"11",X"00",X"00",X"11",X"00",X"44",X"AA",X"B3",X"36",X"90",X"11",X"10",X"46",
		X"F5",X"EA",X"C8",X"99",X"22",X"CC",X"08",X"00",X"CC",X"44",X"88",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"21",X"13",X"13",X"11",X"11",X"50",X"78",X"9C",X"ED",X"75",X"44",
		X"00",X"00",X"E0",X"F0",X"F0",X"B7",X"EC",X"22",X"00",X"00",X"00",X"80",X"08",X"48",X"AC",X"24",
		X"11",X"01",X"11",X"10",X"00",X"00",X"00",X"00",X"54",X"44",X"DD",X"FA",X"C8",X"88",X"44",X"55",
		X"A2",X"22",X"EA",X"C5",X"40",X"A0",X"44",X"00",X"04",X"C8",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"21",X"13",X"02",X"00",X"04",X"74",X"F4",X"3A",X"DE",X"73",X"73",
		X"00",X"02",X"E2",X"F2",X"C5",X"B7",X"EC",X"EC",X"00",X"00",X"00",X"00",X"80",X"48",X"8C",X"04",
		X"00",X"11",X"01",X"00",X"00",X"00",X"00",X"00",X"54",X"44",X"35",X"5D",X"AA",X"24",X"44",X"22",
		X"A2",X"22",X"CA",X"23",X"77",X"42",X"22",X"44",X"00",X"88",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"13",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"20",X"01",X"13",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",
		X"01",X"13",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"41",X"13",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"8C",X"18",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"8C",X"08",
		X"13",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"82",X"27",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"13",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",
		X"00",X"00",X"04",X"4E",X"04",X"10",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"8C",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"27",X"02",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"21",X"31",X"13",X"11",
		X"00",X"00",X"00",X"40",X"48",X"C8",X"8C",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"00",X"10",X"00",X"00",X"00",
		X"88",X"88",X"88",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"01",X"01",X"11",
		X"00",X"00",X"80",X"80",X"1C",X"AC",X"EC",X"8C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"31",X"33",X"33",X"25",X"36",X"02",X"00",X"00",
		X"08",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"11",
		X"00",X"00",X"00",X"00",X"40",X"84",X"DE",X"EC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"00",X"33",X"77",X"EE",X"CC",X"88",X"00",X"00",X"00",
		X"8C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"13",
		X"00",X"00",X"00",X"00",X"10",X"60",X"4F",X"CE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"13",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"82",X"08",X"00",X"00",X"00",X"00",X"00",
		X"DA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"34",X"EF",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EF",X"34",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"31",X"31",
		X"00",X"00",X"00",X"00",X"00",X"40",X"C8",X"C8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"01",
		X"00",X"00",X"00",X"00",X"80",X"6C",X"EC",X"C8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"31",X"02",X"11",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"01",
		X"00",X"00",X"00",X"00",X"00",X"80",X"0C",X"AC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"13",X"05",X"02",X"00",X"00",X"00",X"00",X"00",
		X"48",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"13",
		X"00",X"00",X"00",X"00",X"00",X"60",X"C6",X"56",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"46",X"00",X"00",X"00",X"00",X"00",X"00",
		X"68",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"40",X"00",
		X"00",X"44",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"88",X"00",X"00",X"00",
		X"00",X"20",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"11",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"13",X"22",X"70",X"60",X"00",X"30",X"0F",X"FF",X"FF",X"77",X"23",X"46",
		X"00",X"A4",X"3C",X"3C",X"8D",X"CB",X"7F",X"B7",X"00",X"00",X"80",X"08",X"48",X"48",X"2C",X"AC",
		X"51",X"07",X"10",X"00",X"11",X"00",X"00",X"00",X"D7",X"E3",X"D1",X"E0",X"60",X"88",X"33",X"00",
		X"37",X"5D",X"C8",X"14",X"34",X"34",X"BC",X"00",X"AC",X"AC",X"8C",X"8C",X"80",X"80",X"00",X"00",
		X"00",X"00",X"00",X"10",X"30",X"20",X"07",X"44",X"00",X"30",X"C3",X"FF",X"F7",X"33",X"E3",X"56",
		X"00",X"C0",X"3C",X"0F",X"8F",X"DE",X"6D",X"B7",X"00",X"00",X"00",X"08",X"C0",X"C0",X"0E",X"AC",
		X"54",X"30",X"10",X"22",X"11",X"00",X"00",X"00",X"C6",X"A3",X"D1",X"D0",X"02",X"CE",X"12",X"00",
		X"B7",X"5D",X"88",X"80",X"D1",X"E3",X"C0",X"00",X"AC",X"AC",X"8C",X"8C",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"13",X"22",X"44",X"44",X"00",X"30",X"61",X"31",X"19",X"15",X"23",X"57",
		X"00",X"C0",X"3C",X"0F",X"8F",X"EF",X"7F",X"2E",X"00",X"00",X"00",X"80",X"48",X"48",X"E0",X"60",
		X"54",X"30",X"10",X"22",X"00",X"00",X"00",X"00",X"C6",X"E3",X"91",X"44",X"CC",X"20",X"31",X"00",
		X"AF",X"7F",X"BB",X"11",X"11",X"23",X"CC",X"00",X"20",X"0E",X"8C",X"8C",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"13",X"22",X"44",X"44",X"00",X"12",X"C2",X"0E",X"FE",X"77",X"23",X"46",
		X"00",X"C0",X"F0",X"C3",X"87",X"EF",X"7F",X"BF",X"00",X"00",X"00",X"80",X"48",X"48",X"2C",X"AC",
		X"54",X"44",X"20",X"00",X"11",X"00",X"00",X"00",X"D6",X"23",X"99",X"C8",X"80",X"88",X"33",X"00",
		X"37",X"7C",X"8A",X"01",X"11",X"23",X"CC",X"00",X"AC",X"E0",X"C0",X"40",X"08",X"00",X"00",X"00",
		X"00",X"00",X"03",X"D3",X"14",X"13",X"00",X"00",X"00",X"03",X"3F",X"FF",X"C0",X"FC",X"77",X"66",
		X"00",X"0C",X"ED",X"FD",X"02",X"D3",X"CE",X"26",X"00",X"00",X"48",X"F8",X"42",X"C8",X"00",X"00",
		X"00",X"00",X"03",X"D3",X"14",X"13",X"00",X"00",X"76",X"43",X"3F",X"CC",X"F0",X"FC",X"33",X"00",
		X"E2",X"0E",X"ED",X"31",X"C2",X"D3",X"CC",X"00",X"00",X"00",X"48",X"F8",X"42",X"C8",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"01",X"97",X"6E",X"90",X"30",
		X"00",X"00",X"00",X"08",X"DA",X"27",X"94",X"C0",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",
		X"00",X"03",X"D3",X"94",X"13",X"00",X"00",X"00",X"43",X"3F",X"CC",X"F0",X"FD",X"32",X"00",X"00",
		X"2C",X"ED",X"31",X"C2",X"DB",X"C4",X"00",X"00",X"00",X"48",X"F8",X"52",X"C8",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"D3",X"00",X"00",X"00",X"00",X"00",X"03",X"3F",X"DC",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"ED",X"B1",X"00",X"00",X"00",X"00",X"00",X"00",X"48",X"F8",
		X"94",X"13",X"00",X"00",X"00",X"00",X"00",X"00",X"F1",X"FC",X"33",X"00",X"00",X"00",X"00",X"00",
		X"CA",X"D3",X"CC",X"00",X"00",X"00",X"00",X"00",X"52",X"C8",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"D3",X"94",X"13",X"00",X"00",X"00",X"12",X"2E",X"FF",X"C0",X"FC",X"33",
		X"00",X"00",X"84",X"65",X"FD",X"02",X"D3",X"CC",X"00",X"00",X"00",X"48",X"F8",X"52",X"C8",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"86",X"7F",X"90",X"11",X"00",X"00",X"00",
		X"00",X"52",X"AF",X"94",X"88",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"07",X"99",X"40",X"60",X"52",X"43",X"21",X"10",X"00",X"8C",X"46",X"23",X"81",X"E3",X"4E",X"0F",
		X"00",X"20",X"60",X"C0",X"08",X"00",X"88",X"45",X"00",X"00",X"00",X"00",X"00",X"20",X"60",X"C0",
		X"00",X"10",X"20",X"00",X"00",X"00",X"00",X"00",X"B1",X"10",X"00",X"10",X"00",X"10",X"20",X"00",
		X"09",X"6B",X"4E",X"3C",X"96",X"43",X"30",X"00",X"08",X"8C",X"46",X"02",X"23",X"81",X"C1",X"22",
		X"07",X"99",X"40",X"60",X"52",X"43",X"21",X"10",X"00",X"0C",X"46",X"23",X"91",X"C2",X"4A",X"8F",
		X"10",X"30",X"60",X"48",X"08",X"00",X"88",X"45",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B1",X"10",X"00",X"10",X"00",X"10",X"20",X"40",
		X"18",X"6B",X"60",X"3C",X"96",X"43",X"30",X"00",X"08",X"8C",X"46",X"02",X"23",X"81",X"C1",X"22",
		X"07",X"99",X"40",X"60",X"52",X"43",X"21",X"10",X"00",X"0C",X"46",X"33",X"80",X"C0",X"2C",X"87",
		X"00",X"40",X"C8",X"80",X"08",X"00",X"88",X"45",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"88",
		X"32",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"B1",X"10",X"00",X"10",X"00",X"32",X"00",X"00",
		X"19",X"48",X"E0",X"B4",X"96",X"43",X"30",X"00",X"00",X"8C",X"46",X"02",X"23",X"81",X"C1",X"22",
		X"07",X"99",X"40",X"60",X"52",X"43",X"21",X"01",X"00",X"0C",X"46",X"23",X"90",X"E3",X"68",X"0F",
		X"00",X"00",X"00",X"00",X"08",X"00",X"88",X"45",X"00",X"00",X"00",X"00",X"10",X"30",X"60",X"48",
		X"10",X"20",X"40",X"80",X"00",X"00",X"00",X"00",X"B1",X"10",X"00",X"10",X"00",X"00",X"00",X"00",
		X"19",X"48",X"4A",X"BC",X"96",X"43",X"30",X"00",X"08",X"8C",X"46",X"02",X"23",X"81",X"C1",X"22",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"11",X"10",X"30",X"07",X"7F",X"88",
		X"00",X"FF",X"FF",X"80",X"C0",X"2C",X"9E",X"DE",X"88",X"88",X"88",X"77",X"66",X"66",X"66",X"E6",
		X"10",X"00",X"00",X"00",X"E0",X"10",X"10",X"10",X"A8",X"98",X"44",X"33",X"10",X"00",X"00",X"00",
		X"56",X"56",X"46",X"8C",X"80",X"00",X"00",X"00",X"C4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"CE",X"EE",X"EE",X"FE",X"77",X"77",X"77",X"10",X"30",X"07",X"7F",X"88",
		X"FF",X"EF",X"CF",X"80",X"C0",X"2C",X"9E",X"DE",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"80",
		X"FE",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"A8",X"98",X"44",X"33",X"10",X"00",X"00",X"00",
		X"56",X"56",X"46",X"8C",X"80",X"10",X"10",X"10",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"0E",X"1E",X"03",X"43",X"43",X"10",X"30",X"07",X"7F",X"88",
		X"2C",X"68",X"E0",X"80",X"C0",X"2C",X"9E",X"DE",X"00",X"00",X"00",X"00",X"00",X"07",X"60",X"C0",
		X"1E",X"0E",X"E0",X"00",X"00",X"00",X"00",X"00",X"A8",X"DC",X"66",X"33",X"10",X"00",X"00",X"00",
		X"56",X"56",X"46",X"8C",X"80",X"20",X"60",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"10",X"10",X"10",X"30",X"43",X"B7",X"4C",
		X"00",X"00",X"00",X"80",X"C0",X"2C",X"9E",X"DE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A8",X"98",X"44",X"33",X"10",X"00",X"10",X"10",
		X"56",X"56",X"46",X"8C",X"80",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"10",X"00",X"00",X"00",X"10",X"30",X"07",X"7F",X"88",
		X"02",X"02",X"02",X"80",X"C0",X"2C",X"9E",X"DE",X"00",X"00",X"00",X"00",X"00",X"70",X"61",X"C3",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A8",X"98",X"66",X"13",X"10",X"43",X"43",X"43",
		X"56",X"56",X"46",X"8C",X"80",X"2C",X"0E",X"0E",X"C3",X"07",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"30",X"07",X"7F",X"88",
		X"10",X"10",X"10",X"80",X"C0",X"2C",X"9E",X"DE",X"00",X"00",X"00",X"00",X"17",X"17",X"37",X"B7",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A8",X"98",X"44",X"33",X"10",X"77",X"77",X"77",
		X"56",X"56",X"46",X"8C",X"80",X"EF",X"FF",X"FF",X"F7",X"77",X"77",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"44",X"88",X"00",X"00",X"C0",X"00",X"0F",X"FF",X"FF",X"00",X"03",X"F0",X"AD",
		X"00",X"1E",X"DC",X"CC",X"DC",X"2E",X"B4",X"61",X"00",X"08",X"48",X"A4",X"9E",X"00",X"00",X"08",
		X"C0",X"00",X"00",X"B8",X"54",X"33",X"00",X"00",X"AD",X"88",X"30",X"C0",X"F0",X"70",X"88",X"00",
		X"68",X"B5",X"A6",X"54",X"00",X"10",X"FE",X"00",X"88",X"00",X"00",X"EF",X"C6",X"48",X"08",X"00",
		X"00",X"00",X"21",X"16",X"E8",X"00",X"00",X"01",X"00",X"0F",X"FF",X"FF",X"C0",X"47",X"9E",X"6D",
		X"00",X"0F",X"FF",X"EF",X"FC",X"2E",X"97",X"63",X"00",X"00",X"48",X"86",X"70",X"00",X"00",X"08",
		X"11",X"00",X"00",X"B8",X"54",X"33",X"00",X"00",X"61",X"98",X"21",X"D1",X"E0",X"60",X"98",X"10",
		X"68",X"D1",X"48",X"D9",X"40",X"40",X"F3",X"80",X"88",X"00",X"00",X"EF",X"CE",X"8C",X"00",X"00",
		X"00",X"01",X"03",X"44",X"88",X"00",X"00",X"01",X"00",X"C3",X"A1",X"21",X"32",X"47",X"96",X"6D",
		X"00",X"1E",X"EF",X"FF",X"FF",X"0C",X"F0",X"DB",X"00",X"00",X"48",X"AC",X"DE",X"00",X"00",X"30",
		X"11",X"00",X"00",X"B8",X"54",X"23",X"01",X"00",X"61",X"9A",X"56",X"B2",X"30",X"B0",X"C0",X"00",
		X"5B",X"11",X"C0",X"11",X"00",X"00",X"FF",X"00",X"30",X"00",X"00",X"EF",X"CE",X"8C",X"00",X"00",
		X"00",X"00",X"03",X"44",X"88",X"00",X"00",X"01",X"10",X"1E",X"EE",X"EE",X"11",X"03",X"96",X"6D",
		X"80",X"D2",X"63",X"73",X"FB",X"0C",X"D2",X"63",X"00",X"00",X"48",X"AC",X"DE",X"00",X"00",X"08",
		X"11",X"00",X"00",X"E8",X"16",X"33",X"00",X"00",X"E1",X"9E",X"74",X"C0",X"F0",X"70",X"88",X"00",
		X"78",X"97",X"E2",X"11",X"00",X"00",X"FF",X"00",X"88",X"00",X"00",X"70",X"8E",X"8C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"22",X"EE",X"67",X"13",X"13",X"33",X"0C",
		X"00",X"08",X"6E",X"CC",X"08",X"08",X"08",X"8F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",
		X"7F",X"88",X"30",X"00",X"00",X"00",X"00",X"00",X"CC",X"31",X"E0",X"20",X"10",X"FF",X"00",X"00",
		X"BF",X"8C",X"8C",X"88",X"88",X"00",X"00",X"00",X"CE",X"22",X"44",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"22",X"EE",X"67",X"13",X"13",X"33",X"0C",
		X"00",X"08",X"6E",X"CC",X"08",X"08",X"08",X"8F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",
		X"7F",X"88",X"30",X"00",X"00",X"00",X"00",X"00",X"CC",X"31",X"E0",X"20",X"10",X"11",X"00",X"00",
		X"BF",X"8C",X"8C",X"88",X"88",X"EE",X"00",X"00",X"CE",X"22",X"44",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"21",X"43",X"47",X"67",X"77",X"77",X"0F",X"0F",X"78",X"3D",X"1E",X"0F",X"0F",X"8F",
		X"0F",X"0F",X"E1",X"CB",X"87",X"0F",X"0F",X"1E",X"08",X"0C",X"0E",X"0F",X"0F",X"4B",X"C3",X"CB",
		X"77",X"77",X"66",X"44",X"66",X"33",X"11",X"00",X"88",X"00",X"00",X"11",X"33",X"77",X"FF",X"00",
		X"1E",X"0F",X"0F",X"8F",X"CF",X"EF",X"FF",X"00",X"CB",X"C3",X"4B",X"0F",X"2C",X"48",X"80",X"00",
		X"00",X"10",X"21",X"43",X"47",X"67",X"77",X"77",X"0F",X"0F",X"78",X"3D",X"1E",X"1E",X"1E",X"AC",
		X"0F",X"0F",X"E1",X"CB",X"87",X"87",X"87",X"70",X"08",X"0C",X"0E",X"0F",X"0F",X"4B",X"C3",X"CB",
		X"77",X"77",X"66",X"44",X"66",X"33",X"11",X"00",X"8F",X"01",X"01",X"11",X"33",X"77",X"FF",X"00",
		X"16",X"87",X"0F",X"8F",X"CF",X"EF",X"FF",X"00",X"CB",X"C3",X"4B",X"0F",X"2C",X"48",X"80",X"00",
		X"00",X"10",X"21",X"43",X"47",X"67",X"77",X"77",X"0F",X"0F",X"78",X"3D",X"1E",X"1E",X"68",X"8C",
		X"0F",X"0F",X"E1",X"CB",X"C3",X"C3",X"F0",X"70",X"08",X"0C",X"0E",X"0F",X"0F",X"4B",X"C3",X"CB",
		X"77",X"77",X"66",X"44",X"66",X"33",X"11",X"00",X"9D",X"0E",X"03",X"13",X"33",X"77",X"FF",X"00",
		X"30",X"43",X"4B",X"8F",X"CF",X"EF",X"FF",X"00",X"CB",X"C3",X"4B",X"0F",X"2C",X"48",X"80",X"00",
		X"00",X"00",X"01",X"03",X"07",X"9F",X"DC",X"DC",X"03",X"F0",X"78",X"0F",X"FF",X"3F",X"3D",X"B7",
		X"0E",X"E1",X"C3",X"4B",X"ED",X"98",X"19",X"BF",X"00",X"00",X"08",X"0C",X"0E",X"2D",X"E1",X"69",
		X"DC",X"DC",X"DC",X"88",X"00",X"00",X"00",X"00",X"F7",X"95",X"1F",X"3C",X"70",X"00",X"77",X"FF",
		X"FF",X"FB",X"1F",X"97",X"E3",X"03",X"CF",X"EE",X"69",X"69",X"69",X"2C",X"0C",X"08",X"00",X"00",
		X"00",X"00",X"01",X"03",X"07",X"9F",X"DC",X"DC",X"03",X"F0",X"78",X"0F",X"FF",X"3F",X"3D",X"B7",
		X"0E",X"E1",X"C3",X"4B",X"ED",X"98",X"19",X"BF",X"00",X"00",X"08",X"0C",X"0E",X"2D",X"E1",X"69",
		X"DD",X"DC",X"DC",X"88",X"00",X"00",X"00",X"00",X"FF",X"B7",X"1F",X"3D",X"71",X"00",X"77",X"FF",
		X"FF",X"FB",X"1F",X"97",X"E3",X"03",X"CF",X"EE",X"69",X"69",X"69",X"2C",X"0C",X"08",X"00",X"00",
		X"00",X"00",X"01",X"03",X"07",X"9F",X"DD",X"DD",X"03",X"F0",X"78",X"0F",X"FF",X"FF",X"FF",X"FF",
		X"0E",X"E1",X"C3",X"4B",X"ED",X"FE",X"FF",X"FF",X"00",X"00",X"08",X"0C",X"0E",X"2D",X"E1",X"69",
		X"DD",X"DD",X"DD",X"88",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"77",X"00",X"77",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"EF",X"03",X"CF",X"EE",X"69",X"69",X"69",X"2C",X"0C",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"23",X"00",X"9E",X"56",X"76",X"76",X"76",X"76",X"56",
		X"00",X"80",X"08",X"08",X"08",X"08",X"80",X"BC",X"00",X"00",X"00",X"00",X"00",X"20",X"52",X"D6",
		X"77",X"44",X"44",X"44",X"00",X"00",X"00",X"00",X"83",X"A3",X"B2",X"81",X"81",X"81",X"81",X"98",
		X"3F",X"EF",X"80",X"88",X"88",X"00",X"00",X"08",X"20",X"F7",X"63",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"44",X"44",X"67",X"00",X"9E",X"56",X"76",X"76",X"76",X"76",X"56",
		X"00",X"80",X"08",X"08",X"08",X"08",X"80",X"BC",X"00",X"00",X"00",X"00",X"00",X"20",X"52",X"D6",
		X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"83",X"A3",X"B2",X"81",X"81",X"81",X"81",X"98",
		X"3F",X"EF",X"80",X"88",X"88",X"00",X"00",X"08",X"20",X"F7",X"63",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"13",X"32",X"74",X"44",X"00",X"03",X"3F",X"FF",X"FF",X"88",X"92",X"02",
		X"00",X"0C",X"CF",X"FF",X"FF",X"00",X"B4",X"04",X"00",X"00",X"00",X"08",X"8C",X"8C",X"68",X"68",
		X"77",X"55",X"00",X"22",X"11",X"00",X"00",X"00",X"13",X"03",X"00",X"00",X"30",X"98",X"22",X"00",
		X"AE",X"0F",X"00",X"00",X"C0",X"81",X"44",X"00",X"28",X"0E",X"44",X"04",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"00",X"30",X"16",X"0F",X"0F",X"CB",X"C3",X"C3",
		X"00",X"C0",X"E0",X"1E",X"0F",X"0F",X"25",X"25",X"00",X"00",X"00",X"00",X"00",X"08",X"80",X"80",
		X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C3",X"43",X"83",X"63",X"51",X"20",X"33",X"00",
		X"25",X"0F",X"0F",X"0F",X"1E",X"46",X"CC",X"00",X"80",X"08",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"23",X"33",X"33",X"11",
		X"00",X"80",X"C0",X"C0",X"48",X"E0",X"C2",X"42",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"10",X"32",X"00",X"11",X"00",
		X"42",X"42",X"E0",X"48",X"0C",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"00",X"03",X"07",X"F8",X"03",X"E9",X"61",X"01",
		X"00",X"0C",X"0E",X"CF",X"E7",X"73",X"73",X"51",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"08",
		X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"03",X"61",X"61",X"08",X"07",X"30",X"33",X"00",
		X"51",X"51",X"15",X"59",X"E3",X"46",X"8C",X"00",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"00",X"33",X"77",X"77",X"00",X"03",X"0F",X"00",X"8F",X"01",X"01",X"EF",
		X"00",X"48",X"1E",X"0F",X"03",X"8B",X"CD",X"CD",X"00",X"00",X"00",X"80",X"48",X"0C",X"2C",X"2C",
		X"77",X"77",X"33",X"03",X"00",X"00",X"00",X"00",X"8F",X"01",X"01",X"FF",X"0F",X"62",X"00",X"00",
		X"DD",X"DF",X"FF",X"3F",X"77",X"67",X"CC",X"00",X"2C",X"2C",X"0C",X"0C",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"57",X"11",X"11",X"00",X"00",X"00",
		X"06",X"06",X"DF",X"44",X"C4",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"88",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"20",X"01",X"22",X"00",X"01",X"11",
		X"00",X"00",X"0E",X"0D",X"2B",X"CF",X"00",X"C4",X"00",X"00",X"00",X"00",X"80",X"00",X"88",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"10",X"34",X"20",X"32",X"CC",X"46",X"CC",
		X"84",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",
		X"00",X"00",X"46",X"8E",X"1D",X"2A",X"41",X"83",X"00",X"00",X"00",X"00",X"00",X"0C",X"4C",X"88",
		X"00",X"00",X"01",X"02",X"33",X"11",X"00",X"00",X"14",X"A0",X"45",X"A8",X"04",X"08",X"00",X"00",
		X"04",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"26",
		X"00",X"00",X"00",X"45",X"03",X"13",X"AA",X"B3",X"00",X"00",X"80",X"08",X"08",X"00",X"88",X"0C",
		X"10",X"11",X"EE",X"9A",X"00",X"00",X"00",X"00",X"B8",X"51",X"44",X"00",X"00",X"00",X"00",X"00",
		X"44",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"66",X"07",X"CF",
		X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"CF",X"07",X"66",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"66",X"77",X"44",X"00",X"00",X"00",X"33",X"11",X"11",X"99",X"FF",X"33",X"00",
		X"40",X"40",X"40",X"70",X"70",X"40",X"00",X"00",X"00",X"90",X"90",X"90",X"F0",X"F0",X"30",X"00",
		X"33",X"66",X"44",X"66",X"77",X"44",X"00",X"00",X"88",X"CC",X"44",X"44",X"CC",X"FF",X"33",X"00",
		X"30",X"70",X"40",X"40",X"70",X"40",X"00",X"00",X"00",X"B0",X"F0",X"C0",X"80",X"F0",X"30",X"00",
		X"66",X"11",X"00",X"33",X"77",X"66",X"00",X"00",X"00",X"00",X"CC",X"FF",X"33",X"00",X"00",X"00",
		X"30",X"30",X"60",X"40",X"70",X"40",X"00",X"00",X"C0",X"E0",X"30",X"10",X"90",X"F0",X"30",X"00",
		X"00",X"77",X"77",X"66",X"55",X"00",X"00",X"00",X"11",X"FF",X"FF",X"44",X"44",X"CC",X"77",X"00",
		X"00",X"70",X"70",X"60",X"50",X"00",X"00",X"00",X"10",X"F0",X"F0",X"40",X"40",X"C0",X"70",X"00",
		X"33",X"77",X"44",X"44",X"77",X"44",X"00",X"00",X"00",X"BB",X"FF",X"CC",X"88",X"FF",X"33",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"44",X"44",X"77",X"77",X"44",X"00",X"00",X"00",X"99",X"99",X"99",X"FF",X"FF",X"33",X"00",
		X"60",X"10",X"00",X"30",X"70",X"60",X"00",X"00",X"00",X"00",X"C0",X"F0",X"30",X"00",X"00",X"00",
		X"66",X"11",X"00",X"11",X"77",X"11",X"00",X"00",X"00",X"CC",X"77",X"FF",X"CC",X"88",X"77",X"00",
		X"60",X"10",X"10",X"70",X"00",X"10",X"70",X"00",X"00",X"C0",X"F0",X"80",X"40",X"F0",X"80",X"00",
		X"33",X"77",X"44",X"44",X"66",X"33",X"00",X"00",X"88",X"EE",X"33",X"11",X"11",X"FF",X"EE",X"00",
		X"40",X"40",X"60",X"70",X"50",X"40",X"00",X"00",X"00",X"00",X"00",X"C0",X"F0",X"30",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"44",X"44",X"77",X"77",X"44",X"00",X"00",X"00",X"99",X"99",X"99",X"FF",X"FF",X"33",X"00",
		X"30",X"70",X"40",X"40",X"60",X"30",X"00",X"00",X"80",X"E0",X"30",X"10",X"10",X"F0",X"E0",X"00",
		X"7F",X"FF",X"0F",X"CE",X"CE",X"DF",X"5F",X"07",X"EF",X"CE",X"0C",X"00",X"00",X"CE",X"EF",X"0F",
		X"FF",X"7F",X"0F",X"00",X"07",X"7F",X"FF",X"0F",X"EF",X"FF",X"0F",X"37",X"3F",X"BF",X"AF",X"0E",
		X"07",X"7F",X"FF",X"0F",X"00",X"00",X"00",X"00",X"0E",X"CF",X"EF",X"0F",X"00",X"00",X"00",X"00",
		X"07",X"7F",X"FF",X"0F",X"00",X"00",X"00",X"00",X"0E",X"EF",X"FF",X"0F",X"00",X"00",X"00",X"00",
		X"7F",X"FF",X"0F",X"CE",X"CF",X"DF",X"5F",X"07",X"EF",X"CE",X"0C",X"00",X"0C",X"CE",X"EF",X"0F",
		X"FF",X"7F",X"07",X"00",X"00",X"7F",X"FF",X"0F",X"EF",X"FF",X"0F",X"37",X"37",X"BF",X"AF",X"0A",
		X"7F",X"FF",X"0F",X"CE",X"CE",X"CE",X"4E",X"06",X"EF",X"CF",X"1F",X"13",X"13",X"01",X"01",X"01",
		X"00",X"08",X"8C",X"8C",X"8F",X"3F",X"FF",X"0F",X"01",X"13",X"37",X"37",X"3F",X"BF",X"AF",X"0E",
		X"7F",X"FF",X"0F",X"CE",X"CF",X"DF",X"5F",X"05",X"EF",X"CE",X"0C",X"00",X"0C",X"CE",X"EF",X"0E",
		X"FF",X"7F",X"07",X"00",X"07",X"7F",X"FF",X"0F",X"EE",X"FF",X"0F",X"37",X"3F",X"BF",X"AF",X"0A",
		X"07",X"7F",X"FF",X"0F",X"CE",X"CE",X"CE",X"4E",X"0E",X"EF",X"CE",X"1F",X"13",X"13",X"01",X"00",
		X"0F",X"FF",X"3F",X"8F",X"8C",X"8C",X"08",X"00",X"0E",X"EF",X"FF",X"0F",X"37",X"37",X"37",X"27",
		X"77",X"FF",X"0F",X"CE",X"CF",X"DF",X"5F",X"05",X"EF",X"CE",X"0C",X"00",X"0C",X"CE",X"EF",X"0E",
		X"FF",X"7F",X"07",X"00",X"07",X"7F",X"FF",X"0F",X"EF",X"FF",X"0F",X"37",X"3F",X"BF",X"AF",X"0A",
		X"00",X"08",X"8C",X"CE",X"CE",X"CF",X"DF",X"5F",X"00",X"01",X"01",X"13",X"13",X"1F",X"CF",X"EF",
		X"00",X"FF",X"3F",X"8F",X"8C",X"8C",X"8C",X"08",X"00",X"EE",X"FF",X"0F",X"37",X"37",X"37",X"27",
		X"7F",X"FF",X"0F",X"CE",X"CF",X"DF",X"5F",X"07",X"EF",X"CE",X"0C",X"00",X"0C",X"CE",X"EF",X"0E",
		X"FF",X"7F",X"07",X"00",X"07",X"7F",X"FF",X"0F",X"EF",X"FF",X"0F",X"37",X"3F",X"BF",X"AF",X"0E",
		X"7F",X"FF",X"0F",X"CE",X"CF",X"DF",X"5F",X"05",X"CE",X"EF",X"1F",X"13",X"1F",X"EF",X"CE",X"0E",
		X"37",X"7F",X"8F",X"8C",X"8F",X"7F",X"37",X"07",X"EF",X"FF",X"0F",X"37",X"3F",X"BF",X"AF",X"0A",
		X"7F",X"FF",X"0F",X"CE",X"CF",X"DF",X"5F",X"07",X"EF",X"CE",X"0C",X"00",X"0C",X"CE",X"EF",X"0E",
		X"FF",X"7F",X"07",X"00",X"07",X"7F",X"FF",X"0F",X"EF",X"FF",X"0F",X"33",X"3B",X"BF",X"AF",X"0E",
		X"7F",X"FF",X"0F",X"CE",X"CF",X"DF",X"5F",X"05",X"EF",X"CE",X"0C",X"00",X"0C",X"CE",X"EF",X"0E",
		X"FF",X"7F",X"07",X"00",X"07",X"7F",X"FF",X"0F",X"EF",X"FF",X"0F",X"37",X"3F",X"BF",X"AF",X"0A",
		X"00",X"00",X"00",X"01",X"02",X"11",X"11",X"37",X"00",X"01",X"16",X"19",X"77",X"FF",X"FF",X"FF",
		X"00",X"08",X"84",X"CA",X"ED",X"DC",X"CC",X"FF",X"00",X"00",X"00",X"00",X"08",X"84",X"CA",X"42",
		X"33",X"33",X"11",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"00",X"00",
		X"FF",X"EE",X"EE",X"CC",X"CC",X"12",X"04",X"00",X"42",X"84",X"84",X"84",X"84",X"08",X"00",X"00",
		X"00",X"01",X"12",X"02",X"15",X"33",X"77",X"77",X"0F",X"C2",X"11",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0C",X"03",X"DC",X"EE",X"FF",X"FF",X"FF",X"FF",X"00",X"08",X"84",X"42",X"42",X"A9",X"CD",X"A9",
		X"77",X"FF",X"77",X"77",X"33",X"11",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"00",X"70",X"CD",X"CD",X"A9",X"CA",X"04",X"84",X"84",X"08",
		X"00",X"01",X"30",X"00",X"33",X"77",X"77",X"FF",X"49",X"D2",X"20",X"CC",X"FF",X"FF",X"FF",X"FF",
		X"84",X"D2",X"10",X"CC",X"E2",X"F5",X"FE",X"FD",X"00",X"08",X"84",X"C2",X"60",X"43",X"B8",X"02",
		X"FF",X"FF",X"77",X"77",X"73",X"51",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"10",X"61",X"A9",X"98",X"21",X"42",X"40",X"C0",X"84",X"00",
		X"02",X"70",X"10",X"20",X"20",X"20",X"51",X"91",X"01",X"78",X"40",X"33",X"77",X"FF",X"FF",X"FF",
		X"0C",X"E1",X"42",X"CC",X"FF",X"FF",X"FF",X"EE",X"00",X"08",X"86",X"04",X"40",X"42",X"42",X"30",
		X"51",X"11",X"00",X"20",X"20",X"50",X"00",X"00",X"FF",X"FF",X"FF",X"77",X"33",X"C0",X"20",X"10",
		X"EE",X"FF",X"FF",X"EE",X"88",X"70",X"80",X"00",X"21",X"42",X"42",X"40",X"40",X"C2",X"0E",X"02",
		X"00",X"40",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"10",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"20",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A8",X"64",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"40",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"22",X"00",X"22",X"64",X"11",X"00",X"C8",X"80",X"10",X"00",X"00",X"00",
		X"00",X"00",X"31",X"10",X"88",X"80",X"00",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"C4",X"40",
		X"00",X"00",X"22",X"00",X"11",X"00",X"00",X"00",X"64",X"22",X"00",X"00",X"80",X"88",X"11",X"00",
		X"00",X"11",X"00",X"10",X"31",X"00",X"00",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"33",X"32",X"80",X"00",X"00",X"40",X"00",X"00",X"80",X"44",X"04",X"11",
		X"00",X"00",X"00",X"44",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"40",X"88",
		X"20",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"62",X"00",X"00",X"80",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"22",X"00",X"00",X"11",X"00",X"88",X"00",X"00",X"22",X"00",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"44",X"00",
		X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"22",X"00",X"00",X"22",X"00",X"00",
		X"00",X"00",X"00",X"00",X"44",X"00",X"44",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"00",X"11",X"00",X"00",X"22",X"40",X"00",X"22",X"40",X"00",X"98",X"44",X"77",X"77",
		X"00",X"00",X"44",X"80",X"10",X"80",X"60",X"88",X"00",X"00",X"80",X"00",X"00",X"23",X"91",X"00",
		X"00",X"11",X"20",X"00",X"00",X"00",X"10",X"00",X"BB",X"77",X"33",X"11",X"44",X"88",X"00",X"00",
		X"EC",X"DC",X"CC",X"AA",X"11",X"00",X"00",X"10",X"00",X"00",X"40",X"00",X"00",X"88",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"11",X"00",X"00",X"88",X"23",X"F6",X"CC",X"88",X"91",
		X"00",X"00",X"01",X"0C",X"96",X"47",X"67",X"98",X"00",X"00",X"00",X"08",X"04",X"00",X"08",X"08",
		X"11",X"11",X"00",X"20",X"10",X"00",X"00",X"00",X"91",X"20",X"40",X"18",X"33",X"80",X"00",X"00",
		X"98",X"11",X"33",X"E7",X"CC",X"00",X"00",X"00",X"08",X"88",X"00",X"44",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"21",X"74",X"74",X"AD",X"A5",X"E5",
		X"00",X"44",X"48",X"E2",X"E2",X"5B",X"5A",X"7A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"31",X"31",X"20",X"00",X"00",X"00",X"85",X"0C",X"B0",X"B0",X"B0",X"83",X"B0",X"30",
		X"1A",X"03",X"D0",X"D0",X"D0",X"1C",X"D0",X"C0",X"80",X"80",X"C8",X"C8",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"00",X"2C",X"E1",X"E1",X"0F",X"0F",X"87",X"87",
		X"00",X"00",X"00",X"4C",X"26",X"A4",X"0B",X"5A",X"00",X"00",X"00",X"00",X"00",X"88",X"C4",X"48",
		X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"D0",X"E5",X"A4",X"96",X"F0",X"43",X"10",
		X"E1",X"E1",X"A4",X"48",X"00",X"00",X"81",X"80",X"A6",X"C0",X"48",X"48",X"00",X"88",X"00",X"00",
		X"00",X"10",X"00",X"40",X"74",X"03",X"22",X"10",X"00",X"08",X"A6",X"86",X"C3",X"96",X"0F",X"07",
		X"00",X"00",X"00",X"CC",X"D1",X"0F",X"26",X"5B",X"00",X"00",X"00",X"00",X"88",X"C4",X"6A",X"24",
		X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"A5",X"87",X"A5",X"96",X"87",X"43",X"21",X"00",
		X"61",X"F0",X"78",X"AC",X"C4",X"4A",X"2D",X"00",X"8A",X"28",X"04",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"22",X"25",X"34",X"BC",X"47",X"00",X"00",X"00",X"DD",X"1C",X"87",X"1E",X"0F",
		X"00",X"00",X"00",X"BB",X"C3",X"36",X"1D",X"C3",X"00",X"00",X"00",X"08",X"84",X"4A",X"A2",X"28",
		X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"21",X"E2",X"C3",X"61",X"30",X"00",X"00",
		X"F0",X"78",X"A4",X"00",X"0C",X"A6",X"C0",X"00",X"0F",X"01",X"02",X"06",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"43",X"12",X"00",X"00",X"00",X"11",X"74",X"8F",X"0F",X"87",
		X"00",X"00",X"66",X"C3",X"B4",X"0F",X"78",X"38",X"00",X"00",X"00",X"0C",X"CC",X"19",X"91",X"80",
		X"12",X"43",X"00",X"00",X"00",X"00",X"00",X"00",X"87",X"0F",X"70",X"70",X"10",X"00",X"00",X"00",
		X"1A",X"4B",X"0F",X"87",X"C3",X"70",X"00",X"00",X"80",X"78",X"0C",X"0C",X"0C",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"23",X"00",X"31",X"76",X"A9",X"CB",X"C3",X"3C",X"4B",
		X"00",X"62",X"84",X"49",X"86",X"68",X"E0",X"61",X"00",X"00",X"00",X"88",X"46",X"02",X"00",X"08",
		X"16",X"70",X"34",X"07",X"03",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"3C",X"70",X"00",X"00",X"00",
		X"87",X"38",X"07",X"C3",X"F0",X"00",X"00",X"00",X"E0",X"84",X"08",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"23",X"47",X"9E",X"45",X"85",X"96",X"05",
		X"00",X"4E",X"9F",X"0C",X"48",X"E0",X"78",X"25",X"00",X"00",X"00",X"88",X"44",X"20",X"60",X"C2",
		X"00",X"01",X"23",X"16",X"01",X"00",X"00",X"00",X"4B",X"0F",X"96",X"E1",X"96",X"68",X"00",X"00",
		X"DA",X"03",X"0F",X"C3",X"48",X"00",X"00",X"00",X"2C",X"68",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"10",X"11",X"11",X"00",X"56",X"DB",X"BD",X"A5",X"A5",X"D2",X"C2",
		X"08",X"AF",X"19",X"08",X"C0",X"F0",X"E1",X"2D",X"00",X"00",X"88",X"00",X"04",X"48",X"C2",X"0C",
		X"10",X"10",X"00",X"00",X"01",X"00",X"00",X"00",X"87",X"87",X"0F",X"0F",X"69",X"69",X"1E",X"00",
		X"58",X"0D",X"0F",X"3C",X"68",X"80",X"00",X"00",X"E8",X"4A",X"84",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"11",X"31",X"21",X"21",X"30",X"10",X"26",X"15",X"84",X"B4",X"B4",X"A5",X"0E",X"85",
		X"46",X"8A",X"12",X"D2",X"D2",X"5A",X"07",X"1A",X"00",X"00",X"88",X"C8",X"48",X"48",X"C0",X"80",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C5",X"E5",X"A5",X"30",X"12",X"03",X"00",X"00",
		X"3A",X"7A",X"5A",X"C0",X"84",X"0C",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"22",X"70",X"65",X"00",X"10",X"12",X"04",X"91",X"C4",X"10",X"10",
		X"00",X"80",X"84",X"02",X"98",X"32",X"80",X"80",X"00",X"00",X"00",X"00",X"88",X"44",X"E0",X"6A",
		X"61",X"60",X"70",X"70",X"12",X"01",X"00",X"00",X"10",X"10",X"10",X"10",X"01",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"08",X"00",X"00",X"00",X"68",X"E0",X"E0",X"E0",X"84",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"13",X"32",X"20",X"00",X"60",X"60",X"00",X"E7",X"E3",X"B0",X"58",
		X"00",X"00",X"FF",X"20",X"21",X"09",X"0C",X"84",X"00",X"00",X"00",X"88",X"44",X"62",X"62",X"60",
		X"70",X"70",X"70",X"30",X"03",X"01",X"00",X"00",X"7A",X"08",X"80",X"80",X"80",X"0C",X"40",X"00",
		X"84",X"80",X"0C",X"00",X"00",X"00",X"00",X"00",X"60",X"03",X"06",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"30",X"30",X"30",X"21",X"30",X"70",X"00",X"00",X"76",X"93",X"83",X"21",X"78",X"92",
		X"00",X"66",X"F9",X"94",X"CA",X"08",X"08",X"80",X"00",X"00",X"00",X"88",X"C0",X"E0",X"E0",X"42",
		X"71",X"61",X"70",X"30",X"01",X"00",X"00",X"00",X"E3",X"88",X"08",X"C0",X"E0",X"78",X"07",X"00",
		X"C0",X"48",X"00",X"00",X"00",X"00",X"08",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"70",X"70",X"00",X"00",X"00",X"36",X"44",X"88",X"8E",X"C1",X"78",
		X"00",X"EE",X"F1",X"30",X"0C",X"88",X"08",X"00",X"00",X"00",X"00",X"CC",X"C0",X"20",X"00",X"00",
		X"10",X"30",X"10",X"10",X"01",X"01",X"00",X"00",X"03",X"80",X"E0",X"84",X"E0",X"78",X"52",X"00",
		X"C1",X"2C",X"20",X"00",X"08",X"C5",X"B5",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"33",X"44",X"03",X"8C",X"07",X"07",X"30",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"88",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"21",X"10",X"00",X"00",X"00",X"00",X"00",X"C3",X"1E",X"F0",X"C3",X"C3",X"34",X"03",X"00",
		X"1E",X"80",X"00",X"00",X"38",X"F0",X"0F",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"01",X"11",X"00",X"00",X"00",X"01",X"11",X"66",X"88",X"00",X"42",X"A4",X"43",X"1C",
		X"CC",X"33",X"00",X"00",X"00",X"02",X"60",X"C0",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",
		X"02",X"70",X"70",X"30",X"00",X"00",X"00",X"00",X"21",X"86",X"80",X"21",X"34",X"16",X"00",X"00",
		X"08",X"00",X"08",X"78",X"F0",X"C3",X"0C",X"00",X"00",X"00",X"60",X"C0",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"32",X"64",X"61",X"50",X"00",X"64",X"C8",X"80",X"80",X"08",X"88",X"1A",
		X"00",X"00",X"00",X"00",X"23",X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",
		X"41",X"02",X"00",X"10",X"30",X"30",X"00",X"00",X"34",X"4B",X"86",X"85",X"D2",X"3C",X"01",X"00",
		X"80",X"00",X"80",X"86",X"3C",X"E1",X"0E",X"00",X"60",X"E0",X"E0",X"C0",X"08",X"00",X"00",X"00",
		X"00",X"00",X"11",X"32",X"32",X"74",X"60",X"61",X"00",X"40",X"C8",X"84",X"80",X"00",X"00",X"1E",
		X"00",X"00",X"00",X"22",X"08",X"04",X"C2",X"80",X"00",X"00",X"00",X"00",X"22",X"22",X"31",X"60",
		X"21",X"12",X"01",X"00",X"00",X"00",X"00",X"00",X"90",X"10",X"30",X"C3",X"D2",X"70",X"60",X"00",
		X"C4",X"80",X"A0",X"21",X"30",X"86",X"00",X"00",X"60",X"60",X"60",X"C0",X"80",X"00",X"00",X"00",
		X"00",X"00",X"11",X"32",X"74",X"74",X"60",X"60",X"00",X"00",X"11",X"00",X"00",X"10",X"10",X"32",
		X"00",X"00",X"88",X"00",X"00",X"80",X"80",X"C4",X"00",X"00",X"88",X"C4",X"E2",X"E2",X"60",X"60",
		X"70",X"61",X"12",X"01",X"00",X"00",X"00",X"00",X"D4",X"90",X"81",X"29",X"21",X"10",X"10",X"00",
		X"B2",X"90",X"18",X"49",X"48",X"80",X"80",X"00",X"E0",X"68",X"84",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"21",X"21",X"00",X"00",X"00",X"00",X"00",X"C0",X"C8",X"D9",
		X"00",X"00",X"00",X"00",X"00",X"30",X"31",X"B9",X"00",X"00",X"00",X"00",X"00",X"80",X"48",X"48",
		X"21",X"21",X"03",X"74",X"30",X"10",X"00",X"00",X"FA",X"CA",X"7F",X"FD",X"FC",X"FC",X"21",X"00",
		X"7D",X"B5",X"67",X"73",X"F3",X"F3",X"48",X"00",X"48",X"48",X"0C",X"E2",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"22",X"00",X"30",X"71",X"00",X"11",X"00",X"00",X"00",X"13",X"3F",X"92",
		X"00",X"88",X"CC",X"F0",X"7A",X"FA",X"7D",X"F5",X"00",X"00",X"00",X"88",X"C4",X"E2",X"E2",X"C0",
		X"61",X"61",X"30",X"10",X"22",X"00",X"00",X"00",X"9E",X"FB",X"3A",X"A2",X"F3",X"E0",X"00",X"00",
		X"06",X"C9",X"21",X"F0",X"4A",X"84",X"00",X"00",X"E0",X"E8",X"48",X"08",X"88",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"70",X"20",X"10",X"01",X"33",X"1F",
		X"00",X"00",X"91",X"00",X"04",X"82",X"49",X"87",X"00",X"00",X"88",X"CC",X"66",X"22",X"20",X"E8",
		X"30",X"30",X"30",X"10",X"32",X"11",X"00",X"00",X"96",X"69",X"2C",X"86",X"C2",X"F0",X"F8",X"00",
		X"C1",X"B8",X"7C",X"34",X"12",X"01",X"80",X"00",X"2C",X"0C",X"86",X"C0",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"A1",X"34",X"22",X"77",X"36",
		X"00",X"66",X"91",X"E0",X"3C",X"E1",X"CF",X"F0",X"00",X"00",X"88",X"80",X"C0",X"C8",X"0C",X"8E",
		X"01",X"12",X"10",X"01",X"10",X"00",X"00",X"00",X"1E",X"87",X"2D",X"C3",X"F0",X"30",X"10",X"00",
		X"98",X"DC",X"16",X"01",X"80",X"E0",X"C0",X"00",X"E2",X"C0",X"80",X"80",X"88",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"11",X"00",X"00",X"83",X"38",X"33",X"33",
		X"00",X"FF",X"10",X"10",X"2F",X"C3",X"DC",X"48",X"00",X"00",X"80",X"C0",X"0C",X"0E",X"E0",X"E0",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"33",X"03",X"78",X"4B",X"43",X"30",X"10",X"00",
		X"B3",X"0D",X"F3",X"3D",X"3C",X"F0",X"E0",X"00",X"E0",X"2C",X"EE",X"CC",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"10",X"12",X"52",X"00",X"10",X"70",X"F0",X"C2",X"DE",X"3F",X"FE",
		X"00",X"C0",X"E0",X"87",X"AE",X"38",X"F8",X"76",X"00",X"00",X"00",X"08",X"80",X"80",X"C0",X"6A",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"56",X"07",X"02",X"43",X"2D",X"25",X"10",X"00",
		X"21",X"3F",X"3D",X"BC",X"3C",X"F0",X"C0",X"00",X"66",X"CC",X"C8",X"C0",X"80",X"00",X"00",X"00",
		X"00",X"00",X"11",X"33",X"22",X"10",X"30",X"30",X"00",X"FC",X"B8",X"60",X"D3",X"B5",X"2D",X"3E",
		X"00",X"A2",X"EE",X"FC",X"F8",X"F0",X"A3",X"46",X"00",X"00",X"00",X"00",X"80",X"08",X"00",X"20",
		X"12",X"03",X"02",X"00",X"00",X"00",X"00",X"00",X"7F",X"23",X"01",X"10",X"12",X"07",X"00",X"00",
		X"84",X"69",X"C3",X"96",X"B4",X"E0",X"00",X"00",X"60",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"32",X"32",X"54",X"74",X"30",X"00",X"11",X"F3",X"E6",X"A3",X"E2",X"FA",X"EA",
		X"00",X"88",X"C0",X"E0",X"61",X"93",X"55",X"BF",X"00",X"00",X"00",X"08",X"88",X"C8",X"E8",X"E0",
		X"31",X"30",X"03",X"01",X"01",X"00",X"00",X"00",X"7A",X"F7",X"93",X"00",X"00",X"00",X"01",X"00",
		X"84",X"1F",X"3E",X"3E",X"F0",X"0C",X"08",X"00",X"C0",X"C0",X"E2",X"C4",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"30",X"74",X"30",X"21",X"21",X"00",X"74",X"FC",X"FC",X"CE",X"D5",X"6A",X"58",
		X"00",X"E2",X"F3",X"F3",X"37",X"BA",X"65",X"A1",X"00",X"00",X"80",X"C0",X"E2",X"C0",X"48",X"48",
		X"21",X"21",X"10",X"00",X"00",X"00",X"00",X"00",X"48",X"48",X"C0",X"0C",X"04",X"00",X"00",X"00",
		X"21",X"21",X"30",X"03",X"02",X"00",X"00",X"00",X"48",X"48",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"30",X"30",X"54",X"30",X"00",X"22",X"19",X"60",X"F8",X"B8",X"F4",X"21",
		X"00",X"44",X"89",X"60",X"F1",X"D1",X"F2",X"48",X"00",X"00",X"00",X"80",X"C0",X"40",X"A2",X"C0",
		X"70",X"70",X"60",X"60",X"04",X"40",X"00",X"00",X"47",X"66",X"00",X"42",X"00",X"00",X"00",X"00",
		X"2E",X"66",X"00",X"24",X"00",X"00",X"00",X"00",X"E0",X"E0",X"60",X"60",X"02",X"20",X"00",X"00",
		X"00",X"00",X"10",X"12",X"00",X"71",X"71",X"70",X"00",X"B8",X"F4",X"F0",X"F0",X"F0",X"C3",X"8D",
		X"44",X"32",X"F6",X"D4",X"D4",X"0C",X"06",X"4C",X"00",X"00",X"80",X"C4",X"C0",X"E0",X"E0",X"60",
		X"70",X"70",X"70",X"30",X"12",X"01",X"01",X"00",X"0E",X"4C",X"12",X"22",X"00",X"00",X"00",X"00",
		X"20",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"30",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"00",X"55",X"78",X"B8",X"54",X"D1",X"7E",X"12",X"F3",X"E1",X"F1",X"E0",X"5B",X"63",
		X"C0",X"D1",X"F0",X"30",X"DC",X"0C",X"08",X"60",X"00",X"00",X"88",X"C4",X"E2",X"71",X"10",X"00",
		X"F0",X"70",X"70",X"30",X"01",X"00",X"00",X"00",X"CE",X"84",X"B0",X"90",X"80",X"48",X"04",X"20",
		X"31",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"22",X"10",X"70",X"10",X"74",X"F0",X"00",X"70",X"7C",X"26",X"D3",X"E1",X"E0",X"D1",
		X"00",X"E0",X"F0",X"70",X"8C",X"EE",X"48",X"64",X"00",X"00",X"80",X"E0",X"00",X"00",X"00",X"00",
		X"30",X"88",X"70",X"70",X"30",X"00",X"00",X"00",X"0D",X"67",X"92",X"C0",X"E0",X"F0",X"30",X"00",
		X"00",X"00",X"80",X"C0",X"00",X"00",X"C0",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"32",X"10",X"74",X"50",X"00",X"10",X"F0",X"B0",X"3F",X"C3",X"E0",X"E0",
		X"00",X"F0",X"F0",X"C0",X"00",X"7F",X"7C",X"08",X"00",X"C0",X"88",X"00",X"00",X"00",X"00",X"00",
		X"76",X"30",X"10",X"32",X"10",X"00",X"00",X"00",X"E0",X"C2",X"2E",X"B8",X"F0",X"F0",X"10",X"00",
		X"08",X"08",X"38",X"00",X"C0",X"E0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"C0",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
