library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity GFX1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of GFX1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"CC",X"FF",X"FF",X"00",X"00",X"00",X"00",X"EE",X"FF",X"FF",X"FF",
		X"CC",X"EE",X"EE",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"77",X"22",X"88",X"CC",X"FF",X"FF",X"77",X"11",X"CC",X"FF",X"FF",X"FF",
		X"88",X"CC",X"EE",X"EE",X"EE",X"EE",X"CC",X"88",X"33",X"77",X"DF",X"BF",X"BF",X"FF",X"77",X"33",
		X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"33",X"67",X"CF",X"9F",X"FF",X"FF",X"77",X"33",
		X"22",X"88",X"CC",X"CC",X"EE",X"EE",X"FF",X"FF",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"77",X"33",X"11",X"11",X"00",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"3F",X"7F",X"FF",X"FF",X"EE",X"FF",X"FF",X"FF",X"33",X"33",X"33",X"77",X"77",X"77",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"EE",X"CC",X"00",X"CC",X"FF",X"FF",X"FF",X"FF",X"77",X"00",X"EE",X"FF",
		X"00",X"00",X"00",X"00",X"88",X"FF",X"9F",X"3F",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"11",
		X"00",X"88",X"CC",X"EE",X"EE",X"FF",X"FF",X"FF",X"00",X"FF",X"33",X"11",X"11",X"FF",X"3F",X"FF",
		X"CC",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"BF",X"BF",X"FF",X"77",X"77",X"33",X"11",X"00",
		X"FF",X"FF",X"FF",X"EE",X"EE",X"CC",X"88",X"00",X"33",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CC",X"CC",X"FF",X"FF",X"FF",X"FF",X"77",X"77",X"DF",X"DF",
		X"88",X"EE",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"33",
		X"FF",X"FF",X"FF",X"FF",X"EE",X"EE",X"CC",X"00",X"FF",X"FF",X"FF",X"FF",X"77",X"77",X"33",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"23",X"47",X"57",X"57",X"9F",X"BF",X"BF",X"FF",
		X"00",X"00",X"00",X"00",X"33",X"FF",X"9F",X"BF",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",
		X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"33",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"77",X"77",X"33",X"BB",X"99",X"DD",X"CC",X"EE",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"88",X"FF",X"FF",X"00",X"00",X"88",X"88",X"CC",X"DD",X"CC",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",
		X"11",X"33",X"77",X"77",X"77",X"33",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"FF",
		X"FF",X"FF",X"FF",X"33",X"11",X"11",X"11",X"00",X"FF",X"FF",X"FF",X"CC",X"88",X"88",X"88",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"BF",X"7F",X"FF",X"FF",
		X"FF",X"FF",X"77",X"00",X"00",X"00",X"00",X"00",X"FF",X"33",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"33",X"88",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"88",X"88",X"CC",X"CC",X"EE",X"EE",X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",
		X"00",X"00",X"00",X"00",X"33",X"67",X"47",X"DF",X"00",X"00",X"00",X"00",X"CC",X"EE",X"EE",X"EE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"33",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"11",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"BB",X"BB",X"00",X"00",X"00",X"00",X"00",X"66",X"FF",X"FF",X"66",X"00",X"00",
		X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"33",X"CC",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"FF",X"FF",X"FF",X"FF",
		X"99",X"55",X"55",X"33",X"88",X"44",X"22",X"11",X"88",X"55",X"33",X"11",X"00",X"FF",X"88",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"33",X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CC",X"FF",X"FF",X"FF",
		X"FF",X"CC",X"77",X"FF",X"CC",X"77",X"FF",X"FF",X"FF",X"FF",X"EE",X"BB",X"FF",X"EE",X"DD",X"FF",
		X"FF",X"FF",X"44",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"33",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"BB",X"FF",X"EE",X"EE",X"77",X"BB",X"FF",X"FF",X"FF",X"FF",X"33",X"CC",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"11",X"FF",X"FF",
		X"00",X"00",X"EE",X"DD",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"8D",X"8A",X"8D",X"8A",X"8D",X"8A",X"8D",X"8A",
		X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"DD",X"DD",X"00",X"00",X"00",
		X"88",X"CC",X"22",X"22",X"66",X"CC",X"88",X"00",X"33",X"77",X"CC",X"88",X"88",X"77",X"33",X"00",
		X"22",X"22",X"EE",X"EE",X"22",X"22",X"00",X"00",X"00",X"00",X"FF",X"FF",X"44",X"00",X"00",X"00",
		X"22",X"22",X"AA",X"AA",X"EE",X"EE",X"66",X"00",X"66",X"FF",X"BB",X"99",X"99",X"CC",X"44",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"88",X"DD",X"FF",X"BB",X"99",X"88",X"00",X"00",
		X"88",X"EE",X"EE",X"88",X"88",X"88",X"88",X"00",X"00",X"FF",X"FF",X"CC",X"66",X"33",X"11",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"11",X"BB",X"AA",X"AA",X"AA",X"EE",X"EE",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",X"00",X"99",X"99",X"99",X"DD",X"77",X"33",X"00",
		X"00",X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"CC",X"EE",X"BB",X"99",X"88",X"CC",X"CC",X"00",
		X"CC",X"EE",X"AA",X"AA",X"22",X"22",X"CC",X"00",X"00",X"66",X"99",X"99",X"BB",X"FF",X"66",X"00",
		X"88",X"CC",X"66",X"22",X"22",X"22",X"00",X"00",X"77",X"FF",X"99",X"99",X"99",X"FF",X"66",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"33",X"FF",
		X"77",X"99",X"EE",X"FF",X"77",X"FF",X"FF",X"FF",X"FF",X"77",X"BB",X"CC",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"66",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",
		X"C0",X"C8",X"D5",X"FF",X"FF",X"D9",X"C0",X"80",X"30",X"71",X"F0",X"F3",X"F4",X"F0",X"71",X"30",
		X"CC",X"22",X"11",X"55",X"55",X"99",X"22",X"CC",X"33",X"44",X"88",X"AA",X"AA",X"99",X"44",X"33",
		X"EE",X"EE",X"88",X"88",X"88",X"EE",X"EE",X"00",X"33",X"77",X"CC",X"88",X"CC",X"77",X"33",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"EE",X"00",X"66",X"FF",X"99",X"99",X"99",X"FF",X"FF",X"00",
		X"44",X"66",X"22",X"22",X"66",X"CC",X"88",X"00",X"44",X"CC",X"88",X"88",X"CC",X"77",X"33",X"00",
		X"88",X"CC",X"66",X"22",X"22",X"EE",X"EE",X"00",X"33",X"77",X"CC",X"88",X"88",X"FF",X"FF",X"00",
		X"22",X"22",X"22",X"22",X"EE",X"EE",X"00",X"00",X"88",X"99",X"99",X"99",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"00",X"88",X"99",X"99",X"99",X"99",X"FF",X"FF",X"00",
		X"EE",X"EE",X"22",X"22",X"66",X"CC",X"88",X"00",X"99",X"99",X"99",X"88",X"CC",X"77",X"33",X"00",
		X"EE",X"EE",X"00",X"00",X"00",X"EE",X"EE",X"00",X"FF",X"FF",X"11",X"11",X"11",X"FF",X"FF",X"00",
		X"22",X"22",X"EE",X"EE",X"22",X"22",X"00",X"00",X"88",X"88",X"FF",X"FF",X"88",X"88",X"00",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"66",X"EE",X"CC",X"88",X"EE",X"EE",X"00",X"88",X"CC",X"66",X"33",X"11",X"FF",X"FF",X"00",
		X"22",X"22",X"22",X"22",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"EE",X"EE",X"00",X"88",X"00",X"EE",X"EE",X"00",X"FF",X"FF",X"77",X"33",X"77",X"FF",X"FF",X"00",
		X"EE",X"EE",X"CC",X"88",X"00",X"EE",X"EE",X"00",X"FF",X"FF",X"11",X"33",X"77",X"FF",X"FF",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",X"77",X"FF",X"88",X"88",X"88",X"FF",X"77",X"00",
		X"00",X"88",X"88",X"88",X"88",X"EE",X"EE",X"00",X"77",X"FF",X"88",X"88",X"88",X"FF",X"FF",X"00",
		X"AA",X"CC",X"EE",X"AA",X"22",X"EE",X"CC",X"00",X"77",X"FF",X"88",X"88",X"88",X"FF",X"77",X"00",
		X"22",X"66",X"EE",X"CC",X"88",X"EE",X"EE",X"00",X"77",X"FF",X"99",X"88",X"88",X"FF",X"FF",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"00",X"55",X"DD",X"99",X"99",X"FF",X"66",X"00",
		X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"00",X"88",X"88",X"FF",X"FF",X"88",X"88",X"00",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"88",X"CC",X"EE",X"CC",X"88",X"00",X"00",X"FF",X"FF",X"11",X"00",X"11",X"FF",X"FF",X"00",
		X"EE",X"EE",X"CC",X"88",X"CC",X"EE",X"EE",X"00",X"FF",X"FF",X"11",X"33",X"11",X"FF",X"FF",X"00",
		X"66",X"EE",X"CC",X"88",X"CC",X"EE",X"66",X"00",X"CC",X"EE",X"77",X"33",X"77",X"EE",X"CC",X"00",
		X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"00",X"EE",X"FF",X"11",X"11",X"FF",X"EE",X"00",X"00",
		X"22",X"22",X"22",X"AA",X"EE",X"EE",X"66",X"00",X"CC",X"EE",X"FF",X"BB",X"99",X"88",X"88",X"00",
		X"77",X"DD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"88",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CC",X"FF",X"00",X"FF",X"FF",X"FF",
		X"EE",X"11",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"88",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"DD",X"BB",X"FF",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"CC",X"FF",X"FF",X"FF",
		X"01",X"03",X"05",X"0E",X"05",X"0A",X"05",X"0A",X"88",X"88",X"88",X"88",X"89",X"8B",X"8D",X"8E",
		X"00",X"00",X"00",X"0C",X"1F",X"3F",X"7F",X"FF",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"1F",X"3F",X"7F",X"FF",X"00",X"00",X"00",X"00",X"03",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"CC",X"CC",X"EE",X"6E",X"04",X"04",X"06",X"3F",X"FF",X"FF",X"FF",X"CF",
		X"00",X"00",X"00",X"00",X"CC",X"CC",X"EE",X"6E",X"01",X"03",X"06",X"3F",X"FF",X"FF",X"FF",X"CF",
		X"6E",X"EE",X"EE",X"EE",X"EE",X"CC",X"88",X"08",X"8F",X"0F",X"0F",X"0F",X"8F",X"8F",X"CF",X"01",
		X"6E",X"EE",X"EE",X"EE",X"EE",X"CC",X"88",X"00",X"8F",X"0F",X"0F",X"0F",X"1F",X"3F",X"7F",X"00",
		X"DD",X"FF",X"FF",X"77",X"33",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DD",X"FF",X"EF",X"67",X"23",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"11",X"33",X"77",X"FF",X"FF",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"23",X"67",X"EF",X"FF",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"88",X"CC",X"EE",X"EE",X"EE",X"EE",X"6E",X"01",X"CF",X"8F",X"8F",X"0F",X"0F",X"0F",X"8F",
		X"00",X"88",X"CC",X"EE",X"EE",X"EE",X"EE",X"6E",X"00",X"7F",X"3F",X"1F",X"0F",X"0F",X"0F",X"8F",
		X"6E",X"EE",X"CC",X"CC",X"00",X"00",X"00",X"00",X"CF",X"FF",X"FF",X"FF",X"3F",X"06",X"04",X"04",
		X"6E",X"EE",X"CC",X"CC",X"00",X"00",X"00",X"00",X"CF",X"FF",X"FF",X"FF",X"3F",X"06",X"03",X"01",
		X"FF",X"7F",X"3F",X"1F",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",
		X"FF",X"7F",X"3F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"00",X"00",
		X"80",X"C0",X"C0",X"C0",X"C0",X"80",X"A6",X"84",X"76",X"54",X"F0",X"F0",X"D4",X"F6",X"F0",X"78",
		X"C0",X"E0",X"E0",X"E0",X"E0",X"C0",X"D3",X"86",X"00",X"30",X"76",X"54",X"70",X"70",X"54",X"76",
		X"1F",X"0E",X"0E",X"0E",X"0F",X"0F",X"0F",X"06",X"0F",X"07",X"07",X"07",X"03",X"03",X"01",X"00",
		X"1F",X"0F",X"0F",X"0E",X"0E",X"0E",X"0C",X"08",X"01",X"01",X"01",X"03",X"07",X"0F",X"0F",X"07",
		X"06",X"0F",X"0F",X"0F",X"0E",X"0E",X"0E",X"1F",X"00",X"01",X"03",X"03",X"07",X"07",X"07",X"0F",
		X"08",X"0C",X"0E",X"0E",X"0E",X"0F",X"0F",X"1F",X"07",X"0F",X"0F",X"07",X"03",X"01",X"01",X"01",
		X"84",X"A6",X"80",X"C0",X"C0",X"C0",X"C0",X"80",X"78",X"F0",X"F6",X"D4",X"F0",X"F0",X"54",X"76",
		X"86",X"D3",X"C0",X"E0",X"E0",X"E0",X"E0",X"C0",X"76",X"54",X"70",X"70",X"54",X"76",X"30",X"00",
		X"F0",X"98",X"AE",X"8E",X"9F",X"8E",X"8E",X"06",X"31",X"22",X"EE",X"E2",X"22",X"22",X"EE",X"F1",
		X"F0",X"98",X"AE",X"8E",X"9F",X"8E",X"8E",X"06",X"F1",X"EE",X"22",X"22",X"E2",X"EE",X"22",X"31",
		X"06",X"06",X"1F",X"0E",X"3A",X"F8",X"70",X"F0",X"F0",X"F0",X"E0",X"C1",X"83",X"83",X"83",X"C0",
		X"06",X"06",X"06",X"0E",X"0E",X"1C",X"7C",X"70",X"F0",X"F0",X"90",X"06",X"07",X"8F",X"07",X"A2",
		X"F0",X"70",X"F8",X"3A",X"0E",X"1F",X"06",X"06",X"C0",X"83",X"83",X"83",X"C1",X"E0",X"F0",X"F0",
		X"70",X"7C",X"1C",X"0E",X"0E",X"06",X"06",X"06",X"A2",X"07",X"8F",X"07",X"06",X"90",X"F0",X"F0",
		X"06",X"8E",X"8E",X"9F",X"8E",X"AE",X"98",X"F0",X"F1",X"EE",X"22",X"22",X"E2",X"EE",X"22",X"31",
		X"06",X"8E",X"8E",X"9F",X"8E",X"AE",X"98",X"F0",X"31",X"22",X"EE",X"E2",X"22",X"22",X"EE",X"F1",
		X"10",X"0E",X"0F",X"0F",X"8F",X"A2",X"F0",X"F0",X"C0",X"83",X"07",X"07",X"06",X"32",X"F0",X"F0",
		X"F0",X"F0",X"A2",X"8F",X"0F",X"0F",X"0E",X"10",X"F0",X"F0",X"32",X"06",X"07",X"07",X"83",X"C0",
		X"72",X"55",X"DD",X"D5",X"55",X"55",X"DD",X"72",X"E0",X"E0",X"75",X"1C",X"0E",X"0E",X"17",X"80",
		X"72",X"DD",X"55",X"55",X"D5",X"DD",X"55",X"72",X"80",X"17",X"0E",X"0E",X"1C",X"75",X"E0",X"E0",
		X"22",X"88",X"44",X"88",X"22",X"88",X"44",X"88",X"DD",X"EE",X"BB",X"EE",X"DD",X"EE",X"BB",X"EE",
		X"00",X"00",X"00",X"00",X"08",X"0C",X"06",X"0B",X"08",X"0C",X"06",X"0B",X"05",X"0A",X"05",X"0A",
		X"07",X"0A",X"0C",X"08",X"00",X"00",X"00",X"00",X"05",X"0A",X"05",X"0A",X"07",X"0A",X"0C",X"08",
		X"07",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"0A",X"07",X"0C",X"08",X"0C",X"06",X"0B",
		X"00",X"00",X"00",X"00",X"01",X"13",X"37",X"36",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"1F",X"93",X"93",X"D3",X"80",X"00",X"00",X"00",X"00",X"03",X"17",X"9B",X"9B",X"CA",X"80",
		X"80",X"C4",X"0A",X"D6",X"32",X"FC",X"B6",X"7C",X"93",X"82",X"93",X"C7",X"39",X"57",X"33",X"03",
		X"B4",X"B2",X"54",X"BE",X"7A",X"54",X"FA",X"BA",X"37",X"13",X"56",X"36",X"33",X"57",X"32",X"32",
		X"7C",X"B6",X"FC",X"32",X"D6",X"0A",X"C4",X"80",X"03",X"33",X"57",X"39",X"C7",X"93",X"82",X"93",
		X"00",X"00",X"80",X"D3",X"93",X"93",X"1F",X"03",X"80",X"CA",X"9B",X"9B",X"17",X"03",X"00",X"00",
		X"36",X"37",X"13",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DD",X"EA",X"55",X"6A",X"BE",X"5C",X"3A",X"37",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"17",X"3F",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"0C",X"8E",X"CE",X"CE",X"CE",X"00",X"00",X"07",X"3F",X"FF",X"FF",X"FF",X"FF",
		X"CE",X"CE",X"CE",X"8E",X"0C",X"08",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"3F",X"07",X"00",X"00",
		X"3F",X"3F",X"17",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"0A",X"05",X"0A",X"85",X"C2",X"E1",X"F0",X"05",X"0A",X"05",X"0A",X"14",X"38",X"70",X"F0",
		X"F0",X"E0",X"C1",X"82",X"05",X"0A",X"05",X"0A",X"F0",X"78",X"34",X"1A",X"05",X"0A",X"05",X"0A",
		X"14",X"1A",X"34",X"38",X"34",X"78",X"70",X"78",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"0A",
		X"70",X"78",X"70",X"38",X"34",X"38",X"14",X"1A",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"0A",
		X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"85",X"82",X"C1",X"C2",X"C1",X"E0",X"E1",X"E0",
		X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"E1",X"E0",X"E1",X"C2",X"C1",X"C2",X"85",X"82",
		X"14",X"38",X"70",X"F0",X"F0",X"78",X"34",X"1A",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"0A",
		X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"85",X"C2",X"E1",X"F0",X"F0",X"E0",X"C1",X"82",
		X"05",X"0A",X"05",X"0A",X"05",X"78",X"F0",X"F0",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"34",X"F0",
		X"05",X"0A",X"05",X"0A",X"05",X"0A",X"C1",X"F0",X"05",X"0A",X"05",X"0A",X"05",X"E0",X"F0",X"F0",
		X"F0",X"F0",X"70",X"0A",X"05",X"0A",X"05",X"0A",X"F0",X"38",X"05",X"0A",X"05",X"0A",X"05",X"0A",
		X"F0",X"C2",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"F0",X"F0",X"E1",X"0A",X"05",X"0A",X"05",X"0A",
		X"05",X"1B",X"37",X"7F",X"77",X"FF",X"FF",X"FF",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"37",X"7F",
		X"FF",X"CC",X"33",X"FF",X"EF",X"8A",X"05",X"0A",X"FF",X"FF",X"FF",X"DD",X"BB",X"FF",X"EF",X"8A",
		X"EF",X"8A",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"11",X"FF",X"EF",X"8A",X"05",X"0A",X"05",X"0A",
		X"15",X"1B",X"37",X"B3",X"F7",X"7F",X"FF",X"FF",X"85",X"C2",X"F0",X"F0",X"F0",X"F0",X"C1",X"82",
		X"EF",X"CE",X"8D",X"82",X"C1",X"C2",X"E1",X"F0",X"FF",X"FF",X"DD",X"BB",X"76",X"FC",X"F8",X"F0",
		X"FE",X"DC",X"BC",X"38",X"34",X"78",X"70",X"78",X"15",X"1B",X"37",X"3B",X"67",X"4E",X"8D",X"0A",
		X"05",X"0A",X"8D",X"EE",X"77",X"99",X"EE",X"FF",X"8D",X"EE",X"BB",X"DD",X"EE",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"77",X"F7",X"B7",X"3B",X"15",X"1B",X"85",X"C2",X"F0",X"F0",X"F0",X"F0",X"C1",X"82",
		X"F0",X"E0",X"C1",X"C2",X"85",X"8A",X"CD",X"EE",X"F0",X"F8",X"FC",X"76",X"BB",X"DD",X"FF",X"FF",
		X"77",X"BB",X"FF",X"EE",X"77",X"3B",X"15",X"0A",X"77",X"3B",X"15",X"0A",X"05",X"0A",X"05",X"0A",
		X"05",X"0A",X"05",X"0A",X"05",X"0A",X"8D",X"EE",X"05",X"0A",X"05",X"0A",X"8D",X"EE",X"77",X"11",
		X"05",X"0A",X"05",X"0A",X"0D",X"06",X"03",X"01",X"0D",X"06",X"03",X"01",X"00",X"00",X"00",X"00",
		X"C7",X"1F",X"93",X"93",X"13",X"00",X"00",X"00",X"CF",X"E4",X"E7",X"97",X"0A",X"00",X"00",X"00",
		X"00",X"00",X"00",X"13",X"93",X"93",X"1F",X"C7",X"00",X"00",X"00",X"0A",X"97",X"E7",X"E4",X"CF",
		X"93",X"82",X"93",X"82",X"D9",X"E8",X"D9",X"E8",X"11",X"11",X"11",X"11",X"01",X"01",X"01",X"01",
		X"37",X"3A",X"5C",X"BE",X"6A",X"55",X"EA",X"DD",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"15",X"1B",X"37",X"3B",X"77",X"7F",X"FF",X"FF",
		X"FE",X"DC",X"BC",X"38",X"34",X"78",X"70",X"78",X"FF",X"FF",X"FF",X"FF",X"EF",X"CE",X"8D",X"0A",
		X"15",X"1B",X"37",X"3B",X"77",X"7F",X"FF",X"FF",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"0A",
		X"FE",X"FE",X"FC",X"FC",X"BC",X"F8",X"70",X"78",X"15",X"1B",X"37",X"3B",X"77",X"7F",X"FF",X"FF",
		X"70",X"78",X"70",X"38",X"34",X"38",X"14",X"1A",X"EF",X"EE",X"CD",X"CE",X"8D",X"8A",X"05",X"0A",
		X"EF",X"EE",X"CD",X"CE",X"8D",X"8A",X"05",X"0A",X"15",X"1B",X"37",X"3B",X"77",X"7F",X"FF",X"FF",
		X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"EF",X"EE",X"CD",X"CE",X"8D",X"8A",X"05",X"0A",
		X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"8D",X"8A",X"CD",X"CE",X"EF",X"EE",
		X"05",X"0A",X"8D",X"8A",X"CD",X"CE",X"EF",X"EE",X"FF",X"FF",X"77",X"7F",X"37",X"3B",X"15",X"1B",
		X"FF",X"FF",X"77",X"7F",X"37",X"3B",X"15",X"1B",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"0A",
		X"05",X"0A",X"05",X"0A",X"05",X"8A",X"CD",X"EE",X"05",X"8A",X"CD",X"EE",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"7F",X"37",X"3B",X"15",X"1B",
		X"70",X"78",X"70",X"38",X"34",X"B8",X"DC",X"FE",X"05",X"8A",X"CD",X"66",X"BB",X"DD",X"FF",X"FF",
		X"14",X"1A",X"34",X"38",X"34",X"78",X"70",X"78",X"05",X"0A",X"8D",X"8A",X"CD",X"CE",X"EF",X"EE",
		X"70",X"78",X"F8",X"B8",X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",X"77",X"7F",X"37",X"3B",X"15",X"1B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"F0",X"00",X"00",X"00",X"00",X"10",X"30",X"70",X"F0",
		X"F0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"F0",X"70",X"30",X"10",X"00",X"00",X"00",X"00",
		X"10",X"10",X"30",X"30",X"30",X"70",X"70",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"70",X"70",X"30",X"30",X"30",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"C0",X"E0",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"80",X"80",
		X"10",X"30",X"70",X"F0",X"F0",X"70",X"30",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"07",X"0F",X"0F",X"07",X"03",X"01",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"00",X"00",X"00",X"00",X"00",X"70",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"F0",X"00",X"00",X"00",X"00",X"00",X"E0",X"F0",X"F0",
		X"F0",X"F0",X"70",X"00",X"00",X"00",X"00",X"00",X"F0",X"30",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"8F",X"CF",X"EF",X"0F",X"8F",X"CF",X"EF",X"FF",X"FF",X"FF",X"FF",
		X"11",X"33",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"11",X"33",X"77",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"33",X"11",X"FF",X"77",X"33",X"11",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"11",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"33",X"11",X"FF",X"FF",X"FF",X"77",X"11",X"00",X"00",X"00",
		X"CC",X"EE",X"FF",X"FF",X"FF",X"66",X"33",X"11",X"FF",X"77",X"33",X"11",X"00",X"00",X"00",X"00",
		X"77",X"DD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"88",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"11",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",
		X"11",X"33",X"77",X"EE",X"DD",X"BB",X"FF",X"FF",X"00",X"00",X"00",X"11",X"77",X"FF",X"FF",X"FF",
		X"11",X"33",X"77",X"FF",X"FF",X"FF",X"BB",X"77",X"00",X"00",X"00",X"00",X"11",X"33",X"77",X"FF",
		X"FF",X"FF",X"77",X"CC",X"FF",X"77",X"CC",X"FF",X"FF",X"DD",X"EE",X"FF",X"BB",X"EE",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"44",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"33",X"FF",
		X"FF",X"BB",X"77",X"EE",X"EE",X"FF",X"BB",X"FF",X"FF",X"FF",X"FF",X"CC",X"33",X"FF",X"FF",X"FF",
		X"14",X"38",X"F0",X"F0",X"F0",X"F0",X"34",X"1A",X"8D",X"8A",X"CD",X"56",X"76",X"66",X"77",X"33",
		X"05",X"8A",X"8D",X"CE",X"CD",X"66",X"67",X"BB",X"BB",X"DD",X"DD",X"EE",X"66",X"BB",X"FF",X"FF",
		X"FF",X"FF",X"EE",X"FF",X"F7",X"F3",X"F1",X"F0",X"77",X"3B",X"15",X"1A",X"34",X"38",X"70",X"F0",
		X"14",X"38",X"F0",X"F0",X"F0",X"F8",X"FC",X"FE",X"05",X"8A",X"CD",X"76",X"BB",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"3B",X"05",X"0A",X"05",X"0A",X"F7",X"B3",X"C1",X"C2",X"C1",X"E0",X"E1",X"E0",
		X"F0",X"F0",X"70",X"0A",X"05",X"8A",X"CD",X"2A",X"F0",X"B8",X"CD",X"EE",X"FF",X"3B",X"05",X"0A",
		X"EE",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"FF",X"EE",X"88",X"00",X"00",X"00",X"00",
		X"FF",X"CC",X"33",X"FF",X"EE",X"88",X"00",X"00",X"FF",X"FF",X"FF",X"DD",X"BB",X"FF",X"EE",X"88",
		X"11",X"33",X"77",X"FF",X"77",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"11",X"22",X"77",X"FF",
		X"EE",X"CC",X"88",X"80",X"C0",X"C0",X"E0",X"F0",X"FF",X"FF",X"DD",X"BB",X"76",X"FC",X"F8",X"F0",
		X"11",X"11",X"33",X"B3",X"F7",X"77",X"FF",X"FF",X"80",X"C0",X"F0",X"F0",X"F0",X"F0",X"C0",X"80",
		X"FE",X"DC",X"B8",X"30",X"30",X"70",X"70",X"70",X"11",X"11",X"33",X"33",X"66",X"44",X"88",X"00",
		X"70",X"70",X"70",X"30",X"30",X"B8",X"DC",X"FE",X"00",X"88",X"44",X"66",X"33",X"33",X"11",X"11",
		X"FF",X"FF",X"77",X"F7",X"B3",X"33",X"11",X"11",X"80",X"C0",X"F0",X"F0",X"F0",X"F0",X"C0",X"80",
		X"F0",X"E0",X"C0",X"C0",X"80",X"88",X"CC",X"EE",X"F0",X"F8",X"FC",X"76",X"BB",X"DD",X"FF",X"FF",
		X"77",X"BB",X"FF",X"EE",X"FF",X"77",X"33",X"11",X"FF",X"77",X"33",X"11",X"00",X"00",X"00",X"00",
		X"00",X"00",X"88",X"EE",X"77",X"99",X"EE",X"FF",X"88",X"EE",X"BB",X"DD",X"EE",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"EE",X"00",X"00",X"00",X"00",X"88",X"EE",X"77",X"11",
		X"00",X"00",X"00",X"00",X"88",X"EE",X"FF",X"FF",X"88",X"88",X"CC",X"66",X"77",X"33",X"99",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"FF",
		X"99",X"77",X"FF",X"CC",X"00",X"00",X"00",X"00",X"FF",X"FF",X"AA",X"77",X"77",X"EE",X"CC",X"88",
		X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"88",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"88",X"FF",X"BF",X"FF",X"FF",X"FF",X"00",X"00",X"33",X"77",X"CF",X"9F",X"BF",X"BF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"CC",X"00",X"FF",X"77",X"11",X"11",X"77",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"EE",X"CC",X"00",X"CC",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"77",X"77",X"00",
		X"CC",X"EE",X"FF",X"FF",X"FF",X"FF",X"77",X"11",X"77",X"77",X"33",X"33",X"11",X"00",X"00",X"00",
		X"33",X"33",X"99",X"DD",X"CC",X"EE",X"EE",X"FF",X"FF",X"00",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"77",X"77",X"33",X"BB",X"99",X"88",X"CC",X"EE",X"EE",X"FF",X"FF",X"FF",X"FF",X"77",X"77",
		X"07",X"0A",X"0C",X"08",X"00",X"00",X"00",X"00",X"8D",X"8A",X"8D",X"8A",X"8F",X"8A",X"8C",X"88",
		X"00",X"00",X"00",X"00",X"08",X"0C",X"06",X"0B",X"88",X"8C",X"8E",X"8B",X"8D",X"8A",X"8D",X"8A",
		X"00",X"00",X"00",X"00",X"80",X"C0",X"60",X"B0",X"80",X"C0",X"60",X"B0",X"50",X"A0",X"50",X"A0",
		X"70",X"A0",X"C0",X"80",X"00",X"00",X"00",X"00",X"50",X"A0",X"50",X"A0",X"70",X"A0",X"C0",X"80",
		X"01",X"03",X"05",X"0E",X"05",X"0A",X"05",X"0A",X"00",X"00",X"00",X"00",X"01",X"03",X"05",X"0E",
		X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"0A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"0C",X"0E",X"0E",X"0E",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"07",X"0F",X"0F",X"00",X"00",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0E",X"0E",X"0E",X"0E",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"07",X"03",X"01",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"00",X"00",
		X"00",X"00",X"08",X"0C",X"0E",X"0E",X"0E",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"07",X"0F",X"05",X"00",X"00",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0E",X"0E",X"0E",X"0E",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"0F",X"07",X"03",X"01",X"00",X"00",X"00",X"0F",X"07",X"0F",X"0F",X"0F",X"07",X"00",X"00",
		X"00",X"00",X"08",X"0C",X"06",X"0E",X"0E",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"07",X"0F",X"05",X"00",X"00",X"07",X"0F",X"0F",X"0C",X"0B",X"05",
		X"0E",X"0E",X"06",X"0E",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"0F",X"07",X"03",X"01",X"00",X"00",X"00",X"0E",X"06",X"0F",X"0F",X"0F",X"07",X"00",X"00",
		X"00",X"00",X"08",X"0C",X"06",X"0E",X"0E",X"0E",X"00",X"01",X"00",X"08",X"00",X"04",X"00",X"02",
		X"0A",X"08",X"04",X"01",X"E0",X"F0",X"70",X"70",X"00",X"00",X"07",X"0F",X"87",X"C0",X"C3",X"C1",
		X"0E",X"0E",X"06",X"0E",X"0C",X"08",X"00",X"00",X"04",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"5A",X"0F",X"06",X"03",X"01",X"00",X"00",X"00",X"0E",X"06",X"0F",X"0F",X"0F",X"07",X"00",X"00",
		X"02",X"06",X"0A",X"0D",X"07",X"0E",X"0E",X"06",X"00",X"00",X"00",X"70",X"30",X"10",X"10",X"00",
		X"01",X"02",X"01",X"F0",X"F0",X"F0",X"F1",X"F3",X"08",X"00",X"07",X"0F",X"CF",X"BF",X"FF",X"FF",
		X"0A",X"0E",X"06",X"0E",X"0C",X"08",X"00",X"00",X"00",X"01",X"00",X"00",X"02",X"00",X"00",X"00",
		X"F7",X"5D",X"3F",X"03",X"14",X"10",X"34",X"08",X"FF",X"DF",X"E9",X"E1",X"C3",X"87",X"04",X"0D",
		X"0D",X"0B",X"01",X"84",X"0F",X"8E",X"8E",X"8F",X"00",X"00",X"00",X"78",X"34",X"03",X"01",X"00",
		X"09",X"00",X"03",X"F0",X"F0",X"F0",X"78",X"1E",X"09",X"0C",X"0C",X"F0",X"F0",X"E1",X"C3",X"97",
		X"8E",X"8B",X"CD",X"00",X"CD",X"0B",X"07",X"0A",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"CF",X"EF",X"BB",X"77",X"33",X"08",X"01",X"03",X"7F",X"FF",X"FF",X"FF",X"FF",X"0E",X"0E",X"0C",
		X"00",X"08",X"0C",X"4A",X"FD",X"F0",X"FD",X"FB",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"70",
		X"00",X"00",X"11",X"22",X"75",X"F8",X"F0",X"F0",X"00",X"03",X"89",X"EE",X"FF",X"FF",X"F3",X"F0",
		X"F7",X"FB",X"FD",X"F0",X"FD",X"4A",X"0C",X"08",X"F0",X"70",X"10",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F8",X"75",X"22",X"11",X"00",X"F0",X"F0",X"F3",X"FF",X"FF",X"EE",X"89",X"03",
		X"00",X"07",X"0E",X"0C",X"FE",X"FC",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",
		X"00",X"00",X"11",X"22",X"77",X"DE",X"DE",X"9E",X"00",X"00",X"CC",X"EF",X"FF",X"FF",X"7F",X"7F",
		X"FF",X"FF",X"FE",X"FC",X"FE",X"0C",X"0E",X"07",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",
		X"9E",X"9E",X"DE",X"DE",X"77",X"22",X"11",X"00",X"7F",X"7F",X"7F",X"FF",X"FF",X"EF",X"CC",X"00",
		X"00",X"88",X"CC",X"EE",X"2E",X"0E",X"0E",X"0E",X"60",X"10",X"70",X"10",X"60",X"00",X"00",X"03",
		X"00",X"32",X"F1",X"33",X"76",X"77",X"3F",X"1F",X"FF",X"FC",X"F3",X"F5",X"FD",X"CF",X"EF",X"FD",
		X"8E",X"8B",X"03",X"01",X"01",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"06",X"0F",X"0F",X"06",
		X"1F",X"01",X"05",X"01",X"09",X"09",X"01",X"01",X"F8",X"FD",X"7F",X"0E",X"0C",X"08",X"08",X"00",
		X"40",X"40",X"E0",X"80",X"FE",X"FE",X"F9",X"FD",X"00",X"00",X"03",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0E",X"0F",X"03",X"01",X"01",X"20",X"10",X"00",X"77",X"FF",X"FF",X"FF",X"FF",
		X"FA",X"FF",X"7F",X"2E",X"0C",X"0C",X"0E",X"0E",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"1F",X"3F",X"11",X"00",X"00",X"00",X"00",X"EF",X"EB",X"E1",X"EB",X"CF",X"03",X"01",X"00",
		X"40",X"50",X"20",X"B8",X"E6",X"FB",X"F1",X"FB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"0C",X"0E",X"07",X"07",X"13",X"17",X"00",X"00",X"00",X"77",X"FF",X"FF",X"FC",X"FF",
		X"F5",X"FF",X"7F",X"2E",X"4C",X"00",X"00",X"00",X"01",X"07",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"7E",X"FC",X"76",X"33",X"00",X"01",X"07",X"BE",X"8F",X"87",X"8F",X"0F",X"0F",X"0E",X"0C",
		X"00",X"00",X"00",X"00",X"88",X"CC",X"EE",X"EE",X"00",X"07",X"00",X"80",X"40",X"F0",X"73",X"B3",
		X"00",X"0E",X"0F",X"33",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"0C",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EE",X"EE",X"CC",X"88",X"00",X"00",X"00",X"00",X"B3",X"73",X"F0",X"40",X"80",X"00",X"07",X"00",
		X"FF",X"FF",X"FF",X"FF",X"33",X"0F",X"0E",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"0C",X"00",X"00",
		X"0E",X"4A",X"2C",X"F0",X"AC",X"C8",X"88",X"88",X"33",X"33",X"33",X"11",X"00",X"00",X"00",X"00",
		X"BC",X"BC",X"DA",X"69",X"1F",X"27",X"01",X"00",X"A7",X"A7",X"7F",X"FF",X"FF",X"FF",X"7F",X"37",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"6E",X"4C",X"08",X"00",X"00",X"00",X"00",
		X"0C",X"0C",X"0C",X"48",X"B8",X"20",X"50",X"00",X"77",X"77",X"77",X"23",X"01",X"00",X"00",X"00",
		X"AD",X"AD",X"A5",X"D3",X"3F",X"5F",X"13",X"01",X"CF",X"CF",X"EF",X"FF",X"FB",X"FD",X"EE",X"EE",
		X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"6E",X"7F",X"17",X"01",X"00",X"00",X"00",X"00",
		X"0E",X"0E",X"1E",X"AC",X"BC",X"A8",X"98",X"00",X"33",X"33",X"33",X"11",X"00",X"00",X"00",X"00",
		X"BC",X"BC",X"DA",X"69",X"1F",X"27",X"01",X"13",X"A7",X"A7",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"13",X"13",X"37",X"3F",X"6E",X"00",X"00",X"00",X"FF",X"FF",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"08",X"08",X"08",X"80",X"60",X"40",X"A0",X"00",X"FF",X"FF",X"FE",X"56",X"03",X"01",X"00",X"00",
		X"5B",X"5B",X"5B",X"B7",X"7F",X"BF",X"37",X"37",X"8F",X"8F",X"CF",X"EF",X"F7",X"EA",X"CC",X"CC",
		X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"13",X"13",X"01",X"00",X"00",X"00",X"00",X"00",X"CC",X"EE",X"7F",X"17",X"01",X"00",X"00",X"00",
		X"00",X"88",X"88",X"CC",X"CC",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",
		X"01",X"03",X"56",X"76",X"EF",X"CF",X"DE",X"FE",X"08",X"3E",X"B6",X"F6",X"7E",X"3E",X"B6",X"F6",
		X"EE",X"EE",X"EE",X"CE",X"CE",X"8E",X"0E",X"0C",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"77",X"33",X"11",X"00",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",
		X"00",X"00",X"10",X"10",X"F0",X"1C",X"1C",X"0C",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"0F",X"77",X"33",X"11",X"33",X"37",X"3F",X"3F",X"00",X"88",X"CC",X"FF",X"CF",X"8F",X"0F",X"0F",
		X"0C",X"0C",X"0C",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"3F",X"3F",X"37",X"32",X"11",X"33",X"77",X"0F",X"87",X"4B",X"AD",X"F0",X"EC",X"C8",X"80",X"00",
		X"0C",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"10",X"00",X"00",X"30",X"00",X"00",X"10",
		X"01",X"00",X"80",X"40",X"F0",X"40",X"80",X"00",X"0F",X"13",X"17",X"1F",X"3F",X"3F",X"37",X"37",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"0C",X"10",X"00",X"00",X"30",X"00",X"00",X"10",X"00",
		X"00",X"80",X"40",X"F0",X"40",X"80",X"00",X"00",X"37",X"37",X"3F",X"3F",X"1F",X"17",X"13",X"0F",
		X"22",X"26",X"B7",X"3F",X"5F",X"5F",X"CE",X"8C",X"00",X"00",X"00",X"00",X"00",X"13",X"17",X"3F",
		X"00",X"00",X"00",X"11",X"11",X"99",X"BA",X"BB",X"30",X"27",X"4F",X"5A",X"D2",X"5E",X"C7",X"EF",
		X"8C",X"8E",X"CE",X"DF",X"DF",X"5F",X"5F",X"14",X"3F",X"3F",X"1F",X"1F",X"07",X"03",X"00",X"00",
		X"CC",X"CC",X"CC",X"EE",X"FF",X"7F",X"0F",X"07",X"6F",X"EF",X"67",X"75",X"FC",X"DE",X"0C",X"00",
		X"00",X"00",X"00",X"08",X"4C",X"4E",X"2E",X"C3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"32",X"23",X"23",X"74",X"77",X"60",X"4E",X"9F",X"A7",X"A7",X"BF",X"9F",X"DF",
		X"8C",X"C2",X"2E",X"CE",X"8C",X"88",X"00",X"00",X"33",X"77",X"EF",X"DF",X"8F",X"CF",X"77",X"33",
		X"89",X"EE",X"3F",X"CF",X"4C",X"6E",X"EE",X"CC",X"CF",X"EF",X"EF",X"EF",X"7F",X"37",X"00",X"00",
		X"C1",X"DB",X"5B",X"B7",X"5E",X"4E",X"9E",X"BC",X"00",X"00",X"00",X"03",X"07",X"0F",X"1F",X"1F",
		X"00",X"00",X"00",X"4C",X"EE",X"EE",X"EE",X"EE",X"00",X"01",X"13",X"74",X"56",X"57",X"F9",X"FF",
		X"2D",X"D3",X"3F",X"CE",X"0C",X"00",X"00",X"00",X"3F",X"3F",X"1F",X"17",X"17",X"03",X"01",X"00",
		X"DF",X"9F",X"9F",X"DF",X"FF",X"7F",X"0F",X"00",X"1E",X"CF",X"EF",X"9F",X"CF",X"7F",X"0E",X"00",
		X"00",X"00",X"08",X"0C",X"0C",X"0C",X"86",X"4A",X"00",X"00",X"01",X"03",X"12",X"01",X"07",X"07",
		X"00",X"0C",X"0E",X"87",X"4B",X"0F",X"0F",X"0F",X"04",X"04",X"0D",X"4B",X"87",X"0F",X"0F",X"C3",
		X"0C",X"0E",X"0E",X"86",X"0E",X"0C",X"08",X"00",X"07",X"07",X"16",X"03",X"03",X"01",X"00",X"00",
		X"1E",X"2D",X"1E",X"87",X"4B",X"09",X"01",X"00",X"2D",X"1E",X"1E",X"0F",X"1E",X"2D",X"0D",X"00",
		X"00",X"0C",X"C0",X"C0",X"00",X"0C",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"11",X"33",X"77",X"7F",X"7F",X"7F",X"02",X"25",X"AD",X"AD",X"AD",X"2D",X"2D",X"0A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"7F",X"7F",X"77",X"77",X"33",X"11",X"00",X"08",X"08",X"08",X"FF",X"FF",X"EE",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"77",X"FF",X"EE",X"CC",X"CC",X"CC",X"88",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"61",X"07",X"01",X"61",X"61",X"07",X"00",
		X"19",X"95",X"B7",X"B7",X"B7",X"A6",X"84",X"08",X"00",X"88",X"CC",X"88",X"88",X"00",X"00",X"00",
		X"00",X"0C",X"C0",X"C0",X"00",X"0C",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"11",X"33",X"33",X"77",X"77",X"77",X"02",X"25",X"AD",X"AD",X"AD",X"AD",X"25",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"77",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",X"77",X"FF",X"FF",
		X"C0",X"C0",X"0C",X"00",X"C0",X"C0",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"77",X"77",X"33",X"33",X"11",X"00",X"00",X"CE",X"25",X"AD",X"AD",X"AD",X"AD",X"25",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"76",X"76",X"F0",X"F0",X"F6",X"FE",X"F8",X"BC",X"80",X"C0",X"C0",X"C0",X"C0",X"88",X"88",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"8F",X"8F",X"8F",X"0F",X"0F",X"07",X"07",X"03",X"88",X"88",X"88",X"08",X"0C",X"0C",X"0C",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"03",X"07",X"07",X"07",X"07",X"0E",X"0E",X"0E",X"0C",X"0C",X"0C",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"34",X"70",X"76",X"F6",X"F0",X"F0",X"73",X"33",X"00",X"80",X"C0",X"C0",X"C0",X"C0",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"30",X"43",X"07",X"07",X"00",X"00",X"00",X"00",X"80",X"0C",X"0C",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"8F",X"8F",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FB",X"FB",X"00",X"00",X"00",X"00",X"00",X"00",X"84",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"70",X"73",X"33",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"40",X"60",X"20",X"38",X"78",X"1C",X"0C",X"00",X"00",X"00",X"10",X"12",X"47",X"EF",X"FF",
		X"08",X"08",X"05",X"D7",X"B7",X"3F",X"7F",X"EF",X"08",X"08",X"CC",X"CF",X"CF",X"CF",X"EF",X"FF",
		X"1C",X"1C",X"1C",X"78",X"28",X"A8",X"C8",X"00",X"FF",X"FF",X"FF",X"77",X"77",X"33",X"11",X"00",
		X"EF",X"EF",X"DF",X"DF",X"DF",X"DF",X"DF",X"03",X"FD",X"FD",X"FD",X"FB",X"FD",X"FD",X"FE",X"1F",
		X"00",X"00",X"00",X"00",X"28",X"18",X"1C",X"1C",X"00",X"00",X"00",X"10",X"12",X"47",X"EF",X"FF",
		X"05",X"05",X"05",X"D7",X"B7",X"3F",X"7F",X"EF",X"00",X"00",X"8C",X"8F",X"CF",X"CF",X"EF",X"FF",
		X"3C",X"1C",X"1C",X"08",X"08",X"88",X"88",X"00",X"FF",X"FF",X"FF",X"77",X"77",X"33",X"11",X"00",
		X"EF",X"DF",X"DF",X"BF",X"BF",X"BF",X"BF",X"03",X"FD",X"FD",X"FD",X"FB",X"FB",X"FD",X"FE",X"0F",
		X"00",X"00",X"10",X"98",X"F8",X"9C",X"9C",X"8C",X"01",X"00",X"11",X"33",X"77",X"77",X"FF",X"FF",
		X"0F",X"7F",X"EF",X"CF",X"CF",X"EF",X"FF",X"FF",X"0F",X"CC",X"7F",X"3F",X"D3",X"A5",X"AD",X"AD",
		X"8C",X"9C",X"9C",X"F8",X"98",X"10",X"00",X"00",X"FF",X"FF",X"77",X"77",X"33",X"11",X"00",X"01",
		X"FF",X"FF",X"EF",X"CF",X"CF",X"EF",X"7F",X"0F",X"AD",X"AD",X"A5",X"D3",X"3F",X"7F",X"CC",X"0F",
		X"00",X"00",X"18",X"D0",X"F0",X"5C",X"DE",X"CF",X"07",X"11",X"00",X"11",X"33",X"BB",X"FF",X"FF",
		X"0F",X"FF",X"F1",X"FF",X"FF",X"FF",X"FF",X"FF",X"08",X"8C",X"EF",X"CF",X"CF",X"EF",X"FF",X"FF",
		X"CF",X"DE",X"5C",X"F0",X"D0",X"18",X"00",X"00",X"FF",X"FF",X"BB",X"33",X"11",X"00",X"11",X"07",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F1",X"FF",X"0F",X"FF",X"FF",X"EF",X"CF",X"CF",X"EF",X"8C",X"08",
		X"0C",X"0C",X"0C",X"48",X"40",X"40",X"E0",X"50",X"FF",X"FF",X"EF",X"47",X"03",X"01",X"00",X"00",
		X"78",X"78",X"A5",X"D3",X"2F",X"5F",X"13",X"37",X"4F",X"6F",X"FF",X"FF",X"FB",X"EC",X"EE",X"FE",
		X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",
		X"7F",X"7F",X"FF",X"FF",X"7F",X"7F",X"17",X"01",X"EE",X"CC",X"CC",X"88",X"88",X"CC",X"EE",X"0E",
		X"0C",X"0C",X"0C",X"48",X"40",X"30",X"20",X"50",X"FF",X"FF",X"EF",X"47",X"03",X"01",X"00",X"00",
		X"AD",X"AD",X"A5",X"D3",X"2F",X"5F",X"13",X"01",X"CF",X"EF",X"FF",X"FF",X"FB",X"EC",X"EE",X"FF",
		X"40",X"00",X"88",X"88",X"CC",X"EE",X"FF",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"13",X"13",X"13",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"07",X"00",
		X"FF",X"FF",X"DD",X"CC",X"C8",X"A8",X"30",X"30",X"3F",X"37",X"23",X"30",X"30",X"01",X"00",X"00",
		X"FF",X"FF",X"7F",X"3F",X"3F",X"7F",X"13",X"17",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"FF",X"EE",
		X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"13",X"13",X"37",X"37",X"7F",X"0F",
		X"7F",X"FF",X"FF",X"FF",X"FF",X"EE",X"CC",X"00",X"CC",X"CC",X"88",X"88",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"DD",X"CC",X"D8",X"B8",X"10",X"10",X"3F",X"37",X"23",X"30",X"30",X"01",X"00",X"00",
		X"FF",X"FF",X"7F",X"3F",X"3F",X"7F",X"13",X"13",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"FF",X"EE",
		X"10",X"00",X"00",X"88",X"CC",X"CC",X"EE",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"13",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"EE",X"FF",X"FF",X"FF",X"7F",X"7F",X"37",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"0C",X"0C",X"0E",X"00",X"00",X"00",X"10",X"12",X"47",X"EF",X"FF",
		X"08",X"08",X"05",X"D7",X"B7",X"3F",X"7F",X"FF",X"08",X"08",X"CC",X"CF",X"CF",X"CF",X"EF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"0C",X"0C",X"0E",X"00",X"00",X"00",X"10",X"12",X"47",X"EF",X"FF",
		X"05",X"05",X"05",X"D7",X"B7",X"3F",X"7F",X"FF",X"00",X"00",X"8C",X"8F",X"CF",X"CF",X"EF",X"FF",
		X"0E",X"0E",X"0C",X"48",X"28",X"A8",X"B8",X"70",X"FF",X"FF",X"FF",X"77",X"77",X"33",X"11",X"00",
		X"FF",X"EF",X"DF",X"DF",X"DF",X"DF",X"BF",X"37",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FE",X"FF",
		X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"13",X"37",X"0F",
		X"37",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"4C",X"FF",X"FF",X"EE",X"EE",X"CC",X"CC",X"00",X"00",
		X"0E",X"0E",X"0E",X"2C",X"28",X"A8",X"B8",X"30",X"FF",X"FF",X"FF",X"77",X"77",X"33",X"11",X"00",
		X"FF",X"FF",X"FF",X"DF",X"DF",X"DF",X"DF",X"13",X"FF",X"FF",X"FF",X"FF",X"FB",X"FD",X"FE",X"EE",
		X"60",X"00",X"00",X"00",X"88",X"88",X"CC",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"37",X"37",X"13",X"13",X"13",X"01",X"00",X"00",X"EE",X"EE",X"FF",X"FF",X"FF",X"FF",X"7F",X"0F",
		X"00",X"00",X"10",X"10",X"78",X"1C",X"2C",X"0C",X"00",X"00",X"01",X"03",X"56",X"FE",X"FF",X"FF",
		X"0F",X"37",X"5F",X"2F",X"B7",X"F5",X"78",X"78",X"0F",X"EE",X"EC",X"FB",X"FF",X"FF",X"6F",X"4F",
		X"0C",X"1C",X"1C",X"78",X"10",X"20",X"88",X"0C",X"FF",X"FF",X"EF",X"47",X"12",X"10",X"00",X"00",
		X"78",X"78",X"7D",X"3F",X"A7",X"D7",X"13",X"03",X"4F",X"6F",X"FF",X"FF",X"FB",X"EC",X"FF",X"0F",
		X"00",X"00",X"10",X"10",X"78",X"1C",X"1C",X"0C",X"0B",X"11",X"01",X"30",X"74",X"EF",X"FF",X"FF",
		X"0F",X"FF",X"7F",X"3F",X"3F",X"7D",X"78",X"78",X"0C",X"CC",X"CC",X"FB",X"FF",X"FF",X"6F",X"4F",
		X"0C",X"0C",X"0C",X"48",X"20",X"70",X"A0",X"28",X"FF",X"FF",X"EF",X"47",X"0B",X"01",X"04",X"00",
		X"78",X"78",X"7D",X"F3",X"E3",X"5F",X"13",X"07",X"4F",X"6F",X"FF",X"FF",X"FB",X"EC",X"FF",X"0F",
		X"0C",X"0C",X"0C",X"48",X"40",X"40",X"E0",X"50",X"FF",X"FF",X"EF",X"47",X"03",X"01",X"00",X"00",
		X"78",X"78",X"A5",X"D3",X"2F",X"5F",X"13",X"37",X"4F",X"6F",X"FF",X"FF",X"FB",X"EC",X"EE",X"FE",
		X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"13",X"13",X"37",X"0F",
		X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"EE",X"0C",X"EE",X"CC",X"CC",X"88",X"88",X"00",X"00",X"00",
		X"0C",X"0C",X"0C",X"48",X"40",X"30",X"20",X"50",X"0F",X"0F",X"1E",X"07",X"03",X"10",X"0C",X"08",
		X"2D",X"2D",X"2D",X"C3",X"C3",X"2D",X"03",X"01",X"0F",X"0F",X"0F",X"0F",X"4B",X"2C",X"0E",X"0F",
		X"40",X"00",X"08",X"08",X"0C",X"0E",X"0F",X"0F",X"01",X"02",X"00",X"08",X"01",X"02",X"00",X"00",
		X"01",X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"00",
		X"00",X"88",X"88",X"CC",X"CC",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",
		X"10",X"12",X"47",X"67",X"FE",X"DE",X"CF",X"EF",X"80",X"B6",X"3E",X"7E",X"F6",X"B6",X"3E",X"7E",
		X"EE",X"EE",X"EE",X"CE",X"CF",X"8F",X"01",X"01",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"77",X"33",X"11",X"00",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"88",X"88",X"CC",X"CC",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",
		X"01",X"03",X"56",X"76",X"EF",X"CF",X"DE",X"FE",X"08",X"3E",X"B6",X"F6",X"7E",X"3E",X"B6",X"F6",
		X"EE",X"EE",X"EE",X"CE",X"CE",X"8E",X"0E",X"0C",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"77",X"33",X"11",X"00",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",
		X"00",X"00",X"00",X"00",X"88",X"88",X"8C",X"8E",X"00",X"11",X"33",X"17",X"C3",X"C3",X"17",X"77",
		X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"88",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"8E",X"8F",X"8B",X"89",X"01",X"02",X"00",X"00",X"77",X"17",X"C3",X"C3",X"17",X"33",X"11",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"88",
		X"00",X"00",X"00",X"00",X"88",X"88",X"8E",X"8E",X"00",X"00",X"11",X"17",X"C3",X"C3",X"17",X"77",
		X"00",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"88",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"8F",X"8F",X"89",X"88",X"00",X"00",X"00",X"00",X"77",X"17",X"C3",X"C3",X"17",X"11",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"88",X"00",
		X"00",X"88",X"88",X"C4",X"C4",X"2E",X"2E",X"A6",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",
		X"00",X"31",X"56",X"56",X"AD",X"AD",X"1E",X"1E",X"00",X"FA",X"96",X"87",X"4B",X"5A",X"96",X"87",
		X"A6",X"2E",X"2E",X"C4",X"4C",X"4C",X"8F",X"06",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",
		X"2D",X"0F",X"8F",X"8F",X"47",X"23",X"11",X"00",X"4B",X"1E",X"1E",X"0F",X"0F",X"0F",X"FF",X"00",
		X"00",X"88",X"88",X"4C",X"4C",X"2E",X"A6",X"A6",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",
		X"00",X"31",X"56",X"56",X"AD",X"AD",X"1E",X"1E",X"00",X"FA",X"96",X"96",X"5A",X"5A",X"96",X"87",
		X"A6",X"A6",X"A6",X"4E",X"4E",X"8E",X"0C",X"08",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",
		X"2D",X"0F",X"8F",X"8F",X"47",X"23",X"11",X"00",X"4B",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"01",
		X"00",X"00",X"00",X"00",X"00",X"88",X"4C",X"2E",X"00",X"00",X"00",X"00",X"00",X"33",X"43",X"74",
		X"00",X"00",X"00",X"33",X"CF",X"0F",X"C3",X"3C",X"00",X"00",X"00",X"CC",X"3F",X"0F",X"87",X"0F",
		X"2E",X"2E",X"2E",X"2E",X"2F",X"CF",X"03",X"02",X"74",X"43",X"47",X"61",X"76",X"11",X"00",X"00",
		X"3C",X"C3",X"0F",X"69",X"96",X"8F",X"77",X"00",X"0F",X"87",X"0F",X"69",X"96",X"1F",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"88",X"4C",X"2E",X"00",X"00",X"00",X"00",X"00",X"33",X"43",X"74",
		X"00",X"00",X"00",X"33",X"CF",X"0F",X"C3",X"3C",X"00",X"00",X"00",X"CC",X"3F",X"0F",X"87",X"0F",
		X"2E",X"2E",X"2E",X"2F",X"4F",X"8E",X"0C",X"00",X"74",X"43",X"47",X"70",X"67",X"11",X"00",X"00",
		X"3C",X"C3",X"0F",X"E1",X"3C",X"8F",X"77",X"00",X"0F",X"87",X"0F",X"0F",X"E1",X"1F",X"EF",X"00",
		X"00",X"00",X"88",X"88",X"88",X"88",X"88",X"88",X"00",X"00",X"33",X"22",X"22",X"22",X"22",X"22",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"88",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"22",X"22",X"22",X"22",X"33",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"CC",X"22",X"22",X"EE",X"00",X"EE",X"44",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"22",X"22",X"33",X"00",X"33",X"00",X"00",
		X"00",X"EE",X"00",X"22",X"AA",X"AA",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"00",X"22",X"22",X"22",X"33",X"00",
		X"00",X"44",X"44",X"66",X"66",X"EE",X"EE",X"EE",X"00",X"00",X"11",X"11",X"11",X"33",X"33",X"33",
		X"60",X"69",X"0F",X"9F",X"F9",X"69",X"0F",X"9F",X"00",X"88",X"88",X"88",X"88",X"88",X"88",X"CC",
		X"EE",X"EE",X"EE",X"CE",X"CE",X"8E",X"06",X"0C",X"33",X"33",X"11",X"11",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"11",X"00",X"CC",X"DD",X"DD",X"DD",X"FF",X"FF",X"FF",X"00",
		X"00",X"88",X"88",X"CC",X"CC",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",
		X"10",X"12",X"47",X"67",X"FE",X"DE",X"CF",X"EF",X"80",X"B6",X"3E",X"7E",X"F6",X"B6",X"3E",X"7E",
		X"EE",X"EE",X"EE",X"CE",X"CE",X"8E",X"06",X"0C",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"77",X"33",X"11",X"00",X"FE",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"88",X"CC",X"CC",X"EE",X"EE",X"17",X"C3",X"C3",X"17",X"77",X"11",X"00",X"00",
		X"9F",X"C3",X"C3",X"9F",X"FF",X"FF",X"77",X"11",X"88",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EE",X"EE",X"66",X"EE",X"CD",X"8F",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",
		X"00",X"00",X"00",X"00",X"00",X"33",X"FF",X"00",X"77",X"11",X"00",X"11",X"77",X"FF",X"EF",X"00",
		X"00",X"00",X"00",X"00",X"88",X"CC",X"CC",X"EE",X"00",X"00",X"17",X"C3",X"C3",X"17",X"77",X"00",
		X"00",X"77",X"9F",X"C3",X"C3",X"9F",X"FF",X"FF",X"00",X"00",X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EE",X"EE",X"EE",X"EE",X"CD",X"8F",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",
		X"11",X"00",X"00",X"00",X"11",X"FF",X"FF",X"00",X"FF",X"33",X"00",X"33",X"FF",X"FF",X"EF",X"00",
		X"00",X"00",X"00",X"00",X"88",X"CC",X"CC",X"EE",X"00",X"00",X"00",X"33",X"17",X"C3",X"C3",X"17",
		X"00",X"00",X"77",X"FF",X"9F",X"C3",X"C3",X"9F",X"00",X"00",X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EE",X"EE",X"EE",X"EE",X"CD",X"8F",X"0E",X"00",X"77",X"00",X"00",X"00",X"00",X"77",X"11",X"00",
		X"FF",X"11",X"00",X"00",X"77",X"FF",X"FF",X"00",X"FF",X"FF",X"00",X"77",X"FF",X"FF",X"EF",X"00",
		X"00",X"00",X"00",X"88",X"CC",X"CC",X"EE",X"EE",X"00",X"00",X"00",X"11",X"33",X"77",X"17",X"C3",
		X"00",X"00",X"77",X"FF",X"FF",X"FF",X"9F",X"C3",X"00",X"00",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EE",X"EE",X"EE",X"EE",X"CD",X"8F",X"0E",X"00",X"C3",X"17",X"77",X"70",X"77",X"11",X"00",X"00",
		X"C3",X"9F",X"FF",X"F0",X"FF",X"FF",X"77",X"00",X"FF",X"FF",X"FF",X"F0",X"FF",X"FF",X"EF",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
