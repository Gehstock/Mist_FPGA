`define BUILD_DATE "190321"
`define BUILD_TIME "135526"
