library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity squash_program is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of squash_program is
	type rom is array(0 to  12287) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"F3",X"C3",X"91",X"04",X"FF",X"FF",X"FF",X"FF",X"AF",X"32",X"05",X"A0",X"78",X"D3",X"08",X"79",
		X"D3",X"09",X"3E",X"01",X"32",X"05",X"A0",X"C9",X"AF",X"32",X"05",X"A0",X"78",X"D3",X"08",X"DB",
		X"0C",X"4F",X"3E",X"01",X"32",X"05",X"A0",X"C9",X"87",X"85",X"6F",X"7C",X"CE",X"00",X"67",X"7E",
		X"23",X"66",X"6F",X"E9",X"FF",X"FF",X"FF",X"FF",X"F3",X"F5",X"C5",X"D5",X"E5",X"08",X"D9",X"F5",
		X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",X"AF",X"32",X"00",X"A0",X"3A",X"00",X"B8",X"CD",X"EC",
		X"1C",X"CD",X"41",X"04",X"CD",X"17",X"04",X"CD",X"F5",X"04",X"CD",X"5A",X"01",X"CD",X"7E",X"04",
		X"CD",X"10",X"03",X"CD",X"2E",X"03",X"CD",X"B6",X"00",X"CD",X"DE",X"02",X"CD",X"0C",X"02",X"3A",
		X"00",X"B8",X"CD",X"55",X"02",X"CD",X"B1",X"02",X"CD",X"8A",X"01",X"CD",X"CB",X"01",X"CD",X"2A",
		X"01",X"CD",X"5A",X"01",X"CD",X"4C",X"03",X"CD",X"9C",X"03",X"3A",X"31",X"70",X"B7",X"28",X"09",
		X"21",X"9E",X"8B",X"3A",X"14",X"70",X"CD",X"EA",X"03",X"3A",X"00",X"B8",X"3E",X"01",X"32",X"00",
		X"A0",X"32",X"03",X"A0",X"ED",X"56",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"F1",X"D9",X"08",
		X"E1",X"D1",X"C1",X"F1",X"FB",X"C9",X"1E",X"00",X"3A",X"14",X"70",X"FE",X"5A",X"D0",X"DD",X"21",
		X"15",X"70",X"3A",X"00",X"70",X"21",X"10",X"70",X"47",X"AE",X"70",X"A0",X"CB",X"47",X"F5",X"C4",
		X"F5",X"00",X"F1",X"DD",X"23",X"1C",X"CB",X"4F",X"C4",X"F5",X"00",X"DD",X"23",X"1C",X"3A",X"01",
		X"70",X"21",X"11",X"70",X"47",X"AE",X"70",X"A0",X"CB",X"47",X"F5",X"C4",X"F5",X"00",X"F1",X"DD",
		X"23",X"1C",X"CB",X"4F",X"C8",X"3E",X"07",X"32",X"BA",X"70",X"3A",X"02",X"70",X"CB",X"47",X"20",
		X"18",X"16",X"00",X"21",X"15",X"01",X"19",X"7E",X"21",X"05",X"70",X"57",X"86",X"77",X"7A",X"21",
		X"14",X"70",X"86",X"77",X"C9",X"01",X"02",X"03",X"04",X"3E",X"01",X"DD",X"BE",X"00",X"28",X"04",
		X"DD",X"34",X"00",X"C9",X"DD",X"36",X"00",X"00",X"18",X"D7",X"3A",X"2B",X"70",X"B7",X"C8",X"21",
		X"2C",X"70",X"34",X"3E",X"03",X"BE",X"C0",X"36",X"00",X"3A",X"2B",X"70",X"3D",X"32",X"2B",X"70",
		X"B7",X"28",X"0B",X"3A",X"2D",X"70",X"EE",X"01",X"32",X"2D",X"70",X"B7",X"20",X"06",X"3E",X"0D",
		X"32",X"61",X"70",X"C9",X"3E",X"0E",X"32",X"61",X"70",X"C9",X"3A",X"2E",X"70",X"B7",X"C8",X"21",
		X"2F",X"70",X"34",X"3E",X"03",X"BE",X"C0",X"36",X"00",X"3A",X"2E",X"70",X"3D",X"32",X"2E",X"70",
		X"B7",X"28",X"0B",X"3A",X"30",X"70",X"EE",X"01",X"32",X"30",X"70",X"B7",X"20",X"06",X"3E",X"0D",
		X"32",X"7D",X"70",X"C9",X"3E",X"0E",X"32",X"7D",X"70",X"C9",X"3A",X"26",X"70",X"B7",X"C8",X"21",
		X"24",X"70",X"34",X"3E",X"02",X"BE",X"C0",X"36",X"00",X"21",X"25",X"70",X"3A",X"23",X"70",X"B7",
		X"20",X"17",X"3A",X"5A",X"70",X"3C",X"32",X"5A",X"70",X"34",X"3E",X"04",X"BE",X"C0",X"3A",X"23",
		X"70",X"EE",X"01",X"32",X"23",X"70",X"36",X"00",X"C9",X"3E",X"03",X"BE",X"20",X"07",X"3A",X"26",
		X"70",X"3D",X"32",X"26",X"70",X"3A",X"5A",X"70",X"3D",X"18",X"DB",X"3A",X"2A",X"70",X"B7",X"C8",
		X"21",X"28",X"70",X"34",X"3E",X"02",X"BE",X"C0",X"36",X"00",X"21",X"29",X"70",X"3A",X"27",X"70",
		X"B7",X"20",X"17",X"3A",X"76",X"70",X"3C",X"32",X"76",X"70",X"34",X"3E",X"04",X"BE",X"C0",X"3A",
		X"27",X"70",X"EE",X"01",X"32",X"27",X"70",X"36",X"00",X"C9",X"3E",X"03",X"BE",X"20",X"07",X"3A",
		X"2A",X"70",X"3D",X"32",X"2A",X"70",X"3A",X"76",X"70",X"3D",X"18",X"DB",X"3A",X"3D",X"70",X"B7",
		X"C0",X"3A",X"1A",X"70",X"FE",X"02",X"CA",X"49",X"02",X"FE",X"03",X"CA",X"4F",X"02",X"B7",X"C8",
		X"21",X"1D",X"70",X"7E",X"3C",X"77",X"FE",X"14",X"C0",X"36",X"00",X"3A",X"1C",X"70",X"EE",X"01",
		X"32",X"1C",X"70",X"B7",X"28",X"0F",X"3E",X"04",X"32",X"FB",X"70",X"21",X"66",X"02",X"22",X"F9",
		X"70",X"CD",X"2D",X"26",X"C9",X"3E",X"07",X"18",X"EF",X"AF",X"32",X"1A",X"70",X"18",X"E7",X"AF",
		X"32",X"1A",X"70",X"18",X"F0",X"3A",X"3D",X"70",X"B7",X"C0",X"3A",X"1B",X"70",X"FE",X"03",X"CA",
		X"9D",X"02",X"FE",X"04",X"CA",X"A3",X"02",X"FE",X"05",X"CA",X"A9",X"02",X"B7",X"C8",X"21",X"1E",
		X"70",X"34",X"3E",X"14",X"BE",X"C0",X"36",X"00",X"3A",X"1F",X"70",X"EE",X"01",X"32",X"1F",X"70",
		X"B7",X"28",X"2A",X"3A",X"1B",X"70",X"FE",X"02",X"28",X"0F",X"3E",X"05",X"32",X"FB",X"70",X"21",
		X"76",X"02",X"22",X"F9",X"70",X"CD",X"2D",X"26",X"C9",X"3E",X"06",X"18",X"EF",X"AF",X"32",X"1B",
		X"70",X"18",X"F6",X"AF",X"32",X"1B",X"70",X"18",X"E1",X"AF",X"32",X"1B",X"70",X"3E",X"07",X"18",
		X"DB",X"3A",X"20",X"70",X"B7",X"C8",X"21",X"21",X"70",X"34",X"3E",X"14",X"BE",X"C0",X"36",X"00",
		X"3A",X"22",X"70",X"EE",X"01",X"32",X"22",X"70",X"B7",X"28",X"0F",X"3E",X"01",X"32",X"F7",X"70",
		X"21",X"68",X"02",X"22",X"F5",X"70",X"CD",X"D6",X"23",X"C9",X"3E",X"02",X"18",X"EF",X"3A",X"02",
		X"70",X"E6",X"06",X"CB",X"3F",X"5F",X"16",X"00",X"21",X"0C",X"03",X"19",X"7E",X"32",X"19",X"70",
		X"3A",X"02",X"70",X"E6",X"18",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"32",X"96",X"70",X"3A",X"02",
		X"70",X"E6",X"40",X"B7",X"28",X"02",X"3E",X"01",X"32",X"3C",X"70",X"C9",X"07",X"0B",X"0F",X"15",
		X"3A",X"61",X"70",X"21",X"0C",X"70",X"5F",X"AE",X"73",X"A3",X"B7",X"21",X"0E",X"70",X"28",X"09",
		X"3E",X"FF",X"BE",X"C8",X"7E",X"C6",X"05",X"77",X"C9",X"AF",X"BE",X"C8",X"35",X"C9",X"3A",X"7D",
		X"70",X"21",X"0D",X"70",X"5F",X"AE",X"73",X"A3",X"B7",X"21",X"0F",X"70",X"28",X"09",X"3E",X"FF",
		X"BE",X"C8",X"7E",X"C6",X"05",X"77",X"C9",X"AF",X"BE",X"C8",X"35",X"C9",X"3A",X"37",X"70",X"B7",
		X"28",X"13",X"21",X"38",X"70",X"34",X"3E",X"07",X"BE",X"C0",X"36",X"00",X"3A",X"36",X"70",X"EE",
		X"08",X"32",X"36",X"70",X"C9",X"3E",X"05",X"32",X"36",X"70",X"C9",X"FE",X"64",X"D0",X"DD",X"21",
		X"9A",X"03",X"E5",X"16",X"02",X"DD",X"46",X"00",X"0E",X"00",X"90",X"38",X"03",X"0C",X"18",X"FA",
		X"80",X"71",X"CB",X"E4",X"F5",X"3A",X"36",X"70",X"77",X"F1",X"CB",X"A4",X"23",X"15",X"28",X"05",
		X"DD",X"23",X"C3",X"75",X"03",X"E1",X"7E",X"B7",X"C0",X"C9",X"0A",X"01",X"3A",X"3A",X"70",X"B7",
		X"28",X"13",X"21",X"3B",X"70",X"34",X"3E",X"07",X"BE",X"C0",X"36",X"00",X"3A",X"39",X"70",X"EE",
		X"08",X"32",X"39",X"70",X"C9",X"3E",X"05",X"32",X"39",X"70",X"C9",X"FE",X"64",X"D0",X"DD",X"21",
		X"9A",X"03",X"E5",X"16",X"02",X"DD",X"46",X"00",X"0E",X"00",X"90",X"38",X"03",X"0C",X"18",X"FA",
		X"80",X"71",X"CB",X"E4",X"F5",X"3A",X"39",X"70",X"77",X"F1",X"CB",X"A4",X"23",X"15",X"28",X"05",
		X"DD",X"23",X"C3",X"C5",X"03",X"E1",X"7E",X"B7",X"C0",X"C9",X"FE",X"64",X"D0",X"DD",X"21",X"9A",
		X"03",X"E5",X"16",X"02",X"DD",X"46",X"00",X"0E",X"00",X"90",X"38",X"03",X"0C",X"18",X"FA",X"80",
		X"71",X"CB",X"E4",X"F5",X"36",X"05",X"F1",X"CB",X"A4",X"23",X"15",X"28",X"05",X"DD",X"23",X"C3",
		X"F4",X"03",X"E1",X"7E",X"B7",X"C0",X"C9",X"3A",X"03",X"70",X"3C",X"32",X"03",X"70",X"FE",X"09",
		X"C0",X"AF",X"32",X"03",X"70",X"3A",X"04",X"70",X"EE",X"01",X"32",X"04",X"70",X"B7",X"20",X"04",
		X"32",X"04",X"A0",X"C9",X"21",X"05",X"70",X"7E",X"B7",X"C8",X"3E",X"01",X"32",X"04",X"A0",X"35",
		X"C9",X"06",X"0E",X"DF",X"79",X"2F",X"32",X"00",X"70",X"06",X"0F",X"DF",X"79",X"2F",X"32",X"01",
		X"70",X"3A",X"00",X"A8",X"2F",X"32",X"02",X"70",X"CB",X"7F",X"28",X"01",X"C9",X"CD",X"F4",X"05",
		X"21",X"E5",X"98",X"11",X"69",X"04",X"C3",X"D0",X"04",X"40",X"43",X"4F",X"50",X"49",X"41",X"40",
		X"4D",X"41",X"4C",X"40",X"45",X"46",X"45",X"43",X"54",X"55",X"41",X"44",X"41",X"3F",X"3A",X"0B",
		X"70",X"3C",X"32",X"0B",X"70",X"FE",X"10",X"C0",X"AF",X"32",X"0B",X"70",X"3C",X"32",X"4E",X"70",
		X"C9",X"21",X"40",X"88",X"01",X"FF",X"03",X"36",X"10",X"CB",X"E4",X"36",X"00",X"CB",X"A4",X"23",
		X"0B",X"78",X"B1",X"20",X"F2",X"21",X"00",X"98",X"06",X"20",X"36",X"00",X"23",X"10",X"FB",X"21",
		X"00",X"70",X"01",X"FF",X"07",X"3E",X"FF",X"77",X"BE",X"20",X"0F",X"3E",X"00",X"77",X"BE",X"20",
		X"09",X"23",X"0B",X"78",X"B1",X"20",X"EE",X"C3",X"13",X"06",X"21",X"AA",X"89",X"11",X"ED",X"04",
		X"1A",X"FE",X"3F",X"28",X"0D",X"D6",X"30",X"77",X"CB",X"E4",X"36",X"00",X"CB",X"A4",X"23",X"13",
		X"18",X"EE",X"3A",X"00",X"B8",X"3E",X"01",X"32",X"03",X"A0",X"C3",X"E2",X"04",X"42",X"41",X"44",
		X"40",X"52",X"41",X"4D",X"3F",X"3A",X"09",X"70",X"B7",X"C0",X"01",X"25",X"05",X"3A",X"00",X"70",
		X"E6",X"1F",X"21",X"06",X"70",X"5F",X"AE",X"73",X"A3",X"B7",X"C8",X"5F",X"3A",X"0A",X"70",X"6F",
		X"26",X"00",X"09",X"3C",X"32",X"0A",X"70",X"7E",X"FE",X"C9",X"CA",X"2E",X"05",X"A3",X"C0",X"3E",
		X"FF",X"32",X"09",X"70",X"C9",X"01",X"02",X"08",X"08",X"10",X"04",X"01",X"01",X"C9",X"CD",X"F4",
		X"05",X"21",X"C5",X"88",X"11",X"8E",X"05",X"CD",X"7C",X"05",X"21",X"05",X"89",X"11",X"9D",X"05",
		X"CD",X"7C",X"05",X"21",X"45",X"89",X"11",X"A0",X"05",X"CD",X"7C",X"05",X"21",X"85",X"89",X"11",
		X"AE",X"05",X"CD",X"7C",X"05",X"21",X"C5",X"89",X"11",X"BC",X"05",X"CD",X"7C",X"05",X"21",X"05",
		X"8A",X"11",X"C7",X"05",X"CD",X"7C",X"05",X"21",X"45",X"8A",X"11",X"D6",X"05",X"CD",X"7C",X"05",
		X"21",X"85",X"8A",X"11",X"E5",X"05",X"CD",X"7C",X"05",X"C3",X"E2",X"04",X"1A",X"FE",X"FF",X"C8",
		X"3D",X"3D",X"77",X"CB",X"E4",X"36",X"00",X"CB",X"A4",X"23",X"13",X"C3",X"7C",X"05",X"15",X"21",
		X"22",X"2B",X"24",X"1B",X"19",X"1A",X"26",X"12",X"03",X"0B",X"0A",X"06",X"FF",X"14",X"2B",X"FF",
		X"1B",X"26",X"1B",X"25",X"13",X"12",X"22",X"13",X"1E",X"13",X"1F",X"21",X"25",X"FF",X"22",X"24",
		X"21",X"19",X"24",X"13",X"1F",X"13",X"16",X"21",X"24",X"17",X"25",X"FF",X"1A",X"17",X"20",X"1D",
		X"12",X"25",X"22",X"1B",X"26",X"25",X"FF",X"1C",X"21",X"25",X"17",X"22",X"12",X"1F",X"0C",X"12",
		X"22",X"17",X"26",X"1B",X"26",X"FF",X"1C",X"21",X"25",X"17",X"22",X"12",X"1F",X"21",X"24",X"1B",
		X"1E",X"1E",X"13",X"25",X"FF",X"16",X"1B",X"15",X"1B",X"17",X"1F",X"14",X"24",X"17",X"12",X"03",
		X"0B",X"0A",X"06",X"FF",X"21",X"40",X"88",X"01",X"FF",X"03",X"36",X"10",X"CB",X"E4",X"36",X"00",
		X"CB",X"A4",X"23",X"0B",X"78",X"B1",X"20",X"F2",X"21",X"00",X"98",X"06",X"20",X"36",X"00",X"23",
		X"10",X"FB",X"C9",X"31",X"FF",X"77",X"AF",X"32",X"01",X"A0",X"32",X"02",X"A0",X"3A",X"00",X"B8",
		X"3E",X"01",X"32",X"05",X"A0",X"32",X"06",X"A0",X"0E",X"38",X"06",X"07",X"CF",X"CD",X"92",X"1D",
		X"ED",X"56",X"3E",X"01",X"32",X"00",X"A0",X"FB",X"CD",X"1F",X"08",X"3A",X"00",X"B8",X"00",X"CD",
		X"79",X"08",X"CD",X"C3",X"07",X"3E",X"01",X"32",X"31",X"70",X"32",X"20",X"70",X"32",X"3D",X"70",
		X"32",X"6C",X"70",X"32",X"87",X"70",X"AF",X"32",X"33",X"70",X"01",X"00",X"20",X"C5",X"D5",X"16",
		X"13",X"CD",X"B6",X"21",X"CD",X"E1",X"08",X"CD",X"EA",X"0B",X"CD",X"03",X"0E",X"CD",X"A3",X"17",
		X"01",X"00",X"02",X"0B",X"78",X"B1",X"20",X"FB",X"D1",X"C1",X"3A",X"14",X"70",X"B7",X"20",X"05",
		X"0B",X"78",X"B1",X"20",X"D8",X"AF",X"32",X"20",X"70",X"32",X"31",X"70",X"CD",X"F4",X"05",X"F3",
		X"21",X"56",X"03",X"22",X"F5",X"70",X"3E",X"06",X"32",X"F7",X"70",X"3A",X"00",X"B8",X"CD",X"D6",
		X"23",X"FB",X"3A",X"14",X"70",X"B7",X"28",X"5A",X"FE",X"01",X"28",X"28",X"3E",X"01",X"32",X"31",
		X"70",X"F3",X"21",X"43",X"01",X"22",X"F5",X"70",X"3E",X"03",X"32",X"F7",X"70",X"3A",X"00",X"B8",
		X"CD",X"D6",X"23",X"FB",X"3A",X"00",X"70",X"CB",X"57",X"20",X"2A",X"3A",X"01",X"70",X"CB",X"57",
		X"20",X"27",X"18",X"CE",X"F3",X"21",X"43",X"01",X"22",X"F5",X"70",X"3E",X"04",X"32",X"F7",X"70",
		X"3A",X"00",X"B8",X"CD",X"D6",X"23",X"FB",X"3E",X"01",X"32",X"31",X"70",X"3A",X"00",X"70",X"CB",
		X"57",X"20",X"02",X"18",X"AD",X"3E",X"01",X"18",X"02",X"3E",X"02",X"F5",X"3E",X"01",X"32",X"BA",
		X"70",X"F1",X"32",X"33",X"70",X"CD",X"C3",X"07",X"F3",X"21",X"00",X"00",X"22",X"F9",X"70",X"3E",
		X"02",X"32",X"FB",X"70",X"CD",X"2D",X"26",X"FB",X"3A",X"14",X"70",X"B7",X"20",X"47",X"21",X"FF",
		X"3F",X"22",X"34",X"70",X"AF",X"32",X"33",X"70",X"01",X"F0",X"00",X"0B",X"78",X"B1",X"20",X"FB",
		X"CD",X"A3",X"17",X"CD",X"EA",X"0B",X"CD",X"03",X"0E",X"16",X"13",X"CD",X"B6",X"21",X"3A",X"12",
		X"70",X"21",X"EE",X"88",X"CD",X"6B",X"03",X"3A",X"13",X"70",X"21",X"F1",X"88",X"CD",X"BB",X"03",
		X"3A",X"14",X"70",X"B7",X"C2",X"85",X"06",X"2A",X"34",X"70",X"2B",X"22",X"34",X"70",X"7C",X"B5",
		X"20",X"C6",X"C3",X"3E",X"06",X"AF",X"32",X"AF",X"70",X"3E",X"FF",X"32",X"3E",X"70",X"21",X"14",
		X"70",X"3A",X"33",X"70",X"FE",X"01",X"28",X"01",X"35",X"35",X"3A",X"9D",X"70",X"3D",X"20",X"FD",
		X"3A",X"3E",X"70",X"B7",X"28",X"06",X"3D",X"32",X"3E",X"70",X"18",X"03",X"CD",X"A3",X"17",X"CD",
		X"EA",X"0B",X"CD",X"03",X"0E",X"16",X"13",X"CD",X"B6",X"21",X"3A",X"00",X"B8",X"3A",X"12",X"70",
		X"21",X"EE",X"88",X"CD",X"6B",X"03",X"3A",X"13",X"70",X"21",X"F1",X"88",X"CD",X"BB",X"03",X"3A",
		X"AF",X"70",X"B7",X"C2",X"B9",X"07",X"C3",X"7A",X"07",X"3A",X"14",X"70",X"B7",X"CA",X"3E",X"06",
		X"C3",X"85",X"06",X"3E",X"60",X"32",X"5B",X"70",X"3E",X"90",X"32",X"77",X"70",X"3E",X"0C",X"32",
		X"5C",X"70",X"CB",X"F7",X"32",X"78",X"70",X"3E",X"02",X"32",X"64",X"70",X"32",X"80",X"70",X"3E",
		X"38",X"32",X"5A",X"70",X"32",X"76",X"70",X"AF",X"32",X"20",X"70",X"32",X"31",X"70",X"32",X"F2",
		X"70",X"32",X"32",X"70",X"32",X"3D",X"70",X"32",X"61",X"70",X"32",X"7D",X"70",X"32",X"66",X"70",
		X"32",X"82",X"70",X"32",X"37",X"70",X"32",X"3A",X"70",X"CD",X"81",X"1C",X"CD",X"19",X"22",X"3E",
		X"80",X"32",X"9D",X"70",X"3E",X"10",X"32",X"00",X"98",X"3E",X"04",X"32",X"01",X"98",X"C9",X"0E",
		X"16",X"21",X"A0",X"88",X"06",X"20",X"36",X"C4",X"CB",X"E4",X"36",X"04",X"CB",X"A4",X"23",X"10",
		X"F5",X"0D",X"20",X"F0",X"DD",X"21",X"EC",X"89",X"3E",X"C5",X"CD",X"53",X"08",X"DD",X"21",X"90",
		X"89",X"3E",X"C6",X"CD",X"53",X"08",X"DD",X"21",X"F4",X"89",X"3E",X"C7",X"CD",X"53",X"08",X"CD",
		X"C3",X"08",X"C9",X"CD",X"5D",X"08",X"3E",X"06",X"11",X"00",X"10",X"DD",X"19",X"DD",X"77",X"00",
		X"DD",X"77",X"01",X"DD",X"77",X"1F",X"DD",X"77",X"20",X"DD",X"77",X"21",X"DD",X"77",X"FF",X"DD",
		X"77",X"DF",X"DD",X"77",X"E0",X"DD",X"77",X"E1",X"C9",X"CD",X"F4",X"05",X"21",X"49",X"00",X"22",
		X"F9",X"70",X"3E",X"01",X"32",X"FB",X"70",X"CD",X"2D",X"26",X"21",X"2B",X"01",X"22",X"F5",X"70",
		X"3E",X"00",X"32",X"F7",X"70",X"CD",X"D6",X"23",X"21",X"65",X"01",X"22",X"F9",X"70",X"3E",X"00",
		X"32",X"FB",X"70",X"CD",X"2D",X"26",X"21",X"24",X"02",X"22",X"F5",X"70",X"3E",X"07",X"32",X"F7",
		X"70",X"CD",X"D6",X"23",X"21",X"56",X"03",X"22",X"F5",X"70",X"3E",X"06",X"32",X"F7",X"70",X"CD",
		X"D6",X"23",X"C9",X"16",X"04",X"01",X"00",X"00",X"0B",X"78",X"B1",X"20",X"FB",X"15",X"20",X"F5",
		X"C9",X"01",X"02",X"04",X"07",X"0A",X"0D",X"10",X"15",X"18",X"1B",X"1E",X"21",X"24",X"27",X"29",
		X"2C",X"2A",X"52",X"70",X"3A",X"9C",X"70",X"16",X"00",X"5F",X"19",X"22",X"52",X"70",X"7C",X"FE",
		X"01",X"C0",X"AF",X"67",X"22",X"52",X"70",X"CD",X"60",X"0A",X"3A",X"8E",X"70",X"B7",X"20",X"11",
		X"3A",X"44",X"70",X"FE",X"7C",X"3E",X"01",X"38",X"05",X"32",X"B3",X"70",X"18",X"03",X"32",X"B2",
		X"70",X"3A",X"4E",X"70",X"FE",X"01",X"C2",X"36",X"09",X"AF",X"32",X"4E",X"70",X"3A",X"4B",X"70",
		X"B7",X"C8",X"FE",X"07",X"38",X"10",X"08",X"3A",X"48",X"70",X"FE",X"03",X"30",X"08",X"08",X"3D",
		X"32",X"4B",X"70",X"CD",X"54",X"0A",X"CD",X"80",X"0B",X"3A",X"4B",X"70",X"CB",X"07",X"CB",X"07",
		X"CB",X"07",X"CB",X"07",X"2A",X"4C",X"70",X"16",X"00",X"5F",X"19",X"22",X"4C",X"70",X"7C",X"FE",
		X"00",X"C8",X"AF",X"67",X"22",X"4C",X"70",X"CD",X"AB",X"0A",X"3A",X"48",X"70",X"FE",X"01",X"28",
		X"30",X"FE",X"02",X"28",X"4D",X"FE",X"03",X"28",X"14",X"ED",X"5B",X"3F",X"70",X"2A",X"45",X"70",
		X"97",X"ED",X"52",X"22",X"45",X"70",X"7C",X"32",X"02",X"98",X"18",X"45",X"C9",X"ED",X"5B",X"3F",
		X"70",X"2A",X"45",X"70",X"97",X"ED",X"52",X"22",X"45",X"70",X"7C",X"32",X"02",X"98",X"18",X"10",
		X"C9",X"ED",X"5B",X"3F",X"70",X"2A",X"45",X"70",X"19",X"22",X"45",X"70",X"7C",X"32",X"02",X"98",
		X"ED",X"5B",X"41",X"70",X"2A",X"43",X"70",X"97",X"ED",X"52",X"22",X"43",X"70",X"7C",X"32",X"03",
		X"98",X"C9",X"ED",X"5B",X"3F",X"70",X"2A",X"45",X"70",X"19",X"22",X"45",X"70",X"7C",X"32",X"02",
		X"98",X"ED",X"5B",X"41",X"70",X"2A",X"43",X"70",X"19",X"22",X"43",X"70",X"7C",X"32",X"03",X"98",
		X"C9",X"3A",X"8E",X"70",X"B7",X"C0",X"3A",X"4B",X"70",X"B7",X"20",X"0B",X"3A",X"44",X"70",X"FE",
		X"7C",X"DA",X"1C",X"0A",X"C3",X"4B",X"0A",X"3A",X"49",X"70",X"FE",X"03",X"38",X"03",X"C3",X"4B",
		X"0A",X"3A",X"4A",X"70",X"FE",X"03",X"38",X"03",X"C3",X"1C",X"0A",X"3A",X"44",X"70",X"FE",X"7E",
		X"D0",X"FE",X"7A",X"D8",X"3A",X"46",X"70",X"FE",X"39",X"D0",X"FE",X"23",X"D8",X"3A",X"48",X"70",
		X"FE",X"01",X"28",X"37",X"FE",X"02",X"28",X"04",X"FE",X"03",X"28",X"2F",X"3E",X"00",X"32",X"51",
		X"70",X"3E",X"03",X"32",X"48",X"70",X"CD",X"76",X"18",X"3E",X"02",X"32",X"4B",X"70",X"3E",X"1C",
		X"32",X"47",X"70",X"3E",X"01",X"32",X"8E",X"70",X"32",X"A1",X"70",X"2A",X"52",X"70",X"26",X"A0",
		X"22",X"52",X"70",X"AF",X"32",X"49",X"70",X"32",X"4A",X"70",X"C9",X"3E",X"01",X"32",X"51",X"70",
		X"3E",X"04",X"18",X"CF",X"16",X"00",X"5F",X"21",X"D1",X"08",X"19",X"7E",X"32",X"50",X"70",X"C9",
		X"DD",X"21",X"3F",X"70",X"3A",X"47",X"70",X"FE",X"10",X"30",X"18",X"CB",X"07",X"CB",X"07",X"CB",
		X"07",X"CB",X"07",X"DD",X"77",X"00",X"DD",X"36",X"01",X"00",X"DD",X"36",X"02",X"00",X"DD",X"36",
		X"03",X"01",X"C9",X"20",X"0A",X"DD",X"36",X"00",X"00",X"DD",X"36",X"01",X"01",X"18",X"EB",X"47",
		X"3E",X"20",X"90",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"DD",X"77",X"02",X"DD",X"36",
		X"00",X"00",X"DD",X"36",X"01",X"01",X"DD",X"36",X"03",X"00",X"C9",X"21",X"48",X"70",X"3A",X"46",
		X"70",X"FE",X"D6",X"28",X"64",X"FE",X"23",X"28",X"0E",X"3A",X"44",X"70",X"FE",X"0C",X"CA",X"38",
		X"0B",X"FE",X"F4",X"CA",X"54",X"0B",X"C9",X"CD",X"70",X"0B",X"3A",X"44",X"70",X"FE",X"7C",X"38",
		X"0D",X"3A",X"49",X"70",X"3C",X"32",X"49",X"70",X"AF",X"32",X"4A",X"70",X"18",X"0B",X"3A",X"4A",
		X"70",X"3C",X"32",X"4A",X"70",X"AF",X"32",X"49",X"70",X"3A",X"4B",X"70",X"FE",X"07",X"30",X"10",
		X"B7",X"28",X"0D",X"3D",X"F5",X"CD",X"54",X"0A",X"F1",X"32",X"4B",X"70",X"21",X"45",X"70",X"34",
		X"3A",X"48",X"70",X"FE",X"04",X"20",X"07",X"3E",X"02",X"32",X"48",X"70",X"18",X"AB",X"FE",X"03",
		X"20",X"A7",X"3E",X"01",X"32",X"48",X"70",X"18",X"A0",X"CD",X"43",X"0A",X"CD",X"70",X"0B",X"3A",
		X"48",X"70",X"FE",X"02",X"20",X"07",X"3E",X"04",X"32",X"48",X"70",X"18",X"8C",X"FE",X"01",X"20",
		X"88",X"3E",X"03",X"32",X"48",X"70",X"18",X"81",X"CD",X"43",X"0A",X"CD",X"70",X"0B",X"3A",X"48",
		X"70",X"FE",X"03",X"20",X"06",X"3E",X"04",X"32",X"48",X"70",X"C9",X"FE",X"01",X"C0",X"3E",X"02",
		X"32",X"48",X"70",X"C9",X"CD",X"43",X"0A",X"CD",X"70",X"0B",X"3A",X"48",X"70",X"FE",X"02",X"20",
		X"06",X"3E",X"01",X"32",X"48",X"70",X"C9",X"FE",X"04",X"C0",X"3E",X"03",X"32",X"48",X"70",X"C9",
		X"3A",X"BA",X"70",X"B7",X"C0",X"3A",X"33",X"70",X"B7",X"C8",X"3E",X"06",X"32",X"BA",X"70",X"C9",
		X"3A",X"4F",X"70",X"3D",X"28",X"04",X"32",X"4F",X"70",X"C9",X"3A",X"50",X"70",X"32",X"4F",X"70",
		X"3A",X"48",X"70",X"FE",X"03",X"38",X"0B",X"3A",X"47",X"70",X"FE",X"1A",X"C8",X"3C",X"32",X"47",
		X"70",X"C9",X"3A",X"47",X"70",X"B7",X"28",X"05",X"3D",X"32",X"47",X"70",X"C9",X"3A",X"48",X"70",
		X"3C",X"3C",X"32",X"48",X"70",X"C9",X"3E",X"14",X"32",X"47",X"70",X"3E",X"0F",X"32",X"4B",X"70",
		X"3E",X"00",X"32",X"50",X"70",X"32",X"4F",X"70",X"3E",X"01",X"32",X"48",X"70",X"3E",X"80",X"32",
		X"44",X"70",X"3E",X"80",X"32",X"46",X"70",X"3E",X"10",X"32",X"00",X"98",X"3E",X"04",X"32",X"01",
		X"98",X"3E",X"01",X"32",X"87",X"70",X"CD",X"60",X"0A",X"C9",X"CD",X"7F",X"0D",X"CD",X"D2",X"0C",
		X"CD",X"80",X"0C",X"CD",X"4F",X"0D",X"3A",X"61",X"70",X"FE",X"0E",X"28",X"10",X"FE",X"0C",X"28",
		X"14",X"FE",X"0D",X"20",X"20",X"AF",X"32",X"67",X"70",X"3E",X"30",X"18",X"0E",X"AF",X"32",X"67",
		X"70",X"3E",X"32",X"18",X"06",X"AF",X"32",X"67",X"70",X"3E",X"29",X"32",X"58",X"70",X"3E",X"12",
		X"32",X"54",X"70",X"18",X"0A",X"87",X"C6",X"11",X"32",X"58",X"70",X"3C",X"32",X"54",X"70",X"3E",
		X"02",X"32",X"55",X"70",X"3E",X"04",X"32",X"59",X"70",X"3E",X"04",X"32",X"5D",X"70",X"21",X"5A",
		X"70",X"11",X"5E",X"70",X"7E",X"D6",X"11",X"12",X"13",X"23",X"7E",X"12",X"3A",X"6E",X"70",X"B7",
		X"28",X"1E",X"7E",X"11",X"1F",X"98",X"C6",X"0C",X"12",X"1B",X"2B",X"7E",X"D6",X"04",X"12",X"1B",
		X"3E",X"04",X"12",X"1B",X"21",X"7C",X"0C",X"3A",X"6E",X"70",X"4F",X"06",X"00",X"09",X"7E",X"12",
		X"21",X"54",X"70",X"11",X"04",X"98",X"01",X"0C",X"00",X"ED",X"B0",X"C9",X"00",X"2C",X"2B",X"2A",
		X"3A",X"61",X"70",X"FE",X"0F",X"38",X"04",X"AF",X"32",X"61",X"70",X"87",X"21",X"B4",X"0C",X"16",
		X"00",X"5F",X"19",X"DD",X"21",X"5A",X"70",X"11",X"56",X"70",X"CD",X"9D",X"0C",X"7E",X"CB",X"7F",
		X"20",X"09",X"DD",X"86",X"00",X"12",X"13",X"DD",X"23",X"23",X"C9",X"CB",X"BF",X"4F",X"DD",X"7E",
		X"00",X"91",X"18",X"F1",X"90",X"00",X"90",X"8C",X"8C",X"90",X"82",X"90",X"06",X"90",X"0C",X"8E",
		X"10",X"00",X"10",X"0A",X"0A",X"10",X"82",X"10",X"8A",X"0E",X"90",X"08",X"90",X"00",X"90",X"00",
		X"90",X"00",X"3A",X"63",X"70",X"B7",X"C8",X"21",X"5C",X"70",X"DD",X"21",X"5B",X"70",X"11",X"60",
		X"70",X"3A",X"62",X"70",X"B7",X"20",X"37",X"3A",X"6F",X"70",X"B7",X"20",X"06",X"DD",X"7E",X"00",
		X"FE",X"69",X"D0",X"1A",X"3C",X"12",X"47",X"3A",X"64",X"70",X"B8",X"D0",X"AF",X"12",X"3A",X"65",
		X"70",X"EE",X"01",X"32",X"65",X"70",X"20",X"04",X"DD",X"34",X"00",X"C9",X"3E",X"0F",X"BE",X"20",
		X"04",X"36",X"0B",X"18",X"01",X"34",X"DD",X"34",X"00",X"21",X"63",X"70",X"35",X"C9",X"DD",X"7E",
		X"00",X"FE",X"20",X"D8",X"1A",X"3C",X"12",X"47",X"3A",X"64",X"70",X"B8",X"D0",X"AF",X"12",X"3A",
		X"65",X"70",X"EE",X"01",X"32",X"65",X"70",X"20",X"04",X"DD",X"35",X"00",X"C9",X"3E",X"0B",X"BE",
		X"20",X"0A",X"36",X"0F",X"DD",X"35",X"00",X"21",X"63",X"70",X"35",X"C9",X"35",X"18",X"F5",X"3A",
		X"67",X"70",X"B7",X"C8",X"3A",X"68",X"70",X"21",X"69",X"70",X"BE",X"28",X"05",X"3C",X"32",X"68",
		X"70",X"C9",X"AF",X"32",X"68",X"70",X"21",X"61",X"70",X"56",X"3A",X"66",X"70",X"BA",X"20",X"05",
		X"AF",X"32",X"67",X"70",X"C9",X"3A",X"6D",X"70",X"B7",X"CA",X"AD",X"0D",X"C3",X"C9",X"0D",X"3A",
		X"6C",X"70",X"B7",X"C0",X"F3",X"06",X"0E",X"DF",X"79",X"2F",X"FB",X"21",X"63",X"70",X"11",X"61",
		X"70",X"CB",X"5F",X"C4",X"F2",X"0D",X"CB",X"67",X"C4",X"E2",X"0D",X"21",X"6A",X"70",X"5F",X"AE",
		X"73",X"A3",X"CB",X"6F",X"C4",X"AD",X"0D",X"CB",X"77",X"C4",X"C9",X"0D",X"C9",X"F5",X"AF",X"32",
		X"8C",X"70",X"3C",X"32",X"8B",X"70",X"3A",X"61",X"70",X"FE",X"0B",X"28",X"06",X"3C",X"32",X"61",
		X"70",X"F1",X"C9",X"AF",X"32",X"61",X"70",X"F1",X"C9",X"3E",X"01",X"32",X"8C",X"70",X"32",X"8B",
		X"70",X"3A",X"61",X"70",X"B7",X"28",X"05",X"3D",X"32",X"61",X"70",X"C9",X"3E",X"0B",X"32",X"61",
		X"70",X"C9",X"F5",X"3A",X"5B",X"70",X"FE",X"69",X"30",X"17",X"AF",X"32",X"62",X"70",X"36",X"01",
		X"F1",X"C9",X"F5",X"3A",X"5B",X"70",X"FE",X"20",X"38",X"07",X"3E",X"01",X"32",X"62",X"70",X"36",
		X"01",X"F1",X"C9",X"CD",X"A8",X"0F",X"CD",X"F3",X"0E",X"CD",X"A1",X"0E",X"CD",X"78",X"0F",X"3A",
		X"7D",X"70",X"FE",X"0E",X"28",X"10",X"FE",X"0C",X"28",X"14",X"FE",X"0D",X"20",X"24",X"AF",X"32",
		X"83",X"70",X"3E",X"30",X"18",X"0E",X"AF",X"32",X"83",X"70",X"3E",X"32",X"18",X"06",X"AF",X"32",
		X"83",X"70",X"3E",X"29",X"CB",X"F7",X"32",X"74",X"70",X"3E",X"12",X"CB",X"F7",X"32",X"70",X"70",
		X"18",X"0C",X"87",X"C6",X"11",X"CB",X"F7",X"32",X"74",X"70",X"3C",X"32",X"70",X"70",X"3E",X"02",
		X"32",X"71",X"70",X"3E",X"01",X"32",X"75",X"70",X"3E",X"01",X"32",X"79",X"70",X"21",X"76",X"70",
		X"11",X"7A",X"70",X"7E",X"D6",X"10",X"12",X"13",X"23",X"7E",X"12",X"3A",X"89",X"70",X"B7",X"28",
		X"20",X"7E",X"11",X"1F",X"98",X"D6",X"0A",X"12",X"1B",X"2B",X"7E",X"D6",X"04",X"12",X"1B",X"3E",
		X"04",X"12",X"1B",X"21",X"9D",X"0E",X"3A",X"89",X"70",X"4F",X"06",X"00",X"09",X"7E",X"CB",X"F7",
		X"12",X"21",X"70",X"70",X"11",X"10",X"98",X"01",X"0C",X"00",X"ED",X"B0",X"C9",X"00",X"2C",X"2B",
		X"2A",X"3A",X"7D",X"70",X"FE",X"0F",X"38",X"04",X"AF",X"32",X"7D",X"70",X"87",X"21",X"D5",X"0E",
		X"16",X"00",X"5F",X"19",X"DD",X"21",X"76",X"70",X"11",X"72",X"70",X"CD",X"BE",X"0E",X"7E",X"CB",
		X"7F",X"20",X"09",X"DD",X"86",X"00",X"12",X"13",X"DD",X"23",X"23",X"C9",X"CB",X"BF",X"4F",X"DD",
		X"7E",X"00",X"91",X"18",X"F1",X"90",X"00",X"90",X"0C",X"8C",X"10",X"82",X"10",X"06",X"10",X"0C",
		X"0E",X"10",X"00",X"10",X"8A",X"0A",X"90",X"82",X"90",X"8A",X"8E",X"90",X"88",X"90",X"00",X"90",
		X"00",X"90",X"00",X"3A",X"7F",X"70",X"B7",X"C8",X"21",X"78",X"70",X"DD",X"21",X"77",X"70",X"11",
		X"7C",X"70",X"3A",X"7E",X"70",X"B7",X"20",X"35",X"DD",X"7E",X"00",X"FE",X"D7",X"D0",X"1A",X"3C",
		X"12",X"47",X"3A",X"80",X"70",X"B8",X"D0",X"AF",X"12",X"3A",X"81",X"70",X"EE",X"01",X"32",X"81",
		X"70",X"20",X"04",X"DD",X"34",X"00",X"C9",X"3E",X"0B",X"CB",X"F7",X"BE",X"20",X"04",X"36",X"0F",
		X"18",X"01",X"35",X"DD",X"34",X"00",X"CB",X"F6",X"21",X"7F",X"70",X"35",X"C9",X"3A",X"6F",X"70",
		X"B7",X"20",X"06",X"DD",X"7E",X"00",X"FE",X"8D",X"D8",X"1A",X"3C",X"12",X"47",X"3A",X"80",X"70",
		X"B8",X"D0",X"AF",X"12",X"3A",X"81",X"70",X"EE",X"01",X"32",X"81",X"70",X"20",X"04",X"DD",X"35",
		X"00",X"C9",X"3E",X"0F",X"CB",X"F7",X"BE",X"20",X"0C",X"36",X"0B",X"DD",X"35",X"00",X"CB",X"F6",
		X"21",X"7F",X"70",X"35",X"C9",X"34",X"18",X"F3",X"3A",X"83",X"70",X"B7",X"C8",X"3A",X"84",X"70",
		X"21",X"85",X"70",X"BE",X"28",X"05",X"3C",X"32",X"84",X"70",X"C9",X"AF",X"32",X"84",X"70",X"21",
		X"7D",X"70",X"3A",X"82",X"70",X"56",X"BA",X"20",X"05",X"AF",X"32",X"83",X"70",X"C9",X"3A",X"88",
		X"70",X"B7",X"CA",X"D6",X"0F",X"C3",X"F2",X"0F",X"3A",X"87",X"70",X"B7",X"C0",X"F3",X"06",X"0F",
		X"DF",X"79",X"2F",X"FB",X"21",X"7F",X"70",X"11",X"7D",X"70",X"CB",X"5F",X"C4",X"1B",X"10",X"CB",
		X"67",X"C4",X"0B",X"10",X"21",X"86",X"70",X"5F",X"AE",X"73",X"A3",X"CB",X"6F",X"C4",X"D6",X"0F",
		X"CB",X"77",X"C4",X"F2",X"0F",X"C9",X"F5",X"AF",X"32",X"92",X"70",X"3C",X"32",X"91",X"70",X"3A",
		X"7D",X"70",X"FE",X"0B",X"28",X"06",X"3C",X"32",X"7D",X"70",X"F1",X"C9",X"AF",X"32",X"7D",X"70",
		X"F1",X"C9",X"3E",X"01",X"32",X"92",X"70",X"32",X"91",X"70",X"3A",X"7D",X"70",X"B7",X"28",X"05",
		X"3D",X"32",X"7D",X"70",X"C9",X"3E",X"0B",X"32",X"7D",X"70",X"C9",X"F5",X"3A",X"77",X"70",X"FE",
		X"E0",X"30",X"17",X"AF",X"32",X"7E",X"70",X"36",X"01",X"F1",X"C9",X"F5",X"3A",X"77",X"70",X"FE",
		X"85",X"38",X"07",X"3E",X"01",X"32",X"7E",X"70",X"36",X"01",X"F1",X"C9",X"3A",X"8D",X"70",X"B7",
		X"28",X"05",X"3D",X"32",X"8D",X"70",X"C9",X"3A",X"8E",X"70",X"B7",X"C0",X"3A",X"8B",X"70",X"B7",
		X"28",X"0E",X"CD",X"27",X"11",X"B7",X"C4",X"2A",X"12",X"AF",X"32",X"8B",X"70",X"C3",X"9F",X"10",
		X"3A",X"63",X"70",X"B7",X"20",X"EC",X"CD",X"60",X"10",X"B7",X"C4",X"74",X"11",X"C3",X"9F",X"10",
		X"DD",X"21",X"D3",X"12",X"3A",X"61",X"70",X"CB",X"27",X"CB",X"27",X"16",X"00",X"5F",X"DD",X"19",
		X"21",X"46",X"70",X"3A",X"56",X"70",X"DD",X"86",X"00",X"BE",X"38",X"21",X"3A",X"56",X"70",X"DD",
		X"96",X"01",X"BE",X"30",X"18",X"3A",X"57",X"70",X"21",X"44",X"70",X"DD",X"86",X"03",X"BE",X"38",
		X"0C",X"3A",X"57",X"70",X"DD",X"96",X"02",X"BE",X"30",X"03",X"3E",X"01",X"C9",X"AF",X"C9",X"DD",
		X"21",X"1F",X"11",X"CD",X"BC",X"10",X"32",X"8F",X"70",X"B7",X"20",X"3F",X"3A",X"3C",X"70",X"B7",
		X"C8",X"DD",X"21",X"23",X"11",X"CD",X"BC",X"10",X"B7",X"20",X"40",X"C9",X"21",X"46",X"70",X"3A",
		X"5A",X"70",X"DD",X"86",X"00",X"BE",X"38",X"21",X"3A",X"5A",X"70",X"DD",X"96",X"01",X"BE",X"30",
		X"18",X"3A",X"5B",X"70",X"21",X"44",X"70",X"DD",X"86",X"03",X"BE",X"38",X"0C",X"3A",X"5B",X"70",
		X"DD",X"96",X"02",X"BE",X"30",X"03",X"3E",X"01",X"C9",X"AF",X"C9",X"3E",X"0F",X"32",X"2B",X"70",
		X"3A",X"33",X"70",X"B7",X"28",X"05",X"3E",X"08",X"32",X"BA",X"70",X"3E",X"00",X"32",X"4B",X"70",
		X"3E",X"03",X"32",X"48",X"70",X"3E",X"1E",X"32",X"47",X"70",X"3E",X"01",X"32",X"8E",X"70",X"32",
		X"A1",X"70",X"AF",X"32",X"51",X"70",X"3E",X"0E",X"32",X"B5",X"70",X"CD",X"76",X"18",X"C9",X"08",
		X"02",X"06",X"06",X"00",X"0D",X"06",X"06",X"3A",X"8C",X"70",X"B7",X"3A",X"61",X"70",X"20",X"06",
		X"B7",X"20",X"02",X"3E",X"0C",X"3D",X"CB",X"27",X"CB",X"27",X"DD",X"21",X"A3",X"12",X"16",X"00",
		X"5F",X"DD",X"19",X"3A",X"5A",X"70",X"D6",X"19",X"DD",X"86",X"00",X"08",X"3A",X"5B",X"70",X"D6",
		X"19",X"DD",X"86",X"01",X"21",X"44",X"70",X"BE",X"D2",X"9D",X"10",X"DD",X"86",X"02",X"BE",X"DA",
		X"9D",X"10",X"21",X"46",X"70",X"08",X"BE",X"DA",X"9D",X"10",X"DD",X"96",X"03",X"BE",X"D2",X"9D",
		X"10",X"3E",X"01",X"C9",X"CD",X"B7",X"11",X"3A",X"61",X"70",X"FE",X"00",X"CA",X"02",X"12",X"FE",
		X"01",X"CA",X"C7",X"11",X"FE",X"02",X"CA",X"C7",X"11",X"FE",X"03",X"CA",X"13",X"12",X"FE",X"04",
		X"CA",X"ED",X"11",X"FE",X"05",X"CA",X"ED",X"11",X"FE",X"06",X"CA",X"02",X"12",X"FE",X"07",X"CA",
		X"C7",X"11",X"FE",X"08",X"CA",X"C7",X"11",X"FE",X"09",X"CA",X"13",X"12",X"FE",X"0A",X"CA",X"ED",
		X"11",X"FE",X"0B",X"CA",X"ED",X"11",X"C9",X"3A",X"33",X"70",X"B7",X"C8",X"3A",X"BA",X"70",X"B7",
		X"C0",X"3E",X"05",X"32",X"BA",X"70",X"C9",X"3A",X"48",X"70",X"FE",X"04",X"28",X"06",X"FE",X"01",
		X"28",X"06",X"18",X"09",X"3E",X"01",X"18",X"02",X"3E",X"04",X"32",X"48",X"70",X"3A",X"47",X"70",
		X"4F",X"3E",X"20",X"91",X"32",X"47",X"70",X"3E",X"80",X"32",X"8D",X"70",X"C9",X"3A",X"48",X"70",
		X"FE",X"03",X"28",X"06",X"FE",X"02",X"28",X"06",X"18",X"E3",X"3E",X"02",X"18",X"DC",X"3E",X"03",
		X"18",X"D8",X"3A",X"48",X"70",X"FE",X"01",X"28",X"14",X"FE",X"02",X"28",X"17",X"FE",X"03",X"28",
		X"0C",X"18",X"11",X"3A",X"48",X"70",X"FE",X"03",X"38",X"02",X"18",X"07",X"3C",X"3C",X"32",X"48",
		X"70",X"18",X"C4",X"3D",X"3D",X"32",X"48",X"70",X"18",X"BD",X"CD",X"B7",X"11",X"DD",X"21",X"73",
		X"12",X"3A",X"61",X"70",X"CB",X"27",X"CB",X"27",X"16",X"00",X"5F",X"DD",X"19",X"DD",X"7E",X"01",
		X"32",X"47",X"70",X"3A",X"8C",X"70",X"B7",X"20",X"25",X"DD",X"7E",X"00",X"32",X"48",X"70",X"3E",
		X"80",X"32",X"8D",X"70",X"3A",X"0E",X"70",X"C6",X"05",X"FE",X"0E",X"30",X"08",X"FE",X"05",X"30",
		X"06",X"3E",X"05",X"18",X"02",X"3E",X"0F",X"32",X"4B",X"70",X"CD",X"54",X"0A",X"C9",X"DD",X"7E",
		X"02",X"18",X"D9",X"01",X"0A",X"04",X"00",X"01",X"14",X"04",X"00",X"01",X"1E",X"04",X"00",X"02",
		X"14",X"03",X"00",X"02",X"0A",X"03",X"00",X"02",X"05",X"03",X"00",X"04",X"00",X"01",X"00",X"04",
		X"00",X"01",X"00",X"04",X"0A",X"01",X"00",X"03",X"14",X"02",X"00",X"03",X"0A",X"02",X"00",X"01",
		X"05",X"02",X"00",X"0F",X"0D",X"0F",X"0F",X"11",X"01",X"12",X"11",X"1B",X"00",X"14",X"10",X"25",
		X"00",X"14",X"11",X"2F",X"00",X"14",X"11",X"31",X"08",X"15",X"11",X"31",X"14",X"12",X"11",X"31",
		X"1E",X"13",X"13",X"25",X"1F",X"14",X"14",X"19",X"1E",X"15",X"13",X"11",X"1C",X"15",X"12",X"11",
		X"14",X"0F",X"12",X"00",X"08",X"08",X"04",X"02",X"07",X"06",X"04",X"04",X"06",X"05",X"04",X"05",
		X"06",X"0A",X"02",X"09",X"03",X"0A",X"03",X"08",X"03",X"01",X"08",X"09",X"02",X"05",X"03",X"06",
		X"04",X"04",X"05",X"05",X"05",X"09",X"02",X"04",X"07",X"06",X"09",X"01",X"09",X"06",X"06",X"01",
		X"09",X"04",X"06",X"3A",X"93",X"70",X"B7",X"28",X"05",X"3D",X"32",X"93",X"70",X"C9",X"3A",X"8E",
		X"70",X"B7",X"C0",X"3A",X"91",X"70",X"B7",X"28",X"0E",X"CD",X"FA",X"13",X"B7",X"C4",X"ED",X"14",
		X"AF",X"32",X"91",X"70",X"C3",X"76",X"13",X"3A",X"7F",X"70",X"B7",X"20",X"EC",X"CD",X"37",X"13",
		X"B7",X"C4",X"47",X"14",X"C3",X"76",X"13",X"DD",X"21",X"96",X"15",X"3A",X"7D",X"70",X"CB",X"27",
		X"CB",X"27",X"16",X"00",X"5F",X"DD",X"19",X"21",X"46",X"70",X"3A",X"72",X"70",X"DD",X"86",X"00",
		X"BE",X"38",X"21",X"3A",X"72",X"70",X"DD",X"96",X"01",X"BE",X"30",X"18",X"3A",X"73",X"70",X"21",
		X"44",X"70",X"DD",X"86",X"03",X"BE",X"38",X"0C",X"3A",X"73",X"70",X"DD",X"96",X"02",X"BE",X"30",
		X"03",X"3E",X"01",X"C9",X"AF",X"C9",X"DD",X"21",X"F2",X"13",X"CD",X"90",X"13",X"B7",X"20",X"3F",
		X"3A",X"3C",X"70",X"B7",X"C8",X"DD",X"21",X"F6",X"13",X"CD",X"90",X"13",X"B7",X"20",X"40",X"C9",
		X"21",X"46",X"70",X"3A",X"76",X"70",X"DD",X"86",X"00",X"BE",X"38",X"21",X"3A",X"76",X"70",X"DD",
		X"96",X"01",X"BE",X"30",X"18",X"3A",X"77",X"70",X"21",X"44",X"70",X"DD",X"86",X"03",X"BE",X"38",
		X"0C",X"3A",X"77",X"70",X"DD",X"96",X"02",X"BE",X"30",X"03",X"3E",X"01",X"C9",X"AF",X"C9",X"3E",
		X"0F",X"32",X"2E",X"70",X"3A",X"33",X"70",X"B7",X"28",X"05",X"3E",X"08",X"32",X"BA",X"70",X"3E",
		X"00",X"32",X"4B",X"70",X"3E",X"04",X"32",X"48",X"70",X"3E",X"1C",X"32",X"47",X"70",X"3E",X"01",
		X"32",X"8E",X"70",X"32",X"A1",X"70",X"32",X"51",X"70",X"3E",X"0E",X"32",X"B5",X"70",X"CD",X"76",
		X"18",X"C9",X"08",X"02",X"06",X"06",X"00",X"0D",X"06",X"06",X"3A",X"92",X"70",X"B7",X"3A",X"7D",
		X"70",X"20",X"06",X"B7",X"20",X"02",X"3E",X"0C",X"3D",X"CB",X"27",X"CB",X"27",X"DD",X"21",X"66",
		X"15",X"16",X"00",X"5F",X"DD",X"19",X"3A",X"76",X"70",X"D6",X"19",X"DD",X"86",X"00",X"08",X"3A",
		X"77",X"70",X"C6",X"19",X"DD",X"96",X"01",X"21",X"44",X"70",X"BE",X"DA",X"74",X"13",X"DD",X"96",
		X"02",X"BE",X"D2",X"74",X"13",X"21",X"46",X"70",X"08",X"BE",X"DA",X"74",X"13",X"DD",X"96",X"03",
		X"BE",X"D2",X"74",X"13",X"3E",X"01",X"C9",X"CD",X"B7",X"11",X"3A",X"7D",X"70",X"FE",X"00",X"CA",
		X"C5",X"14",X"FE",X"01",X"CA",X"B0",X"14",X"FE",X"02",X"CA",X"B0",X"14",X"FE",X"03",X"CA",X"D6",
		X"14",X"FE",X"04",X"CA",X"8A",X"14",X"FE",X"05",X"CA",X"8A",X"14",X"FE",X"06",X"CA",X"C5",X"14",
		X"FE",X"07",X"CA",X"B0",X"14",X"FE",X"08",X"CA",X"B0",X"14",X"FE",X"09",X"CA",X"D6",X"14",X"FE",
		X"0A",X"CA",X"8A",X"14",X"FE",X"0B",X"CA",X"8A",X"14",X"C9",X"3A",X"48",X"70",X"FE",X"04",X"28",
		X"06",X"FE",X"01",X"28",X"06",X"18",X"09",X"3E",X"01",X"18",X"02",X"3E",X"04",X"32",X"48",X"70",
		X"3A",X"47",X"70",X"4F",X"3E",X"20",X"91",X"32",X"47",X"70",X"3E",X"80",X"32",X"93",X"70",X"C9",
		X"3A",X"48",X"70",X"FE",X"03",X"28",X"06",X"FE",X"02",X"28",X"06",X"18",X"E3",X"3E",X"02",X"18",
		X"DC",X"3E",X"03",X"18",X"D8",X"3A",X"48",X"70",X"FE",X"01",X"28",X"14",X"FE",X"02",X"28",X"17",
		X"FE",X"03",X"28",X"0C",X"18",X"11",X"3A",X"48",X"70",X"FE",X"03",X"38",X"02",X"18",X"07",X"3C",
		X"3C",X"32",X"48",X"70",X"18",X"C4",X"3D",X"3D",X"32",X"48",X"70",X"18",X"BD",X"CD",X"B7",X"11",
		X"DD",X"21",X"36",X"15",X"3A",X"7D",X"70",X"CB",X"27",X"CB",X"27",X"16",X"00",X"5F",X"DD",X"19",
		X"DD",X"7E",X"01",X"32",X"47",X"70",X"3A",X"92",X"70",X"B7",X"28",X"25",X"DD",X"7E",X"02",X"32",
		X"48",X"70",X"3E",X"80",X"32",X"93",X"70",X"3A",X"0F",X"70",X"C6",X"05",X"FE",X"0E",X"30",X"08",
		X"FE",X"05",X"30",X"06",X"3E",X"05",X"18",X"02",X"3E",X"0F",X"32",X"4B",X"70",X"CD",X"54",X"0A",
		X"C9",X"DD",X"7E",X"00",X"18",X"D9",X"02",X"0A",X"03",X"00",X"02",X"14",X"03",X"00",X"02",X"1E",
		X"03",X"00",X"01",X"14",X"04",X"00",X"01",X"0A",X"04",X"00",X"01",X"05",X"04",X"00",X"03",X"00",
		X"02",X"00",X"03",X"00",X"02",X"00",X"03",X"0A",X"02",X"00",X"04",X"14",X"01",X"00",X"04",X"0A",
		X"01",X"00",X"02",X"05",X"01",X"00",X"0F",X"0D",X"0F",X"0F",X"11",X"01",X"12",X"11",X"1B",X"00",
		X"14",X"10",X"25",X"00",X"14",X"11",X"2F",X"00",X"14",X"11",X"31",X"08",X"15",X"11",X"31",X"14",
		X"12",X"11",X"31",X"1E",X"13",X"13",X"25",X"1F",X"14",X"14",X"19",X"1E",X"15",X"13",X"11",X"1C",
		X"15",X"12",X"11",X"14",X"0F",X"12",X"00",X"08",X"08",X"04",X"02",X"07",X"06",X"04",X"04",X"06",
		X"05",X"04",X"05",X"06",X"0A",X"02",X"09",X"03",X"0A",X"03",X"08",X"03",X"01",X"08",X"09",X"02",
		X"05",X"03",X"06",X"04",X"04",X"05",X"05",X"05",X"09",X"02",X"04",X"07",X"06",X"09",X"01",X"09",
		X"06",X"06",X"01",X"09",X"04",X"06",X"CD",X"F6",X"16",X"3A",X"95",X"70",X"B7",X"28",X"05",X"3D",
		X"32",X"95",X"70",X"C9",X"3A",X"44",X"70",X"FE",X"7C",X"DA",X"17",X"16",X"CD",X"7C",X"16",X"FE",
		X"FF",X"28",X"34",X"F5",X"FE",X"05",X"20",X"07",X"3E",X"01",X"32",X"2A",X"70",X"18",X"04",X"FE",
		X"06",X"28",X"F5",X"F1",X"CB",X"27",X"21",X"5B",X"17",X"16",X"00",X"5F",X"19",X"7E",X"32",X"82",
		X"70",X"23",X"7E",X"32",X"88",X"70",X"3E",X"30",X"32",X"95",X"70",X"3A",X"98",X"70",X"32",X"85",
		X"70",X"3E",X"01",X"32",X"83",X"70",X"C9",X"3A",X"46",X"70",X"FE",X"80",X"30",X"11",X"3A",X"97",
		X"70",X"B7",X"20",X"08",X"3A",X"44",X"70",X"FE",X"60",X"DA",X"2F",X"16",X"C3",X"4A",X"16",X"3A",
		X"77",X"70",X"FE",X"B0",X"38",X"05",X"FE",X"B2",X"D8",X"18",X"0B",X"AF",X"32",X"7E",X"70",X"3E",
		X"01",X"32",X"7F",X"70",X"18",X"10",X"3E",X"01",X"18",X"F2",X"3A",X"44",X"70",X"21",X"77",X"70",
		X"BE",X"C8",X"38",X"F2",X"18",X"E5",X"3A",X"44",X"70",X"FE",X"40",X"38",X"0E",X"FE",X"60",X"38",
		X"05",X"3A",X"99",X"70",X"18",X"08",X"3A",X"9A",X"70",X"18",X"03",X"3A",X"9B",X"70",X"32",X"80",
		X"70",X"3E",X"02",X"32",X"82",X"70",X"3E",X"01",X"32",X"83",X"70",X"C9",X"21",X"44",X"70",X"3A",
		X"77",X"70",X"D6",X"19",X"BE",X"D2",X"B3",X"16",X"C6",X"32",X"BE",X"DA",X"B3",X"16",X"21",X"46",
		X"70",X"3A",X"76",X"70",X"C6",X"19",X"BE",X"DA",X"B3",X"16",X"D6",X"32",X"BE",X"D2",X"B3",X"16",
		X"AF",X"06",X"0C",X"C5",X"F5",X"CD",X"B6",X"16",X"B7",X"28",X"03",X"F1",X"C1",X"C9",X"F1",X"C1",
		X"3C",X"10",X"F0",X"3E",X"FF",X"C9",X"CB",X"27",X"CB",X"27",X"DD",X"21",X"2B",X"17",X"16",X"00",
		X"5F",X"DD",X"19",X"3A",X"76",X"70",X"D6",X"19",X"DD",X"86",X"00",X"08",X"3A",X"77",X"70",X"C6",
		X"19",X"DD",X"96",X"01",X"21",X"44",X"70",X"BE",X"DA",X"F4",X"16",X"DD",X"96",X"02",X"BE",X"D2",
		X"F4",X"16",X"21",X"46",X"70",X"08",X"BE",X"DA",X"F4",X"16",X"DD",X"96",X"03",X"BE",X"D2",X"F4",
		X"16",X"3E",X"01",X"C9",X"AF",X"C9",X"3A",X"96",X"70",X"08",X"3A",X"13",X"70",X"47",X"3A",X"12",
		X"70",X"90",X"FE",X"03",X"38",X"22",X"08",X"3C",X"08",X"FE",X"06",X"38",X"1B",X"08",X"3C",X"CB",
		X"27",X"CB",X"27",X"CB",X"27",X"21",X"73",X"17",X"16",X"00",X"5F",X"19",X"11",X"97",X"70",X"06",
		X"07",X"7E",X"12",X"23",X"13",X"10",X"FA",X"C9",X"08",X"18",X"E4",X"0F",X"0D",X"0F",X"0F",X"11",
		X"01",X"12",X"11",X"1B",X"00",X"14",X"10",X"25",X"00",X"14",X"11",X"2F",X"00",X"14",X"11",X"31",
		X"08",X"15",X"11",X"31",X"14",X"12",X"11",X"31",X"1E",X"13",X"13",X"25",X"1F",X"14",X"14",X"19",
		X"1E",X"15",X"13",X"11",X"1C",X"15",X"12",X"11",X"14",X"0F",X"12",X"02",X"00",X"03",X"00",X"04",
		X"00",X"05",X"00",X"06",X"00",X"07",X"00",X"08",X"00",X"06",X"01",X"06",X"01",X"08",X"01",X"09",
		X"01",X"0A",X"01",X"00",X"02",X"02",X"03",X"04",X"90",X"80",X"00",X"00",X"02",X"02",X"02",X"04",
		X"B0",X"80",X"00",X"00",X"02",X"02",X"02",X"03",X"C0",X"80",X"00",X"00",X"02",X"02",X"02",X"03",
		X"FF",X"70",X"00",X"00",X"01",X"01",X"02",X"02",X"FF",X"60",X"00",X"00",X"01",X"01",X"02",X"02",
		X"FF",X"60",X"00",X"3A",X"4B",X"70",X"B7",X"C4",X"E1",X"08",X"3A",X"B4",X"70",X"FE",X"01",X"20",
		X"05",X"CD",X"36",X"18",X"18",X"05",X"FE",X"02",X"CC",X"3F",X"18",X"3A",X"A1",X"70",X"FE",X"00",
		X"28",X"12",X"FE",X"01",X"CA",X"2B",X"19",X"FE",X"02",X"CA",X"55",X"18",X"FE",X"03",X"CA",X"21",
		X"19",X"C3",X"03",X"19",X"CD",X"2C",X"10",X"CD",X"03",X"13",X"3A",X"33",X"70",X"B7",X"20",X"10",
		X"3E",X"01",X"32",X"6C",X"70",X"32",X"87",X"70",X"CD",X"C6",X"15",X"CD",X"67",X"22",X"18",X"14",
		X"FE",X"01",X"C2",X"27",X"18",X"3E",X"01",X"32",X"87",X"70",X"AF",X"32",X"AE",X"70",X"32",X"6C",
		X"70",X"CD",X"C6",X"15",X"21",X"00",X"02",X"22",X"A2",X"70",X"01",X"00",X"04",X"ED",X"43",X"A4",
		X"70",X"01",X"00",X"02",X"ED",X"43",X"A6",X"70",X"3E",X"09",X"32",X"AD",X"70",X"CD",X"D1",X"09",
		X"3A",X"A0",X"70",X"C2",X"21",X"19",X"C9",X"AF",X"32",X"6C",X"70",X"32",X"87",X"70",X"3E",X"01",
		X"32",X"AE",X"70",X"C3",X"04",X"18",X"3A",X"BA",X"70",X"B7",X"C0",X"3E",X"04",X"18",X"07",X"3A",
		X"BA",X"70",X"B7",X"C0",X"3E",X"03",X"08",X"3A",X"33",X"70",X"B7",X"C8",X"08",X"32",X"BA",X"70",
		X"AF",X"32",X"B4",X"70",X"C9",X"CD",X"2B",X"1A",X"ED",X"5B",X"A2",X"70",X"7A",X"B3",X"28",X"06",
		X"1B",X"ED",X"53",X"A2",X"70",X"C9",X"3A",X"F2",X"70",X"B7",X"C0",X"3E",X"03",X"32",X"A1",X"70",
		X"3E",X"01",X"32",X"A0",X"70",X"C9",X"3A",X"51",X"70",X"B7",X"28",X"16",X"3A",X"B2",X"70",X"FE",
		X"01",X"CA",X"AC",X"18",X"3A",X"B0",X"70",X"3C",X"FE",X"03",X"CA",X"AC",X"18",X"32",X"B0",X"70",
		X"18",X"14",X"3A",X"B3",X"70",X"FE",X"01",X"CA",X"BB",X"18",X"3A",X"B1",X"70",X"3C",X"FE",X"03",
		X"CA",X"BB",X"18",X"32",X"B1",X"70",X"3E",X"01",X"32",X"B4",X"70",X"C9",X"21",X"12",X"70",X"3E",
		X"01",X"32",X"37",X"70",X"3E",X"04",X"32",X"26",X"70",X"18",X"0D",X"21",X"13",X"70",X"3E",X"01",
		X"32",X"3A",X"70",X"3E",X"04",X"32",X"2A",X"70",X"34",X"AF",X"32",X"B0",X"70",X"32",X"B1",X"70",
		X"32",X"B2",X"70",X"32",X"B3",X"70",X"3E",X"02",X"32",X"B4",X"70",X"3A",X"AA",X"70",X"B7",X"28",
		X"10",X"3A",X"AB",X"70",X"3C",X"FE",X"03",X"20",X"04",X"AF",X"32",X"AA",X"70",X"32",X"AB",X"70",
		X"C9",X"3A",X"AC",X"70",X"3C",X"FE",X"03",X"20",X"06",X"3E",X"01",X"32",X"AA",X"70",X"AF",X"32",
		X"AC",X"70",X"C9",X"CD",X"2B",X"1A",X"ED",X"5B",X"A2",X"70",X"7A",X"B3",X"28",X"06",X"1B",X"ED",
		X"53",X"A2",X"70",X"C9",X"3E",X"01",X"32",X"AF",X"70",X"AF",X"32",X"37",X"70",X"32",X"3A",X"70",
		X"C9",X"3A",X"AA",X"70",X"B7",X"CA",X"84",X"1A",X"C3",X"95",X"1B",X"3A",X"19",X"70",X"21",X"12",
		X"70",X"BE",X"CA",X"DB",X"19",X"21",X"13",X"70",X"BE",X"CA",X"EC",X"19",X"ED",X"4B",X"A4",X"70",
		X"78",X"B1",X"28",X"60",X"0B",X"ED",X"43",X"A4",X"70",X"3A",X"44",X"70",X"FE",X"7C",X"30",X"09",
		X"FE",X"0F",X"38",X"05",X"3E",X"01",X"32",X"F2",X"70",X"3A",X"4B",X"70",X"B7",X"20",X"38",X"3A",
		X"AD",X"70",X"3D",X"28",X"05",X"32",X"AD",X"70",X"18",X"2D",X"3E",X"09",X"32",X"AD",X"70",X"3A",
		X"B5",X"70",X"B7",X"28",X"06",X"3D",X"32",X"B5",X"70",X"18",X"1C",X"3A",X"46",X"70",X"FE",X"13",
		X"28",X"09",X"3D",X"32",X"46",X"70",X"32",X"02",X"98",X"18",X"0C",X"3A",X"44",X"70",X"FE",X"0F",
		X"38",X"05",X"3E",X"01",X"32",X"F2",X"70",X"3A",X"2B",X"70",X"B7",X"C0",X"3A",X"2E",X"70",X"B7",
		X"C0",X"3E",X"01",X"C9",X"3A",X"51",X"70",X"B7",X"28",X"0C",X"3E",X"0D",X"32",X"7D",X"70",X"3E",
		X"0C",X"32",X"61",X"70",X"18",X"0A",X"3E",X"0C",X"32",X"7D",X"70",X"3E",X"0D",X"32",X"61",X"70",
		X"ED",X"4B",X"A6",X"70",X"78",X"B1",X"28",X"06",X"0B",X"ED",X"43",X"A6",X"70",X"C9",X"3E",X"02",
		X"32",X"A1",X"70",X"AF",X"32",X"7D",X"70",X"32",X"61",X"70",X"C9",X"3E",X"06",X"32",X"61",X"70",
		X"3E",X"0A",X"32",X"26",X"70",X"3E",X"0D",X"32",X"7D",X"70",X"18",X"0F",X"3E",X"06",X"32",X"7D",
		X"70",X"3E",X"0A",X"32",X"2A",X"70",X"3E",X"0D",X"32",X"61",X"70",X"3E",X"04",X"32",X"A1",X"70",
		X"3E",X"01",X"32",X"6C",X"70",X"32",X"87",X"70",X"3E",X"02",X"32",X"BA",X"70",X"3E",X"01",X"32",
		X"4B",X"70",X"AF",X"32",X"B4",X"70",X"21",X"2C",X"02",X"22",X"F5",X"70",X"3E",X"05",X"32",X"F7",
		X"70",X"CD",X"D6",X"23",X"21",X"00",X"09",X"22",X"A2",X"70",X"C9",X"3A",X"AA",X"70",X"B7",X"20",
		X"2B",X"3E",X"05",X"32",X"64",X"70",X"3E",X"01",X"32",X"6C",X"70",X"01",X"01",X"00",X"ED",X"43",
		X"9E",X"70",X"3A",X"5B",X"70",X"FE",X"30",X"38",X"03",X"FE",X"32",X"D8",X"3E",X"01",X"32",X"63",
		X"70",X"38",X"04",X"32",X"62",X"70",X"C9",X"AF",X"32",X"62",X"70",X"C9",X"3E",X"05",X"32",X"80",
		X"70",X"3E",X"01",X"32",X"87",X"70",X"3A",X"77",X"70",X"FE",X"C7",X"C8",X"38",X"0C",X"FE",X"CA",
		X"D8",X"3E",X"01",X"32",X"7F",X"70",X"32",X"7E",X"70",X"C9",X"AF",X"32",X"7E",X"70",X"3E",X"01",
		X"32",X"7F",X"70",X"C9",X"ED",X"4B",X"9E",X"70",X"0B",X"ED",X"43",X"9E",X"70",X"78",X"B1",X"C0",
		X"3A",X"A0",X"70",X"FE",X"01",X"CA",X"DA",X"1A",X"FE",X"02",X"CA",X"FB",X"1A",X"FE",X"03",X"CA",
		X"06",X"1B",X"FE",X"04",X"CA",X"16",X"1B",X"FE",X"05",X"CA",X"31",X"1B",X"FE",X"06",X"CA",X"4C",
		X"1B",X"21",X"90",X"00",X"22",X"9E",X"70",X"21",X"A0",X"70",X"36",X"00",X"AF",X"32",X"1F",X"98",
		X"32",X"1E",X"98",X"32",X"6E",X"70",X"32",X"89",X"70",X"32",X"37",X"70",X"32",X"3A",X"70",X"3E",
		X"03",X"32",X"1A",X"70",X"3E",X"05",X"32",X"1B",X"70",X"C9",X"3A",X"33",X"70",X"FE",X"02",X"20",
		X"04",X"AF",X"32",X"87",X"70",X"3A",X"33",X"70",X"B7",X"28",X"05",X"3E",X"01",X"32",X"1A",X"70",
		X"3E",X"02",X"32",X"89",X"70",X"21",X"18",X"00",X"C3",X"8D",X"1B",X"3E",X"03",X"32",X"89",X"70",
		X"21",X"90",X"00",X"C3",X"8D",X"1B",X"AF",X"32",X"89",X"70",X"32",X"1F",X"98",X"32",X"1E",X"98",
		X"21",X"90",X"00",X"C3",X"8D",X"1B",X"3E",X"01",X"32",X"6E",X"70",X"3E",X"32",X"32",X"46",X"70",
		X"32",X"02",X"98",X"3E",X"3C",X"32",X"44",X"70",X"32",X"03",X"98",X"21",X"90",X"00",X"C3",X"8D",
		X"1B",X"3E",X"02",X"32",X"6E",X"70",X"3E",X"36",X"32",X"46",X"70",X"32",X"02",X"98",X"3E",X"3E",
		X"32",X"44",X"70",X"32",X"03",X"98",X"21",X"18",X"00",X"C3",X"8D",X"1B",X"3E",X"03",X"32",X"6E",
		X"70",X"3E",X"1C",X"32",X"47",X"70",X"3E",X"04",X"32",X"4B",X"70",X"3E",X"04",X"32",X"50",X"70",
		X"32",X"4F",X"70",X"3E",X"34",X"32",X"46",X"70",X"3E",X"42",X"32",X"44",X"70",X"3E",X"01",X"32",
		X"48",X"70",X"AF",X"32",X"49",X"70",X"32",X"4A",X"70",X"32",X"8E",X"70",X"32",X"A1",X"70",X"21",
		X"18",X"00",X"32",X"6C",X"70",X"3E",X"02",X"32",X"64",X"70",X"32",X"80",X"70",X"22",X"9E",X"70",
		X"21",X"A0",X"70",X"34",X"C9",X"ED",X"4B",X"9E",X"70",X"0B",X"ED",X"43",X"9E",X"70",X"78",X"B1",
		X"C0",X"3A",X"A0",X"70",X"FE",X"01",X"CA",X"C5",X"1B",X"FE",X"02",X"CA",X"EC",X"1B",X"FE",X"03",
		X"CA",X"F7",X"1B",X"FE",X"04",X"CA",X"07",X"1C",X"FE",X"05",X"CA",X"22",X"1C",X"FE",X"06",X"CA",
		X"3D",X"1C",X"C3",X"B1",X"1A",X"3A",X"33",X"70",X"B7",X"28",X"12",X"3A",X"AE",X"70",X"B7",X"28",
		X"07",X"3E",X"01",X"32",X"1B",X"70",X"18",X"05",X"3E",X"02",X"32",X"1B",X"70",X"3E",X"02",X"32",
		X"6E",X"70",X"21",X"18",X"00",X"AF",X"32",X"6C",X"70",X"C3",X"8D",X"1B",X"3E",X"03",X"32",X"6E",
		X"70",X"21",X"90",X"00",X"C3",X"8D",X"1B",X"AF",X"32",X"6E",X"70",X"32",X"1F",X"98",X"32",X"1E",
		X"98",X"21",X"90",X"00",X"C3",X"8D",X"1B",X"3E",X"01",X"32",X"89",X"70",X"3E",X"32",X"32",X"46",
		X"70",X"32",X"02",X"98",X"3E",X"BD",X"32",X"44",X"70",X"32",X"03",X"98",X"21",X"90",X"00",X"C3",
		X"8D",X"1B",X"3E",X"02",X"32",X"89",X"70",X"3E",X"36",X"32",X"46",X"70",X"32",X"02",X"98",X"3E",
		X"BB",X"32",X"44",X"70",X"32",X"03",X"98",X"21",X"18",X"00",X"C3",X"8D",X"1B",X"3E",X"03",X"32",
		X"89",X"70",X"3E",X"1C",X"32",X"47",X"70",X"3E",X"04",X"32",X"4B",X"70",X"3E",X"04",X"32",X"50",
		X"70",X"32",X"4F",X"70",X"3E",X"34",X"32",X"46",X"70",X"3E",X"B8",X"32",X"44",X"70",X"3E",X"02",
		X"32",X"48",X"70",X"AF",X"32",X"49",X"70",X"32",X"4A",X"70",X"32",X"8E",X"70",X"32",X"A1",X"70",
		X"21",X"18",X"00",X"32",X"6C",X"70",X"3E",X"02",X"32",X"64",X"70",X"32",X"80",X"70",X"C3",X"8D",
		X"1B",X"3E",X"02",X"32",X"A1",X"70",X"3E",X"01",X"32",X"A0",X"70",X"AF",X"32",X"AB",X"70",X"32",
		X"AC",X"70",X"32",X"50",X"70",X"32",X"4F",X"70",X"32",X"13",X"70",X"32",X"12",X"70",X"32",X"4B",
		X"70",X"32",X"AA",X"70",X"32",X"B4",X"70",X"32",X"6E",X"70",X"32",X"89",X"70",X"32",X"AB",X"70",
		X"32",X"AC",X"70",X"32",X"61",X"70",X"32",X"7D",X"70",X"32",X"B0",X"70",X"32",X"B1",X"70",X"32",
		X"B2",X"70",X"32",X"B3",X"70",X"3E",X"10",X"32",X"00",X"98",X"3E",X"04",X"32",X"01",X"98",X"21",
		X"00",X"02",X"22",X"A2",X"70",X"01",X"00",X"04",X"ED",X"43",X"A4",X"70",X"01",X"00",X"02",X"ED",
		X"43",X"A6",X"70",X"3E",X"09",X"32",X"AD",X"70",X"C3",X"F6",X"16",X"C9",X"06",X"07",X"0E",X"38",
		X"CF",X"3A",X"B8",X"70",X"B7",X"28",X"07",X"AF",X"32",X"B6",X"70",X"32",X"BB",X"70",X"3A",X"BA",
		X"70",X"FE",X"09",X"30",X"3C",X"FE",X"00",X"28",X"05",X"FE",X"09",X"DC",X"42",X"1D",X"3A",X"B7",
		X"70",X"B7",X"3A",X"B6",X"70",X"28",X"05",X"CD",X"7B",X"1D",X"18",X"03",X"CD",X"6D",X"1D",X"3A",
		X"B9",X"70",X"B7",X"3A",X"B8",X"70",X"CA",X"75",X"1F",X"B7",X"28",X"15",X"DD",X"21",X"BE",X"70",
		X"CD",X"BB",X"1D",X"DD",X"21",X"C9",X"70",X"CD",X"BB",X"1D",X"DD",X"21",X"D4",X"70",X"CD",X"BB",
		X"1D",X"C9",X"4F",X"FE",X"07",X"38",X"14",X"3A",X"BB",X"70",X"B7",X"C0",X"79",X"D6",X"06",X"32",
		X"B6",X"70",X"AF",X"32",X"B7",X"70",X"3C",X"32",X"BB",X"70",X"C9",X"3A",X"BC",X"70",X"B7",X"C0",
		X"79",X"32",X"B8",X"70",X"AF",X"32",X"B9",X"70",X"3C",X"32",X"BC",X"70",X"C9",X"21",X"C9",X"1F",
		X"EF",X"79",X"B7",X"20",X"0F",X"21",X"B7",X"70",X"36",X"01",X"C9",X"B7",X"C8",X"21",X"CF",X"1F",
		X"EF",X"79",X"B7",X"C8",X"21",X"B6",X"70",X"AF",X"77",X"23",X"77",X"32",X"BA",X"70",X"32",X"BB",
		X"70",X"C9",X"0E",X"00",X"06",X"08",X"CF",X"06",X"09",X"CF",X"06",X"0A",X"C3",X"08",X"00",X"06",
		X"00",X"4D",X"CF",X"06",X"01",X"4C",X"CF",X"29",X"06",X"02",X"4D",X"CF",X"06",X"03",X"4C",X"CF",
		X"29",X"06",X"04",X"4D",X"CF",X"06",X"05",X"4C",X"C3",X"08",X"00",X"DD",X"35",X"01",X"C0",X"3A",
		X"BD",X"70",X"DD",X"77",X"01",X"DD",X"35",X"00",X"28",X"18",X"DD",X"CB",X"00",X"46",X"C8",X"DD",
		X"7E",X"08",X"B7",X"C8",X"DD",X"86",X"07",X"C8",X"DD",X"77",X"07",X"DD",X"46",X"0A",X"4F",X"C3",
		X"08",X"00",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"7E",X"57",X"E6",X"E0",X"23",X"28",X"48",X"DD",
		X"75",X"02",X"DD",X"74",X"03",X"07",X"07",X"07",X"21",X"2F",X"1E",X"06",X"00",X"4F",X"09",X"7E",
		X"DD",X"77",X"00",X"7A",X"E6",X"1F",X"C8",X"3D",X"07",X"4F",X"DD",X"6E",X"04",X"DD",X"66",X"05",
		X"09",X"7E",X"23",X"66",X"6F",X"DD",X"4E",X"09",X"ED",X"42",X"DD",X"4E",X"06",X"DD",X"71",X"07",
		X"DD",X"46",X"0A",X"CF",X"78",X"D6",X"08",X"87",X"47",X"4D",X"CF",X"04",X"4C",X"C3",X"08",X"00",
		X"00",X"01",X"02",X"04",X"08",X"10",X"20",X"7A",X"5D",X"54",X"23",X"DD",X"75",X"02",X"DD",X"74",
		X"03",X"21",X"49",X"1E",X"E6",X"0E",X"C3",X"29",X"00",X"57",X"1E",X"69",X"1E",X"73",X"1E",X"7A",
		X"1E",X"81",X"1E",X"88",X"1E",X"94",X"1E",X"1A",X"87",X"4F",X"06",X"00",X"21",X"B5",X"1E",X"09",
		X"DD",X"75",X"04",X"DD",X"74",X"05",X"C3",X"E2",X"1D",X"1A",X"32",X"BD",X"70",X"DD",X"77",X"01",
		X"C3",X"E2",X"1D",X"1A",X"DD",X"77",X"06",X"C3",X"E2",X"1D",X"1A",X"DD",X"77",X"08",X"C3",X"E2",
		X"1D",X"1A",X"DD",X"77",X"09",X"C3",X"E2",X"1D",X"1A",X"DD",X"77",X"02",X"13",X"1A",X"DD",X"77",
		X"03",X"C3",X"E2",X"1D",X"1B",X"DD",X"73",X"02",X"DD",X"72",X"03",X"DD",X"36",X"00",X"01",X"DD",
		X"36",X"01",X"01",X"E1",X"CD",X"92",X"1D",X"21",X"00",X"01",X"22",X"B8",X"70",X"AF",X"32",X"BA",
		X"70",X"32",X"BC",X"70",X"C9",X"5D",X"0D",X"9C",X"0C",X"E7",X"0B",X"3C",X"0B",X"9B",X"0A",X"02",
		X"0A",X"73",X"09",X"EB",X"08",X"6B",X"08",X"F2",X"07",X"80",X"07",X"14",X"07",X"AE",X"06",X"4E",
		X"06",X"F4",X"05",X"9E",X"05",X"4D",X"05",X"01",X"05",X"B9",X"04",X"75",X"04",X"35",X"04",X"F9",
		X"03",X"C0",X"03",X"8A",X"03",X"57",X"03",X"27",X"03",X"FA",X"02",X"CF",X"02",X"A7",X"02",X"81",
		X"02",X"5D",X"02",X"3B",X"02",X"1B",X"02",X"FC",X"01",X"E0",X"01",X"C5",X"01",X"AC",X"01",X"94",
		X"01",X"7D",X"01",X"68",X"01",X"53",X"01",X"40",X"01",X"2E",X"01",X"1D",X"01",X"0D",X"01",X"FE",
		X"00",X"F0",X"00",X"E2",X"00",X"D6",X"00",X"CA",X"00",X"BE",X"00",X"B4",X"00",X"AA",X"00",X"A0",
		X"00",X"97",X"00",X"8F",X"00",X"87",X"00",X"7F",X"00",X"78",X"00",X"71",X"00",X"6B",X"00",X"65",
		X"00",X"5F",X"00",X"5A",X"00",X"55",X"00",X"50",X"00",X"4C",X"00",X"47",X"00",X"43",X"00",X"40",
		X"00",X"3C",X"00",X"39",X"00",X"35",X"00",X"32",X"00",X"30",X"00",X"2D",X"00",X"2A",X"00",X"28",
		X"00",X"26",X"00",X"24",X"00",X"22",X"00",X"20",X"00",X"1E",X"00",X"1C",X"00",X"1B",X"00",X"19",
		X"00",X"18",X"00",X"16",X"00",X"15",X"00",X"14",X"00",X"13",X"00",X"12",X"00",X"11",X"00",X"10",
		X"00",X"0F",X"00",X"0E",X"00",X"21",X"A8",X"1F",X"11",X"BE",X"70",X"01",X"21",X"00",X"ED",X"B0",
		X"87",X"4F",X"87",X"81",X"4F",X"06",X"00",X"21",X"D5",X"1F",X"09",X"11",X"C0",X"70",X"ED",X"A0",
		X"ED",X"A0",X"11",X"CB",X"70",X"ED",X"A0",X"ED",X"A0",X"11",X"D6",X"70",X"ED",X"A0",X"ED",X"A0",
		X"3E",X"01",X"32",X"B9",X"70",X"C3",X"2C",X"1D",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"08",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"09",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"0A",X"92",X"1D",X"FF",X"1F",X"38",X"20",X"7A",
		X"1D",X"1B",X"20",X"4A",X"20",X"DA",X"20",X"DA",X"20",X"DA",X"20",X"DB",X"20",X"FF",X"20",X"1E",
		X"21",X"31",X"21",X"46",X"21",X"58",X"21",X"67",X"21",X"72",X"21",X"77",X"21",X"80",X"21",X"88",
		X"21",X"8D",X"21",X"92",X"21",X"9A",X"21",X"9F",X"21",X"A4",X"21",X"AC",X"21",X"B1",X"21",X"AF",
		X"21",X"E1",X"70",X"36",X"0A",X"2D",X"36",X"00",X"2C",X"35",X"28",X"0D",X"4E",X"CD",X"94",X"1D",
		X"21",X"00",X"00",X"22",X"E2",X"70",X"C3",X"9F",X"1D",X"4F",X"C9",X"21",X"E0",X"70",X"34",X"7E",
		X"FE",X"0C",X"28",X"E2",X"5F",X"E6",X"01",X"20",X"0C",X"16",X"00",X"2A",X"E2",X"70",X"19",X"22",
		X"E2",X"70",X"CD",X"9F",X"1D",X"AF",X"4F",X"C9",X"3E",X"02",X"32",X"E4",X"70",X"21",X"7F",X"00",
		X"CD",X"9F",X"1D",X"0E",X"0B",X"CD",X"94",X"1D",X"18",X"EB",X"3A",X"E4",X"70",X"3D",X"32",X"E4",
		X"70",X"28",X"0F",X"FE",X"FF",X"28",X"28",X"FE",X"02",X"38",X"02",X"18",X"D8",X"CD",X"92",X"1D",
		X"18",X"D3",X"3E",X"0C",X"32",X"E5",X"70",X"3E",X"0A",X"32",X"E6",X"70",X"4F",X"CD",X"94",X"1D",
		X"21",X"7F",X"00",X"22",X"E7",X"70",X"CD",X"9F",X"1D",X"AF",X"32",X"E4",X"70",X"4F",X"C9",X"3A",
		X"E5",X"70",X"3D",X"32",X"E5",X"70",X"FE",X"07",X"38",X"0F",X"2A",X"E7",X"70",X"2B",X"2B",X"2B",
		X"2B",X"22",X"E7",X"70",X"CD",X"9F",X"1D",X"18",X"E0",X"FE",X"06",X"28",X"12",X"B7",X"28",X"1D",
		X"2A",X"E7",X"70",X"23",X"23",X"23",X"23",X"22",X"E7",X"70",X"CD",X"9F",X"1D",X"18",X"CA",X"3A",
		X"E6",X"70",X"3D",X"32",X"E6",X"70",X"4F",X"CD",X"94",X"1D",X"79",X"18",X"E0",X"3A",X"E6",X"70",
		X"3D",X"32",X"E6",X"70",X"4F",X"28",X"10",X"CD",X"94",X"1D",X"21",X"00",X"00",X"CD",X"9F",X"1D",
		X"3E",X"0C",X"32",X"E5",X"70",X"18",X"A8",X"0E",X"FF",X"C9",X"0D",X"01",X"24",X"03",X"04",X"05",
		X"09",X"07",X"00",X"71",X"07",X"FF",X"51",X"51",X"71",X"6F",X"8D",X"8A",X"07",X"00",X"6F",X"07",
		X"FF",X"4F",X"4F",X"6F",X"6D",X"8C",X"88",X"6A",X"6C",X"6D",X"6F",X"91",X"8F",X"8D",X"0D",X"01",
		X"24",X"05",X"08",X"07",X"00",X"69",X"07",X"FF",X"49",X"49",X"69",X"69",X"8A",X"80",X"07",X"00",
		X"67",X"07",X"FF",X"49",X"47",X"67",X"67",X"88",X"80",X"80",X"80",X"80",X"86",X"85",X"01",X"18",
		X"05",X"08",X"85",X"89",X"8A",X"80",X"83",X"87",X"88",X"80",X"66",X"68",X"6A",X"6C",X"8D",X"88",
		X"81",X"01",X"24",X"03",X"04",X"05",X"09",X"71",X"72",X"73",X"74",X"79",X"76",X"79",X"78",X"7B",
		X"99",X"A0",X"74",X"99",X"C0",X"0D",X"01",X"24",X"05",X"08",X"6D",X"6F",X"70",X"71",X"60",X"72",
		X"60",X"74",X"60",X"91",X"A0",X"60",X"91",X"C0",X"01",X"24",X"05",X"08",X"61",X"63",X"64",X"85",
		X"86",X"88",X"81",X"A0",X"68",X"81",X"C0",X"01",X"30",X"03",X"04",X"05",X"0A",X"8D",X"8D",X"8D",
		X"8D",X"0D",X"05",X"00",X"0B",X"7C",X"21",X"05",X"00",X"0B",X"7C",X"21",X"60",X"0B",X"7C",X"21",
		X"01",X"0C",X"03",X"04",X"05",X"0A",X"ED",X"0D",X"01",X"0C",X"05",X"0A",X"F1",X"01",X"0C",X"05",
		X"0A",X"F4",X"01",X"24",X"03",X"01",X"05",X"0F",X"47",X"0D",X"05",X"00",X"0B",X"7C",X"21",X"05",
		X"00",X"0B",X"7C",X"21",X"01",X"24",X"03",X"02",X"05",X"0F",X"41",X"0D",X"05",X"00",X"0B",X"7C",
		X"21",X"05",X"00",X"0B",X"7C",X"21",X"3A",X"F2",X"70",X"B7",X"C8",X"AF",X"32",X"6E",X"70",X"32",
		X"89",X"70",X"3A",X"03",X"98",X"DD",X"21",X"EE",X"70",X"DD",X"BE",X"00",X"28",X"09",X"DD",X"72",
		X"FF",X"DD",X"36",X"FE",X"01",X"18",X"05",X"3E",X"01",X"32",X"F3",X"70",X"21",X"F1",X"70",X"34",
		X"3E",X"06",X"BE",X"C0",X"36",X"00",X"3A",X"F0",X"70",X"EE",X"01",X"32",X"F0",X"70",X"B7",X"20",
		X"3A",X"3A",X"F3",X"70",X"B7",X"20",X"05",X"DD",X"35",X"00",X"18",X"5C",X"DD",X"34",X"00",X"DD",
		X"7E",X"00",X"32",X"03",X"98",X"DD",X"35",X"FF",X"DD",X"7E",X"FF",X"32",X"02",X"98",X"FE",X"00",
		X"28",X"07",X"DD",X"7E",X"00",X"FE",X"0F",X"30",X"3F",X"AF",X"32",X"F2",X"70",X"32",X"F3",X"70",
		X"32",X"ED",X"70",X"32",X"EE",X"70",X"32",X"03",X"98",X"18",X"2D",X"FD",X"21",X"EB",X"70",X"21",
		X"64",X"22",X"3A",X"EF",X"70",X"3C",X"FE",X"03",X"20",X"01",X"AF",X"32",X"EF",X"70",X"5F",X"16",
		X"00",X"19",X"56",X"3A",X"F3",X"70",X"B7",X"20",X"0A",X"CB",X"F2",X"FD",X"72",X"00",X"DD",X"35",
		X"00",X"18",X"05",X"FD",X"72",X"00",X"18",X"A4",X"21",X"EB",X"70",X"11",X"1C",X"98",X"01",X"04",
		X"00",X"ED",X"B0",X"C9",X"2D",X"2F",X"2E",X"00",X"3A",X"F4",X"70",X"B7",X"28",X"05",X"3D",X"32",
		X"F4",X"70",X"C9",X"CD",X"14",X"23",X"FE",X"FF",X"28",X"34",X"F5",X"FE",X"05",X"20",X"07",X"3E",
		X"01",X"32",X"26",X"70",X"18",X"04",X"FE",X"06",X"28",X"F5",X"F1",X"CB",X"27",X"21",X"BE",X"23",
		X"16",X"00",X"5F",X"19",X"7E",X"32",X"66",X"70",X"23",X"7E",X"32",X"6D",X"70",X"3E",X"30",X"32",
		X"F4",X"70",X"3A",X"98",X"70",X"32",X"69",X"70",X"3E",X"01",X"32",X"67",X"70",X"C9",X"3A",X"46",
		X"70",X"FE",X"80",X"30",X"11",X"3A",X"97",X"70",X"B7",X"20",X"08",X"3A",X"44",X"70",X"FE",X"80",
		X"D2",X"C6",X"22",X"C3",X"E2",X"22",X"3A",X"5B",X"70",X"FE",X"40",X"38",X"05",X"FE",X"42",X"D8",
		X"18",X"0C",X"3E",X"00",X"32",X"62",X"70",X"3E",X"01",X"32",X"63",X"70",X"18",X"10",X"3E",X"01",
		X"18",X"F2",X"3A",X"44",X"70",X"21",X"5B",X"70",X"BE",X"C8",X"38",X"F2",X"18",X"E4",X"3A",X"44",
		X"70",X"FE",X"40",X"38",X"0E",X"FE",X"60",X"38",X"05",X"3A",X"99",X"70",X"18",X"08",X"3A",X"9A",
		X"70",X"18",X"03",X"3A",X"9B",X"70",X"32",X"64",X"70",X"3E",X"02",X"32",X"66",X"70",X"3E",X"01",
		X"32",X"67",X"70",X"C9",X"21",X"44",X"70",X"3A",X"5B",X"70",X"D6",X"19",X"BE",X"D2",X"4B",X"23",
		X"C6",X"32",X"BE",X"DA",X"4B",X"23",X"21",X"46",X"70",X"3A",X"5A",X"70",X"C6",X"19",X"BE",X"DA",
		X"4B",X"23",X"D6",X"32",X"BE",X"D2",X"4B",X"23",X"AF",X"06",X"0C",X"C5",X"F5",X"CD",X"4E",X"23",
		X"B7",X"28",X"03",X"F1",X"C1",X"C9",X"F1",X"C1",X"3C",X"10",X"F0",X"3E",X"FF",X"C9",X"CB",X"27",
		X"CB",X"27",X"DD",X"21",X"8E",X"23",X"16",X"00",X"5F",X"DD",X"19",X"3A",X"5A",X"70",X"D6",X"19",
		X"DD",X"86",X"00",X"08",X"3A",X"5B",X"70",X"D6",X"19",X"DD",X"86",X"01",X"21",X"44",X"70",X"BE",
		X"D2",X"8C",X"23",X"DD",X"86",X"02",X"BE",X"DA",X"8C",X"23",X"21",X"46",X"70",X"08",X"BE",X"DA",
		X"8C",X"23",X"DD",X"96",X"03",X"BE",X"D2",X"8C",X"23",X"3E",X"01",X"C9",X"AF",X"C9",X"0F",X"0D",
		X"0F",X"0F",X"11",X"01",X"12",X"11",X"1B",X"00",X"14",X"10",X"25",X"00",X"14",X"11",X"2F",X"00",
		X"14",X"11",X"31",X"08",X"15",X"11",X"31",X"14",X"12",X"11",X"31",X"1E",X"13",X"13",X"25",X"1F",
		X"14",X"14",X"19",X"1E",X"15",X"13",X"11",X"1C",X"15",X"12",X"11",X"14",X"0F",X"12",X"02",X"00",
		X"03",X"00",X"04",X"00",X"05",X"00",X"06",X"00",X"07",X"00",X"08",X"00",X"06",X"01",X"06",X"01",
		X"08",X"01",X"09",X"01",X"0A",X"01",X"21",X"40",X"88",X"ED",X"4B",X"F5",X"70",X"09",X"22",X"F5",
		X"70",X"3A",X"F7",X"70",X"87",X"21",X"16",X"24",X"16",X"00",X"5F",X"19",X"E5",X"DD",X"E1",X"DD",
		X"6E",X"00",X"DD",X"66",X"01",X"3A",X"02",X"70",X"CB",X"6F",X"28",X"04",X"11",X"E9",X"00",X"19",
		X"E5",X"C1",X"2A",X"F5",X"70",X"0A",X"FE",X"2F",X"C8",X"D6",X"30",X"77",X"CB",X"E4",X"36",X"05",
		X"CB",X"A4",X"23",X"03",X"18",X"EF",X"5B",X"24",X"64",X"24",X"74",X"24",X"84",X"24",X"9E",X"24",
		X"B6",X"24",X"C0",X"24",X"C8",X"24",X"20",X"20",X"20",X"20",X"20",X"55",X"4E",X"20",X"42",X"4F",
		X"4E",X"4A",X"4F",X"55",X"52",X"20",X"41",X"20",X"4A",X"41",X"43",X"51",X"55",X"45",X"53",X"20",
		X"44",X"45",X"20",X"50",X"45",X"50",X"45",X"20",X"50",X"45",X"54",X"49",X"54",X"20",X"45",X"54",
		X"20",X"48",X"45",X"4E",X"4B",X"20",X"20",X"20",X"20",X"20",X"20",X"50",X"52",X"45",X"53",X"45",
		X"4E",X"54",X"41",X"2F",X"49",X"4E",X"53",X"45",X"52",X"54",X"45",X"40",X"4D",X"4F",X"4E",X"45",
		X"44",X"41",X"53",X"2F",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"40",X"40",X"40",X"2F",X"50",X"55",X"4C",X"53",X"45",X"40",X"55",X"4E",X"4F",X"40",X"4F",X"40",
		X"44",X"4F",X"53",X"40",X"4A",X"55",X"47",X"41",X"44",X"4F",X"52",X"45",X"53",X"2F",X"40",X"40",
		X"40",X"40",X"50",X"55",X"4C",X"53",X"45",X"40",X"55",X"4E",X"40",X"4A",X"55",X"47",X"41",X"44",
		X"4F",X"52",X"40",X"40",X"40",X"2F",X"47",X"41",X"4D",X"45",X"40",X"4F",X"56",X"45",X"52",X"2F",
		X"43",X"52",X"45",X"44",X"49",X"54",X"53",X"2F",X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",
		X"54",X"40",X"31",X"39",X"38",X"34",X"40",X"42",X"59",X"40",X"49",X"54",X"49",X"53",X"41",X"2F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"50",X"52",X"45",X"53",X"45",X"4E",X"54",X"53",X"2F",X"40",X"40",X"49",
		X"4E",X"53",X"45",X"52",X"54",X"40",X"43",X"4F",X"49",X"4E",X"40",X"40",X"2F",X"40",X"40",X"40",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"2F",X"50",X"55",X"53",
		X"48",X"40",X"4F",X"4E",X"45",X"40",X"4F",X"52",X"40",X"54",X"57",X"4F",X"40",X"50",X"4C",X"41",
		X"59",X"45",X"52",X"53",X"40",X"40",X"2F",X"40",X"40",X"50",X"55",X"53",X"48",X"40",X"4F",X"4E",
		X"4C",X"59",X"40",X"4F",X"4E",X"45",X"40",X"50",X"4C",X"41",X"59",X"45",X"52",X"40",X"2F",X"47",
		X"41",X"4D",X"45",X"40",X"4F",X"56",X"45",X"52",X"2F",X"43",X"52",X"45",X"44",X"49",X"54",X"53",
		X"2F",X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"40",X"31",X"39",X"38",X"34",X"40",
		X"42",X"59",X"40",X"49",X"54",X"49",X"53",X"41",X"2F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3A",X"FB",X"70",
		X"87",X"21",X"B8",X"26",X"16",X"00",X"5F",X"19",X"5E",X"23",X"56",X"ED",X"53",X"FD",X"70",X"DD",
		X"2A",X"FD",X"70",X"DD",X"5E",X"03",X"DD",X"56",X"04",X"2A",X"FD",X"70",X"46",X"23",X"4E",X"23",
		X"7E",X"23",X"B7",X"28",X"31",X"23",X"23",X"08",X"78",X"08",X"D9",X"21",X"40",X"88",X"ED",X"4B",
		X"F9",X"70",X"09",X"E5",X"D9",X"7E",X"23",X"D9",X"77",X"D9",X"1A",X"13",X"D9",X"CB",X"E4",X"77",
		X"CB",X"A4",X"23",X"D9",X"10",X"EF",X"D9",X"E1",X"01",X"20",X"00",X"09",X"D9",X"08",X"47",X"08",
		X"0D",X"D9",X"20",X"DF",X"D9",X"C9",X"00",X"54",X"5D",X"23",X"08",X"78",X"08",X"D9",X"21",X"40",
		X"88",X"ED",X"4B",X"F9",X"70",X"09",X"E5",X"D9",X"7E",X"23",X"D9",X"77",X"D9",X"1A",X"D9",X"CB",
		X"E4",X"77",X"CB",X"A4",X"23",X"D9",X"10",X"F0",X"D9",X"E1",X"01",X"20",X"00",X"09",X"D9",X"08",
		X"47",X"08",X"0D",X"D9",X"20",X"E0",X"D9",X"C9",X"C8",X"26",X"35",X"27",X"87",X"27",X"8C",X"2E",
		X"91",X"2E",X"9A",X"2E",X"A3",X"2E",X"AC",X"2E",X"15",X"05",X"00",X"15",X"9B",X"9C",X"9D",X"AA",
		X"AB",X"AC",X"AD",X"BA",X"00",X"C0",X"AA",X"AB",X"AC",X"AD",X"9B",X"9C",X"9D",X"CC",X"CD",X"CE",
		X"CF",X"9E",X"9F",X"A0",X"AE",X"AF",X"B0",X"B1",X"BB",X"00",X"C1",X"AE",X"AF",X"B0",X"B1",X"9E",
		X"9F",X"A0",X"AE",X"B3",X"B4",X"B1",X"A1",X"A2",X"A3",X"AE",X"B3",X"B4",X"B1",X"BB",X"00",X"C1",
		X"AE",X"C4",X"C8",X"B1",X"A1",X"A2",X"A3",X"AE",X"C4",X"C8",X"B1",X"A4",X"A5",X"A6",X"AE",X"B2",
		X"B5",X"B1",X"BC",X"BE",X"C2",X"AE",X"C6",X"C9",X"B1",X"A4",X"A5",X"A6",X"AE",X"C6",X"C9",X"B1",
		X"A7",X"A8",X"A9",X"B6",X"B7",X"B8",X"B9",X"BD",X"BF",X"C3",X"C5",X"C7",X"CA",X"CB",X"A7",X"A8",
		X"A9",X"C5",X"C7",X"CA",X"CB",X"0D",X"06",X"00",X"1E",X"01",X"02",X"03",X"04",X"05",X"06",X"07",
		X"08",X"09",X"0A",X"0B",X"0C",X"0D",X"0E",X"0F",X"10",X"11",X"12",X"13",X"14",X"15",X"16",X"17",
		X"18",X"19",X"1A",X"1B",X"1C",X"1D",X"1E",X"1F",X"20",X"21",X"22",X"23",X"24",X"25",X"26",X"27",
		X"28",X"29",X"2A",X"2B",X"2C",X"2D",X"2E",X"2F",X"30",X"31",X"32",X"33",X"34",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"35",
		X"36",X"37",X"38",X"39",X"3A",X"3B",X"3C",X"20",X"1C",X"01",X"0C",X"2B",X"3F",X"3F",X"40",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"5B",X"C5",X"3F",X"3F",X"3F",X"40",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"5B",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"40",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"5B",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"41",X"42",X"42",X"42",X"42",X"42",X"46",X"42",X"42",X"42",X"42",X"5F",X"42",X"42",X"42",
		X"42",X"55",X"42",X"42",X"42",X"42",X"42",X"59",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"43",X"8A",X"8A",X"8A",X"8A",X"8A",X"47",X"8A",X"49",X"4F",X"57",X"53",X"57",X"52",X"51",
		X"8A",X"56",X"8A",X"8A",X"8A",X"8A",X"8A",X"5A",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"43",X"8A",X"8A",X"8A",X"8A",X"8A",X"47",X"8A",X"4A",X"00",X"00",X"4D",X"00",X"00",X"54",
		X"8A",X"56",X"8A",X"8A",X"8A",X"8A",X"8A",X"5A",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"44",X"45",X"45",X"45",X"45",X"45",X"47",X"8A",X"4B",X"4C",X"4C",X"4E",X"4C",X"4C",X"50",
		X"8A",X"56",X"45",X"45",X"45",X"45",X"45",X"5C",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"43",X"8A",X"8A",X"8A",X"8A",X"8A",X"48",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",
		X"45",X"58",X"8A",X"8A",X"8A",X"8A",X"8A",X"5A",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"43",X"8A",X"8A",X"8A",X"8A",X"8A",X"47",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",
		X"8A",X"56",X"8A",X"8A",X"8A",X"8A",X"8A",X"5A",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"43",X"8A",X"8A",X"8A",X"8A",X"8A",X"47",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",
		X"8A",X"56",X"8A",X"8A",X"8A",X"8A",X"8A",X"5A",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"43",X"8A",X"8A",X"8A",X"8A",X"8A",X"47",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",
		X"8A",X"56",X"8A",X"8A",X"8A",X"8A",X"8A",X"5A",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"43",X"8A",X"8D",X"8E",X"8F",X"8A",X"47",X"8A",X"8A",X"8A",X"93",X"94",X"95",X"96",X"8A",
		X"8A",X"56",X"8A",X"8D",X"8E",X"8F",X"8A",X"5A",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"43",X"8A",X"90",X"91",X"92",X"8A",X"47",X"8A",X"8A",X"8A",X"97",X"98",X"99",X"9A",X"8A",
		X"8A",X"56",X"8A",X"90",X"91",X"92",X"8A",X"5A",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"43",X"8A",X"8A",X"8A",X"8A",X"8A",X"47",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",
		X"8A",X"56",X"8A",X"8A",X"8A",X"8A",X"8A",X"5A",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"43",X"8A",X"8A",X"8A",X"8A",X"8A",X"47",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",
		X"8A",X"56",X"8A",X"8A",X"8A",X"8A",X"8A",X"5A",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"43",X"8A",X"8A",X"8A",X"8A",X"8A",X"60",X"61",X"61",X"61",X"61",X"61",X"61",X"61",X"61",
		X"61",X"62",X"8A",X"8A",X"8A",X"8A",X"8A",X"5A",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"5D",X"5E",X"5E",X"5E",X"5E",X"5E",X"47",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",
		X"8A",X"56",X"5E",X"5E",X"5E",X"5E",X"5E",X"63",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"43",X"8A",X"8A",X"8A",X"8A",X"8A",X"47",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",
		X"8A",X"56",X"8A",X"8A",X"8A",X"8A",X"8A",X"5A",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"43",X"8A",X"8A",X"8A",X"8A",X"8A",X"47",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",
		X"8A",X"56",X"8A",X"8A",X"8A",X"8A",X"8A",X"5A",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"43",X"66",X"66",X"66",X"66",X"66",X"74",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"66",X"79",X"66",X"66",X"66",X"66",X"66",X"5A",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"43",X"66",X"66",X"66",X"66",X"66",X"74",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"66",X"79",X"66",X"66",X"66",X"66",X"66",X"5A",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"64",X"73",X"73",X"73",X"73",X"73",X"72",X"73",X"73",X"73",X"73",X"73",X"73",X"73",X"73",
		X"73",X"78",X"73",X"73",X"73",X"73",X"73",X"80",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"65",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"85",X"66",X"66",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"7F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"65",
		X"66",X"68",X"69",X"69",X"69",X"69",X"69",X"69",X"69",X"69",X"69",X"69",X"81",X"69",X"69",X"69",
		X"69",X"69",X"69",X"69",X"69",X"69",X"69",X"7A",X"66",X"7F",X"3F",X"3F",X"3F",X"3F",X"65",X"66",
		X"6B",X"6A",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"82",X"66",X"66",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"7B",X"7C",X"66",X"7F",X"3F",X"3F",X"65",X"66",X"6B",
		X"6A",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"82",X"66",X"66",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"7B",X"7C",X"66",X"7F",X"65",X"66",X"6B",X"6A",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"84",X"66",X"66",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"7B",X"7C",X"66",X"66",X"6C",X"6D",X"6E",
		X"6E",X"6E",X"6E",X"6E",X"6E",X"6E",X"6E",X"6E",X"6E",X"6E",X"6E",X"71",X"83",X"77",X"6E",X"6E",
		X"6E",X"6E",X"6E",X"6E",X"6E",X"6E",X"6E",X"6E",X"6E",X"6E",X"7D",X"7E",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"00",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",
		X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",
		X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",
		X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",
		X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",
		X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",
		X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",
		X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",
		X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"13",X"13",X"1B",X"1B",X"1B",X"13",X"13",X"13",X"13",X"13",X"1B",X"1B",X"1B",X"1B",X"13",
		X"13",X"13",X"13",X"1B",X"1B",X"1B",X"13",X"13",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"13",X"13",X"1B",X"1B",X"1B",X"13",X"13",X"13",X"13",X"13",X"1F",X"1F",X"1F",X"1F",X"13",
		X"13",X"13",X"13",X"1B",X"1B",X"1B",X"13",X"13",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",
		X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",
		X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",
		X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",
		X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",
		X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",
		X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"13",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",
		X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"13",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"13",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",
		X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"13",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",
		X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1A",X"1F",X"1F",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1A",X"1F",X"1F",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1A",X"1F",X"1F",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1A",X"1F",X"1F",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"01",X"01",X"00",X"00",
		X"00",X"05",X"01",X"00",X"1C",X"D0",X"D1",X"D2",X"D3",X"D4",X"05",X"01",X"00",X"1C",X"D0",X"D1",
		X"D2",X"D3",X"D5",X"05",X"01",X"00",X"1C",X"D6",X"D7",X"D8",X"D9",X"DA",X"05",X"01",X"00",X"1C",
		X"66",X"66",X"66",X"66",X"66",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
