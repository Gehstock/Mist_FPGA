library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_OBJ_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_OBJ_1 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",X"00",X"02",X"02",X"FE",X"FE",X"42",X"02",X"00",X"00",
		X"62",X"F2",X"BA",X"9A",X"9E",X"CE",X"46",X"00",X"8C",X"DE",X"F2",X"B2",X"92",X"86",X"04",X"00",
		X"08",X"FE",X"FE",X"C8",X"68",X"38",X"18",X"00",X"1C",X"BE",X"A2",X"A2",X"A2",X"E6",X"E4",X"00",
		X"0C",X"9E",X"92",X"92",X"D2",X"7E",X"3C",X"00",X"C0",X"E0",X"B0",X"9E",X"8E",X"C0",X"C0",X"00",
		X"0C",X"6E",X"9A",X"9A",X"B2",X"F2",X"6C",X"00",X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",X"00",
		X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",
		X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",X"44",X"C6",X"82",X"82",X"C6",X"7C",X"38",X"00",
		X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",X"82",X"92",X"92",X"92",X"FE",X"FE",X"00",X"00",
		X"80",X"90",X"90",X"90",X"90",X"FE",X"FE",X"00",X"9E",X"9E",X"92",X"82",X"C6",X"7C",X"38",X"00",
		X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",X"82",X"82",X"FE",X"FE",X"82",X"82",X"00",X"00",
		X"FC",X"FE",X"02",X"02",X"02",X"06",X"04",X"00",X"82",X"C6",X"6E",X"3C",X"18",X"FE",X"FE",X"00",
		X"02",X"02",X"02",X"02",X"FE",X"FE",X"00",X"00",X"FE",X"FE",X"70",X"38",X"70",X"FE",X"FE",X"00",
		X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",X"00",
		X"70",X"F8",X"88",X"88",X"88",X"FE",X"FE",X"00",X"7A",X"FC",X"8E",X"8A",X"82",X"FE",X"7C",X"00",
		X"72",X"F6",X"9E",X"8C",X"88",X"FE",X"FE",X"00",X"0C",X"5E",X"D2",X"92",X"92",X"F6",X"64",X"00",
		X"80",X"80",X"FE",X"FE",X"80",X"80",X"00",X"00",X"FC",X"FE",X"02",X"02",X"02",X"FE",X"FC",X"00",
		X"F0",X"F8",X"1C",X"0E",X"1C",X"F8",X"F0",X"00",X"F8",X"FE",X"1C",X"38",X"1C",X"FE",X"F8",X"00",
		X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",X"C0",X"F0",X"1E",X"1E",X"F0",X"C0",X"00",X"00",
		X"C2",X"E2",X"F2",X"BA",X"9E",X"8E",X"86",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"00",
		X"00",X"00",X"00",X"01",X"0B",X"0F",X"0F",X"0F",X"00",X"00",X"80",X"C0",X"E8",X"F8",X"F8",X"F8",
		X"07",X"00",X"02",X"03",X"00",X"00",X"00",X"00",X"F0",X"80",X"20",X"60",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"1C",X"1C",X"1C",X"0F",X"03",X"07",X"00",X"F0",X"38",X"38",X"38",X"F0",X"C0",X"E0",
		X"0B",X"08",X"1C",X"1F",X"0F",X"07",X"00",X"00",X"D0",X"10",X"38",X"F8",X"F0",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"05",X"0F",X"07",X"07",X"00",X"00",X"80",X"80",X"D0",X"B8",X"D0",X"E0",
		X"07",X"07",X"07",X"0F",X"05",X"00",X"00",X"00",X"E0",X"E0",X"D0",X"F8",X"D0",X"80",X"80",X"00",
		X"00",X"01",X"00",X"08",X"19",X"0F",X"07",X"07",X"00",X"00",X"80",X"88",X"CC",X"B8",X"D0",X"E0",
		X"07",X"07",X"07",X"0F",X"19",X"09",X"00",X"00",X"E0",X"E0",X"D0",X"F8",X"CC",X"C8",X"80",X"80",
		X"00",X"00",X"00",X"00",X"01",X"0F",X"07",X"07",X"00",X"40",X"80",X"80",X"C0",X"B8",X"D0",X"E0",
		X"07",X"07",X"0F",X"0F",X"01",X"01",X"00",X"00",X"E0",X"E0",X"D8",X"F8",X"C0",X"C0",X"80",X"80",
		X"00",X"08",X"08",X"00",X"20",X"23",X"06",X"04",X"04",X"24",X"44",X"00",X"00",X"9C",X"A5",X"00",
		X"04",X"44",X"42",X"00",X"06",X"E4",X"48",X"00",X"42",X"40",X"06",X"04",X"26",X"22",X"00",X"06",
		X"04",X"06",X"23",X"48",X"08",X"00",X"00",X"00",X"00",X"A5",X"39",X"00",X"08",X"48",X"40",X"00",
		X"00",X"28",X"CC",X"00",X"40",X"46",X"06",X"06",X"00",X"02",X"02",X"00",X"10",X"10",X"00",X"00",
		X"7F",X"6F",X"57",X"EF",X"FD",X"7A",X"3D",X"EF",X"FE",X"FE",X"DE",X"AE",X"DE",X"FF",X"F6",X"6A",
		X"56",X"6F",X"FF",X"FE",X"6D",X"56",X"EF",X"7F",X"B7",X"7E",X"FA",X"F5",X"7B",X"EE",X"D7",X"EF",
		X"00",X"00",X"40",X"62",X"4C",X"00",X"00",X"00",X"00",X"38",X"7C",X"7C",X"7C",X"38",X"00",X"00",
		X"3C",X"42",X"81",X"A5",X"A5",X"99",X"42",X"3C",X"FF",X"81",X"81",X"81",X"81",X"81",X"81",X"FF",
		X"02",X"72",X"73",X"7A",X"73",X"72",X"01",X"00",X"40",X"4E",X"CE",X"5E",X"CE",X"4E",X"80",X"00",
		X"02",X"33",X"33",X"39",X"30",X"30",X"00",X"00",X"40",X"CC",X"CC",X"9C",X"0C",X"0C",X"00",X"00",
		X"1E",X"1E",X"0F",X"1F",X"1F",X"17",X"1F",X"1F",X"F8",X"F8",X"D8",X"F8",X"10",X"F8",X"F8",X"F8",
		X"1B",X"1B",X"0F",X"0F",X"03",X"00",X"00",X"00",X"E8",X"78",X"68",X"E0",X"C0",X"00",X"00",X"00",
		X"1F",X"1D",X"1F",X"0F",X"1F",X"1B",X"1B",X"1F",X"F8",X"F8",X"F8",X"B8",X"B0",X"B8",X"F8",X"F8",
		X"1F",X"1F",X"1D",X"1F",X"1F",X"0F",X"1F",X"17",X"F8",X"E8",X"E8",X"E8",X"F0",X"78",X"F8",X"F8",
		X"00",X"00",X"00",X"00",X"01",X"07",X"07",X"07",X"00",X"00",X"00",X"00",X"80",X"E0",X"30",X"F8",
		X"11",X"1E",X"1F",X"17",X"1F",X"0F",X"1F",X"1F",X"88",X"38",X"B8",X"F0",X"B8",X"B8",X"F8",X"F8",
		X"07",X"08",X"08",X"08",X"07",X"00",X"07",X"08",X"C0",X"20",X"20",X"20",X"C0",X"00",X"C0",X"20",
		X"08",X"08",X"07",X"00",X"00",X"0F",X"04",X"00",X"20",X"20",X"C0",X"00",X"20",X"E0",X"20",X"00",
		X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"C0",X"20",X"20",X"C0",X"00",X"C0",X"20",X"20",
		X"07",X"00",X"06",X"09",X"08",X"08",X"04",X"00",X"C0",X"00",X"20",X"20",X"A0",X"60",X"20",X"00",
		X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"50",X"D0",X"D0",X"D0",X"D0",X"D0",
		X"01",X"01",X"03",X"03",X"00",X"00",X"01",X"01",X"B0",X"B0",X"F0",X"F0",X"FC",X"FE",X"FE",X"FE",
		X"00",X"00",X"00",X"20",X"21",X"00",X"04",X"02",X"00",X"00",X"00",X"00",X"C0",X"78",X"3C",X"3C",
		X"02",X"04",X"00",X"21",X"20",X"00",X"00",X"00",X"3C",X"3C",X"78",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0B",X"13",X"1F",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",
		X"0F",X"12",X"0B",X"00",X"00",X"00",X"00",X"00",X"A0",X"40",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0B",X"13",X"1F",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",
		X"0F",X"12",X"0B",X"00",X"00",X"00",X"00",X"00",X"A0",X"40",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0B",X"13",X"1F",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",
		X"0F",X"12",X"0B",X"00",X"00",X"00",X"00",X"00",X"A0",X"40",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"A0",
		X"07",X"07",X"01",X"05",X"03",X"00",X"00",X"00",X"A0",X"E0",X"80",X"A0",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"A0",
		X"07",X"07",X"01",X"05",X"03",X"00",X"00",X"00",X"A0",X"E0",X"80",X"A0",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"A0",
		X"07",X"07",X"01",X"05",X"03",X"00",X"00",X"00",X"A0",X"E0",X"80",X"A0",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"07",X"07",X"0F",X"00",X"00",X"00",X"00",X"80",X"E0",X"E0",X"F0",
		X"0F",X"07",X"07",X"01",X"00",X"00",X"00",X"00",X"F0",X"E0",X"E0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",
		X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"07",X"00",X"00",X"00",X"00",X"80",X"40",X"A0",X"A0",
		X"07",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"A0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"05",X"05",X"07",X"03",X"01",X"80",X"C0",X"C0",X"E0",X"D0",X"D0",X"B0",X"B0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"30",X"30",X"10",X"10",X"10",X"10",X"00",
		X"00",X"00",X"30",X"30",X"39",X"33",X"33",X"02",X"00",X"00",X"0C",X"0C",X"9C",X"CC",X"CC",X"40",
		X"00",X"01",X"72",X"73",X"7A",X"73",X"72",X"02",X"00",X"80",X"4E",X"CE",X"5E",X"CE",X"4E",X"40",
		X"00",X"00",X"15",X"00",X"08",X"08",X"0A",X"00",X"00",X"00",X"A8",X"00",X"10",X"10",X"50",X"00",
		X"33",X"0A",X"31",X"01",X"31",X"08",X"30",X"00",X"C0",X"5C",X"80",X"8C",X"80",X"1C",X"00",X"00",
		X"00",X"10",X"10",X"10",X"10",X"00",X"03",X"10",X"00",X"00",X"08",X"08",X"08",X"00",X"C0",X"08",
		X"10",X"10",X"00",X"08",X"07",X"00",X"00",X"00",X"08",X"08",X"00",X"10",X"E0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"0D",X"1F",X"18",X"30",X"38",X"68",X"F0",X"A0",X"C0",X"00",
		X"3F",X"3F",X"3B",X"19",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"08",X"08",X"00",X"08",X"18",X"28",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"A0",X"C0",X"C0",X"A0",X"F0",X"60",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"38",X"18",X"38",X"78",X"60",X"F0",X"C0",X"E0",
		X"07",X"0F",X"0F",X"0E",X"06",X"02",X"00",X"00",X"40",X"80",X"C0",X"C0",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"10",X"10",X"20",X"60",X"40",X"80",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"C0",X"E0",X"20",X"70",X"70",X"58",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"C0",X"C0",X"70",X"70",X"28",X"38",X"30",
		X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"78",X"D8",X"F0",X"F0",X"D0",X"D0",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"C0",X"40",X"20",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"10",X"18",X"18",X"28",X"30",X"50",X"E0",
		X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"F0",X"F0",X"D0",X"F0",X"F0",X"B0",X"F0",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"40",X"E0",X"60",X"20",X"40",X"C0",X"80",X"00",
		X"01",X"03",X"05",X"03",X"01",X"01",X"03",X"07",X"F6",X"F2",X"E0",X"F0",X"F0",X"D0",X"F0",X"F0",
		X"03",X"01",X"01",X"01",X"01",X"03",X"01",X"00",X"7C",X"FE",X"F6",X"FE",X"F2",X"B0",X"F0",X"E0",
		X"00",X"00",X"00",X"00",X"60",X"F0",X"B0",X"78",X"00",X"10",X"10",X"10",X"10",X"10",X"30",X"30",
		X"1C",X"0E",X"07",X"07",X"01",X"01",X"01",X"01",X"10",X"30",X"30",X"F0",X"FC",X"3E",X"7E",X"FE",
		X"00",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",
		X"20",X"20",X"00",X"00",X"00",X"00",X"7F",X"00",X"80",X"80",X"00",X"02",X"02",X"02",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"3C",X"20",X"21",X"20",X"00",X"82",X"82",X"82",X"02",X"02",X"0E",X"08",
		X"20",X"20",X"00",X"00",X"00",X"00",X"7F",X"00",X"08",X"08",X"00",X"02",X"02",X"02",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"3F",X"20",X"20",X"20",X"00",X"08",X"00",X"02",X"F2",X"02",X"02",X"02",
		X"20",X"20",X"00",X"00",X"40",X"00",X"1F",X"00",X"02",X"02",X"02",X"02",X"0E",X"08",X"F8",X"00",
		X"00",X"30",X"70",X"B2",X"B7",X"FF",X"7F",X"1F",X"00",X"00",X"00",X"00",X"C0",X"A0",X"C0",X"E0",
		X"07",X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"60",X"00",
		X"00",X"00",X"00",X"03",X"0C",X"1C",X"1D",X"1F",X"00",X"00",X"00",X"C0",X"F0",X"F8",X"F8",X"F8",
		X"1F",X"1D",X"1C",X"0C",X"03",X"00",X"00",X"00",X"F8",X"E8",X"98",X"F0",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"07",X"18",X"2C",X"09",X"63",X"7F",X"00",X"00",X"C0",X"E0",X"F0",X"F8",X"F8",X"F8",
		X"7F",X"63",X"09",X"2C",X"18",X"07",X"00",X"00",X"F8",X"F8",X"E8",X"90",X"E0",X"C0",X"00",X"00",
		X"00",X"03",X"1F",X"37",X"23",X"60",X"61",X"7F",X"00",X"C0",X"F8",X"FC",X"FC",X"FE",X"FE",X"FE",
		X"7F",X"61",X"60",X"23",X"37",X"1F",X"03",X"00",X"FE",X"FE",X"FE",X"F4",X"CC",X"F8",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"20",X"20",X"20",X"20",X"20",X"21",X"20",X"00",X"02",X"02",X"02",X"F2",X"82",X"82",X"02",
		X"00",X"08",X"40",X"00",X"10",X"00",X"07",X"00",X"02",X"02",X"0E",X"08",X"38",X"20",X"E0",X"00",
		X"00",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"00",X"02",X"02",X"82",X"82",X"82",X"82",X"82",
		X"00",X"00",X"00",X"00",X"7F",X"00",X"00",X"00",X"02",X"02",X"02",X"02",X"FE",X"00",X"00",X"00",
		X"00",X"00",X"00",X"60",X"61",X"00",X"06",X"07",X"00",X"00",X"00",X"00",X"C0",X"78",X"3C",X"3C",
		X"07",X"06",X"00",X"21",X"20",X"00",X"00",X"00",X"3C",X"3C",X"78",X"C0",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
