library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_PGM_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_PGM_1 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"05",X"02",X"00",X"01",X"03",X"06",X"04",X"07",X"08",X"09",X"0B",X"0A",X"0C",X"0E",X"0D",X"08",
		X"0B",X"0F",X"0A",X"10",X"3C",X"80",X"5C",X"81",X"A6",X"82",X"8C",X"83",X"B2",X"84",X"F6",X"85",
		X"BE",X"86",X"02",X"88",X"28",X"89",X"8E",X"8A",X"C6",X"8B",X"44",X"8D",X"AC",X"8E",X"F6",X"8F",
		X"FE",X"90",X"10",X"92",X"7A",X"93",X"7A",X"93",X"7A",X"93",X"7A",X"93",X"01",X"05",X"0F",X"17",
		X"3B",X"17",X"01",X"14",X"0F",X"17",X"3B",X"17",X"00",X"01",X"05",X"38",X"17",X"3A",X"17",X"01",
		X"07",X"38",X"17",X"01",X"02",X"0F",X"17",X"01",X"0B",X"38",X"17",X"3A",X"17",X"38",X"17",X"00",
		X"01",X"05",X"0F",X"17",X"3B",X"17",X"01",X"14",X"0F",X"17",X"3B",X"17",X"00",X"01",X"05",X"0F",
		X"17",X"3B",X"17",X"01",X"14",X"0F",X"17",X"3B",X"17",X"00",X"01",X"05",X"0F",X"17",X"3B",X"17",
		X"01",X"02",X"0F",X"17",X"3B",X"17",X"01",X"0E",X"0F",X"17",X"3B",X"17",X"01",X"02",X"0F",X"17",
		X"3B",X"17",X"00",X"01",X"03",X"38",X"17",X"0F",X"17",X"01",X"04",X"38",X"17",X"3A",X"17",X"38",
		X"17",X"01",X"07",X"0F",X"17",X"01",X"03",X"38",X"17",X"0F",X"17",X"01",X"02",X"38",X"17",X"3A",
		X"17",X"01",X"04",X"38",X"17",X"00",X"01",X"08",X"0F",X"17",X"3B",X"17",X"01",X"0E",X"0F",X"17",
		X"3B",X"17",X"00",X"01",X"08",X"0F",X"17",X"3B",X"17",X"01",X"0E",X"0F",X"17",X"3B",X"17",X"00",
		X"01",X"03",X"0F",X"17",X"3B",X"17",X"01",X"04",X"0F",X"17",X"3B",X"17",X"01",X"0E",X"0F",X"17",
		X"3B",X"17",X"00",X"01",X"03",X"38",X"17",X"3A",X"17",X"01",X"0D",X"38",X"17",X"0F",X"17",X"01",
		X"02",X"38",X"17",X"0F",X"17",X"01",X"07",X"38",X"17",X"00",X"01",X"03",X"0F",X"17",X"3B",X"17",
		X"00",X"01",X"03",X"0F",X"17",X"3B",X"17",X"00",X"01",X"03",X"0F",X"17",X"3B",X"17",X"01",X"02",
		X"0F",X"17",X"3B",X"17",X"01",X"10",X"0F",X"17",X"3B",X"17",X"00",X"01",X"06",X"38",X"17",X"3A",
		X"17",X"01",X"03",X"38",X"17",X"01",X"07",X"0F",X"17",X"01",X"06",X"38",X"17",X"3A",X"17",X"01",
		X"04",X"38",X"17",X"00",X"01",X"06",X"0F",X"17",X"3B",X"17",X"01",X"10",X"0F",X"17",X"3B",X"17",
		X"00",X"01",X"06",X"0F",X"17",X"3B",X"17",X"01",X"10",X"0F",X"17",X"3B",X"17",X"00",X"01",X"06",
		X"0F",X"17",X"3B",X"17",X"01",X"10",X"0F",X"17",X"3B",X"17",X"00",X"FF",X"01",X"02",X"0F",X"17",
		X"3B",X"17",X"01",X"17",X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",X"38",X"17",X"3A",X"17",X"01",
		X"05",X"38",X"17",X"0F",X"17",X"01",X"03",X"38",X"17",X"01",X"04",X"0F",X"17",X"01",X"04",X"38",
		X"17",X"0F",X"17",X"01",X"03",X"38",X"17",X"0F",X"17",X"38",X"17",X"3A",X"17",X"38",X"17",X"00",
		X"01",X"02",X"0F",X"17",X"3B",X"17",X"01",X"17",X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",X"0F",
		X"17",X"3B",X"17",X"01",X"17",X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",X"0F",X"17",X"3B",X"17",
		X"01",X"03",X"0F",X"17",X"3B",X"17",X"01",X"0E",X"0F",X"17",X"3B",X"17",X"01",X"04",X"0F",X"17",
		X"3B",X"17",X"00",X"01",X"06",X"38",X"17",X"3A",X"17",X"01",X"04",X"38",X"17",X"0F",X"17",X"01",
		X"03",X"38",X"17",X"01",X"03",X"0F",X"17",X"01",X"03",X"38",X"17",X"3A",X"17",X"38",X"17",X"0F",
		X"17",X"01",X"04",X"38",X"17",X"00",X"01",X"06",X"0F",X"17",X"3B",X"17",X"01",X"0E",X"0F",X"17",
		X"3B",X"17",X"00",X"01",X"06",X"0F",X"17",X"3B",X"17",X"01",X"0E",X"0F",X"17",X"3B",X"17",X"00",
		X"01",X"02",X"0F",X"17",X"3B",X"17",X"01",X"03",X"0F",X"17",X"3B",X"17",X"01",X"0E",X"0F",X"17",
		X"3B",X"17",X"01",X"02",X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",X"38",X"17",X"3A",X"17",X"01",
		X"0A",X"38",X"17",X"01",X"04",X"0F",X"17",X"01",X"07",X"38",X"17",X"3A",X"17",X"01",X"03",X"38",
		X"17",X"00",X"01",X"02",X"0F",X"17",X"3B",X"17",X"01",X"15",X"0F",X"17",X"3B",X"17",X"00",X"01",
		X"02",X"0F",X"17",X"3B",X"17",X"01",X"15",X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",X"0F",X"17",
		X"3B",X"17",X"01",X"05",X"0F",X"17",X"3B",X"17",X"01",X"0A",X"0F",X"17",X"3B",X"17",X"01",X"04",
		X"0F",X"17",X"3B",X"17",X"00",X"01",X"08",X"38",X"17",X"3A",X"17",X"01",X"04",X"38",X"17",X"01",
		X"03",X"0F",X"17",X"01",X"03",X"38",X"17",X"3A",X"17",X"01",X"08",X"38",X"17",X"00",X"01",X"08",
		X"0F",X"17",X"3B",X"17",X"01",X"0A",X"0F",X"17",X"3B",X"17",X"00",X"01",X"08",X"0F",X"17",X"3B",
		X"17",X"01",X"0A",X"0F",X"17",X"3B",X"17",X"00",X"01",X"08",X"0F",X"17",X"3B",X"17",X"01",X"0A",
		X"0F",X"17",X"3B",X"17",X"00",X"FF",X"01",X"06",X"0F",X"17",X"3B",X"17",X"00",X"01",X"03",X"38",
		X"17",X"0F",X"17",X"01",X"02",X"38",X"17",X"3A",X"17",X"01",X"02",X"38",X"17",X"01",X"02",X"0F",
		X"17",X"01",X"02",X"38",X"17",X"01",X"02",X"0F",X"17",X"01",X"02",X"38",X"17",X"0F",X"17",X"01",
		X"0A",X"38",X"17",X"00",X"01",X"06",X"0F",X"17",X"3B",X"17",X"00",X"01",X"06",X"0F",X"17",X"3B",
		X"17",X"00",X"01",X"06",X"0F",X"17",X"3B",X"17",X"01",X"0A",X"0F",X"17",X"3B",X"17",X"00",X"01",
		X"09",X"38",X"17",X"0F",X"17",X"01",X"07",X"38",X"17",X"3A",X"17",X"01",X"06",X"38",X"17",X"0F",
		X"17",X"01",X"03",X"38",X"17",X"00",X"01",X"11",X"0F",X"17",X"3B",X"17",X"00",X"01",X"11",X"0F",
		X"17",X"3B",X"17",X"00",X"01",X"06",X"0F",X"17",X"3B",X"17",X"01",X"0A",X"0F",X"17",X"3B",X"17",
		X"00",X"01",X"06",X"38",X"17",X"3A",X"17",X"01",X"04",X"38",X"17",X"0F",X"17",X"01",X"08",X"38",
		X"17",X"0F",X"17",X"01",X"02",X"38",X"17",X"0F",X"17",X"01",X"04",X"38",X"17",X"00",X"01",X"06",
		X"0F",X"17",X"3B",X"17",X"00",X"01",X"06",X"0F",X"17",X"3B",X"17",X"00",X"01",X"06",X"0F",X"17",
		X"3B",X"17",X"01",X"08",X"0F",X"17",X"3B",X"17",X"00",X"01",X"03",X"38",X"17",X"0F",X"17",X"01",
		X"06",X"38",X"17",X"0F",X"17",X"01",X"04",X"38",X"17",X"3A",X"17",X"01",X"08",X"38",X"17",X"0F",
		X"17",X"01",X"03",X"38",X"17",X"00",X"01",X"0F",X"0F",X"17",X"3B",X"17",X"00",X"01",X"0F",X"0F",
		X"17",X"3B",X"17",X"00",X"01",X"0F",X"0F",X"17",X"3B",X"17",X"00",X"FF",X"01",X"02",X"0F",X"17",
		X"3B",X"17",X"01",X"14",X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",X"38",X"17",X"3A",X"17",X"01",
		X"09",X"38",X"17",X"01",X"03",X"0F",X"17",X"01",X"02",X"38",X"17",X"01",X"02",X"0F",X"17",X"01",
		X"04",X"38",X"17",X"3A",X"17",X"01",X"04",X"38",X"17",X"00",X"01",X"02",X"0F",X"17",X"3B",X"17",
		X"01",X"14",X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",X"0F",X"17",X"3B",X"17",X"01",X"14",X"0F",
		X"17",X"3B",X"17",X"00",X"01",X"02",X"0F",X"17",X"3B",X"17",X"0F",X"17",X"3B",X"17",X"01",X"10",
		X"0F",X"17",X"3B",X"17",X"0F",X"17",X"3B",X"17",X"00",X"01",X"04",X"38",X"17",X"3A",X"17",X"01",
		X"05",X"38",X"17",X"01",X"07",X"0F",X"17",X"01",X"04",X"38",X"17",X"3A",X"17",X"01",X"06",X"38",
		X"17",X"00",X"01",X"04",X"0F",X"17",X"3B",X"17",X"01",X"10",X"0F",X"17",X"3B",X"17",X"00",X"01",
		X"04",X"0F",X"17",X"3B",X"17",X"01",X"10",X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",X"0F",X"17",
		X"3B",X"17",X"0F",X"17",X"3B",X"17",X"01",X"10",X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",X"38",
		X"17",X"3A",X"17",X"01",X"03",X"38",X"17",X"0F",X"17",X"01",X"02",X"38",X"17",X"0F",X"17",X"01",
		X"02",X"38",X"17",X"0F",X"17",X"01",X"0B",X"38",X"17",X"0F",X"17",X"01",X"03",X"38",X"17",X"00",
		X"01",X"02",X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",
		X"0F",X"17",X"3B",X"17",X"01",X"06",X"0F",X"17",X"3B",X"17",X"01",X"0D",X"0F",X"17",X"3B",X"17",
		X"00",X"01",X"09",X"38",X"17",X"3A",X"17",X"01",X"02",X"38",X"17",X"01",X"05",X"0F",X"17",X"01",
		X"06",X"38",X"17",X"3A",X"17",X"01",X"04",X"38",X"17",X"00",X"01",X"09",X"0F",X"17",X"3B",X"17",
		X"01",X"0D",X"0F",X"17",X"3B",X"17",X"00",X"01",X"09",X"0F",X"17",X"3B",X"17",X"01",X"0D",X"0F",
		X"17",X"3B",X"17",X"00",X"01",X"09",X"0F",X"17",X"3B",X"17",X"01",X"0D",X"0F",X"17",X"3B",X"17",
		X"00",X"FF",X"01",X"08",X"0F",X"17",X"3B",X"17",X"01",X"11",X"0F",X"17",X"3B",X"17",X"00",X"01",
		X"08",X"38",X"17",X"3A",X"17",X"38",X"17",X"01",X"08",X"0F",X"17",X"01",X"03",X"38",X"17",X"0F",
		X"17",X"01",X"02",X"38",X"17",X"0F",X"17",X"38",X"17",X"3A",X"17",X"38",X"17",X"00",X"01",X"08",
		X"0F",X"17",X"3B",X"17",X"01",X"11",X"0F",X"17",X"3B",X"17",X"00",X"01",X"08",X"0F",X"17",X"3B",
		X"17",X"01",X"11",X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",X"0F",X"17",X"3B",X"17",X"01",X"05",
		X"0F",X"17",X"3B",X"17",X"01",X"0A",X"0F",X"17",X"3B",X"17",X"01",X"06",X"0F",X"17",X"3B",X"17",
		X"00",X"01",X"02",X"38",X"17",X"3A",X"17",X"38",X"17",X"0F",X"17",X"01",X"05",X"38",X"17",X"0F",
		X"17",X"01",X"03",X"38",X"17",X"01",X"04",X"0F",X"17",X"38",X"17",X"3A",X"17",X"01",X"03",X"38",
		X"17",X"0F",X"17",X"01",X"04",X"38",X"17",X"00",X"01",X"02",X"0F",X"17",X"3B",X"17",X"01",X"10",
		X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",X"0F",X"17",X"3B",X"17",X"01",X"10",X"0F",X"17",X"3B",
		X"17",X"00",X"01",X"02",X"0F",X"17",X"3B",X"17",X"01",X"06",X"0F",X"17",X"3B",X"17",X"01",X"09",
		X"0F",X"17",X"3B",X"17",X"01",X"04",X"0F",X"17",X"3B",X"17",X"00",X"01",X"09",X"38",X"17",X"3A",
		X"17",X"38",X"17",X"01",X"07",X"0F",X"17",X"01",X"06",X"38",X"17",X"3A",X"17",X"01",X"03",X"38",
		X"17",X"00",X"01",X"09",X"0F",X"17",X"3B",X"17",X"01",X"0E",X"0F",X"17",X"3B",X"17",X"00",X"01",
		X"09",X"0F",X"17",X"3B",X"17",X"01",X"0E",X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",X"0F",X"17",
		X"3B",X"17",X"01",X"06",X"0F",X"17",X"3B",X"17",X"01",X"09",X"0F",X"17",X"3B",X"17",X"01",X"04",
		X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",X"38",X"17",X"3A",X"17",X"01",X"0A",X"38",X"17",X"01",
		X"03",X"0F",X"17",X"01",X"03",X"38",X"17",X"3A",X"17",X"01",X"08",X"38",X"17",X"00",X"01",X"02",
		X"0F",X"17",X"3B",X"17",X"01",X"10",X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",X"0F",X"17",X"3B",
		X"17",X"01",X"10",X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",X"0F",X"17",X"3B",X"17",X"01",X"10",
		X"0F",X"17",X"3B",X"17",X"00",X"FF",X"01",X"0B",X"0F",X"17",X"3B",X"17",X"00",X"01",X"03",X"38",
		X"17",X"0F",X"17",X"01",X"04",X"38",X"17",X"0F",X"17",X"01",X"02",X"38",X"17",X"3A",X"17",X"01",
		X"02",X"38",X"17",X"0F",X"17",X"01",X"0D",X"38",X"17",X"00",X"01",X"0B",X"0F",X"17",X"3B",X"17",
		X"00",X"01",X"0B",X"0F",X"17",X"3B",X"17",X"00",X"01",X"0B",X"0F",X"17",X"3B",X"17",X"01",X"05",
		X"0F",X"17",X"3B",X"17",X"00",X"01",X"07",X"38",X"17",X"0F",X"17",X"01",X"09",X"38",X"17",X"3A",
		X"17",X"01",X"06",X"38",X"17",X"0F",X"17",X"01",X"03",X"38",X"17",X"00",X"01",X"11",X"0F",X"17",
		X"3B",X"17",X"00",X"01",X"11",X"0F",X"17",X"3B",X"17",X"00",X"01",X"11",X"0F",X"17",X"3B",X"17",
		X"01",X"04",X"0F",X"17",X"3B",X"17",X"00",X"01",X"06",X"38",X"17",X"0F",X"17",X"01",X"0D",X"38",
		X"17",X"0F",X"17",X"38",X"17",X"3A",X"17",X"01",X"05",X"38",X"17",X"00",X"01",X"16",X"0F",X"17",
		X"3B",X"17",X"00",X"01",X"16",X"0F",X"17",X"3B",X"17",X"00",X"01",X"0F",X"0F",X"17",X"3B",X"17",
		X"01",X"06",X"0F",X"17",X"3B",X"17",X"00",X"01",X"09",X"38",X"17",X"0F",X"17",X"01",X"05",X"38",
		X"17",X"3A",X"17",X"01",X"0C",X"38",X"17",X"00",X"01",X"0F",X"0F",X"17",X"3B",X"17",X"00",X"01",
		X"0F",X"0F",X"17",X"3B",X"17",X"00",X"01",X"0F",X"0F",X"17",X"3B",X"17",X"00",X"FF",X"01",X"04",
		X"0F",X"17",X"3B",X"17",X"01",X"0D",X"0F",X"17",X"3B",X"17",X"00",X"01",X"04",X"38",X"17",X"3A",
		X"17",X"01",X"03",X"38",X"17",X"0F",X"17",X"01",X"03",X"38",X"17",X"01",X"04",X"0F",X"17",X"01",
		X"02",X"38",X"17",X"3A",X"17",X"01",X"09",X"38",X"17",X"00",X"01",X"04",X"0F",X"17",X"3B",X"17",
		X"01",X"0D",X"0F",X"17",X"3B",X"17",X"00",X"01",X"04",X"0F",X"17",X"3B",X"17",X"01",X"0D",X"0F",
		X"17",X"3B",X"17",X"00",X"01",X"04",X"0F",X"17",X"3B",X"17",X"01",X"07",X"0F",X"17",X"3B",X"17",
		X"01",X"05",X"0F",X"17",X"3B",X"17",X"01",X"07",X"0F",X"17",X"3B",X"17",X"00",X"01",X"0A",X"38",
		X"17",X"0F",X"17",X"38",X"17",X"3A",X"17",X"38",X"17",X"01",X"03",X"0F",X"17",X"01",X"04",X"38",
		X"17",X"0F",X"17",X"01",X"02",X"38",X"17",X"0F",X"17",X"38",X"17",X"3A",X"17",X"38",X"17",X"00",
		X"01",X"0C",X"0F",X"17",X"3B",X"17",X"01",X"0D",X"0F",X"17",X"3B",X"17",X"00",X"01",X"0C",X"0F",
		X"17",X"3B",X"17",X"01",X"0D",X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",X"0F",X"17",X"3B",X"17",
		X"01",X"09",X"0F",X"17",X"3B",X"17",X"01",X"04",X"0F",X"17",X"3B",X"17",X"01",X"08",X"0F",X"17",
		X"3B",X"17",X"00",X"01",X"02",X"38",X"17",X"3A",X"17",X"01",X"02",X"38",X"17",X"01",X"02",X"0F",
		X"17",X"01",X"07",X"38",X"17",X"01",X"02",X"0F",X"17",X"38",X"17",X"3A",X"17",X"01",X"03",X"38",
		X"17",X"0F",X"17",X"01",X"06",X"38",X"17",X"00",X"01",X"02",X"0F",X"17",X"3B",X"17",X"01",X"0E",
		X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",X"0F",X"17",X"3B",X"17",X"01",X"0E",X"0F",X"17",X"3B",
		X"17",X"00",X"01",X"02",X"0F",X"17",X"3B",X"17",X"01",X"06",X"0F",X"17",X"3B",X"17",X"01",X"07",
		X"0F",X"17",X"3B",X"17",X"00",X"01",X"05",X"38",X"17",X"0F",X"17",X"01",X"03",X"38",X"17",X"3A",
		X"17",X"01",X"03",X"38",X"17",X"01",X"03",X"0F",X"17",X"01",X"03",X"38",X"17",X"0F",X"17",X"01",
		X"02",X"38",X"17",X"01",X"02",X"0F",X"17",X"01",X"04",X"38",X"17",X"00",X"01",X"09",X"0F",X"17",
		X"3B",X"17",X"00",X"01",X"09",X"0F",X"17",X"3B",X"17",X"00",X"01",X"09",X"0F",X"17",X"3B",X"17",
		X"00",X"FF",X"01",X"09",X"0F",X"17",X"3B",X"17",X"00",X"01",X"03",X"38",X"17",X"0F",X"17",X"01",
		X"02",X"38",X"17",X"0F",X"17",X"01",X"02",X"38",X"17",X"3A",X"17",X"01",X"02",X"38",X"17",X"0F",
		X"17",X"01",X"02",X"38",X"17",X"01",X"02",X"0F",X"17",X"01",X"02",X"38",X"17",X"0F",X"17",X"01",
		X"08",X"38",X"17",X"00",X"01",X"09",X"0F",X"17",X"3B",X"17",X"00",X"01",X"09",X"0F",X"17",X"3B",
		X"17",X"00",X"01",X"02",X"0F",X"17",X"3B",X"17",X"01",X"06",X"0F",X"17",X"3B",X"17",X"01",X"10",
		X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",X"38",X"17",X"3A",X"17",X"01",X"08",X"38",X"17",X"0F",
		X"17",X"01",X"02",X"38",X"17",X"0F",X"17",X"01",X"02",X"38",X"17",X"01",X"02",X"0F",X"17",X"01",
		X"03",X"38",X"17",X"01",X"02",X"0F",X"17",X"01",X"02",X"38",X"17",X"3A",X"17",X"38",X"17",X"00",
		X"01",X"02",X"0F",X"17",X"3B",X"17",X"01",X"17",X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",X"0F",
		X"17",X"3B",X"17",X"01",X"17",X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",X"0F",X"17",X"3B",X"17",
		X"01",X"0F",X"0F",X"17",X"3B",X"17",X"01",X"07",X"0F",X"17",X"3B",X"17",X"00",X"01",X"07",X"38",
		X"17",X"0F",X"17",X"01",X"04",X"38",X"17",X"0F",X"17",X"01",X"05",X"38",X"17",X"3A",X"17",X"01",
		X"09",X"38",X"17",X"00",X"01",X"12",X"0F",X"17",X"3B",X"17",X"00",X"01",X"12",X"0F",X"17",X"3B",
		X"17",X"00",X"01",X"0D",X"0F",X"17",X"3B",X"17",X"01",X"04",X"0F",X"17",X"3B",X"17",X"00",X"01",
		X"03",X"38",X"17",X"01",X"02",X"0F",X"17",X"01",X"02",X"38",X"17",X"0F",X"17",X"01",X"02",X"38",
		X"17",X"01",X"02",X"0F",X"17",X"38",X"17",X"3A",X"17",X"01",X"02",X"38",X"17",X"0F",X"17",X"01",
		X"03",X"38",X"17",X"01",X"02",X"0F",X"17",X"01",X"02",X"38",X"17",X"0F",X"17",X"01",X"03",X"38",
		X"17",X"00",X"01",X"0D",X"0F",X"17",X"3B",X"17",X"00",X"01",X"0D",X"0F",X"17",X"3B",X"17",X"00",
		X"01",X"0D",X"0F",X"17",X"3B",X"17",X"00",X"FF",X"01",X"09",X"0F",X"17",X"3B",X"17",X"01",X"10",
		X"0F",X"17",X"3B",X"17",X"00",X"01",X"03",X"38",X"17",X"01",X"02",X"0F",X"17",X"01",X"02",X"38",
		X"17",X"0F",X"17",X"38",X"17",X"3A",X"17",X"38",X"17",X"01",X"04",X"0F",X"17",X"01",X"0B",X"38",
		X"17",X"3A",X"17",X"38",X"17",X"00",X"01",X"09",X"0F",X"17",X"3B",X"17",X"01",X"10",X"0F",X"17",
		X"3B",X"17",X"00",X"01",X"09",X"0F",X"17",X"3B",X"17",X"01",X"10",X"0F",X"17",X"3B",X"17",X"00",
		X"01",X"02",X"0F",X"17",X"3B",X"17",X"01",X"06",X"0F",X"17",X"3B",X"17",X"01",X"06",X"0F",X"17",
		X"3B",X"17",X"01",X"09",X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",X"38",X"17",X"3A",X"17",X"38",
		X"17",X"0F",X"17",X"01",X"02",X"38",X"17",X"0F",X"17",X"01",X"03",X"38",X"17",X"0F",X"17",X"01",
		X"02",X"38",X"17",X"0F",X"17",X"38",X"17",X"3A",X"17",X"38",X"17",X"0F",X"17",X"01",X"02",X"38",
		X"17",X"0F",X"17",X"01",X"02",X"38",X"17",X"0F",X"17",X"01",X"03",X"38",X"17",X"00",X"01",X"02",
		X"0F",X"17",X"3B",X"17",X"01",X"0D",X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",X"0F",X"17",X"3B",
		X"17",X"01",X"0D",X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",X"0F",X"17",X"01",X"02",X"3B",X"17",
		X"01",X"0C",X"0F",X"17",X"3B",X"17",X"01",X"09",X"0F",X"17",X"3B",X"17",X"00",X"01",X"03",X"38",
		X"17",X"3A",X"17",X"38",X"17",X"0F",X"17",X"01",X"03",X"38",X"17",X"0F",X"17",X"01",X"02",X"38",
		X"17",X"01",X"03",X"0F",X"17",X"01",X"03",X"38",X"17",X"0F",X"17",X"01",X"05",X"38",X"17",X"0F",
		X"17",X"38",X"17",X"3A",X"17",X"38",X"17",X"00",X"01",X"03",X"0F",X"17",X"3B",X"17",X"01",X"16",
		X"0F",X"17",X"3B",X"17",X"00",X"01",X"03",X"0F",X"17",X"3B",X"17",X"01",X"16",X"0F",X"17",X"3B",
		X"17",X"00",X"01",X"03",X"0F",X"17",X"3B",X"17",X"01",X"04",X"0F",X"17",X"3B",X"17",X"01",X"0C",
		X"0F",X"17",X"3B",X"17",X"01",X"04",X"0F",X"17",X"3B",X"17",X"00",X"01",X"08",X"38",X"17",X"3A",
		X"17",X"38",X"17",X"01",X"05",X"0F",X"17",X"01",X"04",X"38",X"17",X"0F",X"17",X"38",X"17",X"3A",
		X"17",X"01",X"06",X"38",X"17",X"00",X"01",X"08",X"0F",X"17",X"3B",X"17",X"01",X"0C",X"0F",X"17",
		X"3B",X"17",X"00",X"01",X"08",X"0F",X"17",X"3B",X"17",X"01",X"0C",X"0F",X"17",X"3B",X"17",X"00",
		X"01",X"08",X"0F",X"17",X"3B",X"17",X"01",X"0C",X"0F",X"17",X"3B",X"17",X"00",X"FF",X"01",X"04",
		X"0F",X"17",X"3B",X"17",X"01",X"15",X"0F",X"17",X"3B",X"17",X"00",X"01",X"04",X"38",X"17",X"3A",
		X"17",X"01",X"08",X"38",X"17",X"0F",X"17",X"01",X"0A",X"38",X"17",X"0F",X"17",X"38",X"17",X"3A",
		X"17",X"38",X"17",X"00",X"01",X"04",X"0F",X"17",X"3B",X"17",X"01",X"15",X"0F",X"17",X"3B",X"17",
		X"00",X"01",X"04",X"0F",X"17",X"3B",X"17",X"01",X"15",X"0F",X"17",X"3B",X"17",X"00",X"01",X"04",
		X"0F",X"17",X"3B",X"17",X"01",X"08",X"0F",X"17",X"3B",X"17",X"01",X"0C",X"0F",X"17",X"3B",X"17",
		X"00",X"01",X"06",X"38",X"17",X"01",X"03",X"0F",X"17",X"01",X"04",X"38",X"17",X"3A",X"17",X"38",
		X"17",X"01",X"02",X"0F",X"17",X"01",X"03",X"38",X"17",X"01",X"02",X"0F",X"17",X"01",X"06",X"38",
		X"17",X"00",X"01",X"0D",X"0F",X"17",X"3B",X"17",X"00",X"01",X"0D",X"0F",X"17",X"3B",X"17",X"00",
		X"01",X"02",X"0F",X"17",X"3B",X"17",X"01",X"0A",X"0F",X"17",X"3B",X"17",X"01",X"0C",X"0F",X"17",
		X"3B",X"17",X"00",X"01",X"02",X"38",X"17",X"3A",X"17",X"01",X"04",X"38",X"17",X"0F",X"17",X"01",
		X"0A",X"38",X"17",X"01",X"02",X"0F",X"17",X"01",X"04",X"38",X"17",X"0F",X"17",X"38",X"17",X"3A",
		X"17",X"38",X"17",X"00",X"01",X"02",X"0F",X"17",X"3B",X"17",X"01",X"17",X"0F",X"17",X"3B",X"17",
		X"00",X"01",X"02",X"0F",X"17",X"3B",X"17",X"01",X"17",X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",
		X"0F",X"17",X"3B",X"17",X"01",X"03",X"0F",X"17",X"3B",X"17",X"01",X"0C",X"0F",X"17",X"3B",X"17",
		X"01",X"06",X"0F",X"17",X"3B",X"17",X"00",X"01",X"04",X"38",X"17",X"0F",X"17",X"38",X"17",X"3A",
		X"17",X"01",X"06",X"38",X"17",X"01",X"02",X"0F",X"17",X"01",X"02",X"38",X"17",X"0F",X"17",X"38",
		X"17",X"3A",X"17",X"01",X"04",X"38",X"17",X"0F",X"17",X"01",X"03",X"38",X"17",X"00",X"01",X"06",
		X"0F",X"17",X"3B",X"17",X"01",X"0C",X"0F",X"17",X"3B",X"17",X"00",X"01",X"06",X"0F",X"17",X"3B",
		X"17",X"01",X"0C",X"0F",X"17",X"3B",X"17",X"00",X"01",X"06",X"0F",X"17",X"3B",X"17",X"01",X"0C",
		X"0F",X"17",X"3B",X"17",X"00",X"FF",X"01",X"02",X"0F",X"17",X"3B",X"17",X"01",X"0F",X"0F",X"17",
		X"3B",X"17",X"00",X"01",X"02",X"38",X"17",X"3A",X"17",X"38",X"17",X"0F",X"17",X"01",X"02",X"38",
		X"17",X"0F",X"17",X"01",X"02",X"38",X"17",X"0F",X"17",X"01",X"02",X"38",X"17",X"01",X"04",X"0F",
		X"17",X"38",X"17",X"3A",X"17",X"01",X"09",X"38",X"17",X"00",X"01",X"02",X"0F",X"17",X"3B",X"17",
		X"01",X"0F",X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",X"0F",X"17",X"3B",X"17",X"01",X"0F",X"0F",
		X"17",X"3B",X"17",X"00",X"01",X"02",X"0F",X"17",X"3B",X"17",X"01",X"07",X"0F",X"17",X"3B",X"17",
		X"01",X"07",X"0F",X"17",X"3B",X"17",X"01",X"07",X"0F",X"17",X"3B",X"17",X"00",X"01",X"04",X"38",
		X"17",X"0F",X"17",X"01",X"02",X"38",X"17",X"01",X"02",X"0F",X"17",X"38",X"17",X"3A",X"17",X"38",
		X"17",X"01",X"03",X"0F",X"17",X"01",X"05",X"38",X"17",X"01",X"02",X"0F",X"17",X"01",X"02",X"38",
		X"17",X"0F",X"17",X"38",X"17",X"3A",X"17",X"38",X"17",X"00",X"01",X"0A",X"0F",X"17",X"3B",X"17",
		X"01",X"0F",X"0F",X"17",X"3B",X"17",X"00",X"01",X"0A",X"0F",X"17",X"3B",X"17",X"01",X"0F",X"0F",
		X"17",X"3B",X"17",X"00",X"01",X"09",X"0F",X"17",X"01",X"02",X"3B",X"17",X"01",X"08",X"0F",X"17",
		X"3B",X"17",X"01",X"06",X"0F",X"17",X"3B",X"17",X"00",X"01",X"03",X"38",X"17",X"0F",X"17",X"01",
		X"03",X"38",X"17",X"0F",X"17",X"38",X"17",X"3A",X"17",X"01",X"02",X"38",X"17",X"01",X"04",X"0F",
		X"17",X"01",X"03",X"38",X"17",X"3A",X"17",X"38",X"17",X"0F",X"17",X"01",X"02",X"38",X"17",X"0F",
		X"17",X"01",X"03",X"38",X"17",X"00",X"01",X"09",X"0F",X"17",X"3B",X"17",X"01",X"09",X"0F",X"17",
		X"3B",X"17",X"00",X"01",X"09",X"0F",X"17",X"3B",X"17",X"01",X"09",X"0F",X"17",X"3B",X"17",X"00",
		X"01",X"02",X"0F",X"17",X"3B",X"17",X"01",X"06",X"0F",X"17",X"3B",X"17",X"01",X"09",X"0F",X"17",
		X"3B",X"17",X"01",X"05",X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",X"38",X"17",X"3A",X"17",X"38",
		X"17",X"0F",X"17",X"01",X"02",X"38",X"17",X"0F",X"17",X"01",X"03",X"38",X"17",X"0F",X"17",X"38",
		X"17",X"0F",X"17",X"38",X"17",X"0F",X"17",X"38",X"17",X"0F",X"17",X"01",X"03",X"38",X"17",X"0F",
		X"17",X"01",X"03",X"38",X"17",X"3A",X"17",X"01",X"02",X"38",X"17",X"00",X"01",X"02",X"0F",X"17",
		X"3B",X"17",X"01",X"16",X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",X"0F",X"17",X"3B",X"17",X"01",
		X"16",X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",X"0F",X"17",X"3B",X"17",X"01",X"16",X"0F",X"17",
		X"3B",X"17",X"00",X"FF",X"01",X"02",X"0F",X"17",X"3B",X"17",X"01",X"15",X"0F",X"17",X"3B",X"17",
		X"00",X"01",X"02",X"38",X"17",X"3A",X"17",X"01",X"02",X"38",X"17",X"01",X"02",X"0F",X"17",X"01",
		X"03",X"38",X"17",X"0F",X"17",X"38",X"17",X"01",X"03",X"0F",X"17",X"38",X"17",X"0F",X"17",X"01",
		X"02",X"38",X"17",X"0F",X"17",X"01",X"02",X"38",X"17",X"0F",X"17",X"38",X"17",X"3A",X"17",X"01",
		X"03",X"38",X"17",X"00",X"01",X"02",X"0F",X"17",X"3B",X"17",X"01",X"15",X"0F",X"17",X"3B",X"17",
		X"00",X"01",X"02",X"0F",X"17",X"3B",X"17",X"01",X"15",X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",
		X"0F",X"17",X"3B",X"17",X"01",X"05",X"0F",X"17",X"3B",X"17",X"01",X"0F",X"0F",X"17",X"3B",X"17",
		X"0F",X"17",X"3B",X"17",X"00",X"01",X"06",X"38",X"17",X"0F",X"17",X"38",X"17",X"3A",X"17",X"38",
		X"17",X"01",X"03",X"0F",X"17",X"38",X"17",X"01",X"03",X"0F",X"17",X"01",X"02",X"38",X"17",X"0F",
		X"17",X"01",X"02",X"38",X"17",X"0F",X"17",X"01",X"03",X"38",X"17",X"3A",X"17",X"38",X"17",X"00",
		X"01",X"08",X"0F",X"17",X"3B",X"17",X"01",X"11",X"0F",X"17",X"3B",X"17",X"00",X"01",X"08",X"0F",
		X"17",X"3B",X"17",X"01",X"11",X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",X"0F",X"17",X"3B",X"17",
		X"01",X"05",X"0F",X"17",X"3B",X"17",X"01",X"0F",X"0F",X"17",X"3B",X"17",X"0F",X"17",X"3B",X"17",
		X"00",X"01",X"02",X"38",X"17",X"3A",X"17",X"01",X"03",X"38",X"17",X"0F",X"17",X"01",X"05",X"38",
		X"17",X"01",X"03",X"0F",X"17",X"01",X"03",X"38",X"17",X"0F",X"17",X"01",X"02",X"38",X"17",X"01",
		X"02",X"0F",X"17",X"38",X"17",X"3A",X"17",X"01",X"03",X"38",X"17",X"00",X"01",X"02",X"0F",X"17",
		X"3B",X"17",X"01",X"15",X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",X"0F",X"17",X"3B",X"17",X"01",
		X"15",X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",X"0F",X"17",X"3B",X"17",X"01",X"06",X"0F",X"17",
		X"3B",X"17",X"01",X"07",X"0F",X"17",X"3B",X"17",X"01",X"06",X"0F",X"17",X"3B",X"17",X"00",X"01",
		X"09",X"38",X"17",X"3A",X"17",X"38",X"17",X"01",X"05",X"0F",X"17",X"38",X"17",X"3A",X"17",X"01",
		X"0A",X"38",X"17",X"00",X"01",X"09",X"0F",X"17",X"3B",X"17",X"01",X"07",X"0F",X"17",X"3B",X"17",
		X"00",X"01",X"09",X"0F",X"17",X"3B",X"17",X"01",X"07",X"0F",X"17",X"3B",X"17",X"00",X"01",X"09",
		X"0F",X"17",X"3B",X"17",X"01",X"07",X"0F",X"17",X"3B",X"17",X"00",X"FF",X"01",X"03",X"0F",X"17",
		X"3B",X"17",X"00",X"01",X"03",X"38",X"17",X"3A",X"17",X"01",X"02",X"38",X"17",X"0F",X"17",X"38",
		X"17",X"0F",X"17",X"38",X"17",X"0F",X"17",X"38",X"17",X"0F",X"17",X"01",X"03",X"38",X"17",X"0F",
		X"17",X"38",X"17",X"0F",X"17",X"01",X"04",X"38",X"17",X"0F",X"17",X"01",X"04",X"38",X"17",X"00",
		X"01",X"03",X"0F",X"17",X"3B",X"17",X"00",X"01",X"03",X"0F",X"17",X"3B",X"17",X"00",X"01",X"03",
		X"0F",X"17",X"3B",X"17",X"01",X"07",X"0F",X"17",X"3B",X"17",X"01",X"08",X"0F",X"17",X"3B",X"17",
		X"00",X"01",X"05",X"38",X"17",X"0F",X"17",X"38",X"17",X"0F",X"17",X"01",X"03",X"38",X"17",X"3A",
		X"17",X"38",X"17",X"01",X"03",X"0F",X"17",X"01",X"02",X"38",X"17",X"0F",X"17",X"38",X"17",X"3A",
		X"17",X"01",X"03",X"38",X"17",X"0F",X"17",X"01",X"03",X"38",X"17",X"00",X"01",X"0B",X"0F",X"17",
		X"3B",X"17",X"01",X"08",X"0F",X"17",X"3B",X"17",X"00",X"01",X"0B",X"0F",X"17",X"3B",X"17",X"01",
		X"08",X"0F",X"17",X"3B",X"17",X"00",X"01",X"0B",X"0F",X"17",X"3B",X"17",X"01",X"08",X"0F",X"17",
		X"3B",X"17",X"01",X"05",X"0F",X"17",X"3B",X"17",X"00",X"01",X"07",X"38",X"17",X"0F",X"17",X"38",
		X"17",X"0F",X"17",X"01",X"04",X"38",X"17",X"01",X"05",X"0F",X"17",X"01",X"04",X"38",X"17",X"01",
		X"02",X"0F",X"17",X"38",X"17",X"3A",X"17",X"38",X"17",X"00",X"01",X"1A",X"0F",X"17",X"3B",X"17",
		X"00",X"01",X"1A",X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",X"0F",X"17",X"3B",X"17",X"01",X"16",
		X"0F",X"17",X"01",X"02",X"3B",X"17",X"00",X"01",X"02",X"38",X"17",X"3A",X"17",X"38",X"17",X"0F",
		X"17",X"01",X"03",X"38",X"17",X"0F",X"17",X"38",X"17",X"0F",X"17",X"38",X"17",X"01",X"02",X"0F",
		X"17",X"01",X"02",X"38",X"17",X"0F",X"17",X"38",X"17",X"0F",X"17",X"01",X"02",X"38",X"17",X"0F",
		X"17",X"38",X"17",X"0F",X"17",X"38",X"17",X"3A",X"17",X"01",X"02",X"38",X"17",X"00",X"01",X"02",
		X"0F",X"17",X"3B",X"17",X"01",X"16",X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",X"0F",X"17",X"3B",
		X"17",X"01",X"16",X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",X"0F",X"17",X"3B",X"17",X"01",X"16",
		X"0F",X"17",X"3B",X"17",X"00",X"FF",X"01",X"12",X"0F",X"17",X"3B",X"17",X"00",X"01",X"07",X"38",
		X"17",X"0F",X"17",X"38",X"17",X"01",X"03",X"0F",X"17",X"38",X"17",X"0F",X"17",X"38",X"17",X"0F",
		X"17",X"01",X"02",X"38",X"17",X"3A",X"17",X"01",X"03",X"38",X"17",X"0F",X"17",X"38",X"17",X"0F",
		X"17",X"01",X"03",X"38",X"17",X"00",X"01",X"12",X"0F",X"17",X"3B",X"17",X"00",X"01",X"12",X"0F",
		X"17",X"3B",X"17",X"00",X"01",X"0D",X"0F",X"17",X"3B",X"17",X"01",X"04",X"0F",X"17",X"3B",X"17",
		X"00",X"01",X"03",X"38",X"17",X"0F",X"17",X"38",X"17",X"0F",X"17",X"01",X"07",X"38",X"17",X"3A",
		X"17",X"38",X"17",X"01",X"02",X"0F",X"17",X"01",X"03",X"38",X"17",X"0F",X"17",X"38",X"17",X"0F",
		X"17",X"01",X"05",X"38",X"17",X"00",X"01",X"0D",X"0F",X"17",X"3B",X"17",X"00",X"01",X"0D",X"0F",
		X"17",X"3B",X"17",X"00",X"01",X"02",X"0F",X"17",X"3B",X"17",X"01",X"0A",X"0F",X"17",X"3B",X"17",
		X"00",X"01",X"02",X"38",X"17",X"3A",X"17",X"38",X"17",X"01",X"03",X"0F",X"17",X"01",X"03",X"38",
		X"17",X"0F",X"17",X"01",X"04",X"38",X"17",X"0F",X"17",X"01",X"02",X"38",X"17",X"01",X"03",X"0F",
		X"17",X"01",X"07",X"38",X"17",X"00",X"01",X"02",X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",X"0F",
		X"17",X"3B",X"17",X"00",X"01",X"02",X"0F",X"17",X"3B",X"17",X"01",X"06",X"0F",X"17",X"3B",X"17",
		X"00",X"01",X"05",X"38",X"17",X"0F",X"17",X"01",X"03",X"38",X"17",X"3A",X"17",X"01",X"03",X"38",
		X"17",X"01",X"03",X"0F",X"17",X"01",X"03",X"38",X"17",X"0F",X"17",X"01",X"02",X"38",X"17",X"01",
		X"02",X"0F",X"17",X"01",X"04",X"38",X"17",X"00",X"01",X"09",X"0F",X"17",X"3B",X"17",X"00",X"01",
		X"09",X"0F",X"17",X"3B",X"17",X"00",X"01",X"09",X"0F",X"17",X"3B",X"17",X"00",X"FF",X"01",X"09",
		X"0F",X"17",X"3B",X"17",X"00",X"01",X"03",X"38",X"17",X"01",X"02",X"0F",X"17",X"01",X"02",X"38",
		X"17",X"0F",X"17",X"38",X"17",X"3A",X"17",X"38",X"17",X"0F",X"17",X"38",X"17",X"0F",X"17",X"01",
		X"06",X"38",X"17",X"01",X"02",X"38",X"17",X"0F",X"17",X"01",X"05",X"38",X"17",X"00",X"01",X"09",
		X"0F",X"17",X"3B",X"17",X"00",X"01",X"09",X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",X"0F",X"17",
		X"3B",X"17",X"01",X"06",X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",X"38",X"17",X"3A",X"17",X"38",
		X"17",X"0F",X"17",X"01",X"02",X"38",X"17",X"0F",X"17",X"01",X"03",X"38",X"17",X"0F",X"17",X"38",
		X"17",X"01",X"04",X"38",X"17",X"38",X"17",X"0F",X"17",X"01",X"02",X"38",X"17",X"0F",X"17",X"01",
		X"02",X"38",X"17",X"0F",X"17",X"01",X"03",X"38",X"17",X"00",X"01",X"02",X"0F",X"17",X"3B",X"17",
		X"00",X"01",X"02",X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",X"0F",X"17",X"01",X"02",X"3B",X"17",
		X"00",X"01",X"03",X"38",X"17",X"3A",X"17",X"38",X"17",X"0F",X"17",X"38",X"17",X"0F",X"17",X"38",
		X"17",X"01",X"03",X"0F",X"17",X"38",X"17",X"0F",X"17",X"01",X"02",X"38",X"17",X"0F",X"17",X"38",
		X"17",X"01",X"02",X"0F",X"17",X"01",X"02",X"38",X"17",X"01",X"03",X"0F",X"17",X"01",X"03",X"38",
		X"17",X"00",X"01",X"03",X"0F",X"17",X"3B",X"17",X"00",X"01",X"03",X"0F",X"17",X"3B",X"17",X"00",
		X"01",X"03",X"0F",X"17",X"3B",X"17",X"01",X"04",X"0F",X"17",X"3B",X"17",X"00",X"01",X"08",X"38",
		X"17",X"3A",X"17",X"01",X"02",X"38",X"17",X"0F",X"17",X"01",X"07",X"38",X"17",X"0F",X"17",X"01",
		X"03",X"38",X"17",X"0F",X"17",X"01",X"04",X"38",X"17",X"00",X"01",X"08",X"0F",X"17",X"3B",X"17",
		X"00",X"01",X"08",X"0F",X"17",X"3B",X"17",X"00",X"01",X"08",X"0F",X"17",X"3B",X"17",X"00",X"FF",
		X"01",X"02",X"0F",X"17",X"3B",X"17",X"01",X"17",X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",X"38",
		X"17",X"3A",X"17",X"38",X"17",X"01",X"02",X"0F",X"17",X"01",X"04",X"38",X"17",X"0F",X"17",X"38",
		X"17",X"0F",X"17",X"38",X"17",X"0F",X"17",X"38",X"17",X"01",X"02",X"0F",X"17",X"01",X"04",X"38",
		X"17",X"0F",X"17",X"38",X"17",X"0F",X"17",X"38",X"17",X"3A",X"17",X"38",X"17",X"00",X"01",X"02",
		X"0F",X"17",X"3B",X"17",X"01",X"17",X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",X"0F",X"17",X"3B",
		X"17",X"01",X"17",X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",X"0F",X"17",X"3B",X"17",X"01",X"04",
		X"0F",X"17",X"3B",X"17",X"01",X"0B",X"0F",X"17",X"3B",X"17",X"01",X"06",X"0F",X"17",X"3B",X"17",
		X"00",X"01",X"07",X"38",X"17",X"3A",X"17",X"38",X"17",X"0F",X"17",X"38",X"17",X"01",X"02",X"0F",
		X"17",X"01",X"02",X"38",X"17",X"01",X"02",X"0F",X"17",X"01",X"02",X"38",X"17",X"3A",X"17",X"01",
		X"08",X"38",X"17",X"00",X"01",X"07",X"0F",X"17",X"3B",X"17",X"01",X"0B",X"0F",X"17",X"3B",X"17",
		X"00",X"01",X"07",X"0F",X"17",X"3B",X"17",X"01",X"0B",X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",
		X"0F",X"17",X"3B",X"17",X"01",X"04",X"0F",X"17",X"3B",X"17",X"01",X"0B",X"0F",X"17",X"3B",X"17",
		X"01",X"06",X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",X"38",X"17",X"3A",X"17",X"38",X"17",X"01",
		X"02",X"0F",X"17",X"01",X"03",X"38",X"17",X"01",X"02",X"0F",X"17",X"01",X"02",X"38",X"17",X"0F",
		X"17",X"01",X"02",X"38",X"17",X"01",X"02",X"0F",X"17",X"01",X"03",X"38",X"17",X"01",X"03",X"0F",
		X"17",X"01",X"02",X"38",X"17",X"3A",X"17",X"38",X"17",X"00",X"01",X"02",X"0F",X"17",X"3B",X"17",
		X"01",X"17",X"0F",X"17",X"3B",X"17",X"00",X"01",X"02",X"0F",X"17",X"3B",X"17",X"01",X"17",X"0F",
		X"17",X"3B",X"17",X"00",X"01",X"02",X"0F",X"17",X"3B",X"17",X"01",X"0C",X"0F",X"17",X"3B",X"17",
		X"01",X"0A",X"0F",X"17",X"3B",X"17",X"00",X"01",X"04",X"38",X"17",X"0F",X"17",X"01",X"02",X"38",
		X"17",X"0F",X"17",X"38",X"17",X"0F",X"17",X"01",X"05",X"38",X"17",X"3A",X"17",X"38",X"17",X"0F",
		X"17",X"38",X"17",X"0F",X"17",X"01",X"02",X"38",X"17",X"0F",X"17",X"38",X"17",X"0F",X"17",X"01",
		X"03",X"38",X"17",X"00",X"01",X"0F",X"0F",X"17",X"3B",X"17",X"00",X"01",X"0F",X"0F",X"17",X"3B",
		X"17",X"00",X"01",X"0F",X"0F",X"17",X"3B",X"17",X"00",X"FF",X"01",X"0E",X"0F",X"17",X"3B",X"17",
		X"00",X"01",X"03",X"38",X"17",X"0F",X"17",X"38",X"17",X"0F",X"17",X"38",X"17",X"0F",X"17",X"01",
		X"02",X"38",X"17",X"0F",X"17",X"38",X"17",X"0F",X"17",X"38",X"17",X"3A",X"17",X"01",X"02",X"38",
		X"17",X"0F",X"17",X"38",X"17",X"0F",X"17",X"01",X"02",X"38",X"17",X"0F",X"17",X"38",X"17",X"0F",
		X"17",X"01",X"03",X"38",X"17",X"00",X"01",X"0E",X"0F",X"17",X"3B",X"17",X"00",X"01",X"0E",X"0F",
		X"17",X"3B",X"17",X"00",X"01",X"0A",X"0F",X"17",X"3B",X"17",X"01",X"03",X"0F",X"17",X"3B",X"17",
		X"01",X"03",X"0F",X"17",X"3B",X"17",X"00",X"01",X"06",X"38",X"17",X"01",X"02",X"0F",X"17",X"01",
		X"02",X"38",X"17",X"3A",X"17",X"38",X"17",X"0F",X"17",X"01",X"03",X"38",X"17",X"0F",X"17",X"38",
		X"17",X"3A",X"17",X"38",X"17",X"01",X"02",X"0F",X"17",X"01",X"06",X"38",X"17",X"00",X"01",X"0A",
		X"0F",X"17",X"3B",X"17",X"01",X"07",X"0F",X"17",X"3B",X"17",X"00",X"01",X"0A",X"0F",X"17",X"3B",
		X"17",X"01",X"07",X"0F",X"17",X"3B",X"17",X"00",X"01",X"0A",X"0F",X"17",X"3B",X"17",X"01",X"07",
		X"0F",X"17",X"3B",X"17",X"01",X"03",X"0F",X"17",X"3B",X"17",X"00",X"01",X"0D",X"38",X"17",X"01",
		X"03",X"0F",X"17",X"01",X"06",X"38",X"17",X"3A",X"17",X"38",X"17",X"0F",X"17",X"01",X"03",X"38",
		X"17",X"00",X"01",X"16",X"0F",X"17",X"3B",X"17",X"00",X"01",X"16",X"0F",X"17",X"3B",X"17",X"00",
		X"01",X"03",X"0F",X"17",X"3B",X"17",X"01",X"12",X"0F",X"17",X"3B",X"17",X"01",X"02",X"0F",X"17",
		X"3B",X"17",X"00",X"01",X"03",X"38",X"17",X"3A",X"17",X"38",X"17",X"0F",X"17",X"01",X"02",X"38",
		X"17",X"01",X"03",X"0F",X"17",X"01",X"06",X"38",X"17",X"0F",X"17",X"38",X"17",X"01",X"02",X"0F",
		X"17",X"01",X"04",X"38",X"17",X"3A",X"17",X"01",X"02",X"38",X"17",X"00",X"01",X"03",X"0F",X"17",
		X"3B",X"17",X"01",X"15",X"0F",X"17",X"3B",X"17",X"00",X"01",X"03",X"0F",X"17",X"3B",X"17",X"01",
		X"15",X"0F",X"17",X"3B",X"17",X"00",X"01",X"03",X"0F",X"17",X"3B",X"17",X"01",X"15",X"0F",X"17",
		X"3B",X"17",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"70",X"12",X"74",X"0F",X"78",X"15",X"7C",X"15",X"80",
		X"15",X"84",X"0F",X"88",X"03",X"8C",X"17",X"90",X"15",X"94",X"16",X"98",X"0F",X"9C",X"07",X"A0",
		X"17",X"A4",X"0F",X"A8",X"03",X"AC",X"15",X"B0",X"18",X"B4",X"17",X"B8",X"16",X"BC",X"16",X"95",
		X"76",X"95",X"26",X"95",X"36",X"95",X"86",X"95",X"56",X"95",X"96",X"95",X"46",X"95",X"B6",X"95",
		X"A6",X"95",X"66",X"95",X"C6",X"95",X"D6",X"95",X"F6",X"95",X"E6",X"95",X"B6",X"95",X"66",X"95",
		X"06",X"96",X"C6",X"95",X"16",X"96",X"34",X"18",X"07",X"A8",X"34",X"18",X"87",X"A8",X"34",X"18",
		X"07",X"88",X"34",X"18",X"8F",X"48",X"34",X"18",X"8F",X"A8",X"34",X"18",X"8F",X"88",X"34",X"18",
		X"27",X"68",X"34",X"18",X"08",X"48",X"34",X"18",X"AF",X"A8",X"34",X"18",X"3F",X"88",X"34",X"18",
		X"87",X"68",X"34",X"18",X"67",X"28",X"34",X"18",X"97",X"88",X"34",X"18",X"B7",X"68",X"34",X"18",
		X"6F",X"48",X"34",X"18",X"97",X"28",X"34",X"18",X"B7",X"A8",X"34",X"18",X"3F",X"88",X"34",X"18",
		X"97",X"68",X"34",X"18",X"2F",X"48",X"34",X"18",X"9F",X"88",X"34",X"18",X"1F",X"68",X"34",X"18",
		X"9F",X"48",X"34",X"18",X"BF",X"28",X"34",X"18",X"97",X"A8",X"34",X"18",X"07",X"88",X"34",X"18",
		X"C7",X"68",X"34",X"18",X"3F",X"48",X"34",X"18",X"C7",X"A8",X"34",X"18",X"3F",X"88",X"34",X"18",
		X"4F",X"68",X"34",X"18",X"87",X"48",X"34",X"18",X"5F",X"88",X"34",X"18",X"27",X"68",X"34",X"18",
		X"C7",X"48",X"34",X"18",X"27",X"48",X"34",X"18",X"57",X"A8",X"34",X"18",X"8F",X"88",X"34",X"18",
		X"77",X"68",X"34",X"18",X"4F",X"48",X"34",X"18",X"AF",X"88",X"34",X"18",X"27",X"88",X"34",X"18",
		X"B7",X"48",X"34",X"18",X"27",X"48",X"34",X"18",X"AF",X"88",X"34",X"18",X"1F",X"68",X"34",X"18",
		X"AF",X"48",X"34",X"18",X"CF",X"28",X"34",X"18",X"6F",X"A8",X"34",X"18",X"27",X"68",X"34",X"18",
		X"27",X"48",X"34",X"18",X"3F",X"28",X"34",X"18",X"9F",X"A8",X"34",X"18",X"47",X"88",X"34",X"18",
		X"7F",X"68",X"34",X"18",X"2F",X"48",X"34",X"18",X"27",X"88",X"34",X"18",X"27",X"48",X"34",X"18",
		X"5F",X"48",X"34",X"18",X"27",X"28",X"34",X"18",X"9F",X"A8",X"34",X"18",X"1F",X"88",X"34",X"18",
		X"B7",X"88",X"34",X"18",X"67",X"48",X"34",X"18",X"9F",X"A8",X"34",X"18",X"37",X"68",X"34",X"18",
		X"97",X"68",X"34",X"18",X"77",X"48",X"4E",X"96",X"11",X"98",X"8B",X"96",X"D7",X"96",X"58",X"98",
		X"74",X"97",X"A4",X"98",X"23",X"97",X"46",X"99",X"F5",X"98",X"C0",X"97",X"97",X"99",X"E8",X"99",
		X"8A",X"9A",X"39",X"9A",X"7D",X"9B",X"CE",X"9B",X"DB",X"9A",X"1F",X"9C",X"2C",X"9B",X"01",X"25",
		X"41",X"15",X"70",X"01",X"35",X"41",X"15",X"70",X"01",X"B9",X"41",X"15",X"70",X"01",X"28",X"42",
		X"15",X"70",X"01",X"39",X"42",X"15",X"70",X"01",X"A1",X"42",X"15",X"70",X"01",X"B9",X"42",X"15",
		X"70",X"01",X"29",X"43",X"15",X"70",X"00",X"58",X"41",X"0F",X"30",X"00",X"CE",X"41",X"0F",X"30",
		X"00",X"4E",X"42",X"0F",X"30",X"00",X"57",X"43",X"0F",X"30",X"FF",X"01",X"20",X"41",X"0F",X"78",
		X"01",X"2A",X"41",X"0F",X"78",X"01",X"2F",X"41",X"0F",X"78",X"01",X"A0",X"41",X"0F",X"78",X"01",
		X"2D",X"42",X"0F",X"78",X"01",X"A8",X"42",X"0F",X"78",X"01",X"B3",X"42",X"0F",X"78",X"01",X"21",
		X"43",X"0F",X"78",X"00",X"48",X"41",X"0F",X"30",X"00",X"55",X"41",X"0F",X"30",X"00",X"58",X"41",
		X"0F",X"30",X"00",X"4A",X"42",X"0F",X"30",X"00",X"4E",X"43",X"0F",X"30",X"00",X"51",X"43",X"0F",
		X"30",X"00",X"54",X"43",X"0F",X"30",X"FF",X"01",X"25",X"41",X"15",X"7C",X"01",X"31",X"41",X"15",
		X"7C",X"01",X"A3",X"41",X"15",X"7C",X"01",X"AD",X"41",X"15",X"7C",X"01",X"B2",X"41",X"15",X"7C",
		X"01",X"2A",X"42",X"15",X"7C",X"01",X"AA",X"42",X"15",X"7C",X"01",X"B0",X"42",X"15",X"7C",X"00",
		X"44",X"41",X"0F",X"30",X"00",X"44",X"42",X"0F",X"30",X"00",X"C5",X"42",X"0F",X"30",X"00",X"D6",
		X"42",X"0F",X"30",X"00",X"50",X"43",X"0F",X"30",X"00",X"55",X"43",X"0F",X"30",X"00",X"58",X"43",
		X"0F",X"30",X"FF",X"01",X"21",X"41",X"03",X"8C",X"01",X"35",X"41",X"03",X"8C",X"01",X"A4",X"41",
		X"03",X"8C",X"01",X"AF",X"41",X"03",X"8C",X"01",X"34",X"42",X"03",X"8C",X"01",X"A1",X"42",X"03",
		X"8C",X"01",X"B9",X"42",X"03",X"8C",X"01",X"28",X"43",X"03",X"8C",X"00",X"C7",X"41",X"0F",X"30",
		X"00",X"44",X"42",X"0F",X"30",X"00",X"49",X"42",X"0F",X"30",X"00",X"4F",X"42",X"0F",X"30",X"00",
		X"4B",X"43",X"0F",X"30",X"00",X"50",X"43",X"0F",X"30",X"00",X"56",X"43",X"0F",X"30",X"00",X"59",
		X"43",X"0F",X"30",X"FF",X"01",X"2A",X"41",X"15",X"84",X"01",X"34",X"41",X"15",X"84",X"01",X"A1",
		X"41",X"15",X"84",X"01",X"B6",X"41",X"15",X"84",X"01",X"29",X"42",X"15",X"84",X"01",X"AB",X"42",
		X"15",X"84",X"01",X"B8",X"42",X"15",X"84",X"01",X"26",X"43",X"15",X"84",X"00",X"C6",X"41",X"0F",
		X"30",X"00",X"58",X"42",X"0F",X"30",X"00",X"4C",X"43",X"0F",X"30",X"00",X"4F",X"43",X"0F",X"30",
		X"00",X"50",X"43",X"0F",X"30",X"00",X"53",X"43",X"0F",X"30",X"00",X"56",X"43",X"0F",X"30",X"FF",
		X"01",X"28",X"41",X"16",X"98",X"01",X"31",X"41",X"16",X"98",X"01",X"B1",X"41",X"16",X"98",X"01",
		X"2A",X"42",X"16",X"98",X"01",X"2F",X"42",X"16",X"98",X"01",X"A5",X"42",X"16",X"98",X"01",X"B9",
		X"42",X"16",X"98",X"01",X"21",X"43",X"16",X"98",X"00",X"C4",X"42",X"0F",X"30",X"00",X"C7",X"42",
		X"0F",X"30",X"00",X"D3",X"42",X"0F",X"30",X"00",X"D6",X"42",X"0F",X"30",X"00",X"44",X"43",X"0F",
		X"30",X"00",X"47",X"43",X"0F",X"30",X"00",X"4B",X"43",X"0F",X"30",X"00",X"4F",X"43",X"0F",X"30",
		X"FF",X"01",X"21",X"41",X"12",X"74",X"01",X"A3",X"41",X"12",X"74",X"01",X"AB",X"41",X"12",X"74",
		X"01",X"B9",X"41",X"12",X"74",X"01",X"28",X"42",X"12",X"74",X"01",X"A1",X"42",X"12",X"74",X"01",
		X"B9",X"42",X"12",X"74",X"01",X"29",X"43",X"12",X"74",X"00",X"CE",X"41",X"0F",X"30",X"00",X"D3",
		X"41",X"0F",X"30",X"00",X"CD",X"42",X"0F",X"30",X"00",X"D2",X"42",X"0F",X"30",X"00",X"4C",X"43",
		X"0F",X"30",X"00",X"55",X"43",X"0F",X"30",X"FF",X"01",X"2A",X"41",X"15",X"80",X"01",X"2F",X"41",
		X"15",X"80",X"01",X"33",X"41",X"15",X"80",X"01",X"B1",X"41",X"15",X"80",X"01",X"2D",X"42",X"15",
		X"80",X"01",X"39",X"42",X"15",X"80",X"01",X"A4",X"42",X"15",X"80",X"01",X"2F",X"43",X"15",X"80",
		X"00",X"45",X"41",X"0F",X"30",X"00",X"48",X"41",X"0F",X"30",X"00",X"C6",X"41",X"0F",X"30",X"00",
		X"52",X"42",X"0F",X"30",X"00",X"D4",X"42",X"0F",X"30",X"00",X"4C",X"43",X"0F",X"30",X"00",X"53",
		X"43",X"0F",X"30",X"FF",X"01",X"21",X"41",X"0F",X"88",X"01",X"33",X"41",X"0F",X"88",X"01",X"A5",
		X"41",X"0F",X"88",X"01",X"B5",X"41",X"0F",X"88",X"01",X"35",X"42",X"0F",X"88",X"01",X"AB",X"42",
		X"0F",X"88",X"01",X"B0",X"42",X"0F",X"88",X"01",X"24",X"43",X"0F",X"88",X"00",X"45",X"41",X"0F",
		X"30",X"00",X"C4",X"42",X"0F",X"30",X"00",X"C7",X"42",X"0F",X"30",X"00",X"D6",X"42",X"0F",X"30",
		X"00",X"47",X"43",X"0F",X"30",X"00",X"4D",X"43",X"0F",X"30",X"00",X"50",X"43",X"0F",X"30",X"00",
		X"56",X"43",X"0F",X"30",X"FF",X"01",X"20",X"41",X"15",X"94",X"01",X"32",X"41",X"15",X"94",X"01",
		X"A1",X"41",X"15",X"94",X"01",X"AA",X"41",X"15",X"94",X"01",X"28",X"42",X"15",X"94",X"01",X"35",
		X"42",X"15",X"94",X"01",X"A0",X"42",X"15",X"94",X"01",X"B5",X"42",X"15",X"94",X"00",X"46",X"41",
		X"0F",X"30",X"00",X"49",X"41",X"0F",X"30",X"00",X"50",X"41",X"0F",X"30",X"00",X"55",X"41",X"0F",
		X"30",X"00",X"D8",X"41",X"0F",X"30",X"00",X"44",X"42",X"0F",X"30",X"00",X"4B",X"42",X"0F",X"30",
		X"00",X"C8",X"42",X"0F",X"30",X"FF",X"01",X"21",X"41",X"17",X"90",X"01",X"32",X"41",X"17",X"90",
		X"01",X"26",X"42",X"17",X"90",X"01",X"36",X"42",X"17",X"90",X"01",X"A0",X"42",X"17",X"90",X"01",
		X"B0",X"42",X"17",X"90",X"01",X"21",X"43",X"17",X"90",X"01",X"31",X"43",X"17",X"90",X"00",X"55",
		X"41",X"0F",X"30",X"00",X"58",X"41",X"0F",X"30",X"00",X"55",X"42",X"0F",X"30",X"00",X"44",X"43",
		X"0F",X"30",X"00",X"4A",X"43",X"0F",X"30",X"00",X"4D",X"43",X"0F",X"30",X"00",X"50",X"43",X"0F",
		X"30",X"00",X"53",X"43",X"0F",X"30",X"FF",X"01",X"2B",X"41",X"0F",X"9C",X"01",X"39",X"41",X"0F",
		X"9C",X"01",X"A5",X"41",X"0F",X"9C",X"01",X"AF",X"41",X"0F",X"9C",X"01",X"20",X"42",X"0F",X"9C",
		X"01",X"36",X"42",X"0F",X"9C",X"01",X"A5",X"42",X"0F",X"9C",X"01",X"2B",X"43",X"0F",X"9C",X"00",
		X"54",X"41",X"0F",X"30",X"00",X"57",X"41",X"0F",X"30",X"00",X"44",X"43",X"0F",X"30",X"00",X"47",
		X"43",X"0F",X"30",X"00",X"4A",X"43",X"0F",X"30",X"00",X"4D",X"43",X"0F",X"30",X"00",X"50",X"43",
		X"0F",X"30",X"00",X"53",X"43",X"0F",X"30",X"FF",X"01",X"24",X"41",X"07",X"A0",X"01",X"33",X"41",
		X"07",X"A0",X"01",X"39",X"41",X"07",X"A0",X"01",X"A8",X"41",X"07",X"A0",X"01",X"B9",X"41",X"07",
		X"A0",X"01",X"20",X"42",X"07",X"A0",X"01",X"AE",X"42",X"07",X"A0",X"01",X"24",X"43",X"07",X"A0",
		X"00",X"55",X"41",X"0F",X"30",X"00",X"CA",X"41",X"0F",X"30",X"00",X"43",X"42",X"0F",X"30",X"00",
		X"C7",X"42",X"0F",X"30",X"00",X"4C",X"43",X"0F",X"30",X"00",X"4E",X"43",X"0F",X"30",X"00",X"50",
		X"43",X"0F",X"30",X"00",X"52",X"43",X"0F",X"30",X"FF",X"01",X"25",X"41",X"0F",X"A8",X"01",X"39",
		X"41",X"0F",X"A8",X"01",X"A0",X"41",X"0F",X"A8",X"01",X"B9",X"41",X"0F",X"A8",X"01",X"38",X"42",
		X"0F",X"A8",X"01",X"AB",X"42",X"0F",X"A8",X"01",X"B8",X"42",X"0F",X"A8",X"01",X"22",X"43",X"0F",
		X"A8",X"00",X"C7",X"41",X"0F",X"30",X"00",X"D8",X"41",X"0F",X"30",X"00",X"49",X"42",X"0F",X"30",
		X"00",X"D2",X"42",X"0F",X"30",X"00",X"4C",X"43",X"0F",X"30",X"00",X"4F",X"43",X"0F",X"30",X"00",
		X"53",X"43",X"0F",X"30",X"00",X"56",X"43",X"0F",X"30",X"FF",X"01",X"39",X"41",X"17",X"A4",X"01",
		X"B6",X"41",X"17",X"A4",X"01",X"2E",X"42",X"17",X"A4",X"01",X"39",X"42",X"17",X"A4",X"01",X"A0",
		X"42",X"17",X"A4",X"01",X"B0",X"42",X"17",X"A4",X"01",X"B9",X"42",X"17",X"A4",X"01",X"21",X"43",
		X"17",X"A4",X"00",X"4F",X"41",X"0F",X"30",X"00",X"50",X"41",X"0F",X"30",X"00",X"55",X"41",X"0F",
		X"30",X"00",X"CE",X"41",X"0F",X"30",X"00",X"44",X"43",X"0F",X"30",X"00",X"4C",X"43",X"0F",X"30",
		X"00",X"4F",X"43",X"0F",X"30",X"00",X"51",X"43",X"0F",X"30",X"FF",X"01",X"28",X"41",X"18",X"B4",
		X"01",X"32",X"41",X"18",X"B4",X"01",X"AD",X"41",X"18",X"B4",X"01",X"2B",X"42",X"18",X"B4",X"01",
		X"2E",X"42",X"18",X"B4",X"01",X"A5",X"42",X"18",X"B4",X"01",X"B4",X"42",X"18",X"B4",X"01",X"22",
		X"43",X"18",X"B4",X"00",X"D6",X"41",X"0F",X"30",X"00",X"46",X"43",X"0F",X"30",X"00",X"49",X"43",
		X"0F",X"30",X"00",X"51",X"43",X"0F",X"30",X"00",X"52",X"43",X"0F",X"30",X"00",X"55",X"43",X"0F",
		X"30",X"00",X"58",X"43",X"0F",X"30",X"00",X"59",X"43",X"0F",X"30",X"FF",X"01",X"21",X"41",X"16",
		X"BC",X"01",X"39",X"41",X"16",X"BC",X"01",X"A4",X"41",X"16",X"BC",X"01",X"B8",X"41",X"16",X"BC",
		X"01",X"21",X"42",X"16",X"BC",X"01",X"39",X"42",X"16",X"BC",X"01",X"AD",X"42",X"16",X"BC",X"01",
		X"2D",X"43",X"16",X"BC",X"00",X"C8",X"41",X"0F",X"30",X"00",X"D7",X"41",X"0F",X"30",X"00",X"CC",
		X"42",X"0F",X"30",X"00",X"4B",X"43",X"0F",X"30",X"00",X"4C",X"43",X"0F",X"30",X"00",X"4F",X"43",
		X"0F",X"30",X"00",X"50",X"43",X"0F",X"30",X"00",X"51",X"43",X"0F",X"30",X"FF",X"01",X"21",X"41",
		X"03",X"AC",X"01",X"32",X"41",X"03",X"AC",X"01",X"26",X"42",X"03",X"AC",X"01",X"36",X"42",X"03",
		X"AC",X"01",X"A0",X"42",X"03",X"AC",X"01",X"B0",X"42",X"03",X"AC",X"01",X"21",X"43",X"03",X"AC",
		X"01",X"31",X"43",X"03",X"AC",X"00",X"55",X"41",X"0F",X"30",X"00",X"58",X"41",X"0F",X"30",X"00",
		X"55",X"42",X"0F",X"30",X"00",X"44",X"43",X"0F",X"30",X"00",X"4A",X"43",X"0F",X"30",X"00",X"4D",
		X"43",X"0F",X"30",X"00",X"50",X"43",X"0F",X"30",X"00",X"53",X"43",X"0F",X"30",X"FF",X"01",X"28",
		X"41",X"15",X"B0",X"01",X"31",X"41",X"15",X"B0",X"01",X"B1",X"41",X"15",X"B0",X"01",X"2A",X"42",
		X"15",X"B0",X"01",X"2F",X"42",X"15",X"B0",X"01",X"A5",X"42",X"15",X"B0",X"01",X"B9",X"42",X"15",
		X"B0",X"01",X"21",X"43",X"15",X"B0",X"00",X"C4",X"42",X"0F",X"30",X"00",X"C7",X"42",X"0F",X"30",
		X"00",X"D3",X"42",X"0F",X"30",X"00",X"D6",X"42",X"0F",X"30",X"00",X"44",X"43",X"0F",X"30",X"00",
		X"47",X"43",X"0F",X"30",X"00",X"4B",X"43",X"0F",X"30",X"00",X"4F",X"43",X"0F",X"30",X"FF",X"01",
		X"2B",X"41",X"17",X"B8",X"01",X"39",X"41",X"17",X"B8",X"01",X"A5",X"41",X"17",X"B8",X"01",X"AF",
		X"41",X"17",X"B8",X"01",X"20",X"42",X"17",X"B8",X"01",X"36",X"42",X"17",X"B8",X"01",X"A5",X"42",
		X"17",X"B8",X"01",X"2B",X"43",X"17",X"B8",X"00",X"54",X"41",X"0F",X"30",X"00",X"57",X"41",X"0F",
		X"30",X"00",X"44",X"43",X"0F",X"30",X"00",X"47",X"43",X"0F",X"30",X"00",X"4A",X"43",X"0F",X"30",
		X"00",X"4D",X"43",X"0F",X"30",X"00",X"50",X"43",X"0F",X"30",X"00",X"53",X"43",X"0F",X"30",X"FF",
		X"2C",X"9D",X"E2",X"9C",X"98",X"9C",X"BD",X"9C",X"07",X"9D",X"76",X"9D",X"51",X"9D",X"9B",X"9D",
		X"C0",X"9D",X"E5",X"9D",X"2F",X"9E",X"0A",X"9E",X"54",X"9E",X"9E",X"9E",X"79",X"9E",X"C0",X"9D",
		X"2F",X"9E",X"C3",X"9E",X"0A",X"9E",X"E8",X"9E",X"08",X"00",X"21",X"43",X"FF",X"40",X"00",X"A8",
		X"42",X"98",X"00",X"B3",X"42",X"FF",X"68",X"00",X"2D",X"42",X"FF",X"00",X"00",X"A0",X"41",X"FF",
		X"00",X"00",X"20",X"41",X"50",X"00",X"2A",X"41",X"78",X"00",X"2F",X"41",X"FF",X"FF",X"50",X"00",
		X"AA",X"42",X"80",X"00",X"B0",X"42",X"FF",X"50",X"00",X"2A",X"42",X"FF",X"18",X"00",X"A3",X"41",
		X"68",X"00",X"AD",X"41",X"90",X"00",X"B2",X"41",X"FF",X"28",X"00",X"25",X"41",X"88",X"00",X"31",
		X"41",X"FF",X"48",X"00",X"29",X"43",X"FF",X"08",X"00",X"A1",X"42",X"C8",X"00",X"B9",X"42",X"FF",
		X"40",X"00",X"28",X"42",X"FF",X"18",X"00",X"A3",X"41",X"58",X"00",X"AB",X"41",X"C8",X"00",X"B9",
		X"41",X"FF",X"08",X"00",X"21",X"41",X"FF",X"78",X"00",X"2F",X"43",X"FF",X"20",X"00",X"A4",X"42",
		X"FF",X"68",X"00",X"2D",X"42",X"C8",X"00",X"39",X"42",X"FF",X"88",X"00",X"B1",X"41",X"FF",X"50",
		X"00",X"2A",X"41",X"78",X"00",X"2F",X"41",X"98",X"00",X"33",X"41",X"FF",X"48",X"00",X"29",X"43",
		X"FF",X"08",X"00",X"A1",X"42",X"C8",X"00",X"B9",X"42",X"FF",X"40",X"00",X"28",X"42",X"C8",X"00",
		X"39",X"42",X"FF",X"C8",X"00",X"B9",X"41",X"FF",X"28",X"00",X"25",X"41",X"A8",X"00",X"35",X"41",
		X"FF",X"20",X"00",X"24",X"43",X"FF",X"58",X"00",X"AB",X"42",X"80",X"00",X"B0",X"42",X"FF",X"A8",
		X"00",X"35",X"42",X"FF",X"28",X"00",X"A5",X"41",X"A8",X"00",X"B5",X"41",X"FF",X"08",X"00",X"21",
		X"41",X"98",X"00",X"33",X"41",X"FF",X"30",X"00",X"26",X"43",X"FF",X"58",X"00",X"AB",X"42",X"C0",
		X"00",X"B8",X"42",X"FF",X"48",X"00",X"29",X"42",X"FF",X"08",X"00",X"A1",X"41",X"B0",X"00",X"B6",
		X"41",X"FF",X"50",X"00",X"2A",X"41",X"A0",X"00",X"34",X"41",X"FF",X"40",X"00",X"28",X"43",X"FF",
		X"08",X"00",X"A1",X"42",X"C8",X"00",X"B9",X"42",X"FF",X"A0",X"00",X"34",X"42",X"FF",X"20",X"00",
		X"A4",X"41",X"78",X"00",X"AF",X"41",X"FF",X"08",X"00",X"21",X"41",X"A8",X"00",X"35",X"41",X"FF",
		X"08",X"00",X"21",X"43",X"88",X"00",X"31",X"43",X"FF",X"00",X"00",X"A0",X"42",X"80",X"00",X"B0",
		X"42",X"FF",X"30",X"00",X"26",X"42",X"B0",X"00",X"36",X"42",X"FF",X"FF",X"08",X"00",X"21",X"41",
		X"90",X"00",X"32",X"41",X"FF",X"FF",X"00",X"00",X"A0",X"42",X"A8",X"00",X"B5",X"42",X"FF",X"40",
		X"00",X"28",X"42",X"A8",X"00",X"35",X"42",X"FF",X"08",X"00",X"A1",X"41",X"50",X"00",X"AA",X"41",
		X"FF",X"00",X"00",X"20",X"41",X"90",X"00",X"32",X"41",X"FF",X"58",X"00",X"2B",X"43",X"FF",X"28",
		X"00",X"A5",X"42",X"FF",X"00",X"00",X"20",X"42",X"B0",X"00",X"36",X"42",X"FF",X"28",X"00",X"A5",
		X"41",X"78",X"00",X"AF",X"41",X"FF",X"58",X"00",X"2B",X"41",X"C8",X"00",X"39",X"41",X"FF",X"08",
		X"00",X"21",X"43",X"FF",X"28",X"00",X"A5",X"42",X"C8",X"00",X"B9",X"42",X"FF",X"50",X"00",X"2A",
		X"42",X"78",X"00",X"2F",X"42",X"FF",X"88",X"00",X"B1",X"41",X"FF",X"40",X"00",X"28",X"41",X"88",
		X"00",X"31",X"41",X"FF",X"20",X"00",X"24",X"43",X"FF",X"70",X"00",X"AE",X"42",X"FF",X"00",X"00",
		X"20",X"42",X"FF",X"40",X"00",X"A8",X"41",X"C8",X"00",X"B9",X"41",X"FF",X"20",X"00",X"24",X"41",
		X"98",X"00",X"33",X"41",X"C8",X"00",X"39",X"41",X"FF",X"10",X"00",X"22",X"43",X"FF",X"58",X"00",
		X"AB",X"42",X"C0",X"00",X"B8",X"42",X"FF",X"C0",X"00",X"38",X"42",X"FF",X"00",X"00",X"A0",X"41",
		X"C8",X"00",X"B9",X"41",X"FF",X"28",X"00",X"25",X"41",X"C8",X"00",X"39",X"41",X"FF",X"08",X"00",
		X"21",X"43",X"FF",X"00",X"00",X"A0",X"42",X"80",X"00",X"B0",X"42",X"C8",X"00",X"B9",X"42",X"FF",
		X"70",X"00",X"2E",X"42",X"C8",X"00",X"39",X"42",X"FF",X"B0",X"00",X"B6",X"41",X"FF",X"C8",X"00",
		X"39",X"41",X"FF",X"10",X"00",X"22",X"43",X"FF",X"28",X"00",X"A5",X"42",X"A0",X"00",X"B4",X"42",
		X"FF",X"58",X"00",X"2B",X"42",X"70",X"00",X"2E",X"42",X"FF",X"68",X"00",X"AD",X"41",X"FF",X"40",
		X"00",X"28",X"41",X"90",X"00",X"32",X"41",X"FF",X"68",X"00",X"2D",X"43",X"FF",X"68",X"00",X"AD",
		X"42",X"FF",X"08",X"00",X"21",X"42",X"C8",X"00",X"39",X"42",X"FF",X"20",X"00",X"A4",X"41",X"C0",
		X"00",X"B8",X"41",X"FF",X"08",X"00",X"21",X"41",X"C8",X"00",X"39",X"41",X"FF",X"89",X"9F",X"5F",
		X"9F",X"35",X"9F",X"4A",X"9F",X"74",X"9F",X"B3",X"9F",X"9E",X"9F",X"C8",X"9F",X"DD",X"9F",X"F2",
		X"9F",X"1C",X"A0",X"07",X"A0",X"31",X"A0",X"5B",X"A0",X"46",X"A0",X"DD",X"9F",X"1C",X"A0",X"70",
		X"A0",X"07",X"A0",X"85",X"A0",X"FF",X"07",X"33",X"08",X"4C",X"FF",X"27",X"43",X"06",X"4C",X"FF",
		X"8F",X"02",X"04",X"4C",X"FF",X"8F",X"53",X"02",X"4C",X"FF",X"67",X"02",X"08",X"4C",X"FF",X"FF",
		X"87",X"02",X"06",X"4C",X"FF",X"40",X"63",X"04",X"4C",X"FF",X"AF",X"02",X"02",X"4C",X"FF",X"FF",
		X"3F",X"02",X"08",X"4C",X"FF",X"C7",X"53",X"06",X"4C",X"FF",X"08",X"63",X"04",X"4C",X"FF",X"97",
		X"02",X"02",X"4C",X"FF",X"FF",X"87",X"02",X"08",X"4C",X"FF",X"4F",X"33",X"06",X"4C",X"FF",X"3F",
		X"02",X"04",X"4C",X"FF",X"C7",X"43",X"02",X"4C",X"FF",X"FF",X"8F",X"02",X"08",X"4C",X"FF",X"FF",
		X"07",X"53",X"06",X"4C",X"FF",X"87",X"02",X"04",X"4C",X"07",X"63",X"02",X"4C",X"FF",X"FF",X"27",
		X"02",X"08",X"4C",X"CF",X"33",X"06",X"4C",X"FF",X"27",X"43",X"04",X"4C",X"FF",X"5F",X"02",X"02",
		X"4C",X"FF",X"FF",X"FF",X"2F",X"43",X"08",X"4C",X"FF",X"97",X"02",X"06",X"4C",X"FF",X"3F",X"53",
		X"04",X"4C",X"FF",X"B7",X"02",X"02",X"4C",X"FF",X"97",X"02",X"08",X"4C",X"FF",X"6F",X"02",X"06",
		X"4C",X"FF",X"B7",X"33",X"04",X"4C",X"FF",X"97",X"43",X"02",X"4C",X"FF",X"FF",X"FF",X"27",X"43",
		X"08",X"4C",X"B7",X"02",X"06",X"4C",X"FF",X"FF",X"27",X"33",X"04",X"4C",X"AF",X"63",X"02",X"4C",
		X"FF",X"FF",X"FF",X"4F",X"02",X"08",X"4C",X"FF",X"77",X"63",X"06",X"4C",X"FF",X"8F",X"33",X"04",
		X"4C",X"FF",X"57",X"02",X"02",X"4C",X"FF",X"CF",X"02",X"08",X"4C",X"FF",X"AF",X"02",X"06",X"4C",
		X"FF",X"1F",X"02",X"04",X"4C",X"FF",X"AF",X"43",X"02",X"4C",X"FF",X"FF",X"BF",X"02",X"08",X"4C",
		X"FF",X"9F",X"33",X"06",X"4C",X"FF",X"1F",X"43",X"04",X"4C",X"FF",X"9F",X"02",X"02",X"4C",X"FF",
		X"FF",X"3F",X"02",X"08",X"4C",X"FF",X"27",X"02",X"06",X"4C",X"FF",X"27",X"02",X"04",X"4C",X"FF",
		X"FF",X"6F",X"63",X"02",X"4C",X"FF",X"FF",X"2F",X"02",X"08",X"4C",X"FF",X"7F",X"02",X"06",X"4C",
		X"FF",X"47",X"53",X"04",X"4C",X"FF",X"9F",X"02",X"02",X"4C",X"FF",X"27",X"63",X"08",X"4C",X"FF",
		X"5F",X"02",X"06",X"4C",X"27",X"53",X"04",X"4C",X"FF",X"FF",X"27",X"02",X"02",X"4C",X"FF",X"FF",
		X"FF",X"67",X"43",X"08",X"4C",X"FF",X"FF",X"B7",X"63",X"06",X"4C",X"1F",X"63",X"04",X"4C",X"FF",
		X"9F",X"63",X"02",X"4C",X"FF",X"FF",X"77",X"43",X"08",X"4C",X"FF",X"97",X"43",X"06",X"4C",X"37",
		X"43",X"04",X"4C",X"FF",X"FF",X"9F",X"63",X"02",X"4C",X"FF",X"10",X"00",X"20",X"00",X"30",X"00",
		X"50",X"00",X"00",X"01",X"00",X"02",X"00",X"03",X"00",X"05",X"00",X"10",X"00",X"20",X"00",X"30",
		X"00",X"50",X"56",X"A1",X"18",X"A1",X"DA",X"A0",X"F9",X"A0",X"37",X"A1",X"8A",X"A1",X"6B",X"A1",
		X"A9",X"A1",X"BE",X"A1",X"DD",X"A1",X"11",X"A2",X"F2",X"A1",X"30",X"A2",X"6E",X"A2",X"4F",X"A2",
		X"BE",X"A1",X"11",X"A2",X"83",X"A2",X"F2",X"A1",X"F2",X"A1",X"F8",X"17",X"28",X"40",X"01",X"01",
		X"02",X"0A",X"4C",X"02",X"F8",X"18",X"48",X"C8",X"01",X"02",X"03",X"0C",X"4C",X"03",X"F8",X"17",
		X"68",X"C8",X"01",X"01",X"02",X"0E",X"4C",X"02",X"FF",X"F8",X"17",X"28",X"50",X"01",X"01",X"02",
		X"0A",X"4C",X"02",X"F8",X"17",X"48",X"C8",X"01",X"01",X"02",X"0C",X"4C",X"02",X"F8",X"17",X"68",
		X"C8",X"01",X"01",X"02",X"0E",X"4C",X"02",X"FF",X"F8",X"17",X"28",X"08",X"00",X"01",X"02",X"0A",
		X"4C",X"02",X"F8",X"18",X"68",X"08",X"00",X"02",X"03",X"0C",X"4C",X"03",X"F8",X"17",X"A8",X"C8",
		X"01",X"01",X"03",X"0E",X"4C",X"03",X"FF",X"F8",X"17",X"28",X"08",X"00",X"01",X"02",X"0A",X"4C",
		X"02",X"F8",X"18",X"48",X"C8",X"01",X"02",X"03",X"0C",X"4C",X"03",X"F8",X"18",X"88",X"C8",X"00",
		X"02",X"03",X"0E",X"4C",X"03",X"FF",X"F8",X"17",X"68",X"04",X"00",X"01",X"02",X"0A",X"4C",X"02",
		X"F8",X"17",X"A8",X"00",X"01",X"01",X"02",X"0C",X"4C",X"02",X"FF",X"F8",X"17",X"28",X"40",X"01",
		X"01",X"02",X"0A",X"4C",X"02",X"F8",X"18",X"68",X"C8",X"01",X"02",X"03",X"0C",X"4C",X"03",X"F8",
		X"17",X"A8",X"B0",X"01",X"01",X"02",X"0E",X"4C",X"02",X"FF",X"F8",X"18",X"28",X"C0",X"01",X"02",
		X"03",X"0A",X"4C",X"03",X"F8",X"17",X"A8",X"20",X"01",X"01",X"02",X"0C",X"4C",X"02",X"F8",X"18",
		X"A8",X"C8",X"01",X"02",X"03",X"0E",X"4C",X"03",X"FF",X"F8",X"17",X"28",X"C0",X"00",X"01",X"02",
		X"0A",X"4C",X"02",X"F8",X"18",X"A8",X"C8",X"01",X"02",X"03",X"0C",X"4C",X"03",X"FF",X"F8",X"1D",
		X"28",X"B8",X"01",X"02",X"02",X"0A",X"4C",X"02",X"F8",X"1D",X"68",X"50",X"01",X"02",X"02",X"0C",
		X"4C",X"02",X"F8",X"18",X"A8",X"78",X"01",X"02",X"03",X"0E",X"4C",X"03",X"FF",X"F8",X"17",X"48",
		X"78",X"01",X"01",X"02",X"0A",X"4C",X"02",X"F8",X"17",X"A8",X"B0",X"00",X"01",X"02",X"0C",X"4C",
		X"02",X"FF",X"F8",X"17",X"28",X"A8",X"00",X"01",X"02",X"0A",X"4C",X"02",X"F8",X"17",X"68",X"80",
		X"01",X"01",X"02",X"0C",X"4C",X"02",X"F8",X"17",X"A8",X"20",X"00",X"01",X"02",X"0E",X"4C",X"02",
		X"FF",X"F8",X"18",X"28",X"98",X"01",X"02",X"03",X"0A",X"4C",X"03",X"F8",X"17",X"88",X"20",X"01",
		X"01",X"02",X"0C",X"4C",X"02",X"F8",X"1D",X"A8",X"C8",X"00",X"02",X"02",X"0E",X"4C",X"02",X"FF",
		X"F8",X"18",X"28",X"A8",X"01",X"02",X"03",X"0A",X"4C",X"03",X"F8",X"17",X"48",X"98",X"01",X"01",
		X"02",X"0C",X"4C",X"02",X"F8",X"17",X"88",X"B0",X"00",X"01",X"02",X"0E",X"4C",X"02",X"FF",X"F8",
		X"18",X"28",X"C0",X"01",X"02",X"03",X"0A",X"4C",X"03",X"F8",X"17",X"68",X"00",X"01",X"01",X"02",
		X"0C",X"4C",X"02",X"F8",X"17",X"A8",X"10",X"00",X"01",X"02",X"0E",X"4C",X"02",X"FF",X"F8",X"18",
		X"28",X"B8",X"01",X"02",X"03",X"0A",X"4C",X"03",X"F8",X"17",X"A8",X"28",X"00",X"01",X"02",X"0C",
		X"4C",X"02",X"FF",X"F8",X"18",X"28",X"C8",X"01",X"02",X"02",X"0A",X"4C",X"02",X"F8",X"1D",X"68",
		X"C0",X"01",X"02",X"02",X"0C",X"4C",X"02",X"F8",X"18",X"A8",X"30",X"01",X"02",X"03",X"0E",X"4C",
		X"02",X"FF",X"F8",X"17",X"28",X"30",X"00",X"01",X"02",X"0A",X"4C",X"02",X"F8",X"17",X"28",X"A0",
		X"00",X"01",X"02",X"0C",X"4C",X"02",X"F8",X"17",X"A8",X"40",X"00",X"01",X"02",X"0E",X"4C",X"02",
		X"FF",X"F5",X"A2",X"EF",X"A2",X"E9",X"A2",X"EC",X"A2",X"F2",X"A2",X"FB",X"A2",X"F8",X"A2",X"FE",
		X"A2",X"01",X"A3",X"04",X"A3",X"0A",X"A3",X"07",X"A3",X"0D",X"A3",X"13",X"A3",X"10",X"A3",X"01",
		X"A3",X"0A",X"A3",X"16",X"A3",X"07",X"A3",X"19",X"A3",X"01",X"07",X"40",X"01",X"06",X"40",X"01",
		X"06",X"30",X"01",X"05",X"30",X"01",X"05",X"40",X"01",X"05",X"30",X"01",X"06",X"30",X"01",X"06",
		X"40",X"01",X"05",X"30",X"01",X"05",X"30",X"01",X"04",X"30",X"01",X"04",X"30",X"01",X"04",X"30",
		X"01",X"04",X"30",X"01",X"04",X"30",X"01",X"02",X"40",X"01",X"02",X"30",X"34",X"A3",X"3A",X"A3",
		X"55",X"A3",X"37",X"A3",X"43",X"A3",X"3D",X"A3",X"40",X"A3",X"46",X"A3",X"49",X"A3",X"4C",X"A3",
		X"4F",X"A3",X"52",X"A3",X"02",X"02",X"01",X"07",X"03",X"04",X"07",X"04",X"03",X"00",X"04",X"01",
		X"07",X"06",X"03",X"02",X"02",X"02",X"06",X"03",X"02",X"03",X"06",X"00",X"04",X"05",X"01",X"01",
		X"06",X"06",X"01",X"06",X"06",X"00",X"03",X"06",X"70",X"A3",X"7C",X"A3",X"B2",X"A3",X"76",X"A3",
		X"8E",X"A3",X"82",X"A3",X"88",X"A3",X"94",X"A3",X"9A",X"A3",X"A0",X"A3",X"A6",X"A3",X"AC",X"A3",
		X"B8",X"A3",X"42",X"A4",X"B5",X"A4",X"BF",X"A4",X"BB",X"A5",X"8D",X"A6",X"5F",X"A7",X"DD",X"A7",
		X"46",X"A8",X"AF",X"A8",X"EB",X"A8",X"1D",X"A9",X"4F",X"A9",X"85",X"A9",X"8F",X"A9",X"99",X"A9",
		X"6B",X"AA",X"75",X"AA",X"7F",X"AA",X"91",X"AA",X"9B",X"AA",X"A5",X"AA",X"95",X"AB",X"5D",X"AC",
		X"FD",X"AC",X"DB",X"AD",X"E5",X"AD",X"4E",X"AE",X"A8",X"AE",X"F3",X"AE",X"3E",X"AF",X"BC",X"AF",
		X"11",X"B0",X"98",X"B0",X"0A",X"B1",X"69",X"B1",X"04",X"00",X"00",X"00",X"00",X"00",X"04",X"0A",
		X"05",X"03",X"05",X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"04",X"0A",X"05",X"03",X"05",X"04",
		X"04",X"00",X"00",X"00",X"00",X"00",X"04",X"0A",X"05",X"03",X"05",X"04",X"04",X"00",X"00",X"00",
		X"00",X"00",X"04",X"0A",X"05",X"03",X"05",X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"04",X"0A",
		X"05",X"03",X"05",X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"04",X"0A",X"05",X"03",X"05",X"04",
		X"04",X"00",X"00",X"00",X"00",X"00",X"04",X"0A",X"05",X"03",X"05",X"04",X"04",X"00",X"00",X"00",
		X"00",X"00",X"04",X"0A",X"05",X"03",X"05",X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"04",X"0A",
		X"05",X"03",X"05",X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"04",X"0A",X"05",X"03",X"05",X"04",
		X"04",X"00",X"00",X"00",X"00",X"00",X"04",X"0A",X"05",X"03",X"05",X"04",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"03",X"0A",X"06",X"0C",X"05",X"05",X"00",X"00",X"00",X"00",X"03",X"0A",X"06",X"0C",
		X"05",X"05",X"00",X"00",X"00",X"00",X"04",X"0A",X"06",X"0C",X"05",X"04",X"00",X"00",X"00",X"00",
		X"03",X"0A",X"06",X"0C",X"05",X"05",X"00",X"00",X"00",X"00",X"03",X"0A",X"06",X"0C",X"05",X"05",
		X"00",X"00",X"00",X"00",X"04",X"0A",X"06",X"0C",X"05",X"04",X"00",X"00",X"00",X"00",X"03",X"0A",
		X"06",X"0C",X"05",X"05",X"00",X"00",X"00",X"00",X"03",X"0A",X"06",X"0C",X"05",X"05",X"00",X"00",
		X"00",X"00",X"04",X"0A",X"06",X"0C",X"05",X"04",X"00",X"00",X"00",X"00",X"03",X"0A",X"06",X"0C",
		X"05",X"05",X"00",X"00",X"00",X"00",X"03",X"0A",X"06",X"0C",X"05",X"05",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"3C",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"06",
		X"0A",X"01",X"06",X"0C",X"05",X"06",X"0A",X"01",X"08",X"0B",X"05",X"06",X"0A",X"03",X"03",X"0A",
		X"05",X"06",X"0A",X"04",X"05",X"09",X"05",X"06",X"0A",X"04",X"04",X"08",X"05",X"06",X"09",X"00",
		X"02",X"07",X"05",X"06",X"09",X"0F",X"0A",X"06",X"05",X"06",X"09",X"05",X"0A",X"05",X"05",X"06",
		X"09",X"02",X"05",X"04",X"05",X"06",X"09",X"00",X"04",X"03",X"05",X"06",X"08",X"05",X"03",X"02",
		X"05",X"06",X"08",X"00",X"04",X"01",X"05",X"06",X"08",X"03",X"05",X"00",X"05",X"06",X"07",X"00",
		X"00",X"0F",X"04",X"06",X"07",X"09",X"0A",X"0E",X"04",X"06",X"06",X"00",X"00",X"0D",X"04",X"06",
		X"05",X"03",X"03",X"0C",X"04",X"06",X"05",X"00",X"00",X"0B",X"04",X"06",X"05",X"06",X"0E",X"0A",
		X"04",X"06",X"05",X"00",X"00",X"09",X"04",X"06",X"05",X"03",X"0D",X"08",X"04",X"06",X"05",X"00",
		X"0E",X"07",X"04",X"06",X"04",X"01",X"0F",X"06",X"04",X"06",X"04",X"00",X"07",X"05",X"04",X"06",
		X"04",X"02",X"03",X"04",X"04",X"06",X"04",X"05",X"06",X"03",X"04",X"06",X"04",X"09",X"09",X"02",
		X"04",X"06",X"03",X"08",X"06",X"01",X"04",X"06",X"03",X"07",X"02",X"00",X"04",X"06",X"03",X"07",
		X"07",X"0F",X"03",X"06",X"03",X"07",X"0D",X"0E",X"03",X"06",X"03",X"08",X"0B",X"0D",X"03",X"06",
		X"03",X"09",X"0A",X"0C",X"03",X"06",X"03",X"08",X"09",X"0B",X"03",X"06",X"02",X"0B",X"09",X"0A",
		X"03",X"06",X"02",X"0A",X"0A",X"09",X"03",X"06",X"02",X"09",X"0A",X"08",X"03",X"05",X"01",X"06",
		X"0B",X"07",X"03",X"06",X"01",X"03",X"0D",X"06",X"03",X"05",X"01",X"02",X"08",X"05",X"03",X"06",
		X"01",X"0F",X"00",X"04",X"03",X"FF",X"00",X"00",X"00",X"00",X"00",X"07",X"0A",X"07",X"0C",X"05",
		X"06",X"0A",X"08",X"0B",X"05",X"06",X"0A",X"04",X"0A",X"05",X"05",X"0A",X"05",X"09",X"05",X"07",
		X"0A",X"05",X"08",X"05",X"06",X"09",X"02",X"07",X"05",X"06",X"09",X"0B",X"06",X"05",X"05",X"09",
		X"0A",X"05",X"05",X"07",X"09",X"06",X"04",X"05",X"06",X"09",X"03",X"04",X"05",X"06",X"08",X"04",
		X"02",X"05",X"05",X"08",X"05",X"01",X"05",X"07",X"08",X"06",X"00",X"05",X"06",X"07",X"02",X"0F",
		X"04",X"06",X"07",X"0B",X"0E",X"04",X"05",X"03",X"08",X"0D",X"04",X"07",X"02",X"04",X"0C",X"04",
		X"06",X"02",X"01",X"0B",X"04",X"06",X"02",X"0F",X"0A",X"04",X"05",X"02",X"0F",X"09",X"04",X"07",
		X"02",X"0E",X"08",X"04",X"06",X"02",X"08",X"07",X"04",X"06",X"02",X"00",X"07",X"04",X"05",X"02",
		X"09",X"05",X"04",X"07",X"02",X"04",X"04",X"04",X"06",X"02",X"0B",X"03",X"04",X"06",X"02",X"0A",
		X"02",X"04",X"05",X"02",X"05",X"01",X"04",X"07",X"02",X"03",X"00",X"04",X"06",X"02",X"04",X"0F",
		X"03",X"05",X"02",X"0E",X"0E",X"03",X"05",X"02",X"0A",X"0D",X"03",X"07",X"02",X"0B",X"0C",X"03",
		X"06",X"02",X"0A",X"0B",X"03",X"05",X"02",X"0A",X"0A",X"03",X"05",X"02",X"0A",X"09",X"03",X"07",
		X"02",X"0B",X"08",X"03",X"06",X"01",X"0B",X"07",X"03",X"05",X"01",X"0E",X"06",X"03",X"05",X"01",
		X"09",X"05",X"03",X"07",X"01",X"01",X"04",X"03",X"FF",X"00",X"00",X"00",X"00",X"08",X"0A",X"05",
		X"0C",X"05",X"06",X"0A",X"08",X"0B",X"05",X"05",X"0A",X"02",X"0A",X"05",X"05",X"0A",X"05",X"09",
		X"05",X"08",X"0A",X"03",X"08",X"05",X"06",X"09",X"02",X"07",X"05",X"05",X"09",X"09",X"06",X"05",
		X"05",X"09",X"0A",X"05",X"05",X"08",X"09",X"03",X"04",X"05",X"06",X"09",X"03",X"03",X"05",X"05",
		X"08",X"02",X"02",X"05",X"05",X"08",X"01",X"01",X"05",X"08",X"08",X"04",X"00",X"05",X"06",X"07",
		X"06",X"0F",X"04",X"05",X"07",X"09",X"0E",X"04",X"05",X"06",X"06",X"0D",X"04",X"08",X"05",X"02",
		X"0C",X"04",X"06",X"05",X"06",X"0B",X"04",X"05",X"05",X"0D",X"0A",X"04",X"05",X"05",X"0C",X"09",
		X"04",X"08",X"05",X"0C",X"08",X"04",X"06",X"05",X"0D",X"07",X"04",X"05",X"04",X"0E",X"06",X"04",
		X"05",X"04",X"09",X"05",X"04",X"08",X"04",X"02",X"04",X"04",X"05",X"04",X"05",X"03",X"04",X"05",
		X"04",X"08",X"02",X"04",X"05",X"04",X"05",X"01",X"04",X"08",X"04",X"01",X"00",X"04",X"05",X"03",
		X"08",X"0F",X"03",X"05",X"03",X"0C",X"0E",X"03",X"05",X"03",X"04",X"0D",X"03",X"08",X"03",X"09",
		X"0C",X"03",X"05",X"02",X"01",X"09",X"03",X"05",X"02",X"08",X"08",X"03",X"05",X"02",X"08",X"07",
		X"03",X"08",X"02",X"09",X"06",X"03",X"05",X"01",X"03",X"05",X"03",X"05",X"01",X"0C",X"04",X"03",
		X"05",X"01",X"0D",X"02",X"03",X"08",X"01",X"0F",X"01",X"03",X"FF",X"00",X"00",X"00",X"00",X"01",
		X"05",X"0D",X"04",X"03",X"01",X"01",X"06",X"0C",X"08",X"00",X"01",X"01",X"06",X"0C",X"08",X"0D",
		X"00",X"01",X"07",X"06",X"0B",X"0B",X"00",X"01",X"07",X"0A",X"02",X"0B",X"00",X"01",X"08",X"09",
		X"04",X"0C",X"00",X"01",X"09",X"0C",X"08",X"0E",X"00",X"01",X"0B",X"0C",X"0B",X"0F",X"00",X"01",
		X"0D",X"0D",X"04",X"03",X"01",X"01",X"0F",X"04",X"09",X"06",X"01",X"01",X"0D",X"04",X"04",X"03",
		X"01",X"01",X"0B",X"0C",X"0B",X"0F",X"00",X"01",X"09",X"0C",X"08",X"0E",X"00",X"01",X"07",X"09",
		X"04",X"0C",X"00",X"01",X"05",X"0A",X"02",X"0B",X"00",X"01",X"04",X"06",X"0B",X"0B",X"00",X"01",
		X"03",X"04",X"09",X"0A",X"00",X"01",X"03",X"04",X"04",X"0A",X"00",X"01",X"02",X"0C",X"0B",X"09",
		X"00",X"01",X"01",X"0C",X"08",X"09",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"01",X"05",X"05",
		X"0F",X"00",X"01",X"05",X"09",X"0C",X"00",X"01",X"06",X"09",X"09",X"00",X"01",X"06",X"0C",X"07",
		X"00",X"01",X"08",X"03",X"07",X"00",X"01",X"09",X"05",X"08",X"00",X"01",X"0A",X"09",X"09",X"00",
		X"01",X"0C",X"0C",X"0B",X"00",X"01",X"0D",X"05",X"0F",X"00",X"01",X"0F",X"0A",X"02",X"01",X"01",
		X"0D",X"05",X"0F",X"00",X"01",X"0B",X"0C",X"0B",X"00",X"01",X"09",X"09",X"09",X"00",X"01",X"07",
		X"05",X"08",X"00",X"01",X"05",X"03",X"07",X"00",X"01",X"04",X"0C",X"07",X"00",X"01",X"03",X"0A",
		X"06",X"00",X"01",X"03",X"05",X"05",X"00",X"01",X"02",X"0C",X"04",X"00",X"01",X"01",X"0C",X"03",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"01",X"05",X"03",X"01",X"01",X"01",X"05",X"07",X"0E",X"00",
		X"01",X"06",X"07",X"0B",X"00",X"01",X"07",X"0A",X"09",X"00",X"01",X"08",X"01",X"09",X"00",X"01",
		X"09",X"03",X"0A",X"00",X"01",X"0A",X"07",X"0B",X"00",X"01",X"0C",X"0A",X"0D",X"00",X"01",X"0D",
		X"03",X"01",X"01",X"01",X"0F",X"08",X"04",X"01",X"01",X"0D",X"03",X"01",X"01",X"01",X"0B",X"0A",
		X"0D",X"00",X"01",X"09",X"07",X"0B",X"00",X"01",X"07",X"03",X"0A",X"00",X"01",X"05",X"01",X"09",
		X"00",X"01",X"04",X"0A",X"09",X"00",X"01",X"03",X"08",X"08",X"00",X"01",X"03",X"03",X"08",X"00",
		X"01",X"02",X"0A",X"07",X"00",X"01",X"01",X"07",X"07",X"00",X"FF",X"00",X"00",X"00",X"00",X"03",
		X"05",X"02",X"03",X"0E",X"02",X"03",X"05",X"03",X"03",X"0A",X"03",X"03",X"05",X"05",X"03",X"05",
		X"04",X"03",X"05",X"02",X"03",X"0E",X"02",X"03",X"05",X"03",X"03",X"0A",X"03",X"03",X"05",X"05",
		X"03",X"05",X"04",X"03",X"05",X"02",X"03",X"0E",X"02",X"03",X"05",X"03",X"03",X"0A",X"03",X"03",
		X"05",X"05",X"03",X"05",X"04",X"FF",X"00",X"00",X"00",X"00",X"00",X"04",X"05",X"06",X"0C",X"05",
		X"02",X"05",X"06",X"04",X"07",X"03",X"05",X"06",X"0A",X"08",X"04",X"05",X"06",X"0C",X"05",X"02",
		X"05",X"06",X"04",X"07",X"03",X"05",X"06",X"0A",X"08",X"04",X"05",X"06",X"0C",X"05",X"02",X"05",
		X"06",X"04",X"07",X"03",X"05",X"06",X"0A",X"08",X"FF",X"00",X"00",X"00",X"00",X"03",X"0A",X"0C",
		X"05",X"00",X"03",X"0A",X"04",X"07",X"00",X"03",X"0A",X"0A",X"08",X"00",X"03",X"0A",X"0C",X"05",
		X"00",X"03",X"0A",X"04",X"07",X"00",X"03",X"0A",X"0A",X"08",X"00",X"03",X"0A",X"0C",X"05",X"00",
		X"03",X"0A",X"04",X"07",X"00",X"03",X"0A",X"0A",X"08",X"00",X"FF",X"00",X"00",X"00",X"00",X"04",
		X"0A",X"08",X"01",X"07",X"01",X"01",X"0A",X"06",X"01",X"08",X"01",X"04",X"0A",X"0F",X"00",X"0D",
		X"01",X"01",X"0A",X"0C",X"05",X"0E",X"01",X"04",X"0A",X"0B",X"09",X"02",X"02",X"01",X"0A",X"0D",
		X"06",X"03",X"02",X"04",X"0A",X"02",X"03",X"0E",X"02",X"01",X"0A",X"02",X"04",X"0F",X"02",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"14",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"02",X"01",X"06",X"0C",X"05",X"00",X"02",
		X"01",X"06",X"0C",X"05",X"00",X"02",X"02",X"06",X"0C",X"05",X"00",X"02",X"02",X"06",X"0C",X"05",
		X"00",X"02",X"03",X"06",X"0C",X"05",X"00",X"02",X"03",X"06",X"0C",X"05",X"00",X"02",X"04",X"06",
		X"0C",X"05",X"00",X"02",X"04",X"06",X"0C",X"05",X"00",X"02",X"05",X"06",X"0C",X"05",X"00",X"02",
		X"05",X"06",X"0C",X"05",X"00",X"02",X"06",X"06",X"0C",X"05",X"00",X"02",X"06",X"06",X"0C",X"05",
		X"00",X"02",X"07",X"06",X"0C",X"05",X"00",X"02",X"07",X"06",X"0C",X"05",X"00",X"02",X"08",X"06",
		X"0C",X"05",X"00",X"02",X"08",X"06",X"0C",X"05",X"00",X"02",X"09",X"06",X"0C",X"05",X"00",X"02",
		X"09",X"06",X"0C",X"05",X"00",X"02",X"0A",X"06",X"0C",X"05",X"00",X"02",X"0A",X"06",X"0C",X"05",
		X"00",X"02",X"0B",X"06",X"0C",X"05",X"00",X"02",X"0B",X"06",X"0C",X"05",X"00",X"02",X"0C",X"06",
		X"0C",X"05",X"00",X"02",X"0C",X"06",X"0C",X"05",X"00",X"02",X"0D",X"06",X"0C",X"05",X"00",X"02",
		X"0D",X"06",X"0C",X"05",X"00",X"02",X"0E",X"06",X"0C",X"05",X"00",X"02",X"0E",X"06",X"0C",X"05",
		X"00",X"02",X"0F",X"06",X"0C",X"05",X"00",X"02",X"0F",X"06",X"0C",X"05",X"00",X"02",X"0F",X"06",
		X"0C",X"05",X"00",X"02",X"0F",X"06",X"0C",X"05",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"10",
		X"0F",X"0E",X"01",X"06",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"53",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"53",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"03",
		X"08",X"03",X"0D",X"0E",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"06",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"0B",X"0F",X"0F",X"00",X"0D",X"01",X"15",X"00",X"00",X"00",X"00",
		X"00",X"0B",X"0F",X"0F",X"00",X"0D",X"01",X"15",X"00",X"00",X"00",X"00",X"00",X"0B",X"0F",X"0F",
		X"00",X"0D",X"01",X"09",X"00",X"00",X"00",X"00",X"00",X"0B",X"0F",X"0B",X"0E",X"09",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"0B",X"0F",X"0F",X"00",X"0D",X"01",X"09",X"00",X"00",X"00",X"00",
		X"00",X"0B",X"0F",X"03",X"0D",X"0E",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"0B",X"0F",X"0B",
		X"09",X"02",X"02",X"15",X"00",X"00",X"00",X"00",X"00",X"0B",X"0F",X"0B",X"09",X"02",X"02",X"09",
		X"00",X"00",X"00",X"00",X"00",X"0B",X"0F",X"0B",X"09",X"02",X"02",X"01",X"00",X"00",X"00",X"00",
		X"00",X"1F",X"0F",X"0F",X"00",X"0D",X"01",X"21",X"00",X"00",X"00",X"00",X"00",X"0B",X"0F",X"0B",
		X"0E",X"09",X"01",X"15",X"00",X"00",X"00",X"00",X"00",X"0B",X"0F",X"0B",X"0E",X"09",X"01",X"09",
		X"00",X"00",X"00",X"00",X"00",X"0B",X"0F",X"0F",X"00",X"0D",X"01",X"01",X"00",X"00",X"00",X"00",
		X"00",X"0B",X"0F",X"03",X"0D",X"0E",X"01",X"15",X"00",X"00",X"00",X"00",X"00",X"0B",X"0F",X"0F",
		X"00",X"0D",X"01",X"09",X"00",X"00",X"00",X"00",X"00",X"0B",X"0F",X"0B",X"0E",X"09",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"08",X"01",X"07",X"01",X"11",X"00",X"00",X"00",X"00",
		X"00",X"04",X"0F",X"09",X"09",X"0B",X"02",X"0C",X"0F",X"02",X"03",X"0E",X"02",X"10",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"0F",X"08",X"01",X"07",X"01",X"10",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"0B",X"0F",X"01",X"07",X"01",X"15",X"00",X"00",X"00",X"00",X"0B",
		X"0F",X"01",X"07",X"01",X"15",X"00",X"00",X"00",X"00",X"0B",X"0F",X"01",X"07",X"01",X"09",X"00",
		X"00",X"00",X"00",X"0B",X"0F",X"0C",X"05",X"01",X"01",X"00",X"00",X"00",X"00",X"0B",X"0F",X"01",
		X"07",X"01",X"09",X"00",X"00",X"00",X"00",X"0B",X"0F",X"0E",X"09",X"01",X"01",X"00",X"00",X"00",
		X"00",X"0B",X"0F",X"00",X"0D",X"01",X"15",X"00",X"00",X"00",X"00",X"0B",X"0F",X"00",X"0D",X"01",
		X"09",X"00",X"00",X"00",X"00",X"0B",X"0F",X"00",X"0D",X"01",X"01",X"00",X"00",X"00",X"00",X"1F",
		X"0F",X"01",X"07",X"01",X"21",X"00",X"00",X"00",X"00",X"0B",X"0F",X"0C",X"05",X"01",X"15",X"00",
		X"00",X"00",X"00",X"0B",X"0F",X"0C",X"05",X"01",X"09",X"00",X"00",X"00",X"00",X"0B",X"0F",X"01",
		X"07",X"01",X"01",X"00",X"00",X"00",X"00",X"0B",X"0F",X"0E",X"09",X"01",X"15",X"00",X"00",X"00",
		X"00",X"0B",X"0F",X"01",X"07",X"01",X"09",X"00",X"00",X"00",X"00",X"0B",X"0F",X"0C",X"05",X"01",
		X"01",X"00",X"00",X"00",X"00",X"0F",X"0F",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"04",
		X"0F",X"00",X"00",X"00",X"0C",X"0F",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"0F",X"0F",
		X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"0F",X"06",X"08",
		X"0B",X"00",X"11",X"00",X"00",X"00",X"00",X"0F",X"06",X"0A",X"08",X"00",X"11",X"00",X"00",X"00",
		X"00",X"0F",X"06",X"08",X"0B",X"00",X"11",X"00",X"00",X"00",X"00",X"0F",X"06",X"0A",X"08",X"00",
		X"11",X"00",X"00",X"00",X"00",X"0F",X"06",X"08",X"0B",X"00",X"11",X"00",X"00",X"00",X"00",X"0F",
		X"06",X"0A",X"08",X"00",X"11",X"00",X"00",X"00",X"00",X"0F",X"06",X"08",X"0B",X"00",X"11",X"00",
		X"00",X"00",X"00",X"0F",X"06",X"0A",X"08",X"00",X"11",X"00",X"00",X"00",X"00",X"0F",X"06",X"0F",
		X"0C",X"00",X"11",X"00",X"00",X"00",X"00",X"0F",X"06",X"0A",X"08",X"00",X"11",X"00",X"00",X"00",
		X"00",X"0F",X"06",X"0B",X"09",X"00",X"11",X"00",X"00",X"00",X"00",X"0F",X"06",X"0E",X"0A",X"00",
		X"11",X"00",X"00",X"00",X"00",X"0F",X"06",X"08",X"0B",X"00",X"11",X"00",X"00",X"00",X"00",X"0F",
		X"06",X"0A",X"08",X"00",X"11",X"00",X"00",X"00",X"00",X"0F",X"06",X"08",X"0B",X"00",X"01",X"00",
		X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"03",X"0C",X"08",
		X"01",X"07",X"01",X"01",X"0A",X"08",X"01",X"07",X"01",X"01",X"08",X"08",X"01",X"07",X"01",X"01",
		X"06",X"08",X"01",X"07",X"01",X"01",X"04",X"08",X"01",X"07",X"01",X"01",X"02",X"08",X"01",X"07",
		X"01",X"02",X"00",X"00",X"00",X"00",X"00",X"02",X"0C",X"0C",X"06",X"03",X"01",X"01",X"0A",X"0C",
		X"06",X"03",X"01",X"01",X"08",X"0C",X"06",X"03",X"01",X"01",X"06",X"0C",X"06",X"03",X"01",X"02",
		X"0C",X"0D",X"04",X"01",X"01",X"01",X"0A",X"0D",X"04",X"01",X"01",X"01",X"08",X"0D",X"04",X"01",
		X"01",X"01",X"06",X"0D",X"04",X"01",X"01",X"03",X"0C",X"0C",X"08",X"0E",X"00",X"01",X"0A",X"0C",
		X"08",X"0E",X"00",X"01",X"08",X"0C",X"08",X"0E",X"00",X"01",X"06",X"0C",X"08",X"0E",X"00",X"01",
		X"04",X"0C",X"08",X"0E",X"00",X"01",X"02",X"0C",X"08",X"0E",X"00",X"02",X"00",X"00",X"00",X"00",
		X"00",X"03",X"0C",X"05",X"0F",X"0C",X"00",X"01",X"0A",X"05",X"0F",X"0C",X"00",X"01",X"08",X"05",
		X"0F",X"0C",X"00",X"01",X"06",X"05",X"0F",X"0C",X"00",X"01",X"04",X"05",X"0F",X"0C",X"00",X"01",
		X"02",X"05",X"0F",X"0C",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"02",X"0C",X"0C",X"08",X"0B",
		X"00",X"02",X"0A",X"0C",X"08",X"0B",X"00",X"02",X"08",X"0C",X"08",X"0B",X"00",X"02",X"06",X"0C",
		X"08",X"0B",X"00",X"02",X"04",X"0C",X"08",X"0B",X"00",X"02",X"02",X"0C",X"08",X"0B",X"00",X"08",
		X"01",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"3C",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"06",X"05",X"0B",X"07",X"00",X"02",X"04",X"0B",X"07",X"00",X"02",
		X"03",X"0B",X"07",X"00",X"02",X"02",X"0B",X"07",X"00",X"08",X"01",X"0B",X"07",X"00",X"06",X"05",
		X"0A",X"08",X"00",X"02",X"04",X"0A",X"08",X"00",X"02",X"03",X"0A",X"08",X"00",X"02",X"02",X"0A",
		X"08",X"00",X"08",X"01",X"0A",X"08",X"00",X"02",X"05",X"0C",X"05",X"00",X"02",X"05",X"0C",X"05",
		X"00",X"02",X"04",X"0C",X"05",X"00",X"02",X"04",X"0C",X"05",X"00",X"02",X"03",X"0C",X"05",X"00",
		X"02",X"03",X"0C",X"05",X"00",X"02",X"02",X"0C",X"05",X"00",X"02",X"02",X"0C",X"05",X"00",X"02",
		X"01",X"0C",X"05",X"00",X"02",X"01",X"0C",X"05",X"00",X"FF",X"00",X"00",X"00",X"00",X"0C",X"0D",
		X"0C",X"08",X"0B",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"07",X"0D",X"07",X"0A",X"08",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"07",X"0D",X"07",X"0A",X"08",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"0D",X"06",X"0B",X"09",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"0F",X"0D",
		X"07",X"0A",X"08",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"0C",X"0D",X"07",X"0E",X"0A",X"00",
		X"04",X"00",X"00",X"00",X"00",X"00",X"10",X"0D",X"0C",X"08",X"0B",X"00",X"20",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"0C",X"0D",X"01",X"07",X"01",X"04",X"00",X"00",
		X"00",X"00",X"07",X"0D",X"04",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"07",X"0D",X"04",X"01",
		X"01",X"01",X"00",X"00",X"00",X"00",X"0F",X"0D",X"06",X"03",X"01",X"01",X"00",X"00",X"00",X"00",
		X"0F",X"0D",X"04",X"01",X"01",X"11",X"00",X"00",X"00",X"00",X"0C",X"0D",X"0C",X"05",X"01",X"04",
		X"00",X"00",X"00",X"00",X"10",X"0D",X"01",X"07",X"01",X"20",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"0C",X"0D",X"08",X"0B",X"00",X"04",X"00",X"00",X"00",X"00",X"07",X"0D",X"0A",
		X"08",X"00",X"01",X"00",X"00",X"00",X"00",X"07",X"0D",X"0A",X"08",X"00",X"01",X"00",X"00",X"00",
		X"00",X"0F",X"0D",X"0B",X"09",X"00",X"01",X"00",X"00",X"00",X"00",X"0F",X"0D",X"0A",X"08",X"00",
		X"11",X"00",X"00",X"00",X"00",X"0C",X"0D",X"09",X"0B",X"02",X"04",X"00",X"00",X"00",X"00",X"10",
		X"0D",X"03",X"0E",X"02",X"20",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"10",X"0F",
		X"08",X"01",X"07",X"01",X"10",X"00",X"00",X"00",X"00",X"00",X"10",X"0F",X"0F",X"00",X"0D",X"01",
		X"10",X"00",X"00",X"00",X"00",X"00",X"08",X"0F",X"0B",X"09",X"02",X"02",X"08",X"00",X"00",X"00",
		X"00",X"00",X"08",X"0F",X"0F",X"00",X"0D",X"01",X"08",X"00",X"00",X"00",X"00",X"00",X"10",X"0F",
		X"08",X"01",X"07",X"01",X"10",X"00",X"00",X"00",X"00",X"00",X"08",X"0F",X"07",X"0D",X"06",X"02",
		X"08",X"00",X"00",X"00",X"00",X"00",X"08",X"0F",X"0B",X"09",X"02",X"02",X"08",X"00",X"00",X"00",
		X"00",X"00",X"08",X"0F",X"07",X"0D",X"06",X"02",X"08",X"00",X"00",X"00",X"00",X"00",X"08",X"0F",
		X"09",X"09",X"0B",X"02",X"08",X"00",X"00",X"00",X"00",X"00",X"20",X"0F",X"02",X"03",X"0E",X"02",
		X"50",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"10",X"08",X"04",X"01",
		X"01",X"10",X"00",X"00",X"00",X"00",X"10",X"08",X"01",X"07",X"01",X"10",X"00",X"00",X"00",X"00",
		X"08",X"08",X"00",X"0D",X"01",X"08",X"00",X"00",X"00",X"00",X"08",X"08",X"01",X"07",X"01",X"08",
		X"00",X"00",X"00",X"00",X"10",X"08",X"04",X"01",X"01",X"10",X"00",X"00",X"00",X"00",X"10",X"08",
		X"0D",X"0E",X"01",X"10",X"00",X"00",X"00",X"00",X"10",X"08",X"0D",X"0E",X"01",X"10",X"00",X"00",
		X"00",X"00",X"20",X"08",X"00",X"0D",X"01",X"50",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"08",X"08",X"08",X"0B",X"00",X"08",X"00",X"00",X"00",X"00",X"08",X"08",X"04",X"01",X"01",
		X"08",X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"0B",X"00",X"08",X"00",X"00",X"00",X"00",X"08",
		X"08",X"04",X"01",X"01",X"08",X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"0B",X"00",X"08",X"00",
		X"00",X"00",X"00",X"08",X"08",X"04",X"01",X"01",X"08",X"00",X"00",X"00",X"00",X"08",X"08",X"08",
		X"0B",X"00",X"08",X"00",X"00",X"00",X"00",X"08",X"08",X"04",X"01",X"01",X"08",X"00",X"00",X"00",
		X"00",X"08",X"08",X"08",X"0B",X"00",X"08",X"00",X"00",X"00",X"00",X"08",X"08",X"04",X"01",X"01",
		X"08",X"00",X"00",X"00",X"00",X"08",X"08",X"06",X"03",X"01",X"08",X"00",X"00",X"00",X"00",X"08",
		X"08",X"0A",X"08",X"00",X"08",X"00",X"00",X"00",X"00",X"20",X"08",X"08",X"0B",X"00",X"50",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"1F",X"0E",X"02",X"03",X"0E",X"02",X"01",X"00",
		X"00",X"00",X"00",X"00",X"0B",X"0E",X"09",X"09",X"0B",X"02",X"01",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"0E",X"07",X"02",X"09",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"0B",X"0E",X"07",X"0D",
		X"06",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"0A",X"0E",X"0B",X"09",X"02",X"02",X"02",X"00",
		X"00",X"00",X"00",X"00",X"0A",X"0E",X"03",X"0D",X"0E",X"01",X"02",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"0E",X"0F",X"00",X"0D",X"01",X"02",X"00",X"00",X"00",X"00",X"00",X"0A",X"0E",X"0B",X"0E",
		X"09",X"01",X"02",X"00",X"00",X"00",X"00",X"00",X"0B",X"0E",X"08",X"01",X"07",X"01",X"50",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"1F",X"06",X"09",X"02",X"02",X"01",
		X"00",X"00",X"00",X"00",X"0B",X"06",X"09",X"02",X"02",X"01",X"00",X"00",X"00",X"00",X"1F",X"06",
		X"09",X"02",X"02",X"01",X"00",X"00",X"00",X"00",X"0B",X"06",X"0D",X"0E",X"01",X"01",X"00",X"00",
		X"00",X"00",X"0A",X"06",X"0E",X"09",X"01",X"02",X"00",X"00",X"00",X"00",X"0A",X"06",X"0E",X"09",
		X"01",X"02",X"00",X"00",X"00",X"00",X"0A",X"06",X"09",X"04",X"01",X"02",X"00",X"00",X"00",X"00",
		X"0A",X"06",X"0C",X"05",X"01",X"02",X"00",X"00",X"00",X"00",X"0B",X"06",X"01",X"07",X"01",X"50",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"1F",X"06",X"08",X"0B",X"00",X"01",X"00",
		X"00",X"00",X"00",X"0B",X"06",X"0F",X"0C",X"00",X"01",X"00",X"00",X"00",X"00",X"1F",X"06",X"08",
		X"0E",X"00",X"01",X"00",X"00",X"00",X"00",X"0B",X"06",X"06",X"0F",X"00",X"01",X"00",X"00",X"00",
		X"00",X"0A",X"06",X"04",X"01",X"01",X"02",X"00",X"00",X"00",X"00",X"0A",X"06",X"06",X"03",X"01",
		X"02",X"00",X"00",X"00",X"00",X"0A",X"06",X"09",X"04",X"01",X"02",X"00",X"00",X"00",X"00",X"0A",
		X"06",X"0C",X"05",X"01",X"02",X"00",X"00",X"00",X"00",X"0B",X"06",X"01",X"07",X"01",X"50",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"32",X"C0",X"50",X"DD",X"21",X"52",X"B3",X"DD",
		X"6E",X"00",X"DD",X"7E",X"01",X"67",X"B5",X"CA",X"B0",X"B2",X"DD",X"4E",X"02",X"DD",X"46",X"03",
		X"54",X"5D",X"36",X"0F",X"13",X"0B",X"ED",X"B0",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"DD",X"4E",
		X"02",X"DD",X"46",X"03",X"0B",X"32",X"C0",X"50",X"3E",X"55",X"77",X"BE",X"20",X"3E",X"3E",X"AA",
		X"77",X"BE",X"20",X"38",X"78",X"D9",X"47",X"D9",X"79",X"D9",X"4F",X"D9",X"7C",X"D9",X"67",X"D9",
		X"7D",X"D9",X"6F",X"CB",X"28",X"CB",X"19",X"78",X"B1",X"28",X"08",X"23",X"54",X"5D",X"36",X"0F",
		X"13",X"ED",X"B0",X"D9",X"3E",X"AA",X"BE",X"20",X"0D",X"23",X"0B",X"78",X"B1",X"20",X"C6",X"11",
		X"04",X"00",X"DD",X"19",X"18",X"99",X"EB",X"21",X"94",X"B3",X"18",X"04",X"EB",X"21",X"83",X"B3",
		X"D9",X"01",X"FF",X"03",X"21",X"00",X"40",X"11",X"01",X"40",X"36",X"0F",X"ED",X"B0",X"01",X"FF",
		X"03",X"21",X"00",X"44",X"11",X"01",X"44",X"36",X"0F",X"ED",X"B0",X"32",X"C0",X"50",X"D9",X"7A",
		X"D9",X"67",X"D9",X"7B",X"D9",X"6F",X"D9",X"11",X"8A",X"41",X"06",X"11",X"7E",X"12",X"23",X"13",
		X"10",X"FA",X"D9",X"0E",X"04",X"11",X"9B",X"41",X"06",X"04",X"AF",X"CB",X"25",X"CB",X"14",X"CB",
		X"17",X"10",X"F8",X"13",X"FE",X"0A",X"38",X"02",X"C6",X"06",X"12",X"0D",X"20",X"EA",X"01",X"FF",
		X"7F",X"32",X"C0",X"50",X"DD",X"CB",X"00",X"46",X"DD",X"CB",X"00",X"46",X"DD",X"CB",X"00",X"46",
		X"DD",X"CB",X"00",X"46",X"DD",X"CB",X"00",X"46",X"0B",X"78",X"B1",X"20",X"E4",X"C3",X"00",X"00",
		X"01",X"FF",X"03",X"21",X"00",X"40",X"11",X"00",X"40",X"13",X"36",X"0F",X"ED",X"B0",X"01",X"FF",
		X"03",X"21",X"00",X"44",X"11",X"01",X"44",X"36",X"0F",X"ED",X"B0",X"06",X"0C",X"11",X"8A",X"41",
		X"21",X"6B",X"B3",X"7E",X"12",X"13",X"23",X"10",X"FA",X"06",X"08",X"21",X"00",X"00",X"11",X"60",
		X"B3",X"0E",X"00",X"32",X"C0",X"50",X"79",X"86",X"4F",X"2C",X"20",X"F7",X"24",X"7C",X"E6",X"0F",
		X"20",X"F1",X"1A",X"B9",X"20",X"3A",X"13",X"7C",X"FE",X"40",X"20",X"02",X"26",X"80",X"10",X"E1",
		X"11",X"CA",X"41",X"06",X"0C",X"21",X"77",X"B3",X"7E",X"12",X"13",X"23",X"10",X"FA",X"01",X"FF",
		X"7F",X"32",X"C0",X"50",X"DD",X"CB",X"00",X"46",X"DD",X"CB",X"00",X"46",X"DD",X"CB",X"00",X"46",
		X"DD",X"CB",X"00",X"46",X"DD",X"CB",X"00",X"46",X"0B",X"78",X"B1",X"20",X"E4",X"C3",X"A4",X"06",
		X"7C",X"E6",X"F0",X"0F",X"0F",X"0F",X"0F",X"FE",X"0A",X"38",X"02",X"C6",X"06",X"08",X"11",X"CA",
		X"41",X"21",X"A5",X"B3",X"06",X"13",X"7E",X"12",X"23",X"13",X"10",X"FA",X"13",X"08",X"12",X"C3",
		X"91",X"B2",X"00",X"4C",X"00",X"04",X"00",X"40",X"00",X"04",X"00",X"44",X"00",X"04",X"00",X"00",
		X"3A",X"9C",X"D3",X"E9",X"90",X"1A",X"5C",X"00",X"4A",X"FF",X"FF",X"21",X"10",X"1C",X"0A",X"12",
		X"17",X"14",X"12",X"1A",X"0A",X"1E",X"1A",X"21",X"1E",X"1C",X"0A",X"12",X"17",X"14",X"12",X"1A",
		X"0A",X"1E",X"1A",X"21",X"10",X"1C",X"0A",X"12",X"17",X"14",X"12",X"1A",X"0A",X"26",X"21",X"18",
		X"23",X"14",X"0A",X"0A",X"21",X"10",X"1C",X"0A",X"12",X"17",X"14",X"12",X"1A",X"0A",X"11",X"21",
		X"18",X"13",X"16",X"14",X"0A",X"21",X"1E",X"1C",X"0A",X"12",X"17",X"14",X"12",X"1A",X"0A",X"14",
		X"21",X"21",X"1E",X"21",X"0A",X"21",X"1E",X"1C",X"D1",X"E9",X"11",X"B1",X"3B",X"A4",X"85",X"93",
		X"56",X"FF",X"C7",X"2D",X"F8",X"30",X"20",X"9A",X"C1",X"59",X"92",X"69",X"9F",X"E9",X"03",X"DB",
		X"17",X"C3",X"BB",X"94",X"FC",X"19",X"45",X"FF",X"79",X"2B",X"FE",X"FC",X"24",X"B3",X"EB",X"21",
		X"9F",X"E4",X"34",X"E8",X"BB",X"DC",X"AC",X"9E",X"B1",X"3B",X"20",X"81",X"F8",X"A3",X"A9",X"00",
		X"98",X"F5",X"B0",X"E4",X"0F",X"2B",X"30",X"7D",X"BA",X"83",X"4C",X"79",X"FA",X"19",X"A9",X"31",
		X"A6",X"09",X"1E",X"21",X"20",X"B1",X"24",X"A9",X"23",X"91",X"16",X"6A",X"DA",X"7B",X"36",X"51",
		X"30",X"AB",X"0F",X"B3",X"69",X"20",X"36",X"81",X"0F",X"C1",X"A0",X"0D",X"64",X"61",X"72",X"71",
		X"74",X"35",X"39",X"18",X"29",X"C1",X"19",X"A7",X"23",X"50",X"F1",X"55",X"09",X"34",X"67",X"30",
		X"86",X"2C",X"41",X"6C",X"52",X"67",X"41",X"B7",X"07",X"30",X"79",X"05",X"CF",X"20",X"C7",X"41",
		X"31",X"21",X"14",X"E1",X"20",X"5A",X"00",X"A0",X"B4",X"8B",X"50",X"00",X"9D",X"34",X"60",X"25",
		X"A0",X"B0",X"2C",X"02",X"12",X"71",X"4D",X"20",X"BB",X"E2",X"A3",X"09",X"B1",X"00",X"5D",X"B5",
		X"83",X"36",X"52",X"08",X"71",X"10",X"28",X"3C",X"A4",X"55",X"45",X"C1",X"30",X"95",X"19",X"AE",
		X"49",X"68",X"61",X"F0",X"20",X"35",X"26",X"B0",X"71",X"E3",X"81",X"28",X"80",X"3D",X"5B",X"08",
		X"CC",X"1F",X"A1",X"FE",X"6F",X"F4",X"4B",X"5F",X"A4",X"8F",X"FC",X"DC",X"3F",X"FB",X"97",X"FB",
		X"42",X"1E",X"AE",X"BA",X"D7",X"57",X"9F",X"7A",X"BC",X"E3",X"FE",X"1E",X"5F",X"CD",X"8A",X"C8",
		X"D3",X"23",X"FE",X"26",X"0B",X"B2",X"94",X"DC",X"CA",X"0A",X"B3",X"FE",X"56",X"A3",X"E2",X"F4",
		X"F6",X"CD",X"56",X"87",X"5C",X"76",X"D4",X"B8",X"D4",X"AF",X"DF",X"F4",X"B4",X"5F",X"42",X"FD",
		X"EB",X"F1",X"AB",X"07",X"D5",X"D5",X"3C",X"72",X"9B",X"FF",X"BA",X"71",X"BB",X"7F",X"75",X"37",
		X"55",X"3D",X"54",X"9C",X"DF",X"53",X"6F",X"F6",X"67",X"0A",X"BC",X"4B",X"4D",X"2D",X"95",X"96",
		X"BD",X"B9",X"1C",X"6D",X"96",X"F7",X"BD",X"5F",X"7D",X"77",X"9F",X"0A",X"DB",X"56",X"92",X"DE",
		X"FF",X"59",X"FF",X"4B",X"57",X"E6",X"95",X"B3",X"7A",X"F3",X"49",X"52",X"2E",X"55",X"6E",X"93",
		X"B9",X"05",X"7B",X"0C",X"48",X"BC",X"E0",X"BE",X"51",X"CD",X"29",X"11",X"D9",X"E9",X"01",X"70",
		X"04",X"70",X"05",X"81",X"A1",X"99",X"59",X"B4",X"A0",X"6A",X"10",X"31",X"43",X"71",X"AC",X"2A",
		X"33",X"05",X"89",X"B7",X"B1",X"31",X"1F",X"63",X"08",X"25",X"73",X"A9",X"30",X"30",X"7F",X"81",
		X"8D",X"14",X"AB",X"02",X"91",X"73",X"1B",X"71",X"85",X"EA",X"0E",X"28",X"55",X"58",X"39",X"50",
		X"94",X"11",X"05",X"E0",X"DC",X"0A",X"20",X"03",X"10",X"46",X"14",X"10",X"C1",X"C0",X"E8",X"1B",
		X"2A",X"A9",X"A4",X"E1",X"D2",X"19",X"87",X"01",X"A0",X"80",X"25",X"26",X"73",X"D8",X"73",X"A8",
		X"41",X"65",X"E4",X"30",X"A0",X"20",X"89",X"B1",X"30",X"A0",X"88",X"52",X"6A",X"25",X"38",X"25",
		X"E0",X"22",X"44",X"B5",X"60",X"8C",X"9C",X"5C",X"B2",X"84",X"43",X"05",X"A2",X"34",X"05",X"28",
		X"4A",X"3F",X"69",X"D3",X"3E",X"DF",X"D3",X"4C",X"CD",X"D0",X"3F",X"DA",X"5F",X"5E",X"BE",X"F7",
		X"67",X"D3",X"2F",X"ED",X"D3",X"5C",X"9A",X"ED",X"52",X"C6",X"56",X"FF",X"76",X"DC",X"BB",X"EF",
		X"C7",X"9F",X"EC",X"CA",X"7D",X"1E",X"79",X"F4",X"8A",X"02",X"3C",X"D7",X"BF",X"76",X"B8",X"54",
		X"E9",X"E9",X"FC",X"02",X"66",X"FF",X"FC",X"E0",X"AA",X"AD",X"9E",X"F8",X"EB",X"1F",X"C9",X"77",
		X"98",X"F7",X"3F",X"8F",X"E6",X"55",X"AA",X"93",X"4C",X"6F",X"DF",X"D9",X"93",X"CB",X"7C",X"3F",
		X"B5",X"97",X"2E",X"83",X"CF",X"FF",X"F5",X"CE",X"E5",X"1F",X"7B",X"3B",X"77",X"D6",X"C2",X"4F",
		X"7F",X"0C",X"BE",X"EF",X"BB",X"67",X"DF",X"EE",X"5A",X"AF",X"1F",X"3E",X"37",X"FF",X"C6",X"5E",
		X"DF",X"EF",X"BF",X"D7",X"92",X"6F",X"D5",X"7F",X"FE",X"EE",X"6B",X"D9",X"77",X"4F",X"DE",X"6B",
		X"DE",X"D3",X"87",X"5E",X"A6",X"D7",X"04",X"46",X"5A",X"44",X"2E",X"80",X"26",X"76",X"69",X"2F",
		X"D6",X"FB",X"C7",X"07",X"16",X"05",X"96",X"45",X"4B",X"E2",X"CF",X"04",X"0C",X"AC",X"2F",X"5E",
		X"D1",X"32",X"9F",X"C3",X"BE",X"26",X"2F",X"6A",X"62",X"36",X"C2",X"02",X"76",X"E7",X"0F",X"BE",
		X"97",X"2E",X"DE",X"2D",X"1F",X"4F",X"A3",X"DF",X"6B",X"5F",X"0F",X"8B",X"C2",X"42",X"27",X"05",
		X"2C",X"81",X"01",X"2E",X"86",X"0C",X"4E",X"EB",X"65",X"04",X"56",X"5E",X"16",X"89",X"82",X"A2",
		X"74",X"C4",X"3A",X"97",X"8E",X"B8",X"47",X"3E",X"24",X"C1",X"AB",X"26",X"0B",X"AC",X"E7",X"32",
		X"21",X"7E",X"42",X"57",X"82",X"A3",X"5B",X"05",X"1F",X"CA",X"03",X"EF",X"A6",X"04",X"80",X"46",
		X"92",X"2E",X"86",X"02",X"B3",X"4A",X"4B",X"0F",X"E7",X"AB",X"80",X"9E",X"2A",X"56",X"87",X"4D",
		X"B0",X"79",X"75",X"5C",X"A3",X"2C",X"11",X"CF",X"7E",X"D9",X"72",X"B9",X"D8",X"3D",X"BE",X"E8",
		X"B1",X"F5",X"79",X"F1",X"78",X"B0",X"F8",X"A0",X"D2",X"39",X"F9",X"F8",X"3C",X"72",X"FC",X"E1",
		X"C9",X"E9",X"B1",X"DE",X"B1",X"C4",X"AD",X"B9",X"2B",X"60",X"D3",X"C8",X"EC",X"B5",X"FB",X"F9",
		X"70",X"69",X"1A",X"FD",X"7D",X"DB",X"A9",X"39",X"9D",X"29",X"BA",X"B1",X"00",X"BD",X"3E",X"99",
		X"74",X"F0",X"23",X"A9",X"BB",X"34",X"8B",X"F5",X"F0",X"B5",X"68",X"F0",X"53",X"30",X"F1",X"E7",
		X"A7",X"82",X"FD",X"31",X"B8",X"82",X"D0",X"FF",X"EE",X"D0",X"1A",X"A0",X"F1",X"6D",X"ED",X"F1",
		X"18",X"E7",X"D8",X"F2",X"A1",X"A5",X"FE",X"ED",X"FB",X"D0",X"D9",X"F9",X"F8",X"BB",X"7C",X"4B",
		X"75",X"85",X"74",X"20",X"25",X"66",X"95",X"79",X"69",X"69",X"DF",X"A8",X"31",X"31",X"31",X"DB",
		X"26",X"5B",X"71",X"6F",X"8E",X"16",X"C6",X"63",X"23",X"27",X"43",X"53",X"96",X"46",X"07",X"D6",
		X"58",X"EE",X"CE",X"C4",X"42",X"43",X"04",X"45",X"4F",X"42",X"15",X"46",X"DF",X"07",X"37",X"24",
		X"22",X"6A",X"56",X"41",X"05",X"17",X"D1",X"0F",X"02",X"0B",X"46",X"ED",X"E1",X"AF",X"04",X"D7",
		X"27",X"0E",X"02",X"96",X"17",X"0F",X"07",X"4F",X"0E",X"EC",X"D5",X"4F",X"4A",X"E7",X"E5",X"37",
		X"8A",X"4C",X"8B",X"8D",X"26",X"F5",X"6A",X"15",X"E7",X"97",X"17",X"2E",X"94",X"EB",X"89",X"42",
		X"1C",X"8F",X"06",X"8C",X"2F",X"50",X"37",X"FE",X"2A",X"8F",X"B1",X"05",X"CF",X"10",X"7E",X"E9",
		X"06",X"C7",X"62",X"2F",X"9C",X"56",X"CE",X"6D",X"77",X"0F",X"D2",X"22",X"9B",X"3E",X"2E",X"8B",
		X"76",X"DF",X"92",X"8E",X"44",X"4F",X"D0",X"0E",X"0B",X"AE",X"54",X"5A",X"48",X"56",X"40",X"47",
		X"7E",X"88",X"7D",X"B8",X"92",X"3A",X"FB",X"E8",X"71",X"FF",X"58",X"F9",X"85",X"E9",X"91",X"F7",
		X"AC",X"C5",X"20",X"2F",X"CB",X"F0",X"5C",X"70",X"70",X"BA",X"51",X"B9",X"11",X"A1",X"AC",X"B2",
		X"BD",X"59",X"35",X"58",X"EB",X"21",X"B9",X"B0",X"AC",X"FA",X"C9",X"7D",X"29",X"6A",X"39",X"59",
		X"8C",X"58",X"B4",X"21",X"C0",X"F1",X"76",X"BB",X"F1",X"69",X"5B",X"C8",X"D8",X"79",X"9C",X"F4",
		X"0E",X"2A",X"A9",X"7F",X"35",X"39",X"C9",X"28",X"B7",X"F2",X"38",X"78",X"9A",X"BA",X"E1",X"39",
		X"FD",X"A0",X"A9",X"65",X"FC",X"B9",X"E1",X"1C",X"39",X"D1",X"E1",X"B5",X"85",X"F0",X"C4",X"73",
		X"AE",X"F8",X"37",X"B1",X"78",X"90",X"B1",X"51",X"7F",X"21",X"A8",X"76",X"D9",X"BC",X"FD",X"B8",
		X"EC",X"48",X"3D",X"B7",X"B4",X"99",X"82",X"18",X"FA",X"B1",X"5B",X"7B",X"39",X"8D",X"A9",X"FD",
		X"DF",X"E6",X"FF",X"5E",X"42",X"F7",X"7B",X"CB",X"E7",X"FF",X"F7",X"CF",X"DD",X"AF",X"D7",X"DE",
		X"47",X"6F",X"CF",X"9F",X"67",X"F5",X"1B",X"AD",X"63",X"47",X"DF",X"BF",X"C5",X"FD",X"DF",X"CD",
		X"EB",X"F7",X"87",X"9F",X"DF",X"F3",X"1F",X"FB",X"FF",X"EF",X"FF",X"F5",X"EF",X"9B",X"6F",X"9E",
		X"89",X"6F",X"B4",X"AE",X"F3",X"AB",X"F5",X"9F",X"5B",X"7B",X"4B",X"BF",X"EF",X"7F",X"EF",X"DF",
		X"FF",X"FC",X"1B",X"FD",X"FD",X"EE",X"48",X"FE",X"DF",X"FA",X"E3",X"17",X"77",X"9D",X"7F",X"D5",
		X"F9",X"DD",X"E4",X"D9",X"FA",X"FC",X"D3",X"CD",X"CF",X"AC",X"EB",X"EF",X"CB",X"8F",X"FD",X"F3",
		X"F7",X"F3",X"C3",X"5F",X"CF",X"DC",X"CA",X"DF",X"DA",X"7F",X"FB",X"9F",X"FF",X"B6",X"AF",X"FF",
		X"FF",X"FA",X"DD",X"FD",X"E3",X"D5",X"B7",X"6E",X"D7",X"9D",X"9C",X"E7",X"4B",X"49",X"FE",X"FF",
		X"5A",X"19",X"20",X"70",X"37",X"30",X"C0",X"66",X"90",X"38",X"20",X"20",X"A0",X"C9",X"80",X"00",
		X"0A",X"84",X"04",X"1A",X"0C",X"B2",X"08",X"18",X"00",X"49",X"E4",X"52",X"5C",X"75",X"0C",X"10",
		X"30",X"28",X"D7",X"12",X"1A",X"40",X"02",X"A2",X"00",X"90",X"88",X"24",X"10",X"E8",X"78",X"C8",
		X"82",X"08",X"20",X"00",X"8C",X"21",X"01",X"48",X"99",X"AA",X"EC",X"31",X"46",X"26",X"70",X"CC",
		X"05",X"80",X"B8",X"63",X"C1",X"18",X"00",X"30",X"32",X"00",X"10",X"00",X"A1",X"23",X"22",X"04",
		X"0A",X"C4",X"67",X"00",X"89",X"15",X"00",X"82",X"62",X"80",X"A2",X"50",X"00",X"3E",X"20",X"A3",
		X"32",X"CC",X"2F",X"3C",X"80",X"10",X"81",X"A5",X"01",X"18",X"03",X"75",X"41",X"51",X"56",X"28",
		X"04",X"A0",X"3D",X"6A",X"21",X"54",X"D5",X"15",X"3A",X"9A",X"A3",X"18",X"19",X"98",X"32",X"B0",
		X"F7",X"FD",X"EF",X"4B",X"DA",X"5F",X"A3",X"DB",X"FF",X"EB",X"FB",X"DF",X"C7",X"EE",X"C7",X"F7",
		X"FD",X"BF",X"C9",X"C7",X"63",X"9F",X"F5",X"FF",X"6F",X"1A",X"FE",X"DE",X"7F",X"5F",X"FD",X"FF",
		X"F9",X"95",X"F9",X"EB",X"81",X"3B",X"5D",X"D3",X"DF",X"A3",X"E7",X"CF",X"BE",X"AF",X"8F",X"7E",
		X"34",X"B5",X"1D",X"CB",X"69",X"6F",X"F1",X"93",X"B4",X"EF",X"E7",X"0D",X"FF",X"3D",X"DB",X"AE",
		X"33",X"BB",X"6F",X"5F",X"05",X"83",X"E7",X"9F",X"FB",X"E6",X"BB",X"D1",X"E5",X"D9",X"D7",X"A7",
		X"BF",X"FB",X"7F",X"ED",X"5F",X"7D",X"13",X"D7",X"CC",X"FB",X"DC",X"97",X"FF",X"BD",X"75",X"7F",
		X"C6",X"16",X"FA",X"C8",X"EE",X"E8",X"A3",X"E7",X"FD",X"A7",X"C6",X"0F",X"E3",X"D4",X"EB",X"04",
		X"D1",X"1B",X"C8",X"17",X"C5",X"9F",X"A7",X"77",X"D8",X"A8",X"DF",X"9E",X"3F",X"DB",X"F2",X"FF",
		X"00",X"D1",X"C1",X"28",X"1C",X"18",X"00",X"92",X"60",X"20",X"01",X"6A",X"20",X"C0",X"23",X"1A",
		X"AB",X"5A",X"D0",X"B2",X"1B",X"10",X"91",X"D1",X"D8",X"02",X"44",X"B0",X"82",X"02",X"6C",X"80",
		X"22",X"BC",X"B2",X"38",X"78",X"01",X"20",X"80",X"02",X"9C",X"34",X"A0",X"80",X"30",X"8D",X"A4",
		X"52",X"10",X"24",X"D4",X"C8",X"80",X"B0",X"06",X"1C",X"00",X"54",X"40",X"E4",X"68",X"04",X"48",
		X"09",X"28",X"01",X"40",X"4A",X"0B",X"EA",X"C0",X"20",X"35",X"80",X"C4",X"13",X"10",X"84",X"9A",
		X"C7",X"82",X"34",X"31",X"95",X"38",X"18",X"2A",X"1C",X"DC",X"92",X"A3",X"98",X"00",X"2C",X"7D",
		X"96",X"A4",X"B0",X"38",X"27",X"A2",X"C1",X"20",X"94",X"AD",X"0B",X"82",X"1C",X"A1",X"08",X"00",
		X"A8",X"81",X"20",X"05",X"20",X"A8",X"A4",X"A8",X"27",X"88",X"02",X"88",X"48",X"CB",X"32",X"80",
		X"9F",X"FC",X"74",X"A8",X"D9",X"F9",X"C9",X"FD",X"FB",X"3F",X"FB",X"E8",X"F5",X"F8",X"B8",X"99",
		X"58",X"F9",X"E8",X"6B",X"D3",X"2B",X"7B",X"DE",X"D9",X"FB",X"30",X"F9",X"16",X"7B",X"F9",X"7D",
		X"F0",X"D9",X"7C",X"FB",X"D9",X"71",X"51",X"BA",X"CD",X"F1",X"FC",X"FB",X"FB",X"F7",X"F9",X"F9",
		X"DA",X"E6",X"F8",X"79",X"44",X"AB",X"99",X"58",X"78",X"F5",X"FD",X"E9",X"F9",X"1A",X"9A",X"F5",
		X"FC",X"F1",X"FB",X"7A",X"77",X"B8",X"51",X"31",X"39",X"9B",X"A9",X"F5",X"70",X"79",X"93",X"FD",
		X"39",X"6B",X"DB",X"F1",X"BA",X"B9",X"D9",X"F6",X"9F",X"FC",X"F9",X"E9",X"F1",X"B8",X"DE",X"F9",
		X"E9",X"3C",X"B9",X"B1",X"79",X"F9",X"71",X"B1",X"F2",X"79",X"FC",X"EF",X"F8",X"69",X"E1",X"31",
		X"ED",X"B8",X"99",X"B0",X"E9",X"F3",X"29",X"FB",X"F8",X"FB",X"71",X"BA",X"F9",X"B8",X"3D",X"19",
		X"06",X"03",X"06",X"C4",X"62",X"2C",X"50",X"86",X"12",X"5C",X"06",X"87",X"07",X"48",X"04",X"60",
		X"46",X"D6",X"9F",X"5C",X"44",X"D7",X"A4",X"C7",X"42",X"23",X"8A",X"06",X"07",X"2C",X"21",X"02",
		X"08",X"42",X"97",X"2F",X"87",X"10",X"45",X"5A",X"8C",X"0C",X"14",X"44",X"04",X"06",X"A7",X"E0",
		X"86",X"A1",X"46",X"26",X"02",X"06",X"47",X"2B",X"83",X"4E",X"E6",X"AC",X"B2",X"84",X"56",X"97",
		X"44",X"04",X"AC",X"46",X"0E",X"42",X"66",X"86",X"06",X"A5",X"46",X"1E",X"46",X"D6",X"86",X"06",
		X"02",X"42",X"16",X"01",X"21",X"06",X"3B",X"46",X"12",X"42",X"D6",X"06",X"A3",X"0F",X"77",X"86",
		X"42",X"16",X"86",X"86",X"0A",X"8B",X"05",X"37",X"2D",X"F2",X"C4",X"0E",X"3E",X"D7",X"87",X"06",
		X"C4",X"46",X"85",X"8E",X"4A",X"B0",X"03",X"E6",X"0F",X"C6",X"86",X"D6",X"42",X"08",X"8F",X"65",
		X"3F",X"ED",X"69",X"F9",X"59",X"AB",X"7D",X"B5",X"70",X"FD",X"FD",X"BB",X"3F",X"35",X"39",X"EB",
		X"7E",X"F8",X"BB",X"7C",X"F1",X"F9",X"FD",X"FD",X"ED",X"F9",X"F9",X"61",X"B9",X"DA",X"D0",X"FF",
		X"6D",X"71",X"3F",X"BB",X"D8",X"F5",X"C9",X"68",X"3D",X"F7",X"40",X"F1",X"F8",X"EC",X"A0",X"A8",
		X"67",X"B9",X"DE",X"7F",X"98",X"3C",X"DE",X"E9",X"79",X"89",X"3B",X"B0",X"E9",X"F9",X"88",X"F9",
		X"F0",X"B7",X"FC",X"E8",X"D8",X"F5",X"B6",X"FD",X"B9",X"F0",X"DC",X"52",X"59",X"B9",X"D9",X"E3",
		X"D5",X"F9",X"11",X"B1",X"F9",X"F5",X"E9",X"F8",X"FC",X"79",X"39",X"FB",X"FD",X"B1",X"A0",X"7F",
		X"39",X"FF",X"B5",X"F8",X"33",X"FB",X"D3",X"F8",X"F9",X"EB",X"E9",X"79",X"BD",X"7B",X"F9",X"A0",
		X"D4",X"B7",X"F8",X"F8",X"19",X"51",X"48",X"7A",X"E1",X"B1",X"DC",X"E8",X"30",X"D9",X"74",X"39",
		X"23",X"0E",X"08",X"94",X"06",X"6C",X"32",X"06",X"86",X"86",X"63",X"A6",X"C7",X"84",X"CD",X"C8",
		X"32",X"0F",X"8D",X"0E",X"41",X"0C",X"66",X"06",X"E6",X"02",X"88",X"46",X"44",X"77",X"8E",X"A4",
		X"9E",X"46",X"5E",X"0A",X"6E",X"87",X"82",X"88",X"02",X"1C",X"8D",X"9D",X"02",X"97",X"6A",X"66",
		X"F3",X"A4",X"03",X"81",X"46",X"9A",X"1E",X"34",X"05",X"BD",X"43",X"02",X"03",X"8A",X"A7",X"CC",
		X"02",X"5C",X"2E",X"0A",X"07",X"57",X"14",X"C4",X"08",X"0E",X"26",X"A8",X"6F",X"C6",X"03",X"0E",
		X"92",X"0E",X"A1",X"26",X"37",X"8A",X"86",X"0E",X"02",X"66",X"C1",X"85",X"42",X"52",X"8C",X"66",
		X"86",X"86",X"46",X"0E",X"86",X"E7",X"9E",X"1E",X"C6",X"0B",X"08",X"C6",X"46",X"C6",X"0C",X"44",
		X"40",X"84",X"17",X"85",X"46",X"67",X"46",X"8C",X"46",X"67",X"8D",X"95",X"4E",X"C5",X"40",X"06",
		X"7B",X"BF",X"FD",X"77",X"DF",X"FF",X"27",X"72",X"FE",X"4E",X"7F",X"DB",X"9B",X"67",X"1F",X"F7",
		X"DF",X"BD",X"AF",X"FE",X"F5",X"F5",X"CC",X"36",X"F3",X"FD",X"53",X"6D",X"EF",X"D8",X"BE",X"D5",
		X"BF",X"AB",X"1D",X"F2",X"CB",X"BC",X"FC",X"BD",X"6D",X"03",X"FF",X"BF",X"93",X"FF",X"AF",X"FB",
		X"A3",X"4F",X"C6",X"7D",X"DB",X"79",X"F5",X"7B",X"7D",X"EB",X"FD",X"EB",X"CD",X"A1",X"F1",X"0E",
		X"D2",X"D5",X"AE",X"EB",X"FC",X"EE",X"8D",X"A9",X"FF",X"DF",X"1F",X"F4",X"E2",X"DD",X"36",X"F7",
		X"7F",X"13",X"7D",X"AD",X"F6",X"0E",X"DF",X"CF",X"F7",X"64",X"C3",X"7B",X"F5",X"BE",X"EB",X"39",
		X"AE",X"9F",X"FE",X"EB",X"FD",X"9B",X"56",X"85",X"EB",X"7F",X"59",X"1F",X"3E",X"62",X"C0",X"5F",
		X"7B",X"ED",X"DF",X"F6",X"65",X"79",X"2B",X"FE",X"E7",X"CF",X"7F",X"ED",X"1D",X"FF",X"AF",X"57",
		X"88",X"64",X"4B",X"22",X"C0",X"10",X"A4",X"10",X"19",X"22",X"7A",X"AE",X"0A",X"26",X"A0",X"B4",
		X"18",X"4D",X"B8",X"81",X"29",X"88",X"31",X"70",X"A0",X"F6",X"00",X"14",X"10",X"F0",X"10",X"70",
		X"86",X"80",X"12",X"3E",X"52",X"02",X"B6",X"C9",X"08",X"C0",X"A0",X"70",X"52",X"D8",X"00",X"20",
		X"12",X"08",X"50",X"0D",X"02",X"20",X"8C",X"F3",X"28",X"80",X"90",X"80",X"90",X"16",X"78",X"92",
		X"20",X"22",X"24",X"58",X"2A",X"4D",X"2D",X"85",X"10",X"30",X"01",X"39",X"00",X"00",X"09",X"33",
		X"3F",X"99",X"B0",X"80",X"42",X"72",X"42",X"00",X"11",X"22",X"23",X"A1",X"04",X"08",X"92",X"A3",
		X"B1",X"15",X"10",X"5A",X"A8",X"0A",X"40",X"92",X"A5",X"C4",X"92",X"1B",X"20",X"A0",X"00",X"30",
		X"42",X"59",X"F2",X"1C",X"0C",X"D0",X"C6",X"CA",X"B0",X"AA",X"1A",X"19",X"5A",X"84",X"BF",X"3D",
		X"7D",X"3F",X"EF",X"4D",X"9D",X"99",X"67",X"5B",X"67",X"EB",X"7D",X"D9",X"4D",X"FF",X"D5",X"3D",
		X"9F",X"B4",X"9F",X"C7",X"1D",X"49",X"7D",X"B6",X"A7",X"3E",X"CF",X"AB",X"45",X"EF",X"DD",X"EF",
		X"FF",X"7D",X"C7",X"BB",X"63",X"E7",X"F3",X"BF",X"6F",X"F6",X"EF",X"DF",X"DB",X"DB",X"A7",X"DF",
		X"FB",X"BE",X"AD",X"4B",X"1B",X"5A",X"FF",X"DF",X"3F",X"E7",X"DF",X"87",X"BF",X"ED",X"FD",X"F7",
		X"CF",X"D5",X"FF",X"EB",X"B3",X"F1",X"FF",X"83",X"E5",X"D9",X"DE",X"EC",X"EB",X"CD",X"FF",X"33",
		X"D7",X"CD",X"79",X"B7",X"F7",X"DE",X"CE",X"EF",X"6B",X"A7",X"BD",X"FE",X"FF",X"E3",X"F6",X"9F",
		X"B3",X"FC",X"6B",X"D3",X"79",X"F2",X"D9",X"CF",X"AB",X"8F",X"E7",X"BB",X"F9",X"EE",X"BF",X"B5",
		X"E7",X"8A",X"B3",X"FB",X"3E",X"6F",X"6F",X"6C",X"56",X"EF",X"EB",X"CB",X"D3",X"81",X"F5",X"B1",
		X"60",X"6B",X"4A",X"98",X"10",X"A8",X"E9",X"28",X"98",X"1D",X"98",X"A0",X"08",X"BC",X"1A",X"8D",
		X"86",X"38",X"5D",X"01",X"60",X"A8",X"A2",X"16",X"02",X"64",X"00",X"00",X"A7",X"91",X"03",X"00",
		X"70",X"3A",X"00",X"30",X"18",X"25",X"02",X"90",X"50",X"06",X"80",X"88",X"52",X"80",X"10",X"00",
		X"E8",X"ED",X"A2",X"12",X"00",X"23",X"A4",X"0B",X"84",X"C4",X"80",X"60",X"20",X"82",X"20",X"0C",
		X"88",X"CE",X"2B",X"3E",X"80",X"B7",X"01",X"44",X"10",X"22",X"90",X"03",X"23",X"88",X"11",X"03",
		X"81",X"42",X"00",X"39",X"18",X"DA",X"5A",X"36",X"78",X"80",X"48",X"00",X"84",X"0E",X"20",X"00",
		X"16",X"82",X"66",X"81",X"30",X"14",X"08",X"10",X"84",X"01",X"51",X"A8",X"09",X"04",X"B3",X"00",
		X"4C",X"41",X"40",X"20",X"16",X"C0",X"5A",X"D0",X"02",X"92",X"02",X"19",X"48",X"02",X"80",X"0C",
		X"F9",X"99",X"D5",X"79",X"F0",X"79",X"E8",X"B3",X"97",X"6B",X"39",X"FF",X"FF",X"F9",X"B9",X"3A",
		X"F1",X"79",X"B3",X"A9",X"A0",X"E9",X"7A",X"B1",X"95",X"30",X"A9",X"9D",X"F9",X"30",X"FD",X"72",
		X"5C",X"FC",X"B1",X"F2",X"B9",X"F9",X"59",X"C9",X"73",X"BB",X"3A",X"FA",X"DB",X"98",X"F2",X"D5",
		X"51",X"E8",X"7D",X"FB",X"F9",X"5D",X"F9",X"FF",X"32",X"75",X"FE",X"71",X"B1",X"68",X"F4",X"B9",
		X"FF",X"F9",X"FD",X"B9",X"B1",X"BA",X"59",X"B9",X"BE",X"E8",X"B8",X"F1",X"F7",X"B8",X"F1",X"49",
		X"6D",X"F1",X"9E",X"35",X"E1",X"78",X"E0",X"F9",X"B9",X"F9",X"B0",X"BC",X"D4",X"61",X"63",X"59",
		X"F0",X"87",X"D9",X"B9",X"58",X"72",X"D8",X"EB",X"8A",X"F1",X"35",X"33",X"B5",X"79",X"79",X"FD",
		X"D0",X"6D",X"39",X"F9",X"FF",X"F9",X"54",X"F9",X"7B",X"F9",X"FB",X"E9",X"AD",X"F8",X"79",X"F0",
		X"77",X"07",X"30",X"5D",X"8F",X"C7",X"A5",X"07",X"04",X"A7",X"8D",X"44",X"86",X"C6",X"A0",X"45",
		X"18",X"07",X"D4",X"7F",X"1F",X"03",X"04",X"05",X"07",X"4E",X"66",X"05",X"6E",X"06",X"06",X"4E",
		X"07",X"2E",X"47",X"46",X"06",X"26",X"06",X"46",X"76",X"06",X"02",X"01",X"97",X"D3",X"C6",X"87",
		X"A2",X"87",X"00",X"2A",X"37",X"32",X"A4",X"87",X"66",X"76",X"41",X"1E",X"7E",X"63",X"14",X"89",
		X"BE",X"06",X"0F",X"53",X"CA",X"8E",X"06",X"02",X"46",X"26",X"07",X"87",X"4F",X"44",X"04",X"0A",
		X"96",X"EC",X"10",X"4E",X"0A",X"0C",X"A6",X"A6",X"0E",X"4F",X"C7",X"86",X"02",X"8E",X"06",X"AC",
		X"D6",X"00",X"9B",X"23",X"45",X"2E",X"0C",X"67",X"07",X"22",X"83",X"43",X"62",X"C7",X"0C",X"0E",
		X"87",X"06",X"14",X"66",X"BD",X"16",X"E7",X"0E",X"8F",X"06",X"64",X"0F",X"86",X"0F",X"06",X"86",
		X"FF",X"D1",X"99",X"78",X"5D",X"69",X"F9",X"71",X"DB",X"71",X"3B",X"9B",X"ED",X"7D",X"F8",X"79",
		X"9C",X"F9",X"DB",X"F6",X"EB",X"41",X"77",X"43",X"D9",X"59",X"FB",X"33",X"FF",X"F5",X"B9",X"39",
		X"A8",X"C9",X"31",X"A3",X"5D",X"B4",X"71",X"69",X"78",X"7B",X"BE",X"FD",X"78",X"BD",X"73",X"39",
		X"F4",X"F9",X"BC",X"B1",X"F9",X"64",X"22",X"3C",X"9B",X"5A",X"B9",X"74",X"5C",X"99",X"6B",X"F9",
		X"7F",X"90",X"F9",X"78",X"F8",X"B9",X"3B",X"B1",X"39",X"F9",X"6F",X"F8",X"DE",X"FF",X"B1",X"D8",
		X"A9",X"96",X"E8",X"DA",X"F5",X"7A",X"A4",X"39",X"B9",X"F9",X"DD",X"4B",X"DB",X"FA",X"D8",X"7B",
		X"F5",X"C1",X"B9",X"FC",X"D8",X"79",X"9E",X"90",X"E9",X"50",X"34",X"99",X"A1",X"59",X"FD",X"69",
		X"A1",X"FB",X"1B",X"B8",X"77",X"B9",X"14",X"1B",X"27",X"48",X"FF",X"08",X"F8",X"EB",X"B0",X"F8",
		X"B9",X"66",X"03",X"46",X"0F",X"47",X"75",X"C6",X"47",X"02",X"07",X"02",X"0C",X"24",X"2F",X"02",
		X"8C",X"43",X"82",X"D5",X"2A",X"0F",X"9C",X"02",X"28",X"0C",X"03",X"8D",X"36",X"04",X"23",X"86",
		X"42",X"D2",X"A4",X"46",X"CF",X"8C",X"76",X"96",X"C7",X"05",X"86",X"80",X"5B",X"66",X"46",X"0E",
		X"16",X"4C",X"4E",X"46",X"52",X"07",X"A7",X"C5",X"03",X"0F",X"44",X"A3",X"0E",X"46",X"46",X"64",
		X"0E",X"27",X"26",X"0B",X"07",X"4E",X"82",X"C6",X"07",X"06",X"D6",X"46",X"4E",X"C2",X"A4",X"06",
		X"07",X"47",X"17",X"87",X"58",X"15",X"57",X"07",X"44",X"97",X"0C",X"42",X"04",X"86",X"06",X"57",
		X"03",X"44",X"06",X"46",X"D2",X"0E",X"0F",X"43",X"47",X"56",X"AC",X"4C",X"06",X"06",X"37",X"86",
		X"06",X"56",X"B4",X"07",X"6E",X"28",X"54",X"07",X"C6",X"86",X"07",X"83",X"1E",X"88",X"46",X"AD");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
