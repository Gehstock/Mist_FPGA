library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity wacko_sp_bits_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of wacko_sp_bits_1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"09",
		X"00",X"00",X"99",X"99",X"00",X"90",X"A9",X"93",X"00",X"99",X"9F",X"93",X"00",X"33",X"9F",X"9B",
		X"00",X"93",X"FF",X"9B",X"00",X"93",X"F9",X"93",X"00",X"B9",X"99",X"9B",X"00",X"B9",X"33",X"9B",
		X"00",X"39",X"39",X"39",X"00",X"93",X"33",X"39",X"00",X"99",X"93",X"33",X"00",X"09",X"99",X"33",
		X"00",X"00",X"99",X"33",X"00",X"90",X"33",X"39",X"00",X"99",X"99",X"99",X"00",X"39",X"B9",X"90",
		X"00",X"33",X"99",X"99",X"00",X"93",X"9B",X"39",X"90",X"99",X"93",X"33",X"09",X"00",X"33",X"33",
		X"00",X"00",X"33",X"99",X"00",X"00",X"33",X"99",X"00",X"99",X"93",X"33",X"09",X"33",X"93",X"33",
		X"00",X"33",X"33",X"33",X"00",X"99",X"33",X"33",X"00",X"99",X"39",X"33",X"09",X"99",X"99",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"22",X"99",X"00",X"99",X"99",X"9D",
		X"99",X"99",X"99",X"DD",X"9D",X"22",X"99",X"DD",X"99",X"DD",X"99",X"DD",X"49",X"9D",X"22",X"DD",
		X"9D",X"9D",X"22",X"9D",X"92",X"D2",X"99",X"9D",X"99",X"22",X"99",X"99",X"00",X"99",X"95",X"22",
		X"00",X"59",X"95",X"29",X"00",X"99",X"99",X"22",X"00",X"99",X"99",X"92",X"00",X"99",X"59",X"22",
		X"00",X"99",X"99",X"22",X"00",X"99",X"29",X"29",X"00",X"D2",X"22",X"99",X"00",X"22",X"99",X"22",
		X"00",X"22",X"99",X"22",X"00",X"29",X"99",X"22",X"00",X"99",X"9A",X"22",X"00",X"29",X"99",X"29",
		X"00",X"22",X"99",X"2A",X"00",X"99",X"22",X"29",X"00",X"9A",X"22",X"29",X"00",X"99",X"22",X"22",
		X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"99",X"99",X"00",X"00",X"22",X"99",X"00",X"99",X"99",X"9D",X"99",X"99",X"99",X"DD",
		X"9D",X"22",X"99",X"DD",X"99",X"DD",X"99",X"DD",X"99",X"9D",X"22",X"DD",X"9D",X"9D",X"22",X"9D",
		X"92",X"D2",X"99",X"9D",X"99",X"22",X"99",X"99",X"00",X"99",X"95",X"22",X"09",X"59",X"95",X"29",
		X"09",X"99",X"99",X"22",X"09",X"22",X"22",X"92",X"00",X"29",X"22",X"22",X"00",X"22",X"92",X"22",
		X"00",X"99",X"22",X"29",X"00",X"D9",X"22",X"99",X"00",X"D9",X"99",X"22",X"00",X"29",X"DD",X"22",
		X"00",X"29",X"99",X"22",X"00",X"29",X"9A",X"22",X"00",X"29",X"99",X"29",X"00",X"22",X"99",X"2A",
		X"00",X"99",X"22",X"29",X"00",X"9A",X"22",X"29",X"00",X"99",X"22",X"22",X"00",X"99",X"22",X"22",
		X"00",X"99",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",
		X"00",X"22",X"22",X"22",X"00",X"22",X"99",X"22",X"00",X"22",X"9A",X"22",X"00",X"22",X"99",X"22",
		X"00",X"22",X"99",X"99",X"99",X"92",X"22",X"A9",X"92",X"99",X"22",X"99",X"92",X"22",X"22",X"99",
		X"92",X"99",X"99",X"22",X"92",X"00",X"91",X"29",X"92",X"00",X"92",X"29",X"99",X"99",X"99",X"29",
		X"09",X"29",X"09",X"29",X"00",X"29",X"09",X"29",X"00",X"99",X"09",X"19",X"00",X"90",X"09",X"99",
		X"00",X"90",X"00",X"90",X"00",X"90",X"00",X"90",X"99",X"00",X"00",X"90",X"92",X"00",X"00",X"90",
		X"99",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"99",
		X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"99",X"99",
		X"00",X"22",X"22",X"99",X"00",X"22",X"22",X"A9",X"00",X"22",X"22",X"99",X"00",X"22",X"29",X"92",
		X"00",X"22",X"99",X"29",X"00",X"22",X"92",X"29",X"00",X"22",X"22",X"99",X"00",X"22",X"99",X"99",
		X"00",X"92",X"9A",X"22",X"00",X"99",X"99",X"22",X"00",X"2D",X"29",X"22",X"00",X"22",X"22",X"22",
		X"00",X"22",X"22",X"29",X"00",X"22",X"99",X"99",X"00",X"22",X"90",X"99",X"00",X"29",X"00",X"92",
		X"00",X"99",X"00",X"22",X"00",X"90",X"00",X"22",X"00",X"90",X"00",X"22",X"00",X"90",X"00",X"22",
		X"00",X"99",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"D2",X"00",X"22",
		X"00",X"DD",X"00",X"22",X"00",X"2D",X"00",X"22",X"99",X"22",X"00",X"22",X"92",X"2D",X"00",X"99",
		X"92",X"2D",X"00",X"00",X"92",X"22",X"00",X"00",X"99",X"29",X"00",X"00",X"09",X"99",X"00",X"00",
		X"00",X"09",X"09",X"09",X"00",X"09",X"99",X"90",X"00",X"09",X"99",X"99",X"00",X"09",X"99",X"99",
		X"00",X"09",X"44",X"9B",X"99",X"09",X"99",X"BB",X"9B",X"9B",X"BB",X"BB",X"9B",X"B9",X"BB",X"BB",
		X"99",X"B9",X"BB",X"BB",X"99",X"B9",X"99",X"BB",X"09",X"BB",X"99",X"BB",X"09",X"99",X"99",X"BB",
		X"00",X"95",X"99",X"BB",X"00",X"95",X"99",X"BB",X"00",X"4F",X"99",X"BB",X"00",X"99",X"BB",X"BB",
		X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"B9",X"44",X"BB",X"99",X"90",X"04",X"99",X"BB",X"90",
		X"00",X"00",X"BB",X"90",X"00",X"00",X"BB",X"90",X"00",X"00",X"BB",X"99",X"00",X"09",X"99",X"BB",
		X"00",X"99",X"77",X"BB",X"00",X"9B",X"77",X"BB",X"00",X"BB",X"77",X"BB",X"00",X"B9",X"99",X"BB",
		X"00",X"99",X"11",X"BB",X"00",X"99",X"77",X"BB",X"00",X"19",X"97",X"BB",X"00",X"71",X"11",X"BB",
		X"00",X"00",X"00",X"00",X"00",X"09",X"09",X"00",X"00",X"09",X"99",X"90",X"00",X"09",X"99",X"99",
		X"00",X"09",X"99",X"99",X"00",X"09",X"43",X"9B",X"99",X"09",X"99",X"BB",X"9B",X"9B",X"BB",X"BB",
		X"9B",X"B9",X"BB",X"BB",X"94",X"B9",X"BB",X"BB",X"99",X"B9",X"BB",X"BB",X"09",X"BB",X"99",X"BB",
		X"09",X"BB",X"99",X"BB",X"00",X"99",X"99",X"BB",X"00",X"95",X"99",X"BB",X"00",X"4F",X"99",X"BB",
		X"00",X"49",X"99",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"B9",X"00",X"BB",X"99",X"90",
		X"00",X"99",X"BB",X"90",X"00",X"00",X"BB",X"90",X"00",X"00",X"BB",X"90",X"00",X"00",X"BB",X"99",
		X"00",X"09",X"99",X"B9",X"00",X"99",X"77",X"B9",X"00",X"9B",X"77",X"BB",X"00",X"BB",X"77",X"BB",
		X"00",X"B9",X"99",X"BB",X"00",X"99",X"11",X"BB",X"00",X"99",X"77",X"BB",X"00",X"19",X"97",X"BB",
		X"00",X"77",X"77",X"BB",X"00",X"99",X"77",X"BB",X"00",X"11",X"17",X"BB",X"00",X"77",X"77",X"BB",
		X"00",X"77",X"79",X"BB",X"00",X"99",X"79",X"BB",X"00",X"11",X"99",X"B9",X"00",X"77",X"9B",X"B9",
		X"00",X"77",X"BB",X"B9",X"00",X"99",X"B9",X"B9",X"00",X"11",X"99",X"B9",X"00",X"77",X"1B",X"BB",
		X"00",X"77",X"99",X"BB",X"00",X"77",X"BB",X"9B",X"00",X"99",X"BB",X"9B",X"00",X"11",X"BB",X"99",
		X"00",X"77",X"BB",X"19",X"09",X"77",X"BB",X"99",X"09",X"99",X"9B",X"BB",X"09",X"B9",X"99",X"BB",
		X"09",X"99",X"9B",X"99",X"09",X"90",X"9B",X"99",X"00",X"B9",X"9B",X"90",X"00",X"BB",X"9B",X"99",
		X"00",X"BB",X"99",X"9B",X"00",X"BB",X"09",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"BB",
		X"09",X"99",X"00",X"99",X"99",X"90",X"00",X"09",X"9B",X"90",X"00",X"9B",X"99",X"00",X"00",X"99",
		X"00",X"71",X"11",X"BB",X"00",X"79",X"77",X"BB",X"00",X"99",X"77",X"BB",X"00",X"BB",X"99",X"BB",
		X"00",X"BB",X"BB",X"BB",X"00",X"99",X"BB",X"B9",X"00",X"99",X"BB",X"99",X"00",X"19",X"BB",X"00",
		X"00",X"79",X"99",X"00",X"00",X"77",X"BB",X"00",X"00",X"99",X"BB",X"00",X"00",X"11",X"BB",X"00",
		X"00",X"77",X"BB",X"00",X"00",X"77",X"BB",X"09",X"00",X"77",X"BB",X"99",X"00",X"99",X"BB",X"9B",
		X"00",X"11",X"BB",X"BB",X"00",X"77",X"BB",X"BB",X"00",X"77",X"BB",X"BB",X"00",X"99",X"9B",X"BB",
		X"00",X"09",X"99",X"BB",X"00",X"00",X"BB",X"99",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"99",X"BB",X"00",X"00",X"9B",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"99",X"BB",X"00",
		X"00",X"9B",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"99",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"66",X"00",
		X"00",X"99",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"90",
		X"99",X"99",X"66",X"99",X"9E",X"9E",X"66",X"69",X"9E",X"E9",X"66",X"66",X"9E",X"E9",X"99",X"99",
		X"99",X"E9",X"9C",X"66",X"09",X"EE",X"CC",X"66",X"09",X"EE",X"CC",X"66",X"99",X"EE",X"CC",X"66",
		X"99",X"E9",X"99",X"66",X"99",X"99",X"99",X"66",X"99",X"99",X"CC",X"66",X"99",X"99",X"9C",X"66",
		X"99",X"49",X"9C",X"66",X"99",X"99",X"9C",X"66",X"9C",X"CC",X"CC",X"66",X"9C",X"C9",X"CC",X"66",
		X"9C",X"99",X"CC",X"66",X"99",X"99",X"CC",X"66",X"09",X"99",X"C9",X"66",X"09",X"99",X"99",X"66",
		X"09",X"F9",X"9D",X"66",X"00",X"99",X"DD",X"66",X"00",X"CC",X"D6",X"66",X"00",X"99",X"66",X"66",
		X"00",X"99",X"99",X"00",X"00",X"96",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"00",
		X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"90",X"00",X"99",X"66",X"99",X"09",X"9E",X"66",X"69",
		X"09",X"E9",X"66",X"66",X"09",X"E9",X"99",X"99",X"09",X"E9",X"9C",X"66",X"00",X"EE",X"CC",X"66",
		X"09",X"EE",X"CC",X"66",X"99",X"EE",X"CC",X"66",X"9C",X"E9",X"99",X"66",X"99",X"99",X"99",X"66",
		X"99",X"99",X"CC",X"66",X"99",X"99",X"9C",X"66",X"99",X"49",X"9C",X"66",X"99",X"99",X"9C",X"66",
		X"9C",X"CC",X"CC",X"66",X"9C",X"C9",X"CC",X"66",X"9C",X"99",X"CC",X"66",X"99",X"99",X"CC",X"66",
		X"09",X"99",X"C9",X"66",X"09",X"99",X"99",X"66",X"09",X"99",X"9D",X"66",X"00",X"CC",X"DD",X"66",
		X"00",X"99",X"D6",X"66",X"00",X"DD",X"66",X"66",X"00",X"66",X"66",X"66",X"00",X"66",X"66",X"66",
		X"00",X"66",X"66",X"66",X"00",X"66",X"66",X"66",X"00",X"66",X"66",X"66",X"00",X"66",X"66",X"66",
		X"00",X"66",X"66",X"66",X"00",X"66",X"66",X"66",X"00",X"99",X"66",X"66",X"00",X"55",X"99",X"66",
		X"00",X"99",X"9D",X"66",X"00",X"99",X"DD",X"66",X"00",X"99",X"DD",X"66",X"00",X"55",X"D9",X"66",
		X"00",X"99",X"99",X"66",X"00",X"66",X"66",X"66",X"00",X"66",X"66",X"66",X"00",X"66",X"66",X"66",
		X"00",X"D6",X"66",X"66",X"00",X"DD",X"99",X"66",X"99",X"66",X"99",X"66",X"99",X"66",X"9D",X"66",
		X"99",X"66",X"DD",X"66",X"97",X"66",X"D6",X"99",X"97",X"66",X"D6",X"CC",X"97",X"66",X"96",X"CC",
		X"97",X"69",X"96",X"C9",X"97",X"99",X"99",X"CC",X"97",X"00",X"97",X"CC",X"99",X"00",X"97",X"9C",
		X"99",X"00",X"99",X"9C",X"09",X"00",X"79",X"99",X"09",X"00",X"77",X"9C",X"09",X"00",X"99",X"99",
		X"00",X"66",X"66",X"66",X"00",X"66",X"66",X"66",X"00",X"66",X"66",X"66",X"00",X"66",X"66",X"66",
		X"00",X"99",X"66",X"66",X"00",X"55",X"99",X"66",X"00",X"99",X"9D",X"66",X"00",X"99",X"DD",X"66",
		X"00",X"99",X"DD",X"66",X"00",X"55",X"D9",X"66",X"00",X"99",X"99",X"66",X"00",X"66",X"66",X"66",
		X"00",X"66",X"66",X"66",X"00",X"66",X"66",X"66",X"00",X"66",X"66",X"66",X"00",X"66",X"69",X"66",
		X"00",X"99",X"69",X"66",X"00",X"DD",X"69",X"66",X"00",X"6D",X"69",X"66",X"09",X"66",X"69",X"99",
		X"09",X"66",X"69",X"CC",X"09",X"66",X"69",X"CC",X"09",X"99",X"69",X"CC",X"00",X"77",X"69",X"CC",
		X"00",X"99",X"99",X"CC",X"00",X"99",X"79",X"CC",X"00",X"97",X"99",X"CC",X"00",X"77",X"99",X"9C",
		X"00",X"77",X"99",X"9C",X"00",X"77",X"00",X"9C",X"00",X"99",X"00",X"99",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"B9",X"00",X"00",X"00",X"9E",X"00",
		X"00",X"00",X"9E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9E",X"00",
		X"00",X"00",X"9E",X"00",X"00",X"00",X"99",X"90",X"00",X"09",X"9E",X"99",X"00",X"09",X"99",X"E9",
		X"00",X"09",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"9E",X"99",X"E9",X"00",X"9E",X"99",X"E9",
		X"00",X"EE",X"9E",X"99",X"00",X"99",X"99",X"B9",X"00",X"EE",X"97",X"B9",X"00",X"9E",X"99",X"99",
		X"00",X"99",X"99",X"B9",X"00",X"E9",X"99",X"99",X"00",X"9B",X"E9",X"EE",X"00",X"9B",X"99",X"E9",
		X"00",X"9E",X"9E",X"E9",X"00",X"9E",X"9E",X"E9",X"00",X"9E",X"9E",X"99",X"00",X"9B",X"99",X"B9",
		X"00",X"9B",X"99",X"E9",X"09",X"99",X"E9",X"EB",X"09",X"E9",X"E9",X"EB",X"09",X"49",X"E9",X"B9",
		X"00",X"00",X"B9",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"99",X"90",
		X"00",X"09",X"9E",X"99",X"00",X"09",X"99",X"E9",X"00",X"09",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"9E",X"99",X"E9",X"00",X"9E",X"99",X"E9",X"00",X"E9",X"9E",X"99",X"00",X"99",X"99",X"B9",
		X"00",X"E9",X"97",X"B9",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"B9",X"00",X"E9",X"99",X"99",
		X"00",X"9B",X"99",X"EE",X"00",X"9B",X"99",X"E9",X"00",X"9E",X"99",X"E9",X"00",X"9E",X"9E",X"E9",
		X"00",X"9E",X"9E",X"99",X"00",X"9B",X"99",X"B9",X"00",X"9B",X"9E",X"E9",X"09",X"99",X"EE",X"EB",
		X"09",X"E9",X"EE",X"EB",X"09",X"49",X"9E",X"B9",X"00",X"9E",X"99",X"EE",X"00",X"9E",X"E9",X"EE",
		X"09",X"99",X"99",X"EE",X"09",X"9E",X"9E",X"EE",X"00",X"9E",X"9E",X"9E",X"09",X"9E",X"99",X"99",
		X"09",X"99",X"E9",X"99",X"09",X"EB",X"E9",X"9E",X"09",X"BE",X"99",X"99",X"09",X"B9",X"9E",X"EE",
		X"00",X"99",X"9E",X"99",X"00",X"E9",X"E9",X"99",X"00",X"E9",X"49",X"99",X"00",X"E9",X"E9",X"E9",
		X"00",X"E9",X"9E",X"9E",X"00",X"9E",X"9E",X"99",X"00",X"E9",X"9E",X"EE",X"00",X"E9",X"9E",X"99",
		X"00",X"99",X"9E",X"99",X"00",X"B9",X"99",X"00",X"00",X"B9",X"EE",X"00",X"00",X"E9",X"9E",X"00",
		X"00",X"EE",X"9E",X"90",X"00",X"EE",X"9E",X"90",X"00",X"9E",X"99",X"90",X"00",X"99",X"9E",X"99",
		X"00",X"E9",X"9E",X"B9",X"00",X"E9",X"9E",X"99",X"00",X"E9",X"99",X"EE",X"09",X"99",X"E9",X"9E",
		X"09",X"EE",X"EE",X"99",X"09",X"99",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"9E",X"E9",X"99",X"09",X"9E",X"E9",X"EE",X"09",X"99",X"99",X"EE",X"09",X"9E",X"99",X"E9",
		X"00",X"9E",X"99",X"99",X"00",X"9E",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"EB",X"E9",X"99",
		X"00",X"B9",X"99",X"99",X"00",X"B9",X"9E",X"E9",X"00",X"99",X"9E",X"99",X"00",X"E9",X"EE",X"99",
		X"00",X"E9",X"4E",X"90",X"00",X"E9",X"99",X"90",X"00",X"EB",X"E9",X"99",X"09",X"BB",X"E9",X"E9",
		X"09",X"B9",X"99",X"EE",X"99",X"99",X"EE",X"99",X"9E",X"99",X"EE",X"E9",X"99",X"90",X"99",X"E9",
		X"99",X"00",X"00",X"9B",X"9E",X"00",X"00",X"9E",X"99",X"99",X"00",X"99",X"09",X"E9",X"00",X"E9",
		X"00",X"EE",X"00",X"E9",X"09",X"9E",X"00",X"E9",X"09",X"9E",X"00",X"E9",X"99",X"9E",X"00",X"99",
		X"9E",X"99",X"00",X"E9",X"99",X"B9",X"00",X"99",X"9E",X"B9",X"00",X"9B",X"99",X"99",X"00",X"99",
		X"99",X"00",X"09",X"00",X"9A",X"00",X"99",X"00",X"99",X"00",X"79",X"99",X"09",X"00",X"79",X"77",
		X"09",X"99",X"77",X"77",X"00",X"97",X"79",X"77",X"00",X"97",X"79",X"97",X"00",X"97",X"97",X"99",
		X"00",X"97",X"97",X"44",X"00",X"77",X"99",X"99",X"00",X"79",X"49",X"77",X"00",X"99",X"04",X"77",
		X"09",X"F9",X"00",X"97",X"09",X"99",X"00",X"99",X"09",X"99",X"00",X"E9",X"09",X"99",X"40",X"E9",
		X"09",X"97",X"90",X"79",X"00",X"97",X"94",X"79",X"00",X"97",X"99",X"79",X"00",X"79",X"79",X"79",
		X"00",X"99",X"77",X"79",X"00",X"90",X"77",X"79",X"00",X"09",X"77",X"79",X"00",X"99",X"77",X"79",
		X"00",X"97",X"77",X"79",X"00",X"77",X"77",X"79",X"00",X"77",X"77",X"79",X"00",X"77",X"77",X"99",
		X"00",X"99",X"97",X"77",X"00",X"91",X"99",X"77",X"00",X"91",X"99",X"77",X"00",X"99",X"11",X"77",
		X"00",X"00",X"00",X"99",X"99",X"00",X"99",X"99",X"9A",X"00",X"77",X"99",X"9A",X"00",X"79",X"99",
		X"9A",X"00",X"79",X"77",X"9A",X"90",X"77",X"97",X"99",X"99",X"77",X"99",X"09",X"79",X"99",X"99",
		X"09",X"77",X"97",X"99",X"09",X"77",X"99",X"99",X"09",X"77",X"00",X"77",X"09",X"99",X"00",X"79",
		X"09",X"99",X"00",X"79",X"99",X"99",X"00",X"79",X"97",X"97",X"00",X"79",X"97",X"77",X"00",X"79",
		X"97",X"77",X"00",X"79",X"97",X"79",X"00",X"79",X"97",X"99",X"00",X"79",X"99",X"99",X"90",X"79",
		X"00",X"09",X"90",X"79",X"00",X"09",X"90",X"79",X"00",X"99",X"99",X"79",X"00",X"97",X"79",X"79",
		X"00",X"97",X"79",X"79",X"00",X"97",X"77",X"79",X"00",X"97",X"77",X"79",X"00",X"77",X"77",X"99",
		X"00",X"99",X"97",X"77",X"00",X"91",X"99",X"77",X"00",X"91",X"99",X"77",X"00",X"99",X"11",X"77",
		X"00",X"49",X"99",X"77",X"00",X"99",X"11",X"77",X"00",X"91",X"11",X"77",X"00",X"99",X"99",X"77",
		X"00",X"94",X"49",X"77",X"00",X"94",X"49",X"77",X"00",X"19",X"44",X"77",X"00",X"19",X"99",X"77",
		X"00",X"99",X"11",X"77",X"00",X"91",X"11",X"77",X"00",X"91",X"11",X"77",X"00",X"99",X"99",X"77",
		X"00",X"49",X"49",X"77",X"00",X"99",X"49",X"77",X"00",X"99",X"49",X"77",X"00",X"99",X"99",X"77",
		X"00",X"94",X"97",X"77",X"00",X"94",X"97",X"99",X"00",X"94",X"97",X"00",X"00",X"99",X"77",X"00",
		X"00",X"91",X"77",X"00",X"00",X"91",X"77",X"00",X"00",X"99",X"77",X"00",X"00",X"11",X"77",X"00",
		X"00",X"99",X"77",X"00",X"00",X"11",X"77",X"90",X"00",X"11",X"77",X"99",X"00",X"99",X"77",X"77",
		X"00",X"94",X"99",X"77",X"00",X"79",X"19",X"77",X"00",X"79",X"91",X"77",X"00",X"99",X"99",X"99",
		X"00",X"49",X"99",X"77",X"00",X"99",X"11",X"77",X"00",X"91",X"11",X"77",X"00",X"99",X"99",X"77",
		X"00",X"94",X"49",X"77",X"09",X"94",X"49",X"77",X"09",X"19",X"44",X"77",X"09",X"19",X"99",X"77",
		X"09",X"99",X"11",X"77",X"00",X"91",X"11",X"77",X"00",X"91",X"11",X"77",X"00",X"99",X"99",X"97",
		X"00",X"49",X"49",X"97",X"00",X"99",X"49",X"99",X"00",X"99",X"49",X"00",X"00",X"99",X"99",X"00",
		X"00",X"94",X"97",X"00",X"00",X"94",X"97",X"00",X"00",X"94",X"97",X"00",X"00",X"99",X"77",X"00",
		X"00",X"91",X"77",X"00",X"00",X"91",X"77",X"99",X"00",X"99",X"77",X"97",X"00",X"11",X"77",X"77",
		X"00",X"99",X"77",X"77",X"00",X"11",X"77",X"77",X"00",X"11",X"77",X"77",X"00",X"99",X"77",X"79",
		X"00",X"94",X"99",X"99",X"00",X"79",X"19",X"90",X"00",X"99",X"91",X"00",X"00",X"00",X"99",X"00",
		X"00",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"92",X"99",X"09",X"00",X"99",X"99",X"99",X"09",X"99",X"99",X"99",X"09",X"92",X"22",X"99",
		X"99",X"92",X"29",X"99",X"99",X"92",X"99",X"99",X"09",X"92",X"94",X"99",X"09",X"99",X"94",X"99",
		X"00",X"99",X"44",X"99",X"90",X"99",X"49",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"22",X"99",
		X"99",X"99",X"92",X"99",X"99",X"99",X"59",X"99",X"99",X"99",X"59",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"09",X"99",X"99",X"99",X"09",X"99",X"29",X"99",X"09",X"99",X"22",X"99",
		X"09",X"99",X"29",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"92",X"99",X"09",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"09",X"92",X"22",X"99",
		X"99",X"99",X"29",X"99",X"99",X"99",X"99",X"99",X"09",X"99",X"94",X"99",X"09",X"99",X"94",X"99",
		X"00",X"99",X"44",X"99",X"90",X"99",X"49",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"22",X"99",
		X"99",X"99",X"92",X"99",X"99",X"99",X"59",X"99",X"99",X"99",X"59",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"59",X"99",X"09",X"99",X"99",X"99",X"09",X"99",X"29",X"99",X"09",X"99",X"22",X"99",
		X"09",X"99",X"29",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"92",X"00",X"99",X"99",X"92",X"00",X"99",X"99",X"92",X"00",X"99",X"99",X"92",
		X"00",X"99",X"99",X"92",X"00",X"99",X"99",X"D9",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"09",X"99",X"99",X"00",X"09",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"09",X"99",X"22",X"99",X"09",X"99",X"22",X"99",X"09",X"99",X"22",X"99",
		X"09",X"99",X"22",X"9D",X"09",X"99",X"29",X"D9",X"09",X"99",X"99",X"99",X"00",X"99",X"22",X"99",
		X"00",X"99",X"22",X"99",X"00",X"99",X"22",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"09",X"99",X"99",X"99",X"09",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"09",X"99",X"99",X"99",X"00",X"09",X"99",X"99",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"E9",X"99",X"00",X"09",X"EE",X"93",X"00",X"99",X"3E",X"39",X"00",X"39",X"99",X"39",
		X"00",X"99",X"FF",X"99",X"00",X"99",X"99",X"90",X"00",X"9F",X"99",X"90",X"00",X"9F",X"99",X"90",
		X"00",X"99",X"AA",X"99",X"00",X"39",X"F9",X"39",X"00",X"33",X"99",X"39",X"00",X"33",X"33",X"99",
		X"00",X"33",X"99",X"90",X"00",X"33",X"39",X"00",X"00",X"93",X"39",X"00",X"99",X"93",X"94",X"00",
		X"93",X"99",X"99",X"99",X"93",X"09",X"99",X"39",X"93",X"09",X"B3",X"39",X"99",X"99",X"33",X"39",
		X"00",X"33",X"33",X"39",X"00",X"99",X"39",X"99",X"00",X"00",X"39",X"90",X"00",X"00",X"39",X"00",
		X"00",X"00",X"39",X"00",X"00",X"90",X"33",X"00",X"00",X"99",X"93",X"00",X"00",X"39",X"93",X"00",
		X"00",X"39",X"93",X"00",X"00",X"33",X"93",X"00",X"00",X"33",X"93",X"00",X"00",X"99",X"99",X"00",
		X"99",X"00",X"00",X"99",X"09",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"90",X"00",X"9D",
		X"09",X"99",X"00",X"D9",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"09",X"99",
		X"99",X"D9",X"09",X"99",X"99",X"99",X"09",X"99",X"99",X"D9",X"94",X"99",X"99",X"9D",X"44",X"99",
		X"99",X"99",X"44",X"99",X"99",X"9D",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"F9",X"99",
		X"99",X"99",X"D9",X"99",X"90",X"99",X"D9",X"09",X"90",X"99",X"D9",X"09",X"90",X"90",X"99",X"00",
		X"00",X"90",X"99",X"00",X"00",X"90",X"99",X"00",X"00",X"90",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"99",
		X"00",X"00",X"09",X"9D",X"00",X"90",X"99",X"D9",X"00",X"99",X"99",X"99",X"09",X"99",X"94",X"99",
		X"99",X"D9",X"49",X"99",X"99",X"9D",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"FD",X"99",X"99",X"99",X"3D",X"99",X"99",X"99",X"DD",X"99",X"99",X"99",X"D9",X"99",
		X"99",X"9D",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"9D",X"90",X"99",X"99",X"99",X"00",X"99",X"90",X"90",X"00",
		X"99",X"90",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"99",X"00",X"00",X"90",X"99",X"90",X"00",X"99",X"95",X"99",X"00",X"99",X"95",X"99",
		X"00",X"99",X"59",X"99",X"00",X"99",X"99",X"99",X"00",X"D9",X"99",X"99",X"00",X"D9",X"FD",X"99",
		X"00",X"DD",X"3D",X"99",X"00",X"9D",X"DD",X"99",X"00",X"9D",X"D9",X"99",X"00",X"9D",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"D9",X"90",X"00",X"99",X"99",X"00",X"00",X"90",X"99",X"00",X"00",X"90",X"09",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"A0",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"AA",X"A0",X"00",X"00",X"FF",X"FA",X"00",X"00",X"AF",X"FA",X"00",X"00",X"AA",X"FF",
		X"00",X"0A",X"FF",X"FF",X"00",X"0A",X"FA",X"FF",X"00",X"AA",X"FF",X"FF",X"00",X"FA",X"AA",X"FF",
		X"00",X"AA",X"FA",X"AF",X"00",X"AF",X"FF",X"AF",X"00",X"AF",X"FF",X"FF",X"00",X"AA",X"FF",X"FF",
		X"00",X"FA",X"AF",X"FF",X"00",X"FA",X"AA",X"FF",X"00",X"FA",X"FF",X"FF",X"00",X"FA",X"FF",X"FA",
		X"00",X"FA",X"AF",X"FF",X"00",X"AF",X"AF",X"FF",X"00",X"AF",X"AA",X"AF",X"00",X"AF",X"FA",X"AA",
		X"00",X"AF",X"AA",X"FA",X"00",X"AF",X"FF",X"FA",X"00",X"FF",X"FF",X"AA",X"00",X"FF",X"FF",X"FF",
		X"00",X"AA",X"FF",X"FF",X"00",X"FF",X"FF",X"AA",X"00",X"AF",X"FF",X"00",X"00",X"0A",X"AA",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",
		X"00",X"00",X"00",X"AA",X"0A",X"00",X"00",X"FF",X"0A",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"A0",X"AF",X"00",X"00",X"AA",X"AF",
		X"00",X"00",X"FF",X"AA",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FA",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"FF",X"00",X"0A",
		X"AA",X"FF",X"00",X"AA",X"AF",X"FF",X"00",X"AF",X"AF",X"FF",X"00",X"AF",X"AA",X"FF",X"00",X"FF",
		X"00",X"AF",X"00",X"AA",X"00",X"0A",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"A0",X"00",X"00",X"0A",X"A0",X"A0",X"00",X"00",X"0A",X"A0",X"00",X"00",X"0A",X"A0",X"00",
		X"00",X"00",X"A0",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"A0",X"0A",X"00",X"00",X"00",X"00",
		X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"0F",X"F0",X"00",X"3F",X"F3",X"30",
		X"00",X"0F",X"F0",X"00",X"AA",X"F3",X"F0",X"00",X"00",X"30",X"F0",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"3F",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"0A",X"00",X"00",X"00",X"0A",X"00",X"00",
		X"00",X"A0",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"9F",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"90",X"00",X"00",X"FF",X"90",X"00",X"00",X"FF",X"90",X"00",X"00",X"FF",X"90",
		X"00",X"00",X"FF",X"90",X"00",X"00",X"FF",X"90",X"00",X"00",X"FF",X"90",X"00",X"00",X"FF",X"90",
		X"00",X"00",X"FF",X"90",X"00",X"00",X"FF",X"90",X"00",X"00",X"FF",X"90",X"00",X"00",X"FF",X"90",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"99",X"FF",X"00",
		X"00",X"95",X"99",X"00",X"00",X"95",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"95",X"00",X"90",
		X"00",X"55",X"00",X"90",X"00",X"99",X"99",X"90",X"00",X"00",X"95",X"90",X"00",X"00",X"99",X"90",
		X"00",X"00",X"99",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"9F",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"F9",X"90",X"00",X"00",X"FF",X"90",
		X"00",X"00",X"FF",X"90",X"00",X"00",X"F9",X"90",X"00",X"00",X"F9",X"90",X"00",X"00",X"FF",X"90",
		X"00",X"00",X"FF",X"90",X"00",X"00",X"FF",X"90",X"00",X"00",X"FF",X"90",X"00",X"00",X"FF",X"90",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"99",X"FF",X"00",
		X"00",X"95",X"99",X"00",X"00",X"95",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"95",X"00",X"90",
		X"00",X"55",X"00",X"90",X"00",X"99",X"99",X"90",X"00",X"00",X"95",X"90",X"00",X"00",X"99",X"90",
		X"00",X"00",X"99",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"9F",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"F9",X"00",
		X"00",X"00",X"F9",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"F9",X"90",X"00",X"00",X"FF",X"90",
		X"00",X"00",X"FF",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"F9",X"90",X"00",X"00",X"F9",X"90",
		X"00",X"00",X"F9",X"90",X"00",X"00",X"9F",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"9F",X"90",
		X"00",X"00",X"99",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"FF",X"00",
		X"00",X"95",X"99",X"00",X"00",X"95",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"95",X"00",X"90",
		X"00",X"55",X"00",X"90",X"00",X"99",X"99",X"90",X"00",X"00",X"95",X"90",X"00",X"00",X"99",X"90",
		X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"F9",X"00",X"50",
		X"00",X"99",X"0E",X"00",X"00",X"90",X"99",X"00",X"00",X"90",X"E9",X"00",X"00",X"00",X"99",X"00",
		X"00",X"0A",X"99",X"00",X"00",X"0A",X"99",X"00",X"00",X"0A",X"99",X"0A",X"00",X"0A",X"99",X"00",
		X"00",X"0A",X"99",X"00",X"00",X"0A",X"99",X"00",X"00",X"05",X"99",X"00",X"00",X"0A",X"99",X"83",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"77",X"00",X"00",X"90",X"E9",X"00",
		X"00",X"90",X"99",X"00",X"00",X"90",X"77",X"00",X"00",X"00",X"E7",X"10",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9F",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"99",X"00",X"59",X"00",X"95",X"00",X"95",X"00",X"59",X"00",X"95",X"00",X"59",
		X"00",X"95",X"99",X"59",X"00",X"95",X"99",X"59",X"00",X"95",X"99",X"59",X"09",X"99",X"99",X"99",
		X"09",X"A9",X"44",X"9A",X"99",X"AA",X"99",X"AA",X"9A",X"3A",X"99",X"33",X"9A",X"33",X"99",X"5A",
		X"9A",X"33",X"99",X"35",X"9A",X"5A",X"44",X"33",X"9A",X"3A",X"44",X"AA",X"9A",X"99",X"44",X"AA",
		X"9A",X"90",X"99",X"9A",X"9A",X"90",X"99",X"99",X"93",X"90",X"99",X"09",X"93",X"90",X"99",X"09",
		X"9A",X"00",X"99",X"09",X"9A",X"00",X"99",X"09",X"9A",X"00",X"99",X"09",X"93",X"00",X"44",X"00",
		X"9A",X"00",X"99",X"00",X"9A",X"09",X"00",X"90",X"9A",X"99",X"00",X"99",X"9A",X"95",X"00",X"59",
		X"9A",X"59",X"00",X"95",X"9A",X"99",X"00",X"99",X"9A",X"99",X"00",X"99",X"99",X"00",X"00",X"00",
		X"00",X"99",X"00",X"99",X"00",X"59",X"00",X"95",X"00",X"95",X"00",X"59",X"00",X"95",X"00",X"59",
		X"00",X"95",X"99",X"59",X"00",X"95",X"99",X"59",X"00",X"95",X"99",X"59",X"00",X"99",X"99",X"99",
		X"00",X"99",X"44",X"99",X"00",X"9A",X"99",X"A9",X"00",X"9A",X"99",X"39",X"00",X"93",X"99",X"39",
		X"00",X"93",X"99",X"A9",X"00",X"9A",X"44",X"A9",X"00",X"93",X"44",X"39",X"00",X"93",X"44",X"A9",
		X"00",X"9A",X"99",X"A9",X"00",X"9A",X"99",X"39",X"00",X"9A",X"99",X"A9",X"00",X"9A",X"99",X"A9",
		X"00",X"9A",X"99",X"39",X"00",X"93",X"99",X"39",X"00",X"93",X"99",X"A9",X"00",X"93",X"44",X"99",
		X"00",X"9A",X"99",X"90",X"00",X"99",X"00",X"90",X"00",X"09",X"00",X"99",X"00",X"95",X"00",X"59",
		X"00",X"95",X"00",X"59",X"00",X"95",X"00",X"59",X"00",X"A9",X"00",X"99",X"00",X"9A",X"00",X"90",
		X"00",X"99",X"00",X"99",X"00",X"59",X"00",X"95",X"00",X"95",X"00",X"59",X"00",X"95",X"00",X"59",
		X"00",X"95",X"99",X"59",X"00",X"95",X"99",X"59",X"00",X"95",X"99",X"59",X"00",X"99",X"99",X"99",
		X"00",X"99",X"44",X"90",X"00",X"9A",X"99",X"99",X"00",X"9A",X"99",X"A9",X"00",X"93",X"99",X"3A",
		X"00",X"93",X"99",X"AA",X"00",X"A3",X"44",X"A3",X"00",X"A3",X"44",X"A3",X"00",X"AA",X"44",X"A3",
		X"00",X"3A",X"99",X"AA",X"00",X"3A",X"99",X"3A",X"00",X"3A",X"99",X"3A",X"00",X"AA",X"99",X"A3",
		X"00",X"3A",X"99",X"A3",X"00",X"3A",X"99",X"A3",X"00",X"3A",X"99",X"3A",X"00",X"3A",X"44",X"3A",
		X"00",X"AA",X"99",X"AA",X"00",X"A9",X"00",X"9A",X"00",X"99",X"00",X"99",X"00",X"95",X"00",X"59",
		X"00",X"95",X"00",X"59",X"00",X"95",X"00",X"59",X"00",X"99",X"00",X"99",X"00",X"09",X"00",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"44",X"00",
		X"00",X"94",X"99",X"99",X"00",X"44",X"22",X"49",X"00",X"49",X"99",X"44",X"00",X"99",X"AA",X"44",
		X"99",X"99",X"9A",X"11",X"91",X"59",X"99",X"51",X"9E",X"11",X"99",X"55",X"99",X"11",X"11",X"55",
		X"09",X"11",X"71",X"55",X"00",X"E9",X"79",X"EE",X"00",X"EE",X"77",X"99",X"00",X"99",X"99",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"44",X"00",
		X"00",X"94",X"99",X"99",X"00",X"44",X"22",X"49",X"00",X"49",X"99",X"44",X"00",X"92",X"AA",X"44",
		X"99",X"99",X"9A",X"11",X"91",X"79",X"99",X"71",X"9E",X"11",X"99",X"77",X"99",X"11",X"11",X"77",
		X"09",X"11",X"51",X"77",X"00",X"E9",X"59",X"EE",X"00",X"EE",X"55",X"99",X"00",X"99",X"99",X"90",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"9E",X"09",X"00",X"00",X"F9",X"09",
		X"00",X"00",X"FF",X"99",X"00",X"90",X"FF",X"93",X"00",X"99",X"F4",X"93",X"00",X"33",X"FF",X"9B",
		X"00",X"93",X"FF",X"9B",X"00",X"93",X"FF",X"93",X"00",X"B9",X"4F",X"9B",X"00",X"B9",X"99",X"9B",
		X"00",X"39",X"39",X"39",X"00",X"93",X"33",X"39",X"00",X"99",X"93",X"33",X"00",X"09",X"99",X"33",
		X"00",X"00",X"99",X"33",X"00",X"A0",X"33",X"39",X"04",X"AA",X"99",X"99",X"04",X"05",X"B9",X"90",
		X"00",X"95",X"99",X"00",X"00",X"94",X"93",X"91",X"00",X"49",X"93",X"91",X"40",X"79",X"43",X"15",
		X"00",X"99",X"44",X"11",X"00",X"5A",X"34",X"59",X"00",X"11",X"94",X"11",X"70",X"A5",X"A1",X"55",
		X"00",X"15",X"11",X"91",X"00",X"50",X"A1",X"00",X"04",X"00",X"11",X"00",X"47",X"07",X"10",X"07",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"09",
		X"00",X"00",X"99",X"99",X"00",X"90",X"A9",X"93",X"00",X"99",X"FF",X"93",X"00",X"33",X"FF",X"9B",
		X"00",X"93",X"9F",X"9B",X"00",X"93",X"9F",X"93",X"00",X"B9",X"F9",X"9B",X"00",X"B9",X"99",X"9B",
		X"00",X"39",X"33",X"39",X"00",X"93",X"39",X"39",X"00",X"99",X"33",X"33",X"00",X"09",X"99",X"33",
		X"00",X"00",X"B9",X"33",X"00",X"00",X"33",X"39",X"00",X"00",X"99",X"99",X"00",X"00",X"B9",X"90",
		X"00",X"09",X"33",X"00",X"00",X"99",X"39",X"00",X"00",X"93",X"33",X"00",X"00",X"33",X"33",X"00",
		X"00",X"39",X"39",X"00",X"00",X"39",X"33",X"90",X"00",X"39",X"33",X"99",X"00",X"99",X"33",X"39",
		X"00",X"00",X"33",X"99",X"00",X"00",X"93",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"90",X"00",X"00",X"FF",X"90",X"00",X"00",X"FF",X"90",X"00",X"00",X"FF",X"90",
		X"00",X"00",X"FF",X"90",X"00",X"00",X"FF",X"90",X"00",X"00",X"FF",X"90",X"00",X"00",X"FF",X"90",
		X"00",X"00",X"FF",X"90",X"00",X"00",X"FF",X"90",X"00",X"00",X"FF",X"90",X"00",X"00",X"FF",X"90",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"99",X"FF",X"00",
		X"00",X"95",X"99",X"00",X"00",X"95",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"95",X"00",X"90",
		X"00",X"55",X"00",X"90",X"00",X"99",X"99",X"90",X"00",X"00",X"95",X"90",X"00",X"00",X"99",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"99",X"90",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"94",X"00",X"00",X"9B",X"94",X"90",
		X"09",X"99",X"99",X"99",X"09",X"E9",X"99",X"B9",X"99",X"EE",X"B9",X"BB",X"91",X"9E",X"BB",X"9B",
		X"91",X"99",X"99",X"9B",X"91",X"11",X"59",X"BB",X"91",X"EE",X"59",X"99",X"91",X"EE",X"99",X"95",
		X"91",X"EE",X"99",X"99",X"91",X"E1",X"99",X"B9",X"91",X"11",X"99",X"99",X"91",X"19",X"BB",X"9B",
		X"91",X"99",X"9B",X"B9",X"91",X"9B",X"99",X"00",X"91",X"9B",X"B7",X"00",X"91",X"BB",X"BB",X"00",
		X"91",X"B9",X"BB",X"00",X"91",X"99",X"BB",X"00",X"91",X"90",X"19",X"00",X"91",X"90",X"99",X"90",
		X"91",X"00",X"B9",X"99",X"91",X"00",X"B9",X"B9",X"91",X"00",X"B9",X"BB",X"91",X"00",X"B9",X"BB",
		X"99",X"00",X"B9",X"BB",X"00",X"00",X"B9",X"9B",X"00",X"00",X"B9",X"9B",X"00",X"00",X"99",X"99",
		X"00",X"99",X"00",X"00",X"00",X"E9",X"99",X"00",X"00",X"99",X"93",X"00",X"00",X"9B",X"93",X"90",
		X"00",X"99",X"99",X"99",X"00",X"19",X"99",X"B9",X"00",X"E9",X"B9",X"BB",X"00",X"E1",X"BB",X"9B",
		X"00",X"EE",X"99",X"9B",X"00",X"1E",X"59",X"BB",X"00",X"11",X"59",X"99",X"00",X"11",X"99",X"95",
		X"00",X"11",X"99",X"99",X"00",X"11",X"BB",X"B9",X"00",X"99",X"BB",X"99",X"00",X"BB",X"99",X"BB",
		X"00",X"9B",X"B7",X"B9",X"00",X"99",X"B7",X"99",X"00",X"91",X"B7",X"00",X"00",X"91",X"BB",X"00",
		X"00",X"91",X"BB",X"00",X"00",X"99",X"BB",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"99",X"90",
		X"00",X"00",X"B9",X"99",X"00",X"00",X"B9",X"B9",X"00",X"00",X"B9",X"BB",X"00",X"00",X"B9",X"BB",
		X"00",X"00",X"B9",X"9B",X"00",X"00",X"B9",X"9B",X"00",X"00",X"B9",X"99",X"00",X"00",X"99",X"09",
		X"00",X"00",X"99",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"66",X"00",X"00",X"99",X"66",X"00",
		X"00",X"66",X"66",X"00",X"00",X"99",X"66",X"00",X"00",X"EE",X"66",X"00",X"00",X"EE",X"6D",X"00",
		X"00",X"99",X"6D",X"90",X"00",X"94",X"99",X"90",X"00",X"44",X"C9",X"90",X"00",X"99",X"C9",X"90",
		X"00",X"CC",X"99",X"90",X"00",X"CC",X"9D",X"90",X"00",X"C9",X"9D",X"90",X"00",X"99",X"DD",X"90",
		X"00",X"99",X"99",X"90",X"00",X"95",X"99",X"90",X"00",X"99",X"99",X"90",X"00",X"CC",X"99",X"90",
		X"00",X"CC",X"96",X"90",X"00",X"99",X"96",X"90",X"00",X"66",X"66",X"90",X"00",X"69",X"66",X"00",
		X"00",X"99",X"66",X"00",X"00",X"90",X"96",X"00",X"00",X"90",X"99",X"00",X"00",X"09",X"C9",X"00",
		X"00",X"09",X"99",X"00",X"00",X"09",X"77",X"00",X"00",X"09",X"77",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",
		X"00",X"99",X"66",X"00",X"00",X"EE",X"66",X"90",X"00",X"EE",X"66",X"90",X"00",X"99",X"6D",X"90",
		X"00",X"94",X"99",X"90",X"00",X"94",X"C9",X"90",X"00",X"99",X"C9",X"90",X"00",X"CC",X"99",X"90",
		X"00",X"CC",X"9D",X"90",X"00",X"C9",X"9D",X"99",X"00",X"99",X"DD",X"69",X"00",X"99",X"DD",X"69",
		X"00",X"95",X"DD",X"69",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"CC",X"99",X"99",
		X"00",X"99",X"66",X"69",X"00",X"00",X"66",X"69",X"00",X"99",X"69",X"69",X"00",X"96",X"99",X"99",
		X"00",X"96",X"90",X"99",X"00",X"66",X"99",X"99",X"00",X"66",X"9C",X"99",X"00",X"99",X"99",X"66",
		X"00",X"77",X"00",X"66",X"00",X"77",X"00",X"99",X"00",X"99",X"00",X"97",X"00",X"00",X"00",X"99",
		X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"E9",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"9A",X"00",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"9E",X"00",X"E9",X"99",X"EE",X"00",X"E9",X"9E",X"9E",X"00",X"99",X"E9",X"99",
		X"99",X"9E",X"99",X"9B",X"9E",X"9E",X"99",X"9B",X"9E",X"EE",X"99",X"BB",X"99",X"EE",X"99",X"99",
		X"91",X"9E",X"99",X"9E",X"91",X"9E",X"EE",X"9E",X"99",X"99",X"99",X"9E",X"00",X"9E",X"E9",X"99",
		X"00",X"EE",X"E9",X"90",X"00",X"99",X"9E",X"00",X"00",X"19",X"9B",X"00",X"00",X"E1",X"9B",X"00",
		X"00",X"E9",X"9B",X"00",X"00",X"99",X"99",X"90",X"00",X"B9",X"EE",X"99",X"00",X"BE",X"EE",X"9E",
		X"09",X"99",X"99",X"EE",X"09",X"09",X"09",X"EE",X"09",X"09",X"09",X"99",X"09",X"00",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"E9",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"9A",X"00",X"00",X"99",X"9A",X"00",
		X"00",X"91",X"99",X"00",X"00",X"E9",X"99",X"90",X"00",X"E9",X"9E",X"99",X"00",X"B9",X"E9",X"EE",
		X"09",X"9B",X"99",X"99",X"09",X"99",X"99",X"19",X"99",X"E9",X"99",X"99",X"9E",X"E9",X"99",X"E9",
		X"9E",X"99",X"99",X"EE",X"9E",X"9E",X"99",X"EE",X"99",X"99",X"99",X"99",X"9E",X"9E",X"E9",X"9B",
		X"9E",X"9E",X"E9",X"9B",X"99",X"99",X"9E",X"99",X"00",X"B9",X"9B",X"09",X"00",X"EE",X"9B",X"00",
		X"00",X"99",X"9B",X"90",X"09",X"9E",X"09",X"99",X"09",X"EE",X"00",X"E9",X"99",X"99",X"09",X"99",
		X"9E",X"E9",X"09",X"E9",X"9E",X"E9",X"09",X"E9",X"99",X"E9",X"00",X"EE",X"00",X"99",X"00",X"99",
		X"09",X"99",X"00",X"99",X"99",X"77",X"00",X"79",X"93",X"77",X"09",X"79",X"99",X"77",X"09",X"77",
		X"97",X"77",X"09",X"97",X"97",X"77",X"09",X"99",X"97",X"99",X"09",X"99",X"97",X"99",X"99",X"99",
		X"97",X"90",X"77",X"79",X"97",X"99",X"77",X"99",X"99",X"77",X"77",X"99",X"00",X"77",X"77",X"77",
		X"00",X"77",X"77",X"77",X"09",X"77",X"77",X"77",X"99",X"77",X"99",X"97",X"97",X"94",X"49",X"97",
		X"97",X"94",X"49",X"97",X"97",X"99",X"44",X"49",X"97",X"94",X"99",X"49",X"97",X"99",X"11",X"A9",
		X"97",X"09",X"11",X"99",X"94",X"00",X"11",X"79",X"94",X"00",X"99",X"77",X"0A",X"00",X"19",X"77",
		X"09",X"00",X"19",X"97",X"09",X"00",X"99",X"97",X"00",X"00",X"99",X"97",X"00",X"00",X"00",X"97",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",
		X"09",X"99",X"00",X"99",X"99",X"77",X"00",X"99",X"99",X"77",X"09",X"99",X"93",X"77",X"09",X"79",
		X"93",X"77",X"09",X"97",X"99",X"77",X"09",X"99",X"97",X"79",X"09",X"99",X"97",X"79",X"99",X"99",
		X"97",X"79",X"77",X"99",X"97",X"90",X"77",X"77",X"99",X"99",X"77",X"99",X"00",X"77",X"77",X"90",
		X"00",X"77",X"77",X"99",X"00",X"77",X"77",X"77",X"00",X"97",X"99",X"77",X"00",X"97",X"49",X"77",
		X"00",X"97",X"49",X"77",X"00",X"99",X"44",X"77",X"00",X"97",X"99",X"77",X"00",X"99",X"11",X"77",
		X"00",X"49",X"11",X"79",X"00",X"44",X"11",X"47",X"00",X"74",X"99",X"49",X"00",X"79",X"19",X"79",
		X"00",X"77",X"19",X"79",X"00",X"79",X"00",X"A9",X"00",X"99",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"99",X"00",X"92",X"09",X"99",X"00",X"92",X"99",X"99",
		X"00",X"92",X"22",X"99",X"00",X"22",X"29",X"90",X"00",X"29",X"99",X"90",X"00",X"29",X"99",X"99",
		X"00",X"92",X"94",X"99",X"00",X"99",X"99",X"99",X"09",X"99",X"99",X"99",X"09",X"99",X"99",X"99",
		X"09",X"99",X"95",X"90",X"09",X"99",X"99",X"90",X"09",X"99",X"95",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"D9",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"90",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"00",X"99",X"99",
		X"00",X"00",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"22",X"99",X"00",X"92",X"22",X"99",X"00",X"92",X"29",X"99",X"00",X"92",X"99",X"99",
		X"00",X"99",X"99",X"90",X"00",X"99",X"99",X"90",X"00",X"99",X"99",X"09",X"00",X"99",X"59",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"59",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"DD",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"09",X"99",X"99",X"00",X"09",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"93",X"00",
		X"00",X"99",X"34",X"00",X"00",X"92",X"99",X"00",X"00",X"29",X"22",X"00",X"00",X"24",X"22",X"00",
		X"09",X"22",X"92",X"00",X"09",X"99",X"99",X"09",X"99",X"95",X"99",X"99",X"92",X"99",X"99",X"22",
		X"92",X"29",X"99",X"22",X"92",X"99",X"92",X"29",X"99",X"99",X"22",X"99",X"00",X"99",X"29",X"9D",
		X"00",X"92",X"99",X"2D",X"00",X"99",X"92",X"D2",X"00",X"D9",X"22",X"DD",X"00",X"2D",X"22",X"DD",
		X"00",X"DD",X"22",X"2D",X"00",X"DD",X"22",X"D9",X"00",X"DD",X"22",X"99",X"00",X"D2",X"22",X"00",
		X"00",X"DD",X"A2",X"00",X"00",X"99",X"22",X"99",X"00",X"09",X"99",X"22",X"00",X"09",X"99",X"22",
		X"00",X"99",X"99",X"92",X"00",X"92",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"99",X"00",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"94",X"00",
		X"00",X"99",X"44",X"00",X"00",X"92",X"99",X"00",X"00",X"29",X"22",X"00",X"00",X"29",X"22",X"00",
		X"00",X"22",X"92",X"00",X"00",X"99",X"99",X"00",X"00",X"95",X"99",X"00",X"00",X"99",X"95",X"00",
		X"00",X"29",X"99",X"00",X"00",X"22",X"92",X"90",X"00",X"99",X"29",X"90",X"00",X"99",X"99",X"90",
		X"00",X"9D",X"9D",X"90",X"00",X"9D",X"9D",X"90",X"00",X"92",X"9D",X"99",X"00",X"9D",X"9D",X"D9",
		X"00",X"9D",X"99",X"D9",X"00",X"9D",X"29",X"D9",X"00",X"99",X"29",X"D9",X"00",X"09",X"29",X"D9",
		X"00",X"09",X"99",X"99",X"00",X"09",X"22",X"90",X"00",X"09",X"92",X"00",X"00",X"00",X"92",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"09",
		X"00",X"00",X"99",X"99",X"00",X"90",X"F9",X"93",X"00",X"99",X"FF",X"93",X"00",X"33",X"A9",X"9B",
		X"00",X"93",X"99",X"9B",X"00",X"93",X"99",X"93",X"00",X"B9",X"99",X"9B",X"00",X"B9",X"33",X"9B",
		X"00",X"39",X"39",X"39",X"00",X"93",X"33",X"39",X"00",X"99",X"33",X"33",X"00",X"09",X"93",X"33",
		X"00",X"00",X"99",X"33",X"00",X"00",X"33",X"39",X"00",X"00",X"99",X"99",X"00",X"00",X"B9",X"90",
		X"00",X"99",X"99",X"90",X"00",X"94",X"93",X"99",X"00",X"49",X"93",X"49",X"00",X"99",X"33",X"44",
		X"99",X"99",X"33",X"11",X"91",X"59",X"33",X"51",X"9E",X"11",X"99",X"55",X"99",X"11",X"11",X"55",
		X"09",X"11",X"71",X"55",X"00",X"E9",X"79",X"EE",X"00",X"EE",X"77",X"99",X"00",X"99",X"99",X"90",
		X"00",X"00",X"9E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"09",X"00",X"00",X"99",X"99",
		X"00",X"90",X"F9",X"93",X"00",X"99",X"99",X"93",X"00",X"33",X"99",X"9B",X"00",X"93",X"99",X"9B",
		X"00",X"93",X"F9",X"93",X"00",X"B9",X"99",X"9B",X"00",X"B9",X"33",X"9B",X"00",X"39",X"39",X"39",
		X"00",X"93",X"33",X"39",X"00",X"99",X"33",X"33",X"00",X"09",X"93",X"33",X"00",X"00",X"99",X"33",
		X"00",X"00",X"33",X"39",X"00",X"00",X"99",X"99",X"00",X"00",X"B9",X"90",X"00",X"00",X"99",X"00",
		X"00",X"99",X"93",X"90",X"00",X"94",X"93",X"99",X"00",X"49",X"33",X"49",X"00",X"99",X"33",X"44",
		X"99",X"99",X"33",X"11",X"91",X"79",X"33",X"71",X"9E",X"11",X"99",X"77",X"99",X"11",X"11",X"77",
		X"09",X"11",X"51",X"77",X"00",X"E9",X"59",X"EE",X"00",X"EE",X"55",X"99",X"00",X"99",X"99",X"90",
		X"00",X"00",X"99",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"9F",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"49",X"00",
		X"00",X"00",X"F9",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"F9",X"90",X"00",X"00",X"FF",X"90",
		X"00",X"00",X"9F",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"49",X"90",X"00",X"00",X"F9",X"90",
		X"00",X"00",X"F9",X"90",X"00",X"00",X"9F",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"49",X"90",
		X"00",X"00",X"99",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"FF",X"00",
		X"00",X"95",X"99",X"00",X"00",X"95",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"95",X"00",X"90",
		X"00",X"55",X"00",X"90",X"00",X"99",X"99",X"90",X"00",X"00",X"95",X"90",X"00",X"00",X"99",X"90",
		X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"F9",X"04",X"00",X"00",X"F9",X"00",X"50",
		X"00",X"99",X"0E",X"00",X"00",X"90",X"99",X"00",X"00",X"90",X"E9",X"00",X"00",X"00",X"99",X"00",
		X"00",X"0A",X"9A",X"00",X"00",X"0A",X"49",X"00",X"00",X"0A",X"44",X"0A",X"00",X"0A",X"4A",X"00",
		X"00",X"0A",X"A4",X"00",X"00",X"0A",X"A4",X"00",X"00",X"05",X"49",X"00",X"00",X"0A",X"9A",X"83",
		X"00",X"00",X"A4",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"74",X"00",X"00",X"90",X"E9",X"00",
		X"00",X"90",X"9A",X"00",X"00",X"90",X"77",X"00",X"00",X"00",X"E7",X"10",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9F",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
