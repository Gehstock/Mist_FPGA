library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_PGM is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_PGM is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"3A",X"00",X"B0",X"31",X"00",X"88",X"3E",X"9B",X"32",X"03",X"98",X"AF",X"21",X"00",X"A8",X"06",
		X"08",X"77",X"23",X"10",X"FC",X"21",X"00",X"90",X"06",X"7D",X"77",X"23",X"10",X"FC",X"21",X"00",
		X"88",X"0E",X"04",X"CD",X"B7",X"00",X"CD",X"6C",X"09",X"21",X"10",X"8B",X"FD",X"21",X"13",X"01",
		X"06",X"09",X"CD",X"3D",X"0B",X"31",X"20",X"88",X"21",X"00",X"80",X"0E",X"08",X"CD",X"B7",X"00",
		X"31",X"00",X"88",X"21",X"10",X"8B",X"FD",X"21",X"1C",X"01",X"06",X"09",X"CD",X"3D",X"0B",X"21",
		X"00",X"00",X"CD",X"A0",X"00",X"21",X"F0",X"8A",X"36",X"15",X"21",X"00",X"10",X"CD",X"A0",X"00",
		X"3A",X"00",X"98",X"18",X"04",X"00",X"C3",X"4D",X"12",X"E6",X"0A",X"FE",X"0A",X"CA",X"56",X"01",
		X"11",X"06",X"00",X"FD",X"21",X"25",X"01",X"01",X"07",X"06",X"21",X"10",X"8B",X"3A",X"00",X"98",
		X"E6",X"0A",X"CA",X"56",X"01",X"3A",X"00",X"98",X"07",X"38",X"08",X"CD",X"3D",X"0B",X"3A",X"00",
		X"B0",X"18",X"DD",X"FD",X"19",X"0D",X"20",X"F0",X"CD",X"3D",X"0B",X"3A",X"00",X"B0",X"18",X"D0",
		X"01",X"10",X"00",X"AF",X"86",X"23",X"10",X"FC",X"08",X"3A",X"00",X"B0",X"08",X"0D",X"20",X"F4",
		X"B7",X"C8",X"3A",X"00",X"B0",X"18",X"FB",X"70",X"7E",X"B8",X"3A",X"00",X"B0",X"20",X"FB",X"10",
		X"F6",X"51",X"36",X"00",X"23",X"10",X"FB",X"3A",X"00",X"B0",X"0D",X"20",X"F5",X"4A",X"11",X"55",
		X"00",X"CD",X"FB",X"00",X"11",X"AA",X"55",X"CD",X"E3",X"00",X"11",X"FF",X"AA",X"CD",X"FB",X"00",
		X"11",X"00",X"FF",X"C5",X"7E",X"BA",X"3A",X"00",X"B0",X"20",X"FB",X"73",X"7E",X"BB",X"3A",X"00",
		X"B0",X"20",X"FB",X"23",X"10",X"EE",X"0D",X"20",X"EB",X"C1",X"C9",X"C5",X"2B",X"7E",X"BA",X"3A",
		X"00",X"B0",X"20",X"FB",X"73",X"7E",X"BB",X"3A",X"00",X"B0",X"20",X"FB",X"10",X"EE",X"0D",X"20",
		X"EB",X"C1",X"C9",X"22",X"11",X"1D",X"10",X"01",X"17",X"18",X"1A",X"1B",X"02",X"13",X"10",X"22",
		X"1F",X"1D",X"10",X"10",X"10",X"13",X"1F",X"19",X"1E",X"10",X"01",X"13",X"1F",X"19",X"1E",X"10",
		X"02",X"1C",X"15",X"16",X"24",X"10",X"10",X"22",X"19",X"17",X"18",X"24",X"10",X"20",X"1C",X"11",
		X"29",X"10",X"02",X"10",X"10",X"10",X"10",X"10",X"10",X"20",X"1C",X"11",X"29",X"10",X"01",X"10",
		X"10",X"10",X"10",X"10",X"10",X"E6",X"3A",X"00",X"B0",X"3E",X"80",X"32",X"A4",X"80",X"21",X"00",
		X"88",X"11",X"01",X"88",X"01",X"FF",X"03",X"36",X"10",X"ED",X"B0",X"3E",X"88",X"32",X"03",X"A0",
		X"3E",X"55",X"32",X"CB",X"80",X"32",X"78",X"80",X"32",X"03",X"A8",X"21",X"01",X"A8",X"71",X"0D",
		X"71",X"0E",X"3D",X"11",X"40",X"90",X"21",X"C7",X"10",X"ED",X"B0",X"FD",X"21",X"B8",X"0F",X"21",
		X"A0",X"8B",X"06",X"1B",X"CD",X"3D",X"0B",X"21",X"A1",X"8B",X"06",X"1A",X"CD",X"3D",X"0B",X"21",
		X"A2",X"8B",X"06",X"17",X"CD",X"3D",X"0B",X"3E",X"04",X"CD",X"2F",X"0D",X"3E",X"0A",X"11",X"CE",
		X"80",X"21",X"87",X"0F",X"01",X"0A",X"00",X"ED",X"B0",X"3D",X"20",X"F5",X"11",X"55",X"81",X"21",
		X"87",X"0F",X"0E",X"06",X"ED",X"B0",X"3D",X"20",X"F6",X"21",X"A9",X"80",X"11",X"AA",X"80",X"01",
		X"0D",X"00",X"36",X"00",X"ED",X"B0",X"18",X"49",X"CD",X"53",X"09",X"3A",X"A4",X"80",X"87",X"20",
		X"40",X"06",X"00",X"3A",X"A8",X"80",X"21",X"AB",X"80",X"CD",X"CF",X"0A",X"CD",X"84",X"0A",X"3A",
		X"A8",X"80",X"CB",X"3F",X"C4",X"81",X"0A",X"3E",X"01",X"CD",X"2C",X"0D",X"3A",X"A8",X"80",X"CB",
		X"3F",X"28",X"06",X"CD",X"FB",X"0B",X"CD",X"08",X"0D",X"CD",X"FB",X"0B",X"3E",X"04",X"CD",X"18",
		X"09",X"32",X"A8",X"80",X"3E",X"84",X"32",X"A4",X"80",X"3E",X"0C",X"CD",X"18",X"09",X"CD",X"2C",
		X"0D",X"3E",X"84",X"32",X"A4",X"80",X"3A",X"00",X"98",X"E6",X"2A",X"20",X"38",X"CD",X"6C",X"09",
		X"21",X"A8",X"8B",X"DD",X"21",X"A9",X"80",X"FD",X"21",X"3F",X"0F",X"CD",X"2A",X"0B",X"21",X"AA",
		X"8B",X"CD",X"2A",X"0B",X"21",X"AC",X"8B",X"CD",X"2A",X"0B",X"21",X"AE",X"8B",X"CD",X"2A",X"0B",
		X"21",X"B0",X"8B",X"CD",X"10",X"0B",X"21",X"B2",X"8B",X"CD",X"10",X"0B",X"3A",X"00",X"98",X"E6",
		X"0A",X"FE",X"0A",X"20",X"F7",X"21",X"75",X"80",X"7E",X"B7",X"20",X"02",X"36",X"10",X"CB",X"16",
		X"CD",X"6C",X"09",X"21",X"40",X"8A",X"CD",X"61",X"09",X"21",X"41",X"8A",X"3A",X"A8",X"80",X"D6",
		X"02",X"28",X"02",X"3E",X"10",X"CD",X"62",X"09",X"21",X"91",X"0F",X"11",X"37",X"80",X"01",X"27",
		X"00",X"ED",X"B0",X"AF",X"32",X"70",X"80",X"3A",X"02",X"98",X"E6",X"08",X"0F",X"0F",X"6F",X"3E",
		X"05",X"95",X"6F",X"3A",X"A4",X"80",X"87",X"7D",X"CA",X"44",X"03",X"3E",X"01",X"CD",X"2C",X"0D",
		X"3E",X"FF",X"32",X"CB",X"80",X"CD",X"4A",X"0B",X"21",X"AC",X"8B",X"06",X"1C",X"CD",X"8D",X"0B",
		X"06",X"1B",X"CD",X"8D",X"0B",X"06",X"15",X"CD",X"8D",X"0B",X"06",X"18",X"CD",X"8D",X"0B",X"06",
		X"1A",X"CD",X"8D",X"0B",X"06",X"10",X"CD",X"8D",X"0B",X"2C",X"06",X"1B",X"CD",X"8D",X"0B",X"06",
		X"1B",X"CD",X"8D",X"0B",X"06",X"1A",X"CD",X"8D",X"0B",X"06",X"1A",X"CD",X"8D",X"0B",X"2C",X"06",
		X"17",X"CD",X"8D",X"0B",X"06",X"19",X"CD",X"8D",X"0B",X"06",X"0D",X"CD",X"8D",X"0B",X"06",X"17",
		X"CD",X"8D",X"0B",X"06",X"1A",X"CD",X"8D",X"0B",X"06",X"1C",X"CD",X"8D",X"0B",X"3E",X"55",X"32",
		X"CB",X"80",X"3E",X"08",X"CD",X"18",X"09",X"CD",X"6C",X"09",X"CD",X"4A",X"0B",X"CD",X"91",X"09",
		X"3E",X"10",X"CD",X"18",X"09",X"AF",X"CD",X"2C",X"0D",X"3E",X"81",X"32",X"A4",X"80",X"21",X"68",
		X"1D",X"22",X"A6",X"80",X"3E",X"03",X"32",X"58",X"80",X"21",X"80",X"11",X"22",X"5A",X"80",X"3E",
		X"01",X"32",X"B8",X"80",X"32",X"B7",X"80",X"32",X"41",X"88",X"21",X"37",X"80",X"11",X"79",X"80",
		X"0E",X"27",X"ED",X"B0",X"C3",X"09",X"05",X"CD",X"26",X"09",X"CD",X"6C",X"09",X"CD",X"53",X"09",
		X"CD",X"C4",X"09",X"CD",X"FF",X"08",X"E5",X"D1",X"CD",X"48",X"08",X"47",X"BE",X"38",X"2E",X"20",
		X"10",X"3A",X"80",X"88",X"23",X"BE",X"38",X"25",X"20",X"07",X"3A",X"40",X"88",X"23",X"BE",X"38",
		X"1C",X"3A",X"B8",X"80",X"1B",X"12",X"13",X"78",X"12",X"3A",X"80",X"88",X"13",X"12",X"3A",X"40",
		X"88",X"13",X"12",X"3E",X"05",X"CD",X"2C",X"0D",X"3E",X"07",X"CD",X"C6",X"09",X"21",X"40",X"88",
		X"11",X"F1",X"88",X"01",X"20",X"00",X"3E",X"0C",X"F5",X"7E",X"12",X"09",X"EB",X"F1",X"FE",X"08",
		X"20",X"03",X"09",X"09",X"09",X"09",X"EB",X"3D",X"20",X"EE",X"21",X"53",X"8B",X"FD",X"21",X"04",
		X"10",X"06",X"14",X"CD",X"3D",X"0B",X"21",X"74",X"89",X"06",X"05",X"CD",X"3D",X"0B",X"AF",X"32",
		X"F6",X"88",X"32",X"16",X"89",X"3A",X"A0",X"88",X"32",X"76",X"89",X"3A",X"80",X"88",X"32",X"56",
		X"89",X"3A",X"40",X"88",X"32",X"36",X"89",X"21",X"58",X"80",X"34",X"2A",X"5A",X"80",X"23",X"23",
		X"7E",X"23",X"66",X"6F",X"22",X"5A",X"80",X"3E",X"08",X"CD",X"18",X"09",X"21",X"53",X"8B",X"3A",
		X"59",X"80",X"BE",X"28",X"3C",X"34",X"21",X"73",X"89",X"CD",X"19",X"04",X"21",X"76",X"89",X"CD",
		X"19",X"04",X"3E",X"04",X"CD",X"2C",X"0D",X"18",X"DE",X"01",X"00",X"05",X"B7",X"3E",X"05",X"38",
		X"01",X"AF",X"5F",X"7E",X"CB",X"3F",X"F5",X"FE",X"08",X"28",X"08",X"83",X"20",X"09",X"B1",X"3E",
		X"00",X"20",X"04",X"3E",X"10",X"18",X"01",X"0C",X"77",X"11",X"E0",X"FF",X"19",X"F1",X"10",X"DD",
		X"C9",X"21",X"79",X"89",X"FD",X"21",X"18",X"10",X"06",X"05",X"CD",X"3D",X"0B",X"21",X"B6",X"89",
		X"06",X"07",X"7E",X"11",X"05",X"00",X"19",X"77",X"11",X"DB",X"FF",X"19",X"10",X"F4",X"21",X"18",
		X"8A",X"FD",X"21",X"95",X"10",X"11",X"0A",X"00",X"43",X"3A",X"77",X"80",X"32",X"31",X"90",X"D6",
		X"04",X"F5",X"28",X"04",X"30",X"04",X"FD",X"19",X"FD",X"19",X"CD",X"3D",X"0B",X"F1",X"3C",X"F5",
		X"06",X"07",X"21",X"FB",X"88",X"F5",X"7E",X"FE",X"10",X"20",X"01",X"AF",X"5F",X"F1",X"7B",X"8F",
		X"D6",X"0A",X"30",X"02",X"C6",X"0A",X"77",X"3F",X"F5",X"11",X"20",X"00",X"19",X"10",X"E7",X"F1",
		X"F1",X"D6",X"01",X"30",X"DA",X"21",X"BB",X"89",X"01",X"00",X"07",X"CD",X"1C",X"04",X"3E",X"0A",
		X"CD",X"18",X"09",X"26",X"8A",X"3A",X"B8",X"80",X"C6",X"3F",X"6F",X"11",X"FB",X"88",X"06",X"07",
		X"F5",X"1A",X"FE",X"10",X"20",X"01",X"AF",X"4F",X"F1",X"79",X"8E",X"FE",X"0A",X"38",X"02",X"D6",
		X"0A",X"3F",X"77",X"F5",X"C5",X"01",X"20",X"00",X"09",X"EB",X"09",X"EB",X"C1",X"10",X"E2",X"F1",
		X"11",X"E0",X"FF",X"19",X"11",X"02",X"8B",X"06",X"07",X"1A",X"BE",X"38",X"0F",X"20",X"1A",X"C5",
		X"01",X"E0",X"FF",X"09",X"EB",X"09",X"EB",X"C1",X"10",X"EF",X"18",X"0D",X"7E",X"12",X"C5",X"01",
		X"E0",X"FF",X"09",X"EB",X"09",X"EB",X"C1",X"10",X"F3",X"3E",X"FF",X"32",X"59",X"80",X"3A",X"58",
		X"80",X"B7",X"CA",X"BE",X"05",X"E6",X"03",X"C2",X"BE",X"05",X"CD",X"70",X"0A",X"BB",X"20",X"05",
		X"7E",X"FE",X"0E",X"28",X"35",X"3E",X"04",X"CD",X"54",X"09",X"21",X"70",X"80",X"35",X"3A",X"A4",
		X"80",X"87",X"28",X"0B",X"3E",X"84",X"32",X"A4",X"80",X"21",X"8D",X"1D",X"22",X"A6",X"80",X"C3",
		X"C0",X"17",X"21",X"70",X"80",X"34",X"CD",X"26",X"09",X"3A",X"A4",X"80",X"87",X"28",X"0B",X"3E",
		X"82",X"32",X"A4",X"80",X"21",X"E9",X"1D",X"22",X"A6",X"80",X"3A",X"58",X"80",X"E6",X"0F",X"28",
		X"08",X"E6",X"07",X"20",X"59",X"21",X"41",X"88",X"34",X"21",X"57",X"80",X"3A",X"02",X"98",X"E6",
		X"02",X"C6",X"04",X"86",X"77",X"18",X"47",X"CD",X"0C",X"1E",X"CD",X"26",X"09",X"21",X"41",X"88",
		X"35",X"3A",X"A8",X"80",X"CB",X"3F",X"28",X"31",X"7E",X"B7",X"FD",X"21",X"57",X"10",X"21",X"44",
		X"8B",X"06",X"11",X"CC",X"0F",X"09",X"CD",X"08",X"0D",X"7E",X"B7",X"28",X"19",X"FD",X"21",X"68",
		X"10",X"21",X"44",X"8B",X"06",X"09",X"CD",X"3D",X"0B",X"FD",X"21",X"60",X"10",X"06",X"08",X"CD",
		X"0F",X"09",X"3A",X"41",X"88",X"B7",X"CC",X"08",X"0D",X"7E",X"B7",X"CA",X"D8",X"01",X"31",X"00",
		X"88",X"21",X"A4",X"80",X"CB",X"FE",X"CD",X"6C",X"09",X"21",X"4C",X"0D",X"11",X"19",X"80",X"01",
		X"1C",X"00",X"ED",X"B0",X"21",X"00",X"90",X"3A",X"58",X"80",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",
		X"06",X"03",X"71",X"23",X"77",X"23",X"10",X"FA",X"5F",X"CD",X"53",X"09",X"77",X"23",X"73",X"21",
		X"D3",X"10",X"11",X"00",X"80",X"0E",X"10",X"ED",X"B0",X"2A",X"5A",X"80",X"3A",X"A4",X"80",X"87",
		X"3A",X"57",X"80",X"20",X"07",X"5F",X"3A",X"02",X"98",X"E6",X"04",X"83",X"86",X"32",X"60",X"80",
		X"23",X"7E",X"CE",X"00",X"32",X"61",X"80",X"23",X"23",X"23",X"11",X"62",X"80",X"01",X"07",X"00",
		X"ED",X"B0",X"E5",X"0E",X"05",X"ED",X"B0",X"3A",X"6C",X"80",X"32",X"1F",X"80",X"CD",X"7F",X"17",
		X"3A",X"6D",X"80",X"32",X"25",X"80",X"22",X"35",X"80",X"21",X"59",X"80",X"34",X"28",X"07",X"3A",
		X"A8",X"80",X"FE",X"02",X"20",X"29",X"3E",X"02",X"CD",X"2C",X"0D",X"21",X"44",X"8B",X"FD",X"21",
		X"74",X"0F",X"06",X"07",X"CD",X"3D",X"0B",X"3A",X"58",X"80",X"3C",X"CD",X"03",X"0B",X"06",X"08",
		X"FD",X"21",X"71",X"10",X"CD",X"3D",X"0B",X"CD",X"C4",X"09",X"3E",X"06",X"CD",X"18",X"09",X"3A",
		X"02",X"98",X"E6",X"04",X"47",X"3A",X"58",X"80",X"E6",X"F8",X"0F",X"80",X"0F",X"0F",X"FE",X"03",
		X"38",X"02",X"3E",X"02",X"87",X"57",X"3A",X"63",X"80",X"92",X"30",X"02",X"C6",X"0A",X"32",X"80",
		X"88",X"3A",X"62",X"80",X"DE",X"00",X"32",X"A0",X"88",X"AF",X"32",X"40",X"88",X"CD",X"6C",X"09",
		X"3A",X"58",X"80",X"CD",X"54",X"09",X"E1",X"E5",X"11",X"28",X"80",X"0E",X"03",X"ED",X"B0",X"E1",
		X"7E",X"23",X"5E",X"23",X"56",X"23",X"E5",X"21",X"00",X"00",X"18",X"13",X"C1",X"21",X"00",X"00",
		X"B7",X"ED",X"42",X"FA",X"CB",X"06",X"01",X"20",X"00",X"18",X"03",X"01",X"E0",X"FF",X"09",X"E5",
		X"19",X"36",X"2B",X"EB",X"3D",X"20",X"E5",X"C1",X"E1",X"23",X"23",X"7E",X"B7",X"20",X"D2",X"21",
		X"1F",X"88",X"11",X"20",X"00",X"43",X"36",X"2B",X"19",X"10",X"FB",X"3A",X"68",X"80",X"C6",X"14",
		X"87",X"CB",X"10",X"87",X"CB",X"10",X"4F",X"ED",X"42",X"06",X"05",X"36",X"10",X"19",X"10",X"FB",
		X"3E",X"05",X"21",X"76",X"80",X"77",X"23",X"77",X"3C",X"CD",X"2C",X"0D",X"AF",X"32",X"73",X"80",
		X"32",X"72",X"80",X"32",X"C9",X"80",X"32",X"CA",X"80",X"32",X"CC",X"80",X"21",X"11",X"80",X"77",
		X"2B",X"36",X"04",X"11",X"12",X"80",X"0E",X"06",X"ED",X"B0",X"EB",X"77",X"3D",X"32",X"71",X"80",
		X"21",X"A4",X"80",X"CB",X"BE",X"21",X"18",X"80",X"3A",X"72",X"80",X"B7",X"C2",X"77",X"05",X"3A",
		X"A4",X"80",X"CD",X"2C",X"09",X"CB",X"66",X"C4",X"50",X"08",X"CB",X"6E",X"C4",X"D0",X"07",X"CB",
		X"76",X"C4",X"7E",X"07",X"CB",X"7E",X"C4",X"D5",X"08",X"18",X"DD",X"21",X"A4",X"80",X"7E",X"B7",
		X"3A",X"C1",X"80",X"28",X"17",X"35",X"20",X"0F",X"36",X"04",X"23",X"23",X"5E",X"23",X"56",X"1A",
		X"13",X"72",X"2B",X"73",X"2B",X"77",X"2B",X"23",X"7E",X"0F",X"0F",X"77",X"47",X"C9",X"CD",X"5B",
		X"07",X"11",X"04",X"11",X"21",X"2B",X"80",X"4E",X"69",X"26",X"00",X"19",X"5E",X"7B",X"CB",X"60",
		X"28",X"09",X"23",X"0C",X"7E",X"B7",X"F2",X"B3",X"07",X"18",X"21",X"CB",X"68",X"28",X"09",X"2B",
		X"0D",X"7E",X"B7",X"F2",X"B3",X"07",X"18",X"14",X"B7",X"28",X"11",X"FE",X"06",X"30",X"03",X"0D",
		X"18",X"01",X"0C",X"21",X"2B",X"80",X"3E",X"FF",X"32",X"C9",X"80",X"71",X"7B",X"32",X"27",X"80",
		X"AF",X"32",X"C9",X"80",X"2A",X"31",X"80",X"22",X"14",X"80",X"21",X"18",X"80",X"CB",X"B6",X"C9",
		X"3A",X"C8",X"80",X"B7",X"28",X"66",X"DD",X"21",X"00",X"80",X"3A",X"19",X"80",X"47",X"17",X"3E",
		X"FF",X"32",X"CA",X"80",X"DD",X"7E",X"01",X"30",X"0A",X"FE",X"30",X"28",X"0E",X"FE",X"F3",X"28",
		X"0A",X"18",X"29",X"FE",X"3C",X"28",X"04",X"FE",X"FF",X"20",X"21",X"EE",X"CC",X"DD",X"4E",X"0D",
		X"DD",X"77",X"0D",X"3E",X"CC",X"A9",X"DD",X"77",X"01",X"DD",X"7E",X"05",X"EE",X"CC",X"DD",X"4E",
		X"09",X"DD",X"77",X"09",X"3E",X"CC",X"A9",X"DD",X"77",X"05",X"18",X"1C",X"DD",X"7E",X"01",X"80",
		X"DD",X"77",X"01",X"DD",X"7E",X"05",X"80",X"DD",X"77",X"05",X"DD",X"7E",X"09",X"80",X"DD",X"77",
		X"09",X"DD",X"7E",X"0D",X"80",X"DD",X"77",X"0D",X"AF",X"32",X"CA",X"80",X"2A",X"2F",X"80",X"22",
		X"12",X"80",X"21",X"18",X"80",X"CB",X"AE",X"C9",X"3A",X"A0",X"88",X"FE",X"10",X"C0",X"AF",X"C9",
		X"3A",X"40",X"88",X"3D",X"F2",X"C6",X"08",X"CD",X"48",X"08",X"67",X"3A",X"80",X"88",X"6F",X"ED",
		X"5B",X"64",X"80",X"E5",X"37",X"9B",X"30",X"02",X"C6",X"0A",X"6F",X"7C",X"9A",X"67",X"F2",X"88",
		X"08",X"E1",X"E5",X"ED",X"5B",X"66",X"80",X"37",X"7D",X"9B",X"30",X"02",X"C6",X"0A",X"6F",X"7C",
		X"9A",X"67",X"F2",X"88",X"08",X"E1",X"E5",X"37",X"7D",X"DE",X"02",X"7C",X"DE",X"00",X"F2",X"9A",
		X"08",X"3A",X"77",X"80",X"3D",X"32",X"76",X"80",X"18",X"06",X"3A",X"76",X"80",X"32",X"77",X"80",
		X"E1",X"3A",X"80",X"88",X"3D",X"F2",X"C1",X"08",X"3A",X"A0",X"88",X"3D",X"28",X"0C",X"FE",X"0F",
		X"20",X"0A",X"32",X"72",X"80",X"21",X"FF",X"7F",X"18",X"12",X"3E",X"10",X"32",X"A0",X"88",X"3E",
		X"09",X"32",X"80",X"88",X"3E",X"09",X"32",X"40",X"88",X"2A",X"2D",X"80",X"22",X"10",X"80",X"21",
		X"18",X"80",X"CB",X"A6",X"C9",X"DD",X"21",X"00",X"80",X"21",X"78",X"80",X"CB",X"06",X"2A",X"33",
		X"80",X"3A",X"76",X"80",X"38",X"04",X"3A",X"77",X"80",X"29",X"DD",X"77",X"02",X"DD",X"77",X"06",
		X"DD",X"77",X"0A",X"DD",X"77",X"0E",X"22",X"16",X"80",X"21",X"18",X"80",X"CB",X"BE",X"C9",X"3A",
		X"58",X"80",X"6F",X"26",X"00",X"4D",X"44",X"29",X"09",X"29",X"01",X"58",X"81",X"09",X"C9",X"CD",
		X"3D",X"0B",X"3A",X"B8",X"80",X"77",X"3E",X"08",X"10",X"FE",X"0D",X"20",X"FB",X"F5",X"CD",X"26",
		X"09",X"F1",X"3D",X"20",X"F3",X"C9",X"21",X"A4",X"80",X"CB",X"FE",X"7E",X"87",X"C8",X"3A",X"A8",
		X"80",X"B7",X"C8",X"3E",X"80",X"32",X"A4",X"80",X"32",X"75",X"80",X"3E",X"55",X"32",X"CB",X"80",
		X"AF",X"21",X"48",X"90",X"06",X"05",X"77",X"23",X"23",X"23",X"23",X"10",X"F9",X"CD",X"2C",X"0D",
		X"C3",X"26",X"02",X"AF",X"06",X"1C",X"21",X"06",X"90",X"36",X"00",X"23",X"77",X"23",X"10",X"F9",
		X"C9",X"AF",X"06",X"07",X"11",X"20",X"00",X"77",X"19",X"10",X"FC",X"C9",X"11",X"00",X"88",X"3E",
		X"20",X"13",X"13",X"13",X"21",X"01",X"00",X"19",X"EB",X"01",X"1B",X"00",X"36",X"10",X"ED",X"B0",
		X"13",X"3D",X"20",X"ED",X"C9",X"3E",X"10",X"32",X"32",X"81",X"32",X"33",X"81",X"32",X"34",X"81",
		X"C9",X"CD",X"85",X"09",X"E5",X"C5",X"0E",X"0A",X"11",X"CE",X"80",X"21",X"EB",X"8A",X"06",X"03",
		X"CD",X"55",X"0A",X"7D",X"C6",X"C0",X"6F",X"06",X"07",X"CD",X"55",X"0A",X"3E",X"82",X"85",X"6F",
		X"24",X"0D",X"20",X"EA",X"2D",X"06",X"03",X"CD",X"55",X"0A",X"3E",X"01",X"0E",X"50",X"CD",X"18",
		X"09",X"C1",X"E1",X"C9",X"3E",X"01",X"32",X"1D",X"90",X"06",X"1C",X"FD",X"21",X"79",X"10",X"21",
		X"A7",X"8B",X"CD",X"3D",X"0B",X"21",X"69",X"89",X"06",X"05",X"CD",X"7B",X"0B",X"21",X"6A",X"89",
		X"06",X"04",X"CD",X"7B",X"0B",X"21",X"6B",X"89",X"06",X"03",X"CD",X"7B",X"0B",X"21",X"AE",X"8B",
		X"06",X"11",X"CD",X"3D",X"0B",X"21",X"09",X"8A",X"3E",X"0C",X"77",X"2C",X"77",X"2C",X"77",X"21",
		X"E9",X"89",X"AF",X"77",X"2C",X"77",X"2C",X"77",X"32",X"2B",X"8A",X"21",X"29",X"8A",X"ED",X"4B",
		X"64",X"80",X"CD",X"63",X"0A",X"21",X"2A",X"8A",X"ED",X"4B",X"66",X"80",X"CD",X"63",X"0A",X"CD",
		X"FF",X"08",X"23",X"23",X"7E",X"32",X"4E",X"88",X"3E",X"0C",X"32",X"6E",X"88",X"2B",X"7E",X"32",
		X"8E",X"88",X"2B",X"7E",X"B7",X"20",X"02",X"3E",X"10",X"32",X"AE",X"88",X"2B",X"EB",X"1A",X"FE",
		X"03",X"30",X"03",X"11",X"C6",X"10",X"1B",X"1B",X"06",X"03",X"21",X"2E",X"89",X"CD",X"55",X"0A",
		X"3E",X"08",X"C3",X"18",X"09",X"1A",X"77",X"13",X"3E",X"E0",X"85",X"6F",X"3E",X"FF",X"8C",X"67",
		X"10",X"F3",X"C9",X"11",X"20",X"00",X"71",X"78",X"B7",X"20",X"02",X"06",X"10",X"19",X"70",X"C9",
		X"21",X"3B",X"80",X"11",X"05",X"00",X"43",X"AF",X"4E",X"CB",X"11",X"CE",X"00",X"19",X"10",X"F8",
		X"C9",X"CD",X"08",X"0D",X"3A",X"58",X"80",X"21",X"B5",X"80",X"BE",X"38",X"01",X"77",X"CD",X"F1",
		X"0A",X"21",X"AE",X"80",X"CD",X"D0",X"0A",X"CD",X"70",X"0A",X"21",X"B1",X"80",X"CD",X"CF",X"0A",
		X"21",X"B6",X"80",X"BE",X"38",X"01",X"77",X"FE",X"05",X"C0",X"CD",X"2C",X"0D",X"FD",X"21",X"83",
		X"0E",X"06",X"09",X"21",X"63",X"8A",X"CD",X"3D",X"0B",X"21",X"BB",X"80",X"3E",X"01",X"86",X"27",
		X"30",X"02",X"3E",X"99",X"77",X"3E",X"08",X"CD",X"18",X"09",X"21",X"B4",X"80",X"3E",X"01",X"48",
		X"F5",X"07",X"07",X"07",X"07",X"CB",X"38",X"1F",X"CB",X"38",X"1F",X"CB",X"38",X"1F",X"CB",X"38",
		X"1F",X"86",X"27",X"77",X"2B",X"7E",X"89",X"27",X"77",X"2B",X"7E",X"CE",X"00",X"27",X"77",X"F1",
		X"C9",X"01",X"FF",X"FF",X"0C",X"D6",X"64",X"30",X"FB",X"C6",X"64",X"04",X"D6",X"0A",X"30",X"FB",
		X"C6",X"0A",X"C9",X"CD",X"F1",X"0A",X"11",X"E0",X"FF",X"71",X"19",X"70",X"19",X"77",X"19",X"C9",
		X"DD",X"7E",X"00",X"DD",X"23",X"CD",X"03",X"0B",X"18",X"20",X"4F",X"CB",X"3F",X"CB",X"3F",X"CB",
		X"3F",X"CB",X"3F",X"77",X"79",X"E6",X"0F",X"19",X"77",X"C9",X"06",X"03",X"11",X"E0",X"FF",X"DD",
		X"7E",X"00",X"DD",X"23",X"CD",X"1A",X"0B",X"19",X"10",X"F5",X"19",X"06",X"0C",X"11",X"E0",X"FF",
		X"FD",X"7E",X"00",X"77",X"19",X"FD",X"23",X"10",X"F7",X"C9",X"3E",X"05",X"32",X"09",X"90",X"32",
		X"0D",X"90",X"32",X"11",X"90",X"32",X"13",X"90",X"21",X"C4",X"8A",X"06",X"0A",X"FD",X"21",X"68",
		X"0D",X"CD",X"3D",X"0B",X"06",X"17",X"21",X"A6",X"8B",X"CD",X"3D",X"0B",X"06",X"18",X"21",X"A8",
		X"8B",X"CD",X"3D",X"0B",X"06",X"1C",X"21",X"A9",X"8B",X"18",X"C2",X"3E",X"1D",X"90",X"90",X"4F",
		X"78",X"06",X"90",X"02",X"01",X"07",X"00",X"FD",X"09",X"06",X"03",X"18",X"B0",X"7D",X"E6",X"1F",
		X"87",X"5F",X"16",X"00",X"DD",X"21",X"00",X"90",X"DD",X"19",X"DD",X"36",X"00",X"E0",X"0E",X"1C",
		X"11",X"DF",X"00",X"ED",X"53",X"12",X"80",X"11",X"E0",X"FF",X"FD",X"7E",X"00",X"77",X"C5",X"3A",
		X"12",X"80",X"47",X"DD",X"77",X"00",X"CD",X"2E",X"09",X"3A",X"12",X"80",X"B8",X"28",X"F7",X"3E",
		X"07",X"A0",X"20",X"EB",X"C1",X"19",X"FD",X"23",X"0D",X"10",X"DF",X"FD",X"2B",X"06",X"01",X"20",
		X"DD",X"11",X"81",X"03",X"19",X"FD",X"23",X"C9",X"21",X"51",X"81",X"3A",X"58",X"80",X"47",X"04",
		X"3A",X"B8",X"80",X"23",X"23",X"23",X"23",X"23",X"23",X"BE",X"C8",X"10",X"F6",X"C9",X"7E",X"12",
		X"1B",X"7D",X"C6",X"20",X"6F",X"30",X"01",X"24",X"10",X"F4",X"C9",X"0E",X"09",X"CD",X"85",X"09",
		X"11",X"D1",X"80",X"06",X"07",X"26",X"8B",X"3A",X"B8",X"80",X"3D",X"6F",X"1A",X"BE",X"38",X"22",
		X"20",X"0B",X"13",X"3E",X"E0",X"85",X"6F",X"3E",X"FF",X"8C",X"67",X"10",X"EF",X"78",X"C6",X"03",
		X"83",X"5F",X"30",X"01",X"14",X"0D",X"F2",X"03",X"0C",X"CD",X"D8",X"0B",X"C0",X"11",X"34",X"81",
		X"18",X"20",X"AF",X"B1",X"11",X"31",X"81",X"28",X"0C",X"87",X"87",X"81",X"87",X"4F",X"06",X"00",
		X"21",X"27",X"81",X"ED",X"B8",X"06",X"07",X"26",X"8A",X"3A",X"B8",X"80",X"C6",X"3F",X"6F",X"CD",
		X"EE",X"0B",X"D5",X"CD",X"6C",X"09",X"32",X"4C",X"90",X"32",X"50",X"90",X"32",X"54",X"90",X"32",
		X"58",X"90",X"FD",X"21",X"1D",X"10",X"21",X"A4",X"8B",X"06",X"0F",X"CD",X"3D",X"0B",X"06",X"08",
		X"FD",X"E5",X"FD",X"21",X"60",X"10",X"CD",X"3D",X"0B",X"FD",X"E1",X"3A",X"B8",X"80",X"77",X"21",
		X"46",X"8B",X"06",X"15",X"CD",X"3D",X"0B",X"21",X"47",X"8B",X"06",X"16",X"CD",X"3D",X"0B",X"E1",
		X"CD",X"B1",X"0C",X"F2",X"99",X"0C",X"23",X"10",X"FD",X"2B",X"11",X"34",X"81",X"01",X"03",X"00",
		X"ED",X"B8",X"CD",X"D8",X"0B",X"C0",X"EB",X"21",X"34",X"81",X"01",X"03",X"00",X"ED",X"B8",X"18",
		X"F1",X"36",X"10",X"2B",X"36",X"10",X"2B",X"06",X"03",X"36",X"0A",X"11",X"84",X"03",X"ED",X"53",
		X"10",X"80",X"CD",X"94",X"09",X"3A",X"11",X"80",X"B7",X"F8",X"3A",X"C1",X"80",X"CB",X"67",X"28",
		X"0E",X"7E",X"3C",X"FE",X"2B",X"30",X"16",X"FE",X"0B",X"20",X"14",X"3E",X"11",X"18",X"10",X"CB",
		X"6F",X"28",X"0F",X"7E",X"3D",X"FE",X"10",X"30",X"06",X"3E",X"2A",X"18",X"02",X"3E",X"10",X"77",
		X"18",X"D0",X"E6",X"0A",X"28",X"CC",X"7E",X"FE",X"0A",X"20",X"02",X"36",X"10",X"3A",X"C1",X"80",
		X"E6",X"0A",X"20",X"F9",X"23",X"10",X"B2",X"C9",X"21",X"37",X"80",X"11",X"79",X"80",X"06",X"2B",
		X"1A",X"4E",X"77",X"79",X"12",X"23",X"13",X"10",X"F7",X"21",X"B8",X"80",X"3E",X"03",X"AE",X"77",
		X"21",X"41",X"88",X"46",X"11",X"B7",X"80",X"1A",X"77",X"78",X"12",X"C9",X"32",X"CD",X"80",X"F5",
		X"3A",X"75",X"80",X"B7",X"28",X"04",X"F1",X"C6",X"07",X"F5",X"F1",X"F3",X"32",X"00",X"A0",X"AF",
		X"32",X"01",X"A0",X"E3",X"E3",X"3E",X"08",X"32",X"01",X"A0",X"FB",X"C9",X"04",X"00",X"00",X"00",
		X"00",X"00",X"6C",X"00",X"00",X"00",X"00",X"00",X"1F",X"00",X"00",X"11",X"48",X"8A",X"06",X"00",
		X"03",X"00",X"09",X"00",X"02",X"00",X"02",X"00",X"23",X"20",X"15",X"15",X"14",X"10",X"13",X"1F",
		X"19",X"1E",X"0B",X"01",X"09",X"08",X"04",X"10",X"23",X"24",X"15",X"22",X"1E",X"10",X"15",X"1C",
		X"15",X"13",X"24",X"22",X"1F",X"1E",X"19",X"13",X"23",X"20",X"22",X"1F",X"17",X"22",X"11",X"1D",
		X"1D",X"15",X"14",X"10",X"12",X"29",X"10",X"1B",X"15",X"19",X"24",X"18",X"10",X"15",X"1E",X"17",
		X"15",X"17",X"11",X"1D",X"15",X"10",X"13",X"1F",X"1E",X"13",X"15",X"20",X"24",X"10",X"12",X"29",
		X"10",X"24",X"18",X"1F",X"1D",X"11",X"23",X"10",X"12",X"11",X"22",X"1F",X"1E",X"11",X"16",X"24",
		X"15",X"22",X"10",X"15",X"26",X"15",X"22",X"29",X"10",X"16",X"1F",X"25",X"22",X"24",X"18",X"10",
		X"23",X"13",X"22",X"15",X"15",X"1E",X"10",X"19",X"23",X"11",X"10",X"12",X"1F",X"1E",X"25",X"23",
		X"10",X"23",X"13",X"22",X"15",X"15",X"1E",X"10",X"14",X"25",X"22",X"19",X"1E",X"17",X"10",X"27",
		X"18",X"19",X"13",X"18",X"1E",X"1F",X"10",X"13",X"1F",X"19",X"1E",X"23",X"10",X"13",X"11",X"1E",
		X"10",X"12",X"15",X"10",X"1C",X"1F",X"23",X"24",X"0C",X"24",X"18",X"15",X"10",X"1A",X"1F",X"29",
		X"23",X"24",X"19",X"13",X"1B",X"10",X"14",X"19",X"22",X"15",X"13",X"24",X"23",X"10",X"24",X"18",
		X"15",X"12",X"11",X"1C",X"1C",X"10",X"12",X"29",X"10",X"23",X"1C",X"19",X"14",X"19",X"1E",X"17",
		X"10",X"24",X"18",X"15",X"10",X"23",X"24",X"19",X"13",X"1B",X"23",X"1F",X"25",X"24",X"10",X"1F",
		X"16",X"10",X"19",X"24",X"23",X"10",X"20",X"11",X"24",X"18",X"0C",X"11",X"10",X"12",X"1F",X"1E",
		X"25",X"23",X"10",X"13",X"1F",X"19",X"1E",X"10",X"19",X"23",X"10",X"11",X"27",X"11",X"22",X"14",
		X"15",X"14",X"10",X"16",X"1F",X"22",X"24",X"18",X"15",X"10",X"12",X"11",X"1C",X"1C",X"10",X"18",
		X"19",X"24",X"24",X"19",X"1E",X"17",X"10",X"13",X"1F",X"19",X"1E",X"10",X"27",X"1F",X"22",X"14",
		X"0C",X"11",X"10",X"16",X"22",X"15",X"15",X"10",X"20",X"1C",X"11",X"29",X"10",X"19",X"23",X"10",
		X"11",X"27",X"11",X"22",X"14",X"15",X"14",X"10",X"16",X"1F",X"22",X"15",X"26",X"15",X"1E",X"24",
		X"25",X"11",X"1C",X"1C",X"29",X"10",X"23",X"20",X"15",X"1C",X"1C",X"19",X"1E",X"17",X"10",X"23",
		X"24",X"15",X"22",X"1E",X"0C",X"24",X"18",X"15",X"10",X"16",X"1F",X"22",X"13",X"15",X"10",X"1F",
		X"16",X"10",X"17",X"22",X"11",X"26",X"19",X"24",X"29",X"10",X"19",X"23",X"19",X"1E",X"13",X"22",
		X"15",X"11",X"23",X"15",X"14",X"10",X"11",X"16",X"24",X"15",X"22",X"10",X"15",X"26",X"15",X"22",
		X"29",X"10",X"02",X"1E",X"14",X"12",X"1F",X"1E",X"25",X"23",X"10",X"23",X"13",X"22",X"15",X"15",
		X"1E",X"0C",X"11",X"10",X"12",X"1F",X"1E",X"25",X"23",X"10",X"13",X"1F",X"19",X"1E",X"10",X"19",
		X"23",X"10",X"11",X"27",X"11",X"22",X"14",X"15",X"14",X"11",X"16",X"24",X"15",X"22",X"10",X"24",
		X"18",X"15",X"10",X"02",X"1E",X"14",X"10",X"12",X"1F",X"1E",X"25",X"23",X"10",X"23",X"13",X"22",
		X"15",X"15",X"1E",X"11",X"1E",X"14",X"10",X"15",X"26",X"15",X"22",X"29",X"10",X"04",X"24",X"18",
		X"10",X"1F",X"1E",X"15",X"10",X"24",X"18",X"15",X"22",X"15",X"11",X"16",X"24",X"15",X"22",X"17",
		X"11",X"1D",X"15",X"23",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"23",X"13",X"22",X"15",X"15",
		X"1E",X"23",X"10",X"10",X"10",X"10",X"10",X"1C",X"15",X"24",X"24",X"15",X"22",X"23",X"10",X"10",
		X"10",X"10",X"10",X"16",X"22",X"15",X"15",X"10",X"17",X"11",X"1D",X"15",X"23",X"10",X"10",X"12",
		X"15",X"23",X"24",X"10",X"23",X"13",X"22",X"15",X"15",X"1E",X"10",X"12",X"15",X"23",X"24",X"10",
		X"1C",X"15",X"24",X"24",X"15",X"22",X"23",X"25",X"22",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"0E",X"0F",X"10",X"23",X"10",X"84",X"0F",X"10",X"24",X"10",X"84",X"0F",X"10",X"15",
		X"10",X"84",X"0F",X"10",X"22",X"10",X"84",X"0F",X"10",X"1E",X"10",X"84",X"0F",X"8A",X"8B",X"0E",
		X"0E",X"00",X"00",X"FF",X"11",X"11",X"23",X"19",X"01",X"23",X"24",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"0E",X"0E",X"10",X"23",X"15",X"13",X"1F",X"1E",X"14",X"23",X"10",
		X"10",X"10",X"0C",X"02",X"1E",X"14",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"0E",X"0E",X"10",X"13",X"1F",X"19",X"1E",X"23",X"10",X"1C",X"15",X"16",X"24",X"18",X"19",X"17",
		X"18",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"0E",X"0E",X"10",X"13",X"22",X"15",
		X"14",X"19",X"24",X"23",X"00",X"10",X"13",X"1F",X"19",X"1E",X"23",X"10",X"1C",X"1F",X"23",X"24",
		X"10",X"10",X"28",X"10",X"01",X"00",X"00",X"00",X"0A",X"0A",X"0A",X"0A",X"0A",X"13",X"1F",X"1E",
		X"17",X"22",X"11",X"24",X"25",X"1C",X"11",X"24",X"19",X"1F",X"1E",X"23",X"23",X"24",X"19",X"13",
		X"1B",X"10",X"13",X"18",X"11",X"1E",X"17",X"15",X"23",X"10",X"19",X"1E",X"19",X"24",X"19",X"11",
		X"1C",X"12",X"25",X"24",X"24",X"1F",X"1E",X"10",X"23",X"15",X"1C",X"15",X"13",X"24",X"23",X"10",
		X"19",X"1E",X"19",X"24",X"19",X"11",X"1C",X"17",X"11",X"1D",X"15",X"10",X"1F",X"26",X"15",X"22",
		X"10",X"20",X"1C",X"11",X"29",X"15",X"22",X"10",X"17",X"15",X"24",X"10",X"22",X"15",X"11",X"14",
		X"29",X"10",X"19",X"23",X"10",X"1E",X"15",X"28",X"24",X"24",X"19",X"1D",X"15",X"10",X"1C",X"15",
		X"16",X"24",X"10",X"11",X"12",X"1F",X"26",X"15",X"10",X"10",X"10",X"1D",X"25",X"1C",X"24",X"19",
		X"20",X"1C",X"19",X"15",X"22",X"27",X"18",X"19",X"24",X"15",X"10",X"10",X"28",X"10",X"04",X"10",
		X"12",X"1C",X"25",X"15",X"10",X"10",X"28",X"10",X"02",X"10",X"10",X"22",X"15",X"14",X"10",X"10",
		X"28",X"10",X"01",X"13",X"25",X"22",X"22",X"15",X"1E",X"24",X"10",X"12",X"15",X"23",X"24",X"10",
		X"24",X"19",X"1D",X"15",X"1E",X"15",X"27",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"00",X"00",X"30",X"05",X"1F",X"00",X"31",X"05",X"2F",X"00",X"32",X"05",X"1F",X"00",
		X"33",X"05",X"2F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"0A",X"09",X"08",X"07",X"06",X"00",X"01",X"02",X"03",X"04",X"05",
		X"FF",X"07",X"00",X"36",X"11",X"03",X"00",X"05",X"01",X"01",X"01",X"A4",X"11",X"68",X"8A",X"64",
		X"1F",X"11",X"8D",X"89",X"9C",X"47",X"11",X"72",X"8A",X"64",X"6F",X"11",X"97",X"89",X"9C",X"97",
		X"0D",X"9C",X"8A",X"5C",X"BF",X"00",X"07",X"00",X"5B",X"11",X"02",X"05",X"01",X"01",X"08",X"00",
		X"B4",X"0D",X"48",X"8A",X"6C",X"1F",X"0D",X"AD",X"89",X"94",X"47",X"0D",X"52",X"8A",X"6C",X"6F",
		X"0D",X"B7",X"89",X"94",X"97",X"0D",X"5C",X"8A",X"6C",X"BF",X"00",X"07",X"00",X"80",X"11",X"02",
		X"00",X"00",X"01",X"07",X"00",X"94",X"05",X"48",X"8A",X"6C",X"1F",X"05",X"AD",X"89",X"94",X"47",
		X"05",X"52",X"8A",X"6C",X"6F",X"05",X"B7",X"89",X"94",X"97",X"05",X"5C",X"8A",X"6C",X"BF",X"00",
		X"07",X"00",X"A5",X"11",X"02",X"00",X"01",X"01",X"08",X"00",X"D4",X"11",X"48",X"8A",X"6C",X"1F",
		X"0D",X"8D",X"89",X"9C",X"47",X"0B",X"52",X"8A",X"6C",X"6F",X"05",X"17",X"8B",X"3C",X"97",X"09",
		X"DC",X"89",X"8C",X"BF",X"00",X"07",X"00",X"CA",X"11",X"02",X"00",X"04",X"01",X"01",X"01",X"9C",
		X"05",X"88",X"8A",X"5C",X"1F",X"0D",X"6C",X"8A",X"64",X"3F",X"05",X"F0",X"88",X"C4",X"5F",X"05",
		X"F2",X"89",X"84",X"6F",X"05",X"96",X"8A",X"5C",X"8F",X"00",X"07",X"00",X"F9",X"11",X"02",X"05",
		X"05",X"01",X"02",X"01",X"A4",X"09",X"48",X"8A",X"6C",X"1F",X"05",X"2A",X"89",X"B4",X"2F",X"0D",
		X"AE",X"89",X"94",X"4F",X"05",X"10",X"8B",X"3C",X"5F",X"0D",X"75",X"89",X"A4",X"87",X"05",X"18",
		X"8B",X"3C",X"9F",X"03",X"FC",X"89",X"84",X"BF",X"00",X"07",X"00",X"23",X"12",X"02",X"08",X"03",
		X"02",X"09",X"01",X"74",X"09",X"A8",X"8A",X"54",X"1F",X"05",X"4B",X"89",X"AC",X"37",X"05",X"4E",
		X"8A",X"6C",X"4F",X"03",X"30",X"8B",X"34",X"5F",X"05",X"54",X"8A",X"6C",X"7F",X"05",X"38",X"89",
		X"B4",X"9F",X"00",X"07",X"00",X"11",X"11",X"02",X"08",X"01",X"02",X"02",X"01",X"3C",X"09",X"E8",
		X"8A",X"44",X"1F",X"09",X"0A",X"89",X"BC",X"2F",X"09",X"ED",X"8A",X"44",X"47",X"07",X"10",X"89",
		X"BC",X"5F",X"07",X"15",X"8B",X"3C",X"87",X"03",X"99",X"8A",X"5C",X"A7",X"00",X"08",X"3A",X"00",
		X"B0",X"3A",X"01",X"98",X"E6",X"01",X"20",X"F6",X"D9",X"DD",X"E5",X"32",X"01",X"A8",X"3D",X"32",
		X"01",X"A8",X"3A",X"CB",X"80",X"07",X"32",X"CB",X"80",X"D2",X"02",X"15",X"3A",X"CC",X"80",X"B7",
		X"C2",X"81",X"15",X"3A",X"A4",X"80",X"B7",X"FA",X"A4",X"14",X"3E",X"FF",X"32",X"CC",X"80",X"3A",
		X"70",X"80",X"B7",X"FA",X"86",X"15",X"C2",X"99",X"14",X"3A",X"C9",X"80",X"B7",X"C2",X"A4",X"14",
		X"2A",X"1E",X"80",X"ED",X"5B",X"1C",X"80",X"19",X"22",X"1E",X"80",X"CD",X"7E",X"17",X"FE",X"E0",
		X"38",X"07",X"11",X"00",X"00",X"ED",X"53",X"1C",X"80",X"3A",X"6C",X"80",X"94",X"47",X"F2",X"B3",
		X"12",X"ED",X"44",X"4F",X"2A",X"35",X"80",X"3A",X"2C",X"80",X"B7",X"FA",X"DE",X"12",X"3A",X"69",
		X"80",X"CB",X"3F",X"87",X"87",X"87",X"C6",X"0C",X"91",X"32",X"2C",X"80",X"F2",X"63",X"13",X"7E",
		X"B7",X"CA",X"63",X"13",X"AF",X"32",X"71",X"80",X"32",X"27",X"80",X"C3",X"63",X"13",X"7E",X"B7",
		X"28",X"28",X"3A",X"2B",X"80",X"E6",X"7F",X"6F",X"26",X"00",X"CD",X"11",X"17",X"ED",X"5B",X"1C",
		X"80",X"3A",X"25",X"80",X"BC",X"DA",X"63",X"13",X"3A",X"74",X"80",X"B7",X"28",X"D6",X"AF",X"32",
		X"74",X"80",X"32",X"2C",X"80",X"2A",X"1E",X"80",X"18",X"9F",X"3A",X"73",X"80",X"B7",X"3A",X"25",
		X"80",X"20",X"2A",X"FE",X"DF",X"38",X"CB",X"2A",X"1E",X"80",X"3A",X"68",X"80",X"94",X"F2",X"23",
		X"13",X"ED",X"44",X"FE",X"08",X"30",X"35",X"AF",X"32",X"1C",X"80",X"32",X"1D",X"80",X"3D",X"32",
		X"73",X"80",X"3A",X"68",X"80",X"32",X"1F",X"80",X"CD",X"83",X"17",X"18",X"26",X"FE",X"DF",X"38",
		X"04",X"FE",X"EF",X"38",X"1E",X"AF",X"DD",X"21",X"4C",X"90",X"DD",X"77",X"00",X"DD",X"77",X"04",
		X"DD",X"77",X"08",X"DD",X"77",X"0C",X"32",X"CC",X"80",X"C3",X"57",X"03",X"AF",X"32",X"CC",X"80",
		X"C3",X"77",X"05",X"2A",X"1A",X"80",X"B7",X"ED",X"5A",X"22",X"1C",X"80",X"3E",X"04",X"F2",X"79",
		X"13",X"3E",X"FC",X"EB",X"21",X"00",X"00",X"ED",X"52",X"32",X"19",X"80",X"7C",X"B5",X"32",X"C8",
		X"80",X"28",X"18",X"1E",X"00",X"29",X"38",X"03",X"1C",X"20",X"FA",X"7B",X"87",X"83",X"D6",X"0F",
		X"21",X"01",X"00",X"28",X"03",X"38",X"01",X"6F",X"22",X"2F",X"80",X"3A",X"2C",X"80",X"B7",X"F2",
		X"C8",X"13",X"21",X"00",X"00",X"22",X"1A",X"80",X"2A",X"24",X"80",X"ED",X"5B",X"22",X"80",X"19",
		X"22",X"24",X"80",X"7C",X"2A",X"20",X"80",X"19",X"22",X"22",X"80",X"2A",X"60",X"80",X"29",X"29",
		X"29",X"29",X"22",X"20",X"80",X"C3",X"00",X"14",X"3A",X"2B",X"80",X"E6",X"7F",X"6F",X"26",X"00",
		X"E5",X"11",X"A8",X"17",X"19",X"7E",X"ED",X"5B",X"60",X"80",X"21",X"00",X"00",X"22",X"22",X"80",
		X"22",X"20",X"80",X"B7",X"F2",X"ED",X"13",X"ED",X"52",X"EB",X"21",X"00",X"00",X"E6",X"7F",X"28",
		X"04",X"19",X"3D",X"20",X"FC",X"22",X"1A",X"80",X"E1",X"CD",X"11",X"17",X"22",X"24",X"80",X"7C",
		X"DD",X"77",X"03",X"DD",X"77",X"0B",X"C6",X"10",X"DD",X"77",X"07",X"DD",X"77",X"0F",X"06",X"00",
		X"3A",X"26",X"80",X"87",X"4F",X"21",X"92",X"17",X"09",X"5E",X"23",X"56",X"EB",X"DD",X"2A",X"29",
		X"80",X"3A",X"28",X"80",X"47",X"23",X"5E",X"23",X"56",X"23",X"DD",X"19",X"DD",X"36",X"00",X"10",
		X"7E",X"23",X"B7",X"20",X"F1",X"10",X"EE",X"3A",X"27",X"80",X"32",X"26",X"80",X"87",X"4F",X"21",
		X"92",X"17",X"09",X"5E",X"23",X"56",X"EB",X"DD",X"2A",X"6A",X"80",X"DD",X"22",X"29",X"80",X"3A",
		X"69",X"80",X"32",X"28",X"80",X"47",X"7E",X"23",X"5E",X"23",X"56",X"23",X"DD",X"19",X"DD",X"77",
		X"00",X"7E",X"23",X"B7",X"20",X"F2",X"10",X"EE",X"21",X"71",X"80",X"7E",X"B7",X"20",X"24",X"34",
		X"2A",X"35",X"80",X"7E",X"B7",X"28",X"1C",X"E5",X"11",X"28",X"80",X"01",X"03",X"00",X"ED",X"B0",
		X"E1",X"11",X"69",X"80",X"0E",X"05",X"ED",X"B0",X"22",X"35",X"80",X"3E",X"06",X"32",X"2B",X"80",
		X"32",X"74",X"80",X"3A",X"CA",X"80",X"B7",X"20",X"0B",X"21",X"00",X"80",X"11",X"4C",X"90",X"01",
		X"10",X"00",X"ED",X"B0",X"21",X"10",X"80",X"06",X"04",X"35",X"23",X"20",X"01",X"35",X"4E",X"CB",
		X"11",X"1F",X"23",X"10",X"F4",X"B6",X"77",X"21",X"BF",X"80",X"11",X"00",X"98",X"CD",X"02",X"17",
		X"CD",X"02",X"17",X"CD",X"02",X"17",X"3A",X"A8",X"80",X"B7",X"20",X"36",X"21",X"BB",X"80",X"3A",
		X"01",X"98",X"E6",X"02",X"4F",X"B6",X"28",X"2A",X"3A",X"C1",X"80",X"CB",X"4F",X"20",X"05",X"CB",
		X"5F",X"28",X"1F",X"04",X"04",X"79",X"B7",X"20",X"06",X"7E",X"90",X"27",X"38",X"14",X"77",X"78",
		X"32",X"A8",X"80",X"3E",X"01",X"32",X"B8",X"80",X"7E",X"21",X"62",X"88",X"11",X"E0",X"FF",X"CD",
		X"1A",X"0B",X"21",X"B9",X"80",X"7E",X"23",X"46",X"A8",X"4F",X"3A",X"00",X"98",X"2F",X"E6",X"C0",
		X"77",X"2B",X"70",X"A1",X"23",X"23",X"47",X"AF",X"CB",X"10",X"CE",X"00",X"CB",X"10",X"CE",X"00",
		X"47",X"86",X"27",X"30",X"02",X"3E",X"99",X"77",X"23",X"7E",X"80",X"77",X"78",X"B7",X"2B",X"7E",
		X"11",X"E0",X"FF",X"21",X"62",X"88",X"C4",X"1A",X"0B",X"21",X"BD",X"80",X"7E",X"B7",X"20",X"1F",
		X"2B",X"7E",X"B7",X"28",X"38",X"35",X"23",X"3A",X"CB",X"80",X"3C",X"3E",X"05",X"20",X"01",X"87",
		X"77",X"3E",X"FF",X"32",X"02",X"A8",X"23",X"77",X"3E",X"04",X"CD",X"2F",X"0D",X"18",X"1E",X"35",
		X"20",X"1B",X"23",X"7E",X"B7",X"3A",X"CD",X"80",X"CC",X"2C",X"0D",X"28",X"10",X"34",X"2B",X"3A",
		X"CB",X"80",X"3C",X"3E",X"0D",X"20",X"01",X"87",X"77",X"AF",X"32",X"02",X"A8",X"AF",X"32",X"CC",
		X"80",X"08",X"D9",X"DD",X"E1",X"C9",X"2A",X"1E",X"80",X"ED",X"5B",X"1C",X"80",X"19",X"3E",X"10",
		X"BC",X"30",X"05",X"3E",X"E0",X"BC",X"30",X"12",X"3E",X"03",X"CD",X"2C",X"0D",X"21",X"00",X"00",
		X"ED",X"52",X"EB",X"26",X"11",X"F2",X"AA",X"15",X"26",X"DF",X"22",X"1E",X"80",X"ED",X"53",X"1C",
		X"80",X"2A",X"24",X"80",X"ED",X"5B",X"22",X"80",X"19",X"22",X"24",X"80",X"3E",X"E8",X"BC",X"DA",
		X"85",X"16",X"ED",X"4B",X"35",X"80",X"0A",X"B7",X"28",X"44",X"3A",X"6D",X"80",X"BC",X"CB",X"7A",
		X"28",X"06",X"38",X"3A",X"D6",X"10",X"18",X"02",X"30",X"34",X"C6",X"11",X"CB",X"3F",X"CB",X"3F",
		X"CB",X"3F",X"CE",X"00",X"5F",X"3A",X"1F",X"80",X"C6",X"17",X"CD",X"E2",X"16",X"20",X"2F",X"01",
		X"20",X"00",X"09",X"7E",X"FE",X"10",X"20",X"26",X"3A",X"1F",X"80",X"C6",X"08",X"CD",X"E2",X"16",
		X"20",X"1C",X"B7",X"ED",X"5B",X"22",X"80",X"2A",X"5E",X"80",X"ED",X"5A",X"18",X"1E",X"ED",X"5B",
		X"22",X"80",X"2A",X"5E",X"80",X"ED",X"5A",X"38",X"13",X"22",X"22",X"80",X"18",X"58",X"3E",X"03",
		X"CD",X"2C",X"0D",X"ED",X"5B",X"22",X"80",X"21",X"00",X"00",X"ED",X"52",X"22",X"22",X"80",X"2A",
		X"35",X"80",X"FA",X"55",X"16",X"7E",X"B7",X"23",X"20",X"FB",X"22",X"35",X"80",X"7E",X"B7",X"28",
		X"35",X"32",X"6D",X"80",X"C6",X"11",X"1F",X"1F",X"1F",X"4F",X"06",X"00",X"21",X"35",X"81",X"09",
		X"22",X"6A",X"80",X"18",X"1E",X"2B",X"2B",X"7E",X"B7",X"20",X"FB",X"23",X"22",X"35",X"80",X"7E",
		X"B7",X"28",X"13",X"C6",X"10",X"32",X"6D",X"80",X"3C",X"1F",X"1F",X"1F",X"4F",X"06",X"00",X"21",
		X"35",X"81",X"09",X"22",X"6E",X"80",X"3A",X"1F",X"80",X"32",X"48",X"90",X"3A",X"25",X"80",X"32",
		X"4B",X"90",X"C3",X"A4",X"14",X"01",X"84",X"00",X"3A",X"1F",X"80",X"D6",X"09",X"04",X"0C",X"D6",
		X"28",X"30",X"FA",X"21",X"5F",X"8C",X"11",X"60",X"FF",X"19",X"10",X"FD",X"1E",X"E0",X"06",X"0E",
		X"70",X"19",X"70",X"19",X"7E",X"FE",X"0E",X"28",X"0D",X"FE",X"8B",X"20",X"08",X"3A",X"41",X"88",
		X"3C",X"32",X"41",X"88",X"48",X"71",X"19",X"70",X"19",X"70",X"CD",X"C4",X"16",X"AF",X"32",X"CC",
		X"80",X"C3",X"42",X"05",X"21",X"A4",X"80",X"CB",X"FE",X"21",X"1F",X"88",X"FD",X"21",X"56",X"80",
		X"11",X"20",X"00",X"43",X"7E",X"FD",X"77",X"00",X"19",X"FD",X"2B",X"10",X"F7",X"AF",X"32",X"48",
		X"90",X"C9",X"2A",X"6E",X"80",X"96",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"0E",X"00",X"CB",X"3F",
		X"CB",X"19",X"1F",X"CB",X"19",X"1F",X"CB",X"19",X"47",X"26",X"8C",X"6B",X"ED",X"42",X"7E",X"FE",
		X"10",X"C9",X"4E",X"23",X"7E",X"2B",X"77",X"23",X"1A",X"2F",X"77",X"A1",X"23",X"77",X"23",X"13",
		X"C9",X"11",X"B4",X"17",X"19",X"7E",X"5F",X"21",X"00",X"00",X"E6",X"7F",X"28",X"4D",X"0E",X"00",
		X"FE",X"05",X"28",X"20",X"FE",X"03",X"28",X"18",X"30",X"0C",X"FE",X"01",X"20",X"04",X"CB",X"28",
		X"CB",X"19",X"CB",X"28",X"CB",X"19",X"CB",X"28",X"CB",X"19",X"CB",X"28",X"CB",X"19",X"18",X"29",
		X"CB",X"28",X"CB",X"19",X"CB",X"28",X"CB",X"19",X"CB",X"28",X"CB",X"19",X"60",X"69",X"CB",X"28",
		X"CB",X"19",X"CB",X"28",X"CB",X"19",X"ED",X"4A",X"CB",X"28",X"CB",X"19",X"CB",X"28",X"CB",X"19",
		X"09",X"CB",X"28",X"CB",X"19",X"CB",X"28",X"CB",X"19",X"ED",X"4A",X"7B",X"B7",X"FA",X"76",X"17",
		X"EB",X"21",X"00",X"00",X"ED",X"52",X"3A",X"6D",X"80",X"57",X"1E",X"00",X"19",X"C9",X"7C",X"DD",
		X"21",X"00",X"80",X"DD",X"77",X"00",X"DD",X"77",X"04",X"D6",X"10",X"DD",X"77",X"08",X"DD",X"77",
		X"0C",X"C9",X"8B",X"19",X"CF",X"19",X"25",X"1A",X"7B",X"1A",X"D7",X"1A",X"33",X"1B",X"9B",X"1B",
		X"F1",X"1B",X"47",X"1C",X"A6",X"1C",X"05",X"1D",X"FF",X"85",X"84",X"83",X"82",X"81",X"00",X"01",
		X"02",X"03",X"04",X"05",X"FF",X"85",X"84",X"83",X"82",X"81",X"00",X"01",X"02",X"03",X"04",X"05",
		X"21",X"FF",X"8B",X"06",X"20",X"FD",X"21",X"37",X"80",X"CD",X"3D",X"0B",X"31",X"00",X"88",X"CD",
		X"6C",X"09",X"11",X"35",X"81",X"21",X"01",X"00",X"19",X"EB",X"0E",X"1F",X"70",X"ED",X"B0",X"2A",
		X"5C",X"80",X"11",X"60",X"80",X"1A",X"86",X"32",X"5E",X"80",X"23",X"13",X"1A",X"86",X"32",X"5F",
		X"80",X"23",X"4E",X"23",X"46",X"ED",X"43",X"5C",X"80",X"23",X"13",X"7E",X"12",X"23",X"13",X"7E",
		X"12",X"23",X"23",X"23",X"22",X"35",X"80",X"EB",X"21",X"49",X"90",X"36",X"20",X"21",X"00",X"00",
		X"22",X"1A",X"80",X"22",X"20",X"80",X"22",X"22",X"80",X"21",X"00",X"04",X"22",X"1C",X"80",X"3E",
		X"10",X"32",X"1F",X"80",X"32",X"48",X"90",X"32",X"25",X"80",X"32",X"4B",X"90",X"1A",X"32",X"6D",
		X"80",X"F5",X"C6",X"11",X"1F",X"1F",X"1F",X"4F",X"06",X"00",X"21",X"35",X"81",X"09",X"22",X"6A",
		X"80",X"22",X"6E",X"80",X"F1",X"01",X"E0",X"FF",X"26",X"8B",X"C6",X"11",X"1F",X"1F",X"1F",X"C6",
		X"E0",X"6F",X"13",X"1A",X"B7",X"28",X"11",X"36",X"2B",X"09",X"3D",X"20",X"FA",X"13",X"1A",X"B7",
		X"28",X"06",X"09",X"3D",X"20",X"FC",X"18",X"EA",X"13",X"1A",X"B7",X"20",X"DB",X"3A",X"62",X"80",
		X"32",X"A0",X"88",X"3A",X"63",X"80",X"32",X"80",X"88",X"AF",X"32",X"40",X"88",X"32",X"72",X"80",
		X"32",X"CC",X"80",X"21",X"11",X"80",X"77",X"2B",X"36",X"04",X"11",X"12",X"80",X"01",X"06",X"00",
		X"ED",X"B0",X"EB",X"77",X"21",X"A4",X"80",X"CB",X"BE",X"21",X"18",X"80",X"3A",X"72",X"80",X"B7",
		X"28",X"06",X"CD",X"C4",X"16",X"C3",X"42",X"05",X"3A",X"A4",X"80",X"CD",X"2C",X"09",X"CB",X"66",
		X"C4",X"E8",X"18",X"CB",X"76",X"C4",X"BA",X"18",X"18",X"E2",X"CD",X"5B",X"07",X"2A",X"6A",X"80",
		X"E5",X"11",X"35",X"81",X"B7",X"ED",X"52",X"29",X"26",X"90",X"D1",X"1A",X"CB",X"60",X"28",X"04",
		X"C6",X"04",X"18",X"06",X"CB",X"68",X"28",X"04",X"D6",X"04",X"77",X"12",X"21",X"01",X"00",X"22",
		X"14",X"80",X"21",X"18",X"80",X"CB",X"B6",X"C9",X"3A",X"40",X"88",X"3D",X"F2",X"14",X"19",X"3A",
		X"80",X"88",X"3D",X"F2",X"0F",X"19",X"3A",X"A0",X"88",X"3D",X"28",X"0C",X"FE",X"0F",X"20",X"0A",
		X"32",X"72",X"80",X"21",X"FF",X"7F",X"18",X"12",X"3E",X"10",X"32",X"A0",X"88",X"3E",X"09",X"32",
		X"80",X"88",X"3E",X"09",X"32",X"40",X"88",X"2A",X"2D",X"80",X"22",X"10",X"80",X"21",X"18",X"80",
		X"CB",X"A6",X"C9",X"19",X"00",X"56",X"19",X"03",X"05",X"00",X"00",X"1F",X"04",X"08",X"02",X"07",
		X"05",X"06",X"00",X"3F",X"02",X"06",X"04",X"08",X"04",X"08",X"00",X"67",X"03",X"0A",X"02",X"05",
		X"03",X"09",X"00",X"7F",X"02",X"04",X"02",X"04",X"04",X"08",X"04",X"04",X"00",X"9F",X"04",X"06",
		X"02",X"06",X"06",X"08",X"00",X"00",X"19",X"00",X"23",X"19",X"03",X"00",X"00",X"00",X"1F",X"02",
		X"06",X"03",X"08",X"02",X"0B",X"00",X"37",X"03",X"04",X"05",X"04",X"03",X"05",X"04",X"04",X"00",
		X"6F",X"05",X"08",X"02",X"06",X"03",X"08",X"00",X"8F",X"05",X"08",X"02",X"06",X"03",X"08",X"00",
		X"B7",X"02",X"06",X"03",X"07",X"02",X"04",X"03",X"05",X"00",X"00",X"2B",X"00",X"00",X"00",X"2B",
		X"E0",X"FF",X"00",X"2B",X"40",X"00",X"00",X"2B",X"A0",X"FF",X"00",X"2B",X"80",X"00",X"00",X"2B",
		X"60",X"FF",X"00",X"2B",X"C0",X"00",X"00",X"2B",X"20",X"FF",X"00",X"2B",X"00",X"01",X"00",X"2B",
		X"E0",X"FE",X"00",X"2B",X"40",X"01",X"00",X"2B",X"A0",X"FE",X"00",X"2B",X"80",X"01",X"00",X"2B",
		X"60",X"FE",X"00",X"2B",X"C0",X"01",X"00",X"2B",X"20",X"FE",X"00",X"2B",X"00",X"02",X"00",X"4B",
		X"00",X"00",X"00",X"4C",X"E0",X"FF",X"00",X"60",X"40",X"00",X"5A",X"FF",X"FF",X"00",X"4D",X"A1",
		X"FF",X"00",X"5F",X"80",X"00",X"59",X"FF",X"FF",X"00",X"4E",X"61",X"FF",X"00",X"5E",X"C0",X"00",
		X"58",X"FF",X"FF",X"00",X"4F",X"21",X"FF",X"00",X"5D",X"00",X"01",X"57",X"FF",X"FF",X"00",X"50",
		X"E1",X"FE",X"00",X"5C",X"40",X"01",X"56",X"FF",X"FF",X"00",X"51",X"A1",X"FE",X"00",X"5B",X"80",
		X"01",X"55",X"FF",X"FF",X"00",X"52",X"61",X"FE",X"00",X"54",X"BF",X"01",X"00",X"53",X"21",X"FE",
		X"00",X"53",X"FF",X"01",X"00",X"2C",X"00",X"00",X"00",X"2D",X"E0",X"FF",X"00",X"36",X"40",X"00",
		X"33",X"FF",X"FF",X"00",X"2E",X"A1",X"FF",X"00",X"35",X"80",X"00",X"32",X"FF",X"FF",X"00",X"2F",
		X"61",X"FF",X"00",X"34",X"C0",X"00",X"31",X"FF",X"FF",X"00",X"30",X"21",X"FF",X"00",X"30",X"FF",
		X"00",X"00",X"31",X"E1",X"FE",X"34",X"01",X"00",X"00",X"2F",X"3E",X"01",X"00",X"32",X"A1",X"FE",
		X"35",X"01",X"00",X"00",X"2E",X"7E",X"01",X"00",X"33",X"61",X"FE",X"36",X"01",X"00",X"00",X"2D",
		X"BE",X"01",X"00",X"2C",X"22",X"FE",X"00",X"2C",X"FE",X"01",X"00",X"37",X"00",X"00",X"00",X"38",
		X"E0",X"FF",X"00",X"3F",X"40",X"00",X"3C",X"FF",X"FF",X"00",X"39",X"A1",X"FF",X"00",X"3E",X"80",
		X"00",X"3B",X"FF",X"FF",X"00",X"3A",X"61",X"FF",X"3D",X"01",X"00",X"00",X"3D",X"BF",X"00",X"3A",
		X"FF",X"FF",X"00",X"3B",X"21",X"FF",X"3E",X"01",X"00",X"00",X"39",X"FE",X"00",X"00",X"3C",X"E1",
		X"FE",X"3F",X"01",X"00",X"00",X"38",X"3E",X"01",X"00",X"37",X"A2",X"FE",X"00",X"37",X"7E",X"01",
		X"00",X"38",X"62",X"FE",X"00",X"3F",X"BE",X"01",X"3C",X"FF",X"FF",X"00",X"39",X"23",X"FE",X"00",
		X"3E",X"FE",X"01",X"3B",X"FF",X"FF",X"00",X"40",X"00",X"00",X"00",X"41",X"E0",X"FF",X"00",X"45",
		X"40",X"00",X"43",X"FF",X"FF",X"00",X"42",X"A1",X"FF",X"44",X"01",X"00",X"00",X"44",X"7F",X"00",
		X"42",X"FF",X"FF",X"00",X"43",X"61",X"FF",X"45",X"01",X"00",X"00",X"41",X"BE",X"00",X"00",X"40",
		X"22",X"FF",X"00",X"40",X"FE",X"00",X"00",X"41",X"E2",X"FE",X"00",X"45",X"3E",X"01",X"43",X"FF",
		X"FF",X"00",X"42",X"A3",X"FE",X"44",X"01",X"00",X"00",X"44",X"7D",X"01",X"42",X"FF",X"FF",X"00",
		X"43",X"63",X"FE",X"45",X"01",X"00",X"00",X"41",X"BC",X"01",X"00",X"40",X"24",X"FE",X"00",X"40",
		X"FC",X"01",X"00",X"46",X"00",X"00",X"00",X"47",X"E0",X"FF",X"49",X"01",X"00",X"00",X"4A",X"3F",
		X"00",X"48",X"FF",X"FF",X"00",X"48",X"A1",X"FF",X"4A",X"01",X"00",X"00",X"49",X"7F",X"00",X"47",
		X"FF",X"FF",X"00",X"46",X"62",X"FF",X"00",X"46",X"BE",X"00",X"00",X"47",X"22",X"FF",X"49",X"01",
		X"00",X"00",X"4A",X"FD",X"00",X"48",X"FF",X"FF",X"00",X"48",X"E3",X"FE",X"4A",X"01",X"00",X"00",
		X"49",X"3D",X"01",X"47",X"FF",X"FF",X"00",X"46",X"A4",X"FE",X"00",X"46",X"7C",X"01",X"00",X"47",
		X"64",X"FE",X"49",X"01",X"00",X"00",X"4A",X"BB",X"01",X"48",X"FF",X"FF",X"00",X"48",X"25",X"FE",
		X"4A",X"01",X"00",X"00",X"49",X"FB",X"01",X"47",X"FF",X"FF",X"00",X"4C",X"00",X"00",X"00",X"4B",
		X"E0",X"FF",X"00",X"4D",X"40",X"00",X"00",X"60",X"A0",X"FF",X"5A",X"FF",X"FF",X"00",X"4E",X"81",
		X"00",X"00",X"5F",X"60",X"FF",X"59",X"FF",X"FF",X"00",X"4F",X"C1",X"00",X"00",X"5E",X"20",X"FF",
		X"58",X"FF",X"FF",X"00",X"50",X"01",X"01",X"00",X"5D",X"E0",X"FE",X"57",X"FF",X"FF",X"00",X"51",
		X"41",X"01",X"00",X"5C",X"A0",X"FE",X"56",X"FF",X"FF",X"00",X"52",X"81",X"01",X"00",X"5B",X"60",
		X"FE",X"55",X"FF",X"FF",X"00",X"53",X"C1",X"01",X"00",X"54",X"1F",X"FE",X"00",X"54",X"01",X"02",
		X"00",X"65",X"00",X"00",X"00",X"66",X"E0",X"FF",X"69",X"FF",X"FF",X"00",X"64",X"41",X"00",X"00",
		X"67",X"A0",X"FF",X"6A",X"FF",X"FF",X"00",X"63",X"81",X"00",X"00",X"68",X"60",X"FF",X"6B",X"FF",
		X"FF",X"00",X"62",X"C1",X"00",X"00",X"61",X"1F",X"FF",X"00",X"61",X"01",X"01",X"00",X"62",X"DF",
		X"FE",X"00",X"6B",X"41",X"01",X"68",X"01",X"00",X"00",X"63",X"9E",X"FE",X"00",X"6A",X"81",X"01",
		X"67",X"01",X"00",X"00",X"64",X"5E",X"FE",X"00",X"69",X"C1",X"01",X"66",X"01",X"00",X"00",X"65",
		X"1E",X"FE",X"00",X"65",X"02",X"02",X"00",X"6F",X"00",X"00",X"72",X"FF",X"FF",X"00",X"70",X"E1",
		X"FF",X"73",X"FF",X"FF",X"00",X"6E",X"41",X"00",X"00",X"71",X"A0",X"FF",X"74",X"FF",X"FF",X"00",
		X"6D",X"81",X"00",X"00",X"6C",X"5F",X"FF",X"00",X"6C",X"C1",X"00",X"00",X"6D",X"1F",X"FF",X"00",
		X"74",X"01",X"01",X"71",X"01",X"00",X"00",X"6E",X"DE",X"FE",X"00",X"73",X"41",X"01",X"70",X"01",
		X"00",X"00",X"6F",X"9E",X"FE",X"72",X"FF",X"FF",X"00",X"72",X"82",X"01",X"6F",X"01",X"00",X"00",
		X"70",X"5E",X"FE",X"73",X"FF",X"FF",X"00",X"6E",X"C3",X"01",X"00",X"71",X"1E",X"FE",X"74",X"FF",
		X"FF",X"00",X"6D",X"03",X"02",X"00",X"77",X"00",X"00",X"79",X"FF",X"FF",X"00",X"78",X"E1",X"FF",
		X"7A",X"FF",X"FF",X"00",X"76",X"41",X"00",X"00",X"75",X"9F",X"FF",X"00",X"75",X"81",X"00",X"00",
		X"76",X"5F",X"FF",X"00",X"7A",X"C1",X"00",X"78",X"01",X"00",X"00",X"77",X"1E",X"FF",X"79",X"FF",
		X"FF",X"00",X"79",X"02",X"01",X"77",X"01",X"00",X"00",X"78",X"DE",X"FE",X"7A",X"FF",X"FF",X"00",
		X"76",X"43",X"01",X"00",X"75",X"9D",X"FE",X"00",X"75",X"83",X"01",X"00",X"76",X"5D",X"FE",X"00",
		X"7A",X"C3",X"01",X"78",X"01",X"00",X"00",X"77",X"1C",X"FE",X"79",X"FF",X"FF",X"00",X"79",X"04",
		X"02",X"77",X"01",X"00",X"00",X"7C",X"00",X"00",X"7E",X"FF",X"FF",X"00",X"7D",X"E1",X"FF",X"7F",
		X"FF",X"FF",X"00",X"7B",X"41",X"00",X"00",X"7B",X"9F",X"FF",X"00",X"7F",X"81",X"00",X"7D",X"01",
		X"00",X"00",X"7C",X"5E",X"FF",X"00",X"7E",X"C1",X"00",X"7C",X"01",X"00",X"00",X"7D",X"1E",X"FF",
		X"7F",X"FF",X"FF",X"00",X"7B",X"03",X"01",X"00",X"7B",X"DD",X"FE",X"00",X"7F",X"43",X"01",X"7D",
		X"01",X"00",X"00",X"7C",X"9C",X"FE",X"7E",X"FF",X"FF",X"00",X"7E",X"84",X"01",X"7C",X"01",X"00",
		X"00",X"7D",X"5C",X"FE",X"7F",X"FF",X"FF",X"00",X"7B",X"C5",X"01",X"00",X"7B",X"1B",X"FE",X"00",
		X"7F",X"05",X"02",X"7D",X"01",X"00",X"00",X"FE",X"00",X"10",X"55",X"41",X"00",X"20",X"8A",X"00",
		X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"8A",X"00",X"55",X"55",X"00",X"15",X"41",X"00",X"00",X"00",
		X"14",X"55",X"55",X"45",X"00",X"00",X"28",X"AA",X"AA",X"80",X"10",X"55",X"40",X"00",X"00",X"00",
		X"14",X"55",X"55",X"55",X"41",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"14",X"55",X"55",X"00",X"10",X"00",X"15",X"55",X"55",
		X"55",X"55",X"55",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",X"88",X"00",X"00",X"00",
		X"10",X"55",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"55",X"45",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"28",X"8A",
		X"00",X"00",X"2A",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",X"10",X"55",X"40",X"00",X"00",X"2A",
		X"AA",X"AA",X"82",X"00",X"55",X"55",X"41",X"00",X"00",X"15",X"00",X"00",X"28",X"AA",X"AA",X"80",
		X"0A",X"00",X"00",X"00",X"80",X"14",X"55",X"55",X"55",X"55",X"55",X"45",X"21",X"70",X"80",X"34",
		X"11",X"19",X"80",X"21",X"B2",X"1E",X"01",X"0D",X"00",X"ED",X"B0",X"11",X"04",X"00",X"21",X"00",
		X"80",X"7E",X"D6",X"10",X"FE",X"E0",X"38",X"0C",X"FE",X"F0",X"3E",X"DF",X"38",X"01",X"AF",X"43",
		X"77",X"19",X"10",X"FC",X"21",X"03",X"80",X"43",X"3E",X"DF",X"BE",X"30",X"01",X"77",X"19",X"10",
		X"F7",X"21",X"04",X"00",X"22",X"16",X"80",X"01",X"00",X"04",X"DD",X"21",X"1A",X"80",X"FD",X"21",
		X"00",X"80",X"11",X"04",X"00",X"FD",X"7E",X"00",X"FE",X"E0",X"38",X"0B",X"DD",X"7E",X"00",X"ED",
		X"44",X"DD",X"77",X"00",X"FD",X"7E",X"00",X"DD",X"86",X"00",X"FD",X"77",X"00",X"DD",X"7E",X"01",
		X"C6",X"96",X"DD",X"77",X"01",X"30",X"03",X"DD",X"34",X"02",X"FD",X"7E",X"03",X"FE",X"F0",X"30",
		X"07",X"DD",X"86",X"02",X"FD",X"77",X"03",X"0C",X"3A",X"19",X"80",X"FD",X"AE",X"01",X"FD",X"77",
		X"01",X"FD",X"19",X"1D",X"DD",X"19",X"10",X"BA",X"3A",X"19",X"80",X"EE",X"C0",X"32",X"19",X"80",
		X"21",X"18",X"80",X"CB",X"06",X"36",X"00",X"30",X"F7",X"79",X"B7",X"20",X"94",X"21",X"70",X"80",
		X"35",X"C9",X"40",X"04",X"00",X"FC",X"02",X"00",X"FB",X"FD",X"00",X"F9",X"FB",X"00",X"FD",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
