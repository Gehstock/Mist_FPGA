library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_PGM_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_PGM_1 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"FD",X"6E",X"06",X"FD",X"66",X"07",X"29",X"F5",X"11",X"00",X"00",X"ED",X"5A",X"F1",X"FD",X"75",
		X"06",X"FD",X"74",X"07",X"38",X"36",X"FD",X"7E",X"04",X"FE",X"07",X"D8",X"21",X"32",X"25",X"FD",
		X"7E",X"11",X"B7",X"28",X"03",X"FD",X"35",X"11",X"FD",X"46",X"0A",X"FD",X"7E",X"09",X"FE",X"02",
		X"20",X"04",X"78",X"EE",X"02",X"47",X"78",X"CD",X"E1",X"3D",X"D5",X"C1",X"FD",X"66",X"01",X"FD",
		X"6E",X"03",X"CD",X"83",X"3D",X"FD",X"74",X"01",X"FD",X"75",X"03",X"C9",X"FD",X"7E",X"04",X"FE",
		X"07",X"38",X"C9",X"FD",X"7E",X"11",X"E6",X"0F",X"FE",X"01",X"28",X"C0",X"21",X"3A",X"25",X"FD",
		X"35",X"11",X"18",X"BB",X"FD",X"7E",X"0A",X"16",X"00",X"5F",X"19",X"7E",X"FD",X"77",X"00",X"C9",
		X"3A",X"E7",X"49",X"FE",X"09",X"38",X"02",X"3E",X"09",X"16",X"00",X"5F",X"19",X"7E",X"FD",X"77",
		X"04",X"FD",X"77",X"05",X"21",X"69",X"26",X"CD",X"E1",X"3D",X"FD",X"73",X"06",X"FD",X"72",X"07",
		X"C9",X"FD",X"7E",X"04",X"21",X"A3",X"80",X"16",X"00",X"5F",X"19",X"7E",X"FD",X"B6",X"0C",X"FD",
		X"77",X"0C",X"C9",X"10",X"08",X"08",X"07",X"07",X"06",X"06",X"05",X"05",X"05",X"FD",X"7E",X"09",
		X"FE",X"01",X"C8",X"FD",X"7E",X"0C",X"CB",X"BF",X"B7",X"28",X"04",X"FD",X"35",X"0C",X"C9",X"E5",
		X"CD",X"91",X"80",X"E1",X"FD",X"7E",X"0A",X"CD",X"E1",X"3D",X"FD",X"7E",X"00",X"FD",X"CB",X"0C",
		X"7E",X"20",X"0A",X"BA",X"28",X"07",X"FD",X"CB",X"0C",X"BE",X"3C",X"18",X"08",X"BB",X"28",X"F3",
		X"FD",X"CB",X"0C",X"FE",X"3D",X"FD",X"77",X"00",X"C9",X"ED",X"5F",X"5F",X"ED",X"5F",X"6F",X"26",
		X"00",X"54",X"ED",X"5F",X"E6",X"03",X"3C",X"47",X"86",X"19",X"10",X"FC",X"C9",X"FD",X"66",X"01",
		X"FD",X"6E",X"03",X"CD",X"9E",X"0F",X"E6",X"0F",X"21",X"4E",X"81",X"16",X"00",X"5F",X"19",X"4E",
		X"C5",X"21",X"61",X"26",X"06",X"04",X"C5",X"4E",X"23",X"46",X"23",X"E5",X"FD",X"66",X"01",X"FD",
		X"6E",X"03",X"CD",X"83",X"3D",X"CD",X"9E",X"0F",X"FE",X"FF",X"28",X"1F",X"B7",X"28",X"1C",X"E6",
		X"F0",X"28",X"04",X"FE",X"80",X"20",X"14",X"37",X"E1",X"C1",X"CB",X"19",X"10",X"D8",X"CB",X"39",
		X"CB",X"39",X"CB",X"39",X"CB",X"39",X"79",X"C1",X"A1",X"4F",X"C9",X"A7",X"18",X"EA",X"00",X"03",
		X"09",X"06",X"0C",X"05",X"0A",X"07",X"0D",X"0E",X"0B",X"0F",X"0E",X"0F",X"7E",X"23",X"5E",X"23",
		X"56",X"23",X"D5",X"DD",X"E1",X"E5",X"F5",X"DD",X"7E",X"09",X"FE",X"04",X"30",X"0C",X"CD",X"80",
		X"81",X"CD",X"EA",X"81",X"CD",X"60",X"82",X"CD",X"C5",X"82",X"F1",X"E1",X"3D",X"20",X"DF",X"C9",
		X"06",X"0E",X"DD",X"7E",X"0A",X"DF",X"8E",X"81",X"A6",X"81",X"CC",X"81",X"E4",X"81",X"FD",X"7E",
		X"01",X"DD",X"BE",X"01",X"C0",X"FD",X"7E",X"03",X"5F",X"D6",X"11",X"57",X"DD",X"7E",X"03",X"BB",
		X"D0",X"BA",X"D2",X"1E",X"83",X"C9",X"1E",X"0D",X"16",X"10",X"FD",X"7E",X"03",X"6F",X"D6",X"10",
		X"67",X"DD",X"7E",X"03",X"BD",X"D0",X"BC",X"D8",X"DD",X"7E",X"01",X"FD",X"96",X"01",X"38",X"05",
		X"BB",X"D0",X"C3",X"1E",X"83",X"ED",X"44",X"BA",X"D0",X"C3",X"1E",X"83",X"FD",X"7E",X"01",X"DD",
		X"BE",X"01",X"C0",X"FD",X"7E",X"03",X"5F",X"D6",X"10",X"57",X"DD",X"7E",X"03",X"BB",X"D0",X"BA",
		X"D8",X"C3",X"1E",X"83",X"1E",X"10",X"16",X"0D",X"18",X"C0",X"06",X"0D",X"DD",X"7E",X"0A",X"DF",
		X"14",X"82",X"F8",X"81",X"3E",X"82",X"44",X"82",X"FD",X"7E",X"03",X"DD",X"BE",X"03",X"C0",X"FD",
		X"7E",X"01",X"5F",X"C6",X"10",X"30",X"02",X"3E",X"FF",X"57",X"DD",X"7E",X"01",X"BB",X"D8",X"BA",
		X"DA",X"1E",X"83",X"C9",X"1E",X"10",X"16",X"0D",X"FD",X"7E",X"01",X"6F",X"C6",X"10",X"30",X"02",
		X"3E",X"FF",X"67",X"DD",X"7E",X"01",X"BD",X"D8",X"BC",X"D0",X"DD",X"7E",X"03",X"FD",X"96",X"03",
		X"38",X"05",X"BB",X"D0",X"C3",X"1E",X"83",X"ED",X"44",X"BA",X"D0",X"C3",X"1E",X"83",X"1E",X"0D",
		X"16",X"10",X"18",X"D4",X"FD",X"7E",X"03",X"DD",X"BE",X"03",X"C0",X"FD",X"7E",X"01",X"5F",X"C6",
		X"10",X"30",X"02",X"3E",X"FF",X"57",X"DD",X"7E",X"01",X"BB",X"D8",X"BA",X"D0",X"C3",X"1E",X"83",
		X"06",X"0B",X"DD",X"7E",X"0A",X"DF",X"8A",X"82",X"A6",X"82",X"6E",X"82",X"BF",X"82",X"FD",X"7E",
		X"01",X"DD",X"BE",X"01",X"C0",X"FD",X"7E",X"03",X"5F",X"C6",X"11",X"30",X"02",X"3E",X"FF",X"57",
		X"DD",X"7E",X"03",X"BB",X"D8",X"BA",X"DA",X"1E",X"83",X"C9",X"FD",X"7E",X"01",X"DD",X"BE",X"01",
		X"C0",X"FD",X"7E",X"03",X"5F",X"C6",X"10",X"30",X"02",X"3E",X"FF",X"57",X"DD",X"7E",X"03",X"BB",
		X"D8",X"BA",X"D0",X"C3",X"1E",X"83",X"1E",X"0D",X"16",X"10",X"FD",X"7E",X"03",X"6F",X"C6",X"10",
		X"30",X"02",X"3E",X"FF",X"67",X"DD",X"7E",X"03",X"BD",X"D8",X"BC",X"D0",X"C3",X"B8",X"81",X"1E",
		X"10",X"16",X"0D",X"18",X"E5",X"06",X"07",X"DD",X"7E",X"0A",X"DF",X"EB",X"82",X"00",X"83",X"18",
		X"83",X"D3",X"82",X"FD",X"7E",X"03",X"DD",X"BE",X"03",X"C0",X"FD",X"7E",X"01",X"5F",X"D6",X"10",
		X"57",X"DD",X"7E",X"01",X"BB",X"D0",X"BA",X"D2",X"1E",X"83",X"C9",X"1E",X"10",X"16",X"0D",X"FD",
		X"7E",X"01",X"6F",X"D6",X"10",X"67",X"DD",X"7E",X"01",X"BD",X"D0",X"BC",X"D8",X"C3",X"2A",X"82",
		X"FD",X"7E",X"03",X"DD",X"BE",X"03",X"C0",X"FD",X"7E",X"01",X"5F",X"D6",X"1F",X"57",X"DD",X"7E",
		X"01",X"BB",X"D0",X"BA",X"D8",X"C3",X"1E",X"83",X"16",X"0D",X"1E",X"10",X"18",X"D1",X"78",X"A1",
		X"4F",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"21",X"14",X"4A",X"06",X"38",X"CF",X"21",X"7A",
		X"84",X"11",X"14",X"4A",X"01",X"10",X"00",X"ED",X"B0",X"21",X"8A",X"84",X"11",X"34",X"4A",X"01",
		X"04",X"00",X"ED",X"B0",X"21",X"8E",X"84",X"11",X"58",X"4A",X"01",X"0B",X"00",X"ED",X"B0",X"06",
		X"0B",X"21",X"99",X"40",X"11",X"6F",X"84",X"C5",X"D5",X"1A",X"5F",X"01",X"02",X"02",X"3E",X"BC",
		X"CD",X"1E",X"3D",X"D1",X"13",X"C1",X"10",X"EF",X"3E",X"D0",X"1E",X"05",X"01",X"02",X"02",X"21",
		X"15",X"43",X"CD",X"1E",X"3D",X"3E",X"BC",X"1E",X"02",X"01",X"02",X"02",X"21",X"95",X"41",X"CD",
		X"1E",X"3D",X"3E",X"BC",X"1E",X"04",X"01",X"02",X"02",X"21",X"15",X"42",X"CD",X"1E",X"3D",X"3E",
		X"02",X"01",X"50",X"8C",X"FF",X"3E",X"23",X"06",X"01",X"FF",X"FD",X"21",X"14",X"4A",X"FD",X"7E",
		X"0E",X"FE",X"03",X"20",X"14",X"FD",X"E5",X"FD",X"7E",X"21",X"FE",X"C8",X"DC",X"26",X"84",X"FD",
		X"E1",X"FD",X"7E",X"21",X"FE",X"10",X"CA",X"99",X"84",X"CD",X"BB",X"1B",X"FD",X"7E",X"09",X"21",
		X"C5",X"83",X"F7",X"18",X"0A",X"1C",X"84",X"1C",X"84",X"02",X"16",X"1D",X"84",X"57",X"16",X"FD",
		X"7E",X"08",X"21",X"D8",X"83",X"F7",X"18",X"04",X"E1",X"83",X"0A",X"84",X"CD",X"90",X"11",X"18",
		X"B4",X"CD",X"B2",X"1A",X"1E",X"02",X"FD",X"7E",X"21",X"FE",X"E0",X"20",X"10",X"FD",X"7E",X"23",
		X"FE",X"58",X"20",X"02",X"1E",X"03",X"FD",X"73",X"0F",X"CD",X"D6",X"13",X"C9",X"1E",X"01",X"FD",
		X"7E",X"23",X"FE",X"58",X"20",X"F0",X"1E",X"03",X"18",X"EC",X"FD",X"7E",X"10",X"B7",X"28",X"06",
		X"FD",X"35",X"10",X"C3",X"E4",X"83",X"CD",X"7A",X"14",X"C3",X"E4",X"83",X"C9",X"FD",X"7E",X"21",
		X"FE",X"A0",X"D0",X"C3",X"29",X"16",X"FD",X"21",X"58",X"4A",X"FD",X"7E",X"09",X"FE",X"FF",X"C8",
		X"FD",X"7E",X"09",X"B7",X"20",X"0E",X"21",X"A1",X"28",X"CD",X"AD",X"80",X"CD",X"00",X"80",X"CD",
		X"7D",X"1E",X"18",X"1B",X"FE",X"04",X"20",X"14",X"CD",X"AA",X"20",X"FD",X"7E",X"09",X"FE",X"06",
		X"20",X"0D",X"FD",X"36",X"09",X"FF",X"FD",X"36",X"00",X"00",X"18",X"03",X"CD",X"0D",X"21",X"21",
		X"58",X"4A",X"11",X"A2",X"4B",X"01",X"04",X"00",X"ED",X"B0",X"AF",X"32",X"A1",X"4B",X"C9",X"01",
		X"02",X"03",X"04",X"01",X"02",X"03",X"04",X"01",X"02",X"03",X"85",X"10",X"9F",X"38",X"86",X"00",
		X"9F",X"38",X"00",X"00",X"06",X"06",X"FF",X"FF",X"01",X"04",X"9E",X"08",X"9E",X"38",X"AD",X"10",
		X"5B",X"58",X"06",X"06",X"FF",X"FF",X"00",X"00",X"01",X"3E",X"12",X"FF",X"CD",X"57",X"0E",X"3E",
		X"01",X"01",X"78",X"86",X"FF",X"21",X"2C",X"85",X"11",X"88",X"4B",X"01",X"0F",X"00",X"ED",X"B0",
		X"3E",X"23",X"06",X"04",X"FF",X"DD",X"21",X"4A",X"85",X"CD",X"B2",X"3C",X"3E",X"50",X"32",X"63",
		X"48",X"3E",X"23",X"06",X"04",X"FF",X"DD",X"21",X"5C",X"85",X"CD",X"B2",X"3C",X"3E",X"60",X"32",
		X"62",X"48",X"3E",X"23",X"06",X"04",X"FF",X"DD",X"21",X"69",X"85",X"CD",X"B2",X"3C",X"21",X"3B",
		X"85",X"11",X"A1",X"4B",X"01",X"05",X"00",X"ED",X"B0",X"3E",X"23",X"06",X"04",X"FF",X"DD",X"21",
		X"7D",X"85",X"CD",X"B2",X"3C",X"21",X"40",X"85",X"11",X"A6",X"4B",X"01",X"05",X"00",X"ED",X"B0",
		X"3E",X"23",X"06",X"04",X"FF",X"DD",X"21",X"8E",X"85",X"CD",X"B2",X"3C",X"21",X"45",X"85",X"11",
		X"AB",X"4B",X"01",X"05",X"00",X"ED",X"B0",X"3E",X"23",X"06",X"04",X"FF",X"DD",X"21",X"A1",X"85",
		X"CD",X"B2",X"3C",X"3E",X"23",X"06",X"C0",X"FF",X"3E",X"11",X"FF",X"C9",X"00",X"85",X"58",X"9F",
		X"88",X"00",X"86",X"48",X"9F",X"88",X"00",X"9E",X"50",X"9E",X"88",X"00",X"AD",X"50",X"5B",X"B8",
		X"00",X"AD",X"50",X"5D",X"C8",X"00",X"AD",X"50",X"5C",X"D8",X"04",X"0B",X"AF",X"41",X"00",X"06",
		X"56",X"41",X"4E",X"3A",X"56",X"41",X"4E",X"20",X"43",X"41",X"52",X"00",X"04",X"06",X"AD",X"41",
		X"00",X"06",X"45",X"4E",X"45",X"52",X"47",X"59",X"00",X"04",X"0D",X"AB",X"41",X"00",X"06",X"42",
		X"4F",X"4E",X"55",X"53",X"20",X"42",X"41",X"4C",X"4C",X"4F",X"4F",X"4E",X"00",X"04",X"0A",X"A9",
		X"41",X"00",X"06",X"52",X"45",X"44",X"20",X"4B",X"49",X"4C",X"4C",X"45",X"52",X"00",X"04",X"0C",
		X"A7",X"41",X"00",X"06",X"47",X"52",X"45",X"45",X"4E",X"20",X"4B",X"49",X"4C",X"4C",X"45",X"52",
		X"00",X"04",X"0B",X"A5",X"41",X"00",X"06",X"42",X"4C",X"55",X"45",X"20",X"4B",X"49",X"4C",X"4C",
		X"45",X"52",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"31",X"E0",X"4E",X"DD",X"21",X"0F",X"86",X"21",
		X"7F",X"40",X"3A",X"01",X"48",X"CB",X"6F",X"28",X"07",X"21",X"BF",X"42",X"DD",X"21",X"18",X"86",
		X"DD",X"E5",X"E5",X"CD",X"B2",X"3C",X"3E",X"23",X"06",X"18",X"FF",X"E1",X"E5",X"01",X"02",X"01",
		X"3E",X"00",X"CD",X"99",X"3C",X"E1",X"DD",X"E1",X"3E",X"23",X"06",X"10",X"FF",X"18",X"E1",X"00",
		X"02",X"7F",X"40",X"00",X"0D",X"31",X"50",X"00",X"00",X"02",X"BF",X"42",X"00",X"0D",X"32",X"50",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"31",X"F0",X"4D",X"3E",X"23",X"06",X"20",X"FF",
		X"3A",X"02",X"48",X"CB",X"47",X"CB",X"C7",X"32",X"02",X"48",X"21",X"30",X"48",X"7E",X"4F",X"E6",
		X"F0",X"28",X"17",X"FE",X"70",X"30",X"13",X"79",X"E6",X"0F",X"77",X"E5",X"C5",X"CD",X"F4",X"0F",
		X"C1",X"CD",X"02",X"8D",X"E1",X"3E",X"23",X"06",X"0A",X"FF",X"23",X"11",X"02",X"49",X"B7",X"E5",
		X"ED",X"52",X"E1",X"38",X"D8",X"3E",X"23",X"06",X"40",X"FF",X"3E",X"47",X"06",X"10",X"FF",X"3E",
		X"60",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"31",X"30",X"4E",X"21",X"59",X"87",X"3A",X"02",
		X"48",X"CB",X"77",X"28",X"03",X"21",X"8A",X"87",X"11",X"E8",X"4A",X"01",X"31",X"00",X"ED",X"B0",
		X"3E",X"23",X"06",X"01",X"FF",X"06",X"07",X"FD",X"21",X"E8",X"4A",X"C5",X"FD",X"7E",X"02",X"B7",
		X"CC",X"B5",X"86",X"3E",X"23",X"06",X"01",X"FF",X"FD",X"35",X"02",X"01",X"07",X"00",X"FD",X"09",
		X"C1",X"10",X"E8",X"18",X"E0",X"FD",X"7E",X"01",X"CB",X"BF",X"FD",X"77",X"02",X"FD",X"7E",X"00",
		X"FD",X"CB",X"01",X"7E",X"20",X"0B",X"FE",X"02",X"28",X"0B",X"FD",X"CB",X"01",X"BE",X"3C",X"18",
		X"09",X"FE",X"00",X"28",X"F5",X"FD",X"CB",X"01",X"FE",X"3D",X"FD",X"77",X"00",X"FD",X"6E",X"03",
		X"FD",X"66",X"04",X"FD",X"5E",X"05",X"FD",X"56",X"06",X"0E",X"02",X"D5",X"E5",X"06",X"0F",X"C5",
		X"1A",X"47",X"B7",X"28",X"45",X"E6",X"F0",X"28",X"41",X"FE",X"70",X"30",X"3D",X"D5",X"E5",X"FE",
		X"60",X"20",X"14",X"1E",X"06",X"0E",X"21",X"FD",X"7E",X"00",X"87",X"87",X"81",X"E1",X"E5",X"01",
		X"02",X"02",X"CD",X"1E",X"3D",X"18",X"21",X"FE",X"50",X"20",X"06",X"1E",X"05",X"0E",X"D0",X"18",
		X"E6",X"CD",X"4B",X"0F",X"D5",X"FD",X"7E",X"00",X"21",X"53",X"87",X"CD",X"E1",X"3D",X"D5",X"DD",
		X"E1",X"D1",X"E1",X"E5",X"78",X"CD",X"50",X"89",X"E1",X"D1",X"C1",X"13",X"23",X"23",X"10",X"AF",
		X"E1",X"11",X"C0",X"01",X"19",X"D1",X"C5",X"EB",X"01",X"69",X"00",X"09",X"EB",X"C1",X"0D",X"C2",
		X"EB",X"86",X"C9",X"FB",X"89",X"27",X"8A",X"53",X"8A",X"01",X"01",X"05",X"41",X"40",X"30",X"48",
		X"01",X"82",X"03",X"81",X"40",X"3F",X"48",X"01",X"01",X"01",X"C1",X"40",X"4E",X"48",X"01",X"82",
		X"04",X"01",X"41",X"5D",X"48",X"01",X"01",X"02",X"41",X"41",X"6C",X"48",X"01",X"82",X"03",X"81",
		X"41",X"7B",X"48",X"01",X"01",X"04",X"C1",X"41",X"8A",X"48",X"01",X"02",X"02",X"41",X"40",X"30",
		X"48",X"01",X"02",X"02",X"81",X"40",X"3F",X"48",X"01",X"02",X"02",X"C1",X"40",X"4E",X"48",X"01",
		X"02",X"02",X"01",X"41",X"5D",X"48",X"01",X"02",X"02",X"41",X"41",X"6C",X"48",X"01",X"02",X"02",
		X"81",X"41",X"7B",X"48",X"01",X"02",X"02",X"C1",X"41",X"8A",X"48",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"21",X"20",X"4B",X"06",X"28",X"CF",X"3E",X"08",X"32",X"20",X"4B",X"DD",X"21",X"21",X"4B",X"FD",
		X"7E",X"0A",X"CD",X"EB",X"3D",X"CB",X"FF",X"DD",X"77",X"00",X"FD",X"7E",X"01",X"DD",X"77",X"01",
		X"FD",X"7E",X"03",X"DD",X"77",X"03",X"CD",X"78",X"88",X"DD",X"77",X"04",X"CD",X"9B",X"88",X"28",
		X"51",X"DD",X"77",X"02",X"47",X"3A",X"20",X"4B",X"3D",X"CA",X"6B",X"88",X"32",X"20",X"4B",X"FE",
		X"07",X"30",X"11",X"FD",X"7E",X"0F",X"DD",X"BE",X"01",X"20",X"09",X"FD",X"7E",X"10",X"DD",X"BE",
		X"03",X"CA",X"6B",X"88",X"78",X"2F",X"E6",X"0F",X"DD",X"A6",X"04",X"DD",X"77",X"04",X"78",X"DD",
		X"66",X"01",X"DD",X"6E",X"03",X"CD",X"F7",X"3D",X"CD",X"37",X"89",X"DD",X"74",X"06",X"DD",X"75",
		X"08",X"DD",X"7E",X"02",X"DD",X"77",X"05",X"DD",X"36",X"07",X"00",X"01",X"05",X"00",X"DD",X"09",
		X"18",X"A4",X"DD",X"CB",X"00",X"7E",X"20",X"2D",X"DD",X"7E",X"00",X"E6",X"0F",X"2F",X"E6",X"0F",
		X"DD",X"A6",X"FF",X"DD",X"77",X"FF",X"DD",X"E5",X"E1",X"06",X"05",X"CF",X"01",X"FB",X"FF",X"DD",
		X"09",X"3A",X"20",X"4B",X"3C",X"32",X"20",X"4B",X"C3",X"EC",X"87",X"3A",X"23",X"4B",X"FD",X"36",
		X"11",X"10",X"C3",X"5E",X"23",X"C3",X"14",X"23",X"DD",X"66",X"01",X"DD",X"6E",X"03",X"CD",X"9E",
		X"0F",X"FE",X"FF",X"28",X"14",X"E6",X"F0",X"28",X"04",X"FE",X"80",X"20",X"0C",X"7E",X"E6",X"0F",
		X"21",X"4E",X"81",X"16",X"00",X"5F",X"19",X"7E",X"C9",X"AF",X"C9",X"3E",X"05",X"DD",X"A6",X"00",
		X"20",X"3E",X"FD",X"7E",X"03",X"FD",X"BE",X"10",X"20",X"28",X"3E",X"02",X"FD",X"BE",X"08",X"20",
		X"18",X"DD",X"CB",X"00",X"4E",X"28",X"0A",X"DD",X"7E",X"01",X"FD",X"BE",X"0F",X"38",X"0A",X"18",
		X"11",X"DD",X"7E",X"01",X"FD",X"BE",X"0F",X"38",X"09",X"DD",X"7E",X"00",X"E6",X"0F",X"DD",X"A6",
		X"04",X"C0",X"06",X"01",X"FD",X"7E",X"03",X"FD",X"BE",X"10",X"30",X"40",X"06",X"04",X"18",X"3C",
		X"FD",X"7E",X"01",X"FD",X"BE",X"0F",X"20",X"28",X"3E",X"02",X"FD",X"BE",X"08",X"20",X"18",X"DD",
		X"CB",X"00",X"46",X"20",X"0A",X"DD",X"7E",X"03",X"FD",X"BE",X"10",X"38",X"0A",X"18",X"11",X"DD",
		X"7E",X"03",X"FD",X"BE",X"10",X"38",X"09",X"DD",X"7E",X"00",X"E6",X"0F",X"DD",X"A6",X"04",X"C0",
		X"06",X"02",X"FD",X"7E",X"01",X"FD",X"BE",X"0F",X"38",X"02",X"06",X"08",X"78",X"DD",X"A6",X"04",
		X"C0",X"DD",X"7E",X"00",X"E6",X"0F",X"DD",X"A6",X"04",X"C0",X"78",X"CD",X"F7",X"3D",X"EE",X"02",
		X"CD",X"EB",X"3D",X"DD",X"A6",X"04",X"C9",X"E5",X"21",X"61",X"26",X"CD",X"E1",X"3D",X"E1",X"D5",
		X"C1",X"CD",X"83",X"3D",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E6",X"0F",X"3D",X"87",X"87",X"06",X"00",X"4F",X"DD",X"09",X"01",X"02",X"02",X"C5",X"E5",X"DD",
		X"7E",X"00",X"77",X"CB",X"D4",X"73",X"CB",X"94",X"23",X"DD",X"23",X"10",X"F2",X"E1",X"01",X"20",
		X"00",X"09",X"C1",X"0D",X"20",X"E7",X"C9",X"61",X"60",X"62",X"63",X"64",X"67",X"65",X"66",X"68",
		X"69",X"6A",X"6B",X"6C",X"6D",X"6E",X"6F",X"70",X"70",X"71",X"71",X"73",X"72",X"73",X"72",X"70",
		X"70",X"6A",X"63",X"6C",X"67",X"71",X"71",X"6C",X"72",X"6A",X"72",X"73",X"67",X"73",X"63",X"6C",
		X"67",X"6A",X"63",X"82",X"79",X"7E",X"77",X"7C",X"75",X"80",X"7B",X"78",X"83",X"76",X"7F",X"74",
		X"7D",X"7A",X"81",X"78",X"79",X"7A",X"7B",X"7C",X"7D",X"7E",X"7F",X"78",X"79",X"76",X"77",X"74",
		X"75",X"7A",X"7B",X"74",X"7D",X"76",X"7F",X"7C",X"75",X"7E",X"77",X"74",X"75",X"76",X"77",X"92",
		X"89",X"8E",X"87",X"8C",X"85",X"90",X"8B",X"88",X"93",X"86",X"8F",X"84",X"8D",X"8A",X"91",X"88",
		X"89",X"8A",X"8B",X"8C",X"8D",X"8E",X"8F",X"88",X"89",X"86",X"87",X"84",X"85",X"8A",X"8B",X"84",
		X"8D",X"86",X"8F",X"8C",X"85",X"8E",X"87",X"84",X"85",X"86",X"87",X"9A",X"95",X"9C",X"97",X"9A",
		X"95",X"9F",X"99",X"94",X"9B",X"96",X"9D",X"94",X"9B",X"98",X"9E",X"94",X"95",X"98",X"99",X"9A",
		X"9B",X"9C",X"9D",X"94",X"95",X"96",X"97",X"94",X"95",X"98",X"99",X"94",X"9B",X"96",X"9D",X"9A",
		X"95",X"9C",X"97",X"94",X"95",X"96",X"97",X"AE",X"A5",X"AA",X"A3",X"A8",X"A1",X"AF",X"A7",X"A4",
		X"AC",X"A2",X"AB",X"A0",X"A9",X"A6",X"AD",X"A4",X"A5",X"A6",X"A7",X"A8",X"A9",X"AA",X"AB",X"A4",
		X"A5",X"A2",X"A3",X"A0",X"A1",X"A6",X"A7",X"A0",X"A9",X"A2",X"AB",X"A8",X"A1",X"AA",X"A3",X"A0",
		X"A1",X"A2",X"A3",X"BB",X"B5",X"B8",X"B3",X"B6",X"B1",X"B8",X"B3",X"B4",X"BA",X"B2",X"B9",X"B0",
		X"B7",X"B2",X"B9",X"B4",X"B5",X"B2",X"B3",X"B6",X"B7",X"B8",X"B9",X"B4",X"B5",X"B2",X"B3",X"B0",
		X"B1",X"B2",X"B3",X"B6",X"B7",X"B2",X"B9",X"B6",X"B1",X"B8",X"B3",X"B0",X"B1",X"B2",X"B3",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"11",X"0F",X"48",X"3A",X"01",X"48",X"CB",X"6F",X"28",X"03",X"11",X"15",X"48",X"06",X"1E",X"21",
		X"60",X"4C",X"0E",X"01",X"C5",X"E5",X"D5",X"06",X"06",X"CD",X"71",X"3D",X"D1",X"E1",X"C1",X"FE",
		X"02",X"28",X"0A",X"C5",X"01",X"08",X"00",X"09",X"C1",X"0C",X"10",X"E8",X"C9",X"79",X"F5",X"FE",
		X"1E",X"28",X"19",X"3E",X"1E",X"91",X"21",X"08",X"00",X"3D",X"28",X"06",X"01",X"08",X"00",X"09",
		X"18",X"F7",X"E5",X"C1",X"21",X"47",X"4D",X"11",X"4F",X"4D",X"ED",X"B8",X"F1",X"F5",X"3D",X"21",
		X"60",X"4C",X"4F",X"87",X"87",X"87",X"06",X"00",X"4F",X"09",X"11",X"0F",X"48",X"3A",X"01",X"48",
		X"CB",X"6F",X"28",X"03",X"11",X"15",X"48",X"EB",X"01",X"06",X"00",X"ED",X"B0",X"EB",X"3A",X"E8",
		X"49",X"77",X"23",X"3A",X"E9",X"49",X"77",X"DD",X"21",X"0D",X"8C",X"CD",X"B2",X"3C",X"DD",X"21",
		X"2C",X"8C",X"CD",X"B2",X"3C",X"3E",X"23",X"06",X"30",X"FF",X"F1",X"F5",X"21",X"00",X"01",X"22",
		X"14",X"4A",X"21",X"60",X"4C",X"FE",X"0B",X"38",X"14",X"11",X"50",X"00",X"19",X"D6",X"0A",X"E5",
		X"2A",X"14",X"4A",X"11",X"01",X"00",X"19",X"22",X"14",X"4A",X"E1",X"18",X"E8",X"CD",X"A9",X"8B",
		X"F1",X"FE",X"0B",X"38",X"04",X"D6",X"0A",X"18",X"F8",X"21",X"D6",X"44",X"3D",X"28",X"04",X"2B",
		X"2B",X"18",X"F9",X"06",X"3C",X"1E",X"0B",X"C5",X"E5",X"06",X"13",X"73",X"CD",X"4D",X"3D",X"10",
		X"FA",X"3E",X"23",X"06",X"03",X"FF",X"1C",X"7B",X"FE",X"10",X"38",X"02",X"1E",X"0B",X"E1",X"C1",
		X"10",X"E5",X"C9",X"DD",X"21",X"0D",X"8C",X"CD",X"B2",X"3C",X"DD",X"21",X"2C",X"8C",X"CD",X"B2",
		X"3C",X"21",X"00",X"01",X"22",X"14",X"4A",X"21",X"60",X"4C",X"CD",X"A9",X"8B",X"3E",X"23",X"06",
		X"80",X"FF",X"21",X"B0",X"4C",X"CD",X"A9",X"8B",X"3E",X"23",X"06",X"80",X"FF",X"21",X"00",X"4D",
		X"CD",X"A9",X"8B",X"3E",X"23",X"06",X"80",X"FF",X"C9",X"E5",X"DD",X"E1",X"21",X"F6",X"40",X"06",
		X"0A",X"C5",X"DD",X"E5",X"E5",X"DD",X"21",X"14",X"4A",X"1E",X"0C",X"06",X"02",X"0E",X"00",X"CD",
		X"8A",X"3D",X"E1",X"DD",X"E1",X"DD",X"E5",X"E5",X"01",X"C0",X"00",X"09",X"1E",X"0D",X"06",X"06",
		X"0E",X"00",X"CD",X"8A",X"3D",X"E1",X"DD",X"E1",X"DD",X"E5",X"E5",X"01",X"00",X"02",X"09",X"01",
		X"06",X"00",X"DD",X"09",X"1E",X"0A",X"06",X"02",X"0E",X"00",X"CD",X"8A",X"3D",X"3E",X"23",X"06",
		X"02",X"FF",X"11",X"15",X"4A",X"21",X"0C",X"8C",X"06",X"02",X"CD",X"54",X"3D",X"E1",X"DD",X"E1",
		X"2B",X"2B",X"01",X"08",X"00",X"DD",X"09",X"C1",X"10",X"A7",X"C9",X"00",X"01",X"00",X"18",X"9C",
		X"40",X"00",X"0B",X"54",X"4F",X"44",X"41",X"59",X"3B",X"53",X"20",X"48",X"49",X"5F",X"53",X"43",
		X"4F",X"52",X"45",X"20",X"42",X"45",X"53",X"54",X"20",X"33",X"30",X"00",X"00",X"05",X"D8",X"40",
		X"00",X"0C",X"4F",X"52",X"44",X"45",X"52",X"05",X"D8",X"41",X"00",X"0D",X"53",X"43",X"4F",X"52",
		X"45",X"05",X"D8",X"42",X"00",X"0A",X"4C",X"45",X"56",X"45",X"4C",X"00",X"FF",X"FF",X"FF",X"FF",
		X"31",X"20",X"4F",X"21",X"50",X"4D",X"06",X"1E",X"CF",X"1E",X"3C",X"3E",X"23",X"06",X"01",X"FF",
		X"3A",X"01",X"48",X"CB",X"57",X"20",X"0C",X"1D",X"20",X"09",X"1E",X"3C",X"3A",X"DC",X"49",X"3C",
		X"32",X"DC",X"49",X"D5",X"FD",X"21",X"50",X"4D",X"06",X"05",X"C5",X"FD",X"7E",X"00",X"FD",X"B6",
		X"01",X"C4",X"90",X"8C",X"01",X"06",X"00",X"FD",X"09",X"C1",X"10",X"EE",X"D1",X"C3",X"5B",X"8C",
		X"FD",X"7E",X"03",X"B7",X"28",X"04",X"FD",X"35",X"03",X"C9",X"FD",X"36",X"03",X"04",X"FD",X"6E",
		X"00",X"FD",X"66",X"01",X"01",X"02",X"02",X"FD",X"7E",X"02",X"FE",X"00",X"20",X"2E",X"3A",X"02",
		X"48",X"CB",X"77",X"C2",X"EF",X"8C",X"3A",X"02",X"48",X"CB",X"47",X"28",X"0C",X"3E",X"14",X"CB",
		X"D4",X"5E",X"CB",X"94",X"CD",X"1E",X"3D",X"18",X"0C",X"FD",X"7E",X"04",X"1E",X"03",X"DD",X"21",
		X"77",X"89",X"CD",X"50",X"89",X"FD",X"E5",X"E1",X"06",X"06",X"CF",X"C9",X"CB",X"D4",X"5E",X"CB",
		X"94",X"FD",X"7E",X"02",X"F5",X"CD",X"1E",X"3D",X"F1",X"D6",X"04",X"FD",X"77",X"02",X"C9",X"E5",
		X"FD",X"7E",X"04",X"E6",X"0F",X"21",X"60",X"8D",X"CD",X"E1",X"3D",X"E1",X"7A",X"CD",X"1E",X"3D",
		X"18",X"D3",X"FD",X"21",X"50",X"4D",X"06",X"05",X"FD",X"7E",X"00",X"FD",X"B6",X"01",X"28",X"08",
		X"11",X"06",X"00",X"FD",X"19",X"10",X"F1",X"C9",X"FD",X"75",X"00",X"FD",X"74",X"01",X"FD",X"71",
		X"04",X"FD",X"36",X"02",X"0C",X"79",X"0E",X"04",X"FE",X"50",X"38",X"02",X"0E",X"10",X"21",X"59",
		X"8D",X"3A",X"02",X"48",X"CB",X"47",X"28",X"11",X"21",X"5F",X"8D",X"79",X"E5",X"16",X"00",X"1E",
		X"00",X"CD",X"20",X"2C",X"E1",X"CD",X"04",X"3E",X"C9",X"E5",X"C5",X"3E",X"04",X"CD",X"8E",X"2C",
		X"C1",X"E1",X"18",X"E7",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",
		X"11",X"E0",X"12",X"E4",X"13",X"E8",X"11",X"DC",X"13",X"E0",X"12",X"E4",X"15",X"E8",X"00",X"00",
		X"11",X"EC",X"16",X"E4",X"12",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
