library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity rom_char_u is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of rom_char_u is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7C",X"18",X"30",X"78",X"F8",X"7C",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"7F",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",
		X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"E0",X"E0",X"E0",X"F0",X"F0",X"F0",
		X"F8",X"FC",X"36",X"36",X"36",X"36",X"FC",X"F8",X"F0",X"E0",X"C0",X"80",X"80",X"00",X"00",X"00",
		X"00",X"C0",X"F0",X"F8",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"87",X"FF",X"86",X"FF",
		X"FF",X"FF",X"86",X"86",X"86",X"86",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"7E",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"DB",X"C3",X"FF",X"F7",X"FF",X"E7",X"FF",X"FF",X"FF",X"81",X"81",X"81",X"81",X"FF",X"FF",
		X"FF",X"FF",X"C3",X"FF",X"C3",X"C3",X"FF",X"FF",X"C3",X"FF",X"FF",X"C3",X"C3",X"FF",X"FF",X"C3",
		X"00",X"03",X"0F",X"1F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E1",X"FF",X"61",X"FF",
		X"FF",X"FF",X"61",X"61",X"61",X"61",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"03",X"03",X"07",X"07",X"07",X"0F",X"0F",X"0F",X"1F",X"3F",X"6C",X"6C",X"6C",X"6C",X"3F",X"1F",
		X"0F",X"07",X"03",X"01",X"01",X"00",X"00",X"00",X"42",X"7E",X"C3",X"7E",X"7E",X"C3",X"7E",X"42",
		X"C0",X"60",X"F0",X"58",X"7C",X"C6",X"7F",X"42",X"03",X"06",X"0F",X"1A",X"3E",X"63",X"FE",X"62",
		X"00",X"00",X"00",X"00",X"C0",X"70",X"FC",X"47",X"C0",X"70",X"FC",X"47",X"7F",X"C0",X"7F",X"42",
		X"03",X"0E",X"3F",X"E2",X"FE",X"03",X"FE",X"42",X"00",X"00",X"00",X"00",X"03",X"0E",X"3F",X"E2",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"80",X"C0",X"E0",X"70",X"B8",X"DC",
		X"EE",X"E7",X"E7",X"CF",X"9C",X"3B",X"77",X"EF",X"00",X"FF",X"FF",X"EF",X"CC",X"BB",X"77",X"EF",
		X"CF",X"CF",X"E7",X"73",X"B9",X"DC",X"EE",X"F7",X"00",X"FF",X"FF",X"F7",X"3B",X"DD",X"EE",X"F7",
		X"F3",X"F3",X"E7",X"CE",X"9D",X"3B",X"77",X"EF",X"00",X"00",X"01",X"03",X"07",X"0E",X"1D",X"3B",
		X"77",X"E7",X"E7",X"F3",X"39",X"DC",X"EE",X"F7",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"A0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"F0",X"E0",X"C0",X"80",X"00",X"00",
		X"78",X"78",X"70",X"F0",X"E0",X"E0",X"C0",X"C0",X"C0",X"E0",X"F8",X"3C",X"1C",X"0C",X"0C",X"0C",
		X"00",X"00",X"00",X"00",X"40",X"E0",X"E8",X"FC",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"7B",X"7F",X"FF",X"FF",X"FC",X"10",X"10",X"10",X"38",X"38",X"38",X"7D",X"7D",
		X"80",X"C1",X"F7",X"77",X"3E",X"1C",X"1C",X"1C",X"00",X"00",X"00",X"00",X"02",X"07",X"17",X"3F",
		X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DE",X"FE",X"FF",X"FF",X"3F",
		X"08",X"08",X"08",X"1C",X"1C",X"1C",X"3E",X"3E",X"01",X"83",X"EF",X"EE",X"7C",X"38",X"38",X"38",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"05",X"0F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"0F",X"0F",X"07",X"03",X"01",X"00",X"00",X"1E",X"1E",X"0E",X"0F",X"07",X"07",X"03",X"03",
		X"03",X"07",X"1F",X"3C",X"38",X"30",X"30",X"30",X"23",X"11",X"11",X"08",X"48",X"48",X"44",X"60",
		X"44",X"49",X"23",X"27",X"8F",X"9F",X"3F",X"7F",X"22",X"82",X"C2",X"E1",X"F1",X"F8",X"FC",X"FE",
		X"20",X"29",X"49",X"43",X"43",X"27",X"27",X"0F",X"4F",X"5F",X"1F",X"3F",X"3F",X"7F",X"7F",X"7F",
		X"4F",X"4F",X"6F",X"2F",X"2F",X"AF",X"8F",X"0F",X"F1",X"F9",X"F9",X"FC",X"FC",X"FE",X"FE",X"FE",
		X"24",X"90",X"92",X"C2",X"CA",X"EA",X"E1",X"F1",X"F2",X"F2",X"F4",X"F4",X"FF",X"F2",X"F2",X"F1",
		X"B2",X"92",X"88",X"88",X"C4",X"C4",X"D0",X"E3",X"BD",X"81",X"3C",X"81",X"81",X"3C",X"81",X"BD",
		X"3F",X"1F",X"0F",X"A7",X"83",X"39",X"80",X"BD",X"FC",X"F9",X"F0",X"E5",X"C1",X"9C",X"01",X"BD",
		X"FF",X"FF",X"FF",X"FF",X"3F",X"8F",X"03",X"38",X"3F",X"0F",X"03",X"B8",X"80",X"3F",X"80",X"BD",
		X"FC",X"F1",X"C0",X"1D",X"01",X"FC",X"01",X"BD",X"FF",X"FF",X"FF",X"FF",X"FC",X"F1",X"C0",X"1D",
		X"81",X"E7",X"7F",X"3A",X"38",X"FA",X"FF",X"FF",X"80",X"B0",X"E0",X"6C",X"38",X"3A",X"FE",X"FF",
		X"01",X"0D",X"07",X"36",X"1C",X"5C",X"7D",X"FF",X"00",X"00",X"00",X"00",X"B0",X"E0",X"FA",X"FF",
		X"80",X"F0",X"E2",X"FC",X"FD",X"FF",X"FF",X"FF",X"01",X"0F",X"26",X"3C",X"B8",X"F3",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"0D",X"07",X"5F",X"FF",X"80",X"80",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",
		X"00",X"00",X"FC",X"FC",X"C0",X"00",X"00",X"00",X"00",X"C0",X"F0",X"F8",X"FC",X"FE",X"FE",X"FF",
		X"FF",X"F6",X"FA",X"FB",X"FD",X"FE",X"FF",X"FF",X"00",X"00",X"03",X"0F",X"7F",X"FC",X"F0",X"E0",
		X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",
		X"7E",X"FF",X"99",X"99",X"99",X"81",X"81",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"81",X"C3",X"E7",X"E7",X"E7",X"FF",X"7E",X"3C",X"18",X"18",X"18",
		X"00",X"7E",X"FF",X"FF",X"FF",X"FF",X"3C",X"00",X"00",X"03",X"0F",X"1F",X"3F",X"7F",X"7F",X"FF",
		X"FF",X"AF",X"EF",X"DF",X"DF",X"BF",X"FF",X"FF",X"00",X"00",X"C0",X"F0",X"FE",X"3F",X"0F",X"07",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",
		X"01",X"01",X"03",X"03",X"07",X"07",X"0F",X"0F",X"00",X"00",X"3F",X"3F",X"03",X"00",X"00",X"00",
		X"01",X"0B",X"0E",X"04",X"04",X"0E",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"1B",X"0E",X"4C",X"7C",X"3E",X"67",X"C3",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"1E",X"1E",X"3E",X"3C",X"7C",X"78",X"F8",X"F0",X"F0",X"E0",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"60",X"60",X"70",X"30",X"B8",X"B8",X"9C",X"DE",X"CF",X"E7",X"F3",X"00",
		X"FF",X"FF",X"FF",X"FC",X"FC",X"F8",X"F8",X"F8",X"F0",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EE",X"EE",X"EE",X"DC",X"DC",X"D8",X"D8",X"D8",X"D8",X"D8",X"FF",X"FF",X"FF",X"FF",X"D8",X"D8",
		X"00",X"00",X"00",X"00",X"66",X"66",X"E7",X"E7",X"E7",X"C3",X"C3",X"C3",X"C3",X"81",X"81",X"00",
		X"FF",X"FF",X"FF",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7E",X"7E",X"7E",X"BD",X"BD",X"BD",X"BD",X"BD",X"BD",X"BD",X"FF",X"FF",X"FF",X"FF",X"BD",X"BD",
		X"00",X"00",X"00",X"00",X"06",X"06",X"0E",X"0C",X"1D",X"1D",X"39",X"7B",X"F3",X"E7",X"CF",X"00",
		X"FF",X"FF",X"FF",X"3F",X"3F",X"1F",X"1F",X"1F",X"0F",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"77",X"77",X"77",X"3B",X"3B",X"1B",X"1B",X"1B",X"1B",X"1B",X"FF",X"FF",X"FF",X"FF",X"1B",X"1B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"78",X"78",X"7C",X"3C",X"3E",
		X"1E",X"1F",X"0F",X"0F",X"07",X"01",X"01",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"80",X"C0",X"E0",X"F0",X"F8",X"FC",X"FE",X"FF",X"01",X"03",X"07",X"0F",X"1F",X"3F",X"7F",X"FF",
		X"FF",X"FE",X"FC",X"F8",X"F0",X"E0",X"C0",X"80",X"FF",X"7F",X"3F",X"1F",X"0F",X"07",X"03",X"01",
		X"7F",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"7F",X"3F",X"0F",X"07",X"03",X"01",X"00",X"FF",X"FF",X"FF",X"7F",X"3F",X"0F",X"07",X"01",
		X"FF",X"FF",X"F0",X"80",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",
		X"F0",X"F0",X"E0",X"C0",X"80",X"80",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"FC",X"FC",X"F8",X"F0",X"E0",X"E0",X"C0",X"80",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FC",X"F0",X"F0",X"E0",X"E0",X"C0",X"C0",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FC",X"F8",X"F0",X"E0",X"C0",
		X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FC",X"F8",X"E0",X"C0",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"03",X"1F",X"7F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"07",X"1F",X"3F",X"3F",X"7F",X"7F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",
		X"1F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"01",X"01",X"03",X"07",X"0F",
		X"1F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"01",X"03",X"07",X"0F",X"1F",
		X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"03",X"07",X"07",X"0F",X"1F",X"1F",
		X"3F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"C0",X"C0",X"E0",X"E0",X"E0",X"F0",X"F0",X"F8",X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"E0",X"F0",X"F0",X"F8",X"FE",X"FF",X"FF",
		X"00",X"00",X"00",X"E0",X"F8",X"FC",X"FE",X"FF",X"00",X"3C",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"03",X"03",X"07",X"1F",X"1F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"E7",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"C0",X"E0",X"E0",X"E0",X"F0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"F0",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"0F",X"1F",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"07",X"0F",X"0F",X"1F",X"7F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"07",X"1F",X"3F",X"7F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"81",X"C7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"C0",X"C0",X"E0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"03",X"0F",X"3F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",
		X"03",X"03",X"07",X"07",X"0F",X"0F",X"1F",X"1F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"03",X"07",X"0F",X"0F",X"1F",X"1F",X"3F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"80",X"C0",X"E0",X"F0",X"F9",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"80",X"C0",X"C0",X"C0",X"E0",X"F0",X"F0",X"F8",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"80",X"C0",X"C0",X"E0",X"E0",X"E0",X"F0",X"F0",X"F8",X"FC",X"FE",X"FF",X"FF",
		X"C0",X"C0",X"C0",X"E0",X"F0",X"F0",X"F8",X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"01",X"07",X"1F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"01",X"01",X"01",X"03",X"07",X"0F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"07",X"0F",X"0F",X"1F",X"3F",X"7F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"01",X"03",X"03",X"07",X"07",X"0F",X"1F",X"1F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"01",X"03",X"07",X"8F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"80",X"C0",X"F0",X"F8",X"F8",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"F8",X"FC",X"FE",X"FF",X"FF",
		X"00",X"00",X"00",X"03",X"07",X"07",X"0F",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"80",X"C0",X"C0",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F0",X"FC",X"FE",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"E0",X"F0",X"F0",
		X"F8",X"F8",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"FC",X"FE",X"FE",X"FE",X"FE",X"FF",X"FF",X"01",X"03",X"03",X"03",X"07",X"07",X"07",X"07",
		X"07",X"0F",X"0F",X"0F",X"1F",X"FF",X"FF",X"FF",X"00",X"00",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",
		X"00",X"00",X"03",X"07",X"1F",X"3F",X"3F",X"3F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"03",X"0F",X"1F",X"1F",X"3F",X"FF",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"E1",
		X"F3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"C0",X"E0",X"F8",X"FC",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"F0",X"F8",X"F8",X"FC",X"FF",
		X"00",X"00",X"00",X"7F",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",
		X"07",X"0F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",
		X"07",X"0F",X"1F",X"3F",X"7F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"07",X"0F",X"1F",X"3F",X"7F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"83",
		X"87",X"CF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"80",X"80",X"80",X"C0",X"E0",X"F8",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"E0",X"F0",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"F0",X"F8",X"F8",X"FC",X"FE",X"FE",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"80",X"C0",X"F0",X"F8",X"F8",X"FC",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"FF",
		X"00",X"00",X"00",X"E0",X"F8",X"FF",X"FF",X"FF",X"C0",X"C0",X"C0",X"E1",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"1F",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"3F",X"1F",X"0F",X"03",X"00",X"00",X"FF",X"7F",X"7F",X"3F",X"3F",X"1F",X"0F",X"07",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"1F",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",
		X"1F",X"1F",X"07",X"03",X"03",X"01",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"7F",X"3F",X"1F",X"1F",X"0F",X"0F",X"07",X"03",X"01",X"01",X"01",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",X"3F",X"1F",X"0F",X"07",X"07",X"03",X"01",X"01",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"3F",X"1F",X"1F",X"0F",X"0F",X"07",X"07",X"03",X"03",X"01",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",
		X"3F",X"1F",X"1F",X"0F",X"0F",X"07",X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"7F",X"3F",X"1F",X"1F",X"1F",X"07",X"03",X"01",X"01",X"01",X"00",X"00",X"00",X"00",
		X"FF",X"3F",X"1F",X"1E",X"1E",X"00",X"00",X"00",X"FF",X"FE",X"FC",X"FC",X"F8",X"F8",X"F8",X"F8",
		X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",
		X"FE",X"FC",X"F8",X"F8",X"F0",X"E0",X"E0",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"FC",X"F8",X"F8",X"F0",X"E0",X"E0",X"C0",X"C0",X"80",X"80",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FE",X"FC",X"FC",X"F8",X"F8",X"F0",
		X"E0",X"E0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",
		X"FC",X"FC",X"F8",X"F8",X"F0",X"E0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"7E",X"3C",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",
		X"3F",X"1F",X"1F",X"0F",X"07",X"07",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"1F",X"0F",X"0F",X"07",X"03",X"01",X"01",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"1F",X"0F",X"0F",X"07",X"03",X"01",X"01",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FD",X"F8",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FE",X"FC",X"FC",X"F8",X"F8",X"F0",X"F0",X"E0",X"C0",X"C0",X"80",X"80",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",X"F0",
		X"E0",X"E0",X"E0",X"C0",X"C0",X"80",X"80",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FE",X"FC",X"F8",X"F8",X"F0",X"F0",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",
		X"7F",X"7F",X"7F",X"3F",X"1F",X"1F",X"0F",X"03",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"3F",X"1F",X"0F",X"07",X"07",X"07",X"0F",X"0F",X"0F",X"07",X"03",X"03",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",X"1F",X"0F",X"0F",X"1F",X"1F",X"1F",X"1F",X"07",
		X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"1F",X"0F",
		X"0F",X"07",X"07",X"03",X"03",X"03",X"03",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",X"1F",X"0F",X"0F",X"0F",X"07",X"07",X"07",X"07",
		X"07",X"03",X"03",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"F9",X"F1",X"E0",X"C0",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FC",X"F0",X"C0",X"80",X"80",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",X"F0",X"F0",X"E0",X"C0",X"C0",X"C0",X"80",X"80",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",X"F8",X"F0",
		X"E0",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"FE",X"FE",X"FC",X"F8",X"F8",X"F0",X"F0",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"80",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",X"F0",
		X"F0",X"F0",X"F0",X"E0",X"E0",X"C0",X"80",X"80",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FE",X"FC",X"FC",X"F8",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FE",X"FC",X"F8",X"F8",X"F0",X"E0",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FE",X"FC",X"F8",X"E0",X"80",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"07",X"0F",X"0F",X"1F",X"1F",X"1F",X"3F",X"3F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"03",X"03",X"07",X"07",X"07",X"07",X"07",X"07",
		X"0F",X"0F",X"0F",X"0F",X"1F",X"1F",X"3F",X"3F",X"3F",X"3F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"01",X"01",X"01",X"03",X"03",X"03",X"07",
		X"07",X"07",X"07",X"0F",X"0F",X"0F",X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",X"3F",X"3F",X"3F",X"7F",
		X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"01",X"81",X"81",
		X"C3",X"C3",X"C3",X"E3",X"E7",X"E7",X"FF",X"FF",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"E0",X"E0",
		X"E0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",X"FE",
		X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"80",X"80",X"C0",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FE",
		X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E0",X"E0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"FC",X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"7F",X"7F",X"3F",X"1F",X"0F",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"7F",X"7F",X"3F",X"3F",X"1F",X"1F",X"0F",X"0F",X"07",X"07",X"07",X"03",X"01",X"01",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",
		X"3F",X"3F",X"1F",X"1F",X"0F",X"0F",X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"01",X"01",X"01",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",
		X"3F",X"3F",X"3F",X"1F",X"1F",X"1F",X"0F",X"0F",X"0F",X"07",X"07",X"03",X"03",X"03",X"03",X"03",
		X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"CF",X"03",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FE",X"FC",X"F8",X"F8",X"F0",X"F0",X"E0",X"E0",X"C0",X"C0",X"C0",X"80",X"80",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FC",X"FC",X"FC",X"F8",
		X"F8",X"F8",X"F0",X"F0",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",X"F0",
		X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",X"F8",X"F0",X"E0",X"C0",X"C0",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
