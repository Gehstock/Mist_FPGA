library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity fg_sp_graphx_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of fg_sp_graphx_1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"90",X"10",X"FC",X"16",X"1E",X"16",X"FF",X"97",X"1E",X"16",X"1E",X"14",X"10",X"10",X"00",
		X"03",X"06",X"06",X"1F",X"9F",X"FE",X"FE",X"1F",X"1F",X"0F",X"7F",X"7F",X"5F",X"06",X"16",X"0C",
		X"00",X"10",X"10",X"14",X"1E",X"16",X"FE",X"97",X"1F",X"16",X"1E",X"16",X"1C",X"10",X"90",X"00",
		X"0C",X"16",X"06",X"1F",X"5E",X"7E",X"7F",X"1F",X"1F",X"0F",X"FF",X"FF",X"9F",X"06",X"06",X"03",
		X"00",X"10",X"10",X"F4",X"1E",X"16",X"1E",X"F7",X"1F",X"16",X"1E",X"F6",X"1C",X"10",X"90",X"00",
		X"0C",X"16",X"06",X"5B",X"7A",X"7E",X"1F",X"1F",X"1E",X"FE",X"FB",X"9B",X"1F",X"06",X"06",X"03",
		X"00",X"90",X"10",X"F4",X"1E",X"16",X"1E",X"F7",X"1F",X"16",X"1E",X"F6",X"1C",X"10",X"10",X"00",
		X"03",X"06",X"06",X"9B",X"FA",X"FE",X"1F",X"1F",X"1E",X"7E",X"7B",X"5B",X"1F",X"06",X"16",X"0C",
		X"00",X"E0",X"10",X"1E",X"16",X"FF",X"97",X"1E",X"16",X"1E",X"14",X"10",X"10",X"00",X"00",X"00",
		X"00",X"1F",X"9F",X"FE",X"FE",X"1F",X"1F",X"0F",X"7F",X"7F",X"5F",X"06",X"16",X"0C",X"00",X"00",
		X"00",X"00",X"F8",X"CA",X"8F",X"8B",X"8F",X"8B",X"8E",X"08",X"48",X"80",X"00",X"00",X"00",X"00",
		X"00",X"3F",X"3F",X"0F",X"0F",X"07",X"7F",X"7F",X"4F",X"03",X"03",X"01",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"E0",X"C6",X"C5",X"C7",X"C5",X"84",X"84",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"07",X"03",X"1F",X"1F",X"17",X"01",X"05",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"E0",X"E2",X"E3",X"C2",X"D2",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"1F",X"1F",X"13",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"D2",X"C2",X"7E",X"42",X"C0",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"13",X"1F",X"1F",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"84",X"84",X"FD",X"87",X"85",X"C6",X"F8",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"05",X"01",X"16",X"1E",X"1F",X"07",X"07",X"07",X"00",
		X"00",X"00",X"00",X"00",X"80",X"48",X"08",X"FA",X"0F",X"0B",X"8F",X"FB",X"0E",X"08",X"80",X"00",
		X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"4D",X"7D",X"7F",X"0F",X"0F",X"0F",X"3F",X"3D",X"00",
		X"00",X"00",X"00",X"10",X"10",X"F4",X"1E",X"16",X"1E",X"F7",X"1F",X"16",X"1E",X"F0",X"00",X"00",
		X"00",X"00",X"0C",X"16",X"06",X"5B",X"7A",X"7E",X"1F",X"1F",X"1E",X"FE",X"FB",X"9B",X"1F",X"00",
		X"C0",X"60",X"E1",X"FB",X"DE",X"DC",X"78",X"78",X"F8",X"F8",X"7C",X"5E",X"DB",X"E1",X"60",X"C0",
		X"00",X"01",X"00",X"07",X"0F",X"08",X"08",X"08",X"0F",X"08",X"08",X"08",X"0F",X"00",X"01",X"00",
		X"00",X"80",X"C0",X"B0",X"B1",X"FF",X"FF",X"F0",X"F0",X"FF",X"BF",X"B1",X"F0",X"C0",X"80",X"00",
		X"00",X"07",X"01",X"1F",X"10",X"10",X"11",X"1F",X"10",X"10",X"11",X"1F",X"0F",X"01",X"07",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"2C",X"8C",X"56",X"92",X"E4",X"4E",X"9A",X"9C",X"58",X"28",X"00",
		X"F0",X"DC",X"92",X"FC",X"14",X"19",X"10",X"F1",X"10",X"10",X"11",X"F2",X"18",X"91",X"DC",X"F0",
		X"00",X"01",X"07",X"1B",X"9A",X"FE",X"FF",X"1F",X"1E",X"FE",X"FB",X"9B",X"1F",X"07",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"00",X"C0",X"20",X"30",X"20",X"10",X"20",X"20",X"20",X"40",X"80",X"00",X"00",
		X"80",X"40",X"A9",X"98",X"1C",X"2A",X"34",X"12",X"3D",X"0C",X"16",X"8D",X"14",X"8C",X"42",X"80",
		X"01",X"03",X"07",X"1B",X"9A",X"FE",X"FF",X"1F",X"1E",X"FE",X"FB",X"9B",X"1F",X"07",X"03",X"01",
		X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"00",X"80",X"40",X"00",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"09",X"34",X"31",X"6A",X"49",X"27",X"72",X"59",X"39",X"1A",X"14",X"00",X"00",
		X"00",X"00",X"30",X"00",X"98",X"44",X"86",X"44",X"A2",X"84",X"C4",X"A4",X"88",X"90",X"40",X"00",
		X"00",X"00",X"01",X"03",X"03",X"05",X"06",X"02",X"07",X"01",X"02",X"01",X"02",X"01",X"00",X"00",
		X"00",X"00",X"81",X"00",X"80",X"20",X"00",X"80",X"20",X"00",X"00",X"00",X"81",X"80",X"00",X"00",
		X"00",X"00",X"00",X"1B",X"36",X"14",X"48",X"B0",X"C4",X"28",X"24",X"32",X"0B",X"04",X"00",X"00",
		X"58",X"0E",X"21",X"09",X"1A",X"20",X"00",X"00",X"00",X"00",X"28",X"04",X"06",X"21",X"02",X"18",
		X"04",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"90",X"04",X"88",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"A4",X"40",X"82",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"01",X"10",X"04",X"42",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"02",X"42",X"A6",X"8B",X"D3",X"EE",X"58",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"06",X"02",X"00",X"01",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"90",X"48",X"68",X"60",X"A0",X"28",
		X"F0",X"0C",X"F2",X"FD",X"C3",X"BF",X"41",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"0C",X"13",X"17",X"0F",X"2F",X"5F",X"5E",X"5E",X"5D",X"1D",X"1D",X"1D",X"1D",X"5D",X"5D",
		X"F0",X"0C",X"F2",X"FD",X"C3",X"BF",X"41",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"0C",X"13",X"17",X"2F",X"2F",X"1F",X"1E",X"1E",X"1D",X"5D",X"5D",X"5D",X"5D",X"1D",X"1D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"5D",X"5D",X"1D",X"1D",X"1D",X"1D",X"5D",X"5D",X"5D",X"5D",X"1D",X"1D",X"1D",X"1D",X"5D",X"5D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1D",X"1D",X"5D",X"5D",X"5D",X"5D",X"1D",X"1D",X"1D",X"1D",X"5D",X"5D",X"5D",X"5D",X"1D",X"1D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"E0",X"FC",X"FE",X"FC",X"F8",X"E0",X"F8",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",
		X"C0",X"30",X"08",X"04",X"02",X"02",X"01",X"01",X"01",X"01",X"02",X"02",X"04",X"08",X"30",X"C0",
		X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"F8",X"E0",X"E0",X"F8",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",
		X"00",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"00",
		X"00",X"00",X"03",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"03",X"00",X"00",
		X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",X"1F",X"07",X"07",X"1F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"03",X"4C",X"50",X"D0",X"78",X"58",X"78",X"DC",X"7C",X"58",X"78",X"D8",X"70",X"50",X"4C",X"03",
		X"0C",X"DA",X"D8",X"EF",X"E8",X"F8",X"FC",X"FF",X"F8",X"F8",X"EC",X"EF",X"FC",X"D8",X"DA",X"0C",
		X"00",X"00",X"03",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"03",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"05",X"01",X"81",X"01",X"02",X"04",X"08",X"90",X"30",X"48",X"88",X"04",X"04",X"14",X"04",
		X"02",X"09",X"01",X"00",X"00",X"00",X"00",X"01",X"03",X"01",X"00",X"00",X"01",X"02",X"44",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"9C",X"38",X"80",X"C0",X"60",X"60",X"60",X"60",X"C0",X"80",X"38",X"9C",X"80",X"00",
		X"3F",X"C0",X"01",X"01",X"01",X"02",X"0C",X"1C",X"1C",X"0C",X"02",X"01",X"01",X"01",X"C0",X"3F",
		X"F0",X"0C",X"30",X"40",X"B8",X"70",X"80",X"80",X"80",X"80",X"70",X"B8",X"40",X"30",X"0C",X"F0",
		X"0F",X"60",X"10",X"00",X"0F",X"3E",X"37",X"7F",X"7F",X"37",X"3E",X"0F",X"00",X"10",X"60",X"0F",
		X"C0",X"20",X"67",X"4E",X"60",X"B0",X"18",X"18",X"18",X"18",X"B0",X"60",X"4E",X"67",X"20",X"C0",
		X"0F",X"30",X"00",X"00",X"00",X"00",X"03",X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"30",X"0F",
		X"FC",X"03",X"0C",X"10",X"EE",X"9C",X"E0",X"E0",X"E0",X"E0",X"9C",X"EE",X"10",X"0C",X"03",X"FC",
		X"03",X"18",X"04",X"00",X"03",X"0F",X"0D",X"1F",X"1F",X"0D",X"0F",X"03",X"00",X"04",X"18",X"03",
		X"F0",X"F8",X"B8",X"3C",X"7E",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"7E",X"0C",X"5C",X"3C",X"18",
		X"01",X"B2",X"F8",X"F8",X"FC",X"DF",X"0F",X"07",X"07",X"07",X"07",X"07",X"1F",X"3E",X"1C",X"0E",
		X"18",X"3C",X"5C",X"0E",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"7C",X"38",X"B8",X"F8",X"F0",
		X"0E",X"1C",X"3E",X"1F",X"07",X"07",X"07",X"07",X"07",X"0F",X"DF",X"FC",X"F8",X"F8",X"B2",X"01",
		X"18",X"3C",X"5C",X"0E",X"7E",X"E6",X"AE",X"BE",X"AE",X"E6",X"FE",X"7C",X"3C",X"B8",X"F8",X"F0",
		X"0E",X"1C",X"3E",X"1F",X"0F",X"07",X"07",X"07",X"07",X"0F",X"DF",X"FC",X"F8",X"F8",X"B2",X"01",
		X"F0",X"F8",X"B8",X"3C",X"7E",X"F2",X"D7",X"DF",X"D7",X"F3",X"FE",X"7E",X"0C",X"5C",X"3C",X"18",
		X"01",X"B2",X"F8",X"F8",X"FC",X"DF",X"0F",X"07",X"07",X"07",X"07",X"0F",X"1F",X"3E",X"1C",X"0E",
		X"8A",X"4E",X"1F",X"3F",X"3F",X"F2",X"F0",X"E0",X"E0",X"E3",X"E7",X"FF",X"FF",X"7D",X"38",X"00",
		X"0F",X"1F",X"1D",X"3C",X"7E",X"3F",X"A7",X"E7",X"A7",X"3F",X"7F",X"7E",X"30",X"B0",X"60",X"80",
		X"00",X"38",X"7D",X"FF",X"FF",X"E7",X"E3",X"E0",X"E0",X"F0",X"F2",X"3F",X"3F",X"1F",X"4E",X"8A",
		X"80",X"60",X"B0",X"30",X"7E",X"7F",X"3F",X"A7",X"E7",X"A7",X"3F",X"7E",X"3C",X"1D",X"1F",X"0F",
		X"00",X"40",X"F8",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"18",X"B8",X"78",X"30",X"00",X"00",
		X"00",X"F0",X"F8",X"BF",X"1F",X"0F",X"0F",X"0F",X"0F",X"0E",X"3E",X"7C",X"38",X"1C",X"00",X"00",
		X"00",X"C0",X"F8",X"FE",X"FF",X"FF",X"FE",X"7C",X"38",X"B8",X"F8",X"F0",X"00",X"00",X"00",X"00",
		X"00",X"07",X"07",X"07",X"07",X"0F",X"DF",X"FC",X"F8",X"F8",X"B2",X"01",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"F8",X"FE",X"FF",X"BF",X"86",X"2E",X"1E",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"03",X"03",X"03",X"03",X"0F",X"1F",X"0E",X"07",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"F8",X"1E",X"0E",X"2E",X"BE",X"7C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"37",X"3F",X"3E",X"3E",X"2C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7C",X"BE",X"2E",X"0F",X"1E",X"F8",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2C",X"3E",X"3E",X"3F",X"37",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"1E",X"2E",X"87",X"BF",X"F3",X"D6",X"D8",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"0E",X"1F",X"0F",X"07",X"03",X"03",X"03",X"03",X"00",
		X"00",X"00",X"00",X"00",X"F0",X"F8",X"B8",X"3C",X"7E",X"F2",X"D7",X"DF",X"D6",X"F0",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"01",X"B2",X"F8",X"F8",X"FC",X"DF",X"0F",X"07",X"07",X"07",X"07",X"00",
		X"00",X"00",X"30",X"78",X"B8",X"1C",X"FC",X"CC",X"5C",X"7C",X"5C",X"CC",X"FC",X"F8",X"40",X"00",
		X"00",X"00",X"1C",X"38",X"7C",X"3E",X"1E",X"0F",X"0F",X"0F",X"0F",X"1F",X"BF",X"F8",X"F0",X"00",
		X"80",X"A0",X"00",X"40",X"80",X"50",X"64",X"E0",X"E0",X"60",X"20",X"30",X"20",X"80",X"00",X"80",
		X"01",X"0F",X"03",X"6E",X"3E",X"7F",X"5E",X"5B",X"46",X"76",X"5F",X"4C",X"0F",X"0B",X"15",X"0B",
		X"C0",X"20",X"80",X"70",X"D4",X"20",X"70",X"F0",X"60",X"30",X"F0",X"E0",X"A0",X"D0",X"40",X"80",
		X"04",X"2B",X"63",X"68",X"63",X"17",X"8D",X"1D",X"1D",X"DF",X"E6",X"D3",X"E1",X"90",X"08",X"16",
		X"E0",X"E0",X"70",X"78",X"FC",X"E4",X"AE",X"BE",X"AE",X"E6",X"FC",X"FC",X"18",X"B8",X"78",X"20",
		X"03",X"25",X"41",X"EC",X"D6",X"BF",X"8F",X"0F",X"0F",X"8F",X"55",X"FE",X"CA",X"AC",X"A0",X"10",
		X"C0",X"30",X"80",X"20",X"40",X"80",X"80",X"00",X"00",X"00",X"00",X"08",X"30",X"00",X"30",X"C0",
		X"07",X"1E",X"30",X"37",X"66",X"7C",X"6C",X"68",X"62",X"6A",X"6D",X"34",X"33",X"10",X"0E",X"07",
		X"80",X"60",X"80",X"20",X"30",X"10",X"10",X"00",X"00",X"10",X"10",X"A0",X"60",X"00",X"E0",X"80",
		X"0F",X"05",X"03",X"0F",X"2C",X"5F",X"56",X"44",X"56",X"5F",X"7F",X"2E",X"2E",X"03",X"1F",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"58",X"E0",X"C8",X"0C",X"C0",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"00",X"03",X"0B",X"17",X"15",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"18",X"40",X"90",X"20",X"40",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0F",X"18",X"1B",X"33",X"3E",X"36",X"34",X"00",
		X"00",X"00",X"00",X"00",X"80",X"60",X"80",X"20",X"30",X"10",X"10",X"00",X"00",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"05",X"03",X"0F",X"2C",X"5F",X"56",X"44",X"56",X"5F",X"7F",X"00",
		X"00",X"00",X"00",X"80",X"60",X"00",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"3C",X"61",X"6E",X"CC",X"F9",X"D9",X"D0",X"C4",X"D4",X"DA",X"68",X"00",
		X"80",X"60",X"00",X"20",X"10",X"00",X"00",X"00",X"00",X"20",X"40",X"80",X"C0",X"E0",X"C0",X"80",
		X"0F",X"1C",X"20",X"66",X"68",X"DA",X"D4",X"C4",X"D0",X"D9",X"F9",X"ED",X"6F",X"77",X"3F",X"0F",
		X"80",X"60",X"00",X"40",X"80",X"00",X"20",X"00",X"00",X"00",X"10",X"80",X"E0",X"60",X"E0",X"80",
		X"0F",X"3C",X"61",X"6E",X"CC",X"F9",X"D9",X"D0",X"C4",X"D4",X"DB",X"6F",X"67",X"3E",X"1C",X"0F",
		X"00",X"30",X"00",X"20",X"40",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"30",X"00",
		X"06",X"12",X"30",X"30",X"02",X"04",X"0C",X"08",X"62",X"62",X"48",X"34",X"33",X"10",X"0E",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"12",X"10",X"10",X"00",X"00",X"00",X"00",X"40",X"60",X"40",X"20",X"01",X"00",X"08",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",
		X"00",X"04",X"20",X"20",X"00",X"00",X"04",X"30",X"80",X"C0",X"80",X"40",X"00",X"00",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1C",X"7E",X"F3",X"C3",X"C0",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"E0",X"F3",X"F3",X"7E",X"1C",
		X"00",X"00",X"B1",X"F9",X"FF",X"FF",X"FF",X"1F",X"1F",X"3F",X"3F",X"3F",X"39",X"31",X"00",X"00",
		X"FE",X"F6",X"F0",X"E0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"E0",X"E0",X"F0",X"F6",X"FE",
		X"00",X"01",X"31",X"39",X"3F",X"3F",X"3F",X"1F",X"1F",X"FF",X"FF",X"FF",X"F9",X"B1",X"01",X"00",
		X"1C",X"7E",X"F3",X"E3",X"90",X"08",X"08",X"08",X"98",X"F8",X"F0",X"E0",X"F3",X"F3",X"7E",X"1C",
		X"00",X"00",X"31",X"39",X"3F",X"3D",X"3D",X"1D",X"1F",X"FF",X"FF",X"FF",X"F9",X"B1",X"00",X"00",
		X"FE",X"F6",X"F0",X"E0",X"90",X"08",X"08",X"08",X"98",X"F8",X"F0",X"E0",X"E0",X"F0",X"F6",X"FE",
		X"00",X"01",X"B1",X"F9",X"FF",X"FD",X"FD",X"1D",X"1F",X"3F",X"3F",X"3F",X"39",X"31",X"01",X"00",
		X"00",X"00",X"8C",X"99",X"FF",X"FF",X"FF",X"BF",X"B8",X"B8",X"FC",X"FC",X"BC",X"9E",X"0E",X"1E",
		X"98",X"7E",X"DF",X"4F",X"07",X"0F",X"19",X"10",X"10",X"10",X"59",X"CF",X"47",X"B7",X"3E",X"0C",
		X"21",X"1F",X"1F",X"BF",X"FF",X"FC",X"FD",X"7D",X"5E",X"5F",X"DA",X"F9",X"B8",X"B8",X"38",X"78",
		X"00",X"1E",X"3F",X"B7",X"47",X"CF",X"5C",X"18",X"18",X"18",X"1C",X"0F",X"47",X"CF",X"7E",X"98",
		X"00",X"C0",X"C0",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"E0",X"F3",X"F3",X"7E",X"1C",X"00",X"00",
		X"00",X"F9",X"FF",X"FF",X"FF",X"1F",X"1F",X"3F",X"3F",X"3F",X"39",X"31",X"00",X"00",X"00",X"00",
		X"00",X"E0",X"F8",X"FC",X"FC",X"FC",X"F8",X"F0",X"F0",X"F8",X"FB",X"7F",X"00",X"00",X"00",X"00",
		X"00",X"1F",X"1F",X"0F",X"0F",X"7F",X"7F",X"7F",X"7C",X"58",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"F8",X"FE",X"FC",X"F8",X"7D",X"7D",X"1F",X"06",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"07",X"0F",X"0F",X"0F",X"0E",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"F8",X"FC",X"3C",X"3C",X"3D",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"1F",X"1F",X"1F",X"1F",X"16",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"3D",X"3C",X"38",X"F2",X"A0",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"16",X"1F",X"1F",X"1F",X"1F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"1F",X"7D",X"79",X"E4",X"42",X"42",X"40",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0E",X"0F",X"0F",X"0F",X"07",X"07",X"00",
		X"00",X"00",X"00",X"00",X"7F",X"FB",X"F8",X"F0",X"C8",X"84",X"84",X"84",X"CC",X"F8",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"58",X"7C",X"7F",X"7E",X"7E",X"0E",X"0F",X"1F",X"1F",X"00",
		X"00",X"00",X"1C",X"7E",X"F3",X"E3",X"90",X"08",X"08",X"08",X"98",X"F8",X"F0",X"E0",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"31",X"39",X"3F",X"3D",X"3D",X"1D",X"1F",X"FF",X"FF",X"FF",X"F9",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"E0",X"60",X"20",X"20",X"60",X"E0",X"C0",X"00",X"00",X"80",X"00",
		X"00",X"82",X"C4",X"FE",X"7F",X"FF",X"7E",X"7C",X"FC",X"7E",X"7F",X"FF",X"7E",X"C3",X"80",X"00",
		X"00",X"00",X"80",X"00",X"F0",X"F8",X"98",X"08",X"08",X"98",X"F8",X"F0",X"80",X"C0",X"00",X"00",
		X"00",X"80",X"D3",X"FF",X"FF",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"D1",X"80",X"00",
		X"00",X"30",X"E0",X"E0",X"90",X"08",X"08",X"08",X"98",X"F8",X"F0",X"E0",X"E0",X"E0",X"30",X"00",
		X"00",X"80",X"F0",X"79",X"7F",X"7D",X"3D",X"3D",X"3F",X"7F",X"7F",X"7F",X"79",X"F0",X"80",X"00",
		X"00",X"00",X"00",X"00",X"80",X"F0",X"98",X"08",X"08",X"98",X"F0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"20",X"38",X"1C",X"7F",X"1F",X"7F",X"3F",X"3F",X"7F",X"1F",X"7F",X"1C",X"38",X"20",X"00",
		X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"40",X"40",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"24",X"4C",X"F8",X"FC",X"7F",X"7F",X"FC",X"78",X"F8",X"FC",X"7F",X"7F",X"7C",X"DC",X"84",X"42",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"13",X"3E",X"3F",X"1F",X"1F",X"3F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"F8",X"CC",X"80",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"1C",X"0E",X"3F",X"0F",X"3F",X"1F",X"1F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"40",X"40",X"C0",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"24",X"4C",X"F8",X"FC",X"7F",X"7F",X"FC",X"78",X"F8",X"FC",X"7F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"30",X"10",X"10",X"30",X"E0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"40",X"70",X"38",X"FF",X"3F",X"FF",X"7E",X"7E",X"FF",X"3F",X"FF",X"38",X"00",
		X"08",X"84",X"EC",X"F8",X"F8",X"F8",X"FC",X"7C",X"78",X"FC",X"F8",X"F8",X"FC",X"7C",X"88",X"90",
		X"01",X"00",X"00",X"00",X"07",X"0F",X"0C",X"08",X"08",X"0C",X"0F",X"07",X"00",X"00",X"00",X"00",
		X"40",X"20",X"64",X"FE",X"FA",X"F9",X"FC",X"7C",X"78",X"FC",X"F8",X"F8",X"75",X"66",X"20",X"10",
		X"00",X"00",X"00",X"00",X"07",X"0F",X"0C",X"08",X"08",X"0C",X"0F",X"07",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"24",X"4C",X"F8",X"FC",X"7B",X"7C",X"E6",X"42",X"C2",X"E6",X"7D",X"7F",X"7C",X"DC",X"84",X"42",
		X"00",X"00",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"80",X"00",
		X"16",X"59",X"7F",X"BE",X"3B",X"12",X"00",X"20",X"A0",X"E0",X"F0",X"79",X"5E",X"33",X"0D",X"05",
		X"00",X"00",X"C0",X"80",X"08",X"00",X"00",X"40",X"00",X"00",X"10",X"80",X"04",X"00",X"00",X"00",
		X"04",X"49",X"34",X"48",X"A3",X"B0",X"20",X"20",X"A0",X"20",X"D0",X"08",X"54",X"33",X"08",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"FC",X"FE",X"E1",X"C0",X"C4",X"F8",X"F8",X"C4",X"C0",X"E1",X"FE",X"FC",X"E0",X"00",X"00",
		X"3F",X"FF",X"07",X"8F",X"FF",X"1F",X"0F",X"07",X"0F",X"3F",X"2F",X"07",X"FF",X"3F",X"00",X"00",
		X"00",X"E0",X"FC",X"E3",X"C0",X"C4",X"F8",X"F8",X"C4",X"C0",X"E3",X"FC",X"E0",X"00",X"00",X"00",
		X"00",X"3F",X"FF",X"2F",X"3F",X"0F",X"0F",X"07",X"1F",X"FF",X"8F",X"FF",X"3F",X"00",X"00",X"00",
		X"E0",X"FC",X"FE",X"E1",X"C0",X"C0",X"F8",X"F8",X"C0",X"C0",X"E1",X"FE",X"FC",X"E0",X"00",X"00",
		X"3F",X"FF",X"07",X"8F",X"FF",X"1F",X"07",X"07",X"0F",X"3F",X"2F",X"07",X"FF",X"3F",X"00",X"00",
		X"00",X"E0",X"FC",X"E3",X"C0",X"C0",X"F8",X"F8",X"C0",X"C0",X"E3",X"FC",X"E0",X"00",X"00",X"00",
		X"00",X"3F",X"FF",X"2F",X"3F",X"0F",X"07",X"07",X"1F",X"FF",X"8F",X"FF",X"3F",X"01",X"00",X"00",
		X"F8",X"FE",X"E0",X"40",X"F0",X"44",X"1C",X"F0",X"E0",X"E0",X"F0",X"D8",X"E8",X"BF",X"5E",X"00",
		X"00",X"0D",X"1C",X"3F",X"60",X"98",X"2E",X"47",X"0F",X"0F",X"03",X"03",X"97",X"7F",X"0F",X"00",
		X"00",X"5C",X"BB",X"EC",X"1A",X"30",X"E0",X"E0",X"F0",X"1C",X"44",X"F0",X"40",X"E0",X"FE",X"F8",
		X"00",X"0F",X"7F",X"97",X"03",X"03",X"0F",X"0F",X"07",X"4E",X"B8",X"60",X"3F",X"1C",X"0D",X"00",
		X"00",X"C0",X"80",X"88",X"F0",X"F0",X"88",X"80",X"C2",X"FC",X"F8",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"9F",X"FF",X"3F",X"1F",X"0F",X"1F",X"7F",X"5F",X"0F",X"FF",X"7F",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"F8",X"F8",X"C4",X"C0",X"E3",X"FC",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"0F",X"07",X"1F",X"FF",X"8F",X"FF",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"E0",X"E0",X"F0",X"FF",X"FE",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"07",X"1F",X"17",X"03",X"7F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"F8",X"FE",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"3F",X"23",X"3F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"FF",X"F8",X"F0",X"F0",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"3F",X"0B",X"0F",X"03",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"FE",X"FF",X"F0",X"E0",X"E0",X"FC",X"F8",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"7F",X"03",X"47",X"7F",X"0F",X"03",X"03",X"07",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"FC",X"E3",X"C0",X"C0",X"F8",X"F8",X"C0",X"C0",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"3F",X"FF",X"2F",X"3F",X"0F",X"07",X"07",X"1F",X"FF",X"8F",X"00",
		X"00",X"00",X"C0",X"F8",X"FC",X"C2",X"80",X"80",X"F0",X"F0",X"80",X"80",X"C2",X"F8",X"C0",X"00",
		X"00",X"00",X"7F",X"FF",X"0F",X"9F",X"FF",X"3F",X"0F",X"0F",X"1F",X"7F",X"5F",X"0F",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"E0",X"FC",X"FF",X"F8",X"F8",X"FF",X"FC",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"3F",X"FF",X"07",X"07",X"FF",X"3F",X"07",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"F8",X"FC",X"C3",X"C0",X"F8",X"F8",X"C3",X"FE",X"FC",X"E0",X"00",X"00",X"00",
		X"00",X"00",X"3F",X"7F",X"EF",X"3F",X"0F",X"07",X"07",X"1F",X"FF",X"7F",X"1F",X"00",X"00",X"00",
		X"00",X"E0",X"FC",X"FE",X"E1",X"C0",X"C0",X"F8",X"F8",X"C1",X"C2",X"FE",X"FC",X"E0",X"00",X"00",
		X"00",X"3F",X"FF",X"07",X"8F",X"FF",X"1F",X"07",X"07",X"0F",X"3F",X"EF",X"7F",X"3F",X"00",X"00",
		X"00",X"00",X"FC",X"F8",X"F6",X"FE",X"FC",X"F8",X"F0",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"07",X"0F",X"1F",X"3F",X"3F",X"7F",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"F0",X"F8",X"FC",X"FE",X"F6",X"F8",X"FC",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"7F",X"7F",X"7F",X"3F",X"3F",X"1F",X"0F",X"07",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"1F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"FE",X"FD",X"FF",X"FE",X"F8",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"0F",X"0F",X"1F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"F0",X"F8",X"F8",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"7F",X"7F",X"3F",X"3F",X"1F",X"00",
		X"00",X"00",X"00",X"00",X"F8",X"F0",X"EC",X"FC",X"F8",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"0F",X"1F",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"F8",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"07",X"1F",X"3F",X"77",X"9F",X"1F",X"2F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"C0",X"F8",X"FC",X"FE",X"FE",X"FF",X"E7",X"F8",X"FC",X"FE",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"2F",X"1F",X"87",X"77",X"3B",X"3F",X"1F",X"07",X"01",X"00",X"00",X"00",
		X"40",X"C0",X"C0",X"80",X"0C",X"3C",X"38",X"C0",X"E0",X"C0",X"00",X"80",X"A0",X"70",X"F0",X"78",
		X"00",X"00",X"03",X"05",X"10",X"37",X"7E",X"79",X"F7",X"FD",X"FE",X"0F",X"07",X"02",X"00",X"00",
		X"C0",X"A0",X"00",X"04",X"08",X"40",X"F0",X"80",X"40",X"30",X"00",X"00",X"C0",X"88",X"20",X"10",
		X"00",X"91",X"25",X"4D",X"38",X"72",X"70",X"C2",X"4B",X"B9",X"B8",X"5C",X"0C",X"02",X"40",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",
		X"00",X"01",X"10",X"40",X"20",X"A0",X"C0",X"58",X"10",X"45",X"90",X"00",X"60",X"28",X"0C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"8A",X"CC",X"9F",X"7F",X"7E",X"40",X"14",X"14",X"5D",X"7F",X"7F",X"9E",X"C0",X"80",X"00",
		X"7F",X"1F",X"0F",X"07",X"07",X"07",X"46",X"00",X"00",X"26",X"07",X"07",X"07",X"0F",X"1F",X"7F",
		X"00",X"14",X"94",X"DD",X"8F",X"7F",X"7E",X"00",X"38",X"7E",X"6F",X"8F",X"CC",X"8A",X"0A",X"00",
		X"00",X"00",X"1F",X"07",X"07",X"07",X"26",X"00",X"00",X"46",X"07",X"07",X"07",X"1F",X"00",X"00",
		X"0A",X"8A",X"CF",X"99",X"79",X"FE",X"C0",X"14",X"14",X"DF",X"F9",X"79",X"9E",X"C0",X"80",X"00",
		X"7F",X"1F",X"0F",X"01",X"00",X"01",X"41",X"00",X"00",X"21",X"01",X"00",X"01",X"0F",X"1F",X"7F",
		X"00",X"14",X"D4",X"9F",X"09",X"F9",X"FE",X"00",X"70",X"FE",X"D9",X"09",X"8F",X"CA",X"0A",X"00",
		X"00",X"00",X"1F",X"07",X"00",X"01",X"21",X"00",X"00",X"41",X"01",X"00",X"07",X"1F",X"00",X"00",
		X"02",X"1C",X"7C",X"F8",X"F0",X"70",X"74",X"20",X"00",X"22",X"70",X"70",X"E0",X"EC",X"F0",X"C0",
		X"40",X"78",X"68",X"58",X"78",X"3B",X"1F",X"0E",X"00",X"1F",X"2F",X"FC",X"2D",X"1B",X"03",X"01",
		X"08",X"F0",X"E0",X"C0",X"70",X"70",X"22",X"00",X"20",X"74",X"70",X"F0",X"F0",X"78",X"3C",X"0F",
		X"00",X"01",X"1B",X"2D",X"FC",X"2F",X"1F",X"00",X"0E",X"1F",X"3B",X"78",X"58",X"68",X"78",X"40",
		X"00",X"00",X"F8",X"FC",X"80",X"28",X"28",X"BA",X"FE",X"FE",X"3C",X"80",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"0E",X"0E",X"4C",X"00",X"00",X"4C",X"0E",X"0E",X"0F",X"1F",X"3F",X"FE",X"00",X"00",
		X"00",X"40",X"78",X"00",X"38",X"7E",X"6F",X"8F",X"CC",X"8A",X"0A",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"26",X"00",X"00",X"46",X"07",X"07",X"07",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"2E",X"BF",X"BF",X"CF",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"13",X"03",X"03",X"03",X"07",X"0F",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"D8",X"E2",X"F3",X"E2",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"01",X"01",X"01",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"F5",X"E7",X"02",X"78",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"01",X"00",X"00",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"85",X"C5",X"E7",X"C9",X"39",X"FF",X"E0",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"0F",X"07",X"00",X"00",X"00",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"14",X"D4",X"9F",X"09",X"F9",X"FE",X"00",X"70",X"F8",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"07",X"00",X"01",X"21",X"00",X"00",X"41",X"01",X"00",
		X"00",X"00",X"14",X"14",X"9E",X"32",X"F2",X"FC",X"80",X"28",X"28",X"BE",X"F2",X"F0",X"00",X"00",
		X"00",X"00",X"FE",X"3F",X"1F",X"03",X"00",X"03",X"43",X"00",X"00",X"03",X"23",X"00",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"44",X"CC",X"8C",X"98",X"08",X"00",X"40",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"02",X"10",X"10",X"33",X"37",X"62",X"4B",X"1C",X"1E",X"06",X"00",X"00",X"00",X"00",
		X"50",X"50",X"48",X"88",X"08",X"92",X"00",X"A0",X"80",X"F8",X"48",X"88",X"F0",X"02",X"00",X"00",
		X"18",X"30",X"1E",X"0C",X"0B",X"65",X"28",X"00",X"20",X"48",X"08",X"03",X"0C",X"56",X"38",X"10",
		X"00",X"28",X"A8",X"3E",X"12",X"F2",X"FC",X"00",X"E0",X"FC",X"B2",X"12",X"1E",X"94",X"14",X"00",
		X"00",X"00",X"17",X"0F",X"40",X"0B",X"03",X"50",X"20",X"23",X"23",X"88",X"0F",X"1F",X"00",X"00",
		X"00",X"38",X"18",X"10",X"80",X"C4",X"CC",X"8C",X"18",X"18",X"00",X"C0",X"C0",X"80",X"00",X"00",
		X"03",X"07",X"02",X"00",X"00",X"31",X"33",X"60",X"48",X"18",X"18",X"00",X"00",X"01",X"01",X"00",
		X"00",X"00",X"80",X"C0",X"C0",X"00",X"18",X"18",X"8C",X"CC",X"C4",X"80",X"10",X"18",X"38",X"00",
		X"00",X"01",X"01",X"00",X"00",X"18",X"18",X"48",X"60",X"33",X"31",X"00",X"00",X"02",X"07",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"18",X"0C",X"0C",X"80",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"CE",X"86",X"04",X"20",X"71",X"F3",X"22",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"0C",X"0C",X"18",X"12",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"60",X"60",X"00",X"0C",X"0C",X"46",X"E0",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0C",X"24",X"30",X"19",X"18",X"00",
		X"00",X"00",X"00",X"38",X"18",X"10",X"80",X"C4",X"CC",X"8C",X"18",X"18",X"00",X"C0",X"C0",X"00",
		X"00",X"00",X"03",X"07",X"02",X"00",X"00",X"31",X"33",X"60",X"48",X"18",X"18",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"40",X"10",X"38",X"10",X"00",X"00",X"00",X"40",X"60",X"00",X"80",X"00",X"00",
		X"00",X"00",X"04",X"1C",X"18",X"02",X"03",X"03",X"19",X"18",X"1C",X"08",X"03",X"03",X"00",X"00",
		X"00",X"00",X"80",X"00",X"60",X"40",X"00",X"00",X"00",X"10",X"38",X"10",X"40",X"C0",X"00",X"00",
		X"00",X"00",X"03",X"03",X"08",X"1C",X"18",X"19",X"03",X"03",X"02",X"18",X"1C",X"04",X"00",X"00",
		X"00",X"00",X"80",X"C0",X"40",X"00",X"08",X"18",X"8C",X"CC",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"08",X"08",X"42",X"63",X"05",X"22",X"00",X"10",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"C0",X"60",X"60",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"04",X"04",X"22",X"40",X"40",X"10",X"1C",X"2C",X"00",X"00",X"80",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"80",X"00",X"10",X"30",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"30",X"80",X"20",X"40",X"80",X"80",X"00",X"00",X"00",X"00",X"08",X"30",X"00",X"30",X"C0",
		X"07",X"1E",X"30",X"37",X"66",X"7C",X"6C",X"68",X"62",X"6A",X"6D",X"34",X"33",X"10",X"0E",X"07",
		X"C0",X"30",X"80",X"20",X"40",X"80",X"80",X"00",X"00",X"00",X"00",X"08",X"30",X"00",X"30",X"C0",
		X"07",X"1E",X"30",X"37",X"66",X"7C",X"6C",X"68",X"62",X"6A",X"6D",X"34",X"33",X"10",X"0E",X"07",
		X"C0",X"30",X"80",X"20",X"40",X"80",X"80",X"00",X"00",X"00",X"00",X"08",X"30",X"00",X"30",X"C0",
		X"07",X"1E",X"30",X"37",X"66",X"7C",X"6C",X"68",X"62",X"6A",X"6D",X"34",X"33",X"10",X"0E",X"07",
		X"C0",X"30",X"80",X"20",X"40",X"80",X"80",X"00",X"00",X"00",X"00",X"08",X"30",X"00",X"30",X"C0",
		X"07",X"1E",X"30",X"37",X"66",X"7C",X"6C",X"68",X"62",X"6A",X"6D",X"34",X"33",X"10",X"0E",X"07",
		X"C0",X"30",X"80",X"20",X"40",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"30",X"C0",
		X"07",X"1E",X"30",X"37",X"66",X"7C",X"6C",X"68",X"62",X"6A",X"6D",X"34",X"33",X"10",X"0E",X"07",
		X"C0",X"20",X"80",X"20",X"40",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"20",X"C0",
		X"07",X"1E",X"30",X"37",X"66",X"7C",X"6C",X"68",X"62",X"6A",X"6D",X"34",X"33",X"10",X"0E",X"07",
		X"C0",X"00",X"80",X"00",X"40",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"07",X"1E",X"30",X"37",X"66",X"7C",X"6C",X"68",X"62",X"6A",X"6D",X"34",X"33",X"10",X"0E",X"07",
		X"80",X"00",X"80",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"07",X"1E",X"30",X"37",X"66",X"7C",X"6C",X"68",X"62",X"6A",X"6D",X"34",X"33",X"10",X"0E",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"1E",X"30",X"37",X"66",X"7C",X"6C",X"68",X"62",X"6A",X"6D",X"34",X"33",X"10",X"0E",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"1E",X"30",X"36",X"66",X"7C",X"6C",X"68",X"62",X"6A",X"6C",X"34",X"32",X"10",X"0E",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"1C",X"30",X"34",X"64",X"7C",X"6C",X"68",X"60",X"68",X"6C",X"34",X"30",X"10",X"0C",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"18",X"30",X"30",X"60",X"78",X"68",X"68",X"60",X"68",X"68",X"30",X"30",X"10",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"30",X"30",X"60",X"70",X"60",X"60",X"60",X"60",X"60",X"30",X"30",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"20",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"20",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"F0",X"98",X"08",X"08",X"98",X"F0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"20",X"38",X"1C",X"7F",X"1F",X"7F",X"3F",X"3F",X"7F",X"1F",X"7F",X"1C",X"38",X"20",X"00",
		X"00",X"00",X"00",X"00",X"80",X"F0",X"98",X"08",X"08",X"98",X"F0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"20",X"38",X"1C",X"7F",X"1F",X"7F",X"3F",X"3F",X"7F",X"1F",X"7F",X"1C",X"38",X"20",X"00",
		X"00",X"00",X"00",X"00",X"80",X"F0",X"98",X"08",X"08",X"98",X"F0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"20",X"38",X"1C",X"7F",X"1F",X"7F",X"3F",X"3F",X"7F",X"1F",X"7F",X"1C",X"38",X"20",X"00",
		X"00",X"00",X"00",X"00",X"80",X"F0",X"98",X"08",X"08",X"98",X"F0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"20",X"38",X"1C",X"7F",X"1F",X"7F",X"3F",X"3F",X"7F",X"1F",X"7F",X"1C",X"38",X"20",X"00",
		X"00",X"00",X"00",X"00",X"80",X"F0",X"90",X"00",X"00",X"90",X"F0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"20",X"38",X"1C",X"7F",X"1F",X"7F",X"3F",X"3F",X"7F",X"1F",X"7F",X"1C",X"38",X"20",X"00",
		X"00",X"00",X"00",X"00",X"80",X"E0",X"80",X"00",X"00",X"80",X"E0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"20",X"38",X"1C",X"7F",X"1F",X"7F",X"3F",X"3F",X"7F",X"1F",X"7F",X"1C",X"38",X"20",X"00",
		X"00",X"00",X"00",X"00",X"80",X"C0",X"80",X"00",X"00",X"80",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"20",X"38",X"1C",X"7F",X"1F",X"7F",X"3F",X"3F",X"7F",X"1F",X"7F",X"1C",X"38",X"20",X"00",
		X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"20",X"38",X"1C",X"7F",X"1F",X"7F",X"3F",X"3F",X"7F",X"1F",X"7F",X"1C",X"38",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"20",X"38",X"1C",X"7F",X"1F",X"7F",X"3F",X"3F",X"7F",X"1F",X"7F",X"1C",X"38",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"20",X"38",X"1C",X"7E",X"1E",X"7E",X"3E",X"3E",X"7E",X"1E",X"7E",X"1C",X"38",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"20",X"38",X"1C",X"7C",X"1C",X"7C",X"3C",X"3C",X"7C",X"1C",X"7C",X"1C",X"38",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"20",X"38",X"18",X"78",X"18",X"78",X"38",X"38",X"78",X"18",X"78",X"18",X"38",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"20",X"30",X"10",X"70",X"10",X"70",X"30",X"30",X"70",X"10",X"70",X"10",X"30",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"20",X"20",X"00",X"60",X"00",X"60",X"20",X"20",X"60",X"00",X"60",X"00",X"20",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"00",X"40",X"00",X"00",X"40",X"00",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FC",X"F8",X"F6",X"FE",X"FC",X"F8",X"F0",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"07",X"0F",X"1F",X"3F",X"3F",X"7F",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FC",X"F8",X"F6",X"FE",X"FC",X"F8",X"F0",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"07",X"0F",X"1F",X"3F",X"3F",X"7F",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FC",X"F8",X"F4",X"FC",X"FC",X"F8",X"F0",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"07",X"0F",X"1F",X"3F",X"3F",X"7F",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F8",X"F8",X"F0",X"F8",X"F8",X"F8",X"F0",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"07",X"0F",X"1F",X"3F",X"3F",X"7F",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"07",X"0F",X"1F",X"3F",X"3F",X"7F",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"07",X"0F",X"1F",X"3F",X"3F",X"7F",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"07",X"0F",X"1F",X"3F",X"3F",X"7F",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"07",X"0F",X"1F",X"3F",X"3F",X"7F",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"07",X"0F",X"1F",X"3F",X"3F",X"7F",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"06",X"0E",X"1E",X"3E",X"3E",X"7E",X"7E",X"7E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"0C",X"1C",X"3C",X"3C",X"7C",X"7C",X"7C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"18",X"38",X"38",X"78",X"78",X"78",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"30",X"70",X"70",X"70",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"60",X"60",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"38",X"18",X"10",X"80",X"C4",X"CC",X"8C",X"18",X"18",X"00",X"C0",X"C0",X"80",X"00",X"00",
		X"03",X"07",X"02",X"00",X"00",X"31",X"33",X"60",X"48",X"18",X"18",X"00",X"00",X"01",X"01",X"00",
		X"00",X"38",X"18",X"10",X"80",X"C4",X"CC",X"8C",X"18",X"18",X"00",X"C0",X"C0",X"80",X"00",X"00",
		X"03",X"07",X"02",X"00",X"00",X"31",X"33",X"60",X"48",X"18",X"18",X"00",X"00",X"01",X"01",X"00",
		X"00",X"38",X"18",X"10",X"80",X"C4",X"CC",X"8C",X"18",X"18",X"00",X"C0",X"C0",X"80",X"00",X"00",
		X"03",X"07",X"02",X"00",X"00",X"31",X"33",X"60",X"48",X"18",X"18",X"00",X"00",X"01",X"01",X"00",
		X"00",X"38",X"18",X"10",X"80",X"C0",X"C8",X"88",X"18",X"18",X"00",X"C0",X"C0",X"80",X"00",X"00",
		X"03",X"07",X"02",X"00",X"00",X"31",X"33",X"60",X"48",X"18",X"18",X"00",X"00",X"01",X"01",X"00",
		X"00",X"30",X"10",X"10",X"80",X"C0",X"C0",X"80",X"10",X"10",X"00",X"C0",X"C0",X"80",X"00",X"00",
		X"03",X"07",X"02",X"00",X"00",X"31",X"33",X"60",X"48",X"18",X"18",X"00",X"00",X"01",X"01",X"00",
		X"00",X"20",X"00",X"00",X"80",X"C0",X"C0",X"80",X"00",X"00",X"00",X"C0",X"C0",X"80",X"00",X"00",
		X"03",X"07",X"02",X"00",X"00",X"31",X"33",X"60",X"48",X"18",X"18",X"00",X"00",X"01",X"01",X"00",
		X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"80",X"00",X"00",X"00",X"C0",X"C0",X"80",X"00",X"00",
		X"03",X"07",X"02",X"00",X"00",X"31",X"33",X"60",X"48",X"18",X"18",X"00",X"00",X"01",X"01",X"00",
		X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"80",X"80",X"80",X"00",X"00",
		X"03",X"07",X"02",X"00",X"00",X"31",X"33",X"60",X"48",X"18",X"18",X"00",X"00",X"01",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"07",X"02",X"00",X"00",X"31",X"33",X"60",X"48",X"18",X"18",X"00",X"00",X"01",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"06",X"02",X"00",X"00",X"30",X"32",X"60",X"48",X"18",X"18",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"00",X"00",X"00",X"30",X"30",X"60",X"48",X"18",X"18",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"30",X"30",X"60",X"48",X"18",X"18",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"30",X"30",X"60",X"40",X"10",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"60",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
