module keyboard(
	input [2:0]	Addr,
	input 		JOY_SEL_n,
	input 		KB_SEL_n,
	output 		Kb_Out,
	input 		RD_n,
	input 		WR_n,
	input 		CON,//not sure
	input  		IORQ_n,
	input  		ps2_kbd_clk,
	input  		ps2_kbd_data
);


endmodule 