library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity bg_graphx_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of bg_graphx_1 is
	type rom is array(0 to  1935) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"8A",X"8A",X"8A",X"8A",X"8A",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"8A",X"8A",X"8A",X"8A",X"8A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",
		X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",
		X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",
		X"60",X"60",X"60",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"60",X"60",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"60",X"60",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"60",X"60",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"00",X"00",X"00",X"8A",X"8A",X"8A",X"8A",X"8A",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"8A",X"8A",X"8A",X"8A",X"8A",X"00",X"00",X"00",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7E",X"12",X"1E",X"00",X"7E",X"5A",X"5A",X"00",
		X"7E",X"12",X"1E",X"00",X"7E",X"12",X"1E",X"00",X"7E",X"5A",X"5A",X"00",X"7E",X"12",X"2E",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"10",X"00",X"22",X"00",X"10",X"04",X"00",X"00",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"00",X"00",X"10",X"00",X"48",X"00",X"00",X"20",X"00",X"08",X"40",X"00",X"10",X"04",
		X"00",X"00",X"00",X"01",X"00",X"10",X"00",X"00",X"02",X"00",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",
		X"02",X"00",X"24",X"00",X"08",X"41",X"04",X"00",X"09",X"01",X"04",X"90",X"04",X"20",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"80",X"00",X"00",X"00",X"00",X"80",X"00",X"10",X"80",X"00",X"00",X"20",X"00",X"80",X"00",
		X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"80",X"04",X"00",X"20",X"05",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",
		X"10",X"00",X"41",X"08",X"00",X"20",X"81",X"00",X"10",X"00",X"00",X"82",X"00",X"04",X"00",X"20",
		X"00",X"00",X"24",X"00",X"04",X"01",X"10",X"00",X"02",X"00",X"00",X"00",X"00",X"01",X"00",X"00",
		X"04",X"40",X"08",X"20",X"02",X"00",X"20",X"04",X"80",X"01",X"08",X"20",X"02",X"00",X"04",X"01",
		X"00",X"00",X"00",X"00",X"01",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",
		X"00",X"00",X"10",X"00",X"04",X"00",X"01",X"00",X"04",X"00",X"00",X"09",X"00",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C6",X"92",X"FE",X"00",X"FE",X"82",X"FE",X"00",X"FE",X"82",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FE",X"92",X"F6",X"00",X"FE",X"82",X"FE",X"00",X"FE",X"82",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"DE",X"92",X"FE",X"00",X"FE",X"82",X"FE",X"00",X"FE",X"82",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"DE",X"92",X"F2",X"00",X"FE",X"82",X"FE",X"00",X"FE",X"82",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"FE",X"00",X"FE",X"82",X"FE",X"00",X"FE",X"82",X"FE",X"00",X"FE",X"82",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"FE",X"00",X"DE",X"92",X"F2",X"00",X"FE",X"82",X"FE",X"00",X"FE",X"82",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"50",X"60",X"F0",X"D4",X"5A",X"88",X"A8",X"50",X"A0",X"CC",X"70",X"78",X"40",X"00",
		X"00",X"00",X"00",X"00",X"01",X"02",X"07",X"04",X"06",X"04",X"03",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"38",X"6E",X"76",X"7F",X"5D",X"7F",X"77",X"7F",X"5E",X"76",X"38",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"F8",X"CC",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"CC",X"F8",X"20",X"10",X"10",X"E0",
		X"30",X"79",X"77",X"EF",X"EF",X"DF",X"DF",X"DF",X"EF",X"EF",X"77",X"79",X"31",X"02",X"01",X"00",
		X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"00",X"00",X"00",X"10",X"5C",X"54",X"74",X"10",X"00",
		X"00",X"00",X"7C",X"20",X"7C",X"64",X"7C",X"00",X"00",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",
		X"00",X"03",X"1F",X"11",X"1B",X"11",X"1F",X"03",X"00",X"00",X"00",X"00",X"00",X"10",X"70",X"80",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"80",X"70",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"00",X"00",X"80",X"60",X"60",X"00",X"00",X"00",
		X"00",X"0C",X"02",X"A2",X"12",X"12",X"0C",X"00",X"00",X"00",X"BE",X"00",X"00",X"BE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"FE",X"00",X"FE",X"82",X"FE",X"00",X"FE",X"82",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"E6",X"B2",X"9E",X"00",X"FE",X"82",X"FE",X"00",X"FE",X"82",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C6",X"92",X"FE",X"00",X"FE",X"82",X"FE",X"00",X"FE",X"82",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"9E",X"92",X"F2",X"00",X"FE",X"82",X"FE",X"00",X"FE",X"82",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"FE",X"00",X"FE",X"82",X"FE",X"00",X"FE",X"82",X"FE",X"00",X"FE",X"82",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E6",X"B2",X"9E",X"00",X"FE",X"82",X"FE",X"00",X"FE",X"82",X"FE",X"00",X"FE",X"82",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"38",X"24",X"FE",X"20",X"00",X"FE",X"82",X"FE",X"00",X"FE",X"82",X"FE",X"00",X"FE",X"82",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"92",X"FE",X"00",X"FE",X"82",X"FE",X"00",X"FE",X"82",X"FE",X"00",X"FE",X"82",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"FE",X"00",X"FE",X"92",X"F6",X"00",X"FE",X"82",X"FE",X"82",X"FE",X"82",X"FE",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
