library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity MOONCR_1K is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of MOONCR_1K is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",X"00",X"02",X"02",X"FE",X"FE",X"42",X"02",X"00",X"00",
		X"62",X"F2",X"BA",X"9A",X"9E",X"CE",X"46",X"00",X"8C",X"DE",X"F2",X"B2",X"92",X"86",X"04",X"00",
		X"08",X"FE",X"FE",X"C8",X"68",X"38",X"18",X"00",X"1C",X"BE",X"A2",X"A2",X"A2",X"E6",X"E4",X"00",
		X"0C",X"9E",X"92",X"92",X"D2",X"7E",X"3C",X"00",X"C0",X"E0",X"B0",X"9E",X"8E",X"C0",X"C0",X"00",
		X"0C",X"6E",X"9A",X"9A",X"B2",X"F2",X"6C",X"00",X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",X"00",
		X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",
		X"44",X"C6",X"82",X"82",X"C6",X"7C",X"38",X"00",X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",
		X"82",X"92",X"92",X"92",X"FE",X"FE",X"00",X"00",X"80",X"90",X"90",X"90",X"90",X"FE",X"FE",X"00",
		X"9E",X"9E",X"92",X"82",X"C6",X"7C",X"38",X"00",X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",
		X"82",X"82",X"FE",X"FE",X"82",X"82",X"00",X"00",X"FC",X"FE",X"02",X"02",X"02",X"06",X"04",X"00",
		X"82",X"C6",X"6E",X"3C",X"18",X"FE",X"FE",X"00",X"02",X"02",X"02",X"02",X"FE",X"FE",X"00",X"00",
		X"FE",X"FE",X"70",X"38",X"70",X"FE",X"FE",X"00",X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",
		X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",X"00",X"70",X"F8",X"88",X"88",X"88",X"FE",X"FE",X"00",
		X"7A",X"FC",X"8E",X"8A",X"82",X"FE",X"7C",X"00",X"72",X"F6",X"9E",X"8C",X"88",X"FE",X"FE",X"00",
		X"0C",X"5E",X"D2",X"92",X"92",X"F6",X"64",X"00",X"80",X"80",X"FE",X"FE",X"80",X"80",X"00",X"00",
		X"FC",X"FE",X"02",X"02",X"02",X"FE",X"FC",X"00",X"F0",X"F8",X"1C",X"0E",X"1C",X"F8",X"F0",X"00",
		X"F8",X"FE",X"1C",X"38",X"1C",X"FE",X"F8",X"00",X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",
		X"C0",X"F0",X"1E",X"1E",X"F0",X"C0",X"00",X"00",X"C2",X"E2",X"F2",X"BA",X"9E",X"8E",X"86",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"F0",X"FB",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"D0",X"00",X"00",
		X"81",X"42",X"24",X"18",X"18",X"24",X"42",X"81",X"00",X"18",X"18",X"18",X"18",X"18",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",X"00",
		X"00",X"28",X"28",X"28",X"28",X"28",X"00",X"00",X"00",X"41",X"FF",X"FF",X"41",X"00",X"68",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"0E",X"0E",X"0C",X"1D",X"3F",X"E1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"1D",X"0C",X"0E",X"0E",X"07",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"06",X"0E",X"1C",X"3E",X"AD",X"E1",X"ED",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E1",X"AD",X"3E",X"1C",X"0E",X"06",X"03",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"0F",X"03",X"01",X"01",X"03",X"FF",X"FC",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",
		X"03",X"07",X"07",X"0F",X"3B",X"F8",X"FB",X"F8",X"E0",X"E0",X"F0",X"FC",X"EE",X"0F",X"EF",X"0F",
		X"FB",X"F8",X"3B",X"0F",X"07",X"07",X"03",X"03",X"EF",X"0F",X"EE",X"FC",X"F0",X"E0",X"E0",X"E0",
		X"01",X"01",X"03",X"0F",X"03",X"01",X"00",X"00",X"E0",X"F0",X"F0",X"F0",X"F0",X"FC",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"29",X"26",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"18",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"2B",X"66",X"C1",X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"48",
		X"46",X"39",X"0A",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"10",X"12",X"0A",X"1D",X"00",X"00",X"04",X"00",X"10",X"04",X"88",X"00",
		X"18",X"20",X"11",X"00",X"02",X"00",X"00",X"00",X"00",X"44",X"20",X"10",X"40",X"20",X"00",X"00",
		X"00",X"40",X"80",X"20",X"40",X"11",X"19",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"16",X"10",X"00",X"18",X"0E",X"06",X"03",X"33",X"20",X"21",X"7E",X"7F",X"09",X"06",X"00",X"10",
		X"33",X"00",X"10",X"38",X"3C",X"66",X"6A",X"31",X"3D",X"3D",X"11",X"3F",X"3E",X"10",X"00",X"40",
		X"11",X"40",X"80",X"20",X"56",X"10",X"7F",X"7F",X"80",X"20",X"40",X"10",X"38",X"3C",X"6E",X"66",
		X"10",X"16",X"00",X"00",X"01",X"09",X"3B",X"0F",X"33",X"11",X"00",X"18",X"0E",X"06",X"03",X"33",
		X"06",X"00",X"0C",X"0C",X"0C",X"0C",X"0C",X"40",X"33",X"00",X"28",X"28",X"7F",X"7E",X"28",X"28",
		X"80",X"23",X"4F",X"1E",X"38",X"00",X"1E",X"07",X"00",X"0C",X"02",X"09",X"00",X"08",X"00",X"20",
		X"00",X"08",X"04",X"06",X"03",X"7F",X"7F",X"00",X"40",X"10",X"26",X"0C",X"18",X"7F",X"7F",X"00",
		X"00",X"00",X"00",X"03",X"06",X"2D",X"1F",X"0F",X"20",X"40",X"C8",X"FC",X"FE",X"F4",X"F0",X"F8",
		X"1F",X"1F",X"4D",X"37",X"07",X"0D",X"07",X"02",X"FC",X"FC",X"FA",X"F0",X"F4",X"DC",X"08",X"20",
		X"00",X"00",X"00",X"00",X"05",X"03",X"07",X"07",X"00",X"00",X"00",X"00",X"20",X"80",X"E0",X"C0",
		X"07",X"07",X"02",X"09",X"00",X"00",X"00",X"00",X"E0",X"E0",X"D0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"20",X"10",X"0D",X"07",X"03",X"00",X"00",X"08",X"10",X"40",X"84",X"F8",X"C0",
		X"09",X"35",X"46",X"05",X"08",X"00",X"00",X"00",X"80",X"C0",X"A0",X"80",X"40",X"40",X"00",X"00",
		X"10",X"88",X"04",X"21",X"01",X"0F",X"E7",X"3F",X"14",X"84",X"18",X"30",X"D0",X"C0",X"E0",X"F0",
		X"0F",X"0F",X"17",X"07",X"47",X"0D",X"10",X"20",X"FC",X"F3",X"F0",X"F4",X"B0",X"50",X"08",X"04",
		X"3C",X"42",X"81",X"A5",X"A5",X"99",X"42",X"3C",X"20",X"10",X"0E",X"10",X"20",X"0E",X"14",X"24",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"14",X"0E",X"00",X"3E",X"10",X"08",X"10",X"3E",
		X"01",X"02",X"06",X"0C",X"1C",X"19",X"3B",X"37",X"80",X"40",X"20",X"00",X"00",X"80",X"00",X"A0",
		X"37",X"3B",X"19",X"1C",X"0C",X"06",X"02",X"01",X"A0",X"00",X"80",X"00",X"00",X"20",X"40",X"80",
		X"00",X"01",X"07",X"0E",X"1E",X"1D",X"3B",X"3F",X"40",X"A0",X"10",X"00",X"00",X"80",X"C0",X"00",
		X"37",X"33",X"31",X"18",X"08",X"08",X"05",X"06",X"A0",X"00",X"80",X"00",X"00",X"80",X"00",X"00",
		X"00",X"00",X"03",X"0F",X"1E",X"3D",X"3B",X"3F",X"00",X"30",X"E8",X"88",X"08",X"80",X"C0",X"80",
		X"37",X"32",X"31",X"30",X"10",X"12",X"1C",X"00",X"80",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"0F",X"1F",X"1D",X"3B",X"3F",X"00",X"00",X"FC",X"E4",X"04",X"84",X"C0",X"A0",
		X"37",X"32",X"31",X"20",X"20",X"3C",X"00",X"00",X"80",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"0F",X"1F",X"1D",X"3B",X"37",X"00",X"00",X"F0",X"FE",X"02",X"82",X"C4",X"A0",
		X"37",X"22",X"60",X"40",X"78",X"00",X"00",X"00",X"80",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"0F",X"1F",X"3D",X"3B",X"67",X"00",X"00",X"E0",X"F0",X"1C",X"83",X"C1",X"E2",
		X"46",X"82",X"40",X"20",X"00",X"00",X"00",X"00",X"A4",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"0F",X"1E",X"39",X"63",X"87",X"00",X"00",X"C0",X"F0",X"78",X"9C",X"C6",X"E1",
		X"85",X"40",X"21",X"00",X"00",X"00",X"00",X"00",X"A1",X"02",X"84",X"00",X"00",X"00",X"00",X"00",
		X"01",X"02",X"06",X"0C",X"1C",X"19",X"3B",X"37",X"80",X"40",X"20",X"00",X"00",X"80",X"00",X"80",
		X"37",X"3B",X"19",X"1C",X"0C",X"06",X"02",X"01",X"80",X"00",X"80",X"00",X"00",X"20",X"40",X"80",
		X"00",X"01",X"02",X"06",X"0C",X"0C",X"1D",X"1B",X"00",X"80",X"40",X"00",X"00",X"00",X"80",X"80",
		X"1B",X"1D",X"0C",X"0C",X"06",X"02",X"01",X"00",X"80",X"80",X"00",X"00",X"00",X"40",X"80",X"00",
		X"00",X"00",X"01",X"02",X"04",X"0C",X"1D",X"1B",X"00",X"00",X"80",X"40",X"00",X"00",X"80",X"80",
		X"1B",X"1D",X"0C",X"04",X"02",X"01",X"00",X"00",X"80",X"80",X"00",X"00",X"40",X"80",X"00",X"00",
		X"00",X"00",X"00",X"01",X"02",X"06",X"0D",X"0F",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",
		X"0F",X"0D",X"06",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"02",X"04",X"0F",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",
		X"0F",X"04",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",
		X"07",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"07",X"0C",X"00",X"03",X"0F",X"1C",X"30",X"61",X"63",X"C3",
		X"08",X"10",X"30",X"20",X"1C",X"08",X"05",X"09",X"C7",X"AF",X"07",X"31",X"7C",X"7E",X"FF",X"FF",
		X"08",X"18",X"38",X"1D",X"0E",X"03",X"00",X"00",X"F7",X"7F",X"FF",X"F3",X"7F",X"9F",X"FB",X"2C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0E",X"1F",X"0F",X"06",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"18",X"0D",X"C2",X"24",
		X"00",X"02",X"02",X"01",X"00",X"01",X"01",X"02",X"62",X"27",X"10",X"E6",X"9A",X"1C",X"68",X"20",
		X"05",X"04",X"02",X"01",X"00",X"01",X"01",X"01",X"C1",X"20",X"18",X"08",X"C8",X"C4",X"FF",X"8A",
		X"01",X"06",X"08",X"00",X"00",X"00",X"00",X"00",X"72",X"11",X"20",X"20",X"13",X"0C",X"00",X"00",
		X"00",X"00",X"01",X"02",X"04",X"09",X"19",X"19",X"00",X"00",X"80",X"F3",X"7F",X"FF",X"FF",X"DF",
		X"1B",X"07",X"07",X"09",X"0F",X"0F",X"05",X"0D",X"37",X"8F",X"C7",X"82",X"01",X"87",X"E1",X"F9",
		X"0E",X"07",X"07",X"0B",X"0F",X"3F",X"7F",X"3D",X"FF",X"7F",X"EF",X"F6",X"74",X"8D",X"8B",X"8E",
		X"3D",X"19",X"33",X"07",X"07",X"01",X"00",X"00",X"DF",X"F7",X"FB",X"DF",X"8B",X"8B",X"04",X"02",
		X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"04",X"A8",X"08",X"10",X"05",X"02",
		X"01",X"00",X"00",X"28",X"02",X"00",X"00",X"00",X"01",X"06",X"4F",X"AF",X"6F",X"BF",X"BF",X"7F",
		X"02",X"0C",X"88",X"20",X"00",X"00",X"00",X"02",X"7F",X"7F",X"3A",X"1D",X"2F",X"84",X"03",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"16",X"09",X"17",X"20",X"00",X"80",X"00",
		X"00",X"10",X"FB",X"7D",X"30",X"11",X"80",X"38",X"00",X"00",X"00",X"80",X"40",X"20",X"10",X"10",
		X"DE",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"08",X"08",X"14",X"94",X"28",X"48",X"90",X"B8",
		X"FF",X"E2",X"78",X"FE",X"FF",X"FF",X"99",X"FC",X"7C",X"68",X"10",X"01",X"48",X"F0",X"C0",X"80",
		X"3D",X"39",X"19",X"C2",X"24",X"18",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"61",X"13",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"12",X"04",X"F1",X"52",X"31",X"36",X"05",X"84",X"C0",X"20",X"A0",X"60",X"30",X"48",X"48",X"90",
		X"40",X"21",X"22",X"40",X"20",X"C8",X"0C",X"02",X"60",X"F8",X"30",X"28",X"14",X"18",X"30",X"60",
		X"33",X"4F",X"E3",X"A4",X"28",X"10",X"00",X"00",X"70",X"D0",X"10",X"0C",X"04",X"00",X"00",X"00",
		X"00",X"0C",X"32",X"47",X"9F",X"EF",X"9F",X"FF",X"00",X"60",X"60",X"50",X"04",X"CE",X"BE",X"78",
		X"9C",X"2C",X"74",X"F8",X"F1",X"A3",X"0F",X"CF",X"76",X"6A",X"FC",X"E0",X"E0",X"C0",X"C0",X"E0",
		X"EF",X"EF",X"7F",X"2F",X"8F",X"9F",X"3F",X"7E",X"E0",X"D0",X"F0",X"F8",X"F8",X"F0",X"A4",X"80",
		X"6F",X"3F",X"DF",X"F8",X"31",X"30",X"C0",X"00",X"88",X"F0",X"F0",X"E0",X"E0",X"C0",X"00",X"00",
		X"00",X"01",X"00",X"02",X"04",X"01",X"84",X"20",X"00",X"20",X"00",X"40",X"00",X"00",X"00",X"00",
		X"22",X"90",X"C1",X"35",X"F8",X"F6",X"7E",X"F8",X"00",X"80",X"20",X"10",X"62",X"10",X"00",X"00",
		X"F8",X"FC",X"ED",X"BC",X"C8",X"74",X"0A",X"02",X"00",X"00",X"40",X"10",X"00",X"40",X"20",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"40",X"02",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"00",X"07",X"00",X"01",X"7F",X"08",X"30",X"C0",X"18",X"E0",X"0C",X"D8",X"00",
		X"01",X"00",X"07",X"00",X"03",X"00",X"00",X"00",X"C0",X"0C",X"E0",X"18",X"C0",X"30",X"08",X"00",
		X"00",X"01",X"00",X"02",X"01",X"61",X"1F",X"03",X"00",X"00",X"D8",X"20",X"CC",X"30",X"CC",X"C0",
		X"01",X"0C",X"03",X"0C",X"03",X"00",X"00",X"00",X"98",X"00",X"D8",X"40",X"20",X"80",X"40",X"00",
		X"00",X"00",X"00",X"21",X"18",X"04",X"02",X"01",X"00",X"00",X"20",X"98",X"46",X"30",X"CC",X"E0",
		X"0D",X"02",X"09",X"04",X"02",X"02",X"01",X"00",X"CC",X"B0",X"00",X"A0",X"90",X"40",X"00",X"00",
		X"00",X"00",X"00",X"10",X"08",X"04",X"02",X"01",X"00",X"00",X"00",X"20",X"90",X"4C",X"A2",X"D8",
		X"0B",X"05",X"12",X"09",X"05",X"04",X"02",X"00",X"84",X"00",X"28",X"14",X"20",X"90",X"00",X"00",
		X"00",X"00",X"10",X"08",X"08",X"04",X"02",X"11",X"00",X"00",X"00",X"00",X"A0",X"90",X"4C",X"A2",
		X"13",X"0B",X"25",X"14",X"12",X"0A",X"08",X"00",X"D8",X"84",X"50",X"48",X"80",X"80",X"00",X"00",
		X"00",X"04",X"04",X"02",X"02",X"02",X"13",X"4F",X"00",X"00",X"00",X"00",X"50",X"50",X"28",X"A8",
		X"2B",X"2B",X"24",X"24",X"2A",X"0A",X"00",X"00",X"A4",X"32",X"08",X"50",X"50",X"00",X"00",X"00",
		X"00",X"01",X"01",X"01",X"01",X"09",X"29",X"2B",X"00",X"00",X"00",X"00",X"00",X"20",X"28",X"A8",
		X"2B",X"2B",X"48",X"51",X"95",X"04",X"00",X"00",X"A8",X"A8",X"24",X"04",X"42",X"40",X"00",X"00",
		X"00",X"00",X"03",X"00",X"07",X"00",X"00",X"00",X"08",X"30",X"C0",X"18",X"E0",X"0C",X"00",X"18",
		X"00",X"00",X"07",X"00",X"03",X"00",X"00",X"00",X"00",X"0C",X"E0",X"18",X"C0",X"30",X"08",X"00",
		X"00",X"00",X"06",X"00",X"0D",X"00",X"00",X"00",X"04",X"18",X"C0",X"0C",X"B2",X"28",X"00",X"00",
		X"00",X"00",X"0D",X"00",X"06",X"00",X"00",X"00",X"00",X"28",X"B2",X"0C",X"C0",X"18",X"04",X"00",
		X"00",X"08",X"04",X"80",X"0A",X"00",X"00",X"00",X"0C",X"50",X"86",X"09",X"50",X"84",X"00",X"0A",
		X"00",X"00",X"0A",X"10",X"04",X"08",X"00",X"00",X"00",X"84",X"50",X"09",X"86",X"50",X"0C",X"02",
		X"10",X"08",X"20",X"16",X"00",X"00",X"00",X"00",X"50",X"82",X"0C",X"20",X"12",X"00",X"00",X"05",
		X"00",X"00",X"00",X"16",X"20",X"08",X"10",X"00",X"00",X"00",X"12",X"20",X"0C",X"82",X"50",X"00",
		X"08",X"48",X"14",X"00",X"00",X"00",X"00",X"00",X"82",X"0C",X"31",X"00",X"00",X"00",X"00",X"02",
		X"00",X"00",X"00",X"00",X"04",X"48",X"08",X"10",X"00",X"00",X"00",X"00",X"31",X"0C",X"82",X"00",
		X"60",X"24",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"30",X"02",X"00",X"00",X"00",X"00",X"05",
		X"00",X"00",X"00",X"00",X"00",X"24",X"60",X"00",X"00",X"00",X"00",X"00",X"02",X"30",X"06",X"01",
		X"20",X"84",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"10",X"00",X"04",X"00",X"00",X"00",X"0A",
		X"00",X"00",X"00",X"00",X"00",X"84",X"20",X"40",X"00",X"00",X"00",X"04",X"00",X"10",X"20",X"04",
		X"04",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"00",X"00",X"14",
		X"00",X"00",X"00",X"00",X"40",X"00",X"04",X"00",X"00",X"00",X"08",X"00",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"0A",X"14",X"00",X"21",X"EA",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"02",X"14",X"00",X"20",X"00",X"01",X"94",X"80",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"04",
		X"00",X"00",X"00",X"00",X"10",X"02",X"01",X"08",X"10",X"00",X"41",X"08",X"40",X"00",X"00",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"08",X"10",X"00",X"80",
		X"00",X"00",X"00",X"20",X"04",X"02",X"00",X"10",X"01",X"10",X"00",X"80",X"00",X"00",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"08",X"10",X"00",X"80",X"00",X"01",
		X"40",X"00",X"00",X"02",X"00",X"00",X"20",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"08",X"00",X"80",X"00",X"00",X"00",X"21",X"00",
		X"00",X"08",X"00",X"00",X"01",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"80",X"00",X"00",X"01",X"40",X"00",X"00",
		X"00",X"00",X"00",X"02",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"05",X"2F",X"3C",X"7F",X"37",X"66",X"00",X"90",X"34",X"BE",X"F4",X"F4",X"FA",X"7F",
		X"FC",X"7C",X"7F",X"3F",X"5F",X"2F",X"14",X"02",X"3E",X"0C",X"20",X"94",X"FA",X"FE",X"64",X"40",
		X"00",X"02",X"02",X"17",X"0F",X"3E",X"1B",X"33",X"00",X"C0",X"80",X"D4",X"FE",X"F4",X"FA",X"1F",
		X"7E",X"3E",X"1F",X"1F",X"0F",X"14",X"02",X"00",X"16",X"20",X"94",X"F8",X"FC",X"68",X"40",X"00",
		X"00",X"00",X"02",X"03",X"0F",X"07",X"1D",X"19",X"00",X"00",X"C0",X"C8",X"FC",X"F8",X"74",X"FE",
		X"3F",X"1E",X"1F",X"0F",X"04",X"02",X"00",X"00",X"2C",X"40",X"28",X"F0",X"50",X"40",X"00",X"00",
		X"00",X"00",X"00",X"02",X"05",X"03",X"0F",X"0D",X"00",X"00",X"00",X"80",X"90",X"F8",X"E0",X"3C",
		X"0F",X"07",X"0B",X"02",X"01",X"00",X"00",X"00",X"40",X"20",X"F8",X"50",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"05",X"00",X"00",X"00",X"40",X"90",X"F0",X"F0",X"18",
		X"07",X"03",X"00",X"01",X"00",X"00",X"00",X"00",X"50",X"E0",X"D0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"03",X"03",X"00",X"00",X"00",X"00",X"40",X"E0",X"E0",X"B0",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"C0",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"A0",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"01",X"07",X"06",X"00",X"00",X"C0",X"C0",X"B0",X"70",X"60",X"00",
		X"00",X"06",X"07",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"60",X"70",X"B0",X"C0",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"07",X"06",X"00",X"00",X"00",X"60",X"E0",X"D8",X"B8",X"20",X"00",
		X"0C",X"0C",X"02",X"02",X"03",X"01",X"01",X"00",X"00",X"00",X"C0",X"E0",X"60",X"80",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"00",X"00",X"00",X"00",X"38",X"70",X"C8",X"3C",X"38",
		X"0C",X"0E",X"02",X"07",X"06",X"07",X"02",X"00",X"00",X"00",X"80",X"C0",X"C0",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"06",X"00",X"00",X"00",X"00",X"38",X"FC",X"80",X"38",
		X"06",X"06",X"0D",X"0D",X"0D",X"04",X"00",X"00",X"3C",X"00",X"80",X"80",X"80",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"C0",X"DC",X"7E",
		X"06",X"04",X"0C",X"1B",X"1B",X"17",X"12",X"00",X"14",X"38",X"1C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"60",X"64",X"3E",
		X"02",X"0E",X"3D",X"3B",X"06",X"06",X"00",X"00",X"0E",X"18",X"1C",X"0C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"1E",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"3C",
		X"38",X"36",X"0E",X"0C",X"00",X"00",X"00",X"00",X"0E",X"36",X"38",X"18",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"01",X"07",X"06",X"00",X"00",X"C0",X"C0",X"B0",X"70",X"60",X"00",
		X"00",X"06",X"07",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"60",X"70",X"B0",X"C0",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"07",X"06",X"00",X"00",X"00",X"C0",X"C0",X"B0",X"60",X"00",
		X"00",X"06",X"07",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"60",X"B0",X"C0",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"06",X"00",X"00",X"00",X"00",X"C0",X"A0",X"60",X"00",
		X"00",X"06",X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"A0",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"02",X"00",X"00",X"00",X"00",X"C0",X"A0",X"60",X"00",
		X"00",X"02",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"A0",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"02",X"00",X"00",X"00",X"00",X"80",X"40",X"80",X"00",
		X"00",X"02",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"80",
		X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"80",X"B0",X"A0",X"A0",X"A0",X"A0",X"A0",X"FE",X"02",X"1A",X"0A",X"0A",X"0A",X"0A",X"0A",
		X"A0",X"A0",X"A0",X"A0",X"B0",X"80",X"FF",X"00",X"0A",X"0A",X"0A",X"0A",X"1A",X"02",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"2D",X"00",X"00",X"00",X"00",X"00",X"10",X"38",X"40",
		X"2D",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"38",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0A",X"00",X"00",X"00",X"00",X"00",X"08",X"1C",X"A0",
		X"0A",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"1C",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"04",X"0C",X"50",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"0C",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"46",X"A8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A8",X"46",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"23",X"34",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"34",X"23",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"1A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1A",X"11",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"38",X"44",X"7C",X"00",X"7C",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"7C",X"00",X"54",X"54",X"7C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"1E",X"21",X"D1",X"19",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"19",X"D1",X"21",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"1C",X"22",X"D2",X"1A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1A",X"D2",X"22",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"38",X"44",X"A4",X"34",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"34",X"A4",X"44",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"30",X"48",X"88",X"68",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"68",X"88",X"48",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"50",X"90",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"50",X"90",X"50",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"60",X"A0",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"A0",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"A0",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"A0",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
