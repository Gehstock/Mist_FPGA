library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_1J is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_1J is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"3E",X"00",X"32",X"00",X"B0",X"3E",X"00",X"32",X"00",X"9E",X"3E",X"01",X"32",X"00",X"B8",X"31",
		X"00",X"90",X"C3",X"20",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F5",X"3E",X"00",X"32",X"00",X"B0",X"F1",X"C3",X"C0",X"01",
		X"00",X"10",X"00",X"20",X"00",X"30",X"00",X"50",X"00",X"40",X"80",X"8F",X"00",X"8F",X"80",X"8E",
		X"00",X"8E",X"80",X"8D",X"05",X"00",X"20",X"20",X"20",X"20",X"40",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"05",X"00",X"00",X"00",X"00",X"00",X"20",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"05",X"FF",X"40",
		X"40",X"40",X"40",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C3",X"AD",X"01",X"C3",X"18",X"07",X"C3",X"92",X"01",X"C3",X"64",X"08",X"C3",X"50",X"08",X"C3",
		X"1D",X"0B",X"C3",X"41",X"0B",X"C3",X"21",X"0A",X"C3",X"FD",X"09",X"C3",X"82",X"0A",X"C3",X"98",
		X"0A",X"C3",X"EE",X"09",X"C3",X"AC",X"0B",X"C3",X"18",X"06",X"C3",X"B0",X"0B",X"C3",X"E4",X"0B",
		X"C3",X"F2",X"0B",X"C3",X"01",X"0C",X"C3",X"42",X"0C",X"C3",X"4C",X"0C",X"C3",X"0F",X"60",X"C3",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CD",X"C7",X"03",X"CD",X"20",X"07",X"31",X"00",X"90",X"21",X"00",X"80",X"01",X"00",X"08",X"CD",
		X"50",X"08",X"21",X"00",X"88",X"01",X"F6",X"07",X"CD",X"50",X"08",X"21",X"00",X"90",X"01",X"FF",
		X"03",X"CD",X"5A",X"08",X"21",X"00",X"94",X"01",X"FF",X"03",X"CD",X"50",X"08",X"21",X"20",X"98",
		X"01",X"60",X"00",X"CD",X"50",X"08",X"21",X"00",X"9C",X"01",X"00",X"01",X"CD",X"50",X"08",X"21",
		X"00",X"9A",X"01",X"C8",X"00",X"CD",X"50",X"08",X"3E",X"01",X"32",X"00",X"87",X"3E",X"01",X"32",
		X"01",X"87",X"3A",X"04",X"B0",X"32",X"13",X"80",X"3A",X"05",X"B0",X"32",X"14",X"80",X"CD",X"B9",
		X"02",X"CD",X"08",X"09",X"CD",X"18",X"06",X"3E",X"01",X"32",X"8C",X"80",X"21",X"01",X"00",X"22",
		X"22",X"80",X"3E",X"00",X"32",X"00",X"B0",X"3E",X"FF",X"32",X"02",X"80",X"31",X"00",X"90",X"3E",
		X"00",X"32",X"03",X"80",X"21",X"84",X"00",X"CD",X"68",X"03",X"C3",X"05",X"02",X"3E",X"00",X"32",
		X"00",X"B0",X"3E",X"00",X"32",X"03",X"80",X"21",X"90",X"00",X"CD",X"68",X"03",X"C3",X"05",X"02",
		X"F5",X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",X"CD",X"9F",X"02",X"31",X"00",X"90",X"00",X"00",
		X"00",X"CD",X"58",X"09",X"CD",X"AB",X"09",X"CD",X"1B",X"60",X"CD",X"12",X"60",X"CD",X"82",X"03",
		X"CD",X"2F",X"06",X"CD",X"D9",X"5F",X"CD",X"BD",X"02",X"CD",X"64",X"08",X"CD",X"E2",X"09",X"3A",
		X"77",X"80",X"B7",X"20",X"05",X"CD",X"65",X"03",X"18",X"0B",X"3E",X"00",X"32",X"03",X"80",X"21",
		X"84",X"00",X"CD",X"68",X"03",X"3A",X"03",X"80",X"B7",X"C2",X"47",X"02",X"3E",X"FF",X"32",X"02",
		X"80",X"3E",X"00",X"32",X"00",X"B0",X"3E",X"01",X"32",X"00",X"B0",X"06",X"05",X"0E",X"00",X"21",
		X"0E",X"80",X"7E",X"E6",X"30",X"C2",X"2E",X"02",X"7E",X"E6",X"C0",X"C2",X"35",X"02",X"23",X"0C",
		X"10",X"F0",X"C3",X"16",X"02",X"3E",X"00",X"32",X"00",X"B0",X"32",X"02",X"80",X"79",X"32",X"00",
		X"80",X"7E",X"E6",X"80",X"CA",X"68",X"02",X"2A",X"00",X"80",X"29",X"11",X"04",X"80",X"19",X"5E",
		X"23",X"56",X"EB",X"F9",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"3E",X"00",X"32",X"00",X"B0",
		X"3E",X"01",X"32",X"00",X"B0",X"F1",X"ED",X"45",X"36",X"80",X"2A",X"00",X"80",X"29",X"11",X"7A",
		X"00",X"19",X"5E",X"23",X"56",X"EB",X"F9",X"2A",X"00",X"80",X"29",X"11",X"70",X"00",X"19",X"5E",
		X"23",X"56",X"EB",X"3E",X"00",X"32",X"00",X"B0",X"3E",X"01",X"32",X"00",X"B0",X"E9",X"3E",X"00",
		X"32",X"00",X"B0",X"2A",X"00",X"80",X"11",X"0E",X"80",X"19",X"CB",X"BE",X"C3",X"05",X"02",X"3A",
		X"02",X"80",X"FE",X"FF",X"C8",X"2A",X"00",X"80",X"29",X"11",X"04",X"80",X"19",X"EB",X"21",X"00",
		X"00",X"39",X"23",X"23",X"EB",X"73",X"23",X"72",X"C9",X"CD",X"D0",X"5F",X"C9",X"3A",X"02",X"B0",
		X"E6",X"01",X"C2",X"D0",X"02",X"DD",X"21",X"15",X"80",X"26",X"00",X"CD",X"EE",X"02",X"18",X"05",
		X"3E",X"01",X"32",X"15",X"80",X"3A",X"02",X"B0",X"E6",X"02",X"C2",X"E8",X"02",X"DD",X"21",X"82",
		X"80",X"26",X"01",X"CD",X"EE",X"02",X"18",X"05",X"3E",X"01",X"32",X"82",X"80",X"C9",X"DD",X"7E",
		X"00",X"FE",X"00",X"28",X"6F",X"3A",X"17",X"80",X"32",X"90",X"80",X"7C",X"FE",X"00",X"28",X"17",
		X"3A",X"84",X"80",X"FE",X"FF",X"20",X"10",X"3A",X"85",X"80",X"3C",X"32",X"85",X"80",X"FE",X"02",
		X"38",X"4E",X"3E",X"00",X"32",X"85",X"80",X"DD",X"46",X"01",X"3A",X"17",X"80",X"FE",X"99",X"D2",
		X"33",X"03",X"3A",X"17",X"80",X"C6",X"01",X"27",X"32",X"17",X"80",X"05",X"78",X"FE",X"00",X"20",
		X"E9",X"18",X"07",X"3A",X"87",X"80",X"80",X"32",X"87",X"80",X"DD",X"36",X"00",X"00",X"3A",X"70",
		X"80",X"B7",X"C0",X"CD",X"F0",X"00",X"3E",X"10",X"CD",X"FC",X"00",X"3A",X"81",X"80",X"B7",X"28",
		X"07",X"3A",X"90",X"80",X"FE",X"01",X"20",X"0C",X"3E",X"00",X"32",X"03",X"80",X"C3",X"C6",X"00",
		X"DD",X"36",X"00",X"00",X"C9",X"21",X"9D",X"00",X"11",X"0E",X"80",X"46",X"23",X"7E",X"FE",X"FF",
		X"28",X"08",X"23",X"7E",X"12",X"13",X"10",X"FA",X"18",X"07",X"23",X"1A",X"B6",X"12",X"13",X"10",
		X"F9",X"C9",X"F5",X"C5",X"E5",X"21",X"18",X"80",X"3A",X"27",X"80",X"47",X"3A",X"70",X"80",X"B7",
		X"C2",X"98",X"03",X"3A",X"7A",X"80",X"18",X"0A",X"3A",X"00",X"B0",X"CB",X"40",X"28",X"03",X"C3",
		X"E0",X"0F",X"01",X"00",X"05",X"1F",X"30",X"15",X"CB",X"16",X"F5",X"7E",X"FE",X"03",X"28",X"07",
		X"F1",X"23",X"30",X"0B",X"34",X"18",X"09",X"F1",X"23",X"36",X"FF",X"18",X"03",X"71",X"23",X"71",
		X"23",X"10",X"E2",X"E1",X"C1",X"F1",X"C9",X"3E",X"00",X"32",X"8F",X"80",X"CD",X"18",X"06",X"3E",
		X"01",X"32",X"8C",X"80",X"CD",X"AB",X"09",X"21",X"20",X"98",X"01",X"60",X"00",X"CD",X"CC",X"00",
		X"21",X"00",X"90",X"01",X"00",X"04",X"CD",X"CC",X"00",X"21",X"00",X"94",X"01",X"00",X"04",X"CD",
		X"CC",X"00",X"21",X"62",X"C6",X"11",X"C0",X"9C",X"01",X"40",X"00",X"ED",X"B0",X"CD",X"CF",X"00",
		X"B8",X"C5",X"16",X"CD",X"CF",X"00",X"A2",X"C6",X"08",X"FD",X"21",X"56",X"C3",X"FD",X"6E",X"00",
		X"FD",X"66",X"01",X"AF",X"4F",X"57",X"5F",X"06",X"08",X"7E",X"0F",X"30",X"07",X"1C",X"20",X"04",
		X"14",X"20",X"01",X"0C",X"C3",X"10",X"1F",X"E6",X"10",X"C2",X"39",X"05",X"10",X"EC",X"23",X"FD",
		X"7E",X"02",X"BD",X"20",X"E2",X"FD",X"7E",X"03",X"BC",X"20",X"DC",X"CD",X"6C",X"05",X"FD",X"7E",
		X"0C",X"FD",X"A6",X"0D",X"FE",X"FF",X"28",X"07",X"11",X"0C",X"00",X"FD",X"19",X"18",X"BE",X"FD",
		X"21",X"94",X"C3",X"FD",X"6E",X"00",X"FD",X"66",X"01",X"C3",X"20",X"1F",X"E6",X"10",X"C2",X"39",
		X"05",X"3E",X"FF",X"AE",X"77",X"23",X"7D",X"FD",X"BE",X"02",X"20",X"ED",X"7C",X"FD",X"BE",X"03",
		X"20",X"E7",X"FD",X"6E",X"00",X"FD",X"66",X"01",X"11",X"00",X"00",X"D9",X"11",X"00",X"00",X"D9",
		X"06",X"08",X"7E",X"0F",X"30",X"03",X"13",X"18",X"03",X"D9",X"13",X"D9",X"10",X"F5",X"23",X"FD",
		X"7E",X"02",X"BD",X"20",X"EB",X"C3",X"20",X"3F",X"BC",X"20",X"E5",X"FD",X"6E",X"00",X"FD",X"66",
		X"01",X"C3",X"30",X"1F",X"E6",X"10",X"C2",X"39",X"05",X"3E",X"FF",X"AE",X"77",X"23",X"7D",X"FD",
		X"BE",X"02",X"20",X"ED",X"7C",X"FD",X"BE",X"03",X"20",X"E7",X"FD",X"6E",X"00",X"FD",X"66",X"01",
		X"06",X"08",X"7E",X"0F",X"30",X"03",X"13",X"18",X"03",X"D9",X"13",X"D9",X"10",X"F5",X"23",X"FD",
		X"7E",X"02",X"BD",X"20",X"EB",X"C3",X"30",X"3F",X"BC",X"20",X"E5",X"FD",X"4E",X"04",X"FD",X"46",
		X"05",X"D9",X"7B",X"D9",X"BB",X"20",X"06",X"D9",X"7A",X"D9",X"BA",X"28",X"06",X"FD",X"4E",X"06",
		X"FD",X"46",X"07",X"C5",X"DD",X"E1",X"C3",X"E0",X"1F",X"C3",X"C0",X"1F",X"FD",X"19",X"FD",X"7E",
		X"00",X"FD",X"A6",X"01",X"FE",X"FF",X"C2",X"53",X"04",X"21",X"6C",X"84",X"01",X"28",X"00",X"CD",
		X"CC",X"00",X"CD",X"8B",X"05",X"3E",X"01",X"32",X"15",X"80",X"06",X"04",X"C3",X"40",X"1F",X"E6",
		X"10",X"C2",X"39",X"05",X"21",X"FF",X"FF",X"C3",X"40",X"3F",X"20",X"FB",X"10",X"EE",X"C9",X"F5",
		X"3E",X"FF",X"3D",X"FE",X"00",X"20",X"FB",X"F1",X"C9",X"21",X"6C",X"84",X"01",X"28",X"00",X"CD",
		X"CC",X"00",X"DD",X"21",X"48",X"C6",X"CD",X"D2",X"00",X"C3",X"50",X"1F",X"E6",X"10",X"C2",X"56",
		X"05",X"3E",X"00",X"32",X"15",X"80",X"3A",X"15",X"80",X"B7",X"C2",X"65",X"05",X"3A",X"00",X"B0",
		X"E6",X"10",X"C2",X"6B",X"05",X"CD",X"8B",X"05",X"C3",X"49",X"05",X"C9",X"FD",X"6E",X"04",X"FD",
		X"66",X"05",X"B7",X"FD",X"4E",X"06",X"FD",X"46",X"07",X"ED",X"52",X"CA",X"84",X"05",X"FD",X"4E",
		X"08",X"FD",X"46",X"09",X"C5",X"DD",X"E1",X"CD",X"D2",X"00",X"C9",X"DD",X"21",X"81",X"84",X"FD",
		X"21",X"00",X"B0",X"11",X"14",X"00",X"21",X"E4",X"C5",X"06",X"05",X"C5",X"D5",X"E5",X"DD",X"E5",
		X"11",X"6C",X"84",X"01",X"14",X"00",X"ED",X"B0",X"C3",X"F7",X"1F",X"B7",X"CA",X"B9",X"05",X"CD",
		X"CE",X"05",X"DD",X"21",X"6C",X"84",X"CD",X"D2",X"00",X"DD",X"E1",X"E1",X"D1",X"C1",X"78",X"FE",
		X"03",X"C2",X"C6",X"05",X"FD",X"23",X"FD",X"23",X"19",X"DD",X"23",X"10",X"CE",X"C9",X"C5",X"DD",
		X"E5",X"DD",X"21",X"6E",X"84",X"FD",X"E5",X"C1",X"79",X"FE",X"02",X"C2",X"E3",X"05",X"06",X"04",
		X"C3",X"E5",X"05",X"06",X"08",X"FD",X"7E",X"00",X"B7",X"1F",X"D2",X"F4",X"05",X"DD",X"36",X"00",
		X"31",X"C3",X"F8",X"05",X"C3",X"80",X"1F",X"00",X"DD",X"23",X"DD",X"23",X"10",X"EA",X"DD",X"E1",
		X"C1",X"C9",X"DD",X"7E",X"00",X"FD",X"BE",X"00",X"CA",X"16",X"06",X"FD",X"7E",X"00",X"DD",X"77",
		X"00",X"3E",X"01",X"C3",X"17",X"06",X"AF",X"C9",X"11",X"00",X"8C",X"21",X"00",X"D5",X"01",X"00",
		X"01",X"ED",X"B0",X"11",X"00",X"88",X"21",X"1A",X"0F",X"01",X"70",X"00",X"ED",X"B0",X"C9",X"C5",
		X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",X"DD",X"21",X"00",X"88",X"DD",X"7E",X"00",X"FE",X"FF",X"CA",
		X"A8",X"06",X"DD",X"CB",X"00",X"7E",X"C2",X"95",X"06",X"DD",X"7E",X"03",X"DD",X"BE",X"07",X"28",
		X"03",X"D2",X"9D",X"06",X"DD",X"36",X"07",X"00",X"DD",X"66",X"02",X"DD",X"6E",X"01",X"16",X"00",
		X"DD",X"5E",X"08",X"19",X"E5",X"23",X"23",X"0E",X"00",X"23",X"7E",X"FE",X"FF",X"28",X"05",X"DD",
		X"4E",X"08",X"0C",X"0C",X"DD",X"71",X"08",X"E1",X"FD",X"21",X"00",X"00",X"11",X"10",X"00",X"DD",
		X"7E",X"00",X"E6",X"7F",X"FE",X"00",X"28",X"05",X"FD",X"19",X"3D",X"18",X"F7",X"11",X"00",X"8C",
		X"FD",X"19",X"CD",X"B0",X"06",X"11",X"0A",X"00",X"DD",X"19",X"C3",X"3A",X"06",X"DD",X"34",X"07",
		X"11",X"0A",X"00",X"DD",X"19",X"C3",X"3A",X"06",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"C9",
		X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",X"7E",X"32",X"72",X"88",X"23",X"7E",X"32",X"73",X"88",
		X"DD",X"7E",X"05",X"87",X"11",X"00",X"00",X"5F",X"FD",X"19",X"FD",X"E5",X"DD",X"4E",X"06",X"0D",
		X"11",X"02",X"00",X"DD",X"7E",X"04",X"FE",X"01",X"28",X"03",X"11",X"FE",X"FF",X"21",X"74",X"88",
		X"79",X"FE",X"00",X"28",X"0F",X"FD",X"7E",X"00",X"77",X"23",X"FD",X"7E",X"01",X"77",X"23",X"FD",
		X"19",X"0D",X"18",X"EC",X"FD",X"E1",X"21",X"72",X"88",X"DD",X"4E",X"06",X"79",X"FE",X"00",X"28",
		X"0F",X"7E",X"FD",X"77",X"00",X"23",X"7E",X"FD",X"77",X"01",X"23",X"FD",X"19",X"0D",X"18",X"EC",
		X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"C9",X"3A",X"70",X"80",X"B7",X"C2",X"8E",X"02",X"C9",
		X"DD",X"21",X"00",X"90",X"FD",X"21",X"00",X"94",X"01",X"00",X"00",X"78",X"FE",X"10",X"28",X"3A",
		X"79",X"FE",X"10",X"20",X"0A",X"04",X"0E",X"00",X"11",X"20",X"00",X"DD",X"19",X"FD",X"19",X"DD",
		X"36",X"00",X"5C",X"DD",X"36",X"01",X"5D",X"DD",X"36",X"20",X"5E",X"DD",X"36",X"21",X"5F",X"FD",
		X"36",X"00",X"05",X"FD",X"36",X"01",X"05",X"FD",X"36",X"20",X"05",X"FD",X"36",X"21",X"05",X"DD",
		X"23",X"DD",X"23",X"FD",X"23",X"FD",X"23",X"0C",X"18",X"C1",X"06",X"00",X"21",X"FF",X"FF",X"C3",
		X"90",X"1F",X"CB",X"67",X"20",X"0C",X"2B",X"7C",X"B5",X"20",X"F4",X"04",X"78",X"FE",X"03",X"38",
		X"EB",X"C9",X"16",X"FF",X"15",X"7A",X"20",X"FC",X"C3",X"A0",X"1F",X"CB",X"67",X"28",X"F3",X"16",
		X"FF",X"15",X"7A",X"20",X"FC",X"C3",X"B0",X"1F",X"CB",X"67",X"20",X"F3",X"04",X"78",X"FE",X"03",
		X"38",X"E0",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"36",X"00",X"23",X"0B",X"79",X"B0",X"C2",X"50",X"08",X"C9",X"36",X"00",X"23",X"0B",X"79",X"B0",
		X"C2",X"5A",X"08",X"C9",X"D5",X"E5",X"2A",X"24",X"80",X"5D",X"54",X"19",X"19",X"E5",X"2A",X"22",
		X"80",X"5D",X"54",X"CB",X"23",X"CB",X"12",X"19",X"22",X"22",X"80",X"E1",X"ED",X"5A",X"22",X"24",
		X"80",X"E1",X"D1",X"C9",X"07",X"11",X"54",X"05",X"2E",X"05",X"54",X"05",X"FF",X"FF",X"09",X"11",
		X"45",X"05",X"2E",X"05",X"45",X"05",X"FF",X"FF",X"0B",X"11",X"48",X"05",X"2E",X"05",X"48",X"05",
		X"FF",X"FF",X"0D",X"11",X"4B",X"05",X"2E",X"05",X"4B",X"05",X"FF",X"FF",X"0F",X"11",X"41",X"05",
		X"2E",X"05",X"41",X"05",X"FF",X"FF",X"11",X"11",X"4E",X"05",X"2E",X"05",X"4E",X"05",X"FF",X"FF",
		X"13",X"11",X"4C",X"05",X"2E",X"05",X"4C",X"05",X"FF",X"FF",X"15",X"11",X"54",X"05",X"2E",X"05",
		X"54",X"05",X"FF",X"FF",X"17",X"11",X"44",X"05",X"2E",X"05",X"44",X"05",X"FF",X"FF",X"19",X"11",
		X"2E",X"05",X"2E",X"05",X"2E",X"05",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"10",X"00",
		X"00",X"00",X"03",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"05",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"05",X"00",X"21",X"00",X"B0",X"06",X"10",X"36",X"00",X"23",
		X"10",X"FB",X"21",X"84",X"08",X"11",X"32",X"81",X"01",X"64",X"00",X"ED",X"B0",X"11",X"00",X"81",
		X"06",X"0A",X"0E",X"04",X"CD",X"45",X"09",X"ED",X"A0",X"79",X"B7",X"20",X"FA",X"10",X"F3",X"CD",
		X"45",X"09",X"11",X"E2",X"80",X"01",X"04",X"00",X"ED",X"B0",X"21",X"28",X"81",X"06",X"0A",X"36",
		X"01",X"23",X"10",X"FB",X"C9",X"C5",X"D5",X"3A",X"14",X"80",X"E6",X"07",X"21",X"E8",X"08",X"01",
		X"04",X"00",X"CD",X"F6",X"00",X"D1",X"C1",X"C9",X"DD",X"21",X"78",X"98",X"FD",X"21",X"20",X"98",
		X"21",X"00",X"85",X"06",X"0C",X"0E",X"03",X"78",X"FE",X"00",X"28",X"11",X"23",X"7E",X"2B",X"CB",
		X"6F",X"20",X"05",X"CD",X"82",X"09",X"18",X"EF",X"CD",X"96",X"09",X"18",X"EA",X"79",X"32",X"00",
		X"9A",X"C9",X"05",X"C5",X"D5",X"DD",X"E5",X"D1",X"01",X"08",X"00",X"ED",X"B0",X"11",X"F8",X"FF",
		X"B7",X"DD",X"19",X"D1",X"C1",X"C9",X"0C",X"05",X"C5",X"D5",X"FD",X"E5",X"D1",X"01",X"08",X"00",
		X"ED",X"B0",X"11",X"08",X"00",X"B7",X"FD",X"19",X"D1",X"C1",X"C9",X"21",X"40",X"8C",X"11",X"40",
		X"9C",X"01",X"10",X"00",X"ED",X"B0",X"21",X"A0",X"8C",X"11",X"A0",X"9C",X"01",X"60",X"00",X"ED",
		X"B0",X"3A",X"8C",X"80",X"B7",X"C8",X"FE",X"02",X"28",X"12",X"3E",X"00",X"32",X"8C",X"80",X"21",
		X"00",X"8C",X"11",X"00",X"9C",X"01",X"A0",X"00",X"ED",X"B0",X"18",X"05",X"3E",X"00",X"32",X"8C",
		X"80",X"C9",X"2A",X"6E",X"80",X"7D",X"B4",X"28",X"04",X"2B",X"22",X"6E",X"80",X"C9",X"F5",X"ED",
		X"43",X"6E",X"80",X"ED",X"4B",X"6E",X"80",X"79",X"B0",X"20",X"F8",X"F1",X"C9",X"F5",X"C5",X"D5",
		X"E5",X"DD",X"E5",X"FD",X"E5",X"CD",X"8A",X"0B",X"C5",X"E1",X"4E",X"23",X"46",X"23",X"C5",X"DD",
		X"E1",X"CD",X"21",X"0A",X"3D",X"C2",X"0A",X"0A",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"F1",
		X"C9",X"F5",X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",X"CD",X"82",X"0A",X"E5",X"DD",X"7E",X"05",
		X"3D",X"CB",X"2F",X"16",X"00",X"5F",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"19",X"E5",X"D1",X"E1",
		X"0E",X"00",X"DD",X"46",X"05",X"78",X"3D",X"20",X"02",X"0E",X"0F",X"CD",X"59",X"0A",X"10",X"F5",
		X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"F1",X"C9",X"1A",X"CB",X"40",X"C2",X"67",X"0A",X"E6",
		X"F0",X"0F",X"0F",X"0F",X"0F",X"18",X"02",X"E6",X"0F",X"CD",X"07",X"0B",X"77",X"D5",X"11",X"00",
		X"04",X"19",X"DD",X"7E",X"04",X"77",X"11",X"E0",X"FB",X"19",X"D1",X"CB",X"40",X"CA",X"81",X"0A",
		X"1B",X"C9",X"F5",X"DD",X"46",X"01",X"21",X"00",X"94",X"11",X"E0",X"FF",X"04",X"19",X"10",X"FD",
		X"06",X"00",X"DD",X"4E",X"00",X"09",X"F1",X"C9",X"F5",X"C5",X"D5",X"FD",X"E5",X"CB",X"38",X"CB",
		X"38",X"CB",X"38",X"CB",X"39",X"CB",X"39",X"CB",X"39",X"FD",X"21",X"C7",X"0A",X"16",X"00",X"CB",
		X"20",X"58",X"FD",X"19",X"FD",X"5E",X"00",X"FD",X"56",X"01",X"21",X"00",X"94",X"19",X"06",X"00",
		X"09",X"FD",X"E1",X"D1",X"C1",X"F1",X"C9",X"E0",X"FF",X"C0",X"FF",X"A0",X"FF",X"80",X"FF",X"60",
		X"FF",X"40",X"FF",X"20",X"FF",X"00",X"FF",X"E0",X"FE",X"C0",X"FE",X"A0",X"FE",X"80",X"FE",X"60",
		X"FE",X"40",X"FE",X"20",X"FE",X"00",X"FE",X"E0",X"FD",X"C0",X"FD",X"A0",X"FD",X"80",X"FD",X"60",
		X"FD",X"40",X"FD",X"20",X"FD",X"00",X"FD",X"E0",X"FC",X"C0",X"FC",X"A0",X"FC",X"80",X"FC",X"60",
		X"FC",X"40",X"FC",X"20",X"FC",X"00",X"FC",X"B7",X"20",X"07",X"B9",X"20",X"04",X"3E",X"00",X"18",
		X"0B",X"0E",X"0F",X"C6",X"30",X"FE",X"3A",X"DA",X"1C",X"0B",X"C6",X"07",X"C9",X"F5",X"C5",X"D5",
		X"E5",X"DD",X"E5",X"FD",X"E5",X"CD",X"8A",X"0B",X"C5",X"E1",X"4E",X"23",X"46",X"23",X"C5",X"DD",
		X"E1",X"CD",X"41",X"0B",X"3D",X"C2",X"2A",X"0B",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"F1",
		X"C9",X"F5",X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",X"CD",X"82",X"0A",X"DD",X"23",X"DD",X"23",
		X"DD",X"5E",X"00",X"DD",X"56",X"01",X"3E",X"FF",X"BA",X"CA",X"65",X"0B",X"CD",X"D3",X"5F",X"CD",
		X"9F",X"0B",X"C3",X"4C",X"0B",X"BB",X"CA",X"81",X"0B",X"7B",X"DD",X"23",X"DD",X"23",X"DD",X"5E",
		X"00",X"DD",X"56",X"01",X"CD",X"D3",X"5F",X"CD",X"9F",X"0B",X"3D",X"C2",X"77",X"0B",X"C3",X"4C",
		X"0B",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"F1",X"C9",X"21",X"0E",X"00",X"39",X"5E",X"23",
		X"56",X"E5",X"EB",X"4E",X"23",X"46",X"23",X"7E",X"23",X"EB",X"E1",X"72",X"2B",X"73",X"C9",X"73",
		X"C5",X"01",X"00",X"04",X"09",X"72",X"01",X"E0",X"FB",X"09",X"C1",X"C9",X"CD",X"1E",X"60",X"C9",
		X"87",X"16",X"00",X"5F",X"19",X"5E",X"23",X"56",X"EB",X"E9",X"C5",X"D5",X"E5",X"DD",X"E5",X"DD",
		X"21",X"00",X"94",X"21",X"00",X"90",X"5F",X"16",X"00",X"19",X"DD",X"19",X"11",X"20",X"00",X"06",
		X"20",X"36",X"00",X"DD",X"36",X"00",X"0A",X"DD",X"19",X"19",X"05",X"C2",X"D1",X"0B",X"DD",X"E1",
		X"E1",X"D1",X"C1",X"C9",X"F5",X"C5",X"78",X"CD",X"BA",X"0B",X"3C",X"0D",X"C2",X"E7",X"0B",X"C1",
		X"F1",X"C9",X"DD",X"21",X"12",X"C8",X"CD",X"D2",X"00",X"DD",X"21",X"22",X"C8",X"CD",X"D5",X"00",
		X"C9",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",X"11",X"8A",X"0F",X"29",X"19",X"5E",X"23",X"56",X"26",
		X"00",X"6F",X"19",X"7E",X"DD",X"77",X"02",X"DD",X"36",X"03",X"05",X"3A",X"AC",X"81",X"16",X"00",
		X"5F",X"21",X"A8",X"0F",X"19",X"7E",X"FD",X"77",X"04",X"FD",X"36",X"05",X"05",X"DD",X"7E",X"04",
		X"C6",X"10",X"FD",X"77",X"06",X"DD",X"7E",X"05",X"FD",X"77",X"07",X"FD",X"E1",X"DD",X"E1",X"E1",
		X"D1",X"C9",X"B7",X"CA",X"4B",X"0C",X"09",X"3D",X"C2",X"46",X"0C",X"C9",X"B7",X"CA",X"55",X"0C",
		X"09",X"3D",X"C2",X"50",X"0C",X"5E",X"23",X"56",X"EB",X"C9",X"3A",X"00",X"B0",X"E6",X"20",X"CA",
		X"92",X"0C",X"3A",X"02",X"B0",X"E6",X"04",X"C2",X"62",X"0C",X"3A",X"00",X"B0",X"E6",X"20",X"CA",
		X"92",X"0C",X"3A",X"02",X"B0",X"E6",X"04",X"C2",X"7D",X"0C",X"C3",X"6A",X"0C",X"06",X"FF",X"3E",
		X"1C",X"3D",X"C2",X"81",X"0C",X"10",X"F8",X"3A",X"02",X"B0",X"E6",X"04",X"C2",X"92",X"0C",X"C3",
		X"6A",X"0C",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"FF",X"02",X"FF",X"04",X"FF",X"06",X"FF",X"08",X"FF",X"0A",X"FF",X"0C",X"FF",X"0F",
		X"CC",X"0F",X"AA",X"0F",X"88",X"0F",X"66",X"0F",X"44",X"0F",X"22",X"0F",X"00",X"0F",X"02",X"0F",
		X"04",X"0F",X"06",X"0F",X"08",X"0F",X"0A",X"0F",X"0C",X"0F",X"0F",X"0F",X"0F",X"0C",X"0F",X"0A",
		X"0F",X"08",X"0F",X"06",X"0F",X"04",X"0F",X"02",X"0F",X"00",X"2F",X"00",X"4F",X"00",X"6F",X"00",
		X"8F",X"00",X"AF",X"00",X"CF",X"00",X"FF",X"FF",X"0F",X"00",X"2F",X"00",X"4F",X"00",X"6F",X"00",
		X"8F",X"00",X"AF",X"00",X"CF",X"00",X"FF",X"00",X"FC",X"00",X"FA",X"00",X"F8",X"00",X"F6",X"00",
		X"F4",X"00",X"F2",X"00",X"F0",X"00",X"F0",X"02",X"F0",X"04",X"F0",X"06",X"F0",X"08",X"F0",X"0A",
		X"F0",X"0C",X"F0",X"0F",X"C0",X"0F",X"A0",X"0F",X"80",X"0F",X"60",X"0F",X"40",X"0F",X"20",X"0F",
		X"00",X"0F",X"02",X"0F",X"04",X"0F",X"06",X"0F",X"08",X"0F",X"0A",X"0F",X"0C",X"0F",X"0F",X"0F",
		X"0F",X"0C",X"0F",X"0A",X"0F",X"08",X"0F",X"06",X"0F",X"04",X"0F",X"02",X"FF",X"FF",X"00",X"0F",
		X"22",X"0F",X"44",X"0F",X"66",X"0F",X"88",X"0F",X"AA",X"0F",X"CC",X"0F",X"EE",X"0F",X"FF",X"FF",
		X"0F",X"00",X"2F",X"02",X"4F",X"04",X"6F",X"06",X"8F",X"08",X"AF",X"0A",X"CF",X"0C",X"EF",X"0E",
		X"FF",X"FF",X"0F",X"0F",X"2F",X"0F",X"4F",X"0F",X"6F",X"0F",X"8F",X"0F",X"AF",X"0F",X"CF",X"0F",
		X"EF",X"0F",X"FF",X"FF",X"F0",X"00",X"F2",X"02",X"F4",X"04",X"F6",X"06",X"F8",X"08",X"FA",X"0A",
		X"FC",X"0C",X"FE",X"0E",X"FF",X"FF",X"F0",X"0F",X"F2",X"0F",X"F4",X"0F",X"F6",X"0F",X"F8",X"0F",
		X"FA",X"0F",X"FC",X"0F",X"FE",X"0F",X"FF",X"FF",X"FF",X"00",X"FF",X"02",X"FF",X"04",X"FF",X"06",
		X"FF",X"08",X"FF",X"0A",X"FF",X"0C",X"FF",X"0E",X"FF",X"FF",X"FF",X"0F",X"EE",X"0E",X"DD",X"0D",
		X"CC",X"0C",X"BB",X"0B",X"AA",X"0A",X"99",X"09",X"88",X"08",X"FF",X"FF",X"0F",X"00",X"00",X"00",
		X"9F",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"0F",X"00",X"00",X"0F",X"00",X"00",X"00",
		X"9F",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"0F",X"00",X"00",X"0F",X"00",X"00",X"00",
		X"9F",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"9F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"08",X"00",X"FF",X"FF",X"0F",X"0F",X"00",X"00",X"0F",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0C",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"0D",X"00",X"0B",X"00",X"09",X"00",X"07",X"00",X"05",X"00",X"03",X"00",X"01",X"00",
		X"00",X"00",X"00",X"FF",X"CC",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"0F",X"FF",X"FF",X"00",X"0F",X"22",X"0F",X"44",X"0F",X"66",X"0F",X"88",X"0F",X"AA",X"0F",
		X"CC",X"0F",X"FF",X"0F",X"FF",X"FF",X"FF",X"00",X"FF",X"02",X"FF",X"04",X"FF",X"06",X"FF",X"08",
		X"FF",X"0A",X"FF",X"0C",X"FF",X"0F",X"FF",X"FF",X"0F",X"00",X"2F",X"02",X"4F",X"04",X"6F",X"06",
		X"8F",X"08",X"AF",X"0A",X"CF",X"0C",X"FF",X"0F",X"FF",X"FF",X"99",X"00",X"AA",X"00",X"BB",X"00",
		X"CC",X"00",X"DD",X"00",X"EE",X"00",X"FF",X"00",X"FF",X"FF",X"84",X"D0",X"0F",X"03",X"01",X"05",
		X"03",X"02",X"00",X"00",X"8A",X"00",X"00",X"04",X"01",X"01",X"06",X"00",X"00",X"00",X"8B",X"0A",
		X"0F",X"01",X"07",X"07",X"07",X"01",X"00",X"00",X"0C",X"C4",X"0E",X"02",X"01",X"07",X"01",X"00",
		X"00",X"00",X"0D",X"1C",X"0E",X"01",X"01",X"01",X"01",X"02",X"00",X"00",X"0D",X"46",X"0E",X"01",
		X"01",X"02",X"01",X"02",X"00",X"00",X"0D",X"70",X"0E",X"01",X"01",X"03",X"01",X"02",X"00",X"00",
		X"0D",X"9A",X"0E",X"04",X"01",X"04",X"01",X"02",X"00",X"00",X"0E",X"48",X"0D",X"02",X"07",X"07",
		X"07",X"04",X"00",X"00",X"0F",X"00",X"0D",X"02",X"07",X"07",X"07",X"02",X"00",X"00",X"04",X"BB",
		X"0F",X"03",X"01",X"01",X"01",X"03",X"00",X"00",X"FF",X"FF",X"92",X"0F",X"9A",X"0F",X"9D",X"0F",
		X"9F",X"0F",X"00",X"70",X"71",X"72",X"74",X"76",X"78",X"7A",X"77",X"79",X"7B",X"71",X"73",X"70",
		X"71",X"72",X"74",X"76",X"78",X"7A",X"7A",X"7A",X"00",X"7C",X"7D",X"7E",X"7F",X"FF",X"00",X"FB",
		X"00",X"F8",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"00",X"0C",X"00",X"08",
		X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"08",X"00",X"0C",X"00",X"FF",X"FF",X"FF",X"FF",X"00",
		X"B0",X"0F",X"80",X"0F",X"50",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"3A",X"13",X"80",X"CB",X"77",X"C2",X"EE",X"0F",X"3A",X"01",X"B0",X"C3",X"A2",X"03",X"3A",X"00",
		X"B0",X"C3",X"A2",X"03",X"00",X"00",X"00",X"00",X"3A",X"03",X"B0",X"3A",X"00",X"B0",X"C9",X"00",
		X"3A",X"8E",X"80",X"FE",X"00",X"28",X"0B",X"3A",X"28",X"80",X"CB",X"97",X"32",X"28",X"80",X"C3",
		X"C3",X"00",X"DD",X"21",X"28",X"80",X"DD",X"CB",X"00",X"56",X"C2",X"DD",X"12",X"DD",X"CB",X"00",
		X"7E",X"28",X"42",X"DD",X"36",X"02",X"00",X"2A",X"36",X"80",X"2B",X"22",X"36",X"80",X"7C",X"B5",
		X"20",X"14",X"CD",X"F9",X"2F",X"CD",X"E6",X"2F",X"DD",X"CB",X"00",X"BE",X"DD",X"CB",X"00",X"B6",
		X"DD",X"36",X"02",X"00",X"18",X"1F",X"7C",X"B7",X"20",X"1B",X"7D",X"FE",X"39",X"30",X"16",X"E6",
		X"03",X"FE",X"00",X"20",X"10",X"DD",X"CB",X"00",X"76",X"28",X"06",X"DD",X"CB",X"00",X"B6",X"18",
		X"04",X"DD",X"CB",X"00",X"F6",X"DD",X"7E",X"19",X"DD",X"34",X"23",X"CB",X"5F",X"20",X"04",X"DD",
		X"36",X"23",X"00",X"E6",X"0A",X"28",X"0A",X"DD",X"7E",X"0B",X"FE",X"FF",X"28",X"03",X"C3",X"72",
		X"12",X"3A",X"3F",X"80",X"FE",X"00",X"28",X"17",X"3A",X"20",X"80",X"FE",X"03",X"C2",X"CE",X"12",
		X"DD",X"36",X"17",X"00",X"DD",X"36",X"0B",X"00",X"DD",X"36",X"1C",X"00",X"C3",X"72",X"12",X"DD",
		X"CB",X"00",X"4E",X"C2",X"D2",X"10",X"CD",X"DD",X"1A",X"7C",X"B5",X"20",X"1F",X"ED",X"5B",X"40",
		X"80",X"7A",X"B3",X"28",X"17",X"CB",X"5A",X"28",X"05",X"3E",X"11",X"CD",X"FD",X"1B",X"01",X"10",
		X"00",X"CD",X"E4",X"00",X"3A",X"53",X"84",X"F6",X"C0",X"32",X"53",X"84",X"DD",X"74",X"18",X"DD",
		X"75",X"19",X"CD",X"70",X"18",X"CD",X"B7",X"17",X"DD",X"7E",X"12",X"FE",X"FF",X"C2",X"25",X"12",
		X"2A",X"42",X"80",X"7C",X"B5",X"20",X"0A",X"2A",X"31",X"80",X"7C",X"B5",X"20",X"03",X"C3",X"38",
		X"11",X"DD",X"CB",X"00",X"46",X"C2",X"52",X"11",X"3A",X"20",X"80",X"FE",X"03",X"C2",X"1D",X"11",
		X"CD",X"73",X"17",X"3E",X"12",X"CD",X"FD",X"1B",X"DD",X"36",X"0B",X"00",X"DD",X"36",X"1C",X"00",
		X"DD",X"CB",X"19",X"5E",X"28",X"07",X"DD",X"CB",X"00",X"C6",X"C3",X"72",X"12",X"3A",X"41",X"80",
		X"CB",X"5F",X"28",X"11",X"DD",X"CB",X"00",X"46",X"20",X"0B",X"CD",X"73",X"17",X"DD",X"36",X"17",
		X"08",X"DD",X"CB",X"00",X"C6",X"C3",X"A7",X"11",X"3A",X"20",X"80",X"FE",X"03",X"20",X"10",X"3E",
		X"12",X"CD",X"FD",X"1B",X"DD",X"36",X"0B",X"00",X"DD",X"36",X"1C",X"00",X"C3",X"72",X"12",X"C3",
		X"A7",X"11",X"3A",X"20",X"80",X"FE",X"03",X"C2",X"77",X"11",X"CD",X"73",X"17",X"3E",X"12",X"CD",
		X"FD",X"1B",X"DD",X"36",X"0B",X"00",X"DD",X"36",X"1C",X"00",X"DD",X"CB",X"19",X"4E",X"28",X"07",
		X"DD",X"CB",X"00",X"86",X"C3",X"72",X"12",X"3A",X"41",X"80",X"CB",X"4F",X"28",X"11",X"DD",X"CB",
		X"00",X"46",X"28",X"0B",X"CD",X"73",X"17",X"DD",X"36",X"17",X"00",X"DD",X"CB",X"00",X"86",X"2A",
		X"42",X"80",X"CB",X"7C",X"20",X"04",X"7C",X"B5",X"20",X"0A",X"21",X"00",X"00",X"22",X"42",X"80",
		X"DD",X"CB",X"00",X"86",X"C3",X"A7",X"11",X"3A",X"41",X"80",X"CB",X"5F",X"28",X"12",X"2A",X"42",
		X"80",X"7C",X"B5",X"20",X"0B",X"21",X"00",X"00",X"22",X"31",X"80",X"22",X"38",X"80",X"18",X"1E",
		X"CD",X"E3",X"18",X"DD",X"CB",X"00",X"46",X"20",X"0C",X"2A",X"5A",X"80",X"11",X"0A",X"00",X"19",
		X"22",X"31",X"80",X"18",X"09",X"2A",X"5A",X"80",X"CD",X"D9",X"18",X"22",X"31",X"80",X"CD",X"9A",
		X"18",X"2A",X"42",X"80",X"ED",X"5B",X"31",X"80",X"3A",X"1C",X"80",X"FE",X"00",X"20",X"09",X"3A",
		X"1E",X"80",X"FE",X"00",X"20",X"09",X"18",X"0C",X"B7",X"CB",X"2A",X"CB",X"1B",X"18",X"05",X"B7",
		X"CB",X"23",X"CB",X"12",X"19",X"CB",X"7C",X"20",X"09",X"7C",X"B5",X"28",X"05",X"22",X"42",X"80",
		X"18",X"10",X"DD",X"CB",X"00",X"46",X"28",X"0A",X"21",X"00",X"00",X"22",X"42",X"80",X"DD",X"CB",
		X"00",X"86",X"C3",X"72",X"12",X"DD",X"CB",X"00",X"46",X"C2",X"4F",X"12",X"3A",X"20",X"80",X"FE",
		X"03",X"20",X"06",X"CD",X"73",X"17",X"CD",X"0D",X"17",X"3A",X"20",X"80",X"FE",X"FF",X"20",X"03",
		X"CD",X"33",X"17",X"3A",X"20",X"80",X"B7",X"20",X"03",X"CD",X"53",X"17",X"C3",X"1D",X"11",X"3A",
		X"20",X"80",X"FE",X"03",X"20",X"06",X"CD",X"73",X"17",X"CD",X"0D",X"17",X"3A",X"20",X"80",X"FE",
		X"FF",X"20",X"03",X"CD",X"33",X"17",X"3A",X"20",X"80",X"B7",X"20",X"03",X"CD",X"53",X"17",X"C3",
		X"77",X"11",X"DD",X"CB",X"00",X"9E",X"CD",X"8E",X"15",X"DD",X"CB",X"00",X"5E",X"20",X"03",X"CD",
		X"B4",X"14",X"CD",X"51",X"19",X"DD",X"CB",X"00",X"8E",X"3A",X"02",X"85",X"DD",X"BE",X"03",X"20",
		X"0C",X"3A",X"03",X"85",X"DD",X"BE",X"04",X"20",X"04",X"DD",X"CB",X"00",X"CE",X"DD",X"CB",X"00",
		X"7E",X"28",X"04",X"DD",X"36",X"02",X"0E",X"CD",X"F4",X"16",X"3A",X"3A",X"80",X"FE",X"FF",X"28",
		X"1A",X"FE",X"00",X"20",X"0F",X"3A",X"35",X"80",X"3C",X"32",X"35",X"80",X"CD",X"B7",X"17",X"CD",
		X"FC",X"17",X"18",X"07",X"3A",X"3A",X"80",X"3D",X"32",X"3A",X"80",X"C3",X"C3",X"00",X"3E",X"19",
		X"32",X"00",X"85",X"3A",X"3F",X"80",X"3D",X"32",X"3F",X"80",X"C3",X"C3",X"00",X"3A",X"95",X"80",
		X"FE",X"FF",X"28",X"06",X"CD",X"70",X"13",X"C3",X"6D",X"13",X"DD",X"21",X"5E",X"80",X"FD",X"21",
		X"00",X"85",X"3A",X"5F",X"80",X"FE",X"FF",X"28",X"2C",X"3E",X"01",X"CD",X"FC",X"00",X"3E",X"14",
		X"CD",X"FC",X"00",X"DD",X"36",X"00",X"00",X"DD",X"36",X"01",X"FF",X"FD",X"36",X"00",X"A4",X"FD",
		X"36",X"01",X"20",X"FD",X"7E",X"02",X"D6",X"08",X"FD",X"77",X"02",X"FD",X"7E",X"03",X"D6",X"08",
		X"FD",X"77",X"03",X"18",X"48",X"DD",X"7E",X"00",X"FE",X"40",X"D2",X"41",X"13",X"DD",X"34",X"00",
		X"DD",X"7E",X"00",X"FE",X"40",X"D2",X"41",X"13",X"E6",X"0F",X"20",X"31",X"FD",X"34",X"00",X"18",
		X"2C",X"21",X"00",X"00",X"22",X"00",X"85",X"3A",X"88",X"80",X"FE",X"00",X"20",X"1F",X"3A",X"8E",
		X"80",X"FE",X"00",X"20",X"18",X"3E",X"00",X"32",X"95",X"80",X"3A",X"70",X"80",X"FE",X"00",X"20",
		X"07",X"3E",X"01",X"32",X"78",X"80",X"18",X"05",X"3E",X"01",X"32",X"77",X"80",X"C3",X"C3",X"00",
		X"DD",X"21",X"95",X"80",X"DD",X"7E",X"00",X"E6",X"0F",X"FE",X"0F",X"28",X"0A",X"FE",X"07",X"28",
		X"06",X"CD",X"2D",X"14",X"C3",X"2C",X"14",X"21",X"00",X"00",X"22",X"31",X"80",X"CD",X"DD",X"1A",
		X"CB",X"5D",X"28",X"0C",X"DD",X"36",X"00",X"FF",X"3E",X"A7",X"CD",X"FC",X"00",X"C3",X"2C",X"14",
		X"DD",X"7E",X"00",X"FE",X"0F",X"28",X"27",X"DD",X"36",X"00",X"0F",X"2A",X"AA",X"14",X"DD",X"75",
		X"01",X"DD",X"74",X"02",X"DD",X"36",X"03",X"00",X"3A",X"03",X"85",X"DD",X"77",X"04",X"DD",X"36",
		X"05",X"00",X"DD",X"36",X"06",X"00",X"DD",X"36",X"07",X"00",X"DD",X"36",X"08",X"00",X"2A",X"9A",
		X"80",X"11",X"0A",X"00",X"19",X"22",X"9A",X"80",X"ED",X"5B",X"98",X"80",X"19",X"22",X"98",X"80",
		X"DD",X"34",X"07",X"DD",X"7E",X"07",X"FE",X"05",X"38",X"30",X"DD",X"36",X"07",X"00",X"FD",X"21",
		X"AA",X"14",X"16",X"00",X"DD",X"5E",X"08",X"FD",X"19",X"FD",X"7E",X"00",X"FE",X"FF",X"20",X"08",
		X"FD",X"21",X"AA",X"14",X"DD",X"36",X"08",X"00",X"DD",X"34",X"08",X"DD",X"34",X"08",X"FD",X"7E",
		X"00",X"DD",X"77",X"01",X"FD",X"7E",X"01",X"DD",X"77",X"02",X"3A",X"96",X"80",X"32",X"00",X"85",
		X"3A",X"97",X"80",X"32",X"01",X"85",X"3A",X"99",X"80",X"32",X"03",X"85",X"C9",X"DD",X"7E",X"00",
		X"FE",X"03",X"28",X"1F",X"3E",X"01",X"32",X"8D",X"80",X"DD",X"36",X"00",X"03",X"DD",X"36",X"07",
		X"00",X"DD",X"36",X"08",X"00",X"DD",X"36",X"09",X"00",X"3E",X"01",X"CD",X"FC",X"00",X"3E",X"27",
		X"CD",X"FC",X"00",X"DD",X"7E",X"07",X"FE",X"3C",X"38",X"07",X"DD",X"36",X"00",X"07",X"C3",X"9F",
		X"14",X"DD",X"7E",X"09",X"FE",X"03",X"38",X"2B",X"DD",X"36",X"09",X"00",X"FD",X"21",X"A0",X"14",
		X"16",X"00",X"DD",X"5E",X"08",X"B7",X"FD",X"19",X"FD",X"7E",X"00",X"FE",X"FF",X"20",X"08",X"FD",
		X"21",X"A0",X"14",X"DD",X"36",X"08",X"00",X"FD",X"7E",X"00",X"32",X"00",X"85",X"FD",X"7E",X"01",
		X"32",X"01",X"85",X"DD",X"34",X"07",X"DD",X"34",X"08",X"DD",X"34",X"08",X"DD",X"34",X"09",X"C9",
		X"28",X"C0",X"28",X"80",X"28",X"00",X"28",X"40",X"FF",X"FF",X"48",X"00",X"49",X"00",X"4A",X"00",
		X"4B",X"00",X"FF",X"FF",X"E5",X"D5",X"2A",X"2F",X"80",X"ED",X"5B",X"31",X"80",X"7A",X"B3",X"20",
		X"48",X"3A",X"41",X"80",X"CB",X"5F",X"28",X"41",X"7C",X"B5",X"20",X"11",X"3A",X"29",X"80",X"FE",
		X"1B",X"38",X"06",X"FE",X"23",X"30",X"02",X"18",X"5A",X"3E",X"18",X"18",X"56",X"CB",X"7C",X"20",
		X"14",X"DD",X"34",X"22",X"3A",X"4A",X"80",X"FE",X"04",X"DA",X"4B",X"15",X"DD",X"36",X"22",X"00",
		X"CD",X"4E",X"15",X"18",X"4B",X"DD",X"34",X"22",X"3A",X"4A",X"80",X"FE",X"04",X"DA",X"4B",X"15",
		X"DD",X"36",X"22",X"00",X"CD",X"6E",X"15",X"18",X"37",X"CB",X"7A",X"28",X"14",X"7C",X"B5",X"20",
		X"04",X"3E",X"23",X"18",X"1E",X"CB",X"7C",X"20",X"04",X"3E",X"25",X"18",X"16",X"3E",X"27",X"18",
		X"12",X"7C",X"B5",X"20",X"04",X"3E",X"24",X"18",X"0A",X"CB",X"7C",X"20",X"04",X"3E",X"26",X"18",
		X"02",X"3E",X"28",X"32",X"29",X"80",X"32",X"00",X"85",X"3E",X"93",X"CD",X"FD",X"1B",X"18",X"0B",
		X"32",X"29",X"80",X"32",X"00",X"85",X"3E",X"13",X"CD",X"FD",X"1B",X"D1",X"E1",X"C9",X"3A",X"29",
		X"80",X"FE",X"1B",X"F2",X"5A",X"15",X"3E",X"1B",X"18",X"13",X"FE",X"1E",X"28",X"06",X"38",X"04",
		X"3E",X"1B",X"18",X"09",X"3C",X"FE",X"1E",X"28",X"04",X"38",X"02",X"3E",X"1B",X"C9",X"3A",X"29",
		X"80",X"FE",X"1F",X"F2",X"7A",X"15",X"3E",X"1F",X"18",X"13",X"FE",X"22",X"28",X"06",X"38",X"04",
		X"3E",X"1F",X"18",X"09",X"3C",X"FE",X"22",X"28",X"04",X"38",X"02",X"3E",X"1F",X"C9",X"C5",X"D5",
		X"E5",X"DD",X"E5",X"DD",X"21",X"28",X"80",X"DD",X"7E",X"0B",X"FE",X"FF",X"CA",X"EE",X"16",X"DD",
		X"7E",X"1C",X"FE",X"02",X"CA",X"78",X"16",X"FE",X"01",X"CA",X"BC",X"15",X"DD",X"36",X"1D",X"28",
		X"DD",X"36",X"1E",X"00",X"DD",X"36",X"1F",X"00",X"DD",X"36",X"1C",X"01",X"3A",X"4B",X"80",X"FE",
		X"01",X"30",X"2A",X"3A",X"18",X"80",X"FE",X"00",X"20",X"07",X"3A",X"1A",X"80",X"FE",X"00",X"28",
		X"1C",X"DD",X"36",X"1D",X"00",X"DD",X"36",X"1E",X"00",X"DD",X"36",X"1F",X"00",X"DD",X"36",X"1C",
		X"02",X"21",X"00",X"00",X"22",X"42",X"80",X"22",X"31",X"80",X"C3",X"EE",X"16",X"DD",X"CB",X"00",
		X"DE",X"DD",X"7E",X"0B",X"FE",X"10",X"CA",X"3A",X"16",X"DA",X"3A",X"16",X"DD",X"36",X"1D",X"00",
		X"DD",X"36",X"1E",X"28",X"FE",X"20",X"CA",X"53",X"16",X"DA",X"53",X"16",X"DD",X"36",X"1E",X"04",
		X"DD",X"36",X"1C",X"02",X"DD",X"7E",X"19",X"E6",X"0A",X"28",X"0C",X"21",X"00",X"00",X"22",X"42",
		X"80",X"22",X"31",X"80",X"C3",X"6C",X"16",X"DD",X"7E",X"19",X"FE",X"00",X"28",X"06",X"CD",X"98",
		X"17",X"C3",X"6C",X"16",X"CD",X"73",X"17",X"C3",X"6C",X"16",X"DD",X"36",X"1D",X"00",X"DD",X"36",
		X"1E",X"04",X"DD",X"36",X"1F",X"02",X"01",X"FF",X"7F",X"CD",X"7A",X"17",X"DD",X"36",X"1C",X"02",
		X"C3",X"6C",X"16",X"3A",X"20",X"80",X"B7",X"C2",X"6C",X"16",X"DD",X"36",X"1E",X"04",X"DD",X"36",
		X"1F",X"02",X"01",X"00",X"1A",X"CD",X"7A",X"17",X"DD",X"36",X"1C",X"02",X"DD",X"7E",X"0B",X"FE",
		X"50",X"D2",X"78",X"16",X"3C",X"DD",X"77",X"0B",X"DD",X"7E",X"1D",X"FE",X"00",X"CA",X"8F",X"16",
		X"DD",X"36",X"0C",X"01",X"DD",X"36",X"0D",X"00",X"3D",X"DD",X"77",X"1D",X"C3",X"C9",X"16",X"DD",
		X"7E",X"1E",X"FE",X"00",X"CA",X"A6",X"16",X"DD",X"36",X"0C",X"01",X"DD",X"36",X"0D",X"01",X"3D",
		X"DD",X"77",X"1E",X"C3",X"C9",X"16",X"DD",X"7E",X"1F",X"FE",X"00",X"CA",X"BD",X"16",X"DD",X"36",
		X"0C",X"01",X"DD",X"36",X"0D",X"02",X"3D",X"DD",X"77",X"1F",X"C3",X"C9",X"16",X"DD",X"36",X"0C",
		X"00",X"DD",X"36",X"0D",X"00",X"DD",X"36",X"0B",X"FF",X"CD",X"B7",X"17",X"CD",X"FC",X"17",X"3A",
		X"20",X"80",X"FE",X"03",X"C2",X"EE",X"16",X"3E",X"12",X"CD",X"FD",X"1B",X"DD",X"36",X"0B",X"00",
		X"DD",X"36",X"1C",X"00",X"DD",X"7E",X"19",X"E6",X"0A",X"28",X"03",X"CD",X"73",X"17",X"DD",X"E1",
		X"E1",X"D1",X"C1",X"C9",X"3A",X"29",X"80",X"32",X"00",X"85",X"3A",X"2A",X"80",X"32",X"01",X"85",
		X"3A",X"2B",X"80",X"32",X"02",X"85",X"3A",X"2C",X"80",X"32",X"03",X"85",X"C9",X"3A",X"3B",X"80",
		X"CB",X"7F",X"28",X"0E",X"3A",X"3C",X"80",X"32",X"34",X"80",X"3A",X"3D",X"80",X"32",X"35",X"80",
		X"18",X"0A",X"CB",X"57",X"28",X"0C",X"3A",X"3E",X"80",X"32",X"35",X"80",X"CD",X"B7",X"17",X"CD",
		X"FC",X"17",X"C9",X"3A",X"3B",X"80",X"CB",X"77",X"28",X"08",X"3A",X"3D",X"80",X"32",X"34",X"80",
		X"18",X"0A",X"CB",X"4F",X"28",X"0C",X"3A",X"3D",X"80",X"32",X"35",X"80",X"CD",X"B7",X"17",X"CD",
		X"FC",X"17",X"C9",X"3A",X"3B",X"80",X"CB",X"6F",X"28",X"08",X"3A",X"3C",X"80",X"32",X"34",X"80",
		X"18",X"0A",X"CB",X"47",X"28",X"0C",X"3A",X"3C",X"80",X"32",X"35",X"80",X"CD",X"B7",X"17",X"CD",
		X"FC",X"17",X"C9",X"21",X"00",X"00",X"22",X"42",X"80",X"C9",X"E5",X"C5",X"3A",X"41",X"80",X"E6",
		X"0A",X"28",X"12",X"2A",X"42",X"80",X"09",X"CB",X"7C",X"28",X"03",X"21",X"FF",X"7F",X"22",X"42",
		X"80",X"DD",X"CB",X"00",X"C6",X"C1",X"E1",X"C9",X"E5",X"D5",X"21",X"00",X"00",X"3A",X"43",X"80",
		X"6F",X"CD",X"DD",X"17",X"65",X"DD",X"6E",X"1A",X"7C",X"B7",X"FE",X"08",X"30",X"03",X"21",X"00",
		X"00",X"22",X"42",X"80",X"D1",X"E1",X"C9",X"21",X"63",X"1E",X"DD",X"7E",X"0C",X"87",X"5F",X"16",
		X"00",X"19",X"5E",X"23",X"56",X"D5",X"FD",X"E1",X"DD",X"4E",X"0D",X"06",X"00",X"1E",X"07",X"16",
		X"00",X"79",X"B0",X"CA",X"DC",X"17",X"FD",X"19",X"0B",X"C3",X"D1",X"17",X"C9",X"D5",X"54",X"5D",
		X"B7",X"CB",X"15",X"CB",X"14",X"B7",X"CB",X"15",X"CB",X"14",X"19",X"B7",X"CB",X"1C",X"CB",X"1D",
		X"B7",X"CB",X"1C",X"CB",X"1D",X"B7",X"CB",X"1C",X"CB",X"1D",X"D1",X"C9",X"FD",X"7E",X"00",X"DD",
		X"77",X"01",X"FD",X"7E",X"01",X"DD",X"77",X"02",X"FD",X"7E",X"02",X"DD",X"77",X"12",X"FD",X"7E",
		X"03",X"DD",X"77",X"13",X"FD",X"7E",X"04",X"DD",X"77",X"14",X"FD",X"7E",X"05",X"DD",X"77",X"15",
		X"FD",X"7E",X"06",X"DD",X"77",X"16",X"C9",X"E5",X"D5",X"C5",X"DD",X"7E",X"19",X"CB",X"4F",X"CA",
		X"6C",X"18",X"DD",X"7E",X"01",X"B8",X"CA",X"6C",X"18",X"11",X"02",X"00",X"D2",X"42",X"18",X"11",
		X"FE",X"FF",X"D5",X"11",X"00",X"00",X"21",X"00",X"00",X"DD",X"6E",X"01",X"58",X"B7",X"ED",X"52",
		X"CD",X"C7",X"18",X"D1",X"7D",X"21",X"00",X"00",X"FE",X"01",X"28",X"06",X"38",X"04",X"19",X"3D",
		X"18",X"F6",X"11",X"00",X"00",X"DD",X"5E",X"04",X"19",X"DD",X"75",X"04",X"C1",X"D1",X"E1",X"C9",
		X"21",X"00",X"00",X"22",X"2F",X"80",X"3A",X"18",X"80",X"E6",X"03",X"FE",X"03",X"C2",X"89",X"18",
		X"2A",X"A2",X"1E",X"22",X"2F",X"80",X"C3",X"99",X"18",X"3A",X"1A",X"80",X"E6",X"03",X"FE",X"03",
		X"C2",X"99",X"18",X"2A",X"A6",X"1E",X"22",X"2F",X"80",X"C9",X"D5",X"E5",X"3A",X"3F",X"80",X"FE",
		X"00",X"C2",X"C4",X"18",X"2A",X"2F",X"80",X"DD",X"5E",X"05",X"DD",X"56",X"03",X"19",X"DD",X"75",
		X"05",X"DD",X"74",X"03",X"2A",X"31",X"80",X"DD",X"5E",X"06",X"DD",X"56",X"04",X"19",X"DD",X"75",
		X"06",X"DD",X"74",X"04",X"E1",X"D1",X"C9",X"D5",X"EB",X"B7",X"CB",X"7A",X"20",X"03",X"EB",X"18",
		X"06",X"21",X"00",X"00",X"B7",X"ED",X"52",X"D1",X"C9",X"D5",X"EB",X"21",X"00",X"00",X"B7",X"ED",
		X"52",X"D1",X"C9",X"E5",X"DD",X"E5",X"D5",X"21",X"00",X"00",X"22",X"5A",X"80",X"22",X"5C",X"80",
		X"DD",X"21",X"18",X"1C",X"2A",X"42",X"80",X"DD",X"56",X"01",X"DD",X"5E",X"00",X"B7",X"ED",X"52",
		X"CA",X"22",X"19",X"CB",X"7C",X"C2",X"22",X"19",X"DD",X"66",X"01",X"DD",X"6E",X"00",X"22",X"5C",
		X"80",X"DD",X"66",X"03",X"DD",X"6E",X"02",X"22",X"5A",X"80",X"11",X"04",X"00",X"DD",X"19",X"C3",
		X"F4",X"18",X"2A",X"42",X"80",X"ED",X"5B",X"5C",X"80",X"B7",X"ED",X"52",X"CA",X"4C",X"19",X"CB",
		X"7C",X"C2",X"4C",X"19",X"2A",X"5A",X"80",X"11",X"0A",X"00",X"19",X"22",X"5A",X"80",X"2A",X"5C",
		X"80",X"ED",X"5B",X"5A",X"80",X"19",X"22",X"5C",X"80",X"C3",X"22",X"19",X"D1",X"DD",X"E1",X"E1",
		X"C9",X"DD",X"E5",X"FD",X"E5",X"E5",X"D5",X"DD",X"21",X"6A",X"1C",X"3A",X"A1",X"81",X"87",X"11",
		X"00",X"00",X"5F",X"DD",X"19",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"E5",X"DD",X"E1",X"FD",X"21",
		X"43",X"1E",X"3A",X"29",X"80",X"FE",X"19",X"20",X"06",X"FD",X"21",X"4D",X"1E",X"18",X"08",X"FE",
		X"1A",X"20",X"04",X"FD",X"21",X"57",X"1E",X"DD",X"7E",X"00",X"FE",X"FF",X"CA",X"C7",X"1A",X"21",
		X"00",X"00",X"11",X"00",X"00",X"DD",X"6E",X"00",X"FD",X"46",X"03",X"FD",X"4E",X"02",X"09",X"3A",
		X"2B",X"80",X"5F",X"B7",X"ED",X"52",X"CA",X"BF",X"1A",X"D2",X"BF",X"1A",X"CD",X"C7",X"18",X"22",
		X"5E",X"80",X"21",X"00",X"00",X"DD",X"6E",X"01",X"FD",X"46",X"05",X"FD",X"4E",X"04",X"09",X"B7",
		X"ED",X"52",X"CA",X"BF",X"1A",X"DA",X"BF",X"1A",X"22",X"60",X"80",X"21",X"00",X"00",X"DD",X"6E",
		X"02",X"FD",X"46",X"07",X"FD",X"4E",X"06",X"09",X"11",X"00",X"00",X"3A",X"2C",X"80",X"5F",X"B7",
		X"ED",X"52",X"CA",X"BF",X"1A",X"D2",X"BF",X"1A",X"CD",X"C7",X"18",X"22",X"62",X"80",X"21",X"00",
		X"00",X"DD",X"6E",X"03",X"FD",X"46",X"09",X"FD",X"4E",X"08",X"09",X"B7",X"ED",X"52",X"CA",X"BF",
		X"1A",X"DA",X"BF",X"1A",X"22",X"64",X"80",X"2A",X"5E",X"80",X"ED",X"5B",X"60",X"80",X"44",X"4D",
		X"B7",X"ED",X"52",X"38",X"0A",X"42",X"4B",X"21",X"00",X"00",X"22",X"5E",X"80",X"18",X"06",X"21",
		X"00",X"00",X"22",X"60",X"80",X"2A",X"62",X"80",X"ED",X"5B",X"64",X"80",X"B7",X"ED",X"52",X"38",
		X"08",X"21",X"00",X"00",X"22",X"62",X"80",X"18",X"0A",X"ED",X"5B",X"62",X"80",X"21",X"00",X"00",
		X"22",X"64",X"80",X"60",X"69",X"B7",X"ED",X"52",X"38",X"0B",X"21",X"00",X"00",X"22",X"5E",X"80",
		X"22",X"60",X"80",X"18",X"09",X"21",X"00",X"00",X"22",X"62",X"80",X"22",X"64",X"80",X"2A",X"5E",
		X"80",X"7C",X"B5",X"28",X"13",X"21",X"00",X"00",X"DD",X"6E",X"00",X"FD",X"56",X"03",X"FD",X"5E",
		X"02",X"19",X"7D",X"32",X"2B",X"80",X"18",X"5E",X"2A",X"60",X"80",X"7C",X"B5",X"28",X"13",X"21",
		X"00",X"00",X"DD",X"6E",X"01",X"FD",X"56",X"05",X"FD",X"5E",X"04",X"19",X"7D",X"32",X"2B",X"80",
		X"18",X"44",X"2A",X"62",X"80",X"7C",X"B5",X"28",X"13",X"21",X"00",X"00",X"DD",X"6E",X"02",X"FD",
		X"56",X"07",X"FD",X"5E",X"06",X"19",X"7D",X"32",X"2C",X"80",X"18",X"2A",X"21",X"00",X"00",X"DD",
		X"6E",X"03",X"FD",X"56",X"09",X"FD",X"5E",X"08",X"19",X"7D",X"32",X"2C",X"80",X"18",X"17",X"11",
		X"04",X"00",X"DD",X"19",X"C3",X"87",X"19",X"DD",X"7E",X"01",X"FE",X"FF",X"CA",X"D6",X"1A",X"DD",
		X"21",X"31",X"1E",X"C3",X"87",X"19",X"D1",X"E1",X"FD",X"E1",X"DD",X"E1",X"C9",X"C5",X"D5",X"11",
		X"00",X"00",X"3A",X"02",X"85",X"C6",X"04",X"47",X"3A",X"03",X"85",X"C6",X"00",X"4F",X"CD",X"DE",
		X"00",X"7E",X"CD",X"AF",X"1B",X"FE",X"00",X"28",X"02",X"CB",X"CB",X"3A",X"02",X"85",X"C6",X"0C",
		X"47",X"3A",X"03",X"85",X"C6",X"00",X"4F",X"CD",X"DE",X"00",X"7E",X"CD",X"AF",X"1B",X"FE",X"00",
		X"28",X"02",X"CB",X"CB",X"3A",X"02",X"85",X"C6",X"04",X"47",X"3A",X"03",X"85",X"C6",X"0F",X"4F",
		X"CD",X"DE",X"00",X"7E",X"CD",X"AF",X"1B",X"FE",X"00",X"28",X"02",X"CB",X"DB",X"3A",X"02",X"85",
		X"C6",X"0C",X"47",X"3A",X"03",X"85",X"C6",X"0F",X"4F",X"CD",X"DE",X"00",X"7E",X"CD",X"AF",X"1B",
		X"FE",X"00",X"28",X"02",X"CB",X"DB",X"3A",X"02",X"85",X"C6",X"02",X"47",X"3A",X"03",X"85",X"C6",
		X"04",X"4F",X"CD",X"DE",X"00",X"7E",X"CD",X"D8",X"1B",X"FE",X"00",X"28",X"02",X"CB",X"C3",X"3A",
		X"02",X"85",X"C6",X"02",X"47",X"3A",X"03",X"85",X"C6",X"0C",X"4F",X"CD",X"DE",X"00",X"7E",X"CD",
		X"D8",X"1B",X"FE",X"00",X"28",X"02",X"CB",X"C3",X"3A",X"02",X"85",X"C6",X"0D",X"47",X"3A",X"03",
		X"85",X"C6",X"04",X"4F",X"CD",X"DE",X"00",X"7E",X"CD",X"D8",X"1B",X"FE",X"00",X"28",X"02",X"CB",
		X"C3",X"3A",X"02",X"85",X"C6",X"0D",X"47",X"3A",X"03",X"85",X"C6",X"0C",X"4F",X"CD",X"DE",X"00",
		X"7E",X"CD",X"D8",X"1B",X"FE",X"00",X"28",X"02",X"CB",X"C3",X"62",X"6B",X"D1",X"C1",X"C9",X"FE",
		X"60",X"38",X"22",X"FE",X"80",X"38",X"08",X"FE",X"A0",X"38",X"1A",X"FE",X"C0",X"30",X"16",X"E6",
		X"0F",X"FE",X"06",X"38",X"0C",X"FE",X"08",X"38",X"0C",X"FE",X"0C",X"38",X"04",X"FE",X"0E",X"38",
		X"04",X"3E",X"01",X"18",X"02",X"3E",X"00",X"C9",X"FE",X"60",X"38",X"1E",X"FE",X"80",X"38",X"08",
		X"FE",X"A0",X"38",X"16",X"FE",X"C0",X"30",X"12",X"E6",X"0F",X"FE",X"02",X"38",X"08",X"FE",X"04",
		X"38",X"08",X"FE",X"0E",X"30",X"04",X"3E",X"01",X"18",X"02",X"3E",X"00",X"C9",X"C5",X"FE",X"13",
		X"28",X"06",X"FE",X"93",X"28",X"02",X"18",X"08",X"47",X"3A",X"89",X"80",X"B8",X"28",X"07",X"78",
		X"32",X"89",X"80",X"CD",X"FC",X"00",X"C1",X"C9",X"96",X"00",X"32",X"00",X"C2",X"01",X"5A",X"00",
		X"8E",X"03",X"82",X"00",X"FA",X"05",X"AA",X"00",X"06",X"09",X"D2",X"00",X"B2",X"0C",X"FA",X"00",
		X"FE",X"10",X"22",X"01",X"EA",X"15",X"4A",X"01",X"76",X"1B",X"72",X"01",X"A2",X"21",X"9A",X"01",
		X"6E",X"28",X"C2",X"01",X"DA",X"2F",X"EA",X"01",X"E6",X"37",X"12",X"02",X"92",X"40",X"3A",X"02",
		X"DE",X"49",X"62",X"02",X"CA",X"53",X"8A",X"02",X"56",X"5E",X"B2",X"02",X"82",X"69",X"DA",X"02",
		X"4E",X"75",X"02",X"03",X"BA",X"81",X"2A",X"03",X"FF",X"FF",X"8C",X"1C",X"A1",X"1C",X"B2",X"1C",
		X"C7",X"1C",X"E9",X"1C",X"EA",X"1C",X"13",X"1D",X"2C",X"1D",X"3D",X"1D",X"52",X"1D",X"63",X"1D",
		X"94",X"1D",X"AD",X"1D",X"C6",X"1D",X"E7",X"1D",X"00",X"1E",X"FF",X"FF",X"7B",X"BD",X"31",X"46",
		X"33",X"5D",X"49",X"5E",X"63",X"9D",X"91",X"A6",X"1B",X"45",X"A9",X"BE",X"83",X"D5",X"C1",X"D6",
		X"FF",X"53",X"9D",X"31",X"46",X"33",X"45",X"51",X"9E",X"AB",X"BD",X"51",X"9E",X"53",X"9D",X"A9",
		X"BE",X"FF",X"6B",X"9D",X"31",X"46",X"0B",X"55",X"49",X"5E",X"9B",X"CD",X"61",X"76",X"93",X"A5",
		X"61",X"A6",X"33",X"A5",X"91",X"A6",X"FF",X"4B",X"5D",X"21",X"5E",X"93",X"A5",X"21",X"5E",X"23",
		X"5D",X"49",X"5E",X"93",X"CD",X"49",X"5E",X"23",X"55",X"91",X"A6",X"9B",X"CD",X"91",X"A6",X"4B",
		X"5D",X"91",X"CE",X"93",X"A5",X"91",X"CE",X"FF",X"00",X"FF",X"1B",X"45",X"31",X"46",X"63",X"8D",
		X"31",X"46",X"AB",X"D5",X"31",X"46",X"3B",X"6D",X"61",X"76",X"83",X"B5",X"61",X"76",X"1B",X"45",
		X"91",X"A6",X"63",X"8D",X"91",X"A6",X"AB",X"D5",X"91",X"A6",X"3B",X"6D",X"C1",X"D6",X"83",X"B5",
		X"C1",X"D6",X"FF",X"63",X"8D",X"31",X"46",X"33",X"6D",X"61",X"76",X"83",X"BD",X"61",X"76",X"33",
		X"6D",X"79",X"8E",X"83",X"BD",X"79",X"8E",X"63",X"8D",X"A9",X"BE",X"FF",X"23",X"55",X"31",X"46",
		X"9B",X"CD",X"31",X"46",X"23",X"55",X"A9",X"BE",X"9B",X"CD",X"A9",X"BE",X"FF",X"3B",X"6D",X"31",
		X"46",X"83",X"B5",X"31",X"46",X"63",X"8D",X"91",X"A6",X"1B",X"45",X"A9",X"BE",X"AB",X"D5",X"A9",
		X"BE",X"FF",X"3B",X"B5",X"31",X"46",X"33",X"45",X"31",X"9E",X"AB",X"BD",X"31",X"9E",X"63",X"8D",
		X"91",X"A6",X"FF",X"6B",X"85",X"19",X"2E",X"63",X"75",X"19",X"46",X"63",X"8D",X"31",X"46",X"4B",
		X"8D",X"49",X"5E",X"63",X"75",X"49",X"76",X"63",X"8D",X"61",X"76",X"6B",X"BD",X"79",X"8E",X"63",
		X"75",X"79",X"A6",X"63",X"8D",X"91",X"A6",X"1B",X"8D",X"A9",X"BE",X"63",X"75",X"B1",X"D6",X"63",
		X"8D",X"C1",X"D6",X"FF",X"0B",X"3D",X"49",X"5E",X"B3",X"E5",X"49",X"5E",X"23",X"55",X"79",X"8E",
		X"9B",X"CD",X"79",X"8E",X"3B",X"6D",X"A9",X"BE",X"83",X"B5",X"A9",X"BE",X"FF",X"3B",X"85",X"31",
		X"46",X"93",X"B5",X"31",X"46",X"33",X"45",X"31",X"BE",X"AB",X"BD",X"31",X"BE",X"33",X"5D",X"A9",
		X"BE",X"6B",X"BD",X"A9",X"BE",X"FF",X"33",X"85",X"19",X"2E",X"7B",X"8D",X"19",X"5E",X"23",X"5D",
		X"61",X"76",X"1B",X"2D",X"61",X"BE",X"C3",X"D5",X"31",X"8E",X"93",X"D5",X"79",X"8E",X"63",X"75",
		X"91",X"D6",X"63",X"BD",X"C1",X"D6",X"FF",X"B3",X"E5",X"31",X"46",X"0B",X"3D",X"49",X"5E",X"B3",
		X"E5",X"61",X"76",X"0B",X"3D",X"79",X"8E",X"B3",X"E5",X"91",X"A6",X"0B",X"3D",X"A9",X"BE",X"FF",
		X"3B",X"6D",X"19",X"2E",X"83",X"B5",X"19",X"2E",X"1B",X"2D",X"39",X"6E",X"C3",X"D5",X"39",X"6E",
		X"1B",X"2D",X"81",X"B6",X"C3",X"D5",X"81",X"B6",X"63",X"8D",X"49",X"5E",X"4B",X"5D",X"61",X"8E",
		X"93",X"A5",X"61",X"8E",X"63",X"8D",X"91",X"A6",X"3B",X"6D",X"C1",X"D6",X"83",X"B5",X"C1",X"D6",
		X"FF",X"04",X"FD",X"04",X"16",X"04",X"15",X"04",X"FE",X"DB",X"FD",X"04",X"FE",X"04",X"FD",X"D9",
		X"FE",X"FF",X"FF",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"00",X"FF",
		X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"1A",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",
		X"FF",X"FF",X"FF",X"67",X"1E",X"6A",X"1E",X"18",X"00",X"FF",X"1A",X"00",X"20",X"04",X"FF",X"FF",
		X"00",X"19",X"00",X"28",X"04",X"FF",X"FF",X"00",X"18",X"00",X"04",X"04",X"FF",X"FF",X"00",X"18",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"10",X"00",X"08",X"00",X"F0",X"FF",X"F8",X"FF",X"80",X"01",
		X"FF",X"FF",X"08",X"00",X"10",X"00",X"20",X"00",X"30",X"00",X"01",X"00",X"FF",X"FF",X"02",X"00",
		X"FE",X"FF",X"80",X"01",X"00",X"00",X"80",X"FE",X"00",X"00",X"D9",X"00",X"D8",X"00",X"D7",X"00",
		X"D6",X"00",X"33",X"00",X"34",X"00",X"35",X"00",X"D5",X"FF",X"C0",X"FF",X"00",X"FF",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CD",X"9F",X"02",X"3A",X"03",X"B0",X"C3",X"CB",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3A",X"03",X"B0",X"3A",X"00",X"B0",X"C3",X"27",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3A",X"03",X"B0",X"3A",X"00",X"B0",X"C3",X"5C",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3A",X"03",X"B0",X"3A",X"00",X"B0",X"C3",X"A4",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3A",X"03",X"B0",X"3A",X"00",X"B0",X"C3",X"1F",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3A",X"03",X"B0",X"3A",X"00",X"B0",X"C3",X"4C",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3A",X"03",X"B0",X"3A",X"00",X"B0",X"C3",X"60",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"32",X"03",X"B0",X"DD",X"36",X"00",X"30",X"C3",X"F8",X"05",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3A",X"03",X"B0",X"3A",X"00",X"B0",X"C3",X"72",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3A",X"03",X"B0",X"3A",X"00",X"B0",X"C3",X"8B",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3A",X"03",X"B0",X"3A",X"00",X"B0",X"C3",X"98",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3A",X"03",X"B0",X"11",X"08",X"00",X"C3",X"FC",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CD",X"D2",X"00",X"3A",X"03",X"B0",X"C3",X"F9",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C3",X"C7",X"18",X"C3",X"D9",X"18",X"00",X"3A",X"03",X"B0",X"CD",X"02",X"06",X"C3",X"AB",X"05");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
