library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity gfx1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of gfx1 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"CC",X"66",X"33",X"33",X"33",X"22",X"CC",X"00",X"11",X"22",X"66",X"66",X"66",X"33",X"11",X"00",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"FF",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"33",X"00",
		X"EE",X"33",X"77",X"EE",X"CC",X"00",X"FF",X"00",X"33",X"66",X"00",X"11",X"33",X"77",X"77",X"00",
		X"FF",X"66",X"CC",X"EE",X"33",X"33",X"EE",X"00",X"33",X"00",X"00",X"11",X"00",X"66",X"33",X"00",
		X"EE",X"EE",X"66",X"66",X"FF",X"66",X"66",X"00",X"00",X"11",X"33",X"66",X"77",X"00",X"00",X"00",
		X"EE",X"00",X"EE",X"33",X"33",X"33",X"EE",X"00",X"77",X"66",X"77",X"00",X"00",X"66",X"33",X"00",
		X"EE",X"00",X"00",X"EE",X"33",X"33",X"EE",X"00",X"11",X"33",X"66",X"77",X"66",X"66",X"33",X"00",
		X"FF",X"33",X"66",X"CC",X"88",X"88",X"88",X"00",X"77",X"66",X"00",X"00",X"11",X"11",X"11",X"00",
		X"CC",X"22",X"22",X"CC",X"FF",X"33",X"EE",X"00",X"33",X"66",X"77",X"33",X"44",X"44",X"33",X"00",
		X"EE",X"33",X"33",X"FF",X"33",X"66",X"CC",X"00",X"33",X"66",X"66",X"33",X"00",X"00",X"33",X"00",
		X"CC",X"66",X"33",X"33",X"FF",X"33",X"33",X"00",X"11",X"33",X"66",X"66",X"77",X"66",X"66",X"00",
		X"EE",X"33",X"33",X"EE",X"33",X"33",X"EE",X"00",X"77",X"66",X"66",X"77",X"66",X"66",X"77",X"00",
		X"EE",X"33",X"00",X"00",X"00",X"33",X"EE",X"00",X"11",X"33",X"66",X"66",X"66",X"33",X"11",X"00",
		X"CC",X"66",X"33",X"33",X"33",X"66",X"CC",X"00",X"77",X"66",X"66",X"66",X"66",X"66",X"77",X"00",
		X"FF",X"00",X"00",X"EE",X"00",X"00",X"FF",X"00",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"00",
		X"FF",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"77",X"66",X"66",X"77",X"66",X"66",X"66",X"00",
		X"FF",X"00",X"00",X"77",X"33",X"33",X"FF",X"00",X"11",X"33",X"66",X"66",X"66",X"33",X"11",X"00",
		X"33",X"33",X"33",X"FF",X"33",X"33",X"33",X"00",X"66",X"66",X"66",X"77",X"66",X"66",X"66",X"00",
		X"FF",X"CC",X"CC",X"CC",X"CC",X"CC",X"FF",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"33",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"33",X"00",
		X"33",X"66",X"CC",X"88",X"CC",X"EE",X"77",X"00",X"66",X"66",X"66",X"77",X"77",X"66",X"66",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"00",
		X"33",X"77",X"FF",X"FF",X"BB",X"33",X"33",X"00",X"66",X"77",X"77",X"77",X"66",X"66",X"66",X"00",
		X"33",X"33",X"BB",X"FF",X"FF",X"77",X"33",X"00",X"66",X"77",X"77",X"77",X"66",X"66",X"66",X"00",
		X"EE",X"33",X"33",X"33",X"33",X"33",X"EE",X"00",X"33",X"66",X"66",X"66",X"66",X"66",X"33",X"00",
		X"EE",X"33",X"33",X"33",X"EE",X"00",X"00",X"00",X"77",X"66",X"66",X"66",X"77",X"66",X"66",X"00",
		X"EE",X"33",X"33",X"33",X"FF",X"66",X"DD",X"00",X"33",X"66",X"66",X"66",X"66",X"66",X"33",X"00",
		X"EE",X"33",X"33",X"77",X"CC",X"EE",X"77",X"00",X"77",X"66",X"66",X"66",X"77",X"66",X"66",X"00",
		X"CC",X"66",X"00",X"EE",X"33",X"33",X"EE",X"00",X"33",X"66",X"66",X"33",X"00",X"66",X"33",X"00",
		X"FF",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"EE",X"00",X"66",X"66",X"66",X"66",X"66",X"66",X"33",X"00",
		X"33",X"33",X"33",X"77",X"EE",X"CC",X"88",X"00",X"66",X"66",X"66",X"77",X"33",X"11",X"00",X"00",
		X"33",X"33",X"BB",X"FF",X"FF",X"77",X"33",X"00",X"66",X"66",X"66",X"77",X"77",X"77",X"66",X"00",
		X"33",X"77",X"EE",X"CC",X"EE",X"77",X"33",X"00",X"66",X"77",X"33",X"11",X"33",X"77",X"66",X"00",
		X"33",X"33",X"33",X"EE",X"CC",X"CC",X"CC",X"00",X"33",X"33",X"33",X"11",X"00",X"00",X"00",X"00",
		X"FF",X"77",X"EE",X"CC",X"88",X"00",X"FF",X"00",X"77",X"00",X"00",X"11",X"33",X"77",X"77",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"00",
		X"0F",X"69",X"69",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"CC",X"22",X"99",X"11",X"11",X"99",X"22",X"CC",X"33",X"44",X"99",X"AA",X"AA",X"99",X"44",X"33",
		X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"07",X"07",X"00",X"0F",X"0F",X"0C",X"0F",X"0F",X"08",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"01",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"0F",X"0F",X"03",X"0F",X"0F",X"03",X"0F",X"0F",
		X"0F",X"0F",X"09",X"09",X"09",X"09",X"09",X"09",X"0F",X"0F",X"09",X"09",X"09",X"09",X"09",X"09",
		X"0F",X"0F",X"08",X"08",X"08",X"08",X"0F",X"0F",X"00",X"09",X"09",X"09",X"09",X"09",X"09",X"08",
		X"03",X"07",X"06",X"06",X"06",X"06",X"07",X"03",X"0E",X"0E",X"00",X"00",X"00",X"00",X"0E",X"0E",
		X"08",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"08",X"0F",X"0F",X"00",X"00",X"00",X"00",X"0F",X"0F",
		X"00",X"10",X"10",X"10",X"30",X"21",X"61",X"43",X"00",X"00",X"00",X"00",X"00",X"01",X"10",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"81",X"D0",X"58",
		X"D2",X"F0",X"74",X"76",X"30",X"03",X"00",X"00",X"51",X"70",X"71",X"16",X"10",X"00",X"00",X"00",
		X"40",X"C0",X"C0",X"0C",X"00",X"00",X"00",X"00",X"79",X"F0",X"D5",X"DC",X"90",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"00",
		X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"77",X"11",X"11",X"11",X"11",X"11",X"11",X"00",X"FF",X"66",X"66",X"66",X"66",X"66",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"68",X"68",X"68",X"68",X"68",X"F8",X"00",X"E7",X"81",X"81",X"81",X"81",X"81",X"81",X"00",
		X"CF",X"69",X"69",X"69",X"69",X"69",X"CF",X"00",X"3C",X"6D",X"6D",X"6D",X"6D",X"6D",X"3C",X"00",
		X"62",X"62",X"6A",X"EE",X"EE",X"E6",X"62",X"00",X"C2",X"EB",X"FB",X"FB",X"DA",X"CA",X"C2",X"00",
		X"00",X"06",X"06",X"00",X"00",X"60",X"60",X"00",X"00",X"66",X"66",X"00",X"00",X"06",X"06",X"00",
		X"00",X"60",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"66",X"66",X"00",
		X"00",X"00",X"22",X"44",X"88",X"44",X"22",X"00",X"00",X"00",X"22",X"11",X"00",X"11",X"22",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"60",X"80",X"40",X"40",X"20",X"10",X"00",X"00",X"00",
		X"10",X"10",X"10",X"10",X"10",X"10",X"BA",X"FE",X"00",X"80",X"40",X"40",X"60",X"31",X"31",X"10",
		X"00",X"00",X"10",X"10",X"20",X"40",X"40",X"D1",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"C4",
		X"00",X"10",X"20",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"20",X"C8",
		X"30",X"10",X"11",X"00",X"C0",X"30",X"22",X"01",X"00",X"00",X"40",X"30",X"10",X"00",X"00",X"00",
		X"F2",X"F2",X"FB",X"0E",X"05",X"07",X"0F",X"0F",X"10",X"D5",X"F3",X"E9",X"77",X"D5",X"01",X"0F",
		X"F6",X"F9",X"E2",X"E6",X"FF",X"F8",X"F1",X"FF",X"E6",X"F3",X"F4",X"BC",X"3E",X"19",X"07",X"0D",
		X"00",X"60",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"10",X"F8",X"C0",X"88",X"00",X"00",
		X"33",X"F0",X"74",X"11",X"31",X"40",X"80",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"10",X"20",
		X"0F",X"0F",X"03",X"0E",X"1B",X"FB",X"F2",X"F4",X"FF",X"01",X"E7",X"CE",X"EE",X"FF",X"F9",X"F1",
		X"11",X"7F",X"FC",X"7C",X"FB",X"FF",X"F3",X"F1",X"0E",X"0F",X"0B",X"8C",X"E6",X"D5",X"D1",X"F7",
		X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"F0",X"E4",X"CC",X"00",X"80",X"C0",X"B8",
		X"10",X"10",X"31",X"62",X"80",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"30",X"40",X"80",
		X"F4",X"FC",X"B8",X"20",X"20",X"20",X"20",X"00",X"F2",X"BA",X"32",X"64",X"40",X"80",X"00",X"00",
		X"F8",X"FC",X"FF",X"99",X"00",X"80",X"80",X"40",X"F5",X"FC",X"FE",X"32",X"10",X"00",X"00",X"00",
		X"80",X"60",X"00",X"00",X"00",X"80",X"60",X"10",X"00",X"80",X"C0",X"E8",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C4",X"62",X"22",X"31",X"00",X"00",X"00",X"20",X"10",X"00",X"00",X"00",
		X"00",X"00",X"10",X"10",X"31",X"03",X"04",X"5B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"9C",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"57",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"EC",X"C8",X"80",X"00",
		X"00",X"01",X"01",X"01",X"02",X"12",X"89",X"57",X"00",X"00",X"00",X"00",X"00",X"30",X"11",X"00",
		X"99",X"1F",X"09",X"8F",X"52",X"0B",X"97",X"2D",X"2F",X"77",X"74",X"D7",X"4D",X"05",X"4A",X"85",
		X"38",X"3D",X"3F",X"46",X"69",X"CE",X"8B",X"53",X"69",X"4E",X"DD",X"29",X"9F",X"8A",X"1D",X"0F",
		X"00",X"00",X"00",X"20",X"C0",X"00",X"00",X"00",X"00",X"04",X"08",X"19",X"22",X"3A",X"04",X"8A",
		X"25",X"24",X"15",X"2B",X"0A",X"12",X"15",X"37",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"4F",X"2D",X"4F",X"AB",X"06",X"6E",X"BC",X"A6",X"09",X"0E",X"A8",X"67",X"D6",X"E9",X"E2",
		X"8D",X"D7",X"5D",X"CD",X"2E",X"46",X"8D",X"46",X"8E",X"4B",X"3C",X"37",X"4B",X"EF",X"2A",X"15",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"8A",X"06",X"04",X"4E",X"8E",X"08",X"CC",X"44",
		X"12",X"03",X"71",X"F7",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"31",X"40",X"00",
		X"15",X"82",X"1E",X"32",X"32",X"20",X"20",X"00",X"85",X"03",X"0C",X"03",X"00",X"00",X"00",X"00",
		X"4D",X"E9",X"0E",X"00",X"00",X"00",X"00",X"00",X"4D",X"97",X"81",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"C0",X"40",X"00",X"00",X"40",X"C8",X"E8",X"32",X"11",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"62",X"73",X"78",X"80",X"40",X"20",X"10",X"00",X"00",X"04",X"02",
		X"00",X"00",X"00",X"0C",X"94",X"F9",X"4B",X"0F",X"00",X"02",X"01",X"00",X"06",X"3C",X"7B",X"87",
		X"00",X"00",X"00",X"01",X"86",X"E9",X"7C",X"0F",X"80",X"80",X"86",X"C2",X"BC",X"9F",X"0F",X"0F",
		X"10",X"20",X"40",X"80",X"08",X"08",X"08",X"04",X"00",X"02",X"04",X"08",X"15",X"7B",X"E5",X"6D",
		X"7A",X"87",X"4B",X"37",X"4B",X"4B",X"8F",X"87",X"01",X"01",X"00",X"00",X"80",X"40",X"31",X"10",
		X"0F",X"0F",X"1B",X"09",X"0D",X"0F",X"0F",X"07",X"0D",X"0F",X"0F",X"8F",X"4D",X"09",X"0F",X"0F",
		X"1F",X"A7",X"C3",X"4B",X"1E",X"2D",X"0F",X"0F",X"0E",X"0C",X"0D",X"08",X"09",X"0B",X"0B",X"0F",
		X"04",X"08",X"18",X"20",X"40",X"80",X"88",X"00",X"4E",X"2E",X"4E",X"8E",X"4A",X"3C",X"3D",X"BF",
		X"0F",X"0C",X"0F",X"0F",X"C7",X"5B",X"30",X"05",X"10",X"13",X"21",X"31",X"12",X"01",X"00",X"00",
		X"03",X"81",X"0B",X"8E",X"8F",X"0B",X"03",X"0B",X"07",X"4F",X"2F",X"1F",X"0F",X"8F",X"CE",X"8F",
		X"4F",X"8F",X"0F",X"2D",X"4B",X"9F",X"0B",X"09",X"0B",X"11",X"43",X"61",X"3C",X"0F",X"1E",X"0F",
		X"08",X"08",X"84",X"04",X"08",X"08",X"08",X"04",X"1F",X"2F",X"2E",X"5F",X"9F",X"2D",X"1E",X"7E",
		X"09",X"10",X"32",X"76",X"65",X"42",X"80",X"00",X"01",X"02",X"02",X"00",X"00",X"00",X"00",X"10",
		X"0F",X"0F",X"17",X"7E",X"E9",X"2C",X"20",X"20",X"87",X"C7",X"CF",X"BC",X"06",X"01",X"02",X"00",
		X"0F",X"0F",X"EF",X"E3",X"34",X"07",X"00",X"00",X"8F",X"4F",X"3C",X"C2",X"09",X"06",X"00",X"00",
		X"02",X"00",X"00",X"00",X"08",X"80",X"40",X"20",X"6C",X"2C",X"6C",X"E9",X"1E",X"00",X"08",X"00",
		X"00",X"00",X"01",X"16",X"61",X"30",X"C3",X"E1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"80",X"80",X"C0",X"E8",X"00",X"00",X"04",X"C0",X"C0",X"F7",X"FE",X"F3",X"3C",
		X"ED",X"FE",X"FF",X"C3",X"3C",X"80",X"00",X"00",X"71",X"30",X"01",X"10",X"00",X"10",X"30",X"00",
		X"00",X"68",X"C0",X"E0",X"CA",X"C0",X"08",X"60",X"1E",X"0F",X"B4",X"F2",X"B7",X"25",X"10",X"00",
		X"00",X"30",X"F0",X"78",X"3C",X"B4",X"3C",X"D2",X"00",X"00",X"10",X"21",X"70",X"30",X"F0",X"F0",
		X"00",X"E0",X"C0",X"E8",X"88",X"F0",X"2C",X"F0",X"00",X"F6",X"F8",X"79",X"69",X"DE",X"E1",X"96",
		X"85",X"48",X"DE",X"F0",X"A5",X"61",X"30",X"10",X"73",X"74",X"61",X"10",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"68",X"FC",X"E0",X"C0",X"08",X"00",X"2C",X"A1",X"3C",X"B5",X"D2",X"E7",X"F0",X"F0",
		X"52",X"70",X"78",X"F0",X"96",X"F0",X"F0",X"78",X"00",X"00",X"70",X"03",X"34",X"43",X"D2",X"78",
		X"80",X"A4",X"E0",X"F8",X"88",X"78",X"A4",X"D2",X"E1",X"3C",X"F0",X"79",X"E1",X"FC",X"F0",X"F0",
		X"F0",X"78",X"F8",X"A5",X"D2",X"E1",X"D2",X"61",X"73",X"D6",X"34",X"10",X"07",X"21",X"10",X"00",
		X"2C",X"E0",X"E0",X"FC",X"E0",X"C0",X"08",X"00",X"F0",X"E1",X"F0",X"97",X"F0",X"F6",X"B4",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"EE",X"CC",X"88",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"60",X"80",X"40",X"40",X"20",X"10",X"00",X"00",X"00",
		X"10",X"10",X"10",X"10",X"10",X"10",X"BA",X"FE",X"00",X"80",X"40",X"40",X"60",X"31",X"31",X"10",
		X"00",X"00",X"10",X"10",X"20",X"40",X"40",X"D1",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"C4",
		X"00",X"10",X"20",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"20",X"C8",
		X"30",X"10",X"11",X"00",X"C0",X"30",X"22",X"01",X"00",X"00",X"40",X"30",X"10",X"00",X"00",X"00",
		X"F2",X"F2",X"FB",X"0E",X"05",X"07",X"0F",X"0F",X"10",X"D5",X"F3",X"E9",X"77",X"D5",X"01",X"0F",
		X"F6",X"F9",X"E2",X"E6",X"FF",X"F8",X"F1",X"FF",X"E6",X"F3",X"F4",X"BC",X"3E",X"19",X"07",X"0D",
		X"00",X"60",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"10",X"F8",X"C0",X"88",X"00",X"00",
		X"33",X"F0",X"74",X"11",X"31",X"40",X"80",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"10",X"20",
		X"0F",X"0F",X"03",X"0E",X"1B",X"FB",X"F2",X"F4",X"FF",X"01",X"E7",X"CE",X"EE",X"FF",X"F9",X"F1",
		X"11",X"7F",X"FC",X"7C",X"FB",X"FF",X"F3",X"F1",X"0E",X"0F",X"0B",X"8C",X"E6",X"D5",X"D1",X"F7",
		X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"F0",X"E4",X"CC",X"00",X"80",X"C0",X"B8",
		X"10",X"10",X"31",X"62",X"80",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"30",X"40",X"80",
		X"F4",X"FC",X"B8",X"20",X"20",X"20",X"20",X"00",X"F2",X"BA",X"32",X"64",X"40",X"80",X"00",X"00",
		X"F8",X"FC",X"FF",X"99",X"00",X"80",X"80",X"40",X"F5",X"FC",X"FE",X"32",X"10",X"00",X"00",X"00",
		X"80",X"60",X"00",X"00",X"00",X"80",X"60",X"10",X"00",X"80",X"C0",X"E8",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C4",X"62",X"22",X"31",X"00",X"00",X"00",X"20",X"10",X"00",X"00",X"00",
		X"00",X"00",X"10",X"10",X"31",X"03",X"04",X"5B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"9C",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"57",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"EC",X"C8",X"80",X"00",
		X"00",X"01",X"01",X"01",X"02",X"12",X"89",X"57",X"00",X"00",X"00",X"00",X"00",X"30",X"11",X"00",
		X"99",X"1F",X"09",X"8F",X"52",X"0B",X"97",X"2D",X"2F",X"77",X"74",X"D7",X"4D",X"05",X"4A",X"85",
		X"38",X"3D",X"3F",X"46",X"69",X"CE",X"8B",X"53",X"69",X"4E",X"DD",X"29",X"9F",X"8A",X"1D",X"0F",
		X"00",X"00",X"00",X"20",X"C0",X"00",X"00",X"00",X"00",X"04",X"08",X"19",X"22",X"3A",X"04",X"8A",
		X"25",X"24",X"15",X"2B",X"0A",X"12",X"15",X"37",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"4F",X"2D",X"4F",X"AB",X"06",X"6E",X"BC",X"A6",X"09",X"0E",X"A8",X"67",X"D6",X"E9",X"E2",
		X"8D",X"D7",X"5D",X"CD",X"2E",X"46",X"8D",X"46",X"8E",X"4B",X"3C",X"37",X"4B",X"EF",X"2A",X"15",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"8A",X"06",X"04",X"4E",X"8E",X"08",X"CC",X"44",
		X"12",X"03",X"71",X"F7",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"31",X"40",X"00",
		X"15",X"82",X"1E",X"32",X"32",X"20",X"20",X"00",X"85",X"03",X"0C",X"03",X"00",X"00",X"00",X"00",
		X"4D",X"E9",X"0E",X"00",X"00",X"00",X"00",X"00",X"4D",X"97",X"81",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"C0",X"40",X"00",X"00",X"40",X"C8",X"E8",X"32",X"11",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"22",X"11",X"48",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"02",
		X"00",X"00",X"00",X"0C",X"94",X"F9",X"4B",X"0F",X"00",X"02",X"01",X"00",X"06",X"3C",X"7B",X"87",
		X"00",X"00",X"00",X"01",X"86",X"C8",X"4C",X"0C",X"80",X"80",X"86",X"C2",X"BC",X"9F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"04",X"00",X"02",X"04",X"08",X"04",X"19",X"21",X"09",
		X"6A",X"87",X"4B",X"26",X"4B",X"4B",X"8F",X"87",X"01",X"01",X"00",X"00",X"00",X"00",X"11",X"00",
		X"0F",X"0F",X"1B",X"09",X"0D",X"07",X"03",X"00",X"0D",X"07",X"00",X"00",X"00",X"09",X"0F",X"0C",
		X"0C",X"84",X"C0",X"4A",X"16",X"21",X"03",X"07",X"0E",X"08",X"01",X"00",X"00",X"08",X"08",X"03",
		X"04",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"26",X"46",X"8E",X"4A",X"3C",X"2C",X"8C",
		X"07",X"08",X"0C",X"0C",X"C4",X"48",X"20",X"05",X"10",X"13",X"21",X"31",X"12",X"01",X"00",X"00",
		X"02",X"00",X"09",X"8C",X"8D",X"09",X"00",X"0B",X"06",X"4F",X"27",X"17",X"03",X"01",X"88",X"8F",
		X"4C",X"8C",X"0E",X"21",X"01",X"11",X"01",X"09",X"0B",X"11",X"02",X"20",X"08",X"08",X"00",X"0F",
		X"00",X"00",X"04",X"04",X"08",X"08",X"08",X"04",X"02",X"00",X"04",X"5F",X"9F",X"2D",X"1E",X"7E",
		X"09",X"10",X"32",X"66",X"45",X"00",X"00",X"00",X"01",X"02",X"02",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"01",X"00",X"10",X"C9",X"0C",X"00",X"00",X"87",X"C4",X"44",X"BC",X"06",X"01",X"00",X"00",
		X"0F",X"0F",X"EF",X"E3",X"34",X"07",X"00",X"00",X"8F",X"09",X"00",X"00",X"09",X"06",X"00",X"00",
		X"02",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"6C",X"24",X"28",X"C9",X"0E",X"00",X"08",X"00",
		X"00",X"00",X"00",X"00",X"38",X"70",X"F0",X"F0",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"08",X"00",X"80",X"80",X"00",X"08",X"08",X"08",X"68",X"E1",X"F2",X"F3",
		X"F0",X"F0",X"F0",X"71",X"38",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"01",X"00",X"00",
		X"0F",X"88",X"80",X"00",X"08",X"04",X"00",X"00",X"F3",X"F7",X"FF",X"FE",X"E0",X"08",X"08",X"08",
		X"00",X"00",X"00",X"03",X"07",X"4F",X"3C",X"4B",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"00",X"00",X"00",X"00",X"0E",X"2C",X"0E",X"48",X"00",X"00",X"00",X"08",X"3C",X"2D",X"0F",X"0F",
		X"F3",X"79",X"F1",X"F1",X"F4",X"74",X"00",X"00",X"03",X"07",X"34",X"10",X"00",X"00",X"00",X"00",
		X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"0F",X"1F",X"F1",X"F2",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"12",X"34",X"34",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"C0",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"03",X"B6",X"8F",X"1F",X"3C",
		X"4F",X"9F",X"F0",X"F0",X"A0",X"00",X"00",X"00",X"01",X"03",X"03",X"12",X"10",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"F8",X"E0",X"E0",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"07",X"0F",X"0F",X"0F",X"1F",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"01",
		X"00",X"00",X"00",X"00",X"08",X"4C",X"CC",X"88",X"00",X"00",X"00",X"00",X"0B",X"87",X"C3",X"D2",
		X"FF",X"F6",X"3C",X"3C",X"3F",X"77",X"00",X"00",X"17",X"07",X"17",X"33",X"00",X"00",X"00",X"00",
		X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D6",X"FC",X"E8",X"C8",X"88",X"00",X"00",X"00",
		X"07",X"0F",X"0F",X"06",X"0F",X"1F",X"6F",X"8F",X"00",X"01",X"03",X"06",X"07",X"0F",X"0F",X"FF",
		X"8F",X"6F",X"1F",X"0F",X"06",X"0F",X"0F",X"07",X"FF",X"0F",X"0F",X"87",X"86",X"83",X"01",X"00",
		X"FF",X"E1",X"E1",X"D2",X"52",X"1C",X"08",X"00",X"F1",X"E7",X"8F",X"3C",X"24",X"78",X"C3",X"0E",
		X"30",X"78",X"3C",X"16",X"1E",X"0F",X"0F",X"FF",X"0E",X"0F",X"0F",X"06",X"0F",X"8F",X"6F",X"1F",
		X"FF",X"E1",X"E1",X"C2",X"42",X"0C",X"08",X"00",X"F1",X"E7",X"8F",X"3C",X"24",X"78",X"C3",X"0E",
		X"FF",X"E1",X"E1",X"D2",X"52",X"3C",X"78",X"30",X"F1",X"E7",X"8F",X"3C",X"24",X"78",X"C3",X"0E",
		X"00",X"10",X"12",X"16",X"1E",X"1E",X"2D",X"4A",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"0F",
		X"84",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"1E",X"2D",X"4A",X"84",X"00",X"00",X"00",X"00",
		X"30",X"13",X"13",X"13",X"13",X"13",X"13",X"27",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"2D",X"5B",X"D3",X"5B",X"13",X"00",X"80",X"87",X"87",X"E1",X"3C",X"01",X"00",
		X"EF",X"8F",X"06",X"8F",X"8F",X"09",X"0F",X"0F",X"13",X"37",X"6E",X"FF",X"FF",X"99",X"FF",X"FF",
		X"13",X"5B",X"5B",X"D3",X"2D",X"00",X"00",X"00",X"00",X"01",X"0F",X"0F",X"F0",X"87",X"80",X"00",
		X"0F",X"0F",X"09",X"CF",X"CF",X"46",X"EF",X"FC",X"FF",X"FF",X"99",X"FF",X"FF",X"6E",X"37",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"00",X"00",X"00",X"00",X"0C",X"0E",X"0F",X"87",
		X"07",X"30",X"13",X"13",X"13",X"13",X"13",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"0F",X"96",X"5A",X"34",X"12",X"10",X"00",X"4B",X"34",X"03",X"00",X"00",X"00",X"00",X"00",
		X"8F",X"6F",X"1F",X"0F",X"06",X"0F",X"0F",X"87",X"FF",X"0F",X"0F",X"07",X"06",X"43",X"69",X"78",
		X"8F",X"6F",X"1F",X"0F",X"06",X"0F",X"0F",X"87",X"FF",X"0F",X"0F",X"07",X"06",X"03",X"01",X"30",
		X"FF",X"E1",X"E1",X"C2",X"42",X"0C",X"08",X"C0",X"F1",X"E7",X"8F",X"3C",X"24",X"78",X"C3",X"1E",
		X"FF",X"E1",X"E1",X"C2",X"42",X"2C",X"69",X"C3",X"F1",X"E7",X"8F",X"3C",X"24",X"78",X"C3",X"1E",
		X"01",X"03",X"07",X"07",X"0F",X"1E",X"2D",X"4A",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A7",X"2F",X"4E",X"8C",X"8C",X"08",X"00",X"00",
		X"84",X"84",X"84",X"4A",X"4A",X"E0",X"3F",X"6F",X"71",X"03",X"03",X"03",X"01",X"10",X"10",X"01",
		X"00",X"00",X"00",X"00",X"00",X"01",X"2D",X"ED",X"00",X"00",X"00",X"00",X"00",X"00",X"87",X"F7",
		X"FF",X"FF",X"77",X"3F",X"0F",X"07",X"0F",X"0F",X"33",X"17",X"0E",X"0F",X"0F",X"0E",X"0F",X"0F",
		X"84",X"86",X"43",X"E1",X"E1",X"81",X"E1",X"E1",X"FC",X"FC",X"EC",X"FE",X"1E",X"19",X"0F",X"0F",
		X"0E",X"0F",X"87",X"4B",X"25",X"25",X"12",X"01",X"70",X"12",X"01",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"0F",X"E0",X"4A",X"4A",X"84",X"84",X"8C",X"11",X"10",X"10",X"01",X"03",X"03",X"03",X"70",
		X"00",X"10",X"12",X"16",X"3E",X"7E",X"ED",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",
		X"CC",X"FF",X"7F",X"0F",X"07",X"0F",X"0F",X"07",X"3F",X"1F",X"0F",X"87",X"86",X"83",X"01",X"00",
		X"CD",X"69",X"E1",X"D2",X"52",X"1C",X"08",X"00",X"11",X"FF",X"FF",X"FE",X"EC",X"BC",X"0F",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"0E",X"EF",X"00",X"80",X"84",X"86",X"87",X"87",X"4B",X"25",
		X"EE",X"6E",X"04",X"00",X"00",X"00",X"00",X"00",X"12",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"4C",X"EE",X"66",X"6E",X"CC",X"EE",X"FF",X"00",X"01",X"03",X"06",X"07",X"0F",X"3F",X"F1",
		X"FF",X"7F",X"3F",X"3F",X"07",X"0F",X"0F",X"07",X"F1",X"0F",X"0F",X"07",X"06",X"03",X"01",X"00",
		X"00",X"21",X"E9",X"CA",X"C2",X"0C",X"08",X"00",X"00",X"CC",X"CC",X"FF",X"7F",X"78",X"C3",X"0E",
		X"00",X"08",X"0C",X"0E",X"8E",X"8F",X"8F",X"C3",X"06",X"07",X"03",X"33",X"11",X"11",X"77",X"77",
		X"00",X"CC",X"EE",X"CE",X"CA",X"0C",X"08",X"00",X"88",X"DD",X"FF",X"FE",X"FC",X"FC",X"CB",X"0E",
		X"FE",X"E1",X"E1",X"C2",X"42",X"0C",X"08",X"C0",X"FF",X"FF",X"CF",X"BC",X"AC",X"78",X"C3",X"1E",
		X"FF",X"FF",X"3F",X"1F",X"17",X"0F",X"0F",X"87",X"F7",X"0F",X"0F",X"07",X"06",X"03",X"01",X"30",
		X"01",X"13",X"17",X"17",X"0F",X"1E",X"2D",X"4A",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"CE",X"84",X"84",X"08",X"00",X"00",
		X"84",X"08",X"0C",X"06",X"0E",X"0F",X"8F",X"FE",X"1E",X"07",X"8F",X"8E",X"EF",X"77",X"77",X"77",
		X"CF",X"E1",X"E1",X"C2",X"42",X"0C",X"08",X"C0",X"77",X"67",X"EF",X"FC",X"EC",X"F8",X"C3",X"1E",
		X"0F",X"CE",X"E6",X"6A",X"04",X"00",X"00",X"00",X"70",X"12",X"01",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"08",X"0C",X"06",X"0E",X"0F",X"0F",X"FE",X"1E",X"0F",X"0F",X"8E",X"8F",X"CF",X"FF",X"FF",
		X"E1",X"E9",X"CB",X"CA",X"86",X"84",X"08",X"00",X"77",X"77",X"11",X"11",X"33",X"30",X"61",X"06",
		X"EF",X"E5",X"E1",X"D2",X"52",X"1C",X"08",X"00",X"FF",X"EF",X"CF",X"FC",X"2C",X"78",X"C3",X"0E",
		X"F0",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"F0",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"F0",X"EF",X"EF",X"EF",X"EF",X"EF",X"00",X"00",X"F0",X"1F",X"1F",X"1F",X"1F",X"1F",X"00",X"00",
		X"F0",X"EF",X"EF",X"00",X"00",X"00",X"00",X"00",X"F0",X"1F",X"1F",X"00",X"00",X"00",X"00",X"00",
		X"3C",X"3D",X"79",X"F3",X"F3",X"79",X"3D",X"3C",X"00",X"00",X"03",X"1E",X"1E",X"03",X"00",X"00",
		X"F0",X"0F",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"0F",X"0F",X"FF",X"FF",X"33",X"00",X"00",
		X"F0",X"E1",X"E1",X"FF",X"FF",X"CC",X"00",X"00",X"F0",X"1E",X"1E",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"FF",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",
		X"F0",X"E1",X"E1",X"E1",X"E1",X"E1",X"00",X"00",X"F0",X"1E",X"1E",X"1E",X"1E",X"1E",X"FF",X"FF",
		X"1E",X"1E",X"1E",X"FE",X"FE",X"FE",X"FE",X"1E",X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",X"FF",X"0F",
		X"1E",X"1E",X"1E",X"FE",X"FE",X"FE",X"FE",X"1E",X"03",X"03",X"03",X"33",X"33",X"33",X"33",X"03",
		X"16",X"16",X"16",X"76",X"76",X"76",X"76",X"16",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"08",X"0C",X"84",X"87",X"C3",X"F8",X"FE",X"01",X"01",X"03",X"12",X"1E",X"3C",X"F1",X"F7",
		X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"11",X"11",X"33",X"33",X"FF",X"FF",X"FF",X"FF",
		X"9E",X"9E",X"9E",X"F8",X"F8",X"F8",X"F8",X"9E",X"FF",X"FF",X"FF",X"FF",X"33",X"33",X"11",X"11",
		X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"03",X"03",X"03",X"03",X"CF",X"CF",X"CF",X"CF",
		X"1E",X"1E",X"1E",X"F0",X"F0",X"F0",X"F0",X"1E",X"CF",X"CF",X"CF",X"FC",X"30",X"30",X"30",X"03");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
