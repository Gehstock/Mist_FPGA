library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ps04 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ps04 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"18",X"11",X"31",X"45",X"2A",X"29",X"20",X"E5",X"D5",X"FF",X"3E",X"04",X"11",X"01",X"07",X"DF",
		X"D1",X"E1",X"01",X"01",X"18",X"C3",X"AB",X"07",X"2A",X"29",X"20",X"E5",X"01",X"01",X"18",X"CD",
		X"0F",X"09",X"E1",X"FF",X"3E",X"03",X"11",X"01",X"07",X"DF",X"21",X"00",X"00",X"22",X"27",X"20",
		X"21",X"01",X"01",X"22",X"3A",X"20",X"C3",X"6A",X"18",X"21",X"33",X"20",X"AF",X"BE",X"C8",X"23",
		X"34",X"7E",X"E6",X"04",X"C2",X"55",X"18",X"2A",X"35",X"20",X"CD",X"70",X"18",X"11",X"FA",X"45",
		X"06",X"08",X"C3",X"E9",X"03",X"2A",X"35",X"20",X"CD",X"7A",X"18",X"01",X"01",X"08",X"CD",X"0F",
		X"09",X"21",X"00",X"00",X"22",X"33",X"20",X"22",X"35",X"20",X"21",X"0A",X"20",X"36",X"00",X"C9",
		X"E5",X"FF",X"3E",X"06",X"11",X"02",X"03",X"DF",X"E1",X"C9",X"7D",X"FE",X"74",X"3E",X"02",X"D2",
		X"84",X"18",X"3E",X"07",X"E5",X"F5",X"FF",X"F1",X"11",X"02",X"03",X"DF",X"E1",X"C9",X"21",X"2F",
		X"20",X"AF",X"BE",X"C8",X"23",X"34",X"7E",X"E6",X"04",X"C2",X"B1",X"18",X"2A",X"31",X"20",X"E5",
		X"FF",X"3E",X"02",X"11",X"01",X"07",X"DF",X"E1",X"11",X"02",X"46",X"01",X"01",X"18",X"C3",X"AB",
		X"07",X"2A",X"31",X"20",X"3A",X"43",X"20",X"A7",X"C2",X"C3",X"18",X"22",X"46",X"20",X"3E",X"01",
		X"32",X"42",X"20",X"01",X"01",X"18",X"CD",X"0F",X"09",X"21",X"00",X"00",X"22",X"2F",X"20",X"22",
		X"31",X"20",X"C3",X"6A",X"18",X"21",X"0B",X"23",X"AF",X"BE",X"C8",X"21",X"14",X"20",X"34",X"7E",
		X"E6",X"0F",X"C0",X"2E",X"0A",X"AF",X"BE",X"C0",X"2E",X"0D",X"36",X"01",X"C9",X"21",X"05",X"00",
		X"3A",X"0D",X"23",X"A7",X"C8",X"22",X"12",X"23",X"21",X"11",X"23",X"34",X"C3",X"09",X"03",X"21",
		X"38",X"20",X"AF",X"BE",X"C8",X"36",X"00",X"21",X"00",X"00",X"22",X"0D",X"20",X"22",X"0E",X"20",
		X"11",X"B4",X"42",X"2A",X"12",X"20",X"CD",X"ED",X"08",X"21",X"0A",X"20",X"34",X"E7",X"2E",X"00",
		X"AF",X"BE",X"CA",X"75",X"19",X"23",X"0E",X"05",X"22",X"48",X"20",X"AF",X"BE",X"CA",X"36",X"19",
		X"CD",X"58",X"1C",X"D4",X"3F",X"19",X"CD",X"60",X"1C",X"C2",X"2B",X"19",X"C3",X"75",X"19",X"CD",
		X"6B",X"1C",X"D0",X"3A",X"13",X"20",X"23",X"BE",X"D8",X"F5",X"3E",X"20",X"86",X"47",X"F1",X"B8",
		X"D0",X"2B",X"F1",X"E5",X"2E",X"4B",X"34",X"E1",X"2B",X"36",X"00",X"CD",X"09",X"0B",X"22",X"2D",
		X"20",X"01",X"01",X"18",X"CD",X"0F",X"09",X"21",X"2B",X"20",X"34",X"2E",X"F4",X"36",X"15",X"CD",
		X"91",X"1F",X"C3",X"ED",X"18",X"E7",X"2E",X"13",X"AF",X"BE",X"CA",X"B2",X"19",X"23",X"0E",X"05",
		X"22",X"48",X"20",X"AF",X"BE",X"CA",X"8E",X"19",X"CD",X"58",X"1C",X"D4",X"97",X"19",X"CD",X"60",
		X"1C",X"C2",X"83",X"19",X"C3",X"B2",X"19",X"CD",X"6B",X"1C",X"D0",X"3A",X"13",X"20",X"23",X"BE",
		X"D8",X"F5",X"3E",X"20",X"86",X"47",X"F1",X"B8",X"D0",X"2B",X"C1",X"E5",X"2E",X"4C",X"34",X"C3",
		X"57",X"19",X"E7",X"2E",X"39",X"AF",X"BE",X"CA",X"05",X"1A",X"23",X"0E",X"05",X"22",X"48",X"20",
		X"AF",X"BE",X"CA",X"CB",X"19",X"CD",X"58",X"1C",X"D4",X"D4",X"19",X"CD",X"60",X"1C",X"C2",X"C0",
		X"19",X"C3",X"05",X"1A",X"CD",X"6B",X"1C",X"D0",X"3A",X"13",X"20",X"23",X"BE",X"D8",X"F5",X"3E",
		X"14",X"86",X"47",X"F1",X"B8",X"D0",X"2B",X"D1",X"E5",X"2E",X"4A",X"34",X"E1",X"2B",X"36",X"00",
		X"CD",X"09",X"0B",X"22",X"29",X"20",X"01",X"01",X"18",X"CD",X"0F",X"09",X"21",X"27",X"20",X"34",
		X"2E",X"F2",X"36",X"15",X"C9",X"21",X"51",X"20",X"AF",X"BE",X"CA",X"47",X"1A",X"21",X"56",X"20",
		X"CD",X"5B",X"1A",X"D4",X"19",X"1A",X"C3",X"47",X"1A",X"CD",X"64",X"1A",X"D0",X"23",X"7E",X"D6",
		X"08",X"47",X"3A",X"13",X"20",X"B8",X"D8",X"F5",X"3E",X"18",X"86",X"47",X"F1",X"B8",X"D0",X"E1",
		X"2A",X"56",X"20",X"22",X"31",X"20",X"21",X"2F",X"20",X"34",X"2E",X"F5",X"36",X"10",X"21",X"10",
		X"00",X"CD",X"F0",X"18",X"C3",X"24",X"0E",X"21",X"74",X"20",X"AF",X"BE",X"CA",X"B6",X"1A",X"21",
		X"77",X"20",X"CD",X"5B",X"1A",X"D4",X"7C",X"1A",X"C3",X"B6",X"1A",X"7E",X"D6",X"08",X"47",X"3A",
		X"12",X"20",X"B8",X"C9",X"F5",X"3E",X"08",X"C3",X"77",X"1A",X"23",X"7E",X"D6",X"03",X"47",X"3A",
		X"13",X"20",X"B8",X"C9",X"F5",X"3E",X"04",X"86",X"47",X"F1",X"B8",X"C9",X"CD",X"64",X"1A",X"D0",
		X"CD",X"6A",X"1A",X"D8",X"CD",X"74",X"1A",X"D0",X"D1",X"2A",X"77",X"20",X"CD",X"AB",X"1A",X"CD",
		X"15",X"10",X"E7",X"2E",X"4B",X"7E",X"FE",X"06",X"DA",X"A0",X"1A",X"21",X"72",X"20",X"36",X"00",
		X"21",X"F6",X"20",X"36",X"0A",X"21",X"03",X"00",X"C3",X"F0",X"18",X"22",X"35",X"20",X"3E",X"01",
		X"32",X"33",X"20",X"C3",X"6B",X"10",X"21",X"7D",X"20",X"AF",X"BE",X"CA",X"F1",X"1A",X"21",X"80",
		X"20",X"CD",X"5B",X"1A",X"D4",X"CA",X"1A",X"C3",X"F1",X"1A",X"CD",X"64",X"1A",X"D0",X"CD",X"6A",
		X"1A",X"D8",X"CD",X"74",X"1A",X"D0",X"C1",X"2A",X"80",X"20",X"CD",X"AB",X"1A",X"CD",X"A9",X"10",
		X"E7",X"2E",X"4B",X"7E",X"FE",X"06",X"DA",X"A0",X"1A",X"21",X"7B",X"20",X"36",X"00",X"C3",X"A0",
		X"1A",X"21",X"86",X"20",X"AF",X"BE",X"CA",X"2C",X"1B",X"21",X"89",X"20",X"CD",X"5B",X"1A",X"D4",
		X"05",X"1B",X"C3",X"2C",X"1B",X"CD",X"64",X"1A",X"D0",X"CD",X"6A",X"1A",X"D8",X"CD",X"74",X"1A",
		X"D0",X"E1",X"2A",X"89",X"20",X"CD",X"AB",X"1A",X"CD",X"10",X"11",X"E7",X"2E",X"4C",X"7E",X"FE",
		X"06",X"DA",X"A0",X"1A",X"21",X"84",X"20",X"36",X"00",X"C3",X"A0",X"1A",X"21",X"8F",X"20",X"AF",
		X"BE",X"CA",X"67",X"1B",X"21",X"92",X"20",X"CD",X"5B",X"1A",X"D4",X"40",X"1B",X"C3",X"67",X"1B",
		X"CD",X"64",X"1A",X"D0",X"CD",X"6A",X"1A",X"D8",X"CD",X"74",X"1A",X"D0",X"F1",X"2A",X"92",X"20",
		X"CD",X"AB",X"1A",X"CD",X"77",X"11",X"E7",X"2E",X"4C",X"7E",X"FE",X"06",X"DA",X"A0",X"1A",X"21",
		X"8D",X"20",X"36",X"00",X"C3",X"A0",X"1A",X"21",X"AB",X"20",X"AF",X"BE",X"CA",X"A9",X"1B",X"21",
		X"AE",X"20",X"CD",X"5B",X"1A",X"D4",X"7B",X"1B",X"C3",X"A9",X"1B",X"CD",X"64",X"1A",X"D0",X"CD",
		X"6A",X"1A",X"D8",X"CD",X"74",X"1A",X"D0",X"D1",X"2A",X"AE",X"20",X"CD",X"A3",X"1B",X"21",X"A9",
		X"20",X"11",X"A9",X"40",X"06",X"07",X"CD",X"BB",X"04",X"21",X"23",X"20",X"34",X"21",X"01",X"00",
		X"C3",X"F0",X"18",X"22",X"25",X"20",X"C3",X"86",X"13",X"21",X"B2",X"20",X"AF",X"BE",X"CA",X"D9",
		X"1B",X"21",X"B5",X"20",X"CD",X"5B",X"1A",X"D4",X"BD",X"1B",X"C3",X"D9",X"1B",X"CD",X"64",X"1A",
		X"D0",X"CD",X"6A",X"1A",X"D8",X"CD",X"74",X"1A",X"D0",X"C1",X"2A",X"B5",X"20",X"CD",X"A3",X"1B",
		X"21",X"B0",X"20",X"11",X"B0",X"40",X"C3",X"94",X"1B",X"21",X"B9",X"20",X"AF",X"BE",X"CA",X"09",
		X"1C",X"21",X"BC",X"20",X"CD",X"5B",X"1A",X"D4",X"ED",X"1B",X"C3",X"09",X"1C",X"CD",X"64",X"1A",
		X"D0",X"CD",X"6A",X"1A",X"D8",X"CD",X"74",X"1A",X"D0",X"E1",X"2A",X"BC",X"20",X"CD",X"A3",X"1B",
		X"21",X"B7",X"20",X"11",X"B7",X"40",X"C3",X"94",X"1B",X"21",X"E5",X"20",X"AF",X"BE",X"CA",X"55",
		X"1C",X"21",X"EA",X"20",X"CD",X"5B",X"1A",X"D4",X"1D",X"1C",X"C3",X"55",X"1C",X"F5",X"3E",X"18",
		X"86",X"47",X"F1",X"B8",X"CD",X"6A",X"1A",X"D8",X"F5",X"3E",X"18",X"86",X"47",X"F1",X"B8",X"D0",
		X"C1",X"2A",X"EA",X"20",X"22",X"21",X"20",X"01",X"02",X"10",X"CD",X"0F",X"09",X"21",X"01",X"02",
		X"22",X"1F",X"20",X"21",X"F3",X"20",X"36",X"40",X"2E",X"E0",X"11",X"E0",X"40",X"06",X"10",X"CD",
		X"BB",X"04",X"C3",X"6A",X"18",X"C3",X"6A",X"18",X"23",X"3A",X"12",X"20",X"C6",X"08",X"BE",X"C9",
		X"2A",X"48",X"20",X"23",X"23",X"23",X"22",X"48",X"20",X"0D",X"C9",X"F5",X"3E",X"10",X"86",X"47",
		X"F1",X"B8",X"C9",X"21",X"42",X"20",X"97",X"BE",X"C8",X"23",X"BE",X"C2",X"98",X"1C",X"34",X"2A",
		X"46",X"20",X"01",X"00",X"08",X"09",X"22",X"46",X"20",X"3A",X"05",X"20",X"BD",X"21",X"FD",X"01",
		X"D2",X"95",X"1C",X"26",X"FF",X"22",X"44",X"20",X"2A",X"46",X"20",X"E5",X"CD",X"BC",X"0F",X"CD",
		X"F3",X"11",X"E1",X"7C",X"FE",X"F0",X"D2",X"BE",X"1C",X"FE",X"28",X"DA",X"BE",X"1C",X"7D",X"FE",
		X"30",X"DA",X"BE",X"1C",X"21",X"44",X"20",X"EF",X"2A",X"46",X"20",X"C3",X"E5",X"11",X"21",X"42",
		X"20",X"11",X"42",X"40",X"C3",X"1B",X"10",X"CD",X"18",X"1D",X"22",X"15",X"20",X"E7",X"2E",X"26",
		X"97",X"BE",X"C8",X"23",X"0E",X"03",X"C5",X"E5",X"AF",X"BE",X"CA",X"12",X"1D",X"CD",X"09",X"0B",
		X"22",X"17",X"20",X"CD",X"BC",X"0F",X"CD",X"F3",X"11",X"21",X"18",X"20",X"7E",X"FE",X"2B",X"DC",
		X"0A",X"1D",X"21",X"15",X"20",X"EF",X"2A",X"17",X"20",X"E5",X"CD",X"E5",X"11",X"E1",X"EB",X"E1",
		X"23",X"CD",X"15",X"0B",X"C1",X"0D",X"C2",X"D6",X"1C",X"C9",X"36",X"F0",X"C9",X"CD",X"09",X"0B",
		X"EB",X"C9",X"CD",X"0D",X"1D",X"C3",X"FF",X"1C",X"21",X"19",X"20",X"34",X"7E",X"21",X"FF",X"FE",
		X"E6",X"08",X"C8",X"21",X"01",X"FD",X"C9",X"CD",X"73",X"1D",X"22",X"1A",X"20",X"E7",X"2E",X"32",
		X"97",X"BE",X"C8",X"23",X"0E",X"02",X"C5",X"E5",X"AF",X"BE",X"CA",X"6A",X"1D",X"CD",X"09",X"0B",
		X"22",X"1C",X"20",X"CD",X"BC",X"0F",X"CD",X"F3",X"11",X"21",X"1D",X"20",X"7E",X"FE",X"E8",X"D4",
		X"70",X"1D",X"21",X"1A",X"20",X"EF",X"2A",X"1C",X"20",X"E5",X"CD",X"E5",X"11",X"E1",X"EB",X"E1",
		X"23",X"CD",X"15",X"0B",X"C1",X"0D",X"C2",X"36",X"1D",X"C9",X"CD",X"0D",X"1D",X"C3",X"5F",X"1D",
		X"36",X"28",X"C9",X"21",X"1E",X"20",X"34",X"7E",X"E6",X"08",X"21",X"01",X"03",X"C8",X"21",X"FF",
		X"02",X"C9",X"21",X"3B",X"20",X"97",X"BE",X"C8",X"2B",X"BE",X"CA",X"D2",X"1D",X"35",X"CD",X"4B",
		X"16",X"3A",X"39",X"20",X"E6",X"07",X"21",X"EF",X"1D",X"FE",X"00",X"CA",X"B1",X"1D",X"23",X"23",
		X"23",X"FE",X"01",X"CA",X"B1",X"1D",X"23",X"23",X"23",X"FE",X"02",X"CA",X"B1",X"1D",X"23",X"23",
		X"23",X"EB",X"1A",X"6F",X"26",X"00",X"13",X"D5",X"CD",X"F0",X"18",X"2A",X"29",X"20",X"F7",X"D1",
		X"CD",X"E4",X"02",X"3E",X"1C",X"CD",X"F2",X"02",X"21",X"F0",X"20",X"36",X"20",X"2E",X"00",X"36",
		X"00",X"C9",X"2A",X"29",X"20",X"06",X"18",X"CD",X"CA",X"03",X"2A",X"29",X"20",X"FF",X"3E",X"07",
		X"11",X"01",X"07",X"DF",X"21",X"00",X"00",X"22",X"3A",X"20",X"21",X"00",X"20",X"34",X"C9",X"50",
		X"21",X"1C",X"70",X"23",X"1C",X"90",X"25",X"1C",X"30",X"1F",X"1C",X"21",X"E3",X"20",X"97",X"BE",
		X"C8",X"23",X"BE",X"C2",X"20",X"10",X"23",X"BE",X"C2",X"27",X"1E",X"34",X"CD",X"D0",X"1E",X"22",
		X"EA",X"20",X"CD",X"EA",X"1E",X"22",X"E0",X"20",X"EB",X"1A",X"21",X"E6",X"20",X"77",X"23",X"13",
		X"1A",X"77",X"13",X"EB",X"22",X"E0",X"20",X"21",X"E6",X"20",X"AF",X"BE",X"CA",X"90",X"1E",X"35",
		X"3A",X"E7",X"20",X"21",X"9A",X"47",X"A7",X"CA",X"42",X"1E",X"01",X"02",X"00",X"09",X"3D",X"C2",
		X"3A",X"1E",X"5E",X"23",X"56",X"EB",X"22",X"E8",X"20",X"21",X"1A",X"46",X"3A",X"E7",X"20",X"A7",
		X"CA",X"5B",X"1E",X"11",X"20",X"00",X"19",X"3D",X"C2",X"53",X"1E",X"22",X"EC",X"20",X"21",X"EA",
		X"20",X"CD",X"C4",X"04",X"CD",X"56",X"05",X"21",X"EA",X"20",X"7E",X"FE",X"88",X"DA",X"B2",X"1E",
		X"23",X"7E",X"FE",X"28",X"DA",X"B2",X"1E",X"FE",X"E8",X"D2",X"B2",X"1E",X"21",X"E8",X"20",X"EF",
		X"2A",X"EA",X"20",X"FF",X"11",X"03",X"05",X"3E",X"05",X"DF",X"21",X"EA",X"20",X"C3",X"83",X"05",
		X"2A",X"E0",X"20",X"7E",X"FE",X"FF",X"CA",X"30",X"1E",X"E5",X"21",X"EA",X"20",X"CD",X"C4",X"04",
		X"CD",X"56",X"05",X"E1",X"5E",X"23",X"56",X"23",X"22",X"E0",X"20",X"EB",X"22",X"E6",X"20",X"C3",
		X"30",X"1E",X"21",X"E2",X"20",X"AF",X"BE",X"CA",X"C5",X"1E",X"35",X"23",X"23",X"11",X"E4",X"40",
		X"06",X"0C",X"C3",X"BB",X"04",X"11",X"E2",X"40",X"06",X"0E",X"CD",X"BB",X"04",X"C3",X"91",X"1F",
		X"3A",X"0F",X"23",X"E6",X"03",X"A7",X"21",X"E0",X"88",X"C8",X"FE",X"01",X"21",X"B0",X"E0",X"C8",
		X"FE",X"02",X"21",X"D0",X"30",X"C8",X"21",X"E0",X"C0",X"C9",X"3A",X"0F",X"23",X"E6",X"03",X"A7",
		X"21",X"B2",X"47",X"C8",X"FE",X"01",X"21",X"E5",X"47",X"C8",X"FE",X"02",X"21",X"1A",X"48",X"C8",
		X"21",X"59",X"48",X"C9",X"21",X"1F",X"20",X"97",X"BE",X"C8",X"23",X"BE",X"CA",X"82",X"1F",X"35",
		X"7E",X"FE",X"01",X"C2",X"3C",X"1F",X"2A",X"21",X"20",X"7C",X"FE",X"D8",X"DA",X"21",X"1F",X"26",
		X"D0",X"22",X"21",X"20",X"E5",X"FF",X"11",X"05",X"09",X"3E",X"06",X"DF",X"E1",X"11",X"0C",X"49",
		X"01",X"04",X"1E",X"CD",X"AB",X"07",X"21",X"F0",X"20",X"36",X"20",X"C9",X"2A",X"21",X"20",X"01",
		X"04",X"1E",X"E5",X"CD",X"0F",X"09",X"E1",X"F7",X"3A",X"39",X"20",X"E6",X"0F",X"A7",X"01",X"00",
		X"02",X"11",X"08",X"49",X"CA",X"73",X"1F",X"FE",X"01",X"01",X"50",X"01",X"11",X"04",X"49",X"CA",
		X"73",X"1F",X"FE",X"02",X"01",X"00",X"01",X"11",X"00",X"49",X"CA",X"73",X"1F",X"01",X"50",X"00",
		X"11",X"FC",X"48",X"C5",X"0E",X"04",X"CD",X"E6",X"02",X"C1",X"69",X"60",X"CD",X"F0",X"18",X"C3",
		X"36",X"1F",X"2A",X"21",X"20",X"01",X"01",X"20",X"CD",X"CA",X"03",X"21",X"00",X"00",X"22",X"1F",
		X"20",X"E7",X"2E",X"4D",X"34",X"C9",X"3A",X"0A",X"23",X"E6",X"0F",X"21",X"01",X"3D",X"C6",X"1C",
		X"CD",X"F2",X"02",X"3A",X"0A",X"23",X"E6",X"F0",X"0F",X"0F",X"0F",X"0F",X"21",X"01",X"3C",X"C6",
		X"1C",X"C3",X"F2",X"02",X"ED",X"18",X"02",X"00",X"4F",X"C4",X"B0",X"9A",X"48",X"16",X"02",X"00",
		X"5B",X"C4",X"F0",X"C8",X"51",X"09",X"02",X"00",X"5B",X"C4",X"40",X"D3",X"2E",X"09",X"02",X"00",
		X"5F",X"C4",X"F0",X"C8",X"47",X"09",X"02",X"00",X"5F",X"C4",X"60",X"CC",X"3D",X"09",X"02",X"00",
		X"80",X"C4",X"28",X"AF",X"BC",X"00",X"02",X"00",X"80",X"C4",X"50",X"AF",X"D7",X"00",X"02",X"00",
		X"80",X"C4",X"78",X"AF",X"DA",X"00",X"02",X"00",X"80",X"C4",X"A0",X"AF",X"B9",X"01",X"02",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
