library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_OBJ_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_OBJ_1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"7C",X"C6",X"C6",X"82",X"C6",X"C6",X"7C",X"00",X"00",X"06",X"FE",X"FE",X"86",X"00",X"00",
		X"00",X"66",X"F2",X"BA",X"9E",X"8E",X"C6",X"62",X"00",X"7C",X"FE",X"92",X"92",X"92",X"C6",X"44",
		X"00",X"18",X"FE",X"1E",X"1A",X"D8",X"F8",X"F8",X"00",X"9C",X"BE",X"B2",X"B2",X"B2",X"F6",X"F6",
		X"00",X"4C",X"DE",X"92",X"92",X"92",X"FE",X"7C",X"00",X"E0",X"F0",X"98",X"8E",X"86",X"C2",X"E0",
		X"00",X"6C",X"FE",X"92",X"92",X"92",X"FE",X"6C",X"00",X"7C",X"FE",X"92",X"92",X"92",X"F6",X"64",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"14",X"40",X"25",X"A4",X"25",X"98",X"02",X"28",
		X"3E",X"7F",X"F8",X"F8",X"F8",X"C0",X"C1",X"43",X"00",X"00",X"04",X"18",X"18",X"00",X"80",X"C0",
		X"03",X"01",X"00",X"18",X"18",X"20",X"00",X"00",X"C0",X"80",X"00",X"18",X"18",X"04",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7E",X"D6",X"D0",X"D0",X"D0",X"D6",X"7E",
		X"00",X"44",X"EE",X"BA",X"92",X"82",X"FE",X"FE",X"00",X"44",X"C6",X"82",X"82",X"82",X"FE",X"7C",
		X"00",X"7C",X"FE",X"82",X"82",X"BA",X"FE",X"FE",X"00",X"C6",X"C6",X"92",X"92",X"92",X"FE",X"FE",
		X"00",X"C0",X"C0",X"90",X"92",X"96",X"FE",X"FE",X"00",X"6C",X"EE",X"8A",X"8A",X"82",X"FE",X"7C",
		X"00",X"FE",X"FE",X"D0",X"10",X"16",X"FE",X"FE",X"00",X"00",X"C6",X"FE",X"FE",X"FE",X"C6",X"00",
		X"00",X"FC",X"FE",X"C2",X"06",X"0E",X"0C",X"08",X"00",X"82",X"C6",X"EE",X"38",X"92",X"FE",X"FE",
		X"00",X"1E",X"0E",X"06",X"02",X"E2",X"FE",X"FE",X"00",X"FE",X"C6",X"60",X"30",X"60",X"C6",X"FE",
		X"00",X"FE",X"CE",X"9C",X"38",X"72",X"E6",X"FE",X"00",X"7C",X"EE",X"C6",X"C6",X"C6",X"EE",X"7C",
		X"00",X"60",X"F0",X"90",X"90",X"92",X"FE",X"FE",X"00",X"06",X"7E",X"F6",X"CE",X"C6",X"DE",X"7C",
		X"00",X"62",X"F6",X"9E",X"90",X"96",X"FE",X"FE",X"00",X"C4",X"8E",X"9A",X"9A",X"B2",X"F2",X"66",
		X"00",X"F0",X"C2",X"FE",X"FE",X"FE",X"C2",X"F0",X"00",X"FC",X"FE",X"FA",X"02",X"02",X"FE",X"FC",
		X"00",X"C0",X"F8",X"FC",X"0E",X"FC",X"F8",X"C0",X"00",X"FE",X"C6",X"0C",X"18",X"0C",X"C6",X"FE",
		X"00",X"C6",X"C6",X"28",X"10",X"28",X"C6",X"C6",X"00",X"FE",X"FE",X"D2",X"12",X"16",X"F6",X"F6",
		X"00",X"CE",X"E2",X"F2",X"BA",X"9E",X"8E",X"E6",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"88",X"C8",X"30",X"38",X"1E",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",
		X"00",X"00",X"00",X"18",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"04",X"0C",X"00",X"00",
		X"00",X"00",X"18",X"24",X"28",X"18",X"00",X"00",X"00",X"00",X"18",X"0A",X"36",X"08",X"0C",X"00",
		X"00",X"78",X"C8",X"8C",X"A4",X"C8",X"38",X"00",X"38",X"04",X"BC",X"78",X"86",X"64",X"38",X"00",
		X"00",X"A8",X"86",X"02",X"44",X"10",X"14",X"10",X"04",X"10",X"20",X"00",X"00",X"00",X"02",X"0C",
		X"02",X"08",X"10",X"00",X"00",X"00",X"01",X"06",X"05",X"08",X"00",X"00",X"00",X"01",X"00",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"22",X"22",X"22",X"22",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F1",X"11",X"1F",X"11",X"F1",X"11",X"1F",X"11",X"F1",X"11",X"1F",X"11",X"F1",X"11",X"00",X"00",
		X"F1",X"11",X"1F",X"11",X"00",X"00",X"00",X"00",X"F1",X"11",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"38",X"54",X"7C",X"54",X"38",X"81",X"83",X"F0",X"08",X"E4",X"12",X"C9",X"25",X"95",X"D5",
		X"AB",X"A9",X"A4",X"93",X"48",X"27",X"10",X"0F",X"D5",X"95",X"25",X"C9",X"12",X"E4",X"08",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"10",X"08",X"04",X"04",X"04",X"08",X"F0",X"E0",
		X"03",X"07",X"0F",X"07",X"00",X"00",X"00",X"00",X"C0",X"80",X"00",X"00",X"80",X"40",X"40",X"80",
		X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"00",X"00",X"00",X"3C",X"04",X"00",X"00",X"00",X"00",
		X"10",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"84",X"C4",X"64",X"34",X"18",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"04",X"00",X"00",X"00",X"00",
		X"11",X"30",X"04",X"0C",X"18",X"30",X"60",X"00",X"84",X"04",X"04",X"04",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"04",X"00",X"00",X"00",X"80",
		X"10",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"84",X"84",X"04",X"04",X"88",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"43",X"23",X"13",X"0B",X"07",X"03",X"03",X"00",X"FF",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"3C",X"7E",X"7E",X"7E",X"7E",X"00",X"00",X"00",X"00",X"7E",X"7E",X"7E",X"7E",X"3C",X"00",
		X"00",X"00",X"06",X"0E",X"1E",X"3E",X"3C",X"00",X"00",X"3C",X"3E",X"1E",X"0E",X"06",X"00",X"00",
		X"00",X"00",X"7E",X"7E",X"7E",X"7E",X"00",X"00",X"00",X"00",X"60",X"70",X"78",X"7C",X"3C",X"00",
		X"00",X"3C",X"7C",X"78",X"70",X"60",X"00",X"00",X"00",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"00",
		X"12",X"08",X"02",X"00",X"0A",X"00",X"34",X"0A",X"20",X"12",X"0C",X"00",X"48",X"55",X"52",X"94",
		X"44",X"92",X"08",X"14",X"52",X"04",X"0A",X"01",X"80",X"58",X"45",X"32",X"0C",X"60",X"94",X"00",
		X"04",X"48",X"30",X"04",X"38",X"00",X"04",X"18",X"00",X"60",X"14",X"08",X"00",X"18",X"24",X"04",
		X"A4",X"88",X"70",X"10",X"28",X"14",X"20",X"C0",X"18",X"04",X"40",X"34",X"08",X"10",X"64",X"08",
		X"00",X"00",X"44",X"28",X"20",X"10",X"10",X"08",X"00",X"00",X"94",X"44",X"22",X"40",X"20",X"10",
		X"00",X"00",X"48",X"48",X"89",X"15",X"11",X"08",X"00",X"00",X"42",X"84",X"0A",X"09",X"10",X"08",
		X"00",X"00",X"85",X"4A",X"52",X"42",X"00",X"00",X"00",X"00",X"05",X"92",X"62",X"11",X"00",X"00",
		X"10",X"90",X"60",X"24",X"28",X"44",X"00",X"00",X"20",X"10",X"14",X"08",X"6A",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"3C",X"60",X"C0",
		X"01",X"03",X"07",X"0E",X"0E",X"14",X"08",X"00",X"C0",X"80",X"80",X"40",X"20",X"20",X"00",X"00",
		X"FF",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CA",X"90",X"A0",X"C0",X"80",X"80",X"80",X"00",
		X"32",X"62",X"92",X"82",X"82",X"82",X"92",X"A2",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"CF",X"CF",X"CE",X"CC",X"C8",X"00",X"00",X"80",
		X"8B",X"FB",X"FB",X"88",X"8B",X"8B",X"FB",X"FB",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",
		X"8B",X"BB",X"88",X"FB",X"7B",X"1B",X"0B",X"03",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"84",X"C8",X"D0",X"C0",X"C8",X"CC",X"CE",
		X"00",X"00",X"1B",X"3B",X"F8",X"FB",X"8B",X"BB",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"10",X"00",X"00",X"02",X"00",X"20",X"08",
		X"08",X"00",X"10",X"01",X"00",X"08",X"00",X"40",X"00",X"82",X"00",X"00",X"10",X"42",X"00",X"08",
		X"00",X"00",X"08",X"00",X"40",X"01",X"20",X"00",X"20",X"04",X"00",X"00",X"08",X"20",X"02",X"00",
		X"10",X"80",X"00",X"00",X"08",X"00",X"80",X"00",X"08",X"04",X"08",X"10",X"10",X"08",X"04",X"08",
		X"00",X"04",X"00",X"00",X"80",X"04",X"20",X"00",X"20",X"04",X"00",X"00",X"80",X"00",X"00",X"04",
		X"02",X"00",X"48",X"00",X"01",X"10",X"04",X"80",X"20",X"00",X"00",X"00",X"00",X"04",X"00",X"10",
		X"08",X"40",X"00",X"04",X"00",X"80",X"00",X"00",X"00",X"10",X"80",X"02",X"00",X"20",X"08",X"00",
		X"00",X"04",X"40",X"00",X"80",X"00",X"02",X"00",X"04",X"20",X"80",X"02",X"00",X"08",X"00",X"00",
		X"00",X"00",X"00",X"20",X"01",X"00",X"48",X"00",X"00",X"00",X"41",X"00",X"00",X"08",X"42",X"00",
		X"00",X"00",X"00",X"00",X"01",X"40",X"04",X"10",X"00",X"00",X"00",X"00",X"12",X"00",X"00",X"10",
		X"00",X"1F",X"20",X"5C",X"B0",X"B8",X"BC",X"80",X"00",X"F0",X"08",X"04",X"04",X"04",X"84",X"24",
		X"80",X"B0",X"B8",X"BC",X"5C",X"20",X"1F",X"00",X"04",X"84",X"24",X"04",X"04",X"08",X"F0",X"00",
		X"00",X"1F",X"20",X"5C",X"A4",X"AC",X"BC",X"80",X"00",X"F0",X"08",X"04",X"04",X"04",X"04",X"04",
		X"80",X"A4",X"AC",X"BC",X"5C",X"20",X"1F",X"00",X"04",X"04",X"04",X"04",X"04",X"08",X"F0",X"00",
		X"00",X"1F",X"20",X"5C",X"BC",X"AC",X"A4",X"80",X"00",X"F0",X"08",X"04",X"04",X"04",X"04",X"04",
		X"80",X"BC",X"AC",X"A4",X"5C",X"20",X"1F",X"00",X"04",X"04",X"04",X"04",X"04",X"08",X"F0",X"00",
		X"00",X"03",X"07",X"0F",X"1F",X"1F",X"3F",X"3F",X"00",X"C0",X"E0",X"F0",X"F8",X"F8",X"FC",X"FC",
		X"3F",X"3F",X"1F",X"1F",X"0F",X"07",X"03",X"00",X"FC",X"FC",X"F8",X"F8",X"F0",X"E0",X"C0",X"00",
		X"00",X"18",X"34",X"04",X"04",X"04",X"03",X"00",X"00",X"60",X"90",X"90",X"90",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"04",X"03",X"00",X"00",X"60",X"90",X"90",X"90",X"92",X"0C",X"00",
		X"00",X"61",X"92",X"92",X"92",X"92",X"0C",X"00",X"00",X"06",X"09",X"09",X"09",X"01",X"00",X"00",
		X"00",X"18",X"2C",X"20",X"20",X"20",X"C0",X"00",X"00",X"06",X"09",X"09",X"09",X"49",X"30",X"00",
		X"00",X"00",X"00",X"00",X"30",X"20",X"C0",X"00",X"00",X"86",X"49",X"49",X"49",X"49",X"30",X"00",
		X"02",X"02",X"3C",X"40",X"60",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"40",X"40",X"3C",
		X"02",X"02",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"02",X"3C",X"40",X"40",X"3C",
		X"40",X"3C",X"02",X"02",X"3C",X"40",X"40",X"3C",X"3C",X"40",X"40",X"38",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"60",X"40",X"3C",X"02",X"02",X"3C",X"40",X"40",X"3C",X"02",X"02",X"04",X"00",
		X"00",X"00",X"00",X"00",X"08",X"0C",X"02",X"02",X"3C",X"40",X"40",X"3C",X"02",X"02",X"3C",X"40",
		X"3C",X"16",X"17",X"01",X"01",X"17",X"16",X"3C",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"07",X"02",X"05",X"07",X"00",X"00",X"00",X"00",X"80",X"F0",X"70",X"80",X"00",X"00",
		X"00",X"00",X"00",X"E2",X"FE",X"02",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",
		X"3C",X"68",X"E8",X"80",X"80",X"E8",X"68",X"3C",X"00",X"00",X"01",X"0F",X"0E",X"01",X"00",X"00",
		X"00",X"00",X"E0",X"40",X"A0",X"E0",X"00",X"00",X"00",X"00",X"00",X"4E",X"7F",X"40",X"00",X"00",
		X"3C",X"66",X"E7",X"81",X"E7",X"81",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",
		X"34",X"2C",X"34",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"18",X"18",X"2C",
		X"00",X"38",X"10",X"10",X"18",X"18",X"18",X"10",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"81",X"E7",X"81",X"E7",X"66",X"3C",X"2C",X"18",X"18",X"18",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"34",X"2C",X"34",X"10",X"18",X"18",X"18",X"10",X"10",X"38",X"00",
		X"00",X"00",X"06",X"3F",X"3E",X"07",X"00",X"00",X"00",X"00",X"A8",X"10",X"A0",X"58",X"00",X"00",
		X"00",X"00",X"01",X"07",X"07",X"01",X"00",X"00",X"08",X"54",X"EA",X"C0",X"C0",X"EA",X"54",X"08",
		X"2C",X"70",X"E6",X"F8",X"F8",X"E6",X"70",X"2C",X"00",X"00",X"1A",X"05",X"08",X"15",X"00",X"00",
		X"00",X"00",X"E0",X"7C",X"FC",X"60",X"00",X"00",X"10",X"2A",X"57",X"03",X"03",X"57",X"2A",X"10",
		X"00",X"00",X"80",X"E0",X"E0",X"80",X"00",X"00",X"34",X"0E",X"67",X"1F",X"1F",X"67",X"0E",X"34",
		X"28",X"3C",X"3C",X"18",X"18",X"18",X"00",X"00",X"00",X"00",X"00",X"24",X"28",X"14",X"20",X"14",
		X"3C",X"18",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"42",X"A5",X"42",X"24",X"7E",X"3C",
		X"00",X"24",X"A5",X"99",X"5A",X"FF",X"7E",X"3C",X"14",X"20",X"14",X"28",X"24",X"00",X"00",X"00",
		X"00",X"00",X"18",X"18",X"18",X"3C",X"3C",X"28",X"3C",X"7E",X"24",X"42",X"A5",X"42",X"24",X"00",
		X"00",X"00",X"00",X"00",X"00",X"18",X"18",X"3C",X"3C",X"7E",X"FF",X"5A",X"99",X"A5",X"24",X"00",
		X"1C",X"26",X"02",X"03",X"07",X"3E",X"1C",X"00",X"00",X"00",X"40",X"E0",X"20",X"00",X"00",X"00",
		X"00",X"07",X"08",X"00",X"0F",X"07",X"00",X"00",X"00",X"88",X"48",X"F8",X"90",X"10",X"00",X"00",
		X"00",X"01",X"73",X"FE",X"FE",X"73",X"01",X"00",X"00",X"00",X"00",X"04",X"07",X"02",X"00",X"00",
		X"00",X"38",X"7C",X"E0",X"C0",X"40",X"64",X"38",X"00",X"00",X"08",X"09",X"1F",X"13",X"11",X"00",
		X"00",X"00",X"E0",X"F0",X"80",X"10",X"E0",X"00",X"00",X"80",X"CE",X"7F",X"7F",X"CE",X"80",X"00",
		X"30",X"7C",X"E6",X"C2",X"C2",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"18",X"10",
		X"64",X"64",X"64",X"28",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"70",X"10",X"18",X"3C",
		X"E7",X"3C",X"18",X"18",X"3C",X"3C",X"3C",X"18",X"10",X"18",X"30",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"44",X"C2",X"C2",X"E6",X"7C",X"30",X"3C",X"18",X"10",X"70",X"1C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"28",X"64",X"64",X"74",X"18",X"3C",X"3C",X"3C",X"18",X"18",X"3C",X"66",
		X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"D0",X"90",X"90",X"E0",X"C0",X"C0",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",
		X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"C0",X"88",X"90",X"E0",X"C0",X"C0",
		X"01",X"02",X"02",X"04",X"00",X"00",X"00",X"00",X"80",X"40",X"40",X"20",X"00",X"00",X"00",X"00",
		X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"C0",X"88",X"88",X"F0",X"C0",X"C0",
		X"01",X"02",X"04",X"08",X"00",X"00",X"00",X"00",X"80",X"40",X"20",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"C0",
		X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"C0",X"C0",X"C0",X"E0",X"90",X"D0",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"02",X"02",X"01",X"00",X"00",X"00",X"00",X"20",X"40",X"40",X"80",
		X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"C0",X"C0",X"E0",X"90",X"88",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"04",X"02",X"01",X"00",X"00",X"00",X"00",X"10",X"20",X"40",X"80",
		X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"C0",X"C0",X"F0",X"88",X"88",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"FD",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"F4",X"10",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"FD",
		X"00",X"03",X"04",X"00",X"00",X"00",X"00",X"00",X"FE",X"64",X"10",X"08",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"04",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"FD",
		X"00",X"01",X"02",X"04",X"08",X"00",X"00",X"00",X"FE",X"64",X"20",X"20",X"18",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"BF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"7F",X"2F",X"08",X"70",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"BF",X"00",X"00",X"00",X"00",X"00",X"20",X"C0",X"00",
		X"7F",X"26",X"08",X"10",X"20",X"00",X"00",X"00",X"00",X"C0",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"BF",X"00",X"00",X"00",X"10",X"20",X"40",X"80",X"00",
		X"7F",X"26",X"04",X"04",X"18",X"00",X"00",X"00",X"00",X"80",X"40",X"20",X"10",X"00",X"00",X"00",
		X"00",X"01",X"00",X"2C",X"1C",X"1F",X"07",X"03",X"00",X"00",X"80",X"80",X"80",X"00",X"80",X"C0",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"30",X"10",X"08",X"00",X"00",X"00",
		X"00",X"02",X"01",X"2C",X"1C",X"1F",X"07",X"03",X"00",X"00",X"00",X"80",X"80",X"00",X"80",X"C0",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"80",X"40",X"40",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"2C",X"1C",X"1F",X"07",X"03",X"80",X"80",X"80",X"80",X"80",X"00",X"80",X"C0",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"80",X"80",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"08",X"10",X"30",X"E0",X"C0",
		X"03",X"07",X"1F",X"1C",X"2C",X"00",X"01",X"00",X"C0",X"80",X"00",X"80",X"80",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"20",X"40",X"40",X"80",X"B0",
		X"03",X"07",X"1F",X"1C",X"2C",X"01",X"02",X"00",X"C0",X"80",X"00",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"F8",
		X"03",X"07",X"1F",X"1C",X"2C",X"00",X"00",X"00",X"C0",X"80",X"00",X"80",X"80",X"80",X"80",X"80",
		X"00",X"00",X"00",X"10",X"0C",X"06",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"DC",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E2",X"E0",X"60",X"30",X"70",X"00",X"30",X"00",
		X"00",X"00",X"04",X"02",X"32",X"09",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"8C",X"D2",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E2",X"E0",X"60",X"30",X"70",X"00",X"30",X"00",
		X"00",X"00",X"00",X"01",X"01",X"11",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"F0",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E8",X"E4",X"60",X"30",X"70",X"00",X"30",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"30",X"00",X"70",X"30",X"60",X"E0",X"E2",
		X"03",X"07",X"07",X"0C",X"10",X"00",X"00",X"00",X"DC",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"30",X"00",X"70",X"30",X"60",X"E0",X"E2",
		X"03",X"07",X"09",X"32",X"02",X"04",X"00",X"00",X"D2",X"8C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"30",X"00",X"70",X"30",X"60",X"E4",X"E8",
		X"03",X"0F",X"11",X"01",X"01",X"00",X"00",X"00",X"F0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"03",X"01",X"01",X"01",X"03",X"07",X"3F",X"20",X"C0",X"80",X"80",X"80",X"80",X"C0",X"F0",
		X"1F",X"0F",X"07",X"05",X"05",X"07",X"03",X"01",X"E0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",
		X"02",X"03",X"01",X"01",X"01",X"03",X"07",X"1F",X"40",X"C0",X"80",X"80",X"80",X"80",X"C0",X"E0",
		X"0F",X"0F",X"07",X"05",X"05",X"07",X"03",X"01",X"E0",X"40",X"40",X"20",X"20",X"20",X"40",X"00",
		X"00",X"00",X"00",X"01",X"01",X"03",X"07",X"0F",X"00",X"00",X"00",X"80",X"80",X"80",X"C0",X"E0",
		X"0F",X"0F",X"07",X"05",X"05",X"07",X"03",X"01",X"C0",X"40",X"20",X"10",X"10",X"10",X"20",X"00",
		X"01",X"03",X"07",X"05",X"05",X"07",X"0F",X"1F",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"E0",
		X"3F",X"07",X"03",X"01",X"01",X"01",X"03",X"04",X"F0",X"C0",X"80",X"80",X"80",X"80",X"C0",X"20",
		X"01",X"03",X"07",X"05",X"05",X"07",X"0F",X"0F",X"00",X"40",X"20",X"20",X"20",X"40",X"C0",X"E0",
		X"1F",X"07",X"03",X"01",X"01",X"01",X"03",X"02",X"E0",X"C0",X"80",X"80",X"80",X"80",X"C0",X"40",
		X"01",X"03",X"07",X"05",X"05",X"07",X"0F",X"0F",X"00",X"20",X"10",X"10",X"10",X"20",X"40",X"C0",
		X"0F",X"07",X"03",X"01",X"01",X"00",X"00",X"00",X"E0",X"C0",X"80",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"18",X"1F",X"1F",X"00",X"00",X"00",X"20",X"30",X"F8",X"E0",X"C0",
		X"1F",X"2F",X"4F",X"7E",X"7C",X"78",X"30",X"00",X"80",X"80",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"1F",X"1F",X"00",X"00",X"00",X"20",X"30",X"F8",X"E0",X"C0",
		X"1F",X"2F",X"4F",X"7A",X"72",X"62",X"04",X"18",X"80",X"80",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"0F",X"1F",X"00",X"00",X"00",X"10",X"18",X"A0",X"C0",X"C0",
		X"1F",X"2F",X"4F",X"72",X"62",X"42",X"04",X"18",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"30",X"78",X"7C",X"7E",X"4F",X"2F",X"1F",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",X"80",
		X"1F",X"1F",X"18",X"10",X"00",X"00",X"00",X"00",X"C0",X"E0",X"F8",X"30",X"20",X"00",X"00",X"00",
		X"18",X"04",X"62",X"72",X"7A",X"4F",X"2F",X"1F",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",X"80",
		X"1F",X"1F",X"08",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"78",X"30",X"20",X"00",X"00",X"00",
		X"18",X"04",X"42",X"62",X"72",X"4F",X"2F",X"1F",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",
		X"1F",X"0F",X"08",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"A0",X"18",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"0C",X"1E",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"E0",
		X"03",X"03",X"03",X"07",X"0F",X"00",X"00",X"00",X"E0",X"F0",X"F8",X"FC",X"9E",X"5E",X"3C",X"00",
		X"00",X"00",X"00",X"04",X"0C",X"1E",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"E0",
		X"03",X"03",X"03",X"07",X"03",X"00",X"00",X"00",X"E0",X"FC",X"E2",X"F1",X"99",X"5C",X"3C",X"00",
		X"00",X"00",X"00",X"08",X"18",X"04",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",
		X"03",X"03",X"03",X"07",X"01",X"00",X"00",X"00",X"E0",X"FC",X"E2",X"E1",X"91",X"58",X"3C",X"00",
		X"00",X"00",X"00",X"0F",X"07",X"03",X"03",X"03",X"00",X"3C",X"5E",X"9E",X"FC",X"F8",X"F0",X"E0",
		X"03",X"07",X"1E",X"0C",X"04",X"00",X"00",X"00",X"E0",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"07",X"03",X"03",X"03",X"00",X"3C",X"5C",X"99",X"F1",X"E2",X"FC",X"E0",
		X"03",X"07",X"1E",X"0C",X"04",X"00",X"00",X"00",X"E0",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"07",X"03",X"03",X"03",X"00",X"3C",X"58",X"91",X"E1",X"E2",X"FC",X"E0",
		X"03",X"03",X"04",X"18",X"08",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"0F",X"10",X"11",X"8A",X"8A",X"3A",X"FC",X"68",
		X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"68",X"FC",X"3A",X"8A",X"8A",X"11",X"10",X"0F",
		X"00",X"00",X"00",X"00",X"06",X"06",X"03",X"00",X"00",X"08",X"14",X"22",X"11",X"38",X"FF",X"48",
		X"00",X"03",X"06",X"06",X"00",X"00",X"00",X"00",X"48",X"FF",X"38",X"11",X"22",X"14",X"08",X"00",
		X"00",X"00",X"00",X"30",X"30",X"1F",X"00",X"00",X"00",X"20",X"30",X"28",X"14",X"BA",X"79",X"78",
		X"00",X"00",X"1F",X"30",X"30",X"00",X"00",X"00",X"78",X"79",X"BA",X"14",X"28",X"30",X"20",X"00",
		X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"02",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"04",X"05",X"04",X"01",X"00",X"00",X"00",X"80",X"00",X"40",X"00",X"40",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"0B",X"08",X"0B",X"00",X"03",X"00",X"00",X"80",X"30",X"00",X"18",X"00",X"18",
		X"00",X"00",X"02",X"02",X"02",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"04",X"05",X"04",X"00",X"00",X"01",X"00",X"40",X"00",X"40",X"00",X"80",X"00",X"00",
		X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"0B",X"08",X"0B",X"00",X"00",X"01",X"18",X"00",X"18",X"00",X"30",X"80",X"00",X"00",
		X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"10",X"20",X"40",X"80",
		X"01",X"08",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"10",X"20",X"40",X"80",
		X"15",X"08",X"10",X"02",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"10",X"20",X"40",X"80",
		X"29",X"14",X"28",X"12",X"04",X"0A",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"08",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"20",X"00",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"02",X"10",X"08",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"20",X"10",X"00",X"00",X"00",X"00",
		X"00",X"04",X"0A",X"04",X"12",X"28",X"14",X"29",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"20",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"08",X"04",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"40",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"04",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"80",X"10",X"88",X"40",X"A0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"04",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"14",X"4A",X"A4",X"50",X"A0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"40",X"00",X"00",X"80",
		X"01",X"02",X"04",X"08",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"40",X"88",X"10",X"80",
		X"01",X"02",X"04",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"01",X"00",X"A0",X"50",X"A0",X"44",X"0A",X"14",X"00",
		X"02",X"04",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"33",X"0B",X"06",X"00",X"00",X"00",X"00",X"80",X"CC",X"D0",X"60",
		X"05",X"05",X"65",X"1D",X"0E",X"01",X"01",X"02",X"A0",X"A0",X"A6",X"B8",X"70",X"80",X"00",X"00",
		X"00",X"00",X"01",X"03",X"03",X"01",X"01",X"1E",X"00",X"00",X"80",X"C0",X"C0",X"80",X"80",X"78",
		X"25",X"05",X"05",X"05",X"0E",X"11",X"21",X"01",X"A4",X"A0",X"A0",X"A0",X"70",X"88",X"04",X"00",
		X"01",X"03",X"03",X"01",X"01",X"01",X"01",X"06",X"80",X"C0",X"C0",X"80",X"80",X"80",X"80",X"60",
		X"0D",X"15",X"15",X"05",X"06",X"09",X"08",X"08",X"B0",X"A8",X"A8",X"A0",X"60",X"90",X"90",X"50",
		X"02",X"01",X"01",X"0E",X"1D",X"65",X"05",X"05",X"00",X"00",X"80",X"70",X"B8",X"A6",X"A0",X"A0",
		X"06",X"0B",X"33",X"01",X"00",X"00",X"00",X"00",X"60",X"D0",X"CC",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"21",X"11",X"0E",X"05",X"05",X"05",X"25",X"00",X"04",X"88",X"70",X"A0",X"A0",X"A0",X"A4",
		X"1E",X"01",X"01",X"03",X"03",X"01",X"00",X"00",X"78",X"80",X"80",X"C0",X"C0",X"80",X"00",X"00",
		X"08",X"08",X"09",X"06",X"05",X"15",X"15",X"0D",X"50",X"90",X"90",X"60",X"A0",X"A8",X"A8",X"B0",
		X"06",X"01",X"01",X"01",X"01",X"03",X"03",X"01",X"60",X"80",X"80",X"80",X"80",X"C0",X"C0",X"80",
		X"00",X"00",X"04",X"04",X"02",X"01",X"07",X"0E",X"00",X"20",X"20",X"10",X"18",X"F8",X"08",X"F4",
		X"0E",X"07",X"01",X"02",X"04",X"04",X"00",X"00",X"F6",X"09",X"F8",X"18",X"10",X"20",X"20",X"00",
		X"00",X"00",X"00",X"01",X"01",X"01",X"19",X"3E",X"00",X"00",X"82",X"04",X"08",X"F8",X"08",X"F4",
		X"3E",X"19",X"01",X"01",X"01",X"00",X"00",X"00",X"F7",X"08",X"F8",X"08",X"04",X"82",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"61",X"FE",X"00",X"00",X"00",X"60",X"87",X"F8",X"09",X"F6",
		X"FE",X"61",X"01",X"00",X"00",X"00",X"00",X"00",X"F4",X"08",X"F8",X"87",X"60",X"00",X"00",X"00",
		X"00",X"04",X"04",X"08",X"18",X"1F",X"90",X"6F",X"00",X"00",X"20",X"20",X"40",X"80",X"E0",X"70",
		X"2F",X"10",X"1F",X"18",X"08",X"04",X"04",X"00",X"70",X"E0",X"80",X"40",X"20",X"20",X"00",X"00",
		X"00",X"00",X"41",X"20",X"10",X"1F",X"10",X"EF",X"00",X"00",X"00",X"80",X"80",X"80",X"98",X"7C",
		X"2F",X"10",X"1F",X"10",X"20",X"41",X"00",X"00",X"7C",X"98",X"80",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"06",X"E1",X"1F",X"10",X"2F",X"00",X"00",X"00",X"00",X"00",X"80",X"86",X"7F",
		X"6F",X"90",X"1F",X"E1",X"06",X"00",X"00",X"00",X"7F",X"86",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"34",X"3E",X"3F",X"36",X"6F",X"DF",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"30",X"D8",X"6C",X"34",X"1A",X"05",X"03",
		X"00",X"01",X"03",X"00",X"07",X"07",X"01",X"07",X"D6",X"FF",X"EF",X"41",X"EB",X"FB",X"1D",X"67",
		X"07",X"01",X"07",X"07",X"00",X"03",X"01",X"00",X"67",X"19",X"FB",X"EF",X"41",X"EB",X"EB",X"D6",
		X"00",X"00",X"00",X"3C",X"3E",X"00",X"01",X"3F",X"00",X"00",X"00",X"00",X"7C",X"FE",X"FF",X"FF",
		X"01",X"00",X"3E",X"3C",X"00",X"00",X"00",X"00",X"FF",X"FE",X"7C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"02",X"04",X"04",X"24",X"3C",X"07",X"C0",X"EC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"07",X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"FC",X"FC",X"EC",X"CC",X"C0",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"04",X"08",X"00",X"00",X"21",X"00",X"00",X"80",X"20",X"10",X"08",X"00",X"84",
		X"21",X"00",X"10",X"08",X"04",X"01",X"00",X"00",X"84",X"00",X"08",X"00",X"20",X"80",X"00",X"00",
		X"00",X"00",X"00",X"10",X"08",X"00",X"00",X"01",X"00",X"20",X"20",X"00",X"00",X"00",X"C2",X"24",
		X"01",X"00",X"04",X"08",X"00",X"00",X"00",X"00",X"20",X"C0",X"10",X"08",X"04",X"00",X"00",X"00",
		X"00",X"00",X"08",X"04",X"00",X"01",X"02",X"C4",X"00",X"80",X"80",X"02",X"04",X"80",X"40",X"20",
		X"04",X"02",X"01",X"00",X"00",X"00",X"20",X"40",X"20",X"40",X"80",X"00",X"00",X"08",X"04",X"00",
		X"00",X"00",X"06",X"88",X"08",X"20",X"20",X"20",X"40",X"00",X"E0",X"00",X"08",X"44",X"05",X"00",
		X"00",X"20",X"20",X"18",X"00",X"07",X"40",X"00",X"04",X"44",X"04",X"00",X"10",X"60",X"10",X"00",
		X"09",X"10",X"08",X"01",X"80",X"00",X"80",X"08",X"30",X"00",X"04",X"00",X"01",X"01",X"01",X"00",
		X"00",X"00",X"80",X"80",X"40",X"00",X"10",X"2D",X"08",X"80",X"01",X"01",X"02",X"40",X"08",X"30",
		X"00",X"00",X"07",X"0B",X"17",X"29",X"39",X"3E",X"00",X"00",X"E0",X"D0",X"E8",X"94",X"9C",X"7C",
		X"3E",X"39",X"29",X"17",X"0B",X"07",X"00",X"00",X"7C",X"9C",X"94",X"E8",X"D0",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
