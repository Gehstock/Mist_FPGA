library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ps06 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ps06 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"0A",X"03",X"0B",X"04",X"04",X"03",X"05",X"0C",X"06",X"03",X"07",X"04",X"08",X"03",X"07",X"03",
		X"06",X"03",X"05",X"03",X"04",X"03",X"0B",X"20",X"0A",X"FF",X"0E",X"0B",X"02",X"0A",X"07",X"09",
		X"03",X"08",X"03",X"07",X"03",X"06",X"03",X"05",X"08",X"02",X"01",X"05",X"01",X"06",X"08",X"08",
		X"02",X"07",X"02",X"06",X"06",X"04",X"02",X"0B",X"03",X"0A",X"07",X"09",X"03",X"08",X"01",X"07",
		X"01",X"06",X"02",X"00",X"02",X"01",X"0B",X"02",X"03",X"0B",X"03",X"0A",X"03",X"09",X"03",X"08",
		X"03",X"07",X"02",X"06",X"06",X"05",X"08",X"06",X"FF",X"01",X"00",X"01",X"01",X"06",X"02",X"08",
		X"05",X"02",X"07",X"08",X"08",X"02",X"07",X"02",X"06",X"02",X"05",X"07",X"02",X"01",X"05",X"01",
		X"06",X"01",X"07",X"08",X"08",X"02",X"09",X"08",X"0A",X"02",X"0B",X"06",X"03",X"03",X"0B",X"06",
		X"0A",X"02",X"09",X"06",X"08",X"02",X"07",X"04",X"06",X"02",X"05",X"05",X"04",X"03",X"05",X"02",
		X"06",X"02",X"07",X"06",X"08",X"03",X"09",X"05",X"0A",X"03",X"0B",X"04",X"04",X"03",X"05",X"03",
		X"06",X"03",X"07",X"03",X"08",X"04",X"09",X"05",X"0A",X"02",X"0B",X"03",X"04",X"01",X"05",X"01",
		X"06",X"01",X"07",X"04",X"08",X"02",X"07",X"01",X"06",X"01",X"00",X"01",X"01",X"0A",X"02",X"02",
		X"05",X"02",X"06",X"02",X"07",X"02",X"08",X"02",X"09",X"0A",X"0A",X"03",X"0B",X"03",X"04",X"03",
		X"05",X"03",X"06",X"02",X"07",X"02",X"08",X"02",X"08",X"10",X"0A",X"02",X"09",X"02",X"08",X"02",
		X"07",X"03",X"06",X"FF",X"00",X"00",X"60",X"1F",X"60",X"00",X"00",X"00",X"10",X"10",X"10",X"10",
		X"10",X"10",X"28",X"28",X"28",X"28",X"10",X"10",X"10",X"10",X"10",X"10",X"21",X"1C",X"1C",X"1B",
		X"1D",X"1C",X"1C",X"1C",X"1D",X"21",X"1C",X"1C",X"1E",X"1C",X"1C",X"1C",X"00",X"00",X"01",X"00",
		X"00",X"00",X"90",X"60",X"40",X"08",X"41",X"10",X"00",X"10",X"01",X"00",X"00",X"62",X"0D",X"00",
		X"08",X"F4",X"F8",X"11",X"00",X"38",X"B2",X"02",X"60",X"AB",X"C7",X"07",X"40",X"DB",X"DB",X"37",
		X"00",X"FD",X"3F",X"03",X"80",X"3D",X"FE",X"02",X"C1",X"8B",X"F1",X"07",X"E0",X"E7",X"F7",X"0F",
		X"E0",X"EC",X"AE",X"09",X"C0",X"DC",X"76",X"0D",X"80",X"8C",X"B9",X"05",X"80",X"2C",X"DF",X"03",
		X"C0",X"78",X"D3",X"03",X"20",X"59",X"EE",X"03",X"90",X"F9",X"FF",X"01",X"80",X"F1",X"C7",X"04",
		X"84",X"7B",X"17",X"10",X"80",X"F7",X"FB",X"02",X"00",X"2F",X"39",X"04",X"00",X"1E",X"1C",X"00",
		X"00",X"8C",X"01",X"10",X"00",X"80",X"00",X"00",X"00",X"80",X"00",X"41",X"10",X"00",X"04",X"C2",
		X"08",X"80",X"0C",X"00",X"21",X"94",X"20",X"97",X"BE",X"C8",X"23",X"BE",X"C2",X"20",X"10",X"23",
		X"BE",X"C2",X"9B",X"49",X"34",X"CD",X"E5",X"49",X"22",X"99",X"20",X"21",X"99",X"20",X"CD",X"ED",
		X"49",X"21",X"99",X"20",X"7E",X"FE",X"28",X"DA",X"D6",X"49",X"23",X"7E",X"FE",X"2C",X"DA",X"D6",
		X"49",X"FE",X"EC",X"D2",X"D6",X"49",X"3A",X"F7",X"20",X"A7",X"C2",X"C3",X"49",X"CD",X"11",X"4A",
		X"22",X"97",X"20",X"21",X"97",X"20",X"EF",X"2A",X"99",X"20",X"CD",X"09",X"4A",X"21",X"99",X"20",
		X"CD",X"C4",X"04",X"C3",X"AC",X"03",X"21",X"F7",X"20",X"36",X"00",X"2E",X"94",X"11",X"94",X"40",
		X"06",X"0B",X"C3",X"BB",X"04",X"2A",X"EA",X"20",X"01",X"00",X"07",X"09",X"C9",X"E5",X"CD",X"C4",
		X"04",X"7D",X"FE",X"78",X"3E",X"07",X"DA",X"FB",X"49",X"3E",X"02",X"F5",X"FF",X"F1",X"11",X"02",
		X"03",X"DF",X"E1",X"CD",X"C4",X"04",X"C3",X"EF",X"08",X"FF",X"3E",X"04",X"11",X"02",X"03",X"DF",
		X"C9",X"CD",X"37",X"4A",X"DA",X"2F",X"4A",X"CD",X"42",X"4A",X"D2",X"31",X"4A",X"CD",X"4A",X"4A",
		X"D5",X"22",X"9B",X"20",X"21",X"99",X"20",X"CD",X"03",X"4A",X"D1",X"21",X"F7",X"20",X"34",X"EB",
		X"C9",X"CD",X"55",X"4A",X"C3",X"20",X"4A",X"2B",X"3A",X"04",X"20",X"C6",X"05",X"BE",X"11",X"FC",
		X"00",X"C9",X"23",X"3A",X"05",X"20",X"C6",X"0A",X"BE",X"C9",X"2B",X"CD",X"03",X"4A",X"11",X"00",
		X"FC",X"21",X"EC",X"48",X"C9",X"2B",X"CD",X"03",X"4A",X"11",X"00",X"04",X"21",X"F4",X"48",X"C9",
		X"21",X"9F",X"20",X"97",X"BE",X"C8",X"23",X"BE",X"C2",X"72",X"4A",X"34",X"CD",X"E5",X"49",X"22",
		X"A3",X"20",X"21",X"A3",X"20",X"CD",X"ED",X"49",X"21",X"A3",X"20",X"7E",X"FE",X"28",X"DA",X"CF",
		X"4A",X"23",X"7E",X"FE",X"2C",X"DA",X"CF",X"4A",X"FE",X"EC",X"D2",X"CF",X"4A",X"3A",X"F8",X"20",
		X"A7",X"C2",X"BF",X"4A",X"CD",X"37",X"4A",X"DA",X"B2",X"4A",X"CD",X"42",X"4A",X"D2",X"B9",X"4A",
		X"CD",X"4A",X"4A",X"D5",X"22",X"A5",X"20",X"21",X"A3",X"20",X"CD",X"03",X"4A",X"D1",X"21",X"F8",
		X"20",X"34",X"EB",X"22",X"A1",X"20",X"C3",X"BF",X"4A",X"CD",X"55",X"4A",X"C3",X"A3",X"4A",X"21",
		X"A1",X"20",X"EF",X"2A",X"A3",X"20",X"CD",X"09",X"4A",X"21",X"A3",X"20",X"C3",X"D0",X"49",X"21",
		X"F8",X"20",X"36",X"00",X"2E",X"9F",X"11",X"9F",X"40",X"06",X"0A",X"C3",X"BB",X"04",X"21",X"D4",
		X"20",X"AF",X"BE",X"C8",X"23",X"BE",X"C2",X"20",X"10",X"23",X"BE",X"C2",X"F5",X"4A",X"34",X"CD",
		X"E5",X"49",X"22",X"D9",X"20",X"21",X"D9",X"20",X"CD",X"ED",X"49",X"21",X"D9",X"20",X"7E",X"FE",
		X"28",X"DA",X"4F",X"4B",X"23",X"7E",X"FE",X"2C",X"DA",X"4F",X"4B",X"FE",X"EC",X"D2",X"4F",X"4B",
		X"3A",X"F9",X"20",X"A7",X"C2",X"39",X"4B",X"CD",X"37",X"4A",X"DA",X"35",X"4B",X"CD",X"42",X"4A",
		X"D2",X"49",X"4B",X"CD",X"4A",X"4A",X"D5",X"22",X"DB",X"20",X"21",X"D9",X"20",X"CD",X"03",X"4A",
		X"D1",X"21",X"F9",X"20",X"34",X"EB",X"22",X"D7",X"20",X"21",X"D7",X"20",X"EF",X"2A",X"D9",X"20",
		X"CD",X"09",X"4A",X"21",X"D9",X"20",X"C3",X"D0",X"49",X"CD",X"55",X"4A",X"C3",X"26",X"4B",X"21",
		X"F9",X"20",X"36",X"00",X"2E",X"D4",X"11",X"D4",X"40",X"C3",X"E0",X"49",X"21",X"FA",X"20",X"97",
		X"BE",X"C8",X"CD",X"ED",X"0E",X"FE",X"20",X"21",X"00",X"FB",X"D2",X"76",X"4B",X"FE",X"16",X"26",
		X"FC",X"D2",X"76",X"4B",X"26",X"FE",X"22",X"FB",X"20",X"2A",X"FD",X"20",X"E5",X"FF",X"3E",X"07",
		X"11",X"01",X"05",X"DF",X"E1",X"06",X"0E",X"11",X"B7",X"42",X"CD",X"EF",X"08",X"21",X"FE",X"20",
		X"7E",X"FE",X"30",X"DC",X"AE",X"4B",X"21",X"FB",X"20",X"EF",X"2A",X"FD",X"20",X"E5",X"FF",X"3E",
		X"00",X"11",X"01",X"05",X"DF",X"E1",X"06",X"0E",X"11",X"B7",X"42",X"C3",X"AC",X"03",X"36",X"E8",
		X"C9",X"21",X"16",X"2C",X"11",X"04",X"4C",X"0E",X"0B",X"CD",X"54",X"03",X"DB",X"01",X"07",X"DA",
		X"D6",X"4B",X"07",X"07",X"07",X"07",X"DA",X"A0",X"04",X"07",X"DA",X"E9",X"4B",X"07",X"DA",X"F2",
		X"4B",X"D3",X"05",X"C3",X"BC",X"4B",X"CD",X"ED",X"0E",X"C6",X"01",X"27",X"77",X"26",X"22",X"77",
		X"CD",X"85",X"03",X"CD",X"E9",X"0A",X"C3",X"BC",X"4B",X"CD",X"ED",X"18",X"CD",X"85",X"03",X"C3",
		X"BC",X"4B",X"21",X"03",X"23",X"36",X"22",X"E5",X"CD",X"ED",X"18",X"CD",X"85",X"03",X"E1",X"36",
		X"21",X"C3",X"BC",X"4B",X"0F",X"11",X"04",X"12",X"04",X"13",X"1B",X"0C",X"0E",X"03",X"04",X"06",
		X"01",X"21",X"00",X"20",X"70",X"2E",X"4F",X"70",X"2E",X"BE",X"70",X"E7",X"2E",X"4B",X"7E",X"FE",
		X"06",X"DA",X"50",X"4C",X"2E",X"00",X"36",X"00",X"2E",X"4C",X"7E",X"FE",X"06",X"DA",X"5C",X"4C",
		X"2E",X"13",X"36",X"00",X"2E",X"3D",X"AF",X"BE",X"C2",X"68",X"4C",X"2E",X"40",X"AF",X"BE",X"C2",
		X"71",X"4C",X"2E",X"49",X"36",X"00",X"2E",X"26",X"11",X"26",X"41",X"06",X"13",X"C3",X"BB",X"04",
		X"E5",X"21",X"72",X"20",X"70",X"2E",X"7B",X"70",X"E1",X"C3",X"28",X"4C",X"E5",X"21",X"84",X"20",
		X"70",X"2E",X"8D",X"70",X"E1",X"C3",X"34",X"4C",X"E5",X"21",X"C5",X"20",X"70",X"E1",X"C3",X"3B",
		X"4C",X"E5",X"21",X"CC",X"20",X"70",X"E1",X"C3",X"42",X"4C",X"CD",X"A0",X"04",X"CD",X"A8",X"06",
		X"CD",X"92",X"0A",X"21",X"E0",X"20",X"11",X"CE",X"4C",X"06",X"0C",X"CD",X"BB",X"04",X"2E",X"04",
		X"36",X"50",X"21",X"0B",X"23",X"34",X"CD",X"D4",X"01",X"21",X"0D",X"20",X"36",X"00",X"2E",X"EA",
		X"7E",X"FE",X"94",X"D3",X"05",X"D2",X"99",X"4C",X"CD",X"CD",X"4E",X"21",X"12",X"CC",X"11",X"02",
		X"16",X"3E",X"05",X"DF",X"21",X"0B",X"23",X"36",X"00",X"CD",X"85",X"03",X"21",X"12",X"2C",X"11",
		X"FD",X"4C",X"01",X"02",X"58",X"CD",X"A8",X"05",X"CD",X"73",X"03",X"C3",X"F0",X"04",X"DA",X"4C",
		X"00",X"01",X"01",X"01",X"07",X"05",X"00",X"00",X"E0",X"E0",X"07",X"05",X"08",X"06",X"03",X"07",
		X"03",X"08",X"03",X"09",X"03",X"0A",X"03",X"0B",X"03",X"04",X"03",X"05",X"03",X"06",X"03",X"07",
		X"03",X"08",X"03",X"09",X"07",X"0A",X"02",X"0B",X"01",X"04",X"07",X"02",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"C0",X"F3",X"C0",X"F3",X"C0",X"F3",X"C0",X"F3",X"C0",X"FF",X"C0",
		X"FF",X"80",X"7F",X"00",X"3F",X"00",X"00",X"00",X"00",X"FC",X"3F",X"FE",X"7F",X"FF",X"FF",X"FF",
		X"FF",X"03",X"C0",X"03",X"C0",X"FF",X"FF",X"FF",X"FF",X"FE",X"7F",X"FC",X"3F",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"00",X"07",X"00",X"07",X"00",X"07",
		X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"FF",X"0F",X"FF",
		X"3F",X"FF",X"7F",X"FF",X"FF",X"C0",X"E3",X"C0",X"E3",X"C0",X"E3",X"FF",X"FF",X"FF",X"7F",X"FF",
		X"3F",X"FF",X"0F",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C0",
		X"F3",X"E0",X"F3",X"F0",X"F3",X"FC",X"F3",X"FF",X"FF",X"DF",X"FF",X"8F",X"7F",X"07",X"3F",X"00",
		X"00",X"00",X"00",X"01",X"80",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"80",X"00",
		X"00",X"00",X"00",X"3C",X"00",X"3E",X"3E",X"3F",X"7F",X"8F",X"FF",X"87",X"FF",X"C7",X"E3",X"C7",
		X"E3",X"C7",X"E3",X"FF",X"E1",X"FF",X"F1",X"FE",X"FC",X"7C",X"7C",X"00",X"3C",X"FE",X"FF",X"CA",
		X"02",X"4E",X"FE",X"FE",X"CA",X"F7",X"4D",X"21",X"28",X"23",X"36",X"80",X"23",X"77",X"23",X"EB",
		X"21",X"36",X"4E",X"87",X"4F",X"06",X"00",X"09",X"7E",X"23",X"66",X"6F",X"C3",X"DD",X"4D",X"3A",
		X"28",X"23",X"A7",X"C8",X"21",X"2A",X"23",X"35",X"C0",X"EB",X"2A",X"2B",X"23",X"7E",X"A7",X"CA",
		X"02",X"4E",X"FE",X"FF",X"CA",X"F1",X"4D",X"12",X"23",X"7E",X"D3",X"02",X"23",X"22",X"2B",X"23",
		X"C9",X"3A",X"29",X"23",X"F2",X"B7",X"4D",X"3E",X"01",X"32",X"2A",X"23",X"3E",X"80",X"32",X"28",
		X"23",X"C9",X"3E",X"FF",X"D3",X"02",X"AF",X"32",X"28",X"23",X"32",X"4A",X"20",X"C9",X"21",X"26",
		X"23",X"7E",X"3D",X"77",X"C0",X"2B",X"7E",X"23",X"77",X"23",X"7E",X"A7",X"C2",X"22",X"4E",X"C3",
		X"CF",X"4D",X"3A",X"23",X"23",X"CD",X"AD",X"4D",X"AF",X"32",X"27",X"23",X"C9",X"AF",X"32",X"24",
		X"23",X"3C",X"32",X"27",X"23",X"C9",X"5B",X"4E",X"5F",X"4E",X"7F",X"4E",X"CB",X"4E",X"11",X"73",
		X"41",X"21",X"23",X"23",X"06",X"06",X"C3",X"BB",X"04",X"01",X"00",X"05",X"05",X"01",X"00",X"02",
		X"00",X"05",X"05",X"01",X"00",X"03",X"00",X"05",X"05",X"01",X"00",X"01",X"FF",X"00",X"00",X"01",
		X"E6",X"01",X"E9",X"01",X"EB",X"01",X"EC",X"01",X"EE",X"01",X"F0",X"01",X"F2",X"02",X"F3",X"01",
		X"F2",X"01",X"F0",X"01",X"EE",X"01",X"EC",X"01",X"EB",X"01",X"E9",X"01",X"E6",X"00",X"00",X"02",
		X"B9",X"02",X"CC",X"02",X"D7",X"02",X"CC",X"01",X"D7",X"01",X"D9",X"02",X"D7",X"02",X"CC",X"02",
		X"D7",X"01",X"DD",X"01",X"E1",X"02",X"DD",X"02",X"D7",X"02",X"DD",X"01",X"D7",X"01",X"CC",X"01",
		X"D7",X"01",X"D9",X"04",X"CC",X"02",X"B9",X"02",X"CC",X"02",X"D7",X"02",X"CC",X"01",X"D7",X"01",
		X"D9",X"02",X"D7",X"02",X"CC",X"02",X"D7",X"01",X"DD",X"01",X"CC",X"01",X"D7",X"01",X"DD",X"01",
		X"E6",X"01",X"DD",X"01",X"E6",X"01",X"EB",X"04",X"E6",X"00",X"00",X"00",X"00",X"CD",X"15",X"02",
		X"21",X"11",X"2C",X"01",X"04",X"60",X"C3",X"10",X"09",X"2D",X"53",X"50",X"45",X"45",X"44",X"0D",
		X"0A",X"09",X"44",X"42",X"09",X"30",X"30",X"09",X"09",X"3B",X"59",X"2D",X"53",X"50",X"45",X"45",
		X"44",X"0D",X"0A",X"09",X"44",X"42",X"09",X"30",X"42",X"30",X"48",X"09",X"09",X"3B",X"53",X"2D",
		X"CD",X"05",X"04",X"E6",X"F0",X"FE",X"80",X"CA",X"52",X"0C",X"FE",X"40",X"CA",X"78",X"0C",X"FE",
		X"20",X"CA",X"9C",X"0C",X"FE",X"10",X"CA",X"B6",X"0C",X"FE",X"C0",X"CA",X"30",X"4F",X"FE",X"90",
		X"CA",X"58",X"4F",X"FE",X"60",X"CA",X"78",X"4F",X"FE",X"30",X"CA",X"9F",X"4F",X"C3",X"F7",X"0B",
		X"21",X"3E",X"20",X"11",X"04",X"20",X"1A",X"BE",X"D2",X"F7",X"0B",X"23",X"23",X"13",X"1A",X"BE",
		X"DA",X"F7",X"0B",X"CD",X"8B",X"0C",X"CD",X"95",X"0C",X"CD",X"4F",X"4F",X"C3",X"FA",X"0B",X"CD",
		X"62",X"0C",X"2E",X"01",X"D0",X"2E",X"02",X"C9",X"21",X"3E",X"20",X"3A",X"04",X"20",X"BE",X"D2",
		X"F7",X"0B",X"21",X"41",X"20",X"3A",X"05",X"20",X"BE",X"D2",X"F7",X"0B",X"CD",X"C9",X"0C",X"CD",
		X"D3",X"0C",X"CD",X"4F",X"4F",X"C3",X"FA",X"0B",X"21",X"3F",X"20",X"11",X"04",X"20",X"1A",X"BE",
		X"DA",X"F7",X"0B",X"23",X"13",X"1A",X"BE",X"DA",X"F7",X"0B",X"CD",X"AC",X"0C",X"CD",X"96",X"4F",
		X"CD",X"95",X"0C",X"C3",X"FA",X"0B",X"CD",X"62",X"0C",X"26",X"FE",X"D0",X"26",X"FD",X"C9",X"21",
		X"3F",X"20",X"3A",X"04",X"20",X"BE",X"DA",X"F7",X"0B",X"23",X"23",X"3A",X"05",X"20",X"BE",X"D2",
		X"F7",X"0B",X"CD",X"AC",X"0C",X"CD",X"BE",X"4F",X"CD",X"D3",X"0C",X"C3",X"FA",X"0B",X"CD",X"62",
		X"0C",X"26",X"02",X"D0",X"26",X"03",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
