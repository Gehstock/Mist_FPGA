library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity swimmer_big_sprite_tile_bit1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of swimmer_big_sprite_tile_bit1 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"07",X"0F",X"07",X"0F",X"00",X"00",X"00",X"80",X"C0",X"80",X"80",X"90",
		X"0F",X"7E",X"FE",X"FF",X"CF",X"EF",X"EF",X"EF",X"30",X"3E",X"7F",X"FF",X"F3",X"F7",X"F7",X"F7",
		X"00",X"00",X"00",X"00",X"00",X"39",X"38",X"39",X"00",X"00",X"00",X"60",X"F4",X"FA",X"B8",X"B8",
		X"30",X"33",X"3F",X"3F",X"3F",X"01",X"01",X"03",X"F8",X"F8",X"FF",X"FF",X"FF",X"FE",X"FC",X"CC",
		X"00",X"00",X"03",X"07",X"0F",X"07",X"0F",X"0F",X"00",X"00",X"80",X"C0",X"80",X"80",X"90",X"30",
		X"1E",X"3E",X"3F",X"3F",X"3F",X"3E",X"23",X"76",X"38",X"7C",X"FC",X"FC",X"EC",X"67",X"27",X"47",
		X"00",X"00",X"01",X"02",X"02",X"02",X"04",X"05",X"1F",X"CF",X"27",X"13",X"13",X"09",X"C9",X"28",
		X"05",X"05",X"05",X"01",X"00",X"00",X"00",X"00",X"28",X"24",X"14",X"14",X"14",X"14",X"04",X"04",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"31",X"F8",X"E0",X"E2",X"C7",X"FF",X"FF",X"FF",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"1F",X"7F",X"FF",X"FF",X"FF",X"F3",X"31",X"FF",X"3F",X"FF",X"FF",X"FF",X"FF",X"DD",X"D0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"31",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DC",X"10",
		X"01",X"03",X"0E",X"0C",X"1C",X"38",X"F0",X"F8",X"F8",X"E0",X"00",X"07",X"1C",X"38",X"30",X"70",
		X"F0",X"FF",X"FF",X"FE",X"FF",X"DC",X"DF",X"CC",X"70",X"E0",X"80",X"00",X"00",X"0C",X"FF",X"E0",
		X"00",X"00",X"00",X"30",X"30",X"38",X"3B",X"3F",X"00",X"00",X"00",X"0C",X"0C",X"1C",X"9C",X"DC",
		X"3F",X"3F",X"3F",X"3F",X"3E",X"1E",X"1F",X"0F",X"8C",X"9C",X"9C",X"3C",X"3C",X"7C",X"F8",X"F8",
		X"16",X"1B",X"36",X"37",X"6F",X"6E",X"78",X"78",X"40",X"20",X"40",X"60",X"E4",X"EC",X"7C",X"7C",
		X"7C",X"3C",X"1C",X"1C",X"1C",X"00",X"00",X"00",X"3C",X"3C",X"3C",X"3C",X"3C",X"7C",X"7C",X"00",
		X"1F",X"3F",X"3F",X"3B",X"3D",X"3D",X"3C",X"3C",X"E4",X"C4",X"C8",X"EC",X"DC",X"77",X"7F",X"7F",
		X"7C",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"7E",X"78",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"27",X"6E",X"6E",X"7D",X"78",X"78",X"7C",X"6F",X"6F",X"FF",X"FB",X"00",X"00",X"00",X"00",
		X"3C",X"1C",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"60",X"F0",X"F0",X"78",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"7F",
		X"00",X"00",X"40",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"40",X"60",X"78",X"78",X"F0",X"F0",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"60",X"40",X"F8",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"0E",X"1F",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"05",X"07",X"07",X"0F",X"0F",X"E0",X"F7",X"FB",X"FB",
		X"0E",X"0F",X"1F",X"5F",X"DF",X"DF",X"BF",X"BF",X"00",X"04",X"AB",X"D7",X"E7",X"EF",X"EF",X"DF",
		X"BF",X"DF",X"C7",X"81",X"00",X"FC",X"FB",X"F7",X"DF",X"DF",X"BF",X"BF",X"7F",X"7F",X"FF",X"FF",
		X"07",X"07",X"03",X"7B",X"F9",X"FB",X"F7",X"F7",X"F8",X"F8",X"78",X"B0",X"80",X"A2",X"32",X"77",
		X"2F",X"07",X"0F",X"00",X"00",X"00",X"00",X"00",X"77",X"1F",X"0F",X"1F",X"1E",X"1C",X"1C",X"1C",
		X"06",X"04",X"02",X"06",X"27",X"37",X"3E",X"3E",X"68",X"D8",X"6C",X"EC",X"F6",X"76",X"1E",X"1E",
		X"3C",X"3C",X"3C",X"3C",X"3C",X"3E",X"3E",X"00",X"3E",X"3C",X"38",X"38",X"38",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"E0",
		X"60",X"60",X"E0",X"E0",X"E0",X"00",X"00",X"00",X"60",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"78",X"78",X"70",X"60",X"78",X"38",X"1C",X"0C",
		X"80",X"80",X"C0",X"C0",X"00",X"00",X"00",X"00",X"0F",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"1F",X"07",X"01",X"00",X"00",X"0F",X"7F",X"3F",X"DF",X"DF",X"9F",X"1F",X"BF",X"BF",X"BF",X"BF",
		X"9F",X"CF",X"E7",X"F2",X"F8",X"FC",X"FC",X"FC",X"C7",X"87",X"03",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C7",X"83",X"03",X"07",X"0F",X"10",X"00",X"00",X"00",X"00",
		X"83",X"83",X"C7",X"FF",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"80",X"00",X"00",X"00",X"00",X"00",X"FF",X"83",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"3F",X"00",X"00",X"00",X"00",X"01",X"7F",X"FF",X"E0",
		X"FF",X"FF",X"3F",X"0F",X"07",X"03",X"03",X"07",X"BF",X"9F",X"C7",X"F1",X"FC",X"FF",X"FF",X"FE",
		X"07",X"13",X"18",X"3E",X"FC",X"F0",X"80",X"00",X"FC",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"70",X"F8",X"00",X"00",X"00",X"00",X"02",X"07",X"07",X"17",
		X"00",X"00",X"00",X"01",X"03",X"03",X"07",X"07",X"37",X"67",X"EF",X"EF",X"EF",X"EF",X"EF",X"F3",
		X"01",X"03",X"07",X"0B",X"1D",X"3F",X"80",X"DF",X"FC",X"FC",X"FB",X"F7",X"F7",X"EF",X"0F",X"DF",
		X"EF",X"F7",X"FB",X"FD",X"FE",X"FC",X"FB",X"F7",X"DF",X"DF",X"BF",X"3F",X"7F",X"7F",X"FF",X"FF",
		X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"C1",X"E3",X"E7",X"F7",X"F7",X"FB",X"70",X"F0",X"F8",X"FA",X"FB",X"FB",X"FD",X"FD",
		X"FB",X"FB",X"FD",X"FD",X"FE",X"FE",X"FF",X"FF",X"FD",X"E3",X"81",X"00",X"00",X"3F",X"DF",X"EF",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"3F",X"3F",X"DF",X"EF",X"EF",X"F7",X"F0",X"FB",
		X"E0",X"E0",X"F0",X"F0",X"07",X"EF",X"DF",X"DF",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"A0",
		X"80",X"C0",X"E0",X"D0",X"B8",X"FC",X"01",X"FB",X"00",X"00",X"00",X"00",X"40",X"E0",X"E0",X"E8",
		X"FB",X"FB",X"FD",X"FD",X"FE",X"FE",X"FF",X"FF",X"F7",X"EF",X"DF",X"BF",X"7F",X"3F",X"DF",X"EF",
		X"FC",X"FC",X"FE",X"FF",X"F0",X"00",X"FF",X"FF",X"03",X"01",X"00",X"00",X"00",X"00",X"FC",X"FF",
		X"EC",X"EE",X"F7",X"F7",X"F7",X"F7",X"F7",X"CF",X"00",X"00",X"00",X"80",X"C0",X"C0",X"E0",X"E0",
		X"00",X"07",X"18",X"60",X"40",X"81",X"83",X"84",X"00",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",
		X"84",X"82",X"81",X"C0",X"60",X"78",X"3F",X"1F",X"7F",X"3F",X"FF",X"03",X"00",X"00",X"F0",X"F8",
		X"0F",X"0F",X"30",X"27",X"2F",X"2F",X"2F",X"2F",X"E1",X"C0",X"00",X"00",X"F8",X"FF",X"FF",X"FF",
		X"37",X"33",X"35",X"36",X"03",X"03",X"01",X"00",X"FF",X"FF",X"FC",X"00",X"E0",X"EF",X"FF",X"FF",
		X"F7",X"77",X"37",X"2F",X"0F",X"EF",X"CF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"DF",X"DF",X"1F",X"1F",X"BF",X"BF",X"BC",X"B8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"C0",X"80",X"80",X"80",X"9F",X"FF",X"FF",X"FF",X"03",X"01",X"00",X"01",X"F9",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"EF",X"EE",X"F1",X"F3",X"F7",X"F3",X"FB",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E3",X"C1",X"FB",X"F9",X"FA",X"FB",X"FD",X"FD",X"FD",X"FD",
		X"BF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"A0",X"B0",X"B0",X"78",X"78",X"7C",X"FC",X"3E",
		X"F8",X"E0",X"00",X"F0",X"FE",X"FF",X"F1",X"E0",X"1E",X"1E",X"0E",X"06",X"1E",X"1C",X"38",X"30",
		X"00",X"FF",X"01",X"01",X"01",X"F1",X"F1",X"F1",X"00",X"9F",X"91",X"D1",X"D1",X"F1",X"F1",X"F1",
		X"F1",X"F1",X"F1",X"F1",X"F1",X"71",X"31",X"31",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",
		X"00",X"9F",X"90",X"D0",X"D0",X"F1",X"F1",X"F1",X"00",X"FF",X"00",X"00",X"00",X"F1",X"F1",X"F1",
		X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",
		X"00",X"FF",X"30",X"30",X"30",X"F0",X"F0",X"F1",X"00",X"F1",X"0A",X"0A",X"04",X"00",X"00",X"80",
		X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"40",X"A0",X"91",X"9F",X"DF",X"DF",X"FF",X"FF",
		X"01",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"9F",X"CF",X"E7",X"F2",X"F8",X"FC",X"FC",X"FC",
		X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"FD",X"F7",X"EF",X"CF",X"9E",X"BE",X"3E",X"7F",
		X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"3F",X"7F",X"FF",X"07",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"03",X"00",X"00",X"00",X"00",X"80",X"F0",X"FC",X"FE",X"1F",X"03",X"01",X"00",
		X"87",X"C0",X"C0",X"C0",X"E0",X"00",X"00",X"00",X"E1",X"03",X"03",X"03",X"07",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C1",X"C3",X"00",X"07",X"1F",X"3F",X"7F",X"F0",X"E0",X"C0",
		X"C1",X"C1",X"E3",X"FF",X"F0",X"00",X"00",X"00",X"E7",X"E1",X"C0",X"00",X"00",X"00",X"00",X"3C",
		X"03",X"FF",X"FF",X"F6",X"80",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"3F",X"0F",X"07",X"07",X"07",
		X"CF",X"DF",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"70",X"00",X"80",X"80",X"80",X"C0",X"C0",X"E0",
		X"3F",X"87",X"C3",X"F1",X"F8",X"FF",X"FF",X"FE",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"31",X"00",X"F1",X"0A",X"0A",X"04",X"00",X"00",X"80",
		X"51",X"B1",X"31",X"31",X"71",X"71",X"F1",X"F1",X"40",X"20",X"11",X"1F",X"1F",X"1E",X"3F",X"3F",
		X"00",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"00",X"00",X"00",X"F8",X"F8",X"F8",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"F8",X"F8",X"F8",X"18",X"18",X"18",X"F8",X"F8",
		X"00",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"E0",X"18",X"06",X"02",X"81",X"C1",X"21",
		X"FE",X"FC",X"FF",X"00",X"00",X"00",X"FE",X"FE",X"21",X"41",X"81",X"02",X"06",X"38",X"20",X"20",
		X"E1",X"03",X"03",X"03",X"06",X"00",X"07",X"7F",X"7E",X"FC",X"39",X"03",X"00",X"00",X"00",X"00",
		X"05",X"0D",X"0D",X"1E",X"1E",X"3E",X"3F",X"7C",X"FD",X"FE",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",
		X"00",X"00",X"00",X"80",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",
		X"F7",X"F7",X"77",X"8F",X"CF",X"EF",X"CF",X"DF",X"EF",X"EE",X"EC",X"F4",X"F0",X"F7",X"F7",X"FB",
		X"46",X"0E",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"1F",X"00",
		X"81",X"00",X"00",X"00",X"1F",X"FF",X"FF",X"FF",X"F0",X"F0",X"14",X"EC",X"F4",X"F4",X"F4",X"F4",
		X"00",X"00",X"00",X"00",X"07",X"FF",X"FF",X"00",X"0F",X"03",X"1D",X"3E",X"FE",X"F8",X"C0",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"FB",X"F9",X"FA",X"FB",X"FD",X"FD",X"3D",X"1D",
		X"FC",X"F0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"C0",X"C0",X"E0",
		X"FF",X"FF",X"0F",X"F1",X"FE",X"FF",X"F1",X"E0",X"D4",X"BC",X"BC",X"6C",X"C0",X"C0",X"80",X"00",
		X"00",X"FF",X"01",X"01",X"01",X"01",X"01",X"31",X"00",X"3F",X"30",X"70",X"70",X"F1",X"F1",X"F1",
		X"51",X"B1",X"31",X"71",X"71",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F0",X"F0",X"F0",X"F1",X"F1",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"F8",X"F8",X"F8",X"F8",X"18",X"18",X"18",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"F8",X"00",
		X"FE",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"20",X"10",X"08",X"07",X"01",X"01",X"C1",X"FF",
		X"FF",X"FF",X"7F",X"7F",X"3F",X"3F",X"1F",X"00",X"FF",X"FE",X"FC",X"F8",X"F0",X"E0",X"C0",X"00",
		X"0F",X"07",X"03",X"FF",X"80",X"80",X"80",X"FF",X"FC",X"FC",X"F8",X"F0",X"00",X"00",X"03",X"FF",
		X"FF",X"7F",X"3F",X"1F",X"0F",X"07",X"03",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"31",X"30",X"30",X"30",X"78",X"F8",X"FC",X"FF",X"F1",X"E0",X"40",X"00",X"00",X"04",X"1F",X"FF",
		X"FF",X"FF",X"FF",X"FD",X"FC",X"F0",X"C0",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3E",X"00",
		X"F1",X"E1",X"41",X"01",X"03",X"03",X"07",X"FF",X"F1",X"F1",X"F1",X"F1",X"80",X"80",X"80",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"1E",X"00",X"FF",X"FF",X"FF",X"FF",X"BF",X"3F",X"1F",X"00",
		X"F1",X"F1",X"F1",X"F1",X"01",X"01",X"01",X"FF",X"FF",X"FF",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"00",
		X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"FF",X"7F",X"7B",X"03",X"03",X"03",X"03",X"03",X"03",
		X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"FC",X"00",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"00",
		X"F1",X"F1",X"F1",X"F1",X"F0",X"F0",X"F0",X"FF",X"F1",X"F1",X"F1",X"F1",X"00",X"00",X"00",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"07",X"0F",X"07",X"0F",X"00",X"00",X"00",X"80",X"C0",X"80",X"80",X"90",
		X"0F",X"7E",X"FE",X"FF",X"CF",X"EF",X"EF",X"EF",X"30",X"3E",X"7F",X"FF",X"F3",X"F7",X"F7",X"F7",
		X"00",X"00",X"00",X"00",X"00",X"39",X"38",X"39",X"00",X"00",X"00",X"60",X"F4",X"FA",X"B8",X"B8",
		X"30",X"33",X"3F",X"3F",X"3F",X"01",X"01",X"03",X"F8",X"F8",X"FF",X"FF",X"FF",X"FE",X"FC",X"CC",
		X"00",X"00",X"03",X"07",X"0F",X"07",X"0F",X"0F",X"00",X"00",X"80",X"C0",X"80",X"80",X"90",X"30",
		X"1E",X"3E",X"3F",X"3F",X"3F",X"3E",X"23",X"76",X"38",X"7C",X"FC",X"FC",X"EC",X"67",X"27",X"47",
		X"00",X"00",X"01",X"02",X"02",X"02",X"04",X"05",X"1F",X"CF",X"27",X"13",X"13",X"09",X"C9",X"28",
		X"05",X"05",X"05",X"01",X"00",X"00",X"00",X"00",X"28",X"24",X"14",X"14",X"14",X"14",X"04",X"04",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"31",X"F8",X"E0",X"E2",X"C7",X"FF",X"FF",X"FF",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"1F",X"7F",X"FF",X"FF",X"FF",X"F3",X"31",X"FF",X"3F",X"FF",X"FF",X"FF",X"FF",X"DD",X"D0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"31",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DC",X"10",
		X"01",X"03",X"0E",X"0C",X"1C",X"38",X"F0",X"F8",X"F8",X"E0",X"00",X"07",X"1C",X"38",X"30",X"70",
		X"F0",X"FF",X"FF",X"FE",X"FF",X"DC",X"DF",X"CC",X"70",X"E0",X"80",X"00",X"00",X"0C",X"FF",X"E0",
		X"00",X"00",X"00",X"30",X"30",X"38",X"3B",X"3F",X"00",X"00",X"00",X"0C",X"0C",X"1C",X"9C",X"DC",
		X"3F",X"3F",X"3F",X"3F",X"3E",X"1E",X"1F",X"0F",X"8C",X"9C",X"9C",X"3C",X"3C",X"7C",X"F8",X"F8",
		X"16",X"1B",X"36",X"37",X"6F",X"6E",X"78",X"78",X"40",X"20",X"40",X"60",X"E4",X"EC",X"7C",X"7C",
		X"7C",X"3C",X"1C",X"1C",X"1C",X"00",X"00",X"00",X"3C",X"3C",X"3C",X"3C",X"3C",X"7C",X"7C",X"00",
		X"1F",X"3F",X"3F",X"3B",X"3D",X"3D",X"3C",X"3C",X"E4",X"C4",X"C8",X"EC",X"DC",X"77",X"7F",X"7F",
		X"7C",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"7E",X"78",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"27",X"6E",X"6E",X"7D",X"78",X"78",X"7C",X"6F",X"6F",X"FF",X"FB",X"00",X"00",X"00",X"00",
		X"3C",X"1C",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"60",X"F0",X"F0",X"78",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"7F",
		X"00",X"00",X"40",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"40",X"60",X"78",X"78",X"F0",X"F0",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"60",X"40",X"F8",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"0E",X"1F",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"05",X"07",X"07",X"0F",X"0F",X"E0",X"F7",X"FB",X"FB",
		X"0E",X"0F",X"1F",X"5F",X"DF",X"DF",X"BF",X"BF",X"00",X"04",X"AB",X"D7",X"E7",X"EF",X"EF",X"DF",
		X"BF",X"DF",X"C7",X"81",X"00",X"FC",X"FB",X"F7",X"DF",X"DF",X"BF",X"BF",X"7F",X"7F",X"FF",X"FF",
		X"07",X"07",X"03",X"7B",X"F9",X"FB",X"F7",X"F7",X"F8",X"F8",X"78",X"B0",X"80",X"A2",X"32",X"77",
		X"2F",X"07",X"0F",X"00",X"00",X"00",X"00",X"00",X"77",X"1F",X"0F",X"1F",X"1E",X"1C",X"1C",X"1C",
		X"06",X"04",X"02",X"06",X"27",X"37",X"3E",X"3E",X"68",X"D8",X"6C",X"EC",X"F6",X"76",X"1E",X"1E",
		X"3C",X"3C",X"3C",X"3C",X"3C",X"3E",X"3E",X"00",X"3E",X"3C",X"38",X"38",X"38",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"E0",
		X"60",X"60",X"E0",X"E0",X"E0",X"00",X"00",X"00",X"60",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"78",X"78",X"70",X"60",X"78",X"38",X"1C",X"0C",
		X"80",X"80",X"C0",X"C0",X"00",X"00",X"00",X"00",X"0F",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"1F",X"07",X"01",X"00",X"00",X"0F",X"7F",X"3F",X"DF",X"DF",X"9F",X"1F",X"BF",X"BF",X"BF",X"BF",
		X"9F",X"CF",X"E7",X"F2",X"F8",X"FC",X"FC",X"FC",X"C7",X"87",X"03",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C7",X"83",X"03",X"07",X"0F",X"10",X"00",X"00",X"00",X"00",
		X"83",X"83",X"C7",X"FF",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"80",X"00",X"00",X"00",X"00",X"00",X"FF",X"83",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"3F",X"00",X"00",X"00",X"00",X"01",X"7F",X"FF",X"E0",
		X"FF",X"FF",X"3F",X"0F",X"07",X"03",X"03",X"07",X"BF",X"9F",X"C7",X"F1",X"FC",X"FF",X"FF",X"FE",
		X"07",X"13",X"18",X"3E",X"FC",X"F0",X"80",X"00",X"FC",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"70",X"F8",X"00",X"00",X"00",X"00",X"02",X"07",X"07",X"17",
		X"00",X"00",X"00",X"01",X"03",X"03",X"07",X"07",X"37",X"67",X"EF",X"EF",X"EF",X"EF",X"EF",X"F3",
		X"01",X"03",X"07",X"0B",X"1D",X"3F",X"80",X"DF",X"FC",X"FC",X"FB",X"F7",X"F7",X"EF",X"0F",X"DF",
		X"EF",X"F7",X"FB",X"FD",X"FE",X"FC",X"FB",X"F7",X"DF",X"DF",X"BF",X"3F",X"7F",X"7F",X"FF",X"FF",
		X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"C1",X"E3",X"E7",X"F7",X"F7",X"FB",X"70",X"F0",X"F8",X"FA",X"FB",X"FB",X"FD",X"FD",
		X"FB",X"FB",X"FD",X"FD",X"FE",X"FE",X"FF",X"FF",X"FD",X"E3",X"81",X"00",X"00",X"3F",X"DF",X"EF",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"3F",X"3F",X"DF",X"EF",X"EF",X"F7",X"F0",X"FB",
		X"E0",X"E0",X"F0",X"F0",X"07",X"EF",X"DF",X"DF",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"A0",
		X"80",X"C0",X"E0",X"D0",X"B8",X"FC",X"01",X"FB",X"00",X"00",X"00",X"00",X"40",X"E0",X"E0",X"E8",
		X"FB",X"FB",X"FD",X"FD",X"FE",X"FE",X"FF",X"FF",X"F7",X"EF",X"DF",X"BF",X"7F",X"3F",X"DF",X"EF",
		X"FC",X"FC",X"FE",X"FF",X"F0",X"00",X"FF",X"FF",X"03",X"01",X"00",X"00",X"00",X"00",X"FC",X"FF",
		X"EC",X"EE",X"F7",X"F7",X"F7",X"F7",X"F7",X"CF",X"00",X"00",X"00",X"80",X"C0",X"C0",X"E0",X"E0",
		X"00",X"07",X"18",X"60",X"40",X"81",X"83",X"84",X"00",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",
		X"84",X"82",X"81",X"C0",X"60",X"78",X"3F",X"1F",X"7F",X"3F",X"FF",X"03",X"00",X"00",X"F0",X"F8",
		X"0F",X"0F",X"30",X"27",X"2F",X"2F",X"2F",X"2F",X"E1",X"C0",X"00",X"00",X"F8",X"FF",X"FF",X"FF",
		X"37",X"33",X"35",X"36",X"03",X"03",X"01",X"00",X"FF",X"FF",X"FC",X"00",X"E0",X"EF",X"FF",X"FF",
		X"F7",X"77",X"37",X"2F",X"0F",X"EF",X"CF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"DF",X"DF",X"1F",X"1F",X"BF",X"BF",X"BC",X"B8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"C0",X"80",X"80",X"80",X"9F",X"FF",X"FF",X"FF",X"03",X"01",X"00",X"01",X"F9",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"EF",X"EE",X"F1",X"F3",X"F7",X"F3",X"FB",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E3",X"C1",X"FB",X"F9",X"FA",X"FB",X"FD",X"FD",X"FD",X"FD",
		X"BF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"A0",X"B0",X"B0",X"78",X"78",X"7C",X"FC",X"3E",
		X"F8",X"E0",X"00",X"F0",X"FE",X"FF",X"F1",X"E0",X"1E",X"1E",X"0E",X"06",X"1E",X"1C",X"38",X"30",
		X"00",X"FF",X"01",X"01",X"01",X"F1",X"F1",X"F1",X"00",X"9F",X"91",X"D1",X"D1",X"F1",X"F1",X"F1",
		X"F1",X"F1",X"F1",X"F1",X"F1",X"71",X"31",X"31",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",
		X"00",X"9F",X"90",X"D0",X"D0",X"F1",X"F1",X"F1",X"00",X"FF",X"00",X"00",X"00",X"F1",X"F1",X"F1",
		X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",
		X"00",X"FF",X"30",X"30",X"30",X"F0",X"F0",X"F1",X"00",X"F1",X"0A",X"0A",X"04",X"00",X"00",X"80",
		X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"40",X"A0",X"91",X"9F",X"DF",X"DF",X"FF",X"FF",
		X"01",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"9F",X"CF",X"E7",X"F2",X"F8",X"FC",X"FC",X"FC",
		X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"FD",X"F7",X"EF",X"CF",X"9E",X"BE",X"3E",X"7F",
		X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"3F",X"7F",X"FF",X"07",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"03",X"00",X"00",X"00",X"00",X"80",X"F0",X"FC",X"FE",X"1F",X"03",X"01",X"00",
		X"87",X"C0",X"C0",X"C0",X"E0",X"00",X"00",X"00",X"E1",X"03",X"03",X"03",X"07",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C1",X"C3",X"00",X"07",X"1F",X"3F",X"7F",X"F0",X"E0",X"C0",
		X"C1",X"C1",X"E3",X"FF",X"F0",X"00",X"00",X"00",X"E7",X"E1",X"C0",X"00",X"00",X"00",X"00",X"3C",
		X"03",X"FF",X"FF",X"F6",X"80",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"3F",X"0F",X"07",X"07",X"07",
		X"CF",X"DF",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"70",X"00",X"80",X"80",X"80",X"C0",X"C0",X"E0",
		X"3F",X"87",X"C3",X"F1",X"F8",X"FF",X"FF",X"FE",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"31",X"00",X"F1",X"0A",X"0A",X"04",X"00",X"00",X"80",
		X"51",X"B1",X"31",X"31",X"71",X"71",X"F1",X"F1",X"40",X"20",X"11",X"1F",X"1F",X"1E",X"3F",X"3F",
		X"00",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"00",X"00",X"00",X"F8",X"F8",X"F8",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"F8",X"F8",X"F8",X"18",X"18",X"18",X"F8",X"F8",
		X"00",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"E0",X"18",X"06",X"02",X"81",X"C1",X"21",
		X"FE",X"FC",X"FF",X"00",X"00",X"00",X"FE",X"FE",X"21",X"41",X"81",X"02",X"06",X"38",X"20",X"20",
		X"E1",X"03",X"03",X"03",X"06",X"00",X"07",X"7F",X"7E",X"FC",X"39",X"03",X"00",X"00",X"00",X"00",
		X"05",X"0D",X"0D",X"1E",X"1E",X"3E",X"3F",X"7C",X"FD",X"FE",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",
		X"00",X"00",X"00",X"80",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",
		X"F7",X"F7",X"77",X"8F",X"CF",X"EF",X"CF",X"DF",X"EF",X"EE",X"EC",X"F4",X"F0",X"F7",X"F7",X"FB",
		X"46",X"0E",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"1F",X"00",
		X"81",X"00",X"00",X"00",X"1F",X"FF",X"FF",X"FF",X"F0",X"F0",X"14",X"EC",X"F4",X"F4",X"F4",X"F4",
		X"00",X"00",X"00",X"00",X"07",X"FF",X"FF",X"00",X"0F",X"03",X"1D",X"3E",X"FE",X"F8",X"C0",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"FB",X"F9",X"FA",X"FB",X"FD",X"FD",X"3D",X"1D",
		X"FC",X"F0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"C0",X"C0",X"E0",
		X"FF",X"FF",X"0F",X"F1",X"FE",X"FF",X"F1",X"E0",X"D4",X"BC",X"BC",X"6C",X"C0",X"C0",X"80",X"00",
		X"00",X"FF",X"01",X"01",X"01",X"01",X"01",X"31",X"00",X"3F",X"30",X"70",X"70",X"F1",X"F1",X"F1",
		X"51",X"B1",X"31",X"71",X"71",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F0",X"F0",X"F0",X"F1",X"F1",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"F8",X"F8",X"F8",X"F8",X"18",X"18",X"18",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"F8",X"00",
		X"FE",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"20",X"10",X"08",X"07",X"01",X"01",X"C1",X"FF",
		X"FF",X"FF",X"7F",X"7F",X"3F",X"3F",X"1F",X"00",X"FF",X"FE",X"FC",X"F8",X"F0",X"E0",X"C0",X"00",
		X"0F",X"07",X"03",X"FF",X"80",X"80",X"80",X"FF",X"FC",X"FC",X"F8",X"F0",X"00",X"00",X"03",X"FF",
		X"FF",X"7F",X"3F",X"1F",X"0F",X"07",X"03",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"31",X"30",X"30",X"30",X"78",X"F8",X"FC",X"FF",X"F1",X"E0",X"40",X"00",X"00",X"04",X"1F",X"FF",
		X"FF",X"FF",X"FF",X"FD",X"FC",X"F0",X"C0",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3E",X"00",
		X"F1",X"E1",X"41",X"01",X"03",X"03",X"07",X"FF",X"F1",X"F1",X"F1",X"F1",X"80",X"80",X"80",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"1E",X"00",X"FF",X"FF",X"FF",X"FF",X"BF",X"3F",X"1F",X"00",
		X"F1",X"F1",X"F1",X"F1",X"01",X"01",X"01",X"FF",X"FF",X"FF",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"00",
		X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"FF",X"7F",X"7B",X"03",X"03",X"03",X"03",X"03",X"03",
		X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"FC",X"00",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"00",
		X"F1",X"F1",X"F1",X"F1",X"F0",X"F0",X"F0",X"FF",X"F1",X"F1",X"F1",X"F1",X"00",X"00",X"00",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
