library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_OBJ_0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_OBJ_0 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",X"00",X"02",X"02",X"FE",X"FE",X"42",X"02",X"00",X"00",
		X"62",X"F2",X"BA",X"9A",X"9E",X"CE",X"46",X"00",X"8C",X"DE",X"F2",X"B2",X"92",X"86",X"04",X"00",
		X"08",X"FE",X"FE",X"C8",X"68",X"38",X"18",X"00",X"1C",X"BE",X"A2",X"A2",X"A2",X"E6",X"E4",X"00",
		X"0C",X"9E",X"92",X"92",X"D2",X"7E",X"3C",X"00",X"C0",X"E0",X"B0",X"9E",X"8E",X"C0",X"C0",X"00",
		X"0C",X"6E",X"9A",X"9A",X"B2",X"F2",X"6C",X"00",X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",X"00",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"00",X"70",X"F8",X"8D",X"85",X"C0",X"60",X"00",
		X"8E",X"4A",X"2E",X"10",X"E8",X"A4",X"E2",X"00",X"18",X"3C",X"7E",X"FF",X"3C",X"3C",X"3C",X"3C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",
		X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",X"44",X"C6",X"82",X"82",X"C6",X"7C",X"38",X"00",
		X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",X"82",X"92",X"92",X"92",X"FE",X"FE",X"00",X"00",
		X"80",X"90",X"90",X"90",X"90",X"FE",X"FE",X"00",X"9E",X"9E",X"92",X"82",X"C6",X"7C",X"38",X"00",
		X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",X"82",X"82",X"FE",X"FE",X"82",X"82",X"00",X"00",
		X"FC",X"FE",X"02",X"02",X"02",X"06",X"04",X"00",X"82",X"C6",X"6E",X"3C",X"18",X"FE",X"FE",X"00",
		X"02",X"02",X"02",X"02",X"FE",X"FE",X"00",X"00",X"FE",X"FE",X"70",X"38",X"70",X"FE",X"FE",X"00",
		X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",X"00",
		X"70",X"F8",X"88",X"88",X"88",X"FE",X"FE",X"00",X"7A",X"FC",X"8E",X"8A",X"82",X"FE",X"7C",X"00",
		X"72",X"F6",X"9E",X"8C",X"88",X"FE",X"FE",X"00",X"0C",X"5E",X"D2",X"92",X"92",X"F6",X"64",X"00",
		X"80",X"80",X"FE",X"FE",X"80",X"80",X"00",X"00",X"FC",X"FE",X"02",X"02",X"02",X"FE",X"FC",X"00",
		X"F0",X"F8",X"1C",X"0E",X"1C",X"F8",X"F0",X"00",X"F8",X"FE",X"1C",X"38",X"1C",X"FE",X"F8",X"00",
		X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",X"C0",X"F0",X"1E",X"1E",X"F0",X"C0",X"00",X"00",
		X"C2",X"E2",X"F2",X"BA",X"9E",X"8E",X"86",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",
		X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"03",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"15",X"06",X"03",X"00",X"01",X"00",X"00",X"00",X"50",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"16",X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"C0",
		X"05",X"06",X"03",X"00",X"02",X"00",X"00",X"00",X"40",X"D0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"13",X"06",X"00",X"00",X"00",X"00",X"40",X"00",X"80",X"C0",
		X"05",X"06",X"03",X"00",X"04",X"00",X"00",X"00",X"40",X"C0",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"03",X"06",X"00",X"00",X"00",X"00",X"00",X"20",X"80",X"C0",
		X"05",X"06",X"03",X"08",X"00",X"00",X"00",X"00",X"40",X"C0",X"80",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",
		X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"00",
		X"00",X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"00",X"00",X"00",X"78",X"00",X"00",X"04",X"96",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"78",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"0C",X"03",X"00",X"00",X"00",X"00",X"00",X"20",X"18",X"08",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"C0",X"10",X"0C",X"86",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"04",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"08",
		X"00",X"00",X"00",X"02",X"01",X"00",X"00",X"00",X"84",X"00",X"20",X"10",X"08",X"80",X"00",X"00",
		X"00",X"00",X"00",X"04",X"02",X"02",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",
		X"00",X"00",X"00",X"06",X"03",X"00",X"00",X"00",X"98",X"88",X"00",X"40",X"20",X"10",X"00",X"00",
		X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"10",X"10",X"11",X"11",X"01",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"00",X"00",X"00",X"78",X"00",X"00",X"00",X"9C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"78",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"0C",X"03",X"00",X"00",X"00",X"00",X"00",X"20",X"18",X"08",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"C0",X"10",X"10",X"8C",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"04",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"08",
		X"00",X"00",X"00",X"02",X"01",X"00",X"00",X"00",X"84",X"00",X"30",X"28",X"10",X"84",X"00",X"00",
		X"00",X"00",X"00",X"04",X"02",X"02",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",
		X"00",X"00",X"00",X"06",X"03",X"00",X"00",X"00",X"98",X"88",X"00",X"60",X"10",X"30",X"10",X"00",
		X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"10",X"10",X"11",X"12",X"01",X"01",X"00",X"00",X"10",X"10",X"10",X"10",X"80",X"00",X"00",
		X"03",X"05",X"08",X"08",X"04",X"03",X"05",X"09",X"80",X"40",X"20",X"20",X"40",X"80",X"40",X"20",
		X"5A",X"AC",X"5A",X"A9",X"0A",X"0C",X"08",X"1C",X"AA",X"74",X"AA",X"34",X"A0",X"60",X"10",X"38",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"00",
		X"00",X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"08",X"10",X"20",X"20",X"21",X"00",X"00",X"C0",X"00",X"00",X"00",X"10",X"10",
		X"21",X"00",X"04",X"03",X"00",X"00",X"00",X"00",X"10",X"10",X"20",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"3E",X"51",X"60",X"8F",X"90",X"A0",X"C0",X"00",X"18",X"20",X"A0",X"40",X"C0",X"44",X"28",
		X"4C",X"52",X"52",X"2C",X"10",X"0F",X"00",X"00",X"20",X"20",X"20",X"40",X"80",X"00",X"00",X"00",
		X"20",X"07",X"89",X"11",X"11",X"10",X"08",X"07",X"78",X"84",X"00",X"18",X"28",X"30",X"00",X"00",
		X"60",X"80",X"88",X"18",X"30",X"00",X"00",X"00",X"00",X"00",X"04",X"0A",X"04",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"08",X"14",X"08",X"00",X"1C",X"22",X"41",X"49",X"41",X"22",X"1C",X"00",
		X"00",X"00",X"30",X"48",X"48",X"30",X"00",X"00",X"00",X"00",X"38",X"44",X"54",X"44",X"38",X"02",
		X"00",X"1C",X"22",X"41",X"41",X"41",X"22",X"1C",X"00",X"00",X"0E",X"11",X"11",X"11",X"0E",X"00",
		X"00",X"00",X"00",X"31",X"49",X"49",X"30",X"00",X"00",X"70",X"88",X"04",X"04",X"04",X"88",X"70",
		X"00",X"04",X"0A",X"04",X"38",X"44",X"82",X"82",X"00",X"00",X"00",X"38",X"44",X"82",X"92",X"82",
		X"82",X"44",X"38",X"44",X"44",X"44",X"38",X"00",X"44",X"38",X"00",X"0C",X"12",X"12",X"0C",X"00",
		X"00",X"00",X"04",X"0A",X"04",X"20",X"00",X"00",X"02",X"05",X"02",X"00",X"20",X"50",X"20",X"00",
		X"00",X"00",X"00",X"06",X"09",X"09",X"06",X"00",X"00",X"08",X"14",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"14",X"08",X"00",X"38",X"44",X"00",X"60",X"90",X"90",X"60",X"00",X"38",X"44",
		X"44",X"44",X"38",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"04",X"08",X"11",X"00",X"00",X"00",X"00",X"00",X"40",X"20",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"07",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"60",
		X"04",X"04",X"04",X"04",X"00",X"00",X"00",X"00",X"10",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"07",X"06",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",
		X"02",X"02",X"02",X"02",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"02",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0F",X"00",X"00",X"00",X"20",X"40",X"80",X"00",X"20",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"02",X"02",X"00",X"01",X"01",X"01",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",
		X"02",X"04",X"05",X"05",X"05",X"15",X"15",X"10",X"80",X"40",X"40",X"40",X"40",X"50",X"50",X"10",
		X"00",X"00",X"00",X"02",X"03",X"02",X"00",X"09",X"00",X"00",X"00",X"80",X"80",X"80",X"00",X"20",
		X"02",X"04",X"01",X"08",X"00",X"00",X"00",X"00",X"80",X"40",X"00",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"0F",X"00",X"00",X"00",X"00",X"C0",X"E0",X"60",X"00",
		X"21",X"05",X"01",X"00",X"02",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"02",X"02",X"00",X"01",X"01",X"01",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",
		X"02",X"04",X"05",X"04",X"04",X"10",X"10",X"00",X"80",X"40",X"40",X"40",X"40",X"10",X"10",X"00",
		X"01",X"01",X"02",X"02",X"00",X"01",X"01",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",
		X"01",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"19",X"21",X"41",X"01",X"01",X"7C",X"01",X"00",X"48",X"44",X"42",X"42",X"40",X"00",X"BE",
		X"7D",X"00",X"02",X"42",X"42",X"22",X"12",X"00",X"80",X"3E",X"80",X"80",X"82",X"84",X"98",X"00",
		X"00",X"02",X"0A",X"4A",X"45",X"85",X"84",X"01",X"60",X"18",X"00",X"00",X"0C",X"70",X"0E",X"B0",
		X"0D",X"70",X"0E",X"30",X"00",X"00",X"18",X"06",X"80",X"21",X"A1",X"A2",X"52",X"50",X"40",X"00",
		X"07",X"00",X"10",X"28",X"14",X"8A",X"84",X"81",X"E0",X"00",X"08",X"14",X"28",X"51",X"21",X"81",
		X"81",X"84",X"8A",X"14",X"28",X"10",X"00",X"07",X"81",X"A1",X"51",X"28",X"14",X"08",X"00",X"E0",
		X"00",X"00",X"20",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",
		X"00",X"40",X"02",X"00",X"00",X"00",X"20",X"00",X"00",X"08",X"00",X"00",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"10",X"02",X"01",X"06",X"00",X"10",X"00",X"02",X"80",X"70",X"50",X"D0",
		X"A3",X"15",X"07",X"02",X"10",X"02",X"00",X"00",X"B0",X"60",X"E2",X"80",X"90",X"02",X"80",X"10",
		X"00",X"00",X"00",X"00",X"0A",X"0C",X"01",X"20",X"00",X"00",X"00",X"00",X"80",X"00",X"40",X"80",
		X"09",X"14",X"2A",X"00",X"05",X"06",X"00",X"00",X"40",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"18",X"20",X"40",X"43",X"84",X"89",X"8A",X"E0",X"18",X"04",X"02",X"C2",X"21",X"91",X"51",
		X"8A",X"89",X"84",X"43",X"40",X"20",X"18",X"07",X"51",X"91",X"21",X"C2",X"02",X"04",X"18",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"00",X"00",X"00",X"78",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"78",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"0C",X"03",X"00",X"00",X"00",X"00",X"00",X"20",X"18",X"08",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"80",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"04",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"08",
		X"00",X"00",X"00",X"02",X"01",X"00",X"00",X"00",X"84",X"00",X"00",X"00",X"00",X"80",X"00",X"00",
		X"00",X"00",X"00",X"04",X"02",X"02",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",
		X"00",X"00",X"00",X"06",X"03",X"00",X"00",X"00",X"98",X"88",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"10",X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
