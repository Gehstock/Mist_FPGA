library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity obj4 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of obj4 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"C1",X"C0",X"C0",X"C1",X"61",X"01",
		X"00",X"00",X"00",X"06",X"0B",X"01",X"01",X"01",X"00",X"C1",X"C3",X"E0",X"E4",X"7C",X"3C",X"1D",
		X"00",X"00",X"00",X"00",X"00",X"18",X"0C",X"1C",X"1C",X"10",X"06",X"01",X"01",X"09",X"04",X"20",
		X"00",X"00",X"00",X"00",X"0C",X"0C",X"04",X"06",X"02",X"00",X"20",X"10",X"B0",X"F8",X"FC",X"BC",
		X"00",X"00",X"00",X"00",X"00",X"80",X"44",X"C6",X"02",X"03",X"01",X"60",X"E0",X"A0",X"A0",X"50",
		X"00",X"00",X"00",X"0C",X"06",X"0F",X"0F",X"04",X"00",X"10",X"B8",X"F8",X"FC",X"AE",X"A6",X"AA",
		X"00",X"00",X"00",X"0C",X"06",X"0F",X"0F",X"04",X"00",X"10",X"B8",X"F8",X"FC",X"AE",X"A6",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"30",X"98",X"9C",X"9E",X"8E",X"8F",X"8F",X"83",X"80",X"90",X"00",X"20",X"40",
		X"00",X"00",X"00",X"30",X"98",X"9C",X"9E",X"8E",X"8F",X"8F",X"83",X"80",X"88",X"08",X"10",X"80",
		X"00",X"06",X"07",X"03",X"C1",X"C0",X"C0",X"00",X"40",X"00",X"00",X"00",X"1C",X"3C",X"00",X"00",
		X"00",X"06",X"07",X"03",X"C1",X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",X"C0",X"FC",X"FC",X"E0",X"C0",
		X"1E",X"1C",X"00",X"00",X"C0",X"C0",X"E0",X"E3",X"C3",X"A3",X"81",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"1C",X"00",X"00",X"C0",X"C0",X"E0",X"E3",X"E3",X"63",X"E1",X"60",X"60",X"E0",X"E0",X"C0",
		X"06",X"0A",X"92",X"80",X"70",X"E0",X"70",X"30",X"38",X"38",X"7C",X"FC",X"FC",X"9C",X"C8",X"D8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"08",X"10",X"F1",
		X"00",X"00",X"00",X"00",X"03",X"07",X"03",X"01",X"11",X"08",X"0C",X"0E",X"1E",X"BE",X"FE",X"FE",
		X"00",X"00",X"00",X"00",X"10",X"D8",X"2C",X"FE",X"2C",X"D8",X"10",X"00",X"00",X"00",X"00",X"00",
		X"08",X"18",X"B8",X"F8",X"F0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"18",X"10",
		X"80",X"A0",X"A0",X"B0",X"E0",X"C0",X"00",X"20",X"10",X"08",X"A0",X"A0",X"28",X"08",X"18",X"10",
		X"03",X"E7",X"FD",X"F8",X"F8",X"F0",X"F3",X"E7",X"FD",X"FC",X"E0",X"80",X"0C",X"1C",X"1C",X"00",
		X"00",X"30",X"18",X"1C",X"1C",X"3C",X"3C",X"38",X"3C",X"3C",X"1C",X"C0",X"E0",X"C0",X"00",X"00",
		X"00",X"18",X"3C",X"1C",X"0C",X"00",X"CC",X"6E",X"3E",X"BE",X"7A",X"61",X"61",X"01",X"1A",X"04",
		X"00",X"38",X"3C",X"1C",X"1C",X"1E",X"1C",X"1C",X"1C",X"1C",X"3C",X"18",X"00",X"00",X"80",X"80",
		X"00",X"1C",X"3C",X"FC",X"FC",X"3E",X"1E",X"1E",X"0E",X"04",X"08",X"0C",X"0C",X"0C",X"00",X"00",
		X"00",X"18",X"3C",X"FC",X"3C",X"1C",X"1C",X"1C",X"3E",X"3E",X"3C",X"0C",X"00",X"80",X"C0",X"C0",
		X"00",X"00",X"00",X"78",X"FC",X"F8",X"F8",X"F0",X"00",X"00",X"C0",X"E0",X"E0",X"E0",X"E0",X"00",
		X"00",X"60",X"70",X"30",X"B8",X"F8",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"E0",X"80",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F0",X"98",X"E8",X"F4",X"FC",X"FC",X"FC",X"F8",X"F8",X"F0",X"00",X"00",X"00",
		X"E0",X"F0",X"A0",X"F0",X"90",X"32",X"93",X"21",X"20",X"70",X"F0",X"F8",X"F8",X"F0",X"30",X"00",
		X"00",X"00",X"00",X"10",X"7C",X"FC",X"F8",X"78",X"78",X"FC",X"F8",X"78",X"10",X"00",X"00",X"00",
		X"70",X"F0",X"EC",X"DC",X"DE",X"DE",X"DE",X"5E",X"5E",X"5E",X"DE",X"DE",X"DE",X"DC",X"EC",X"F0",
		X"70",X"E8",X"FC",X"EC",X"C6",X"EE",X"FE",X"6E",X"46",X"6E",X"FE",X"EE",X"C6",X"EC",X"FC",X"E8",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"80",X"C0",X"80",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"18",X"08",X"38",X"38",X"18",X"18",X"30",X"18",X"30",X"38",X"10",X"08",
		X"02",X"04",X"EE",X"0C",X"06",X"0C",X"06",X"06",X"0E",X"0A",X"06",X"00",X"00",X"00",X"00",X"00",
		X"10",X"30",X"70",X"70",X"30",X"70",X"50",X"30",X"30",X"70",X"50",X"30",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"E0",X"E0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F4",X"F0",X"F0",X"28",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"80",X"00",X"00",X"00",X"00",X"00",
		X"E1",X"00",X"00",X"00",X"00",X"C0",X"60",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"60",X"20",X"20",X"31",X"38",X"35",X"1F",X"1E",
		X"00",X"00",X"00",X"00",X"03",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"60",X"B0",X"40",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"40",X"00",X"40",X"00",X"00",X"40",X"00",X"40",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"FF",X"03",X"83",X"03",X"83",X"03",X"03",X"83",X"03",X"83",X"23",X"13",X"0B",X"07",X"FE",X"FC",
		X"FC",X"FE",X"07",X"0B",X"13",X"0B",X"0B",X"23",X"03",X"23",X"03",X"03",X"23",X"03",X"23",X"FF",
		X"60",X"F0",X"F8",X"FC",X"FC",X"FE",X"FC",X"EC",X"CE",X"CE",X"C0",X"C0",X"E0",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"72",X"F9",X"FE",X"FF",X"6F",X"9F",X"DF",X"5F",
		X"5F",X"5F",X"6F",X"27",X"0F",X"07",X"00",X"00",X"00",X"00",X"40",X"80",X"00",X"00",X"00",X"00",
		X"03",X"07",X"06",X"0A",X"0C",X"0C",X"08",X"10",X"18",X"14",X"10",X"38",X"30",X"20",X"20",X"60",
		X"50",X"40",X"C0",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"18",X"30",X"F6",X"F7",X"F7",X"F3",X"FB",X"F9",X"FC",X"E4",X"C2",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"30",X"70",X"F0",X"F0",X"E0",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"49",X"2A",X"08",X"7E",X"08",X"2A",X"49",X"80",X"00",X"02",X"09",X"80",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"30",X"78",X"70",X"F0",X"70",X"78",X"30",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"80",X"80",X"80",X"00",X"C0",X"70",X"60",X"60",X"C0",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"80",X"80",X"80",X"80",X"00",X"80",X"60",X"00",X"80",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"14",X"D0",X"4C",X"C4",X"14",X"10",X"24",X"28",X"44",X"48",X"04",
		X"00",X"00",X"00",X"00",X"00",X"14",X"10",X"CC",X"44",X"C8",X"04",X"08",X"04",X"08",X"04",X"0C",
		X"00",X"08",X"A0",X"80",X"C8",X"E0",X"60",X"FC",X"60",X"E4",X"C0",X"90",X"80",X"08",X"40",X"00",
		X"00",X"00",X"80",X"00",X"00",X"80",X"40",X"C0",X"40",X"80",X"00",X"00",X"20",X"00",X"00",X"00",
		X"00",X"C8",X"20",X"10",X"88",X"C4",X"64",X"E4",X"E4",X"64",X"C4",X"88",X"10",X"24",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"82",X"C0",X"60",X"E0",X"E0",X"60",X"C0",X"80",X"00",X"00",X"00",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"F0",X"00",X"00",X"80",X"E0",X"C0",X"00",X"00",X"00",X"E0",X"00",X"00",X"80",X"F0",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"01",X"00",X"F0",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"06",X"0E",X"0E",X"1C",X"1A",X"1A",X"1C",X"0E",X"0E",X"06",X"00",X"00",X"00",X"0E",X"0E",
		X"00",X"06",X"0E",X"0E",X"1C",X"1A",X"1A",X"1C",X"0E",X"0E",X"86",X"80",X"80",X"00",X"00",X"00",
		X"01",X"DF",X"5F",X"5F",X"5F",X"DF",X"5F",X"5F",X"DF",X"5F",X"5F",X"5F",X"DF",X"FF",X"DF",X"01",
		X"00",X"01",X"01",X"81",X"C0",X"00",X"60",X"64",X"64",X"60",X"00",X"C0",X"81",X"01",X"01",X"00",
		X"60",X"70",X"70",X"70",X"70",X"F0",X"70",X"70",X"70",X"F0",X"70",X"70",X"F0",X"70",X"70",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"20",X"60",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"10",X"60",X"80",X"00",X"60",X"10",X"8C",X"80",X"80",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"56",X"AA",X"00",X"00",X"C0",X"40",X"40",X"40",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"80",X"C0",X"F0",X"38",X"0C",X"74",X"74",X"0C",X"38",X"F0",X"C0",X"80",X"00",X"00",
		X"00",X"60",X"F0",X"F0",X"98",X"08",X"0C",X"94",X"94",X"0C",X"08",X"98",X"F0",X"F0",X"60",X"00",
		X"18",X"18",X"18",X"18",X"3C",X"24",X"24",X"24",X"24",X"24",X"24",X"3C",X"18",X"18",X"18",X"18",
		X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"00",X"00",X"04",X"04",X"04",X"04",X"04",X"04",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"1B",X"38",X"20",X"40",X"80",X"00",X"00",X"00",X"80",
		X"80",X"C0",X"C0",X"E0",X"F0",X"F9",X"BD",X"AF",X"AF",X"AB",X"EB",X"FB",X"EB",X"FF",X"EF",X"FF",
		X"EF",X"FF",X"EE",X"FE",X"FC",X"FC",X"F8",X"78",X"F0",X"F0",X"80",X"E0",X"F0",X"F0",X"E0",X"C0",
		X"00",X"00",X"80",X"40",X"20",X"22",X"35",X"38",X"35",X"22",X"20",X"E0",X"E0",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"E0",X"E0",X"20",X"22",X"35",X"38",X"35",X"22",X"20",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"1B",X"38",X"20",X"40",X"80",X"00",X"00",X"00",X"80",
		X"80",X"C0",X"C0",X"E0",X"F0",X"F9",X"BD",X"AF",X"AF",X"AB",X"EB",X"FB",X"EB",X"FF",X"EF",X"FF",
		X"EF",X"FF",X"EE",X"FE",X"E4",X"E8",X"E8",X"DC",X"DE",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"12",X"01",X"81",X"C9",X"25",X"05",X"C5",X"05",X"05",X"35",X"E5",X"C9",X"81",X"12",X"0C",
		X"00",X"08",X"00",X"44",X"CA",X"02",X"02",X"02",X"00",X"02",X"40",X"02",X"0A",X"04",X"20",X"00",
		X"00",X"00",X"E0",X"10",X"08",X"08",X"54",X"F4",X"F4",X"04",X"08",X"08",X"10",X"E0",X"00",X"00",
		X"00",X"00",X"C0",X"20",X"10",X"08",X"08",X"08",X"08",X"08",X"08",X"10",X"20",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"40",X"20",X"20",X"20",X"20",X"40",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"04",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"04",X"80",
		X"0C",X"01",X"03",X"C1",X"76",X"20",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"19",X"08",X"08",X"81",X"81",X"41",X"04",X"05",X"03",X"06",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"61",X"60",X"E0",X"B1",X"B9",X"B1",X"E0",X"80",X"80",X"05",X"07",X"03",X"06",X"00",X"00",
		X"AC",X"A4",X"5C",X"F8",X"F0",X"C0",X"01",X"01",X"13",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"59",X"5F",X"7F",X"FF",X"C6",X"86",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"BE",X"FC",X"F8",X"B8",X"10",X"00",X"04",X"0F",X"0F",X"06",X"0C",X"00",X"00",X"00",X"00",
		X"AA",X"BE",X"FC",X"F8",X"B8",X"10",X"00",X"04",X"0F",X"0F",X"06",X"0C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"C0",X"C0",X"01",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"06",X"02",X"86",X"40",X"58",X"BC",X"AE",X"A6",
		X"AA",X"AA",X"BC",X"58",X"40",X"80",X"00",X"02",X"06",X"0C",X"18",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"5E",X"3F",X"18",X"7A",X"F6",X"04",X"3E",X"12",X"21",X"70",X"F8",X"F8",X"F8",X"FF",X"FF",X"73",
		X"50",X"72",X"46",X"8E",X"9C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"A1",X"A1",X"B1",X"BC",X"70",X"E2",X"00",X"00",X"02",X"02",X"00",X"00",X"00",X"00",
		X"CE",X"CC",X"CD",X"DC",X"DD",X"F8",X"F1",X"C1",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"C0",X"E0",X"F0",X"F0",X"F0",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"81",X"B8",X"BC",X"AE",X"A6",
		X"AA",X"AA",X"BC",X"BA",X"83",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"06",X"02",X"86",X"40",X"58",X"BC",X"AE",X"A6",
		X"C0",X"20",X"20",X"20",X"C0",X"00",X"C0",X"20",X"20",X"20",X"C0",X"00",X"20",X"E0",X"20",X"00",
		X"C0",X"20",X"20",X"C0",X"00",X"C0",X"20",X"20",X"C0",X"00",X"20",X"20",X"A0",X"60",X"20",X"00",
		X"C0",X"20",X"20",X"C0",X"00",X"C0",X"20",X"20",X"C0",X"00",X"C0",X"20",X"20",X"20",X"20",X"00",
		X"C0",X"20",X"20",X"20",X"C0",X"00",X"C0",X"20",X"20",X"20",X"C0",X"00",X"E0",X"40",X"40",X"C0",
		X"C0",X"20",X"20",X"C0",X"00",X"C0",X"20",X"20",X"C0",X"00",X"C0",X"20",X"20",X"20",X"C0",X"00",
		X"C0",X"20",X"C0",X"00",X"C0",X"20",X"C0",X"00",X"20",X"20",X"A0",X"60",X"00",X"E0",X"00",X"00",
		X"C0",X"20",X"C0",X"00",X"C0",X"20",X"C0",X"00",X"C0",X"20",X"20",X"C0",X"00",X"E0",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
