library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity exerion_04 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of exerion_04 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"F3",
		X"00",X"0F",X"00",X"00",X"00",X"61",X"00",X"2C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"8E",X"F1",
		X"00",X"01",X"01",X"00",X"08",X"E1",X"00",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"8C",X"FF",X"F0",
		X"00",X"01",X"02",X"08",X"09",X"E1",X"90",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"0C",X"EF",X"FF",X"FB",
		X"80",X"70",X"04",X"48",X"6F",X"E7",X"D2",X"3E",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"8C",X"F1",X"F8",
		X"C0",X"F0",X"04",X"68",X"6F",X"EF",X"D2",X"3F",X"00",X"CC",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E8",
		X"E8",X"F7",X"14",X"78",X"09",X"EF",X"DF",X"3F",X"00",X"EE",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"F9",
		X"EC",X"FF",X"1E",X"7E",X"09",X"EF",X"DF",X"3F",X"00",X"EE",X"13",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"F3",X"FE",X"F9",X"FF",
		X"EE",X"FF",X"1F",X"7F",X"09",X"EF",X"DF",X"3F",X"00",X"FF",X"13",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"08",X"EF",X"F8",X"FF",X"F1",X"FE",
		X"EE",X"FF",X"15",X"7F",X"09",X"EF",X"DF",X"3F",X"00",X"FF",X"13",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"08",X"FF",X"F1",X"F7",X"F0",X"F8",X"FF",
		X"CC",X"FF",X"04",X"6E",X"6F",X"EF",X"DF",X"3F",X"88",X"FF",X"13",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"CC",X"FF",X"F7",X"FC",X"F0",X"FC",
		X"88",X"77",X"04",X"4C",X"6F",X"EF",X"DF",X"3F",X"88",X"FF",X"37",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"48",X"FF",X"FF",X"F7",X"FC",
		X"00",X"01",X"02",X"08",X"09",X"EF",X"99",X"3F",X"88",X"FF",X"37",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"FC",X"F7",X"FC",
		X"00",X"01",X"01",X"00",X"00",X"88",X"00",X"3F",X"88",X"FF",X"37",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"EE",X"FF",X"11",X"F0",X"00",X"00",X"00",X"00",X"F0",X"F8",X"FF",X"FD",
		X"00",X"0F",X"00",X"80",X"F0",X"70",X"00",X"26",X"88",X"FF",X"37",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"EE",X"CC",X"FF",X"FF",X"33",X"F0",X"00",X"00",X"80",X"FF",X"F0",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"E0",X"F0",X"5A",X"10",X"08",X"88",X"FF",X"37",X"00",X"00",X"00",X"00",X"00",
		X"00",X"88",X"FF",X"FE",X"FF",X"FF",X"FB",X"F1",X"00",X"00",X"FE",X"F6",X"F8",X"FE",X"BE",X"BF",
		X"00",X"00",X"00",X"F0",X"F0",X"5A",X"30",X"0F",X"08",X"FF",X"37",X"00",X"00",X"CC",X"11",X"00",
		X"00",X"CC",X"FF",X"FC",X"F7",X"FF",X"FB",X"F1",X"8E",X"FF",X"FF",X"F3",X"D3",X"FE",X"FE",X"FF",
		X"00",X"00",X"80",X"F0",X"F0",X"78",X"78",X"0F",X"00",X"6F",X"37",X"00",X"00",X"EE",X"13",X"00",
		X"00",X"EE",X"FF",X"FC",X"F7",X"FE",X"FB",X"F1",X"00",X"00",X"84",X"F2",X"D7",X"FF",X"FE",X"FF",
		X"00",X"00",X"C0",X"F8",X"FF",X"5F",X"F0",X"01",X"00",X"8E",X"71",X"00",X"00",X"EE",X"13",X"00",
		X"00",X"EE",X"FF",X"FF",X"F1",X"FE",X"FB",X"F1",X"00",X"00",X"00",X"C0",X"F7",X"FF",X"D7",X"F7",
		X"00",X"00",X"C0",X"FE",X"FF",X"5F",X"F1",X"00",X"00",X"CC",X"F7",X"00",X"00",X"FF",X"37",X"00",
		X"00",X"FF",X"FF",X"F3",X"F0",X"FF",X"FB",X"F1",X"00",X"00",X"C8",X"F7",X"F7",X"F7",X"1F",X"B7",
		X"00",X"00",X"E8",X"FF",X"FF",X"7F",X"F3",X"10",X"00",X"EE",X"F7",X"00",X"00",X"FF",X"37",X"00",
		X"00",X"FF",X"FF",X"F0",X"10",X"00",X"EA",X"F1",X"08",X"ED",X"F7",X"FC",X"F7",X"F7",X"5B",X"E7",
		X"00",X"00",X"EC",X"FF",X"FF",X"5F",X"F7",X"10",X"00",X"FF",X"FF",X"10",X"88",X"FF",X"37",X"00",
		X"00",X"77",X"88",X"10",X"EE",X"FF",X"D9",X"F1",X"87",X"F0",X"F4",X"FD",X"FD",X"F5",X"F3",X"F6",
		X"00",X"00",X"EE",X"FF",X"FF",X"5F",X"FF",X"18",X"00",X"FF",X"FF",X"31",X"88",X"FF",X"37",X"00",
		X"00",X"88",X"77",X"EE",X"FF",X"FF",X"FB",X"F1",X"00",X"80",X"FC",X"F8",X"F9",X"F1",X"F3",X"F6",
		X"00",X"00",X"EE",X"FF",X"FF",X"7F",X"FF",X"1F",X"88",X"FF",X"FF",X"31",X"88",X"FF",X"37",X"00",
		X"00",X"FF",X"F7",X"FF",X"FF",X"FF",X"33",X"F0",X"00",X"00",X"80",X"F7",X"F9",X"B5",X"E3",X"F4",
		X"00",X"00",X"EE",X"FF",X"FF",X"5F",X"FF",X"1F",X"88",X"FF",X"FF",X"31",X"88",X"FF",X"37",X"00",
		X"88",X"FF",X"F7",X"FF",X"F7",X"FF",X"F7",X"F7",X"00",X"00",X"00",X"80",X"EB",X"F3",X"F4",X"F4",
		X"00",X"00",X"EE",X"FF",X"FF",X"5F",X"FF",X"19",X"88",X"FF",X"7F",X"01",X"88",X"FF",X"B7",X"00",
		X"CC",X"FF",X"F7",X"FC",X"F7",X"FE",X"F7",X"FF",X"00",X"00",X"88",X"7F",X"EB",X"FB",X"FC",X"B4",
		X"00",X"00",X"EE",X"FF",X"FF",X"7F",X"FF",X"11",X"88",X"FF",X"FF",X"03",X"88",X"FF",X"C7",X"00",
		X"EE",X"FF",X"F7",X"FE",X"F1",X"FE",X"F7",X"FF",X"00",X"84",X"F6",X"F3",X"EF",X"FB",X"FC",X"B7",
		X"00",X"00",X"EE",X"FF",X"FF",X"5F",X"FF",X"11",X"88",X"FF",X"FF",X"13",X"88",X"FF",X"F7",X"00",
		X"FF",X"FF",X"FF",X"F7",X"F0",X"FE",X"F7",X"FF",X"0C",X"ED",X"F7",X"F0",X"EF",X"BF",X"9F",X"E7",
		X"00",X"00",X"CC",X"FF",X"FF",X"5F",X"FF",X"00",X"88",X"FF",X"FF",X"13",X"88",X"FF",X"F7",X"00",
		X"FF",X"FF",X"FF",X"F1",X"FC",X"FF",X"F7",X"FF",X"00",X"80",X"F0",X"F7",X"F0",X"FB",X"9F",X"6F",
		X"00",X"00",X"CC",X"FF",X"FF",X"7F",X"FF",X"01",X"88",X"FF",X"FF",X"13",X"00",X"FF",X"FF",X"10",
		X"FF",X"FF",X"F7",X"F0",X"FE",X"FF",X"F7",X"FF",X"00",X"00",X"08",X"F0",X"F0",X"F9",X"3F",X"6B",
		X"00",X"00",X"88",X"FF",X"FF",X"5F",X"7F",X"0F",X"00",X"FF",X"FF",X"13",X"00",X"FF",X"FF",X"10",
		X"FF",X"FF",X"F7",X"FC",X"FF",X"FF",X"F7",X"FF",X"00",X"00",X"00",X"00",X"80",X"F8",X"7B",X"3F",
		X"00",X"00",X"00",X"FF",X"FF",X"5F",X"33",X"0F",X"00",X"66",X"FF",X"13",X"00",X"EE",X"FF",X"10",
		X"FF",X"FF",X"F7",X"FE",X"FF",X"FF",X"F7",X"FF",X"00",X"00",X"00",X"08",X"87",X"BE",X"F9",X"F1",
		X"00",X"00",X"00",X"EE",X"FF",X"00",X"00",X"08",X"00",X"80",X"FF",X"13",X"00",X"04",X"FF",X"10",
		X"FF",X"FF",X"F7",X"FE",X"FF",X"FF",X"F7",X"FF",X"00",X"00",X"08",X"87",X"F7",X"9F",X"BF",X"97",
		X"00",X"00",X"00",X"88",X"77",X"F0",X"70",X"0E",X"00",X"88",X"FF",X"13",X"00",X"4C",X"CC",X"10",
		X"CF",X"FF",X"F7",X"FF",X"FF",X"FF",X"B7",X"FF",X"00",X"00",X"87",X"F0",X"FE",X"1F",X"1F",X"C7",
		X"00",X"00",X"00",X"00",X"08",X"F0",X"69",X"0F",X"00",X"88",X"FF",X"01",X"00",X"CC",X"CF",X"10",
		X"8F",X"FF",X"B7",X"FF",X"FF",X"FF",X"97",X"6F",X"00",X"00",X"08",X"C3",X"F8",X"DF",X"3E",X"CF",
		X"00",X"00",X"00",X"00",X"48",X"F0",X"69",X"01",X"00",X"08",X"7F",X"01",X"00",X"CC",X"FF",X"10",
		X"0F",X"EF",X"97",X"EF",X"FF",X"FF",X"4B",X"0F",X"00",X"00",X"00",X"0C",X"C0",X"F8",X"96",X"ED",
		X"00",X"00",X"00",X"00",X"68",X"F0",X"78",X"00",X"00",X"00",X"0F",X"01",X"00",X"88",X"FF",X"10",
		X"0E",X"0F",X"0F",X"8F",X"FF",X"3F",X"69",X"0F",X"00",X"00",X"00",X"00",X"00",X"C0",X"D2",X"F8",
		X"00",X"00",X"00",X"00",X"69",X"FF",X"6F",X"00",X"00",X"00",X"0C",X"00",X"00",X"88",X"FF",X"10",
		X"0E",X"0F",X"0F",X"0F",X"EF",X"0F",X"2D",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",
		X"00",X"00",X"00",X"80",X"6F",X"FF",X"6F",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"10",
		X"0C",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"87",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",
		X"00",X"00",X"00",X"C0",X"6F",X"FF",X"7F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"F7",X"00",
		X"08",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"FC",
		X"00",X"00",X"00",X"EE",X"6F",X"FF",X"6F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",
		X"00",X"0E",X"0F",X"0F",X"0F",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"84",X"E1",X"DE",
		X"00",X"00",X"00",X"CC",X"6F",X"FF",X"6F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"86",
		X"00",X"00",X"00",X"88",X"6F",X"FF",X"7F",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"96",
		X"00",X"00",X"00",X"00",X"6F",X"FF",X"6F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"C3",X"78",X"0F",X"A5",
		X"00",X"00",X"00",X"00",X"6E",X"FF",X"6F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"78",X"5A",X"E5",
		X"00",X"00",X"00",X"00",X"4C",X"FF",X"7F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"E5",
		X"00",X"00",X"00",X"00",X"08",X"FF",X"6F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"F2",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"67",X"0E",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"8C",X"F1",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"E6",X"F8",
		X"00",X"00",X"00",X"00",X"48",X"10",X"00",X"0C",X"00",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",
		X"00",X"00",X"00",X"00",X"68",X"30",X"08",X"3C",X"00",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"CE",X"F0",X"F2",
		X"00",X"00",X"00",X"08",X"78",X"78",X"69",X"3C",X"00",X"00",X"CC",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"0E",X"EF",X"FF",X"F6",
		X"00",X"00",X"00",X"08",X"7C",X"79",X"69",X"3C",X"00",X"00",X"CC",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"EC",X"F6",
		X"00",X"00",X"E1",X"68",X"7E",X"F3",X"7E",X"3C",X"00",X"00",X"EE",X"13",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F6",
		X"00",X"E0",X"E1",X"69",X"7F",X"7F",X"6F",X"3F",X"00",X"00",X"EE",X"13",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"80",X"FF",X"F6",
		X"E0",X"EF",X"EF",X"6F",X"7F",X"7F",X"01",X"00",X"00",X"00",X"FF",X"13",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"EF",X"F3",X"F7",X"F6",
		X"EE",X"EF",X"EF",X"6F",X"7F",X"FF",X"E0",X"3C",X"00",X"00",X"FF",X"13",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"EE",X"77",X"00",X"F0",X"00",X"00",X"00",X"00",X"CE",X"E7",X"FF",X"FF",
		X"00",X"EE",X"EF",X"6F",X"7F",X"77",X"F0",X"3C",X"00",X"88",X"FF",X"13",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"CC",X"FF",X"FF",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"EE",X"FF",X"FF",
		X"00",X"00",X"EF",X"6E",X"7F",X"3B",X"3C",X"0F",X"00",X"88",X"FF",X"13",X"00",X"00",X"00",X"00",
		X"00",X"CC",X"FF",X"FE",X"FB",X"FF",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"FB",
		X"00",X"00",X"00",X"08",X"7F",X"59",X"B4",X"3C",X"00",X"88",X"FF",X"03",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"F2",X"F3",X"FE",X"FE",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EA",
		X"00",X"00",X"00",X"08",X"7F",X"68",X"3C",X"0F",X"00",X"88",X"3F",X"01",X"00",X"00",X"00",X"00",
		X"88",X"FF",X"FF",X"FC",X"F3",X"FE",X"FE",X"F1",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"FE",
		X"00",X"00",X"00",X"00",X"66",X"78",X"F0",X"3C",X"00",X"88",X"FF",X"10",X"00",X"00",X"00",X"00",
		X"CC",X"FF",X"FF",X"FF",X"F0",X"FF",X"FE",X"F1",X"00",X"00",X"00",X"00",X"33",X"E0",X"FB",X"F7",
		X"00",X"00",X"00",X"00",X"08",X"78",X"3C",X"0F",X"00",X"00",X"FF",X"10",X"00",X"00",X"00",X"00",
		X"CC",X"FF",X"FF",X"F3",X"FF",X"FF",X"FE",X"F1",X"00",X"00",X"00",X"00",X"FB",X"F3",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"08",X"78",X"B4",X"3C",X"00",X"00",X"FF",X"10",X"00",X"00",X"00",X"00",
		X"CC",X"FF",X"FF",X"FC",X"FF",X"FF",X"FE",X"F1",X"00",X"00",X"0E",X"0F",X"FE",X"F6",X"F4",X"FC",
		X"00",X"00",X"00",X"00",X"08",X"78",X"3F",X"0F",X"00",X"00",X"EE",X"10",X"00",X"00",X"00",X"00",
		X"CC",X"FF",X"FF",X"FC",X"FF",X"7F",X"FE",X"F1",X"00",X"00",X"00",X"00",X"C8",X"FE",X"F4",X"FC",
		X"00",X"00",X"00",X"00",X"08",X"78",X"FF",X"3F",X"00",X"00",X"EE",X"10",X"00",X"00",X"02",X"00",
		X"CC",X"FF",X"7F",X"DE",X"FF",X"3F",X"DE",X"E1",X"00",X"00",X"00",X"00",X"FB",X"FE",X"F4",X"FD",
		X"00",X"00",X"00",X"00",X"08",X"7E",X"3F",X"0F",X"00",X"00",X"EE",X"10",X"00",X"00",X"2A",X"00",
		X"8C",X"FF",X"3F",X"9E",X"EF",X"1F",X"9E",X"E1",X"00",X"00",X"00",X"CC",X"FD",X"FF",X"F4",X"FF",
		X"00",X"00",X"00",X"00",X"08",X"7F",X"BF",X"3F",X"00",X"00",X"E6",X"10",X"00",X"00",X"BB",X"00",
		X"0C",X"EF",X"1F",X"0F",X"0F",X"87",X"0F",X"E1",X"00",X"00",X"08",X"EF",X"FC",X"F1",X"FC",X"FF",
		X"00",X"00",X"00",X"00",X"08",X"7F",X"3F",X"0F",X"00",X"00",X"E2",X"00",X"00",X"00",X"FF",X"11",
		X"0C",X"00",X"00",X"00",X"0E",X"0F",X"0F",X"E1",X"00",X"00",X"00",X"00",X"88",X"F9",X"FE",X"FF",
		X"00",X"00",X"00",X"00",X"08",X"7F",X"FF",X"3F",X"00",X"00",X"80",X"00",X"00",X"00",X"FF",X"11",
		X"04",X"0F",X"0F",X"0F",X"01",X"00",X"0E",X"E1",X"00",X"00",X"00",X"88",X"F1",X"FF",X"FE",X"FD",
		X"00",X"00",X"00",X"00",X"08",X"7F",X"3F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"13",
		X"08",X"0F",X"0F",X"0F",X"0F",X"0F",X"01",X"F0",X"00",X"0C",X"EF",X"FE",X"F3",X"FF",X"F2",X"F5",
		X"00",X"00",X"00",X"00",X"08",X"7F",X"BF",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"13",
		X"0C",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"E1",X"00",X"00",X"88",X"FD",X"F2",X"FE",X"FA",X"F5",
		X"00",X"00",X"00",X"00",X"08",X"7F",X"3F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"01",
		X"0C",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"C3",X"00",X"00",X"00",X"00",X"C0",X"F6",X"F2",X"F5",
		X"00",X"00",X"01",X"00",X"08",X"7F",X"FF",X"3F",X"00",X"00",X"00",X"00",X"00",X"44",X"FE",X"01",
		X"0E",X"0F",X"87",X"0F",X"FF",X"B7",X"2F",X"C3",X"00",X"00",X"EE",X"F7",X"F0",X"F2",X"F2",X"F5",
		X"00",X"08",X"03",X"00",X"00",X"7F",X"3F",X"0F",X"00",X"00",X"00",X"00",X"00",X"44",X"7E",X"00",
		X"0E",X"CF",X"97",X"FF",X"FF",X"7F",X"3C",X"C3",X"08",X"8F",X"FF",X"F7",X"F2",X"F0",X"F2",X"F9",
		X"00",X"0C",X"07",X"00",X"00",X"6E",X"BF",X"3F",X"00",X"00",X"00",X"00",X"00",X"EE",X"6C",X"00",
		X"0E",X"FF",X"B7",X"FF",X"FF",X"FF",X"AD",X"D3",X"00",X"00",X"C0",X"F1",X"FC",X"F0",X"F8",X"FD",
		X"00",X"8E",X"2F",X"00",X"00",X"4C",X"3F",X"0F",X"00",X"00",X"00",X"00",X"00",X"EE",X"15",X"00",
		X"CE",X"FF",X"F7",X"FE",X"FF",X"FF",X"ED",X"F3",X"00",X"00",X"00",X"F0",X"FC",X"F0",X"FC",X"F9",
		X"00",X"CF",X"6F",X"01",X"08",X"38",X"FF",X"3F",X"00",X"00",X"00",X"00",X"00",X"FF",X"33",X"00",
		X"CE",X"FF",X"F7",X"FC",X"FF",X"FF",X"FD",X"F3",X"00",X"00",X"00",X"0C",X"9F",X"F1",X"FC",X"F9",
		X"00",X"EF",X"EF",X"E1",X"69",X"70",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"FF",X"77",X"00",
		X"EE",X"FF",X"F7",X"F8",X"FC",X"FF",X"FD",X"F3",X"00",X"00",X"00",X"00",X"7F",X"E9",X"F9",X"F9",
		X"00",X"EF",X"EF",X"E1",X"69",X"7F",X"F0",X"12",X"00",X"00",X"00",X"00",X"88",X"FF",X"77",X"00",
		X"EE",X"FF",X"FF",X"F3",X"F0",X"FF",X"FD",X"F3",X"00",X"00",X"08",X"FB",X"FF",X"F5",X"FA",X"F5",
		X"00",X"EF",X"EF",X"01",X"6F",X"7F",X"FF",X"D3",X"00",X"00",X"00",X"00",X"88",X"DF",X"FF",X"00",
		X"EE",X"FF",X"FF",X"FF",X"F3",X"FE",X"FD",X"F3",X"00",X"0E",X"EF",X"FD",X"FF",X"F7",X"F2",X"F1",
		X"00",X"EF",X"EF",X"01",X"6F",X"7F",X"FB",X"D3",X"00",X"00",X"00",X"00",X"CC",X"EF",X"FF",X"11",
		X"EE",X"FF",X"F7",X"FE",X"F7",X"FE",X"FD",X"F3",X"00",X"00",X"00",X"EC",X"F2",X"F7",X"FA",X"F9",
		X"00",X"EF",X"EF",X"E1",X"6F",X"7F",X"FF",X"D3",X"00",X"00",X"00",X"00",X"4C",X"FF",X"FF",X"11",
		X"CC",X"FF",X"F7",X"F8",X"F7",X"FF",X"FD",X"F3",X"88",X"FF",X"FB",X"F4",X"F2",X"F6",X"F0",X"F1",
		X"00",X"EF",X"EF",X"E1",X"6F",X"7F",X"FB",X"D3",X"00",X"00",X"00",X"00",X"4C",X"FF",X"FF",X"11",
		X"88",X"FF",X"F7",X"FF",X"FF",X"FF",X"FD",X"F1",X"EF",X"FD",X"FB",X"F2",X"F3",X"F4",X"F2",X"F9",
		X"00",X"CF",X"6F",X"01",X"08",X"7F",X"FF",X"D3",X"00",X"00",X"00",X"00",X"8C",X"FF",X"FC",X"11",
		X"00",X"EE",X"F7",X"FF",X"FF",X"FF",X"11",X"F0",X"00",X"00",X"F1",X"F7",X"F0",X"F0",X"F1",X"F1",
		X"00",X"8E",X"2F",X"00",X"00",X"08",X"FB",X"D3",X"00",X"00",X"00",X"00",X"8C",X"FF",X"FB",X"00",
		X"00",X"88",X"77",X"EE",X"FF",X"FF",X"11",X"F0",X"00",X"00",X"C8",X"F7",X"F0",X"F4",X"F5",X"F0",
		X"00",X"0C",X"07",X"00",X"F0",X"70",X"CC",X"D3",X"00",X"00",X"00",X"00",X"8C",X"FF",X"F7",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"F0",X"00",X"00",X"00",X"C4",X"F0",X"F4",X"F5",X"F0",
		X"00",X"08",X"03",X"08",X"F0",X"F0",X"01",X"C0",X"00",X"00",X"00",X"00",X"08",X"FF",X"FF",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"88",X"F9",X"F8",X"FC",X"FD",X"FC",
		X"00",X"00",X"01",X"48",X"F0",X"F0",X"2D",X"03",X"00",X"00",X"00",X"00",X"00",X"6F",X"FF",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"CF",X"FF",X"F5",X"F9",X"F1",X"FC",X"FF",X"FC",
		X"00",X"00",X"00",X"68",X"F0",X"F0",X"69",X"00",X"00",X"00",X"00",X"00",X"88",X"9F",X"FF",X"31",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"EE",X"F3",X"F8",X"F3",X"F0",X"FC",X"FD",
		X"00",X"00",X"00",X"69",X"FF",X"FF",X"69",X"00",X"04",X"00",X"00",X"00",X"88",X"FF",X"FF",X"31",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"E0",X"F8",X"FF",X"FB",X"FF",X"FD",
		X"00",X"00",X"80",X"6D",X"FF",X"FF",X"6B",X"90",X"4C",X"00",X"00",X"00",X"CC",X"FF",X"FF",X"31",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"E1",X"FA",X"FB",X"FF",X"FD",
		X"00",X"00",X"C0",X"6F",X"FF",X"FF",X"6F",X"F0",X"6E",X"00",X"00",X"00",X"EE",X"FF",X"FF",X"31",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"08",X"FE",X"FB",X"F3",X"FE",
		X"00",X"00",X"CC",X"6F",X"FF",X"FF",X"6F",X"FF",X"FF",X"01",X"00",X"00",X"EE",X"FF",X"FF",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"8E",X"F3",X"FF",X"FF",X"F1",X"FE",
		X"00",X"00",X"88",X"6F",X"FF",X"FF",X"6F",X"99",X"FF",X"01",X"00",X"00",X"EE",X"FF",X"F7",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"0F",X"8F",X"F5",X"F8",X"FE",X"FC",X"FB",
		X"00",X"00",X"00",X"6F",X"FF",X"FF",X"6F",X"00",X"FF",X"01",X"00",X"00",X"EE",X"FF",X"F3",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"08",X"0F",X"E1",X"F0",X"FC",X"F7",X"FA",X"FF",
		X"00",X"00",X"00",X"6E",X"FF",X"FF",X"6F",X"00",X"FF",X"01",X"00",X"00",X"EE",X"FF",X"B4",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"08",X"F0",X"FF",X"FB",X"F8",X"F3",
		X"00",X"00",X"00",X"4C",X"FF",X"FF",X"2F",X"0F",X"FF",X"01",X"00",X"00",X"CC",X"FF",X"1F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"08",X"80",X"FA",X"F7",X"F1",
		X"00",X"00",X"00",X"08",X"FF",X"FF",X"09",X"0F",X"CE",X"01",X"00",X"00",X"CC",X"FF",X"7F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"C8",X"FF",X"F9",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"64",X"00",X"0C",X"00",X"00",X"00",X"EE",X"FF",X"FF",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"ED",X"CF",X"0C",X"00",X"00",X"00",X"EE",X"FF",X"FF",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"88",X"FF",X"F9",
		X"00",X"00",X"00",X"00",X"FF",X"7B",X"ED",X"CF",X"08",X"00",X"00",X"00",X"CE",X"FF",X"FF",X"03",
		X"00",X"0E",X"0F",X"0F",X"07",X"00",X"00",X"F0",X"00",X"00",X"00",X"08",X"FF",X"F7",X"F2",X"FC",
		X"00",X"00",X"00",X"00",X"FF",X"F3",X"FC",X"CF",X"00",X"00",X"00",X"00",X"CE",X"FF",X"FF",X"13",
		X"08",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"E1",X"00",X"00",X"0C",X"CF",X"F4",X"F2",X"FA",X"FC",
		X"00",X"00",X"00",X"00",X"FF",X"F3",X"FC",X"CF",X"00",X"00",X"00",X"00",X"0E",X"FF",X"FF",X"17",
		X"0C",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"87",X"00",X"0E",X"0F",X"EF",X"F0",X"F2",X"F0",X"FC",
		X"00",X"00",X"00",X"00",X"FF",X"7B",X"ED",X"CF",X"00",X"00",X"00",X"00",X"04",X"F8",X"FF",X"37",
		X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"CF",X"FB",X"F2",X"F1",X"FA",
		X"00",X"00",X"00",X"00",X"FF",X"7B",X"ED",X"CF",X"00",X"00",X"00",X"00",X"80",X"F7",X"FF",X"37",
		X"0E",X"0F",X"0F",X"8F",X"FF",X"1F",X"2D",X"0F",X"00",X"00",X"00",X"00",X"ED",X"FF",X"7F",X"FB",
		X"00",X"00",X"00",X"00",X"FF",X"F3",X"FC",X"CF",X"00",X"00",X"00",X"00",X"C8",X"FF",X"FE",X"37",
		X"0F",X"EF",X"0F",X"EF",X"FF",X"7F",X"4B",X"0F",X"00",X"00",X"00",X"00",X"00",X"EC",X"FF",X"FB",
		X"00",X"00",X"00",X"00",X"FF",X"F3",X"FC",X"CF",X"00",X"00",X"00",X"00",X"CC",X"FF",X"FF",X"37",
		X"0F",X"FF",X"97",X"EF",X"FF",X"FF",X"87",X"4F",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"FB",
		X"00",X"00",X"00",X"00",X"FF",X"7B",X"ED",X"CF",X"00",X"00",X"00",X"00",X"EE",X"FF",X"FF",X"37",
		X"8F",X"FF",X"B7",X"FF",X"FF",X"FF",X"9F",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C8",
		X"00",X"00",X"00",X"00",X"FF",X"7B",X"ED",X"CF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"17",
		X"CF",X"FF",X"F7",X"FF",X"FF",X"FF",X"BF",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"FB",
		X"00",X"00",X"00",X"80",X"FF",X"F3",X"FC",X"CF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"13",
		X"EF",X"FF",X"F7",X"FE",X"FF",X"FF",X"FF",X"FE",X"00",X"00",X"00",X"00",X"00",X"8C",X"F6",X"F8",
		X"00",X"00",X"00",X"E0",X"FF",X"F3",X"FC",X"CF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"03",
		X"FF",X"FF",X"F7",X"FE",X"FF",X"FF",X"FF",X"FE",X"00",X"00",X"00",X"00",X"00",X"88",X"FF",X"F1",
		X"00",X"00",X"00",X"F0",X"EE",X"7B",X"ED",X"CF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"01",
		X"FF",X"FF",X"F7",X"F8",X"FF",X"FF",X"FF",X"FE",X"00",X"00",X"00",X"00",X"0C",X"CF",X"F3",X"F0",
		X"00",X"00",X"80",X"F0",X"FE",X"7B",X"ED",X"CF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"01",
		X"FF",X"FF",X"FF",X"F1",X"FC",X"FF",X"FF",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F4",
		X"00",X"00",X"C0",X"F8",X"DD",X"F3",X"FC",X"01",X"00",X"00",X"00",X"00",X"EE",X"FF",X"FF",X"01",
		X"FF",X"FF",X"FF",X"F7",X"F0",X"FE",X"FF",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"F7",
		X"00",X"00",X"C0",X"FE",X"BB",X"F3",X"FC",X"00",X"00",X"00",X"00",X"00",X"EE",X"FF",X"7F",X"00",
		X"FF",X"FF",X"F7",X"FE",X"F3",X"FC",X"FF",X"FE",X"00",X"00",X"00",X"00",X"00",X"08",X"CF",X"F3",
		X"00",X"00",X"E8",X"FF",X"77",X"7B",X"65",X"10",X"00",X"00",X"00",X"00",X"CC",X"FF",X"7F",X"00",
		X"EE",X"FF",X"F7",X"F8",X"F7",X"FE",X"FF",X"FE",X"00",X"00",X"00",X"00",X"0E",X"0F",X"8F",X"F0",
		X"00",X"00",X"EC",X"FF",X"FF",X"51",X"A0",X"10",X"00",X"00",X"00",X"00",X"CC",X"B9",X"37",X"00",
		X"88",X"FF",X"F7",X"FF",X"F7",X"FF",X"FF",X"F7",X"00",X"00",X"00",X"00",X"00",X"0E",X"FD",X"F0",
		X"00",X"00",X"EE",X"FF",X"FF",X"1B",X"DD",X"18",X"00",X"00",X"00",X"00",X"88",X"73",X"02",X"00",
		X"00",X"EE",X"F7",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"C2",X"F0",
		X"00",X"00",X"EE",X"FF",X"FF",X"7F",X"FF",X"1F",X"00",X"00",X"00",X"00",X"88",X"F7",X"01",X"00",
		X"00",X"88",X"77",X"EE",X"FF",X"FF",X"FF",X"F0",X"00",X"00",X"00",X"00",X"0E",X"0F",X"87",X"F0",
		X"00",X"00",X"EE",X"FF",X"FF",X"5F",X"FF",X"1F",X"00",X"00",X"00",X"00",X"00",X"FF",X"01",X"00",
		X"00",X"00",X"00",X"00",X"EE",X"FF",X"77",X"F0",X"00",X"00",X"00",X"00",X"00",X"0E",X"0F",X"F0",
		X"00",X"00",X"EE",X"FF",X"FF",X"5F",X"FF",X"19",X"00",X"00",X"00",X"CC",X"00",X"7F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"00",X"00",X"EE",X"FF",X"FF",X"7F",X"FF",X"11",X"00",X"00",X"00",X"EE",X"01",X"6E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E1",
		X"00",X"00",X"EE",X"FF",X"FF",X"5F",X"FF",X"11",X"00",X"00",X"00",X"FF",X"13",X"26",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"C3",
		X"00",X"00",X"CC",X"FF",X"FF",X"5F",X"FF",X"00",X"00",X"00",X"00",X"FF",X"37",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"C3",
		X"00",X"00",X"CC",X"FF",X"FF",X"7F",X"FF",X"01",X"00",X"00",X"88",X"FE",X"37",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"EE",X"FF",X"11",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"87",
		X"00",X"00",X"88",X"FF",X"FF",X"5F",X"7F",X"0F",X"00",X"00",X"CC",X"FD",X"37",X"00",X"00",X"00",
		X"00",X"00",X"EE",X"CC",X"FF",X"FF",X"33",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"84",
		X"00",X"00",X"00",X"FF",X"FF",X"5F",X"33",X"0F",X"00",X"00",X"CC",X"F3",X"7F",X"00",X"00",X"00",
		X"00",X"88",X"FF",X"FE",X"FF",X"FF",X"33",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"8C",
		X"00",X"00",X"00",X"EE",X"FF",X"00",X"00",X"00",X"00",X"00",X"CC",X"FF",X"7F",X"00",X"00",X"00",
		X"00",X"CC",X"FF",X"FC",X"F7",X"FF",X"FB",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CE",
		X"00",X"00",X"00",X"88",X"77",X"F0",X"78",X"09",X"00",X"00",X"CC",X"FF",X"7F",X"00",X"00",X"00",
		X"00",X"EE",X"FF",X"FC",X"F7",X"FE",X"FB",X"F1",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"E3",
		X"00",X"00",X"00",X"00",X"08",X"F0",X"69",X"2D",X"00",X"00",X"CC",X"FF",X"7F",X"00",X"00",X"00",
		X"00",X"EE",X"FF",X"FF",X"F1",X"FE",X"FB",X"F1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"00",X"00",X"00",X"00",X"48",X"F0",X"69",X"25",X"00",X"00",X"CC",X"FF",X"34",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"F7",X"F0",X"FF",X"FB",X"F1",X"00",X"00",X"00",X"00",X"00",X"0C",X"FF",X"F1",
		X"00",X"00",X"00",X"00",X"68",X"F0",X"78",X"21",X"00",X"00",X"88",X"FF",X"43",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"F0",X"FE",X"FF",X"DB",X"F1",X"00",X"00",X"00",X"00",X"0E",X"FF",X"F7",X"F8",
		X"00",X"00",X"00",X"00",X"69",X"FF",X"6F",X"21",X"00",X"00",X"88",X"FF",X"B7",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"F8",X"FF",X"FF",X"CB",X"F1",X"00",X"00",X"00",X"00",X"00",X"CF",X"F1",X"F8",
		X"00",X"00",X"00",X"80",X"6F",X"FF",X"6F",X"2B",X"00",X"00",X"00",X"FF",X"B7",X"00",X"00",X"00",
		X"00",X"EF",X"7F",X"FE",X"FF",X"0F",X"4B",X"E1",X"00",X"00",X"00",X"00",X"00",X"00",X"E4",X"F5",
		X"00",X"00",X"00",X"C0",X"6F",X"FF",X"7F",X"2B",X"00",X"00",X"00",X"FF",X"7F",X"10",X"00",X"00",
		X"00",X"0F",X"0F",X"1E",X"0F",X"0F",X"2D",X"E1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E4",
		X"00",X"00",X"00",X"EE",X"6F",X"FF",X"6F",X"2F",X"00",X"00",X"00",X"EE",X"FF",X"21",X"00",X"00",
		X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"1E",X"E1",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"F5",
		X"00",X"00",X"00",X"CC",X"6F",X"FF",X"6F",X"2B",X"00",X"00",X"00",X"2E",X"FF",X"21",X"00",X"00",
		X"00",X"03",X"0C",X"01",X"00",X"00",X"0F",X"E1",X"00",X"00",X"00",X"00",X"00",X"CC",X"FF",X"F1",
		X"00",X"00",X"00",X"88",X"6F",X"FF",X"7F",X"2B",X"00",X"00",X"00",X"CE",X"FF",X"21",X"00",X"00",
		X"00",X"0C",X"03",X"0E",X"0F",X"0F",X"00",X"F0",X"00",X"00",X"00",X"0E",X"8F",X"FF",X"F7",X"F3",
		X"00",X"00",X"00",X"00",X"6F",X"FF",X"6F",X"23",X"00",X"00",X"00",X"FF",X"FF",X"21",X"00",X"00",
		X"00",X"0F",X"4B",X"0F",X"0F",X"0F",X"4B",X"C3",X"00",X"00",X"0E",X"EF",X"F7",X"FF",X"F4",X"F3",
		X"00",X"00",X"00",X"00",X"6E",X"FF",X"6F",X"23",X"00",X"00",X"00",X"FF",X"7F",X"10",X"00",X"00",
		X"08",X"0F",X"4B",X"0F",X"CF",X"7F",X"87",X"87",X"00",X"00",X"00",X"0E",X"FE",X"F0",X"FF",X"F2",
		X"00",X"C0",X"00",X"C2",X"5C",X"FF",X"7F",X"27",X"00",X"00",X"00",X"FF",X"F3",X"00",X"00",X"00",
		X"0C",X"0F",X"C3",X"8F",X"FF",X"FF",X"1F",X"96",X"00",X"00",X"00",X"00",X"C3",X"F1",X"F3",X"FA",
		X"00",X"E0",X"10",X"C3",X"38",X"FF",X"6F",X"2F",X"00",X"00",X"00",X"FF",X"7F",X"00",X"00",X"00",
		X"0E",X"8F",X"D3",X"FF",X"FF",X"FF",X"3F",X"96",X"00",X"00",X"00",X"00",X"00",X"E0",X"F0",X"F8",
		X"00",X"FE",X"D2",X"CF",X"77",X"FF",X"6F",X"09",X"00",X"00",X"00",X"FF",X"7F",X"00",X"00",X"00",
		X"0E",X"FF",X"F3",X"FE",X"FF",X"FF",X"7F",X"D6",X"00",X"00",X"00",X"00",X"00",X"C8",X"F0",X"F1",
		X"00",X"FF",X"DF",X"CF",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"37",X"00",X"00",X"00",
		X"CE",X"FF",X"F3",X"F0",X"FF",X"FE",X"FF",X"F6",X"00",X"00",X"00",X"00",X"CF",X"F7",X"F7",X"F1",
		X"00",X"EE",X"11",X"CF",X"7F",X"EF",X"9F",X"3F",X"00",X"00",X"00",X"EE",X"37",X"00",X"00",X"00",
		X"EE",X"FF",X"F3",X"F0",X"F0",X"FC",X"FF",X"F6",X"00",X"00",X"08",X"CF",X"F7",X"F4",X"F2",X"F4",
		X"00",X"CC",X"00",X"CE",X"7F",X"49",X"8E",X"3F",X"00",X"00",X"00",X"EE",X"37",X"00",X"00",X"00",
		X"EE",X"FF",X"FB",X"FF",X"FF",X"F8",X"FF",X"F6",X"00",X"0C",X"8F",X"F7",X"F7",X"F9",X"F5",X"F6",
		X"00",X"00",X"00",X"00",X"09",X"48",X"8C",X"3F",X"00",X"00",X"00",X"CC",X"13",X"00",X"00",X"00",
		X"EE",X"FF",X"FB",X"FF",X"FF",X"F8",X"FF",X"F6",X"00",X"00",X"08",X"6B",X"F7",X"FB",X"FD",X"F2",
		X"00",X"00",X"00",X"00",X"01",X"48",X"00",X"0C",X"00",X"00",X"00",X"CC",X"13",X"00",X"00",X"00",
		X"EE",X"FF",X"F3",X"F8",X"FF",X"FC",X"FF",X"F6",X"00",X"00",X"00",X"86",X"F9",X"FA",X"FD",X"F2",
		X"00",X"00",X"00",X"0C",X"03",X"48",X"00",X"08",X"00",X"00",X"00",X"88",X"01",X"00",X"00",X"00",
		X"EE",X"FF",X"F3",X"FE",X"FF",X"FE",X"FF",X"F6",X"00",X"08",X"0F",X"CF",X"F9",X"F4",X"F6",X"F7",
		X"00",X"00",X"00",X"00",X"00",X"48",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",
		X"EE",X"FF",X"F3",X"FF",X"FF",X"FF",X"FF",X"F6",X"0C",X"0F",X"8F",X"FF",X"F2",X"F0",X"F6",X"F5",
		X"00",X"00",X"00",X"00",X"00",X"48",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"FF",X"F3",X"FF",X"FF",X"FF",X"FF",X"F6",X"00",X"00",X"0C",X"C7",X"F4",X"F1",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"48",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"FF",X"F3",X"FF",X"FF",X"FF",X"F7",X"F7",X"00",X"00",X"00",X"00",X"00",X"F9",X"E9",X"F2",
		X"00",X"00",X"00",X"00",X"00",X"48",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"FF",X"FB",X"FF",X"FF",X"FF",X"FB",X"F3",X"00",X"00",X"00",X"00",X"00",X"00",X"E5",X"F2",
		X"00",X"00",X"00",X"00",X"00",X"48",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"FB",X"FF",X"FF",X"FF",X"31",X"F0",X"00",X"00",X"00",X"00",X"00",X"FE",X"E7",X"F3",
		X"00",X"00",X"00",X"00",X"00",X"48",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",
		X"00",X"CC",X"33",X"EE",X"FF",X"77",X"00",X"F0",X"00",X"00",X"00",X"00",X"C3",X"7A",X"F6",X"F5",
		X"00",X"00",X"00",X"00",X"00",X"48",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"77",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"0C",X"69",X"FF",X"F4",
		X"00",X"00",X"00",X"00",X"00",X"48",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"F7",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"80",X"F9",X"F4",
		X"00",X"00",X"00",X"00",X"00",X"48",X"00",X"00",X"00",X"88",X"11",X"00",X"00",X"CC",X"FF",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"F4",
		X"00",X"00",X"00",X"00",X"00",X"48",X"00",X"00",X"00",X"88",X"33",X"00",X"00",X"CC",X"FF",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"84",X"F4",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"48",X"00",X"00",X"00",X"CC",X"33",X"00",X"00",X"CC",X"BF",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"0F",X"8F",X"F4",X"FD",
		X"00",X"00",X"00",X"00",X"00",X"48",X"00",X"00",X"00",X"CC",X"73",X"00",X"00",X"CC",X"7F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"0F",X"F8",X"FB",
		X"00",X"00",X"00",X"0E",X"03",X"48",X"00",X"08",X"00",X"EE",X"73",X"00",X"00",X"EE",X"FF",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"CB",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"48",X"00",X"0C",X"00",X"E6",X"73",X"00",X"00",X"EE",X"FF",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E6",
		X"00",X"00",X"00",X"00",X"09",X"48",X"84",X"3C",X"00",X"FF",X"30",X"00",X"00",X"FF",X"FF",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"E8",X"F6",
		X"00",X"C0",X"00",X"C2",X"78",X"49",X"86",X"3C",X"00",X"FF",X"13",X"00",X"80",X"FF",X"FF",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"8E",X"F9",X"F4",
		X"00",X"E0",X"10",X"C3",X"78",X"E1",X"96",X"3C",X"00",X"EF",X"13",X"00",X"80",X"FF",X"7F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"C4",X"F2",
		X"00",X"FE",X"D2",X"CF",X"7F",X"E1",X"9E",X"3F",X"00",X"6F",X"13",X"00",X"80",X"FF",X"17",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"C0",X"F6",X"F1",
		X"00",X"FF",X"DF",X"CF",X"7F",X"EF",X"9F",X"3F",X"00",X"8E",X"13",X"00",X"00",X"FE",X"F3",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"87",X"FE",X"F0",X"F2",X"F5",
		X"00",X"EE",X"11",X"CF",X"7F",X"EF",X"9F",X"3F",X"00",X"EE",X"01",X"00",X"00",X"F9",X"F7",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"C4",X"F4",X"FF",X"F4",
		X"00",X"CC",X"00",X"CE",X"7F",X"01",X"8E",X"3F",X"00",X"CC",X"01",X"00",X"88",X"FF",X"F7",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"C4",X"F9",X"F5",
		X"00",X"00",X"00",X"00",X"09",X"00",X"8C",X"3F",X"00",X"0C",X"00",X"00",X"88",X"FF",X"F7",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"88",X"FF",X"F7",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"FF",
		X"00",X"00",X"00",X"0E",X"03",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"CC",X"FF",X"E7",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"80",X"F2",X"FA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"FF",X"53",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"88",X"F4",X"F2",X"FA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EF",X"37",X"00",
		X"00",X"00",X"00",X"00",X"EE",X"FF",X"11",X"F0",X"00",X"00",X"0C",X"0F",X"EF",X"F0",X"F8",X"F5",
		X"00",X"00",X"00",X"00",X"00",X"00",X"5A",X"18",X"00",X"00",X"00",X"00",X"6E",X"FF",X"37",X"00",
		X"00",X"00",X"CC",X"DD",X"FF",X"FF",X"33",X"F0",X"08",X"0F",X"0F",X"CF",X"F3",X"F1",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"80",X"5A",X"78",X"00",X"00",X"00",X"00",X"6E",X"FF",X"37",X"00",
		X"00",X"00",X"FF",X"FD",X"F7",X"FF",X"33",X"F0",X"00",X"00",X"00",X"86",X"FD",X"F0",X"E1",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"1E",X"3C",X"00",X"00",X"00",X"44",X"6E",X"FF",X"37",X"00",
		X"00",X"88",X"FF",X"F1",X"F7",X"FE",X"FB",X"F0",X"00",X"00",X"00",X"00",X"00",X"F0",X"E5",X"F1",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"5A",X"3C",X"00",X"00",X"00",X"66",X"EE",X"EF",X"37",X"00",
		X"00",X"CC",X"FF",X"F9",X"F7",X"FE",X"FB",X"F0",X"00",X"00",X"08",X"8F",X"F0",X"78",X"F5",X"F5",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"5A",X"3C",X"00",X"00",X"00",X"EE",X"EE",X"DF",X"37",X"00",
		X"00",X"EE",X"FF",X"FF",X"F1",X"FF",X"FB",X"F0",X"00",X"00",X"00",X"C4",X"F0",X"B4",X"F7",X"F7",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"1E",X"78",X"00",X"00",X"00",X"EE",X"DD",X"FF",X"9F",X"00",
		X"00",X"EE",X"FF",X"F7",X"F8",X"FF",X"7B",X"F0",X"00",X"0C",X"ED",X"F1",X"F0",X"D6",X"F6",X"F6",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"5A",X"78",X"00",X"00",X"00",X"EE",X"DD",X"FF",X"9B",X"00",
		X"00",X"0E",X"FF",X"F1",X"1E",X"0F",X"4B",X"F0",X"00",X"00",X"08",X"F2",X"F4",X"E9",X"F2",X"F2",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"5B",X"78",X"00",X"00",X"00",X"FF",X"BB",X"FF",X"CF",X"10",
		X"00",X"0E",X"0F",X"69",X"01",X"00",X"4A",X"F0",X"00",X"00",X"00",X"00",X"3C",X"FB",X"F2",X"F1",
		X"00",X"00",X"00",X"00",X"80",X"F8",X"1F",X"78",X"00",X"00",X"00",X"FF",X"BB",X"3F",X"CD",X"10",
		X"00",X"0E",X"00",X"21",X"EE",X"FF",X"59",X"F0",X"00",X"00",X"00",X"00",X"00",X"C0",X"F0",X"F1",
		X"00",X"00",X"00",X"00",X"80",X"FC",X"5B",X"7F",X"00",X"00",X"00",X"9F",X"73",X"FF",X"EE",X"10",
		X"00",X"02",X"FF",X"CC",X"FF",X"FF",X"7B",X"F0",X"00",X"00",X"00",X"00",X"C0",X"F5",X"F0",X"F1",
		X"00",X"00",X"00",X"00",X"80",X"FE",X"5B",X"3F",X"00",X"00",X"00",X"EF",X"73",X"FF",X"FF",X"10",
		X"00",X"CC",X"FF",X"FE",X"FB",X"FF",X"33",X"F0",X"00",X"00",X"00",X"EE",X"FD",X"78",X"F8",X"F8",
		X"00",X"00",X"00",X"00",X"C0",X"FF",X"1F",X"3F",X"00",X"00",X"88",X"FF",X"73",X"FF",X"FF",X"10",
		X"00",X"FF",X"FF",X"F2",X"F3",X"FE",X"FB",X"F0",X"00",X"0E",X"CF",X"F7",X"F0",X"B4",X"F8",X"FC",
		X"00",X"00",X"00",X"00",X"C0",X"FF",X"5B",X"3F",X"00",X"00",X"CC",X"FF",X"73",X"FF",X"FF",X"10",
		X"88",X"FF",X"FF",X"FC",X"F3",X"FE",X"FB",X"F1",X"00",X"00",X"0E",X"FB",X"F0",X"C7",X"F8",X"FC",
		X"00",X"00",X"00",X"00",X"C8",X"FF",X"5B",X"7F",X"00",X"00",X"CC",X"FF",X"73",X"EE",X"F7",X"00",
		X"CC",X"FF",X"FF",X"FF",X"F0",X"FF",X"FB",X"F1",X"00",X"00",X"00",X"84",X"3C",X"F6",X"F0",X"FD",
		X"00",X"00",X"00",X"00",X"C8",X"FF",X"1F",X"7F",X"00",X"00",X"CC",X"FF",X"73",X"CC",X"F7",X"00",
		X"CC",X"FF",X"FF",X"F3",X"FC",X"FF",X"FB",X"F1",X"00",X"00",X"00",X"00",X"C7",X"F0",X"F0",X"FB",
		X"00",X"00",X"00",X"00",X"CC",X"FF",X"5B",X"7F",X"00",X"00",X"CC",X"FF",X"71",X"CC",X"F7",X"00",
		X"CC",X"FF",X"FF",X"F0",X"FE",X"FF",X"DB",X"F1",X"00",X"00",X"00",X"88",X"F6",X"F4",X"F2",X"F2",
		X"00",X"00",X"00",X"00",X"CC",X"FF",X"5B",X"7F",X"00",X"00",X"EE",X"FF",X"31",X"80",X"F3",X"00",
		X"CC",X"FF",X"FF",X"FC",X"FF",X"FF",X"CB",X"F1",X"00",X"00",X"08",X"EF",X"FF",X"F0",X"F0",X"F2",
		X"00",X"00",X"00",X"00",X"CC",X"FF",X"1F",X"7F",X"00",X"00",X"EE",X"FF",X"10",X"80",X"70",X"00",
		X"CC",X"FF",X"7F",X"FC",X"FF",X"7F",X"ED",X"F1",X"00",X"00",X"00",X"00",X"F6",X"F1",X"F0",X"F2",
		X"00",X"00",X"00",X"00",X"CC",X"FF",X"5B",X"3F",X"00",X"00",X"EE",X"FF",X"13",X"00",X"60",X"00",
		X"8C",X"FF",X"7F",X"9E",X"FF",X"1F",X"9E",X"E1",X"00",X"00",X"88",X"FB",X"FD",X"F1",X"F0",X"F2",
		X"00",X"00",X"00",X"00",X"CC",X"FF",X"5B",X"3F",X"00",X"00",X"CE",X"FF",X"13",X"00",X"20",X"00",
		X"0C",X"FF",X"3F",X"1E",X"0F",X"87",X"0F",X"E1",X"00",X"8F",X"FF",X"F4",X"F9",X"F1",X"F7",X"F3",
		X"00",X"00",X"00",X"00",X"CC",X"FF",X"1F",X"3F",X"00",X"00",X"CE",X"FF",X"37",X"00",X"00",X"00",
		X"0C",X"EF",X"1F",X"0F",X"0F",X"0F",X"0F",X"E1",X"0F",X"FF",X"F7",X"F1",X"F0",X"F9",X"F9",X"F3",
		X"00",X"00",X"00",X"00",X"88",X"FF",X"5B",X"7F",X"00",X"00",X"BF",X"FF",X"37",X"00",X"00",X"00",
		X"0C",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"E1",X"00",X"CC",X"F1",X"FA",X"F0",X"FD",X"F8",X"F3",
		X"00",X"00",X"00",X"00",X"88",X"FF",X"5B",X"7F",X"00",X"00",X"7F",X"FF",X"37",X"00",X"00",X"00",
		X"08",X"07",X"00",X"00",X"00",X"08",X"0F",X"E1",X"00",X"00",X"E0",X"F0",X"F4",X"FD",X"F0",X"F1",
		X"00",X"00",X"00",X"00",X"88",X"FF",X"1F",X"7F",X"00",X"88",X"FF",X"FF",X"37",X"00",X"00",X"00",
		X"00",X"09",X"0F",X"0C",X"0F",X"07",X"00",X"F0",X"0E",X"0F",X"C3",X"F0",X"F6",X"FC",X"F4",X"F1",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"5B",X"7F",X"00",X"88",X"FF",X"FF",X"37",X"00",X"00",X"00",
		X"00",X"0E",X"0F",X"1E",X"0F",X"0F",X"3C",X"E1",X"00",X"00",X"0C",X"F0",X"FA",X"F2",X"F8",X"F1",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"5B",X"7F",X"00",X"88",X"FF",X"FF",X"37",X"00",X"00",X"00",
		X"00",X"0F",X"0F",X"1E",X"FF",X"3F",X"69",X"C3",X"00",X"00",X"00",X"00",X"F9",X"F3",X"F0",X"F5",
		X"00",X"00",X"00",X"00",X"00",X"EE",X"1F",X"3F",X"00",X"88",X"FF",X"FF",X"33",X"00",X"00",X"00",
		X"08",X"EF",X"3F",X"BC",X"FF",X"FF",X"C3",X"C3",X"00",X"00",X"00",X"FF",X"FD",X"F8",X"F2",X"F1",
		X"00",X"00",X"00",X"00",X"00",X"EE",X"5B",X"3F",X"00",X"88",X"FF",X"BF",X"13",X"00",X"00",X"00",
		X"0C",X"FF",X"7F",X"FC",X"FF",X"FF",X"97",X"D3",X"00",X"0F",X"8F",X"FD",X"F6",X"F8",X"FB",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"5B",X"3F",X"00",X"88",X"FF",X"7B",X"01",X"00",X"00",X"00",
		X"8C",X"FF",X"FF",X"F0",X"FE",X"FD",X"B7",X"F3",X"00",X"00",X"0E",X"C3",X"F0",X"F0",X"FA",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"1F",X"7F",X"00",X"88",X"FF",X"F7",X"30",X"00",X"00",X"00",
		X"CC",X"FF",X"FF",X"F0",X"F0",X"F8",X"F7",X"F3",X"00",X"00",X"00",X"0C",X"E1",X"F0",X"FA",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"88",X"5B",X"7F",X"00",X"08",X"FF",X"FF",X"70",X"00",X"00",X"00",
		X"CC",X"FF",X"FF",X"FF",X"FF",X"F8",X"F7",X"F3",X"00",X"00",X"00",X"00",X"00",X"F4",X"F4",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"5B",X"19",X"00",X"00",X"EF",X"FF",X"71",X"00",X"00",X"00",
		X"CC",X"FF",X"FF",X"FF",X"FF",X"F8",X"F7",X"F3",X"00",X"00",X"00",X"00",X"08",X"E9",X"F0",X"F6",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"8E",X"FF",X"71",X"00",X"00",X"00",
		X"CC",X"FF",X"FF",X"F0",X"FE",X"F9",X"F7",X"F3",X"00",X"00",X"00",X"00",X"00",X"80",X"F4",X"F7",
		X"00",X"00",X"00",X"00",X"48",X"10",X"00",X"0C",X"00",X"00",X"FF",X"FF",X"73",X"00",X"00",X"00",
		X"CC",X"FF",X"FF",X"FC",X"FF",X"FD",X"F7",X"F3",X"00",X"00",X"00",X"00",X"00",X"00",X"4C",X"F5",
		X"00",X"00",X"00",X"00",X"68",X"30",X"08",X"3C",X"00",X"88",X"FF",X"FF",X"73",X"00",X"00",X"00",
		X"CC",X"FF",X"FF",X"FC",X"FF",X"FF",X"F7",X"F3",X"00",X"00",X"00",X"00",X"00",X"88",X"7B",X"F7",
		X"00",X"00",X"00",X"00",X"78",X"78",X"69",X"3C",X"00",X"88",X"FF",X"FF",X"73",X"00",X"00",X"00",
		X"88",X"FF",X"FF",X"FC",X"FF",X"FF",X"F7",X"F3",X"00",X"00",X"00",X"00",X"0C",X"EF",X"BD",X"F7",
		X"00",X"00",X"80",X"FF",X"7C",X"79",X"69",X"3C",X"00",X"88",X"FF",X"FF",X"73",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"FC",X"FF",X"FF",X"FB",X"F3",X"00",X"00",X"00",X"00",X"00",X"80",X"BC",X"F3",
		X"04",X"00",X"86",X"0F",X"7E",X"F3",X"7E",X"3C",X"00",X"88",X"FF",X"DF",X"31",X"00",X"44",X"11",
		X"00",X"EE",X"FF",X"FE",X"FF",X"FF",X"FD",X"F1",X"00",X"00",X"00",X"00",X"0E",X"0F",X"DE",X"FB",
		X"0E",X"C2",X"96",X"FF",X"7F",X"7F",X"6F",X"3F",X"00",X"00",X"FF",X"CF",X"31",X"00",X"EE",X"11",
		X"00",X"88",X"FF",X"CC",X"FF",X"FF",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"ED",X"FF",
		X"0F",X"C3",X"96",X"0F",X"7F",X"7F",X"6F",X"3F",X"00",X"00",X"4F",X"ED",X"30",X"00",X"6E",X"31",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",
		X"0F",X"CF",X"97",X"0F",X"7F",X"FF",X"7F",X"3F",X"00",X"00",X"0E",X"F1",X"32",X"00",X"AE",X"31",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"11",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"F7",X"F4",
		X"0E",X"CE",X"97",X"FF",X"7F",X"7F",X"01",X"26",X"00",X"00",X"00",X"F3",X"32",X"00",X"AE",X"31",
		X"00",X"00",X"FF",X"CC",X"FF",X"FF",X"33",X"F0",X"00",X"00",X"00",X"00",X"0C",X"0F",X"F0",X"F4",
		X"04",X"00",X"86",X"0F",X"7F",X"7F",X"A4",X"09",X"00",X"00",X"00",X"EE",X"33",X"00",X"EE",X"31",
		X"00",X"CC",X"FF",X"FE",X"FB",X"FF",X"33",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"F4",
		X"00",X"00",X"80",X"FF",X"7F",X"77",X"B4",X"6F",X"00",X"00",X"00",X"CC",X"11",X"00",X"CC",X"10",
		X"00",X"FF",X"FF",X"F2",X"F3",X"FE",X"FB",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"00",X"00",X"00",X"00",X"7F",X"B3",X"3C",X"2F",X"00",X"00",X"00",X"CC",X"00",X"00",X"CC",X"10",
		X"88",X"FF",X"FF",X"FC",X"F3",X"FE",X"FB",X"F1",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"F3",
		X"00",X"00",X"00",X"00",X"6E",X"B3",X"3C",X"2F",X"00",X"00",X"00",X"88",X"00",X"00",X"88",X"00",
		X"CC",X"FF",X"FF",X"FF",X"F0",X"FF",X"FB",X"F1",X"00",X"00",X"00",X"00",X"00",X"0E",X"0F",X"C3",
		X"00",X"00",X"00",X"00",X"4C",X"D1",X"B4",X"6F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"FF",X"FF",X"F3",X"FF",X"FF",X"FB",X"F1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"B4",X"6F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"FF",X"FF",X"FC",X"FF",X"FF",X"DB",X"F1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E9",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"3C",X"6F",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"FF",X"FF",X"FC",X"FF",X"7F",X"CB",X"F1",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"3C",X"6F",X"00",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"FF",X"7F",X"DE",X"FF",X"3F",X"ED",X"E1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"B4",X"2F",X"00",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"8C",X"FF",X"3F",X"9E",X"FF",X"1F",X"9E",X"E1",X"00",X"00",X"00",X"00",X"00",X"CC",X"F3",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"B7",X"2F",X"00",X"00",X"CC",X"01",X"00",X"00",X"00",X"00",
		X"0C",X"EF",X"1F",X"0F",X"0F",X"87",X"0F",X"E1",X"00",X"00",X"00",X"08",X"8F",X"FF",X"F5",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"FC",X"3F",X"6F",X"00",X"00",X"CC",X"01",X"00",X"00",X"00",X"00",
		X"0C",X"00",X"00",X"00",X"0E",X"0F",X"0F",X"E1",X"00",X"00",X"0C",X"8F",X"FF",X"F3",X"F5",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"FE",X"3F",X"6F",X"00",X"00",X"EE",X"13",X"00",X"00",X"00",X"00",
		X"04",X"0F",X"0F",X"0F",X"01",X"00",X"0E",X"E1",X"00",X"00",X"00",X"08",X"F5",X"F0",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"B7",X"6F",X"00",X"00",X"EE",X"13",X"00",X"00",X"00",X"00",
		X"08",X"0F",X"0F",X"0F",X"0F",X"0F",X"01",X"F0",X"00",X"00",X"00",X"00",X"00",X"F0",X"FF",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"B7",X"6F",X"00",X"00",X"FF",X"13",X"00",X"00",X"00",X"00",
		X"0C",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"E1",X"00",X"00",X"00",X"F7",X"F9",X"F3",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"3F",X"2F",X"00",X"00",X"FF",X"13",X"00",X"00",X"00",X"00",
		X"0C",X"0F",X"0F",X"0F",X"0F",X"4B",X"0F",X"C3",X"00",X"0E",X"EF",X"F7",X"FB",X"FB",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"3F",X"2F",X"00",X"88",X"FF",X"13",X"00",X"00",X"00",X"00",
		X"0E",X"0F",X"87",X"0F",X"CF",X"B7",X"0F",X"C3",X"00",X"00",X"00",X"EE",X"FB",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"B7",X"6F",X"00",X"88",X"FF",X"13",X"00",X"00",X"00",X"00",
		X"0E",X"0F",X"87",X"BF",X"FF",X"7F",X"1E",X"C3",X"00",X"00",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"B7",X"6F",X"00",X"88",X"FF",X"03",X"00",X"00",X"00",X"00",
		X"0E",X"8F",X"B7",X"FF",X"FF",X"FF",X"AD",X"D3",X"0E",X"CF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"3F",X"6F",X"00",X"88",X"3F",X"01",X"00",X"00",X"00",X"00",
		X"0E",X"FF",X"F7",X"FE",X"FF",X"FF",X"EB",X"F3",X"00",X"00",X"CE",X"FD",X"FF",X"FE",X"FE",X"F7",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"3F",X"6F",X"00",X"88",X"FE",X"00",X"00",X"00",X"00",X"00",
		X"CE",X"FF",X"F7",X"FC",X"FF",X"FF",X"FB",X"F3",X"00",X"00",X"00",X"E8",X"FF",X"FE",X"FE",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"B7",X"2F",X"00",X"80",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"FF",X"F7",X"F8",X"FC",X"FF",X"FB",X"F3",X"00",X"00",X"00",X"00",X"FF",X"F4",X"F6",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"B7",X"2F",X"00",X"88",X"FF",X"10",X"00",X"00",X"00",X"00",
		X"EE",X"FF",X"FF",X"F3",X"F0",X"FF",X"FB",X"F3",X"00",X"00",X"0C",X"CB",X"F2",X"F5",X"F0",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"EE",X"3F",X"23",X"00",X"88",X"FF",X"10",X"00",X"00",X"00",X"00",
		X"EE",X"FF",X"FF",X"FF",X"F3",X"FE",X"FB",X"F3",X"00",X"00",X"00",X"0C",X"F7",X"FD",X"F4",X"FD",
		X"00",X"00",X"00",X"00",X"48",X"DC",X"37",X"0C",X"00",X"88",X"FF",X"10",X"00",X"00",X"00",X"00",
		X"EE",X"FF",X"F7",X"FE",X"F7",X"FE",X"FB",X"F3",X"00",X"00",X"FF",X"FE",X"F7",X"FE",X"FF",X"FD",
		X"00",X"00",X"00",X"00",X"68",X"30",X"08",X"3C",X"00",X"88",X"FF",X"10",X"00",X"00",X"00",X"00",
		X"CC",X"FF",X"F7",X"F8",X"F7",X"FF",X"FB",X"F3",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"00",X"00",X"00",X"08",X"78",X"78",X"69",X"3C",X"00",X"88",X"FF",X"10",X"00",X"00",X"00",X"00",
		X"88",X"FF",X"F7",X"FF",X"FF",X"FF",X"FB",X"F1",X"00",X"00",X"EA",X"F9",X"FE",X"FF",X"FB",X"FE",
		X"00",X"00",X"00",X"08",X"7C",X"79",X"69",X"3C",X"00",X"00",X"FF",X"10",X"00",X"00",X"00",X"00",
		X"00",X"EE",X"F7",X"FF",X"FF",X"FF",X"33",X"F0",X"00",X"00",X"00",X"00",X"F9",X"FF",X"FF",X"FE",
		X"00",X"00",X"E1",X"68",X"7E",X"F3",X"7E",X"3C",X"00",X"00",X"F6",X"10",X"00",X"00",X"00",X"00",
		X"00",X"88",X"77",X"EE",X"FF",X"FF",X"33",X"F0",X"00",X"00",X"08",X"C3",X"F3",X"FD",X"FF",X"F7",
		X"00",X"E0",X"E1",X"69",X"7F",X"7F",X"6F",X"3F",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"11",X"F0",X"00",X"0C",X"0F",X"0F",X"F7",X"FB",X"F6",X"F7",
		X"E0",X"EF",X"EF",X"6F",X"7F",X"7F",X"6F",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"8F",X"FB",X"F5",X"F7",
		X"EE",X"EF",X"EF",X"6F",X"7F",X"F7",X"7E",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"CC",X"FF",X"F7",
		X"00",X"EE",X"EF",X"6F",X"7F",X"7F",X"6F",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"EC",X"F7",
		X"00",X"00",X"EF",X"6E",X"7F",X"7F",X"6F",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E2",
		X"00",X"00",X"00",X"08",X"7F",X"F7",X"7E",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"08",X"2F",X"EF",X"FB",
		X"00",X"00",X"00",X"08",X"7F",X"7F",X"6F",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"8E",X"F8",
		X"00",X"00",X"00",X"00",X"6E",X"33",X"08",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"F8",
		X"00",X"00",X"00",X"00",X"4C",X"11",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
