library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity program1x is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of program1x is
	type rom is array(0 to  10239) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"32",X"45",X"40",X"7D",X"32",X"54",X"50",X"7C",X"32",X"57",X"50",X"C9",X"3A",X"43",X"40",X"A7",
		X"20",X"17",X"3A",X"47",X"40",X"A7",X"20",X"11",X"3E",X"01",X"32",X"47",X"40",X"21",X"F1",X"26",
		X"22",X"50",X"50",X"21",X"02",X"A7",X"22",X"52",X"50",X"3A",X"45",X"40",X"A7",X"20",X"17",X"3A",
		X"48",X"40",X"A7",X"20",X"11",X"3E",X"01",X"32",X"48",X"40",X"21",X"F1",X"26",X"22",X"54",X"50",
		X"21",X"02",X"87",X"22",X"56",X"50",X"3A",X"59",X"50",X"FE",X"A8",X"C8",X"3A",X"58",X"50",X"FE",
		X"F0",X"38",X"1C",X"3A",X"47",X"40",X"A7",X"28",X"16",X"3A",X"50",X"50",X"32",X"58",X"50",X"3A",
		X"53",X"50",X"32",X"5B",X"50",X"3E",X"27",X"32",X"59",X"50",X"3E",X"04",X"CD",X"96",X"2C",X"3A",
		X"5C",X"50",X"FE",X"F8",X"D8",X"3A",X"48",X"40",X"A7",X"C8",X"3A",X"54",X"50",X"32",X"5C",X"50",
		X"3A",X"57",X"50",X"32",X"5F",X"50",X"3E",X"27",X"32",X"5D",X"50",X"3E",X"04",X"C3",X"9F",X"2C",
		X"00",X"FE",X"12",X"D2",X"5F",X"3C",X"06",X"04",X"21",X"50",X"50",X"7E",X"C6",X"08",X"93",X"FE",
		X"11",X"38",X"07",X"23",X"23",X"23",X"23",X"10",X"F2",X"C9",X"23",X"23",X"23",X"7E",X"C6",X"02",
		X"92",X"FE",X"0D",X"30",X"F1",X"2B",X"2B",X"7E",X"E6",X"7F",X"FE",X"28",X"28",X"E6",X"3E",X"60",
		X"32",X"40",X"40",X"2B",X"36",X"F9",X"18",X"DB",X"2A",X"02",X"41",X"E5",X"11",X"F4",X"07",X"19",
		X"CD",X"64",X"08",X"7E",X"FE",X"20",X"38",X"0C",X"FE",X"28",X"38",X"37",X"FE",X"E1",X"38",X"04",
		X"FE",X"E8",X"38",X"2F",X"C3",X"D3",X"87",X"FE",X"14",X"20",X"2F",X"7E",X"D6",X"B8",X"FE",X"04",
		X"00",X"38",X"20",X"D1",X"06",X"03",X"21",X"50",X"50",X"7E",X"C6",X"10",X"93",X"FE",X"18",X"38",
		X"07",X"23",X"23",X"23",X"23",X"10",X"F2",X"C9",X"23",X"23",X"23",X"7E",X"92",X"FE",X"0C",X"30",
		X"F3",X"18",X"01",X"E1",X"3E",X"01",X"32",X"14",X"40",X"C9",X"FE",X"0C",X"30",X"44",X"D1",X"3A",
		X"50",X"50",X"C6",X"10",X"93",X"FE",X"18",X"30",X"08",X"3A",X"53",X"50",X"92",X"FE",X"0C",X"38",
		X"E3",X"3A",X"54",X"50",X"C6",X"10",X"93",X"FE",X"18",X"30",X"0A",X"3A",X"57",X"50",X"C6",X"0A",
		X"92",X"FE",X"0E",X"38",X"CF",X"3A",X"58",X"50",X"C6",X"10",X"93",X"FE",X"18",X"D0",X"3A",X"5B",
		X"50",X"C6",X"0A",X"92",X"FE",X"16",X"D0",X"3A",X"59",X"50",X"D6",X"08",X"28",X"B6",X"3D",X"C0",
		X"18",X"B2",X"E1",X"C9",X"00",X"A7",X"28",X"6C",X"FE",X"12",X"30",X"2B",X"7E",X"FE",X"83",X"38",
		X"04",X"FE",X"88",X"38",X"9E",X"D1",X"06",X"04",X"21",X"50",X"50",X"7E",X"C6",X"11",X"93",X"FE",
		X"15",X"38",X"07",X"23",X"23",X"23",X"23",X"10",X"F2",X"C9",X"23",X"C3",X"EE",X"89",X"C6",X"09",
		X"92",X"FE",X"13",X"30",X"F1",X"18",X"C9",X"D1",X"06",X"04",X"21",X"51",X"50",X"7E",X"D6",X"2E",
		X"28",X"21",X"3D",X"28",X"1E",X"2B",X"7E",X"C6",X"15",X"93",X"FE",X"22",X"30",X"10",X"23",X"23",
		X"23",X"7E",X"C6",X"0A",X"92",X"FE",X"0E",X"38",X"A7",X"23",X"23",X"10",X"E0",X"C9",X"23",X"23",
		X"23",X"18",X"F6",X"2B",X"7E",X"C6",X"13",X"93",X"FE",X"18",X"30",X"F2",X"23",X"23",X"23",X"7E",
		X"C6",X"05",X"18",X"E0",X"E1",X"C9",X"31",X"00",X"48",X"3E",X"04",X"32",X"05",X"50",X"3E",X"01",
		X"32",X"03",X"50",X"32",X"01",X"50",X"32",X"3F",X"50",X"C3",X"C3",X"A7",X"00",X"00",X"00",X"CD",
		X"C8",X"80",X"3A",X"14",X"40",X"A7",X"C8",X"00",X"00",X"00",X"3A",X"07",X"41",X"E6",X"08",X"28",
		X"04",X"F1",X"C3",X"38",X"82",X"3A",X"00",X"42",X"CD",X"CE",X"13",X"AF",X"32",X"14",X"40",X"C9",
		X"21",X"17",X"42",X"3A",X"00",X"60",X"E6",X"01",X"28",X"19",X"7E",X"A7",X"C8",X"36",X"00",X"2E",
		X"14",X"7E",X"3C",X"FE",X"0A",X"20",X"0F",X"36",X"00",X"23",X"7E",X"3C",X"FE",X"0A",X"20",X"06",
		X"36",X"00",X"C9",X"36",X"01",X"C9",X"77",X"C9",X"AF",X"32",X"06",X"70",X"32",X"07",X"70",X"CD",
		X"00",X"A5",X"CD",X"55",X"8A",X"3E",X"08",X"32",X"07",X"41",X"21",X"00",X"50",X"06",X"20",X"36",
		X"00",X"23",X"23",X"10",X"FA",X"CD",X"28",X"87",X"C3",X"DA",X"97",X"33",X"4B",X"8E",X"8D",X"8B",
		X"98",X"5E",X"01",X"5E",X"8F",X"8B",X"80",X"98",X"84",X"91",X"5E",X"81",X"94",X"93",X"93",X"8E",
		X"8D",X"FF",X"31",X"4A",X"8F",X"94",X"92",X"87",X"FF",X"53",X"4B",X"01",X"5E",X"8E",X"91",X"5E",
		X"02",X"5E",X"8F",X"8B",X"80",X"98",X"84",X"91",X"92",X"5E",X"81",X"94",X"93",X"93",X"8E",X"8D",
		X"FF",X"3E",X"01",X"32",X"06",X"60",X"32",X"04",X"60",X"AF",X"32",X"02",X"60",X"32",X"03",X"60",
		X"C9",X"3A",X"07",X"41",X"E6",X"08",X"C8",X"2A",X"14",X"42",X"7C",X"B5",X"C8",X"F1",X"CD",X"00",
		X"83",X"CD",X"91",X"82",X"3A",X"15",X"42",X"A7",X"20",X"18",X"3A",X"14",X"42",X"3D",X"20",X"12",
		X"21",X"5B",X"82",X"CD",X"17",X"0A",X"CD",X"B6",X"1F",X"3A",X"00",X"68",X"E6",X"01",X"28",X"E5",
		X"18",X"10",X"21",X"72",X"82",X"CD",X"17",X"0A",X"CD",X"B6",X"1F",X"3A",X"00",X"68",X"E6",X"03",
		X"28",X"F6",X"32",X"18",X"42",X"E6",X"02",X"28",X"03",X"CD",X"19",X"83",X"CD",X"19",X"83",X"CD",
		X"3B",X"8A",X"CD",X"24",X"00",X"C3",X"4A",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"21",X"40",X"50",X"06",X"08",X"36",X"00",X"23",X"23",X"23",X"23",X"10",X"F8",X"2E",X"06",X"06",
		X"36",X"36",X"00",X"23",X"10",X"FB",X"C3",X"3F",X"0D",X"21",X"14",X"42",X"7E",X"A7",X"20",X"09",
		X"23",X"7E",X"A7",X"C8",X"35",X"2B",X"36",X"09",X"C9",X"35",X"C9",X"36",X"0B",X"A7",X"ED",X"52",
		X"36",X"0A",X"ED",X"52",X"3D",X"20",X"F4",X"C9",X"CD",X"3F",X"0D",X"3A",X"00",X"70",X"CD",X"03",
		X"88",X"00",X"32",X"19",X"42",X"47",X"3A",X"18",X"42",X"E6",X"02",X"28",X"01",X"78",X"32",X"1A",
		X"42",X"11",X"20",X"00",X"3A",X"19",X"42",X"A7",X"28",X"09",X"3D",X"28",X"06",X"21",X"A2",X"4B",
		X"CD",X"2B",X"83",X"3A",X"1A",X"42",X"A7",X"C8",X"3D",X"C8",X"21",X"62",X"49",X"C3",X"2B",X"83",
		X"DE",X"04",X"9A",X"05",X"07",X"06",X"66",X"06",X"66",X"06",X"66",X"06",X"66",X"06",X"66",X"06",
		X"66",X"06",X"CB",X"06",X"16",X"07",X"16",X"07",X"16",X"07",X"26",X"07",X"26",X"07",X"C9",X"07",
		X"C9",X"07",X"C9",X"07",X"C9",X"07",X"7F",X"24",X"1A",X"25",X"57",X"25",X"B9",X"25",X"D9",X"25",
		X"D9",X"25",X"B9",X"25",X"F9",X"25",X"F9",X"25",X"F9",X"25",X"F9",X"25",X"F9",X"25",X"F9",X"25",
		X"F9",X"25",X"F9",X"25",X"6C",X"4A",X"86",X"80",X"8C",X"84",X"5E",X"8E",X"95",X"84",X"91",X"FF",
		X"21",X"02",X"48",X"11",X"20",X"00",X"06",X"20",X"36",X"5E",X"19",X"10",X"FB",X"C3",X"51",X"83",
		X"CD",X"28",X"87",X"00",X"00",X"AF",X"32",X"04",X"70",X"C9",X"06",X"EF",X"C5",X"CD",X"6B",X"19",
		X"CD",X"D2",X"1B",X"C1",X"10",X"F6",X"C9",X"2A",X"00",X"41",X"22",X"26",X"41",X"2A",X"02",X"41",
		X"22",X"28",X"41",X"3A",X"04",X"41",X"32",X"2A",X"41",X"3A",X"07",X"41",X"32",X"2B",X"41",X"3A",
		X"0C",X"41",X"32",X"2C",X"41",X"3A",X"17",X"41",X"32",X"4C",X"41",X"2A",X"1F",X"41",X"22",X"2D",
		X"41",X"2A",X"14",X"41",X"22",X"4A",X"41",X"11",X"2F",X"41",X"21",X"07",X"50",X"06",X"1B",X"7E",
		X"12",X"23",X"23",X"13",X"10",X"F9",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"21",X"07",X"41",X"CB",X"C6",X"3A",X"00",X"60",X"E6",X"20",X"C8",X"3E",X"01",X"32",X"07",X"70",
		X"32",X"06",X"70",X"C9",X"CD",X"6B",X"A2",X"CD",X"C3",X"9C",X"CD",X"91",X"82",X"21",X"B4",X"83",
		X"CD",X"1B",X"0A",X"C9",X"00",X"21",X"06",X"50",X"06",X"1B",X"36",X"00",X"23",X"23",X"10",X"FA",
		X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CD",X"C8",X"80",X"3A",X"1B",X"42",X"A7",X"28",X"09",X"3D",X"32",X"1B",X"42",X"AF",X"32",X"14",
		X"40",X"C9",X"C3",X"E0",X"89",X"A7",X"C8",X"CD",X"18",X"9D",X"F1",X"3A",X"07",X"41",X"CB",X"5F",
		X"C2",X"38",X"82",X"0F",X"38",X"5D",X"21",X"19",X"42",X"CD",X"0B",X"88",X"00",X"28",X"72",X"3A",
		X"18",X"42",X"E6",X"02",X"28",X"06",X"3A",X"1A",X"42",X"A7",X"20",X"77",X"CD",X"C0",X"83",X"3A",
		X"15",X"41",X"FE",X"14",X"20",X"07",X"3A",X"00",X"41",X"C3",X"2D",X"88",X"00",X"3E",X"60",X"32",
		X"1B",X"42",X"C3",X"90",X"37",X"21",X"02",X"20",X"22",X"00",X"41",X"CD",X"55",X"84",X"CD",X"12",
		X"9D",X"21",X"39",X"B7",X"22",X"02",X"41",X"3E",X"75",X"32",X"04",X"41",X"3E",X"01",X"32",X"02",
		X"60",X"32",X"04",X"60",X"AF",X"32",X"06",X"60",X"32",X"03",X"60",X"CD",X"00",X"8C",X"06",X"60",
		X"C3",X"3B",X"87",X"21",X"1A",X"42",X"CD",X"0B",X"88",X"00",X"20",X"0C",X"CD",X"DE",X"A0",X"3A",
		X"19",X"42",X"A7",X"20",X"09",X"C3",X"38",X"82",X"3A",X"19",X"42",X"A7",X"28",X"9E",X"AF",X"18",
		X"18",X"CD",X"D6",X"A0",X"3A",X"18",X"42",X"E6",X"02",X"CA",X"38",X"82",X"3A",X"1A",X"42",X"A7",
		X"CA",X"38",X"82",X"3A",X"28",X"41",X"A7",X"28",X"5D",X"08",X"11",X"26",X"43",X"21",X"26",X"41",
		X"01",X"27",X"00",X"ED",X"B0",X"CD",X"E7",X"83",X"21",X"50",X"50",X"06",X"04",X"36",X"F8",X"23",
		X"23",X"23",X"23",X"10",X"F8",X"2A",X"28",X"43",X"22",X"02",X"41",X"3A",X"2A",X"43",X"32",X"04",
		X"41",X"3A",X"2B",X"43",X"32",X"07",X"41",X"3A",X"2C",X"43",X"32",X"0C",X"41",X"2A",X"26",X"43",
		X"22",X"00",X"41",X"2A",X"2D",X"43",X"CD",X"47",X"2C",X"2A",X"4A",X"43",X"CD",X"97",X"87",X"11",
		X"07",X"50",X"21",X"2F",X"43",X"06",X"1B",X"7E",X"12",X"23",X"13",X"13",X"10",X"F9",X"08",X"28",
		X"0D",X"CD",X"30",X"84",X"18",X"14",X"CD",X"E7",X"83",X"CD",X"EA",X"9C",X"18",X"49",X"21",X"07",
		X"41",X"CB",X"86",X"AF",X"32",X"06",X"70",X"32",X"07",X"70",X"CD",X"08",X"36",X"3A",X"2E",X"43",
		X"A7",X"20",X"25",X"3A",X"4B",X"43",X"FE",X"14",X"20",X"2A",X"CD",X"90",X"87",X"FE",X"3C",X"30",
		X"06",X"CD",X"D0",X"83",X"C3",X"C5",X"84",X"D6",X"1E",X"32",X"00",X"41",X"CD",X"D0",X"83",X"CD",
		X"55",X"84",X"CD",X"DA",X"83",X"C3",X"DC",X"84",X"FE",X"03",X"30",X"71",X"C3",X"5D",X"88",X"00",
		X"00",X"00",X"00",X"00",X"A7",X"20",X"14",X"21",X"06",X"50",X"06",X"36",X"36",X"00",X"23",X"10",
		X"FB",X"AF",X"CD",X"93",X"82",X"CD",X"34",X"00",X"C3",X"00",X"87",X"3D",X"CD",X"61",X"87",X"32",
		X"15",X"41",X"07",X"C6",X"70",X"6F",X"26",X"83",X"7E",X"32",X"00",X"41",X"23",X"7E",X"32",X"01",
		X"41",X"CD",X"55",X"84",X"C3",X"35",X"88",X"CD",X"20",X"88",X"2A",X"00",X"41",X"EB",X"2A",X"26",
		X"43",X"A7",X"ED",X"52",X"C2",X"07",X"86",X"3A",X"15",X"41",X"47",X"3A",X"4B",X"43",X"90",X"C2",
		X"07",X"86",X"3A",X"20",X"41",X"A7",X"28",X"0A",X"FE",X"12",X"30",X"0D",X"AF",X"32",X"04",X"70",
		X"18",X"2E",X"3A",X"15",X"41",X"FE",X"14",X"28",X"F3",X"3E",X"01",X"18",X"F0",X"FE",X"12",X"30",
		X"09",X"3D",X"32",X"20",X"41",X"07",X"C6",X"92",X"18",X"AB",X"3E",X"20",X"32",X"23",X"41",X"CD",
		X"55",X"84",X"CD",X"E1",X"88",X"06",X"00",X"C5",X"CD",X"80",X"35",X"C1",X"10",X"F9",X"18",X"D9",
		X"CD",X"28",X"87",X"3E",X"17",X"32",X"49",X"50",X"06",X"08",X"CD",X"56",X"0D",X"C3",X"BD",X"84",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CD",X"3F",X"0D",X"CD",X"08",X"36",X"21",X"60",X"04",X"22",X"00",X"41",X"21",X"89",X"00",X"22",
		X"14",X"41",X"6C",X"22",X"1F",X"41",X"CD",X"28",X"87",X"21",X"19",X"47",X"22",X"02",X"41",X"3E",
		X"80",X"32",X"04",X"41",X"C3",X"63",X"0D",X"00",X"21",X"00",X"40",X"06",X"00",X"36",X"00",X"23",
		X"10",X"FB",X"C9",X"3E",X"01",X"32",X"04",X"70",X"C3",X"0B",X"19",X"CD",X"56",X"0D",X"3E",X"60",
		X"32",X"1B",X"42",X"C3",X"A5",X"8A",X"FE",X"A7",X"20",X"06",X"3E",X"89",X"32",X"14",X"41",X"C9",
		X"FE",X"D2",X"20",X"F8",X"3E",X"B3",X"18",X"F4",X"3E",X"17",X"32",X"49",X"50",X"C3",X"74",X"2C",
		X"00",X"F5",X"FE",X"02",X"3E",X"89",X"38",X"02",X"3E",X"B3",X"32",X"14",X"41",X"F1",X"C9",X"21",
		X"37",X"50",X"06",X"03",X"36",X"04",X"23",X"23",X"10",X"FA",X"21",X"1B",X"48",X"11",X"20",X"00",
		X"0E",X"03",X"E5",X"06",X"20",X"36",X"DE",X"19",X"10",X"FB",X"E1",X"23",X"0D",X"20",X"F3",X"C9",
		X"CD",X"87",X"88",X"3A",X"26",X"43",X"C9",X"22",X"14",X"41",X"3A",X"4C",X"43",X"32",X"17",X"41",
		X"C9",X"3E",X"C7",X"32",X"53",X"50",X"32",X"57",X"50",X"3A",X"44",X"50",X"C9",X"32",X"50",X"50",
		X"32",X"5C",X"50",X"CD",X"28",X"87",X"3E",X"01",X"32",X"04",X"70",X"C9",X"3E",X"01",X"32",X"04",
		X"70",X"3A",X"21",X"41",X"C9",X"AF",X"32",X"04",X"70",X"C3",X"8F",X"1A",X"AF",X"32",X"04",X"70",
		X"C3",X"98",X"3D",X"3A",X"20",X"41",X"A7",X"C2",X"68",X"81",X"3A",X"15",X"41",X"C3",X"E7",X"80",
		X"00",X"00",X"00",X"00",X"00",X"CD",X"AC",X"31",X"3A",X"59",X"50",X"FE",X"A8",X"C0",X"C3",X"0C",
		X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"60",X"C9",X"E6",X"03",X"20",X"01",X"3C",X"C6",X"02",X"C9",X"3A",X"00",X"70",X"E6",X"03",
		X"28",X"02",X"35",X"C9",X"3D",X"C9",X"3A",X"4A",X"40",X"A7",X"CA",X"CB",X"17",X"C3",X"EA",X"11",
		X"3E",X"01",X"32",X"4A",X"40",X"CD",X"6A",X"31",X"AF",X"32",X"4A",X"40",X"C9",X"FE",X"3C",X"D2",
		X"3E",X"87",X"C3",X"C5",X"84",X"CD",X"87",X"88",X"3A",X"20",X"41",X"A7",X"CA",X"07",X"86",X"3A",
		X"2E",X"43",X"47",X"C5",X"CD",X"74",X"88",X"C1",X"3A",X"20",X"41",X"B8",X"20",X"F5",X"2A",X"00",
		X"41",X"EB",X"2A",X"26",X"43",X"A7",X"ED",X"52",X"20",X"E9",X"C3",X"22",X"86",X"3E",X"02",X"32",
		X"2E",X"43",X"32",X"20",X"41",X"21",X"F0",X"23",X"22",X"00",X"41",X"21",X"25",X"24",X"22",X"26",
		X"43",X"C3",X"01",X"86",X"3A",X"20",X"41",X"FE",X"05",X"D2",X"E5",X"87",X"C3",X"93",X"31",X"3A",
		X"20",X"41",X"A7",X"C0",X"C3",X"C1",X"2C",X"CD",X"68",X"89",X"2A",X"02",X"41",X"CD",X"B1",X"02",
		X"3A",X"20",X"41",X"A7",X"20",X"47",X"3A",X"4B",X"43",X"FE",X"04",X"38",X"05",X"CD",X"6F",X"87",
		X"18",X"03",X"CD",X"E1",X"0A",X"3A",X"4B",X"43",X"FE",X"14",X"20",X"0D",X"11",X"50",X"50",X"21",
		X"00",X"2C",X"01",X"0F",X"00",X"ED",X"B0",X"18",X"10",X"21",X"0C",X"07",X"22",X"51",X"50",X"2E",
		X"0A",X"22",X"55",X"50",X"2E",X"08",X"22",X"59",X"50",X"3A",X"4B",X"43",X"FE",X"0B",X"38",X"08",
		X"CD",X"91",X"82",X"AF",X"32",X"06",X"60",X"C9",X"AF",X"CD",X"93",X"82",X"C9",X"FE",X"12",X"38",
		X"4E",X"3E",X"01",X"32",X"37",X"50",X"3E",X"03",X"32",X"39",X"50",X"32",X"3B",X"50",X"11",X"20",
		X"00",X"21",X"1B",X"48",X"E5",X"06",X"20",X"36",X"A4",X"19",X"10",X"FB",X"E1",X"23",X"0E",X"AE",
		X"3E",X"02",X"E5",X"06",X"20",X"71",X"19",X"10",X"FC",X"E1",X"23",X"0C",X"3D",X"20",X"F3",X"CD",
		X"A0",X"36",X"3A",X"20",X"41",X"FE",X"18",X"38",X"03",X"CD",X"14",X"39",X"2A",X"02",X"41",X"7D",
		X"CD",X"3A",X"02",X"3E",X"04",X"32",X"46",X"50",X"21",X"1B",X"48",X"3E",X"01",X"18",X"10",X"CD",
		X"6F",X"87",X"21",X"22",X"02",X"22",X"51",X"50",X"CD",X"DE",X"9C",X"21",X"0B",X"48",X"AF",X"32",
		X"02",X"60",X"22",X"21",X"41",X"AF",X"32",X"06",X"60",X"3E",X"01",X"32",X"03",X"60",X"32",X"04",
		X"60",X"C9",X"7C",X"FE",X"25",X"C2",X"91",X"30",X"79",X"FE",X"06",X"C3",X"83",X"30",X"7C",X"FE",
		X"25",X"C2",X"91",X"30",X"23",X"C3",X"79",X"30",X"CD",X"0A",X"9D",X"FE",X"2F",X"C0",X"3E",X"04",
		X"32",X"41",X"50",X"3C",X"32",X"45",X"50",X"C9",X"32",X"50",X"50",X"32",X"5C",X"50",X"00",X"00",
		X"00",X"3E",X"01",X"32",X"04",X"70",X"01",X"06",X"50",X"21",X"C3",X"4B",X"CD",X"CB",X"0A",X"01",
		X"10",X"02",X"CD",X"45",X"0D",X"C9",X"3E",X"F8",X"32",X"50",X"50",X"32",X"54",X"50",X"32",X"58",
		X"50",X"32",X"5C",X"50",X"C9",X"33",X"4A",X"91",X"84",X"8F",X"8B",X"80",X"98",X"FF",X"CD",X"00",
		X"83",X"CD",X"91",X"82",X"21",X"A5",X"89",X"CD",X"1B",X"0A",X"06",X"F0",X"CD",X"56",X"0D",X"AF",
		X"32",X"0C",X"41",X"32",X"17",X"41",X"3A",X"07",X"41",X"E6",X"01",X"C6",X"50",X"6F",X"26",X"41",
		X"34",X"C3",X"D7",X"85",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3A",X"41",X"50",X"FE",X"3E",X"CA",X"7D",X"84",X"3A",X"14",X"40",X"C3",X"85",X"84",X"7E",X"FE",
		X"28",X"CA",X"84",X"81",X"FE",X"A8",X"CA",X"84",X"81",X"23",X"23",X"7E",X"C3",X"8E",X"81",X"00",
		X"22",X"00",X"41",X"2A",X"53",X"03",X"EB",X"2A",X"D6",X"8D",X"19",X"EB",X"2A",X"3A",X"42",X"19",
		X"11",X"29",X"53",X"A7",X"ED",X"52",X"C9",X"C3",X"E0",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"02",X"42",X"06",X"06",
		X"36",X"00",X"23",X"10",X"FB",X"3A",X"18",X"42",X"E6",X"02",X"00",X"2E",X"0E",X"06",X"06",X"36",
		X"00",X"23",X"10",X"FB",X"C9",X"CD",X"24",X"00",X"AF",X"32",X"18",X"42",X"C3",X"3B",X"8A",X"32",
		X"49",X"40",X"0E",X"03",X"C3",X"64",X"2C",X"E1",X"E5",X"11",X"F3",X"10",X"19",X"CD",X"64",X"08",
		X"7E",X"FE",X"8D",X"38",X"23",X"FE",X"90",X"38",X"12",X"FE",X"A0",X"38",X"1B",X"FE",X"A6",X"30",
		X"17",X"0E",X"08",X"FE",X"A3",X"30",X"06",X"0E",X"05",X"18",X"02",X"0E",X"14",X"C3",X"67",X"37",
		X"CD",X"00",X"0E",X"3E",X"74",X"32",X"04",X"41",X"C3",X"D3",X"02",X"00",X"3A",X"00",X"42",X"E6",
		X"E0",X"C0",X"C3",X"BE",X"3F",X"21",X"00",X"2C",X"11",X"50",X"50",X"01",X"10",X"00",X"ED",X"B0",
		X"C3",X"96",X"37",X"79",X"3D",X"28",X"05",X"3D",X"18",X"05",X"7B",X"C9",X"3E",X"32",X"C9",X"3E",
		X"34",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"01",X"01",X"01",X"02",X"02",X"02",X"02",
		X"02",X"03",X"03",X"03",X"04",X"04",X"04",X"06",X"06",X"06",X"06",X"08",X"08",X"08",X"08",X"08",
		X"08",X"08",X"08",X"08",X"08",X"0A",X"0A",X"0A",X"0A",X"0A",X"00",X"3A",X"41",X"50",X"4F",X"3E",
		X"3A",X"32",X"41",X"50",X"3C",X"CD",X"00",X"97",X"06",X"08",X"E5",X"CD",X"56",X"0D",X"E1",X"79",
		X"32",X"41",X"50",X"3C",X"32",X"45",X"50",X"C9",X"00",X"00",X"3A",X"20",X"41",X"A7",X"28",X"06",
		X"FE",X"12",X"38",X"25",X"18",X"07",X"3A",X"15",X"41",X"FE",X"14",X"20",X"1C",X"3A",X"41",X"50",
		X"5F",X"3E",X"3A",X"0E",X"04",X"32",X"41",X"50",X"3C",X"32",X"45",X"50",X"06",X"10",X"CD",X"56",
		X"0D",X"0D",X"28",X"41",X"CD",X"B3",X"8A",X"18",X"EC",X"3A",X"41",X"50",X"5F",X"3E",X"3A",X"0E",
		X"04",X"06",X"10",X"32",X"41",X"50",X"3C",X"32",X"45",X"50",X"21",X"43",X"50",X"7E",X"FE",X"C7",
		X"30",X"04",X"34",X"2E",X"47",X"34",X"C5",X"06",X"01",X"CD",X"56",X"0D",X"C1",X"10",X"EB",X"0D",
		X"28",X"05",X"CD",X"B3",X"8A",X"18",X"DA",X"3A",X"43",X"50",X"FE",X"C7",X"30",X"04",X"0C",X"04",
		X"18",X"D8",X"32",X"03",X"41",X"06",X"60",X"CD",X"56",X"0D",X"C9",X"CD",X"51",X"2C",X"0F",X"3A",
		X"00",X"68",X"38",X"03",X"3A",X"00",X"60",X"CB",X"57",X"28",X"13",X"E5",X"2D",X"11",X"E9",X"0C",
		X"E5",X"19",X"CD",X"64",X"08",X"7E",X"E1",X"FE",X"E0",X"20",X"0E",X"E1",X"18",X"0C",X"E6",X"08",
		X"28",X"08",X"E5",X"2C",X"11",X"00",X"0D",X"18",X"E7",X"F1",X"C3",X"62",X"2D",X"00",X"00",X"00",
		X"CD",X"CF",X"12",X"2A",X"02",X"41",X"CD",X"A2",X"01",X"3A",X"50",X"40",X"A7",X"20",X"0F",X"3A",
		X"01",X"41",X"FE",X"3C",X"D2",X"57",X"9B",X"45",X"CD",X"D3",X"01",X"68",X"18",X"10",X"24",X"FE",
		X"A0",X"30",X"06",X"25",X"25",X"3C",X"32",X"50",X"40",X"3E",X"00",X"CD",X"B4",X"9C",X"E5",X"F5",
		X"11",X"F7",X"00",X"19",X"CD",X"64",X"08",X"7E",X"FE",X"E0",X"CA",X"A9",X"8C",X"23",X"23",X"7E",
		X"FE",X"90",X"28",X"0C",X"FE",X"91",X"00",X"00",X"FE",X"9A",X"28",X"04",X"FE",X"9B",X"20",X"03",
		X"C3",X"BE",X"1B",X"FE",X"E0",X"28",X"72",X"C3",X"20",X"9D",X"00",X"20",X"20",X"CB",X"57",X"28",
		X"46",X"E5",X"2D",X"11",X"E9",X"0C",X"19",X"CD",X"64",X"08",X"7E",X"FE",X"E0",X"28",X"3B",X"E1",
		X"7D",X"FE",X"39",X"30",X"31",X"FE",X"29",X"38",X"72",X"3E",X"01",X"18",X"21",X"E5",X"2C",X"11",
		X"00",X"0D",X"19",X"CD",X"64",X"08",X"7E",X"FE",X"E0",X"28",X"1F",X"E1",X"7D",X"FE",X"B1",X"38",
		X"12",X"FE",X"DF",X"30",X"56",X"3A",X"00",X"41",X"FE",X"91",X"30",X"07",X"3E",X"00",X"32",X"20",
		X"40",X"18",X"48",X"2C",X"18",X"45",X"2D",X"18",X"42",X"F1",X"3E",X"9D",X"32",X"04",X"41",X"E1",
		X"3E",X"03",X"C3",X"9E",X"8C",X"11",X"F3",X"10",X"19",X"CD",X"64",X"08",X"7E",X"FE",X"E0",X"28",
		X"09",X"06",X"01",X"CD",X"B8",X"1B",X"E1",X"18",X"E7",X"F1",X"11",X"20",X"00",X"2B",X"2B",X"06",
		X"03",X"19",X"7E",X"FE",X"7C",X"28",X"2A",X"FE",X"7E",X"28",X"23",X"C3",X"0C",X"1F",X"00",X"00",
		X"E1",X"3E",X"73",X"32",X"04",X"41",X"3E",X"0F",X"32",X"08",X"41",X"7D",X"FE",X"29",X"30",X"06",
		X"3E",X"29",X"6F",X"C3",X"3A",X"02",X"FE",X"DE",X"38",X"F9",X"3E",X"DE",X"18",X"F4",X"CD",X"3C",
		X"0E",X"36",X"5E",X"19",X"36",X"5E",X"23",X"E5",X"01",X"28",X"04",X"3A",X"01",X"41",X"FE",X"0A",
		X"38",X"11",X"01",X"1E",X"03",X"FE",X"1A",X"38",X"0A",X"01",X"14",X"02",X"FE",X"2A",X"28",X"03",
		X"01",X"0A",X"01",X"70",X"CD",X"3C",X"0E",X"36",X"00",X"CD",X"3C",X"0E",X"36",X"00",X"CD",X"6C",
		X"2C",X"E1",X"EB",X"7B",X"E6",X"1F",X"C6",X"C0",X"6F",X"26",X"4B",X"01",X"3A",X"50",X"D5",X"CD",
		X"CB",X"0A",X"D1",X"A7",X"ED",X"52",X"7D",X"07",X"07",X"07",X"4F",X"7C",X"E6",X"03",X"07",X"07",
		X"07",X"81",X"4F",X"3A",X"00",X"41",X"81",X"21",X"00",X"22",X"06",X"21",X"23",X"23",X"BE",X"28",
		X"04",X"10",X"F9",X"18",X"04",X"26",X"44",X"36",X"01",X"E1",X"7C",X"3C",X"E6",X"F8",X"67",X"C3",
		X"E1",X"8C",X"11",X"FF",X"FF",X"C5",X"7E",X"AB",X"47",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"A8",
		X"4F",X"0F",X"0F",X"0F",X"47",X"E6",X"1F",X"AA",X"5F",X"78",X"E6",X"E0",X"A9",X"57",X"78",X"0F",
		X"E6",X"F0",X"AB",X"5F",X"23",X"C1",X"78",X"BC",X"D8",X"20",X"DA",X"79",X"BD",X"D8",X"18",X"D5",
		X"2A",X"58",X"41",X"06",X"04",X"7E",X"10",X"FD",X"3A",X"3B",X"42",X"86",X"FE",X"5F",X"C9",X"C3",
		X"F0",X"0C",X"2A",X"A0",X"8D",X"EB",X"2A",X"AD",X"8D",X"19",X"7C",X"85",X"FE",X"A9",X"C3",X"6A",
		X"31",X"C3",X"30",X"0E",X"3A",X"0E",X"40",X"A7",X"C0",X"2A",X"58",X"41",X"7E",X"2E",X"14",X"46",
		X"4E",X"3A",X"3A",X"42",X"86",X"D6",X"DD",X"18",X"04",X"32",X"0C",X"41",X"C9",X"3A",X"0E",X"40",
		X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"3A",X"07",X"41",X"E6",X"08",X"28",X"0B",X"CD",X"C9",X"9C",X"06",X"1E",X"36",X"00",
		X"23",X"10",X"FB",X"C9",X"11",X"03",X"68",X"21",X"63",X"40",X"7E",X"A7",X"28",X"07",X"35",X"3E",
		X"01",X"20",X"01",X"AF",X"12",X"23",X"CD",X"18",X"A0",X"00",X"00",X"00",X"3A",X"66",X"40",X"A7",
		X"CA",X"6F",X"92",X"3C",X"FE",X"03",X"20",X"01",X"AF",X"32",X"66",X"40",X"28",X"02",X"3E",X"01",
		X"32",X"05",X"68",X"C3",X"6F",X"92",X"00",X"3A",X"04",X"41",X"BE",X"28",X"0E",X"77",X"23",X"FE",
		X"76",X"38",X"0C",X"FE",X"7D",X"38",X"0C",X"FE",X"90",X"30",X"0D",X"3E",X"FE",X"18",X"0D",X"3E",
		X"10",X"18",X"08",X"7E",X"C6",X"10",X"18",X"03",X"7E",X"D6",X"08",X"77",X"32",X"00",X"78",X"3A",
		X"67",X"40",X"A7",X"28",X"68",X"21",X"00",X"58",X"11",X"00",X"59",X"3C",X"32",X"67",X"40",X"FE",
		X"02",X"28",X"29",X"FE",X"15",X"28",X"42",X"FE",X"80",X"28",X"44",X"3A",X"68",X"40",X"D6",X"06",
		X"4F",X"AF",X"12",X"3A",X"00",X"42",X"E6",X"02",X"28",X"04",X"79",X"C6",X"10",X"4F",X"71",X"3E",
		X"02",X"12",X"79",X"00",X"00",X"00",X"77",X"79",X"32",X"68",X"40",X"C9",X"3E",X"07",X"12",X"36",
		X"27",X"3C",X"12",X"36",X"0F",X"3C",X"12",X"36",X"0F",X"3E",X"01",X"12",X"36",X"01",X"3E",X"03",
		X"12",X"36",X"00",X"3E",X"10",X"32",X"68",X"40",X"C9",X"3E",X"07",X"12",X"36",X"3C",X"C9",X"3E",
		X"07",X"12",X"36",X"38",X"00",X"00",X"00",X"00",X"AF",X"32",X"67",X"40",X"C9",X"11",X"00",X"59",
		X"AF",X"12",X"2E",X"69",X"3A",X"0F",X"40",X"BE",X"28",X"1A",X"77",X"3A",X"53",X"50",X"47",X"00",
		X"00",X"0F",X"0F",X"80",X"21",X"00",X"58",X"77",X"3E",X"01",X"12",X"77",X"3E",X"08",X"12",X"36",
		X"0F",X"C3",X"8D",X"8F",X"3A",X"6A",X"40",X"A7",X"28",X"21",X"3D",X"32",X"6A",X"40",X"CB",X"67",
		X"20",X"08",X"E6",X"0F",X"07",X"07",X"C6",X"D6",X"18",X"06",X"E6",X"0F",X"47",X"3E",X"64",X"90",
		X"21",X"00",X"58",X"77",X"3E",X"01",X"12",X"36",X"00",X"18",X"D1",X"3A",X"6B",X"40",X"A7",X"28",
		X"1C",X"21",X"00",X"58",X"C6",X"30",X"38",X"08",X"77",X"3E",X"01",X"12",X"36",X"00",X"18",X"07",
		X"07",X"77",X"3E",X"01",X"12",X"36",X"01",X"AF",X"32",X"6B",X"40",X"18",X"AF",X"21",X"00",X"58",
		X"3A",X"6C",X"40",X"A7",X"28",X"17",X"3D",X"32",X"6C",X"40",X"28",X"18",X"FE",X"2F",X"28",X"1B",
		X"07",X"4F",X"3E",X"A0",X"91",X"77",X"3E",X"01",X"12",X"36",X"00",X"18",X"20",X"3E",X"08",X"12",
		X"36",X"00",X"18",X"19",X"3E",X"07",X"12",X"36",X"38",X"18",X"12",X"3E",X"0C",X"12",X"36",X"20",
		X"3C",X"12",X"36",X"09",X"3E",X"07",X"12",X"36",X"30",X"3C",X"12",X"36",X"10",X"3E",X"02",X"12",
		X"3A",X"6D",X"40",X"A7",X"28",X"20",X"D6",X"04",X"32",X"6D",X"40",X"FE",X"7C",X"20",X"14",X"77",
		X"3E",X"03",X"12",X"36",X"02",X"3E",X"0C",X"12",X"36",X"20",X"3C",X"12",X"36",X"09",X"3E",X"09",
		X"12",X"36",X"10",X"C3",X"17",X"90",X"3A",X"6E",X"40",X"A7",X"28",X"21",X"3D",X"32",X"6E",X"40",
		X"20",X"07",X"3E",X"07",X"12",X"36",X"38",X"18",X"EA",X"FE",X"0F",X"20",X"E6",X"3E",X"07",X"12",
		X"36",X"2A",X"3E",X"0C",X"12",X"36",X"01",X"3C",X"12",X"36",X"08",X"18",X"D1",X"3A",X"6F",X"40",
		X"A7",X"28",X"12",X"D6",X"20",X"32",X"6F",X"40",X"77",X"3E",X"03",X"12",X"36",X"00",X"3E",X"09",
		X"12",X"36",X"0F",X"18",X"22",X"3A",X"70",X"40",X"A7",X"CA",X"00",X"96",X"D6",X"17",X"77",X"3E",
		X"03",X"12",X"36",X"01",X"AF",X"32",X"70",X"40",X"18",X"E4",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"3E",X"09",X"12",X"36",X"00",X"3E",X"04",X"12",X"3A",X"62",X"40",X"A7",X"28",X"29",
		X"3D",X"32",X"62",X"40",X"FE",X"1F",X"20",X"10",X"3E",X"0C",X"12",X"36",X"20",X"3C",X"12",X"36",
		X"09",X"3E",X"0A",X"12",X"36",X"10",X"18",X"0E",X"E6",X"04",X"3E",X"39",X"20",X"02",X"3E",X"1C",
		X"77",X"3E",X"05",X"12",X"36",X"01",X"C3",X"FA",X"90",X"3A",X"43",X"40",X"47",X"3A",X"45",X"40",
		X"B0",X"28",X"21",X"3A",X"00",X"42",X"E6",X"03",X"28",X"08",X"FE",X"02",X"28",X"08",X"36",X"4C",
		X"18",X"06",X"36",X"71",X"18",X"02",X"36",X"39",X"3E",X"05",X"12",X"36",X"00",X"3E",X"0A",X"12",
		X"36",X"0F",X"18",X"D2",X"3A",X"47",X"40",X"47",X"3A",X"48",X"40",X"B0",X"28",X"23",X"3A",X"00",
		X"42",X"E6",X"3F",X"28",X"0C",X"E6",X"06",X"C6",X"30",X"77",X"3E",X"05",X"12",X"36",X"00",X"18",
		X"B5",X"3E",X"0C",X"12",X"36",X"20",X"3C",X"12",X"36",X"09",X"3E",X"0A",X"12",X"36",X"10",X"18",
		X"A5",X"E5",X"2A",X"3D",X"40",X"7E",X"E1",X"FE",X"93",X"20",X"1C",X"3A",X"20",X"41",X"FE",X"12",
		X"38",X"15",X"3A",X"00",X"42",X"E6",X"0F",X"20",X"8D",X"36",X"CF",X"3E",X"05",X"12",X"36",X"02",
		X"3E",X"0C",X"12",X"36",X"0C",X"18",X"CF",X"3A",X"71",X"40",X"A7",X"28",X"0F",X"D6",X"04",X"32",
		X"71",X"40",X"2F",X"77",X"3E",X"05",X"12",X"36",X"01",X"C3",X"6D",X"90",X"3A",X"72",X"40",X"A7",
		X"28",X"13",X"3D",X"32",X"72",X"40",X"C6",X"C9",X"4F",X"06",X"1B",X"0A",X"77",X"3E",X"05",X"12",
		X"36",X"00",X"C3",X"6D",X"90",X"3E",X"0A",X"12",X"36",X"00",X"3A",X"73",X"40",X"A7",X"28",X"0D",
		X"3D",X"32",X"73",X"40",X"28",X"02",X"3E",X"01",X"32",X"00",X"60",X"18",X"11",X"3A",X"74",X"40",
		X"A7",X"28",X"0B",X"3D",X"32",X"74",X"40",X"28",X"02",X"3E",X"01",X"32",X"01",X"60",X"C9",X"00",
		X"00",X"3A",X"77",X"40",X"A7",X"28",X"05",X"3D",X"32",X"77",X"40",X"C9",X"3A",X"78",X"40",X"4F",
		X"C6",X"03",X"32",X"78",X"40",X"06",X"95",X"0A",X"FE",X"FF",X"20",X"07",X"AF",X"32",X"76",X"40",
		X"F1",X"F1",X"C9",X"CD",X"30",X"93",X"03",X"AF",X"12",X"0A",X"77",X"3E",X"01",X"12",X"03",X"0A",
		X"77",X"3E",X"0C",X"12",X"36",X"20",X"3C",X"12",X"36",X"09",X"3E",X"08",X"12",X"36",X"10",X"C9",
		X"3A",X"79",X"40",X"A7",X"28",X"05",X"3D",X"32",X"79",X"40",X"C9",X"3A",X"7A",X"40",X"4F",X"06",
		X"94",X"0A",X"CB",X"7F",X"20",X"16",X"32",X"79",X"40",X"03",X"3E",X"02",X"12",X"0A",X"77",X"3E",
		X"03",X"12",X"03",X"0A",X"77",X"3E",X"09",X"12",X"36",X"0F",X"18",X"0A",X"E6",X"7F",X"32",X"79",
		X"40",X"3E",X"09",X"12",X"36",X"00",X"79",X"3C",X"32",X"7A",X"40",X"C9",X"00",X"00",X"00",X"00",
		X"3A",X"76",X"40",X"A7",X"C8",X"21",X"00",X"58",X"11",X"00",X"59",X"3D",X"C2",X"33",X"92",X"CD",
		X"21",X"91",X"CD",X"60",X"91",X"3A",X"7B",X"40",X"A7",X"20",X"38",X"3A",X"7C",X"40",X"FE",X"00",
		X"20",X"02",X"3E",X"E0",X"4F",X"06",X"95",X"0A",X"CB",X"7F",X"20",X"16",X"32",X"7B",X"40",X"03",
		X"3E",X"04",X"12",X"0A",X"77",X"3E",X"05",X"12",X"03",X"0A",X"77",X"3E",X"0A",X"12",X"36",X"0F",
		X"18",X"0A",X"E6",X"7F",X"32",X"7B",X"40",X"3E",X"0A",X"12",X"36",X"00",X"79",X"3C",X"32",X"7C",
		X"40",X"18",X"04",X"3D",X"32",X"7B",X"40",X"3A",X"7D",X"40",X"A7",X"28",X"06",X"3D",X"32",X"7D",
		X"40",X"F1",X"C9",X"3A",X"7E",X"40",X"FE",X"DF",X"20",X"02",X"3E",X"D5",X"4F",X"06",X"95",X"0A",
		X"E6",X"3F",X"32",X"7D",X"40",X"0A",X"CB",X"7F",X"20",X"0B",X"CB",X"77",X"3E",X"01",X"20",X"09",
		X"32",X"00",X"60",X"18",X"07",X"AF",X"32",X"00",X"60",X"32",X"01",X"60",X"79",X"3C",X"32",X"7E",
		X"40",X"F1",X"C9",X"3D",X"20",X"08",X"CD",X"21",X"91",X"CD",X"67",X"9F",X"18",X"B9",X"CD",X"21",
		X"91",X"3A",X"79",X"40",X"A7",X"28",X"06",X"3D",X"32",X"79",X"40",X"18",X"AA",X"3A",X"7A",X"40",
		X"4F",X"C6",X"03",X"32",X"7A",X"40",X"06",X"94",X"0A",X"32",X"79",X"40",X"03",X"3E",X"02",X"12",
		X"0A",X"77",X"3E",X"03",X"12",X"03",X"0A",X"77",X"3E",X"09",X"12",X"36",X"10",X"18",X"88",X"3A",
		X"20",X"41",X"FE",X"12",X"18",X"2D",X"3A",X"00",X"42",X"0F",X"30",X"30",X"3A",X"00",X"68",X"E6",
		X"40",X"20",X"06",X"3A",X"07",X"41",X"0F",X"38",X"2B",X"3A",X"00",X"60",X"A7",X"28",X"08",X"E6",
		X"88",X"20",X"32",X"06",X"06",X"18",X"02",X"06",X"02",X"3A",X"65",X"40",X"4F",X"3D",X"FA",X"D3",
		X"92",X"18",X"2D",X"3A",X"04",X"41",X"BE",X"28",X"03",X"77",X"18",X"D0",X"3E",X"FF",X"32",X"00",
		X"78",X"C3",X"6F",X"8E",X"3A",X"00",X"60",X"E6",X"02",X"20",X"0A",X"3A",X"00",X"68",X"A7",X"28",
		X"D6",X"E6",X"08",X"28",X"CE",X"06",X"00",X"3A",X"65",X"40",X"4F",X"A7",X"20",X"1F",X"3E",X"0A",
		X"32",X"65",X"40",X"3A",X"00",X"42",X"A0",X"20",X"D3",X"06",X"9A",X"0A",X"47",X"3A",X"03",X"41",
		X"0F",X"0F",X"E6",X"3F",X"EE",X"3F",X"80",X"32",X"00",X"78",X"C3",X"6F",X"8E",X"3D",X"20",X"E0",
		X"18",X"E1",X"22",X"79",X"40",X"26",X"D5",X"22",X"7D",X"40",X"C9",X"00",X"00",X"00",X"00",X"00",
		X"CD",X"1B",X"0A",X"3E",X"01",X"32",X"76",X"40",X"21",X"00",X"00",X"22",X"77",X"40",X"21",X"00",
		X"00",X"22",X"79",X"40",X"21",X"00",X"E0",X"22",X"7B",X"40",X"21",X"00",X"D5",X"22",X"7D",X"40",
		X"3E",X"07",X"32",X"00",X"59",X"3E",X"38",X"32",X"00",X"58",X"06",X"F0",X"CD",X"56",X"0D",X"C9",
		X"32",X"77",X"40",X"FE",X"40",X"C0",X"3E",X"FF",X"32",X"7B",X"40",X"32",X"7D",X"40",X"C9",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CD",X"96",X"89",X"3E",X"02",X"32",X"76",X"40",X"21",
		X"00",X"28",X"22",X"77",X"40",X"21",X"00",X"34",X"22",X"79",X"40",X"21",X"00",X"D5",X"22",X"7D",
		X"40",X"C9",X"CD",X"56",X"0D",X"3E",X"03",X"32",X"76",X"40",X"21",X"00",X"9B",X"22",X"77",X"40",
		X"21",X"00",X"94",X"C3",X"F2",X"92",X"00",X"FE",X"7D",X"C8",X"FE",X"7F",X"C8",X"FE",X"F5",X"C8",
		X"FE",X"F7",X"C9",X"32",X"04",X"41",X"AF",X"32",X"6A",X"40",X"C3",X"4A",X"93",X"00",X"00",X"00",
		X"3A",X"00",X"42",X"E6",X"40",X"28",X"04",X"3A",X"02",X"41",X"C9",X"3A",X"02",X"41",X"D6",X"20",
		X"C9",X"11",X"20",X"00",X"3A",X"18",X"41",X"A7",X"C8",X"3A",X"15",X"41",X"FE",X"0A",X"30",X"05",
		X"AF",X"32",X"18",X"41",X"C9",X"0E",X"8F",X"C9",X"3A",X"7F",X"40",X"A7",X"CA",X"5A",X"96",X"3D",
		X"32",X"7F",X"40",X"FE",X"2F",X"20",X"11",X"3E",X"0C",X"12",X"36",X"28",X"3C",X"12",X"36",X"09",
		X"3E",X"09",X"12",X"36",X"10",X"C3",X"17",X"90",X"07",X"47",X"3A",X"00",X"42",X"E6",X"03",X"07",
		X"07",X"07",X"C6",X"C0",X"90",X"77",X"3E",X"03",X"12",X"36",X"00",X"C3",X"17",X"90",X"6F",X"06",
		X"06",X"1A",X"FE",X"80",X"C0",X"22",X"95",X"40",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"57",X"03",X"97",X"07",X"57",X"03",X"87",X"07",X"57",X"03",X"87",X"07",X"AC",X"01",X"97",
		X"07",X"AC",X"01",X"87",X"07",X"AC",X"01",X"87",X"07",X"57",X"03",X"97",X"07",X"57",X"03",X"87",
		X"07",X"57",X"03",X"87",X"07",X"AC",X"01",X"97",X"07",X"AC",X"01",X"87",X"07",X"AC",X"01",X"87",
		X"07",X"57",X"03",X"FF",X"07",X"3B",X"02",X"87",X"07",X"FA",X"02",X"87",X"07",X"3B",X"02",X"87",
		X"07",X"FA",X"02",X"87",X"07",X"3B",X"02",X"87",X"07",X"FA",X"02",X"87",X"07",X"3B",X"02",X"87",
		X"07",X"FA",X"02",X"87",X"07",X"FC",X"01",X"87",X"07",X"A7",X"02",X"87",X"07",X"FC",X"01",X"87",
		X"07",X"A7",X"02",X"87",X"07",X"FC",X"01",X"87",X"07",X"A7",X"02",X"87",X"07",X"FC",X"01",X"87",
		X"07",X"A7",X"02",X"87",X"07",X"3B",X"02",X"87",X"07",X"FA",X"02",X"87",X"07",X"3B",X"02",X"87",
		X"07",X"FA",X"02",X"87",X"07",X"3B",X"02",X"87",X"03",X"3B",X"02",X"83",X"03",X"3B",X"02",X"83",
		X"07",X"3B",X"02",X"FF",X"0F",X"57",X"03",X"0F",X"AC",X"01",X"0F",X"57",X"03",X"0F",X"AC",X"01",
		X"0F",X"AC",X"01",X"0F",X"D6",X"00",X"0F",X"AC",X"01",X"0F",X"D6",X"00",X"0F",X"57",X"03",X"0F",
		X"AC",X"01",X"0F",X"57",X"03",X"0F",X"AC",X"01",X"0F",X"AC",X"01",X"0F",X"D6",X"00",X"0F",X"AC",
		X"01",X"0F",X"D6",X"00",X"1F",X"57",X"03",X"1F",X"AC",X"01",X"1F",X"57",X"03",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"D6",X"00",X"0F",X"1D",X"01",X"1F",X"D6",X"00",X"0F",X"D6",X"00",X"0F",X"AA",X"00",X"0F",
		X"8F",X"00",X"1F",X"55",X"00",X"0F",X"6B",X"00",X"1F",X"55",X"00",X"0F",X"6B",X"00",X"0F",X"55",
		X"00",X"0F",X"47",X"00",X"40",X"6B",X"00",X"FF",X"07",X"7D",X"01",X"03",X"7D",X"01",X"03",X"7D",
		X"01",X"07",X"1D",X"01",X"07",X"FE",X"00",X"07",X"E2",X"00",X"07",X"FE",X"00",X"07",X"1D",X"01",
		X"07",X"FE",X"00",X"0F",X"E2",X"00",X"0F",X"1D",X"01",X"1F",X"1D",X"01",X"07",X"53",X"01",X"03",
		X"53",X"01",X"03",X"53",X"01",X"07",X"FE",X"00",X"07",X"E2",X"00",X"07",X"D6",X"00",X"07",X"E2",
		X"00",X"07",X"FE",X"00",X"07",X"E2",X"00",X"07",X"D6",X"00",X"07",X"E2",X"00",X"07",X"FE",X"00",
		X"07",X"E2",X"00",X"1F",X"D6",X"00",X"07",X"7D",X"01",X"03",X"7D",X"01",X"03",X"7D",X"01",X"07",
		X"1D",X"01",X"07",X"FE",X"00",X"07",X"E2",X"00",X"07",X"FE",X"00",X"07",X"1D",X"01",X"07",X"FE",
		X"00",X"0F",X"E2",X"00",X"0F",X"BE",X"00",X"1F",X"8F",X"00",X"FF",X"07",X"6B",X"00",X"0F",X"6B",
		X"00",X"0F",X"6B",X"00",X"0F",X"6B",X"00",X"0F",X"6B",X"00",X"0F",X"6B",X"00",X"0F",X"47",X"00",
		X"0F",X"47",X"00",X"0F",X"6B",X"00",X"0F",X"6B",X"00",X"0F",X"6B",X"00",X"0F",X"6B",X"00",X"0F",
		X"6B",X"00",X"0F",X"6B",X"00",X"0F",X"40",X"00",X"0F",X"40",X"00",X"1F",X"47",X"00",X"1F",X"47",
		X"00",X"1F",X"47",X"00",X"FF",X"00",X"9E",X"40",X"9E",X"00",X"9E",X"40",X"8E",X"40",X"8E",X"FF",
		X"07",X"D6",X"00",X"87",X"07",X"D6",X"00",X"87",X"07",X"6B",X"00",X"87",X"07",X"6B",X"00",X"87",
		X"07",X"D6",X"00",X"87",X"07",X"6B",X"00",X"87",X"07",X"6B",X"00",X"87",X"07",X"6B",X"00",X"87",
		X"3A",X"15",X"41",X"FE",X"14",X"C2",X"B8",X"93",X"3A",X"1B",X"41",X"47",X"3A",X"1A",X"41",X"E6",
		X"7F",X"B8",X"30",X"08",X"3A",X"1A",X"41",X"FE",X"83",X"DA",X"12",X"90",X"2F",X"E6",X"7F",X"C6",
		X"28",X"47",X"3A",X"00",X"42",X"E6",X"07",X"20",X"02",X"3E",X"04",X"3D",X"07",X"07",X"07",X"07",
		X"80",X"47",X"3A",X"00",X"41",X"FE",X"4C",X"38",X"08",X"FE",X"75",X"30",X"04",X"0E",X"0F",X"18",
		X"02",X"0E",X"08",X"70",X"3E",X"03",X"12",X"36",X"00",X"3E",X"09",X"12",X"71",X"C3",X"17",X"90",
		X"00",X"00",X"79",X"32",X"75",X"40",X"11",X"20",X"00",X"C9",X"3A",X"75",X"40",X"A7",X"CA",X"12",
		X"90",X"FE",X"22",X"3E",X"40",X"28",X"02",X"3E",X"AC",X"77",X"AF",X"32",X"75",X"40",X"3E",X"03",
		X"12",X"36",X"00",X"0E",X"0F",X"C3",X"49",X"96",X"26",X"50",X"3E",X"06",X"32",X"74",X"40",X"C3",
		X"30",X"3A",X"32",X"5F",X"50",X"18",X"03",X"32",X"5B",X"50",X"3E",X"08",X"32",X"73",X"40",X"C9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"32",X"45",X"50",X"3E",X"80",X"32",X"6D",X"40",X"C9",X"32",X"49",X"50",X"18",X"F5",X"32",X"45",
		X"50",X"3E",X"10",X"32",X"6E",X"40",X"C9",X"FE",X"11",X"30",X"07",X"7D",X"E6",X"E0",X"C6",X"0B",
		X"18",X"05",X"7D",X"E6",X"E0",X"C6",X"1B",X"6F",X"11",X"20",X"00",X"C9",X"36",X"86",X"3E",X"C0",
		X"32",X"6F",X"40",X"C3",X"FE",X"32",X"36",X"87",X"18",X"F4",X"23",X"77",X"23",X"EB",X"C9",X"0E",
		X"FF",X"18",X"02",X"0E",X"01",X"21",X"50",X"50",X"06",X"03",X"7E",X"FE",X"F8",X"30",X"03",X"79",
		X"86",X"77",X"23",X"23",X"23",X"23",X"10",X"F2",X"21",X"3A",X"50",X"C9",X"CD",X"64",X"08",X"3A",
		X"15",X"41",X"FE",X"14",X"C0",X"F1",X"7E",X"D6",X"B8",X"FE",X"04",X"D2",X"A7",X"3B",X"C6",X"20",
		X"C3",X"63",X"3B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"23",X"78",X"C6",X"8C",X"5F",X"16",X"40",X"1A",X"A7",X"28",X"08",X"7E",X"FE",X"17",
		X"38",X"0F",X"35",X"18",X"0E",X"7E",X"FE",X"DF",X"30",X"03",X"34",X"18",X"06",X"3E",X"01",X"18",
		X"01",X"AF",X"12",X"2B",X"2B",X"3A",X"00",X"42",X"C9",X"32",X"70",X"40",X"77",X"2B",X"2B",X"C9",
		X"34",X"26",X"50",X"2B",X"C3",X"D7",X"30",X"32",X"03",X"40",X"32",X"47",X"40",X"32",X"48",X"40",
		X"C9",X"32",X"54",X"50",X"3E",X"F0",X"32",X"71",X"40",X"C9",X"CD",X"0B",X"36",X"C3",X"60",X"0D",
		X"00",X"00",X"01",X"E4",X"04",X"3E",X"08",X"32",X"73",X"40",X"C9",X"2B",X"3E",X"04",X"32",X"74",
		X"40",X"C3",X"63",X"17",X"36",X"02",X"2B",X"3E",X"02",X"32",X"74",X"40",X"7E",X"FE",X"06",X"D0",
		X"36",X"06",X"C9",X"2A",X"91",X"40",X"7C",X"A7",X"20",X"3A",X"2A",X"00",X"41",X"54",X"5D",X"C3",
		X"80",X"A7",X"ED",X"42",X"28",X"1C",X"62",X"6B",X"01",X"01",X"05",X"ED",X"42",X"28",X"13",X"62",
		X"6B",X"01",X"BE",X"05",X"ED",X"42",X"28",X"0A",X"62",X"6B",X"01",X"62",X"07",X"ED",X"42",X"C2",
		X"30",X"9C",X"C3",X"D8",X"99",X"22",X"91",X"40",X"21",X"9C",X"0F",X"22",X"93",X"40",X"3E",X"06",
		X"DD",X"77",X"02",X"C9",X"2A",X"00",X"41",X"01",X"F8",X"07",X"ED",X"42",X"CA",X"53",X"99",X"2A",
		X"91",X"40",X"2D",X"7D",X"FE",X"03",X"DA",X"5D",X"99",X"EB",X"3A",X"93",X"40",X"6F",X"26",X"01",
		X"4E",X"21",X"94",X"40",X"7E",X"FE",X"F0",X"28",X"05",X"36",X"F0",X"A1",X"18",X"14",X"36",X"0F",
		X"A1",X"0F",X"0F",X"0F",X"0F",X"47",X"3A",X"93",X"40",X"FE",X"9E",X"28",X"04",X"3C",X"32",X"93",
		X"40",X"78",X"EB",X"94",X"2F",X"CD",X"91",X"9C",X"2D",X"E5",X"3A",X"92",X"40",X"BC",X"30",X"54",
		X"11",X"F8",X"10",X"19",X"CD",X"64",X"08",X"11",X"20",X"00",X"7E",X"FE",X"C1",X"28",X"13",X"FE",
		X"80",X"38",X"41",X"FE",X"83",X"30",X"3D",X"2B",X"7E",X"23",X"D6",X"8B",X"30",X"04",X"C6",X"0B",
		X"38",X"32",X"C3",X"8E",X"99",X"CD",X"3C",X"0E",X"1E",X"20",X"0E",X"08",X"19",X"0D",X"28",X"1C",
		X"7E",X"D6",X"A6",X"38",X"F7",X"FE",X"12",X"30",X"F3",X"36",X"5E",X"19",X"36",X"5E",X"19",X"36",
		X"21",X"19",X"36",X"23",X"2B",X"36",X"22",X"CD",X"3C",X"0E",X"36",X"20",X"E1",X"7C",X"E6",X"F8",
		X"3D",X"67",X"18",X"0C",X"E1",X"7C",X"FE",X"C7",X"38",X"10",X"FE",X"D8",X"30",X"0C",X"26",X"C7",
		X"3E",X"73",X"32",X"93",X"40",X"3E",X"30",X"32",X"7F",X"40",X"7D",X"DD",X"77",X"00",X"7C",X"FE",
		X"06",X"30",X"02",X"26",X"01",X"DD",X"74",X"03",X"22",X"91",X"40",X"3A",X"00",X"42",X"E6",X"3F",
		X"FE",X"38",X"18",X"06",X"3E",X"17",X"DD",X"77",X"01",X"C9",X"3E",X"24",X"DD",X"77",X"01",X"3A",
		X"40",X"50",X"C6",X"08",X"95",X"FE",X"1C",X"30",X"10",X"3A",X"43",X"50",X"C6",X"0C",X"94",X"FE",
		X"14",X"30",X"06",X"3E",X"01",X"32",X"14",X"40",X"C9",X"EB",X"2A",X"24",X"41",X"7D",X"FE",X"E1",
		X"D0",X"C6",X"0D",X"93",X"FE",X"11",X"D0",X"7C",X"C6",X"0C",X"92",X"FE",X"0F",X"D0",X"3E",X"60",
		X"C3",X"DD",X"1F",X"3E",X"FE",X"DD",X"77",X"00",X"AF",X"32",X"92",X"40",X"C9",X"3E",X"D9",X"DD",
		X"77",X"03",X"3E",X"A4",X"DD",X"77",X"01",X"DD",X"7E",X"00",X"C6",X"04",X"DD",X"77",X"00",X"FE",
		X"F8",X"D2",X"2E",X"9A",X"C9",X"00",X"00",X"00",X"3A",X"97",X"40",X"A7",X"20",X"0B",X"36",X"06",
		X"23",X"36",X"02",X"3E",X"06",X"32",X"97",X"40",X"C9",X"3D",X"36",X"80",X"18",X"F7",X"DD",X"7E",
		X"00",X"FE",X"31",X"DA",X"DC",X"98",X"2B",X"1E",X"A0",X"C3",X"B5",X"98",X"3A",X"20",X"41",X"A7",
		X"C0",X"DD",X"21",X"5C",X"50",X"CD",X"03",X"98",X"3A",X"15",X"41",X"FE",X"0A",X"D8",X"DD",X"21",
		X"58",X"50",X"21",X"91",X"40",X"11",X"99",X"40",X"06",X"04",X"1A",X"4E",X"77",X"79",X"12",X"23",
		X"13",X"10",X"F7",X"CD",X"03",X"98",X"21",X"91",X"40",X"11",X"99",X"40",X"06",X"04",X"1A",X"4E",
		X"77",X"79",X"12",X"23",X"13",X"10",X"F7",X"C9",X"21",X"98",X"40",X"3A",X"00",X"41",X"4F",X"3A",
		X"15",X"41",X"81",X"BE",X"C8",X"77",X"21",X"F1",X"08",X"C3",X"35",X"98",X"01",X"09",X"08",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"20",X"30",X"40",X"60",X"80",X"60",X"40",X"20",X"00",X"21",X"11",X"4A",X"11",X"20",
		X"00",X"3E",X"04",X"A7",X"01",X"EC",X"99",X"F5",X"0A",X"77",X"ED",X"52",X"D9",X"06",X"20",X"CD",
		X"56",X"0D",X"D9",X"03",X"F1",X"3D",X"20",X"EF",X"06",X"F0",X"CD",X"56",X"0D",X"C9",X"7C",X"D6",
		X"30",X"67",X"2E",X"F9",X"22",X"91",X"40",X"C9",X"CD",X"00",X"0E",X"E5",X"C5",X"3A",X"07",X"41",
		X"E6",X"01",X"C6",X"52",X"4F",X"06",X"41",X"0A",X"3C",X"02",X"C5",X"21",X"DF",X"4A",X"0A",X"D6",
		X"19",X"30",X"03",X"0A",X"2D",X"3D",X"0F",X"0F",X"0F",X"0F",X"47",X"E6",X"E0",X"4F",X"78",X"E6",
		X"03",X"CB",X"60",X"28",X"08",X"47",X"A7",X"ED",X"42",X"36",X"1F",X"18",X"06",X"47",X"A7",X"ED",
		X"42",X"36",X"1E",X"C1",X"0A",X"FE",X"30",X"30",X"03",X"C1",X"E1",X"C9",X"00",X"AF",X"02",X"D5",
		X"3E",X"38",X"32",X"A3",X"40",X"3A",X"07",X"41",X"57",X"E6",X"01",X"3C",X"07",X"5F",X"A2",X"20",
		X"1D",X"7B",X"B2",X"32",X"07",X"41",X"79",X"D6",X"39",X"6F",X"26",X"42",X"34",X"CD",X"08",X"36",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D1",X"C1",X"E1",X"C9",X"21",X"7F",
		X"49",X"06",X"0C",X"36",X"1D",X"11",X"20",X"00",X"19",X"78",X"00",X"00",X"00",X"00",X"00",X"E5",
		X"C5",X"0E",X"0A",X"CD",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C1",X"E1",
		X"10",X"E1",X"CB",X"45",X"28",X"05",X"21",X"7E",X"49",X"18",X"D6",X"00",X"00",X"00",X"00",X"00",
		X"18",X"C3",X"0E",X"02",X"06",X"E0",X"C5",X"CD",X"80",X"35",X"06",X"01",X"CD",X"56",X"0D",X"C1",
		X"10",X"F4",X"0D",X"20",X"EF",X"3A",X"07",X"41",X"47",X"E6",X"01",X"6F",X"3C",X"07",X"B0",X"C8",
		X"3E",X"52",X"85",X"6F",X"26",X"41",X"36",X"00",X"21",X"7F",X"49",X"11",X"20",X"00",X"06",X"0C",
		X"7E",X"FE",X"1D",X"20",X"0B",X"19",X"10",X"F7",X"CB",X"45",X"C8",X"21",X"7E",X"49",X"18",X"ED",
		X"E5",X"C5",X"D5",X"C3",X"B3",X"9A",X"7C",X"92",X"FE",X"1B",X"D0",X"08",X"7D",X"93",X"FE",X"1E",
		X"D0",X"D9",X"47",X"3A",X"3A",X"50",X"0F",X"0F",X"0F",X"E6",X"1F",X"90",X"C6",X"1E",X"0F",X"0F",
		X"0F",X"47",X"E6",X"E0",X"4F",X"78",X"E6",X"07",X"47",X"08",X"2F",X"C6",X"1E",X"6F",X"26",X"48",
		X"09",X"D9",X"78",X"D9",X"77",X"D9",X"C9",X"21",X"06",X"48",X"01",X"02",X"20",X"CD",X"45",X"0D",
		X"21",X"24",X"4B",X"01",X"0A",X"50",X"CD",X"CB",X"0A",X"11",X"75",X"15",X"01",X"1F",X"00",X"1A",
		X"FE",X"FF",X"28",X"06",X"77",X"ED",X"42",X"13",X"18",X"F5",X"3E",X"17",X"32",X"49",X"50",X"06",
		X"0A",X"C5",X"06",X"10",X"CD",X"56",X"0D",X"3E",X"0A",X"CD",X"34",X"0E",X"CD",X"37",X"0A",X"C1",
		X"10",X"EF",X"3E",X"01",X"32",X"50",X"40",X"3E",X"73",X"C3",X"83",X"93",X"00",X"3A",X"20",X"41",
		X"A7",X"C8",X"FE",X"05",X"D0",X"21",X"58",X"50",X"7E",X"FE",X"F8",X"30",X"44",X"D6",X"02",X"77",
		X"3A",X"40",X"50",X"C6",X"26",X"BE",X"30",X"5B",X"06",X"00",X"7E",X"FE",X"A9",X"30",X"06",X"FE",
		X"59",X"38",X"02",X"06",X"01",X"2E",X"5B",X"78",X"86",X"77",X"2E",X"5C",X"7E",X"FE",X"F8",X"D0",
		X"3A",X"00",X"42",X"47",X"0F",X"30",X"01",X"35",X"2E",X"5F",X"7E",X"FE",X"54",X"38",X"06",X"78",
		X"35",X"E6",X"18",X"28",X"03",X"34",X"34",X"34",X"7E",X"FE",X"CF",X"D8",X"2E",X"5C",X"36",X"FF",
		X"C9",X"3A",X"20",X"41",X"3D",X"FE",X"03",X"30",X"D1",X"3A",X"00",X"42",X"A7",X"20",X"CB",X"3E",
		X"60",X"32",X"6A",X"40",X"00",X"00",X"21",X"F1",X"04",X"22",X"58",X"50",X"21",X"02",X"27",X"22",
		X"5A",X"50",X"C9",X"3A",X"5C",X"50",X"FE",X"F8",X"38",X"9E",X"7E",X"32",X"5C",X"50",X"3A",X"5B",
		X"50",X"32",X"5F",X"50",X"21",X"05",X"01",X"22",X"5D",X"50",X"3E",X"30",X"32",X"6C",X"40",X"C9",
		X"3A",X"A1",X"40",X"A7",X"C8",X"3D",X"28",X"1B",X"32",X"A1",X"40",X"E6",X"07",X"20",X"05",X"3E",
		X"06",X"32",X"72",X"40",X"DD",X"36",X"01",X"3E",X"DD",X"7E",X"00",X"FE",X"F8",X"D0",X"3D",X"DD",
		X"77",X"00",X"C9",X"DD",X"36",X"00",X"FF",X"C9",X"32",X"01",X"60",X"3E",X"07",X"32",X"00",X"59",
		X"3E",X"3F",X"32",X"00",X"58",X"C9",X"3A",X"07",X"41",X"E6",X"01",X"C6",X"50",X"6F",X"26",X"41",
		X"7E",X"FE",X"02",X"D2",X"D0",X"37",X"3A",X"00",X"42",X"C3",X"CE",X"37",X"3A",X"07",X"41",X"E6",
		X"01",X"C6",X"50",X"4F",X"06",X"41",X"0A",X"A7",X"CA",X"21",X"98",X"01",X"08",X"07",X"C3",X"12",
		X"98",X"C6",X"05",X"67",X"3A",X"07",X"41",X"E6",X"01",X"C6",X"50",X"4F",X"06",X"41",X"0A",X"FE",
		X"01",X"D8",X"3A",X"93",X"40",X"24",X"FE",X"85",X"D0",X"25",X"25",X"C9",X"36",X"F7",X"2B",X"36",
		X"F6",X"C3",X"B0",X"13",X"32",X"5C",X"50",X"32",X"43",X"40",X"32",X"6A",X"40",X"3E",X"08",X"32",
		X"1B",X"42",X"C9",X"CD",X"BE",X"1F",X"C3",X"00",X"83",X"CD",X"BE",X"1F",X"21",X"62",X"40",X"C9",
		X"CD",X"1B",X"0A",X"3A",X"07",X"41",X"E6",X"08",X"CA",X"03",X"93",X"C3",X"2A",X"93",X"22",X"55",
		X"50",X"3E",X"04",X"32",X"59",X"50",X"C9",X"00",X"00",X"00",X"CD",X"30",X"84",X"AF",X"32",X"0C",
		X"41",X"C9",X"3A",X"15",X"41",X"D6",X"0D",X"FE",X"07",X"30",X"04",X"3E",X"07",X"18",X"02",X"3E",
		X"04",X"32",X"42",X"50",X"32",X"46",X"50",X"C3",X"CF",X"12",X"3A",X"20",X"41",X"A7",X"28",X"E2",
		X"18",X"ED",X"CD",X"24",X"1F",X"C3",X"DA",X"83",X"3E",X"FF",X"32",X"4C",X"50",X"C3",X"58",X"87",
		X"2B",X"2B",X"11",X"20",X"00",X"19",X"7E",X"FE",X"E0",X"CA",X"A9",X"8C",X"23",X"23",X"7E",X"FE",
		X"E0",X"CA",X"C9",X"8C",X"F1",X"E1",X"CB",X"5F",X"C3",X"5B",X"8C",X"BF",X"4B",X"68",X"67",X"65",
		X"6E",X"6B",X"6A",X"1C",X"FF",X"BE",X"4B",X"1B",X"67",X"6E",X"1A",X"6A",X"FF",X"BF",X"4B",X"5E",
		X"5E",X"5E",X"5E",X"0B",X"0A",X"1C",X"FF",X"BE",X"4B",X"5E",X"5E",X"5E",X"5E",X"5E",X"FF",X"00",
		X"A3",X"4A",X"88",X"8D",X"92",X"93",X"91",X"94",X"82",X"93",X"88",X"8E",X"8D",X"92",X"FF",X"A4",
		X"4B",X"9B",X"FF",X"A5",X"4B",X"88",X"8D",X"92",X"84",X"91",X"93",X"5E",X"82",X"8E",X"88",X"8D",
		X"92",X"5E",X"80",X"8D",X"83",X"5E",X"8F",X"91",X"84",X"92",X"92",X"5E",X"92",X"93",X"80",X"91",
		X"93",X"FF",X"A6",X"4B",X"9B",X"FF",X"A7",X"4B",X"82",X"8E",X"8D",X"93",X"91",X"8E",X"8B",X"5E",
		X"82",X"80",X"91",X"5E",X"81",X"98",X"5E",X"91",X"87",X"98",X"93",X"87",X"8C",X"88",X"82",X"80",
		X"8B",X"8B",X"98",X"FF",X"A8",X"4B",X"81",X"8E",X"94",X"8D",X"82",X"88",X"8D",X"86",X"5E",X"88",
		X"93",X"5E",X"96",X"88",X"93",X"87",X"5E",X"89",X"8E",X"98",X"5E",X"92",X"93",X"88",X"82",X"8A",
		X"9D",X"FF",X"A9",X"4B",X"9B",X"FF",X"AA",X"4B",X"92",X"82",X"8E",X"91",X"84",X"5E",X"8F",X"8E",
		X"88",X"8D",X"93",X"92",X"5E",X"80",X"8D",X"83",X"5E",X"91",X"84",X"96",X"80",X"91",X"83",X"92",
		X"5E",X"81",X"98",X"FF",X"4B",X"4A",X"7E",X"7C",X"FF",X"AC",X"4B",X"89",X"94",X"8C",X"8F",X"88",
		X"8D",X"86",X"5E",X"8E",X"8D",X"5E",X"7F",X"7D",X"5E",X"8C",X"8E",X"8D",X"84",X"98",X"5E",X"81",
		X"80",X"86",X"9C",X"FF",X"AD",X"4B",X"F6",X"F4",X"FF",X"AE",X"4B",X"F7",X"F5",X"5E",X"83",X"88",
		X"80",X"8C",X"8E",X"8D",X"83",X"9C",X"8E",X"91",X"5E",X"A3",X"A2",X"A1",X"5E",X"82",X"8B",X"8E",
		X"94",X"83",X"9D",X"FF",X"AF",X"4B",X"9B",X"FF",X"B0",X"4B",X"92",X"82",X"8E",X"91",X"84",X"5E",
		X"8F",X"8E",X"88",X"8D",X"93",X"92",X"5E",X"81",X"98",X"5E",X"92",X"87",X"8E",X"8E",X"93",X"88",
		X"8D",X"86",X"FF",X"B1",X"4B",X"84",X"8D",X"84",X"8C",X"88",X"84",X"92",X"5E",X"9F",X"84",X"97",
		X"93",X"91",X"80",X"5E",X"8F",X"8E",X"88",X"8D",X"93",X"92",X"5E",X"85",X"8E",X"91",X"FF",X"92",
		X"4A",X"A6",X"A4",X"FF",X"B3",X"4B",X"92",X"87",X"8E",X"8E",X"93",X"88",X"8D",X"86",X"5E",X"A7",
		X"A5",X"5E",X"89",X"8E",X"8A",X"84",X"91",X"A0",X"5E",X"FF",X"B4",X"4B",X"9B",X"FF",X"B5",X"4B",
		X"80",X"95",X"8E",X"88",X"83",X"5E",X"8B",X"8E",X"92",X"92",X"5E",X"8E",X"85",X"5E",X"82",X"80",
		X"91",X"5E",X"81",X"98",X"5E",X"84",X"95",X"80",X"83",X"88",X"8D",X"86",X"FF",X"B6",X"4B",X"84",
		X"8D",X"84",X"8C",X"88",X"84",X"92",X"9C",X"8C",X"88",X"92",X"92",X"88",X"8B",X"84",X"92",X"5E",
		X"80",X"8D",X"83",X"FF",X"B7",X"4B",X"84",X"91",X"94",X"8F",X"93",X"88",X"8D",X"86",X"5E",X"95",
		X"8E",X"8B",X"82",X"80",X"8D",X"8E",X"92",X"9D",X"FF",X"B8",X"4B",X"9B",X"FF",X"B9",X"4B",X"86",
		X"80",X"88",X"8D",X"5E",X"8E",X"8D",X"84",X"5E",X"84",X"97",X"93",X"91",X"80",X"5E",X"82",X"80",
		X"91",X"5E",X"85",X"8E",X"91",X"5E",X"04",X"08",X"FF",X"BA",X"4B",X"91",X"84",X"96",X"80",X"91",
		X"83",X"92",X"9E",X"9E",X"93",X"87",X"84",X"8D",X"9C",X"92",X"82",X"8E",X"91",X"84",X"5E",X"81",
		X"8E",X"8D",X"94",X"92",X"FF",X"BB",X"4B",X"8F",X"8E",X"88",X"8D",X"93",X"92",X"5E",X"85",X"8E",
		X"91",X"5E",X"84",X"97",X"93",X"91",X"80",X"5E",X"91",X"84",X"96",X"80",X"91",X"83",X"92",X"9D",
		X"FF",X"2A",X"3C",X"42",X"EB",X"2A",X"3A",X"42",X"19",X"7C",X"85",X"FE",X"9E",X"18",X"03",X"22",
		X"55",X"41",X"EB",X"2A",X"63",X"26",X"19",X"EB",X"2A",X"50",X"26",X"EB",X"2A",X"16",X"8A",X"7C",
		X"85",X"FE",X"8B",X"C3",X"66",X"0B",X"C3",X"10",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CD",X"60",X"91",X"3E",X"0A",X"12",X"36",X"00",X"C9",
		X"3E",X"07",X"32",X"00",X"59",X"3E",X"38",X"32",X"00",X"58",X"3E",X"A0",X"32",X"A2",X"40",X"C9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"3A",X"9D",X"40",X"FE",X"FE",X"D2",X"CC",X"1D",X"3A",X"00",X"42",X"0F",X"D2",X"CC",
		X"1D",X"C9",X"34",X"C3",X"76",X"12",X"77",X"77",X"76",X"76",X"66",X"66",X"65",X"65",X"65",X"55",
		X"55",X"55",X"45",X"55",X"54",X"45",X"45",X"55",X"54",X"54",X"54",X"44",X"45",X"45",X"44",X"44",
		X"44",X"44",X"34",X"44",X"44",X"43",X"44",X"43",X"34",X"44",X"43",X"43",X"43",X"43",X"43",X"43",
		X"33",X"34",X"33",X"34",X"33",X"33",X"32",X"33",X"32",X"23",X"33",X"32",X"32",X"23",X"33",X"32",
		X"6B",X"6B",X"50",X"50",X"40",X"40",X"3C",X"40",X"40",X"40",X"6B",X"6B",X"6B",X"6B",X"78",X"78",
		X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"3A",X"A2",X"40",X"A7",X"CA",X"88",X"A0",X"3D",
		X"32",X"A2",X"40",X"C3",X"D0",X"26",X"4F",X"06",X"A0",X"AF",X"21",X"00",X"58",X"11",X"00",X"59",
		X"12",X"0A",X"77",X"3E",X"01",X"12",X"36",X"00",X"3E",X"08",X"12",X"36",X"0F",X"F1",X"C9",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"03",X"38",X"06",X"3A",X"43",X"40",X"C3",X"8B",X"3E",
		X"3A",X"00",X"42",X"0F",X"38",X"F4",X"C3",X"56",X"3F",X"47",X"3A",X"00",X"68",X"E6",X"40",X"20",
		X"01",X"04",X"78",X"C9",X"00",X"CD",X"59",X"A0",X"32",X"5C",X"50",X"C9",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"FF",X"80",X"FF",X"00",X"00",X"80",X"FF",X"00",X"00",X"80",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"80",X"FF",X"80",X"3A",X"A3",X"40",X"A7",X"CA",X"A0",X"91",X"3D",
		X"32",X"A3",X"40",X"0F",X"E6",X"7F",X"C6",X"6C",X"C3",X"26",X"A0",X"3A",X"50",X"40",X"A7",X"C8",
		X"3A",X"76",X"40",X"A7",X"C0",X"C3",X"4A",X"93",X"10",X"4B",X"91",X"80",X"8D",X"8A",X"5E",X"5E",
		X"92",X"82",X"8E",X"91",X"84",X"5E",X"5E",X"5E",X"8D",X"80",X"8C",X"84",X"FF",X"F2",X"4A",X"01",
		X"92",X"93",X"FF",X"F4",X"4A",X"02",X"8D",X"83",X"FF",X"F6",X"4A",X"03",X"91",X"83",X"FF",X"59",
		X"4A",X"93",X"88",X"8C",X"84",X"FF",X"CD",X"44",X"84",X"21",X"07",X"42",X"18",X"06",X"CD",X"44",
		X"84",X"21",X"13",X"42",X"E5",X"11",X"0D",X"42",X"06",X"06",X"1A",X"BE",X"38",X"2C",X"20",X"04",
		X"2B",X"1B",X"10",X"F6",X"E1",X"E5",X"1E",X"27",X"06",X"06",X"1A",X"BE",X"38",X"3D",X"20",X"04",
		X"2B",X"1B",X"10",X"F6",X"E1",X"E5",X"1E",X"2D",X"06",X"06",X"1A",X"BE",X"38",X"44",X"20",X"04",
		X"2B",X"1B",X"10",X"F6",X"E1",X"06",X"F0",X"C3",X"56",X"0D",X"2E",X"22",X"1E",X"28",X"01",X"06",
		X"00",X"ED",X"B0",X"2E",X"08",X"1E",X"22",X"0E",X"06",X"ED",X"B0",X"2E",X"33",X"1E",X"36",X"0E",
		X"06",X"00",X"00",X"ED",X"B8",X"1E",X"0D",X"3E",X"2E",X"18",X"1B",X"2E",X"22",X"1E",X"28",X"01",
		X"06",X"00",X"ED",X"B0",X"2E",X"31",X"1E",X"34",X"0E",X"03",X"ED",X"B0",X"1E",X"27",X"3E",X"31",
		X"18",X"04",X"1E",X"2D",X"3E",X"34",X"E1",X"01",X"06",X"00",X"ED",X"B8",X"6F",X"CD",X"C9",X"A6",
		X"36",X"5E",X"23",X"36",X"80",X"E5",X"3E",X"04",X"32",X"B9",X"49",X"AF",X"CD",X"F4",X"A7",X"3A",
		X"00",X"42",X"E6",X"0C",X"28",X"05",X"CD",X"2E",X"A2",X"18",X"0D",X"E1",X"7E",X"E5",X"F5",X"36",
		X"5E",X"CD",X"2E",X"A2",X"F1",X"E1",X"77",X"E5",X"21",X"CF",X"A0",X"CD",X"1B",X"0A",X"21",X"A4",
		X"40",X"34",X"7E",X"FE",X"3D",X"20",X"1D",X"36",X"00",X"21",X"99",X"49",X"7E",X"A7",X"20",X"13",
		X"3A",X"B9",X"49",X"A7",X"20",X"09",X"E1",X"CD",X"2E",X"A2",X"06",X"F0",X"C3",X"56",X"0D",X"36",
		X"09",X"2E",X"B9",X"35",X"CD",X"51",X"2C",X"E6",X"01",X"3C",X"47",X"3A",X"00",X"40",X"A0",X"20",
		X"1A",X"21",X"00",X"60",X"CB",X"48",X"28",X"02",X"26",X"68",X"7E",X"21",X"A5",X"40",X"E6",X"0C",
		X"20",X"21",X"36",X"3C",X"06",X"01",X"CD",X"56",X"0D",X"18",X"94",X"AF",X"32",X"00",X"40",X"E1",
		X"7D",X"FE",X"2E",X"28",X"C2",X"FE",X"31",X"28",X"BE",X"FE",X"34",X"28",X"BA",X"2B",X"36",X"80",
		X"E5",X"18",X"E1",X"47",X"7E",X"FE",X"3B",X"38",X"20",X"3E",X"28",X"28",X"01",X"AF",X"77",X"E1",
		X"E5",X"CB",X"50",X"20",X"0A",X"35",X"7E",X"FE",X"80",X"30",X"C9",X"36",X"99",X"18",X"C5",X"34",
		X"7E",X"FE",X"9A",X"38",X"BF",X"36",X"80",X"18",X"BB",X"34",X"18",X"B8",X"06",X"06",X"18",X"02",
		X"06",X"03",X"1A",X"77",X"13",X"C5",X"01",X"20",X"00",X"09",X"C1",X"10",X"F5",X"C9",X"21",X"21",
		X"50",X"06",X"07",X"36",X"01",X"23",X"23",X"10",X"FA",X"21",X"A8",X"A0",X"3E",X"04",X"CD",X"1D",
		X"0A",X"11",X"08",X"42",X"21",X"B2",X"49",X"CD",X"1C",X"A2",X"1E",X"22",X"21",X"B4",X"49",X"CD",
		X"1C",X"A2",X"1E",X"28",X"21",X"B6",X"49",X"CD",X"1C",X"A2",X"21",X"12",X"49",X"CD",X"20",X"A2",
		X"2E",X"14",X"CD",X"20",X"A2",X"2E",X"16",X"CD",X"20",X"A2",X"C9",X"AF",X"32",X"43",X"40",X"32",
		X"45",X"40",X"C9",X"03",X"03",X"04",X"07",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",
		X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"07",X"04",X"03",X"03",X"03",X"03",X"00",X"00",X"83",
		X"4A",X"6A",X"5E",X"61",X"5E",X"63",X"5E",X"6E",X"5E",X"63",X"5E",X"6A",X"FF",X"A5",X"4B",X"01",
		X"61",X"65",X"6B",X"6C",X"5E",X"5E",X"5E",X"5E",X"02",X"68",X"66",X"60",X"65",X"6E",X"5E",X"5E",
		X"5E",X"03",X"80",X"67",X"66",X"61",X"60",X"6E",X"67",X"6A",X"FF",X"66",X"4B",X"87",X"5E",X"5E",
		X"5E",X"5E",X"87",X"5E",X"5E",X"5E",X"87",X"5E",X"85",X"5E",X"5E",X"5E",X"5E",X"5E",X"5E",X"5E",
		X"87",X"FF",X"47",X"4B",X"1F",X"5E",X"0B",X"0A",X"5E",X"5E",X"5E",X"5E",X"5E",X"5E",X"87",X"5E",
		X"5E",X"85",X"5E",X"5E",X"0B",X"0A",X"5E",X"5E",X"91",X"FF",X"88",X"4B",X"1F",X"5E",X"82",X"5E",
		X"5E",X"1F",X"82",X"5E",X"5E",X"87",X"5E",X"0B",X"0A",X"85",X"5E",X"87",X"5E",X"5E",X"5E",X"5E",
		X"5E",X"5E",X"90",X"8A",X"8B",X"FF",X"89",X"4B",X"82",X"85",X"82",X"83",X"85",X"83",X"82",X"5E",
		X"5E",X"5E",X"5E",X"5E",X"5E",X"87",X"5E",X"5E",X"5E",X"5E",X"5E",X"85",X"5E",X"8D",X"8E",X"8F",
		X"8F",X"FF",X"8A",X"4B",X"82",X"84",X"82",X"83",X"84",X"83",X"82",X"5E",X"5E",X"5E",X"89",X"5E",
		X"1F",X"85",X"85",X"5E",X"5E",X"5E",X"8A",X"8B",X"1F",X"8C",X"8F",X"8F",X"8F",X"FF",X"8B",X"4B",
		X"86",X"86",X"86",X"86",X"86",X"86",X"86",X"5E",X"5E",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"5E",X"5E",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"FF",X"AD",X"4B",X"04",X"5E",X"65",X"6E",
		X"5E",X"60",X"5E",X"5E",X"5E",X"5E",X"95",X"96",X"97",X"5E",X"5E",X"5E",X"5E",X"5E",X"5E",X"05",
		X"80",X"67",X"66",X"61",X"60",X"6E",X"67",X"6A",X"FF",X"8E",X"4B",X"68",X"6C",X"69",X"60",X"81",
		X"65",X"62",X"9B",X"9A",X"0B",X"0A",X"A1",X"9E",X"5E",X"5E",X"5E",X"5E",X"5E",X"5E",X"5E",X"5E",
		X"87",X"5E",X"0B",X"0A",X"FF",X"CF",X"4A",X"9C",X"AB",X"A1",X"A2",X"94",X"A5",X"A1",X"9E",X"5E",
		X"5E",X"5E",X"5E",X"5E",X"5E",X"91",X"5E",X"5E",X"5E",X"1F",X"FF",X"F0",X"4A",X"9B",X"9D",X"A1",
		X"A8",X"AA",X"92",X"A6",X"A2",X"A1",X"A3",X"5E",X"5E",X"5E",X"5E",X"5E",X"90",X"5E",X"5E",X"8D",
		X"8E",X"8B",X"FF",X"D1",X"4A",X"AB",X"9F",X"A0",X"A9",X"92",X"A7",X"A1",X"A2",X"A4",X"9E",X"5E",
		X"5E",X"5E",X"8D",X"8E",X"8B",X"85",X"8C",X"8F",X"8F",X"FF",X"F2",X"4A",X"98",X"9F",X"A0",X"AB",
		X"9F",X"92",X"A0",X"AB",X"A1",X"AB",X"9F",X"98",X"5E",X"5E",X"8C",X"8F",X"8F",X"8E",X"8F",X"8F",
		X"8F",X"FF",X"F3",X"4A",X"98",X"5E",X"5E",X"9F",X"A0",X"92",X"AB",X"9F",X"A2",X"AB",X"A2",X"98",
		X"5E",X"5E",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"FF",X"F4",X"4A",X"98",X"99",X"99",X"99",
		X"99",X"93",X"99",X"99",X"99",X"99",X"99",X"98",X"FF",X"B6",X"4B",X"06",X"6A",X"63",X"60",X"5E",
		X"5E",X"5E",X"5E",X"5E",X"07",X"6A",X"18",X"6C",X"5E",X"5E",X"5E",X"5E",X"5E",X"08",X"6F",X"65",
		X"6E",X"65",X"6A",X"64",X"FF",X"77",X"4B",X"B1",X"5E",X"5E",X"5E",X"B3",X"5E",X"5E",X"5E",X"85",
		X"5E",X"5E",X"5E",X"1F",X"5E",X"5E",X"5E",X"5E",X"5E",X"5E",X"5E",X"87",X"FF",X"98",X"4B",X"B6",
		X"B6",X"0B",X"0A",X"B5",X"B4",X"B6",X"5E",X"5E",X"87",X"0B",X"0A",X"5E",X"87",X"5E",X"1F",X"5E",
		X"5E",X"87",X"5E",X"5E",X"5E",X"5E",X"5E",X"87",X"FF",X"99",X"4B",X"B8",X"B0",X"B8",X"B8",X"B8",
		X"B8",X"B8",X"5E",X"5E",X"5E",X"BA",X"5E",X"B9",X"5E",X"5E",X"87",X"FF",X"9A",X"4B",X"B7",X"B7",
		X"B7",X"B2",X"B7",X"90",X"B7",X"5E",X"5E",X"5E",X"BC",X"5E",X"5E",X"B9",X"5E",X"5E",X"5E",X"5E",
		X"5E",X"5E",X"BB",X"0B",X"0A",X"BB",X"BB",X"FF",X"7B",X"4B",X"1F",X"5E",X"5E",X"AC",X"AE",X"AD",
		X"5E",X"5E",X"B6",X"B6",X"B6",X"B6",X"B6",X"BD",X"B6",X"5E",X"5E",X"B6",X"B6",X"86",X"86",X"86",
		X"86",X"86",X"FF",X"9C",X"4B",X"AF",X"AE",X"AF",X"AF",X"AE",X"AE",X"AE",X"5E",X"5E",X"B8",X"B8",
		X"B8",X"B8",X"B8",X"B8",X"B8",X"5E",X"5E",X"B8",X"B8",X"86",X"86",X"86",X"86",X"86",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"CD",X"00",X"83",X"21",X"01",X"01",X"22",X"02",X"60",X"21",X"07",X"50",
		X"11",X"73",X"A2",X"06",X"1A",X"1A",X"77",X"23",X"23",X"13",X"10",X"F9",X"21",X"8F",X"A2",X"3E",
		X"17",X"CD",X"1D",X"0A",X"0E",X"10",X"06",X"20",X"CD",X"56",X"0D",X"0D",X"20",X"F8",X"C9",X"00",
		X"3E",X"08",X"32",X"07",X"41",X"32",X"04",X"70",X"CD",X"5E",X"A6",X"CD",X"18",X"A5",X"CD",X"D4",
		X"A4",X"CD",X"D2",X"A6",X"C9",X"00",X"00",X"00",X"CD",X"00",X"83",X"CD",X"91",X"82",X"21",X"07",
		X"50",X"06",X"19",X"36",X"04",X"23",X"23",X"10",X"FA",X"2E",X"25",X"36",X"06",X"2E",X"07",X"36",
		X"03",X"21",X"60",X"9D",X"3E",X"19",X"CD",X"1D",X"0A",X"0E",X"20",X"C3",X"F6",X"A4",X"00",X"00",
		X"5E",X"5E",X"5E",X"5E",X"89",X"8A",X"5E",X"5E",X"B9",X"5E",X"5E",X"5E",X"81",X"8B",X"8F",X"5E",
		X"5E",X"80",X"83",X"5E",X"88",X"8C",X"90",X"B8",X"5E",X"81",X"84",X"84",X"86",X"8D",X"91",X"5E",
		X"5E",X"81",X"85",X"84",X"87",X"8E",X"5E",X"5E",X"5E",X"82",X"92",X"8C",X"8B",X"8F",X"5E",X"5E",
		X"BA",X"5E",X"A7",X"88",X"8C",X"90",X"B8",X"5E",X"5E",X"93",X"94",X"95",X"96",X"91",X"5E",X"5E",
		X"5E",X"97",X"8C",X"8C",X"9A",X"5E",X"5E",X"5E",X"B9",X"98",X"8C",X"8C",X"9B",X"5E",X"5E",X"5E",
		X"5E",X"97",X"8C",X"8C",X"9C",X"A0",X"B8",X"5E",X"5E",X"99",X"9D",X"9E",X"9F",X"8E",X"5E",X"5E",
		X"5E",X"5E",X"81",X"A1",X"A5",X"5E",X"5E",X"5E",X"5E",X"5E",X"81",X"A2",X"A5",X"5E",X"5E",X"5E",
		X"5E",X"BA",X"A3",X"8C",X"8E",X"5E",X"5E",X"5E",X"5E",X"5E",X"A7",X"A8",X"A9",X"5E",X"5E",X"5E",
		X"B9",X"89",X"84",X"86",X"8B",X"8A",X"5E",X"5E",X"5E",X"81",X"A1",X"8C",X"A1",X"8B",X"8F",X"5E",
		X"5E",X"81",X"A2",X"8C",X"A2",X"8C",X"90",X"B8",X"5E",X"A3",X"AA",X"AB",X"8C",X"8D",X"91",X"5E",
		X"5E",X"AD",X"A4",X"AC",X"A4",X"8E",X"5E",X"5E",X"5E",X"5E",X"5E",X"88",X"8C",X"90",X"5E",X"5E",
		X"5E",X"AE",X"84",X"86",X"8D",X"91",X"5E",X"5E",X"BA",X"99",X"9D",X"B4",X"B5",X"B6",X"5E",X"5E",
		X"5E",X"AF",X"A6",X"B3",X"B7",X"B1",X"5E",X"5E",X"5E",X"97",X"B2",X"AF",X"87",X"A5",X"B8",X"5E",
		X"5E",X"B0",X"B1",X"97",X"AA",X"A5",X"5E",X"5E",X"BA",X"A7",X"82",X"B0",X"A4",X"8E",X"5E",X"5E",
		X"70",X"4A",X"6A",X"5E",X"63",X"5E",X"6D",X"5E",X"60",X"5E",X"FF",X"52",X"4A",X"BC",X"5E",X"01",
		X"09",X"08",X"01",X"FF",X"14",X"4B",X"60",X"66",X"66",X"5E",X"69",X"65",X"6D",X"64",X"6B",X"6A",
		X"5E",X"69",X"63",X"6A",X"63",X"69",X"BD",X"63",X"62",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"D9",X"21",X"0C",X"50",X"7E",X"06",X"08",X"35",X"23",X"23",X"10",X"FB",X"D9",X"C9",X"3E",X"01",
		X"32",X"01",X"70",X"CD",X"91",X"82",X"3E",X"01",X"32",X"03",X"60",X"CD",X"00",X"83",X"21",X"0D",
		X"50",X"01",X"04",X"0A",X"71",X"23",X"23",X"10",X"FB",X"79",X"FE",X"04",X"20",X"05",X"01",X"07",
		X"05",X"18",X"F1",X"21",X"C6",X"4B",X"11",X"40",X"A5",X"0E",X"1C",X"CD",X"50",X"A6",X"E6",X"07",
		X"28",X"09",X"D9",X"06",X"01",X"CD",X"56",X"0D",X"D9",X"18",X"F0",X"06",X"08",X"1A",X"77",X"23",
		X"13",X"10",X"FA",X"D5",X"11",X"28",X"00",X"A7",X"ED",X"52",X"D1",X"0D",X"20",X"E4",X"11",X"20",
		X"01",X"CD",X"50",X"A6",X"06",X"01",X"CD",X"56",X"0D",X"1B",X"7A",X"B3",X"20",X"F3",X"21",X"20",
		X"A6",X"3E",X"03",X"CD",X"1D",X"0A",X"C3",X"F4",X"A4",X"E5",X"CD",X"37",X"0A",X"E1",X"36",X"5E",
		X"23",X"C9",X"CD",X"00",X"83",X"CD",X"91",X"82",X"CD",X"2E",X"A2",X"0E",X"06",X"C3",X"F6",X"A4",
		X"97",X"97",X"97",X"97",X"97",X"97",X"97",X"97",X"97",X"3E",X"05",X"32",X"0B",X"42",X"32",X"25",
		X"42",X"32",X"2B",X"42",X"21",X"E0",X"A6",X"11",X"2E",X"42",X"01",X"09",X"00",X"ED",X"B0",X"C3",
		X"D7",X"A7",X"21",X"17",X"42",X"3A",X"00",X"60",X"0F",X"30",X"0C",X"7E",X"A7",X"C8",X"36",X"00",
		X"2E",X"1D",X"7E",X"A7",X"C2",X"1D",X"82",X"36",X"01",X"C9",X"3A",X"00",X"70",X"E6",X"0C",X"20",
		X"0D",X"CD",X"10",X"82",X"2E",X"1C",X"3A",X"00",X"68",X"E6",X"20",X"C3",X"18",X"82",X"D6",X"08",
		X"38",X"33",X"28",X"1C",X"CD",X"10",X"82",X"2E",X"1C",X"3A",X"00",X"68",X"E6",X"20",X"28",X"0D",
		X"7E",X"A7",X"C8",X"36",X"00",X"06",X"06",X"CD",X"1F",X"82",X"10",X"FB",X"C9",X"36",X"01",X"C9",
		X"CD",X"02",X"A7",X"2E",X"1C",X"3A",X"00",X"68",X"E6",X"20",X"28",X"F1",X"7E",X"A7",X"C8",X"36",
		X"00",X"06",X"03",X"18",X"E2",X"CD",X"02",X"A7",X"2E",X"1C",X"3A",X"00",X"68",X"E6",X"20",X"28",
		X"0C",X"7E",X"A7",X"C8",X"36",X"00",X"2E",X"1D",X"7E",X"A7",X"C2",X"1D",X"82",X"36",X"01",X"C9",
		X"3A",X"00",X"68",X"E6",X"40",X"CA",X"7C",X"9C",X"C3",X"8B",X"9C",X"3A",X"00",X"68",X"E6",X"40",
		X"CA",X"7C",X"9C",X"C3",X"CC",X"1D",X"47",X"3A",X"00",X"68",X"E6",X"40",X"78",X"CA",X"46",X"A0",
		X"3A",X"43",X"40",X"C3",X"8B",X"3E",X"3A",X"00",X"68",X"E6",X"40",X"20",X"04",X"7E",X"D6",X"03",
		X"C9",X"7E",X"D6",X"05",X"C9",X"3A",X"07",X"41",X"E6",X"08",X"C2",X"BD",X"3A",X"CD",X"51",X"2C",
		X"C3",X"B4",X"3A",X"21",X"00",X"B0",X"06",X"03",X"36",X"AA",X"10",X"FC",X"2E",X"04",X"06",X"03",
		X"36",X"55",X"10",X"FC",X"C3",X"00",X"08",X"21",X"00",X"00",X"01",X"FF",X"3F",X"CD",X"72",X"8D",
		X"EB",X"22",X"3A",X"42",X"21",X"00",X"80",X"01",X"00",X"9F",X"CD",X"72",X"8D",X"EB",X"22",X"3C",
		X"42",X"C3",X"42",X"82",X"32",X"99",X"49",X"32",X"00",X"40",X"C9",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
