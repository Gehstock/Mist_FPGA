library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity skyskip_sp_bits_4 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of skyskip_sp_bits_4 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",
		X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",X"00",
		X"08",X"08",X"14",X"32",X"F0",X"68",X"24",X"40",X"10",X"10",X"10",X"10",X"08",X"08",X"08",X"04",
		X"F1",X"FF",X"FF",X"FE",X"FF",X"FF",X"3F",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"3F",X"1F",X"1F",X"DF",X"1F",X"1F",X"3F",X"FF",X"3F",X"9F",X"5F",X"4F",
		X"2F",X"2F",X"0F",X"07",X"03",X"80",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"06",X"0C",X"FC",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FB",X"FF",X"EF",X"1F",X"BF",X"FF",X"FF",X"FC",X"03",X"FF",X"FF",X"7F",X"7F",X"7F",X"3F",X"3F",
		X"01",X"88",X"04",X"02",X"01",X"00",X"80",X"41",X"41",X"E3",X"FF",X"FF",X"3F",X"03",X"00",X"FF",
		X"00",X"03",X"00",X"80",X"C0",X"E0",X"E0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"E0",X"C0",X"80",X"80",X"80",X"C0",X"40",X"00",X"00",X"00",
		X"F0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"80",X"00",X"00",X"80",X"80",X"C0",X"E0",
		X"F0",X"FC",X"FF",X"FF",X"CF",X"BF",X"BF",X"7F",X"7F",X"EF",X"C2",X"99",X"36",X"6E",X"28",X"18",
		X"00",X"40",X"60",X"30",X"00",X"80",X"E0",X"E0",X"C0",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",
		X"00",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"03",X"02",X"00",X"00",X"01",X"03",X"03",X"02",X"05",X"02",X"03",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"80",X"C0",X"E0",X"E0",X"E0",X"F0",X"F8",X"F8",X"F8",X"F8",X"FC",X"FC",X"FC",
		X"7C",X"3C",X"3C",X"1C",X"1E",X"1D",X"0C",X"08",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7C",X"3C",X"3D",X"1F",X"1E",X"1C",X"0E",X"07",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"60",X"F0",X"F0",X"F0",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",
		X"00",X"00",X"0E",X"04",X"00",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"80",X"80",X"00",X"00",X"11",X"0E",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"80",X"80",X"00",X"00",X"11",X"0E",X"20",X"00",X"00",
		X"82",X"03",X"07",X"0F",X"0F",X"6E",X"F6",X"F8",X"FC",X"FC",X"FC",X"FC",X"FC",X"E0",X"00",X"00",
		X"00",X"02",X"03",X"07",X"8F",X"CF",X"E6",X"E0",X"E0",X"E0",X"00",X"00",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"4C",X"84",X"08",X"CC",X"00",X"00",X"00",X"80",X"84",X"00",
		X"00",X"98",X"83",X"41",X"60",X"80",X"00",X"00",X"C3",X"FF",X"FF",X"FF",X"FF",X"FE",X"C0",X"9C",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",X"F2",
		X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"B3",X"C1",X"F8",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"7E",X"3C",X"18",X"00",X"04",X"02",
		X"FE",X"3C",X"CF",X"F1",X"FF",X"FF",X"FB",X"F3",X"F3",X"E3",X"F8",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"7E",X"3C",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"9E",X"EC",X"F5",X"C1",X"C1",X"E3",X"F3",X"FB",X"F9",X"F9",X"F8",X"00",X"A0",X"40",X"A0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"00",X"30",X"78",X"F8",
		X"FC",X"80",X"F0",X"FC",X"FE",X"FE",X"FE",X"FC",X"FE",X"FD",X"FD",X"FF",X"FF",X"FF",X"FB",X"F9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"C0",X"C0",X"E0",X"F0",X"F8",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"F8",X"F8",X"F8",
		X"00",X"00",X"04",X"04",X"04",X"14",X"30",X"30",X"30",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"10",X"00",X"00",X"40",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"90",X"80",X"80",X"40",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"7E",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"FF",X"FF",
		X"EF",X"FE",X"FF",X"FF",X"FB",X"F0",X"E0",X"C0",X"06",X"96",X"16",X"56",X"56",X"50",X"40",X"00",
		X"EF",X"F6",X"F7",X"FF",X"FB",X"F1",X"E1",X"01",X"00",X"80",X"C0",X"C0",X"C0",X"C0",X"60",X"7C",
		X"EF",X"F6",X"F7",X"FF",X"FB",X"F0",X"E0",X"C0",X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"DF",X"8F",X"86",X"86",X"87",X"EF",X"FF",X"FF",
		X"00",X"01",X"04",X"02",X"01",X"05",X"07",X"33",X"4B",X"86",X"86",X"87",X"87",X"CF",X"FF",X"FF",
		X"FE",X"7E",X"3E",X"3E",X"3C",X"78",X"F0",X"E0",X"E8",X"ED",X"8D",X"8D",X"C5",X"E0",X"30",X"98",
		X"7F",X"3F",X"3E",X"3E",X"7C",X"F8",X"F0",X"F0",X"E0",X"C0",X"80",X"80",X"C0",X"E0",X"30",X"98",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"1F",
		X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"77",X"77",X"BB",X"BB",X"B9",X"BC",X"AE",X"A6",
		X"26",X"44",X"0C",X"08",X"19",X"F2",X"F2",X"00",X"01",X"02",X"03",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"3C",X"3C",X"1C",X"18",
		X"00",X"78",X"FC",X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"78",X"78",
		X"78",X"F0",X"F0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"F0",X"FC",X"FE",X"FF",X"FF",X"FF",X"BF",X"3F",X"FF",X"FE",X"F2",X"50",X"08",X"0C",X"0A",X"09",
		X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"C0",X"80",X"00",X"00",X"3C",
		X"04",X"02",X"00",X"00",X"68",X"58",X"D8",X"B8",X"38",X"78",X"F0",X"F0",X"F0",X"30",X"E0",X"E0",
		X"72",X"60",X"30",X"08",X"08",X"40",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"BF",X"1F",X"0F",X"07",X"03",X"01",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"03",
		X"03",X"71",X"D0",X"D8",X"88",X"D8",X"D8",X"D0",X"60",X"00",X"02",X"07",X"07",X"0F",X"0F",X"CF",
		X"83",X"C3",X"31",X"31",X"E3",X"C7",X"47",X"1F",X"FF",X"FC",X"F8",X"F0",X"80",X"40",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"F2",X"FF",X"FF",X"FF",X"FF",X"7F",
		X"FE",X"F7",X"F7",X"E7",X"EF",X"EF",X"FF",X"EC",X"E8",X"E0",X"E0",X"C6",X"8E",X"1E",X"1F",X"3F",
		X"3F",X"FF",X"7F",X"7F",X"7F",X"7F",X"7F",X"7C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"3F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",X"B8",X"30",X"50",X"10",X"80",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"04",X"40",X"10",X"40",X"28",X"00",X"00",X"00",
		X"C0",X"C0",X"C0",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"03",X"01",X"18",X"7C",X"FF",X"FF",X"FF",X"FF",X"FE",X"FD",X"FB",X"E7",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"27",X"67",X"67",X"4F",X"8F",X"0F",X"05",
		X"00",X"00",X"00",X"00",X"00",X"03",X"CF",X"CF",X"CF",X"FF",X"FF",X"FF",X"FF",X"DF",X"8F",X"07",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"F0",X"F0",X"70",X"00",
		X"00",X"1C",X"3E",X"3E",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"38",X"3C",X"3C",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"FC",X"FE",X"FE",X"FC",X"FC",X"FF",X"FE",X"FD",X"FD",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"00",X"71",X"FD",X"BF",X"BF",X"BF",X"DF",X"E0",X"7F",X"01",X"01",X"00",X"00",X"00",X"80",X"C0",
		X"30",X"90",X"D0",X"00",X"80",X"80",X"80",X"0B",X"3C",X"78",X"78",X"78",X"3C",X"9F",X"9F",X"0F",
		X"40",X"C0",X"80",X"80",X"C0",X"60",X"24",X"0C",X"1F",X"3C",X"38",X"38",X"18",X"9C",X"8F",X"0F",
		X"0F",X"1F",X"7F",X"FF",X"F7",X"FC",X"F8",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"1F",X"7F",X"FF",X"FE",X"FC",X"F8",X"E0",X"80",X"00",X"00",X"80",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"7F",X"FF",X"FF",X"FC",X"F8",X"F0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",
		X"E0",X"F0",X"F8",X"FC",X"FE",X"DE",X"3F",X"FF",X"FF",X"FE",X"FC",X"FC",X"F8",X"F8",X"FC",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"E0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F8",
		X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"60",X"80",X"80",X"C0",X"C0",X"E0",X"E0",X"E0",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"E0",X"E0",X"E0",X"C0",X"00",X"00",X"00",
		X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"E0",X"E0",X"C0",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"F8",X"FC",X"FE",X"FC",X"F8",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"00",
		X"FC",X"F8",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"00",
		X"1E",X"BF",X"1F",X"CF",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"E0",
		X"3E",X"FF",X"FF",X"FF",X"FF",X"FF",X"F9",X"F8",X"F1",X"F1",X"E1",X"E3",X"E7",X"E7",X"C7",X"CF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"1F",
		X"7F",X"F1",X"F0",X"E0",X"E0",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F1",X"FF",X"7F",X"1F",X"1F",
		X"FF",X"FF",X"7C",X"BB",X"BB",X"BF",X"BF",X"BD",X"BD",X"BF",X"BF",X"BB",X"BB",X"7C",X"FF",X"FF",
		X"FF",X"FF",X"E0",X"DF",X"BF",X"BF",X"BF",X"B1",X"BF",X"BF",X"BF",X"BF",X"BF",X"CE",X"FF",X"FF",
		X"FF",X"FF",X"E7",X"DB",X"DB",X"DB",X"FB",X"FB",X"DB",X"DB",X"3B",X"FB",X"FB",X"07",X"FF",X"FF",
		X"FF",X"03",X"03",X"F3",X"F3",X"F3",X"FF",X"FF",X"FC",X"F8",X"F0",X"E0",X"C0",X"C0",X"C0",X"C0",
		X"1C",X"3E",X"FE",X"7C",X"7E",X"3E",X"3C",X"1C",X"1C",X"08",X"00",X"0A",X"1B",X"1F",X"3E",X"3C",
		X"78",X"7C",X"FC",X"FE",X"FC",X"F8",X"E8",X"A2",X"A6",X"E6",X"6E",X"6E",X"7C",X"7C",X"38",X"10",
		X"7F",X"3F",X"FF",X"66",X"70",X"30",X"38",X"18",X"18",X"08",X"02",X"0B",X"1B",X"1F",X"3E",X"3C",
		X"78",X"7C",X"FC",X"FE",X"FC",X"F8",X"E8",X"A4",X"A0",X"E0",X"60",X"66",X"7F",X"7F",X"7E",X"38",
		X"00",X"0F",X"1F",X"FF",X"FF",X"FD",X"0D",X"1E",X"A6",X"02",X"02",X"02",X"A6",X"1C",X"0C",X"0C",
		X"1C",X"FC",X"FC",X"7E",X"80",X"FC",X"FE",X"F6",X"F6",X"A6",X"E6",X"CF",X"E7",X"6A",X"62",X"C0",
		X"3F",X"3E",X"38",X"F8",X"FC",X"FC",X"0C",X"1E",X"A6",X"03",X"03",X"03",X"A7",X"1E",X"0C",X"0C",
		X"18",X"F8",X"FC",X"7E",X"80",X"FC",X"F8",X"F0",X"F0",X"A0",X"E0",X"C0",X"60",X"60",X"E0",X"C0",
		X"00",X"10",X"10",X"18",X"BC",X"F6",X"F2",X"F0",X"78",X"38",X"3C",X"1C",X"0C",X"06",X"06",X"06",
		X"06",X"0E",X"0E",X"9F",X"FD",X"FF",X"FB",X"BF",X"BF",X"E6",X"46",X"06",X"04",X"08",X"00",X"00",
		X"3E",X"78",X"60",X"20",X"A0",X"E0",X"F0",X"F0",X"78",X"38",X"3C",X"1C",X"0C",X"06",X"06",X"06",
		X"06",X"0E",X"0E",X"9E",X"FC",X"FC",X"FC",X"F8",X"B8",X"F0",X"40",X"00",X"00",X"00",X"00",X"00",
		X"3C",X"7C",X"FC",X"FC",X"00",X"00",X"20",X"70",X"70",X"50",X"50",X"20",X"00",X"00",X"00",X"00",
		X"7E",X"7E",X"4C",X"00",X"FC",X"FC",X"1C",X"3C",X"78",X"0C",X"04",X"05",X"07",X"07",X"0F",X"1E",
		X"3C",X"00",X"00",X"20",X"70",X"70",X"50",X"50",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"38",X"7C",X"7C",X"48",X"00",X"FC",X"FC",X"1C",X"3C",X"7C",X"0C",X"04",X"06",X"06",X"07",X"0F",
		X"1C",X"38",X"7C",X"FC",X"00",X"00",X"20",X"70",X"70",X"50",X"50",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"E0",X"F0",X"A8",X"0C",X"0E",X"0E",X"1F",X"0E",X"0E",X"04",X"04",X"00",X"00",
		X"00",X"00",X"C0",X"E0",X"F0",X"E8",X"0C",X"0E",X"0E",X"1F",X"0E",X"0E",X"04",X"04",X"00",X"00",
		X"1F",X"38",X"74",X"6C",X"3A",X"14",X"0B",X"00",X"00",X"00",X"04",X"04",X"00",X"00",X"00",X"00",
		X"6C",X"FC",X"0C",X"18",X"04",X"04",X"0E",X"0E",X"0E",X"9F",X"8E",X"0E",X"04",X"04",X"00",X"00",
		X"1F",X"38",X"74",X"6C",X"3A",X"14",X"0B",X"00",X"04",X"04",X"0E",X"0E",X"04",X"00",X"00",X"00",
		X"06",X"00",X"7C",X"FF",X"FF",X"FF",X"C7",X"00",X"00",X"07",X"01",X"03",X"03",X"04",X"03",X"03",
		X"38",X"FE",X"FF",X"FF",X"FF",X"DF",X"18",X"00",X"00",X"07",X"01",X"03",X"03",X"04",X"03",X"03",
		X"C7",X"EF",X"FE",X"FE",X"FF",X"FF",X"FB",X"FD",X"DF",X"8F",X"80",X"80",X"00",X"10",X"01",X"01",
		X"1C",X"0C",X"7F",X"FF",X"FF",X"FF",X"E7",X"00",X"00",X"0F",X"09",X"03",X"03",X"04",X"0B",X"0B",
		X"06",X"00",X"7C",X"FF",X"FF",X"FF",X"C7",X"00",X"00",X"C7",X"C1",X"E3",X"63",X"44",X"0B",X"0B",
		X"CF",X"FF",X"FE",X"FF",X"FF",X"FF",X"7B",X"3D",X"1F",X"0F",X"00",X"00",X"00",X"10",X"01",X"01",
		X"E0",X"E3",X"23",X"21",X"A1",X"E0",X"F0",X"D0",X"90",X"38",X"78",X"E9",X"CB",X"CE",X"84",X"04",
		X"00",X"00",X"03",X"0F",X"1F",X"07",X"03",X"00",X"00",X"80",X"C0",X"C1",X"03",X"06",X"0C",X"08",
		X"00",X"00",X"03",X"0F",X"07",X"01",X"00",X"00",X"80",X"C0",X"C0",X"C1",X"43",X"06",X"0C",X"88",
		X"FF",X"FF",X"E6",X"C0",X"C0",X"E0",X"E0",X"E0",X"7F",X"5E",X"5E",X"77",X"C1",X"62",X"22",X"C1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"C3",X"E6",X"FE",X"FE",X"FC",X"FC",X"F8",X"F0",X"C0",
		X"02",X"03",X"86",X"EC",X"FC",X"FC",X"F8",X"F0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"D8",X"F8",X"F0",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"E4",X"E4",X"3E",X"3E",X"FE",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"00",X"00",X"00",
		X"F8",X"9C",X"9C",X"F2",X"F2",X"FE",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",
		X"F8",X"E4",X"E4",X"3E",X"3E",X"FE",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"02",X"05",X"02",X"00",X"00",
		X"00",X"00",X"E0",X"00",X"F0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"0F",X"00",
		X"AA",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"07",X"00",X"00",X"00",
		X"38",X"00",X"7F",X"00",X"FF",X"00",X"7F",X"00",X"3F",X"00",X"1F",X"00",X"0F",X"00",X"00",X"00",
		X"03",X"00",X"00",X"00",X"60",X"00",X"F8",X"00",X"FF",X"00",X"3F",X"00",X"1C",X"00",X"00",X"00",
		X"50",X"00",X"FC",X"00",X"FE",X"00",X"FF",X"00",X"7F",X"00",X"3F",X"00",X"7F",X"00",X"3F",X"00",
		X"AA",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"EF",X"00",X"F3",X"00",X"FC",X"00",X"FF",X"00",X"FF",X"00",X"1E",X"00",X"00",X"00",
		X"3F",X"00",X"0F",X"00",X"C0",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"1F",X"00",X"0E",X"00",
		X"F8",X"F8",X"7C",X"7C",X"3E",X"3F",X"3F",X"1F",X"1F",X"1F",X"9F",X"9F",X"9F",X"CF",X"CF",X"E7",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"0F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"CF",X"07",X"00",X"00",X"00",X"00",X"00",X"C0",X"F0",X"FF",X"0F",
		X"73",X"7F",X"3F",X"3F",X"1F",X"0F",X"C6",X"00",X"F0",X"00",X"FE",X"00",X"1F",X"00",X"00",X"00",
		X"1F",X"1F",X"1F",X"0F",X"1F",X"1F",X"0F",X"07",X"00",X"00",X"00",X"80",X"F0",X"FC",X"FC",X"EC",
		X"3F",X"3F",X"3F",X"1F",X"1F",X"0F",X"1F",X"1F",X"1F",X"8F",X"C7",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"B7",X"83",X"80",X"C0",X"E0",X"E0",X"F0",X"F9",X"FF",X"7E",X"04",
		X"0C",X"1E",X"1F",X"1F",X"0F",X"0F",X"0F",X"07",X"03",X"01",X"00",X"80",X"00",X"F0",X"00",X"1C",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"07",X"03",X"E1",X"FD",X"FD",X"3D",X"07",
		X"9F",X"CF",X"0F",X"03",X"00",X"00",X"00",X"C0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",
		X"03",X"03",X"01",X"00",X"02",X"03",X"03",X"07",X"0F",X"1F",X"1F",X"3F",X"3F",X"3F",X"1F",X"07",
		X"FC",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"1F",X"03",X"C0",X"F0",X"E0",
		X"FF",X"FF",X"FF",X"3F",X"07",X"01",X"00",X"04",X"04",X"06",X"06",X"07",X"07",X"03",X"03",X"01",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"EF",X"E7",X"F0",X"F8",
		X"3C",X"1F",X"0F",X"07",X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"03",X"01",X"01",X"01",X"00",
		X"FF",X"00",X"40",X"60",X"F0",X"E8",X"8C",X"8E",X"0E",X"1F",X"0E",X"0E",X"04",X"04",X"00",X"00",
		X"FF",X"7C",X"1C",X"18",X"04",X"04",X"0E",X"8E",X"0E",X"1F",X"0E",X"0E",X"04",X"04",X"00",X"00",
		X"1F",X"38",X"74",X"6C",X"3A",X"14",X"0B",X"00",X"00",X"00",X"04",X"04",X"00",X"00",X"00",X"FF",
		X"1F",X"38",X"74",X"6C",X"3A",X"14",X"0B",X"00",X"04",X"04",X"0E",X"0E",X"04",X"00",X"00",X"FF",
		X"00",X"53",X"1E",X"DF",X"DF",X"14",X"00",X"31",X"00",X"07",X"00",X"03",X"03",X"04",X"8B",X"8B",
		X"00",X"FF",X"00",X"43",X"FF",X"FF",X"78",X"00",X"80",X"C7",X"C1",X"E3",X"63",X"47",X"0B",X"0B",
		X"CF",X"FF",X"FE",X"FF",X"FF",X"FF",X"7B",X"3D",X"1F",X"0F",X"00",X"00",X"00",X"10",X"01",X"00",
		X"FF",X"00",X"03",X"0F",X"07",X"01",X"00",X"00",X"80",X"C0",X"C0",X"C1",X"43",X"06",X"0C",X"88",
		X"FF",X"00",X"07",X"1F",X"1F",X"07",X"03",X"00",X"00",X"80",X"C0",X"C1",X"43",X"06",X"0C",X"08",
		X"FF",X"FF",X"E6",X"C0",X"C0",X"E0",X"E0",X"E0",X"7F",X"5F",X"5E",X"77",X"C1",X"E3",X"E3",X"00",
		X"FF",X"FF",X"E6",X"C0",X"C0",X"E0",X"E0",X"E0",X"7F",X"5F",X"5E",X"7F",X"C1",X"E3",X"E3",X"00",
		X"3F",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"3F",X"9F",X"FF",X"F8",X"FC",X"3F",X"0F",X"07",X"07",
		X"07",X"03",X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"9F",X"87",X"83",X"C3",X"03",X"01",X"01",X"01",
		X"C0",X"F0",X"F8",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"F8",X"F0",X"C0",
		X"C0",X"F0",X"F8",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"F8",X"F0",X"C0",
		X"00",X"0E",X"0E",X"0E",X"30",X"30",X"40",X"00",X"00",X"40",X"30",X"30",X"0E",X"0E",X"0E",X"00",
		X"01",X"B0",X"F4",X"E8",X"F4",X"F8",X"F8",X"FE",X"FE",X"FC",X"E8",X"72",X"F2",X"E4",X"E8",X"80",
		X"FF",X"EF",X"BF",X"7F",X"FF",X"FF",X"FD",X"7F",X"3D",X"1D",X"0D",X"00",X"00",X"0C",X"02",X"00",
		X"2F",X"7F",X"7F",X"3F",X"5F",X"1B",X"87",X"41",X"00",X"02",X"01",X"00",X"00",X"20",X"00",X"40",
		X"00",X"20",X"C0",X"0F",X"1F",X"1F",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"10",X"00",X"08",X"0F",X"1F",X"1F",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"88",X"88",X"08",X"08",X"0E",X"0F",X"07",X"07",X"76",X"F6",X"F2",X"FA",X"02",X"02",X"02",X"00",
		X"00",X"00",X"00",X"01",X"01",X"1D",X"3F",X"3F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"7F",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"80",X"C0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"80",X"00",X"00",X"00",X"80",X"C0",X"E0",
		X"F0",X"F0",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"1D",X"3C",X"39",X"38",X"3C",X"7C",X"3E",X"1F",X"1F",X"3E",X"3E",X"5E",X"CF",X"D7",X"12",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"F0",X"FA",X"F9",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"F1",X"F8",X"F8",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"04",X"12",X"09",X"07",X"03",X"03",X"3F",X"7F",X"FF",
		X"E0",X"E0",X"F0",X"F8",X"F8",X"F8",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"F8",X"F6",X"EF",X"E7",X"E5",X"E2",X"E1",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"12",X"1A",X"3F",X"FF",X"FF",
		X"00",X"20",X"20",X"00",X"00",X"10",X"00",X"D0",X"E8",X"60",X"E0",X"E0",X"B0",X"70",X"F0",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C4",X"F0",X"60",X"E0",X"E0",X"B0",X"70",X"F0",X"FC",
		X"F8",X"D8",X"F8",X"FA",X"C0",X"80",X"C2",X"C2",X"C0",X"E0",X"E0",X"F0",X"F0",X"F0",X"E0",X"00",
		X"F8",X"D9",X"F8",X"F9",X"C0",X"80",X"C0",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F0",X"E0",X"00",
		X"7F",X"70",X"E0",X"EC",X"EE",X"EF",X"C5",X"D2",X"85",X"82",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"03",X"03",X"03",X"03",X"07",X"07",X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",X"1F",X"FF",X"0F",X"00",X"1F",X"1F",X"0F",X"C0",X"40",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",X"1F",X"0F",X"0F",X"00",X"1F",X"1F",X"0F",X"08",X"00",X"10",
		X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"07",X"0F",X"1F",X"1F",X"3F",X"3F",X"7F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"F3",X"E3",X"E7",X"E7",X"FF",X"FE",X"FE",X"3E",X"0C",X"00",X"02",X"01",X"00",
		X"FF",X"FF",X"FF",X"F3",X"E3",X"E7",X"E7",X"FF",X"FE",X"FE",X"3E",X"0C",X"00",X"04",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"0F",X"3F",X"DF",X"9E",X"3C",X"7E",
		X"00",X"38",X"68",X"C4",X"84",X"06",X"0C",X"98",X"FA",X"FE",X"8C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"7F",X"BE",X"DC",X"E9",X"F7",X"7B",X"7E",X"B8",X"10",X"00",X"00",X"20",X"10",X"00",X"00",
		X"FF",X"7E",X"BE",X"DC",X"E9",X"F7",X"7B",X"7E",X"B8",X"50",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"E0",X"C0",X"E0",X"38",X"9C",X"9F",X"FF",X"F8",X"C0",X"C0",X"C0",X"E1",X"FF",X"FF",X"F7",
		X"00",X"E0",X"C0",X"E0",X"38",X"9C",X"9F",X"FF",X"F8",X"C0",X"C0",X"C0",X"E1",X"FF",X"FF",X"F7",
		X"00",X"00",X"40",X"C0",X"80",X"F8",X"FC",X"E2",X"86",X"1C",X"E8",X"E0",X"E2",X"F6",X"F4",X"F0",
		X"F1",X"7B",X"3A",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C7",X"8F",X"FF",X"FD",X"F9",X"69",X"09",X"09",X"09",X"08",X"08",X"00",X"00",X"00",X"00",X"00",
		X"C7",X"8F",X"FF",X"FD",X"F9",X"69",X"09",X"09",X"09",X"08",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FC",X"F8",X"78",X"2C",X"2F",X"27",X"FF",X"FF",X"FF",X"E0",X"C0",X"E0",X"FF",X"FF",
		X"00",X"00",X"FC",X"F8",X"78",X"2C",X"2F",X"27",X"FF",X"FF",X"FF",X"E0",X"C0",X"E0",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"E0",X"F0",X"FC",X"81",
		X"C3",X"FE",X"F0",X"F0",X"F0",X"F6",X"F6",X"70",X"70",X"30",X"3E",X"1C",X"00",X"00",X"00",X"00",
		X"FF",X"97",X"F3",X"FF",X"FF",X"FF",X"22",X"22",X"22",X"24",X"44",X"44",X"00",X"FF",X"FE",X"00",
		X"FF",X"97",X"F3",X"FF",X"FF",X"FF",X"22",X"22",X"22",X"24",X"44",X"44",X"00",X"FF",X"FE",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
