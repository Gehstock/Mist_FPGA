library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity galaga_cpu3 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of galaga_cpu3 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"31",X"00",X"9B",X"C3",X"7B",X"00",X"FF",X"FF",X"87",X"30",X"05",X"24",X"18",X"02",X"FF",X"FF",
		X"85",X"6F",X"D0",X"24",X"C9",X"FF",X"FF",X"FF",X"77",X"23",X"10",X"FC",X"C9",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F5",X"C5",X"D5",X"E5",X"3E",X"01",X"32",X"22",X"68",X"AF",
		X"32",X"22",X"68",X"CD",X"B1",X"00",X"E1",X"D1",X"C1",X"F1",X"C9",X"3E",X"01",X"32",X"22",X"68",
		X"11",X"01",X"91",X"1A",X"A7",X"20",X"FC",X"67",X"6F",X"01",X"10",X"00",X"86",X"23",X"10",X"FC",
		X"0D",X"20",X"F9",X"FE",X"FF",X"28",X"02",X"3E",X"21",X"12",X"1A",X"A7",X"20",X"FC",X"AF",X"32",
		X"22",X"68",X"21",X"00",X"9A",X"36",X"00",X"11",X"01",X"9A",X"01",X"FF",X"00",X"ED",X"B0",X"18",
		X"FE",X"3A",X"B8",X"9A",X"A7",X"C2",X"A1",X"06",X"21",X"60",X"9A",X"36",X"00",X"11",X"61",X"9A",
		X"01",X"0F",X"00",X"ED",X"B0",X"3A",X"B7",X"9A",X"A7",X"C2",X"42",X"03",X"3A",X"79",X"9A",X"A7",
		X"28",X"09",X"21",X"A8",X"9A",X"86",X"77",X"AF",X"32",X"79",X"9A",X"3A",X"A0",X"9A",X"A7",X"28",
		X"6F",X"3A",X"11",X"92",X"21",X"80",X"9A",X"BE",X"28",X"20",X"32",X"80",X"9A",X"3C",X"28",X"0C",
		X"21",X"EA",X"06",X"22",X"82",X"9A",X"AF",X"32",X"00",X"9A",X"18",X"09",X"21",X"FA",X"06",X"22",
		X"82",X"9A",X"32",X"00",X"9A",X"32",X"81",X"9A",X"18",X"12",X"21",X"00",X"9A",X"34",X"7E",X"FE",
		X"22",X"20",X"1E",X"36",X"00",X"3A",X"81",X"9A",X"3C",X"32",X"81",X"9A",X"2A",X"82",X"9A",X"CF",
		X"5E",X"23",X"56",X"ED",X"53",X"84",X"9A",X"3E",X"1F",X"D7",X"5E",X"23",X"56",X"ED",X"53",X"86",
		X"9A",X"2A",X"86",X"9A",X"ED",X"5B",X"84",X"9A",X"19",X"22",X"86",X"9A",X"7C",X"32",X"61",X"9A",
		X"0F",X"0F",X"0F",X"0F",X"32",X"62",X"9A",X"3E",X"0A",X"32",X"65",X"9A",X"AF",X"32",X"70",X"9A",
		X"21",X"74",X"9A",X"36",X"13",X"3A",X"B3",X"9A",X"A7",X"28",X"09",X"AF",X"32",X"B3",X"9A",X"CD",
		X"F9",X"03",X"18",X"09",X"3A",X"D3",X"9A",X"A7",X"28",X"03",X"CD",X"4F",X"04",X"21",X"74",X"9A",
		X"36",X"0F",X"3A",X"AF",X"9A",X"A7",X"28",X"09",X"AF",X"32",X"AF",X"9A",X"CD",X"F9",X"03",X"18",
		X"09",X"3A",X"CF",X"9A",X"A7",X"28",X"03",X"CD",X"4F",X"04",X"21",X"74",X"9A",X"36",X"03",X"3A",
		X"A3",X"9A",X"A7",X"28",X"09",X"AF",X"32",X"A3",X"9A",X"CD",X"F9",X"03",X"18",X"09",X"3A",X"C3",
		X"9A",X"A7",X"28",X"03",X"CD",X"4F",X"04",X"21",X"74",X"9A",X"36",X"02",X"3A",X"A2",X"9A",X"A7",
		X"28",X"09",X"AF",X"32",X"A2",X"9A",X"CD",X"F9",X"03",X"18",X"09",X"3A",X"C2",X"9A",X"A7",X"28",
		X"03",X"CD",X"4F",X"04",X"21",X"74",X"9A",X"36",X"04",X"3A",X"A4",X"9A",X"A7",X"28",X"09",X"AF",
		X"32",X"A4",X"9A",X"CD",X"F9",X"03",X"18",X"09",X"3A",X"C4",X"9A",X"A7",X"28",X"03",X"CD",X"4F",
		X"04",X"21",X"74",X"9A",X"36",X"01",X"3A",X"A1",X"9A",X"A7",X"28",X"09",X"AF",X"32",X"A1",X"9A",
		X"CD",X"F9",X"03",X"18",X"09",X"3A",X"C1",X"9A",X"A7",X"28",X"03",X"CD",X"4F",X"04",X"3A",X"B2",
		X"9A",X"A7",X"28",X"08",X"21",X"74",X"9A",X"36",X"12",X"CD",X"A7",X"04",X"3A",X"A5",X"9A",X"A7",
		X"28",X"2C",X"21",X"74",X"9A",X"36",X"05",X"CD",X"7A",X"03",X"21",X"7E",X"9A",X"34",X"3A",X"7E",
		X"9A",X"FE",X"06",X"38",X"11",X"36",X"00",X"3A",X"7C",X"9A",X"FE",X"04",X"38",X"03",X"3D",X"18",
		X"02",X"3E",X"0C",X"32",X"7C",X"9A",X"3A",X"7C",X"9A",X"32",X"6F",X"9A",X"18",X"03",X"32",X"C5",
		X"9A",X"3A",X"A6",X"9A",X"A7",X"28",X"24",X"21",X"74",X"9A",X"36",X"06",X"CD",X"7A",X"03",X"21",
		X"7F",X"9A",X"34",X"7E",X"FE",X"1C",X"20",X"0B",X"AF",X"32",X"7F",X"9A",X"3A",X"7D",X"9A",X"3C",
		X"32",X"7D",X"9A",X"3A",X"7D",X"9A",X"32",X"70",X"9A",X"18",X"03",X"32",X"C6",X"9A",X"3A",X"A9",
		X"9A",X"A7",X"28",X"0A",X"21",X"74",X"9A",X"36",X"09",X"CD",X"7A",X"03",X"18",X"03",X"32",X"C9",
		X"9A",X"3A",X"A7",X"9A",X"A7",X"28",X"0B",X"21",X"74",X"9A",X"36",X"07",X"CD",X"A7",X"04",X"C3",
		X"32",X"03",X"3A",X"B1",X"9A",X"A7",X"28",X"0A",X"21",X"74",X"9A",X"36",X"11",X"CD",X"7A",X"03",
		X"18",X"03",X"32",X"D1",X"9A",X"3A",X"AD",X"9A",X"A7",X"28",X"08",X"21",X"74",X"9A",X"36",X"0D",
		X"CD",X"A7",X"04",X"3A",X"AE",X"9A",X"A7",X"28",X"12",X"21",X"74",X"9A",X"36",X"0E",X"CD",X"A7",
		X"04",X"3E",X"09",X"32",X"6A",X"9A",X"3E",X"06",X"32",X"6F",X"9A",X"3A",X"B4",X"9A",X"A7",X"28",
		X"08",X"21",X"74",X"9A",X"36",X"14",X"CD",X"A7",X"04",X"3A",X"B5",X"9A",X"A7",X"28",X"08",X"21",
		X"74",X"9A",X"36",X"15",X"CD",X"A7",X"04",X"3A",X"AA",X"9A",X"A7",X"28",X"08",X"21",X"74",X"9A",
		X"36",X"0A",X"CD",X"A7",X"04",X"3A",X"AB",X"9A",X"A7",X"28",X"08",X"21",X"74",X"9A",X"36",X"0B",
		X"CD",X"A7",X"04",X"3A",X"B0",X"9A",X"A7",X"28",X"0A",X"21",X"74",X"9A",X"36",X"10",X"CD",X"7A",
		X"03",X"18",X"03",X"32",X"D0",X"9A",X"3A",X"AC",X"9A",X"A7",X"28",X"08",X"21",X"74",X"9A",X"36",
		X"0C",X"CD",X"A7",X"04",X"3A",X"B6",X"9A",X"A7",X"28",X"08",X"21",X"74",X"9A",X"36",X"16",X"CD",
		X"A7",X"04",X"3A",X"A8",X"9A",X"A7",X"28",X"08",X"21",X"74",X"9A",X"36",X"08",X"CD",X"A7",X"04",
		X"18",X"1A",X"21",X"A0",X"9A",X"36",X"00",X"11",X"A1",X"9A",X"01",X"15",X"00",X"ED",X"B0",X"21",
		X"C0",X"9A",X"36",X"00",X"11",X"C1",X"9A",X"01",X"16",X"00",X"ED",X"B0",X"21",X"60",X"9A",X"11",
		X"10",X"68",X"01",X"10",X"00",X"ED",X"B0",X"3A",X"70",X"9A",X"32",X"05",X"68",X"3A",X"71",X"9A",
		X"32",X"0A",X"68",X"3A",X"72",X"9A",X"32",X"0F",X"68",X"C9",X"21",X"74",X"9A",X"7E",X"87",X"86",
		X"21",X"2A",X"07",X"D7",X"11",X"75",X"9A",X"01",X"03",X"00",X"ED",X"B0",X"3A",X"74",X"9A",X"FE",
		X"0E",X"20",X"18",X"3A",X"4C",X"9A",X"A7",X"28",X"0D",X"3D",X"28",X"06",X"3A",X"4D",X"9A",X"A7",
		X"20",X"09",X"3E",X"02",X"18",X"02",X"3E",X"01",X"32",X"76",X"9A",X"21",X"C0",X"9A",X"3A",X"74",
		X"9A",X"85",X"6F",X"7E",X"A7",X"20",X"1B",X"34",X"21",X"76",X"9A",X"46",X"48",X"21",X"30",X"9A",
		X"3A",X"75",X"9A",X"85",X"6F",X"AF",X"DF",X"41",X"21",X"00",X"9A",X"3A",X"75",X"9A",X"85",X"6F",
		X"AF",X"DF",X"CD",X"77",X"05",X"21",X"76",X"9A",X"35",X"28",X"0A",X"21",X"75",X"9A",X"34",X"21",
		X"77",X"9A",X"34",X"18",X"ED",X"3A",X"78",X"9A",X"A7",X"C8",X"AF",X"32",X"78",X"9A",X"21",X"C0",
		X"9A",X"3A",X"74",X"9A",X"85",X"6F",X"36",X"00",X"C9",X"21",X"C0",X"9A",X"3A",X"74",X"9A",X"85",
		X"6F",X"34",X"21",X"74",X"9A",X"7E",X"87",X"86",X"21",X"2A",X"07",X"D7",X"11",X"75",X"9A",X"01",
		X"03",X"00",X"ED",X"B0",X"3A",X"74",X"9A",X"FE",X"0E",X"20",X"18",X"3A",X"4C",X"9A",X"A7",X"28",
		X"0D",X"3D",X"28",X"06",X"3A",X"4D",X"9A",X"A7",X"20",X"09",X"3E",X"02",X"18",X"02",X"3E",X"01",
		X"32",X"76",X"9A",X"21",X"76",X"9A",X"46",X"48",X"21",X"30",X"9A",X"3A",X"75",X"9A",X"85",X"6F",
		X"AF",X"DF",X"41",X"21",X"00",X"9A",X"3A",X"75",X"9A",X"85",X"6F",X"AF",X"DF",X"18",X"31",X"21",
		X"74",X"9A",X"7E",X"87",X"86",X"21",X"2A",X"07",X"D7",X"11",X"75",X"9A",X"01",X"03",X"00",X"ED",
		X"B0",X"3A",X"74",X"9A",X"FE",X"0E",X"20",X"18",X"3A",X"4C",X"9A",X"A7",X"28",X"0D",X"3D",X"28",
		X"06",X"3A",X"4D",X"9A",X"A7",X"20",X"09",X"3E",X"02",X"18",X"02",X"3E",X"01",X"32",X"76",X"9A",
		X"CD",X"77",X"05",X"21",X"76",X"9A",X"35",X"28",X"0A",X"21",X"75",X"9A",X"34",X"21",X"77",X"9A",
		X"34",X"18",X"ED",X"3A",X"78",X"9A",X"A7",X"C8",X"AF",X"32",X"78",X"9A",X"21",X"C0",X"9A",X"3A",
		X"74",X"9A",X"85",X"6F",X"36",X"00",X"C9",X"21",X"74",X"9A",X"7E",X"87",X"86",X"21",X"2A",X"07",
		X"D7",X"11",X"75",X"9A",X"01",X"03",X"00",X"ED",X"B0",X"3A",X"74",X"9A",X"FE",X"0E",X"20",X"18",
		X"3A",X"4C",X"9A",X"A7",X"28",X"0D",X"3D",X"28",X"06",X"3A",X"4D",X"9A",X"A7",X"20",X"09",X"3E",
		X"02",X"18",X"02",X"3E",X"01",X"32",X"76",X"9A",X"21",X"C0",X"9A",X"3A",X"74",X"9A",X"85",X"6F",
		X"7E",X"A7",X"20",X"1B",X"34",X"21",X"76",X"9A",X"46",X"48",X"21",X"30",X"9A",X"3A",X"75",X"9A",
		X"85",X"6F",X"AF",X"DF",X"41",X"21",X"00",X"9A",X"3A",X"75",X"9A",X"85",X"6F",X"AF",X"DF",X"CD",
		X"77",X"05",X"21",X"76",X"9A",X"35",X"28",X"0A",X"21",X"75",X"9A",X"34",X"21",X"77",X"9A",X"34",
		X"18",X"ED",X"3A",X"78",X"9A",X"A7",X"C8",X"AF",X"32",X"78",X"9A",X"21",X"C0",X"9A",X"3A",X"74",
		X"9A",X"85",X"6F",X"36",X"00",X"21",X"A0",X"9A",X"3A",X"74",X"9A",X"85",X"6F",X"3A",X"74",X"9A",
		X"FE",X"08",X"28",X"0F",X"FE",X"0C",X"28",X"0D",X"FE",X"14",X"28",X"15",X"FE",X"07",X"28",X"19",
		X"36",X"00",X"C9",X"35",X"C9",X"35",X"28",X"03",X"CB",X"46",X"C8",X"3E",X"01",X"32",X"B6",X"9A",
		X"C9",X"36",X"00",X"21",X"B3",X"9A",X"36",X"01",X"C9",X"36",X"00",X"21",X"A0",X"9A",X"AF",X"06",
		X"08",X"DF",X"23",X"77",X"23",X"23",X"06",X"0C",X"DF",X"21",X"C0",X"9A",X"06",X"08",X"DF",X"23",
		X"77",X"23",X"23",X"06",X"0C",X"DF",X"C9",X"21",X"00",X"9A",X"3A",X"75",X"9A",X"85",X"6F",X"34",
		X"3A",X"75",X"9A",X"21",X"6F",X"07",X"CF",X"5E",X"23",X"56",X"EB",X"11",X"88",X"9A",X"01",X"03",
		X"00",X"ED",X"B0",X"EB",X"21",X"30",X"9A",X"3A",X"75",X"9A",X"85",X"6F",X"7E",X"EB",X"D7",X"22",
		X"7A",X"9A",X"7E",X"3C",X"CA",X"B2",X"06",X"11",X"D0",X"06",X"2A",X"7A",X"9A",X"7E",X"E6",X"0F",
		X"EB",X"CF",X"4E",X"23",X"46",X"EB",X"7E",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"28",X"07",X"CB",
		X"38",X"CB",X"19",X"3D",X"20",X"F9",X"3A",X"77",X"9A",X"A7",X"28",X"0D",X"3D",X"28",X"05",X"21",
		X"6B",X"9A",X"18",X"08",X"21",X"66",X"9A",X"18",X"03",X"21",X"61",X"9A",X"71",X"7E",X"0F",X"0F",
		X"0F",X"0F",X"23",X"77",X"23",X"70",X"7E",X"0F",X"0F",X"0F",X"0F",X"23",X"77",X"3A",X"77",X"9A",
		X"A7",X"28",X"0D",X"3D",X"28",X"05",X"11",X"6F",X"9A",X"18",X"08",X"11",X"6A",X"9A",X"18",X"03",
		X"11",X"65",X"9A",X"2A",X"7A",X"9A",X"7E",X"D6",X"0C",X"28",X"44",X"3A",X"88",X"9A",X"A7",X"28",
		X"23",X"3D",X"28",X"10",X"21",X"00",X"9A",X"3A",X"75",X"9A",X"85",X"6F",X"7E",X"FE",X"06",X"30",
		X"13",X"2F",X"18",X"30",X"21",X"00",X"9A",X"3A",X"75",X"9A",X"85",X"6F",X"7E",X"FE",X"06",X"30",
		X"03",X"87",X"18",X"20",X"3A",X"89",X"9A",X"A7",X"28",X"18",X"47",X"21",X"00",X"9A",X"3A",X"75",
		X"9A",X"85",X"6F",X"7E",X"90",X"38",X"0B",X"D6",X"0A",X"30",X"04",X"ED",X"44",X"18",X"05",X"AF",
		X"18",X"02",X"3E",X"0A",X"12",X"21",X"70",X"9A",X"3A",X"77",X"9A",X"85",X"6F",X"3A",X"8A",X"9A",
		X"77",X"21",X"CD",X"07",X"3A",X"74",X"9A",X"D7",X"7E",X"2A",X"7A",X"9A",X"23",X"5E",X"16",X"00",
		X"21",X"00",X"00",X"06",X"08",X"CB",X"3F",X"30",X"01",X"19",X"CB",X"23",X"CB",X"12",X"10",X"F5",
		X"45",X"21",X"00",X"9A",X"3A",X"75",X"9A",X"85",X"6F",X"78",X"BE",X"C0",X"21",X"30",X"9A",X"3A",
		X"75",X"9A",X"85",X"6F",X"34",X"34",X"21",X"00",X"9A",X"3A",X"75",X"9A",X"85",X"6F",X"36",X"00",
		X"C9",X"21",X"00",X"9A",X"36",X"00",X"11",X"01",X"9A",X"01",X"FF",X"00",X"ED",X"B0",X"31",X"00",
		X"9B",X"C9",X"3A",X"77",X"9A",X"A7",X"28",X"0D",X"3D",X"28",X"05",X"21",X"6F",X"9A",X"18",X"08",
		X"21",X"6A",X"9A",X"18",X"03",X"21",X"65",X"9A",X"36",X"00",X"3E",X"01",X"32",X"78",X"9A",X"C9",
		X"50",X"81",X"00",X"89",X"26",X"91",X"C8",X"99",X"EC",X"A2",X"9D",X"AC",X"E0",X"B6",X"C0",X"C1",
		X"45",X"CD",X"7A",X"D9",X"69",X"E6",X"1C",X"F4",X"00",X"00",X"30",X"01",X"68",X"01",X"36",X"01",
		X"A8",X"01",X"68",X"01",X"00",X"02",X"AC",X"01",X"08",X"02",X"00",X"FE",X"58",X"FE",X"08",X"FE",
		X"98",X"FE",X"58",X"FE",X"D0",X"FE",X"98",X"FE",X"D6",X"FE",X"00",X"5B",X"00",X"6C",X"00",X"5B",
		X"00",X"7E",X"00",X"6C",X"00",X"97",X"00",X"81",X"00",X"99",X"00",X"D9",X"00",X"B6",X"00",X"D9",
		X"00",X"97",X"00",X"B6",X"00",X"7E",X"00",X"99",X"00",X"81",X"00",X"01",X"00",X"01",X"01",X"01",
		X"02",X"01",X"01",X"03",X"01",X"01",X"04",X"01",X"01",X"05",X"01",X"00",X"06",X"01",X"00",X"20",
		X"03",X"00",X"0A",X"03",X"00",X"0D",X"03",X"00",X"07",X"03",X"00",X"13",X"03",X"00",X"16",X"03",
		X"00",X"19",X"03",X"00",X"1C",X"03",X"00",X"1F",X"01",X"02",X"2C",X"03",X"00",X"10",X"03",X"00",
		X"23",X"01",X"00",X"24",X"01",X"00",X"25",X"03",X"00",X"28",X"01",X"00",X"29",X"03",X"00",X"E4",
		X"07",X"3B",X"08",X"19",X"08",X"E5",X"07",X"85",X"08",X"9F",X"08",X"B3",X"08",X"F9",X"09",X"09",
		X"0A",X"19",X"0A",X"C3",X"09",X"D5",X"09",X"E7",X"09",X"29",X"0A",X"6D",X"0A",X"B1",X"0A",X"DD",
		X"0A",X"21",X"0B",X"65",X"0B",X"C7",X"08",X"13",X"09",X"5D",X"09",X"83",X"0C",X"11",X"0D",X"5F",
		X"0D",X"8D",X"09",X"9F",X"09",X"B1",X"09",X"C7",X"08",X"C7",X"08",X"C7",X"08",X"2F",X"0C",X"91",
		X"0B",X"C7",X"0B",X"FD",X"0B",X"1B",X"0C",X"2F",X"0C",X"93",X"0D",X"07",X"0E",X"83",X"0E",X"85",
		X"0D",X"07",X"0D",X"55",X"0D",X"7B",X"0D",X"C5",X"0E",X"01",X"0F",X"3D",X"0F",X"04",X"02",X"02",
		X"02",X"02",X"04",X"04",X"0A",X"07",X"0C",X"0B",X"04",X"0A",X"0D",X"04",X"01",X"04",X"0C",X"02",
		X"06",X"05",X"02",X"0A",X"FF",X"00",X"00",X"06",X"71",X"01",X"72",X"01",X"73",X"01",X"75",X"01",
		X"74",X"01",X"73",X"01",X"72",X"01",X"71",X"01",X"70",X"01",X"8B",X"01",X"8A",X"01",X"0C",X"04",
		X"86",X"01",X"87",X"01",X"88",X"01",X"89",X"01",X"8A",X"01",X"89",X"01",X"88",X"01",X"87",X"01",
		X"86",X"01",X"85",X"01",X"84",X"01",X"83",X"01",X"FF",X"00",X"00",X"04",X"88",X"01",X"8A",X"01",
		X"70",X"01",X"71",X"01",X"73",X"01",X"75",X"01",X"77",X"01",X"78",X"01",X"0C",X"06",X"74",X"01",
		X"73",X"01",X"72",X"01",X"71",X"01",X"70",X"01",X"8B",X"01",X"FF",X"00",X"00",X"07",X"89",X"01",
		X"8A",X"01",X"8B",X"01",X"0C",X"01",X"70",X"01",X"71",X"01",X"72",X"01",X"0C",X"01",X"73",X"01",
		X"74",X"01",X"75",X"01",X"0C",X"03",X"8B",X"01",X"70",X"01",X"71",X"01",X"0C",X"01",X"72",X"01",
		X"73",X"01",X"74",X"01",X"0C",X"01",X"75",X"01",X"76",X"01",X"77",X"01",X"0C",X"03",X"71",X"01",
		X"72",X"01",X"73",X"01",X"0C",X"01",X"74",X"01",X"75",X"01",X"76",X"01",X"0C",X"01",X"77",X"01",
		X"78",X"01",X"79",X"01",X"FF",X"00",X"00",X"05",X"71",X"01",X"72",X"01",X"73",X"01",X"0C",X"01",
		X"74",X"01",X"75",X"01",X"76",X"01",X"0C",X"01",X"77",X"01",X"78",X"01",X"79",X"01",X"FF",X"00",
		X"00",X"04",X"61",X"01",X"7A",X"01",X"60",X"01",X"78",X"01",X"7A",X"01",X"76",X"01",X"78",X"01",
		X"75",X"01",X"FF",X"00",X"00",X"00",X"76",X"01",X"79",X"01",X"60",X"01",X"63",X"01",X"66",X"01",
		X"63",X"01",X"60",X"01",X"79",X"01",X"FF",X"00",X"00",X"07",X"81",X"08",X"81",X"01",X"86",X"03",
		X"88",X"09",X"8B",X"03",X"8A",X"09",X"86",X"03",X"88",X"09",X"73",X"03",X"71",X"09",X"86",X"03",
		X"88",X"09",X"8B",X"03",X"8A",X"09",X"86",X"03",X"71",X"09",X"75",X"03",X"76",X"09",X"74",X"03",
		X"72",X"09",X"71",X"03",X"8B",X"09",X"89",X"03",X"88",X"09",X"84",X"03",X"74",X"09",X"76",X"03",
		X"74",X"09",X"71",X"03",X"73",X"04",X"8B",X"04",X"88",X"04",X"71",X"04",X"8A",X"04",X"88",X"04",
		X"0C",X"10",X"FF",X"00",X"00",X"06",X"8A",X"09",X"81",X"03",X"88",X"09",X"83",X"03",X"86",X"09",
		X"81",X"03",X"83",X"09",X"85",X"03",X"8A",X"09",X"81",X"03",X"88",X"09",X"83",X"03",X"86",X"09",
		X"81",X"03",X"88",X"09",X"71",X"03",X"72",X"09",X"71",X"03",X"8B",X"09",X"89",X"03",X"88",X"09",
		X"86",X"03",X"84",X"09",X"88",X"03",X"89",X"09",X"8B",X"03",X"89",X"09",X"86",X"03",X"8B",X"04",
		X"88",X"04",X"83",X"04",X"88",X"04",X"85",X"04",X"83",X"04",X"0C",X"10",X"FF",X"00",X"00",X"07",
		X"81",X"0C",X"83",X"09",X"86",X"03",X"85",X"0C",X"81",X"0C",X"86",X"0C",X"88",X"09",X"8B",X"03",
		X"8A",X"0C",X"88",X"0C",X"89",X"0C",X"88",X"09",X"86",X"03",X"84",X"0C",X"89",X"0C",X"74",X"0C",
		X"71",X"09",X"89",X"03",X"88",X"0C",X"71",X"09",X"8A",X"03",X"0C",X"10",X"FF",X"02",X"00",X"03",
		X"78",X"02",X"0C",X"01",X"78",X"01",X"79",X"01",X"7B",X"01",X"61",X"03",X"0C",X"03",X"FF",X"02",
		X"00",X"03",X"73",X"02",X"0C",X"01",X"73",X"01",X"74",X"01",X"76",X"01",X"78",X"03",X"0C",X"02",
		X"FF",X"02",X"00",X"03",X"70",X"02",X"0C",X"01",X"70",X"01",X"71",X"01",X"73",X"01",X"75",X"03",
		X"0C",X"02",X"FF",X"01",X"00",X"04",X"78",X"01",X"7A",X"01",X"63",X"01",X"78",X"01",X"7A",X"01",
		X"63",X"01",X"65",X"03",X"FF",X"01",X"00",X"05",X"73",X"01",X"78",X"01",X"7A",X"01",X"73",X"01",
		X"78",X"01",X"7A",X"01",X"60",X"03",X"FF",X"01",X"00",X"07",X"8A",X"01",X"73",X"01",X"78",X"01",
		X"8A",X"01",X"73",X"01",X"78",X"01",X"7A",X"03",X"FF",X"01",X"06",X"04",X"7A",X"01",X"78",X"01",
		X"7A",X"01",X"61",X"01",X"65",X"01",X"68",X"03",X"FF",X"01",X"06",X"04",X"78",X"01",X"75",X"01",
		X"78",X"01",X"7A",X"01",X"61",X"01",X"65",X"03",X"FF",X"01",X"06",X"04",X"75",X"01",X"71",X"01",
		X"75",X"01",X"78",X"01",X"7A",X"01",X"60",X"03",X"FF",X"02",X"04",X"03",X"7A",X"01",X"76",X"01",
		X"78",X"01",X"75",X"01",X"76",X"01",X"73",X"01",X"75",X"01",X"72",X"01",X"73",X"01",X"8A",X"01",
		X"8B",X"01",X"88",X"01",X"86",X"01",X"85",X"01",X"83",X"01",X"82",X"01",X"83",X"01",X"86",X"01",
		X"85",X"01",X"88",X"01",X"86",X"01",X"8A",X"01",X"88",X"01",X"8B",X"01",X"8A",X"01",X"73",X"01",
		X"72",X"01",X"73",X"01",X"75",X"01",X"8A",X"01",X"70",X"01",X"72",X"01",X"FF",X"02",X"04",X"03",
		X"76",X"01",X"73",X"01",X"75",X"01",X"72",X"01",X"73",X"01",X"70",X"01",X"72",X"01",X"8A",X"01",
		X"8B",X"01",X"86",X"01",X"88",X"01",X"85",X"01",X"83",X"01",X"82",X"01",X"80",X"01",X"9A",X"01",
		X"9A",X"01",X"83",X"01",X"82",X"01",X"85",X"01",X"83",X"01",X"86",X"01",X"85",X"01",X"88",X"01",
		X"86",X"01",X"8A",X"01",X"88",X"01",X"8B",X"01",X"8A",X"01",X"88",X"01",X"86",X"01",X"85",X"01",
		X"FF",X"02",X"10",X"03",X"93",X"02",X"9A",X"02",X"83",X"03",X"9A",X"01",X"98",X"01",X"96",X"01",
		X"95",X"01",X"93",X"02",X"95",X"03",X"96",X"02",X"98",X"02",X"9A",X"02",X"9B",X"02",X"9A",X"02",
		X"98",X"01",X"96",X"01",X"95",X"01",X"92",X"01",X"93",X"01",X"95",X"01",X"FF",X"02",X"04",X"03",
		X"7A",X"01",X"77",X"01",X"78",X"01",X"75",X"01",X"77",X"01",X"73",X"01",X"75",X"01",X"72",X"01",
		X"73",X"01",X"8A",X"01",X"80",X"01",X"88",X"01",X"87",X"01",X"85",X"01",X"83",X"01",X"82",X"01",
		X"83",X"01",X"87",X"01",X"85",X"01",X"88",X"01",X"87",X"01",X"8A",X"01",X"88",X"01",X"80",X"01",
		X"8A",X"01",X"73",X"01",X"72",X"01",X"73",X"01",X"75",X"01",X"8A",X"01",X"70",X"01",X"72",X"01",
		X"FF",X"02",X"04",X"03",X"77",X"01",X"73",X"01",X"75",X"01",X"72",X"01",X"73",X"01",X"70",X"01",
		X"72",X"01",X"8A",X"01",X"80",X"01",X"87",X"01",X"88",X"01",X"85",X"01",X"83",X"01",X"82",X"01",
		X"80",X"01",X"9A",X"01",X"9A",X"01",X"83",X"01",X"82",X"01",X"85",X"01",X"83",X"01",X"87",X"01",
		X"85",X"01",X"88",X"01",X"87",X"01",X"8A",X"01",X"88",X"01",X"80",X"01",X"8A",X"01",X"88",X"01",
		X"87",X"01",X"85",X"01",X"FF",X"02",X"10",X"03",X"93",X"02",X"9A",X"02",X"83",X"03",X"9A",X"01",
		X"98",X"01",X"97",X"01",X"95",X"01",X"93",X"02",X"95",X"03",X"97",X"02",X"98",X"02",X"9A",X"02",
		X"90",X"02",X"9A",X"02",X"98",X"01",X"97",X"01",X"95",X"01",X"92",X"01",X"93",X"01",X"95",X"01",
		X"FF",X"02",X"04",X"03",X"7A",X"01",X"76",X"01",X"78",X"01",X"75",X"01",X"76",X"01",X"73",X"01",
		X"75",X"01",X"72",X"01",X"73",X"01",X"8A",X"01",X"8A",X"01",X"88",X"01",X"86",X"01",X"85",X"01",
		X"83",X"01",X"82",X"01",X"83",X"01",X"85",X"01",X"86",X"01",X"88",X"01",X"86",X"01",X"8A",X"01",
		X"70",X"01",X"72",X"01",X"73",X"04",X"FF",X"02",X"04",X"03",X"76",X"01",X"73",X"01",X"75",X"01",
		X"72",X"01",X"73",X"01",X"70",X"01",X"72",X"01",X"8A",X"01",X"8A",X"01",X"86",X"01",X"86",X"01",
		X"85",X"01",X"83",X"01",X"82",X"01",X"80",X"01",X"9A",X"01",X"9A",X"01",X"8B",X"01",X"80",X"01",
		X"82",X"01",X"83",X"01",X"85",X"01",X"86",X"01",X"88",X"01",X"8A",X"04",X"FF",X"02",X"10",X"03",
		X"73",X"02",X"75",X"02",X"76",X"02",X"75",X"02",X"73",X"02",X"72",X"02",X"70",X"02",X"72",X"02",
		X"73",X"02",X"8B",X"02",X"8A",X"02",X"86",X"02",X"83",X"04",X"FF",X"00",X"00",X"04",X"71",X"04",
		X"73",X"04",X"71",X"04",X"73",X"04",X"76",X"04",X"78",X"04",X"76",X"04",X"78",X"04",X"FF",X"00",
		X"00",X"06",X"56",X"01",X"55",X"01",X"54",X"01",X"53",X"01",X"52",X"01",X"51",X"01",X"50",X"01",
		X"6B",X"01",X"6A",X"01",X"69",X"01",X"68",X"01",X"67",X"01",X"66",X"01",X"65",X"01",X"64",X"01",
		X"63",X"01",X"62",X"01",X"61",X"01",X"60",X"01",X"7B",X"01",X"7A",X"01",X"79",X"01",X"78",X"01",
		X"77",X"01",X"76",X"01",X"75",X"01",X"74",X"01",X"73",X"01",X"72",X"01",X"71",X"01",X"70",X"01",
		X"8B",X"01",X"8A",X"01",X"89",X"01",X"88",X"01",X"87",X"01",X"86",X"01",X"85",X"01",X"84",X"01",
		X"83",X"01",X"FF",X"02",X"04",X"05",X"60",X"01",X"78",X"01",X"75",X"01",X"71",X"01",X"60",X"01",
		X"78",X"01",X"75",X"01",X"71",X"01",X"60",X"01",X"78",X"01",X"75",X"01",X"71",X"01",X"60",X"01",
		X"78",X"01",X"75",X"01",X"71",X"01",X"60",X"01",X"78",X"01",X"75",X"01",X"71",X"01",X"60",X"01",
		X"78",X"01",X"75",X"01",X"71",X"01",X"60",X"01",X"0C",X"01",X"78",X"01",X"7A",X"01",X"75",X"01",
		X"78",X"01",X"73",X"01",X"75",X"01",X"61",X"01",X"7A",X"01",X"76",X"01",X"73",X"01",X"61",X"01",
		X"7A",X"01",X"76",X"01",X"73",X"01",X"61",X"01",X"7A",X"01",X"76",X"01",X"73",X"01",X"61",X"01",
		X"7A",X"01",X"76",X"01",X"73",X"01",X"61",X"01",X"79",X"01",X"76",X"01",X"73",X"01",X"61",X"01",
		X"79",X"01",X"76",X"01",X"73",X"01",X"61",X"01",X"0C",X"01",X"79",X"01",X"61",X"01",X"78",X"01",
		X"79",X"01",X"75",X"01",X"78",X"01",X"FF",X"02",X"02",X"05",X"60",X"01",X"60",X"01",X"60",X"01",
		X"FF",X"02",X"04",X"05",X"61",X"02",X"78",X"02",X"78",X"02",X"61",X"02",X"78",X"02",X"78",X"02",
		X"61",X"02",X"78",X"02",X"78",X"02",X"61",X"02",X"78",X"02",X"78",X"02",X"61",X"02",X"78",X"02",
		X"7A",X"02",X"75",X"02",X"63",X"02",X"7A",X"02",X"7A",X"02",X"63",X"02",X"7A",X"02",X"7A",X"02",
		X"63",X"02",X"7A",X"02",X"79",X"02",X"63",X"02",X"79",X"02",X"79",X"02",X"63",X"02",X"79",X"02",
		X"76",X"02",X"73",X"02",X"FF",X"02",X"02",X"05",X"78",X"01",X"78",X"01",X"78",X"01",X"FF",X"02",
		X"10",X"05",X"85",X"06",X"85",X"06",X"85",X"06",X"85",X"06",X"85",X"04",X"85",X"04",X"86",X"06",
		X"86",X"06",X"86",X"06",X"86",X"06",X"86",X"04",X"86",X"04",X"FF",X"02",X"04",X"05",X"81",X"01",
		X"81",X"01",X"81",X"01",X"FF",X"02",X"00",X"07",X"65",X"01",X"0C",X"01",X"61",X"01",X"0C",X"01",
		X"63",X"01",X"FF",X"02",X"00",X"05",X"7A",X"05",X"0C",X"01",X"7A",X"01",X"0C",X"01",X"7A",X"03",
		X"0C",X"01",X"78",X"07",X"0C",X"01",X"78",X"07",X"0C",X"01",X"78",X"03",X"0C",X"01",X"7B",X"05",
		X"0C",X"01",X"7B",X"01",X"0C",X"01",X"7B",X"03",X"0C",X"01",X"7A",X"07",X"0C",X"01",X"7A",X"07",
		X"0C",X"01",X"7A",X"03",X"0C",X"01",X"7B",X"01",X"0C",X"01",X"7B",X"01",X"0C",X"03",X"7B",X"01",
		X"0C",X"01",X"7B",X"03",X"0C",X"01",X"61",X"01",X"0C",X"01",X"61",X"01",X"0C",X"03",X"61",X"01",
		X"0C",X"01",X"61",X"03",X"0C",X"01",X"61",X"03",X"0C",X"01",X"61",X"03",X"0C",X"01",X"63",X"01",
		X"0C",X"01",X"63",X"01",X"0C",X"03",X"63",X"01",X"0C",X"01",X"63",X"03",X"0C",X"01",X"63",X"03",
		X"0C",X"01",X"63",X"03",X"0C",X"01",X"FF",X"02",X"00",X"03",X"86",X"02",X"8A",X"02",X"71",X"02",
		X"76",X"02",X"86",X"02",X"8A",X"02",X"71",X"02",X"76",X"02",X"86",X"02",X"8A",X"02",X"71",X"02",
		X"76",X"02",X"86",X"02",X"8A",X"02",X"71",X"02",X"76",X"02",X"86",X"02",X"8A",X"02",X"71",X"02",
		X"76",X"02",X"86",X"02",X"8A",X"02",X"71",X"02",X"76",X"02",X"86",X"02",X"8A",X"02",X"71",X"02",
		X"76",X"02",X"86",X"02",X"8A",X"02",X"71",X"02",X"76",X"02",X"77",X"01",X"0C",X"01",X"77",X"01",
		X"0C",X"03",X"77",X"01",X"0C",X"01",X"77",X"03",X"0C",X"01",X"69",X"01",X"0C",X"01",X"69",X"01",
		X"0C",X"03",X"69",X"01",X"0C",X"01",X"69",X"03",X"0C",X"01",X"69",X"03",X"0C",X"01",X"69",X"03",
		X"0C",X"01",X"8B",X"02",X"73",X"02",X"76",X"02",X"7B",X"02",X"7B",X"02",X"76",X"02",X"73",X"02",
		X"8B",X"02",X"FF",X"00",X"00",X"02",X"86",X"08",X"81",X"08",X"86",X"08",X"81",X"08",X"86",X"08",
		X"81",X"08",X"86",X"08",X"81",X"08",X"82",X"01",X"0C",X"01",X"82",X"01",X"0C",X"03",X"82",X"01",
		X"0C",X"01",X"82",X"03",X"0C",X"01",X"84",X"01",X"0C",X"01",X"84",X"01",X"0C",X"03",X"84",X"01",
		X"0C",X"01",X"84",X"03",X"0C",X"01",X"84",X"03",X"0C",X"01",X"84",X"03",X"0C",X"01",X"7B",X"08",
		X"76",X"04",X"8B",X"04",X"FF",X"00",X"0C",X"05",X"75",X"0C",X"71",X"0C",X"8A",X"0C",X"86",X"0C",
		X"0C",X"09",X"75",X"03",X"71",X"09",X"8A",X"03",X"86",X"04",X"8A",X"04",X"71",X"04",X"89",X"04",
		X"70",X"04",X"73",X"04",X"8B",X"0C",X"73",X"0C",X"76",X"0C",X"78",X"0C",X"0C",X"09",X"79",X"03",
		X"76",X"09",X"72",X"03",X"8B",X"04",X"89",X"04",X"86",X"04",X"72",X"04",X"89",X"04",X"76",X"04",
		X"FF",X"00",X"0C",X"05",X"71",X"0C",X"8A",X"0C",X"86",X"0C",X"85",X"0C",X"0C",X"09",X"81",X"03",
		X"8A",X"09",X"86",X"03",X"85",X"04",X"86",X"04",X"8A",X"04",X"86",X"04",X"89",X"04",X"8B",X"04",
		X"88",X"0C",X"8B",X"0C",X"73",X"0C",X"76",X"0C",X"0C",X"09",X"76",X"03",X"72",X"09",X"8B",X"03",
		X"8A",X"04",X"86",X"04",X"82",X"04",X"8B",X"04",X"89",X"04",X"82",X"04",X"FF",X"00",X"00",X"03",
		X"75",X"18",X"75",X"18",X"75",X"18",X"71",X"0C",X"75",X"0C",X"73",X"18",X"73",X"18",X"72",X"18",
		X"76",X"0C",X"78",X"0C",X"FF",X"FB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
