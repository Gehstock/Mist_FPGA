library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity romg is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of romg is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"D8",X"00",X"F8",X"00",X"FE",X"03",X"B8",X"00",X"F8",X"01",X"F8",X"00",X"60",X"00",X"F0",
		X"00",X"FC",X"07",X"FE",X"7F",X"FF",X"00",X"F9",X"00",X"F9",X"00",X"F9",X"00",X"FE",X"01",X"FE",
		X"01",X"02",X"11",X"50",X"00",X"D8",X"00",X"F8",X"00",X"FE",X"03",X"B8",X"00",X"F8",X"01",X"F8",
		X"00",X"60",X"00",X"F0",X"E0",X"FC",X"3F",X"FE",X"03",X"FF",X"00",X"F9",X"00",X"F9",X"00",X"F9",
		X"00",X"FE",X"01",X"FE",X"01",X"02",X"11",X"50",X"00",X"D8",X"00",X"F8",X"00",X"FE",X"03",X"B8",
		X"00",X"F8",X"01",X"F8",X"00",X"60",X"00",X"F0",X"70",X"FC",X"1F",X"FE",X"07",X"FF",X"00",X"F9",
		X"00",X"F9",X"00",X"F9",X"00",X"FE",X"01",X"FE",X"01",X"02",X"11",X"50",X"00",X"D8",X"00",X"F8",
		X"00",X"FE",X"03",X"B8",X"00",X"F8",X"01",X"F8",X"00",X"60",X"E0",X"F0",X"1C",X"FC",X"07",X"FE",
		X"03",X"FF",X"00",X"F9",X"00",X"F9",X"00",X"F9",X"00",X"FE",X"01",X"FE",X"01",X"02",X"11",X"50",
		X"00",X"D8",X"00",X"F8",X"00",X"FE",X"03",X"B8",X"40",X"F8",X"61",X"F8",X"30",X"60",X"18",X"F0",
		X"0C",X"FC",X"07",X"FE",X"03",X"FF",X"00",X"F9",X"00",X"F9",X"00",X"F9",X"00",X"FE",X"01",X"FE",
		X"01",X"02",X"09",X"FC",X"01",X"F8",X"03",X"98",X"03",X"18",X"07",X"1C",X"07",X"8E",X"03",X"86",
		X"01",X"C7",X"01",X"9E",X"07",X"02",X"09",X"FC",X"01",X"F8",X"01",X"F8",X"01",X"F0",X"01",X"E0",
		X"01",X"E0",X"00",X"C0",X"00",X"E0",X"00",X"C0",X"03",X"02",X"09",X"FC",X"00",X"F8",X"01",X"F0",
		X"03",X"C8",X"07",X"9C",X"07",X"0E",X"03",X"06",X"03",X"87",X"03",X"3E",X"0F",X"02",X"0F",X"28",
		X"00",X"68",X"00",X"78",X"00",X"FE",X"01",X"58",X"00",X"F8",X"00",X"78",X"00",X"30",X"00",X"FC",
		X"00",X"FE",X"01",X"7F",X"03",X"79",X"04",X"79",X"08",X"79",X"10",X"7E",X"00",X"02",X"0F",X"28",
		X"00",X"68",X"00",X"78",X"00",X"FE",X"01",X"58",X"00",X"F8",X"00",X"78",X"00",X"30",X"00",X"FC",
		X"00",X"FE",X"03",X"7F",X"0F",X"79",X"38",X"79",X"00",X"79",X"00",X"7E",X"00",X"02",X"0F",X"28",
		X"00",X"68",X"00",X"78",X"00",X"FE",X"01",X"58",X"00",X"F8",X"00",X"78",X"00",X"30",X"00",X"FC",
		X"07",X"FE",X"3F",X"7F",X"00",X"79",X"00",X"79",X"00",X"79",X"00",X"7E",X"00",X"02",X"0F",X"28",
		X"00",X"68",X"00",X"78",X"00",X"FE",X"01",X"58",X"00",X"F8",X"00",X"78",X"00",X"30",X"78",X"FC",
		X"0F",X"FE",X"00",X"7F",X"00",X"79",X"00",X"79",X"00",X"79",X"00",X"7E",X"00",X"02",X"0F",X"28",
		X"00",X"68",X"00",X"78",X"00",X"FE",X"01",X"58",X"00",X"F8",X"00",X"78",X"18",X"30",X"0E",X"FC",
		X"07",X"FE",X"01",X"7F",X"00",X"79",X"00",X"79",X"00",X"79",X"00",X"7E",X"00",X"02",X"0F",X"28",
		X"00",X"68",X"00",X"78",X"00",X"FE",X"01",X"58",X"00",X"F8",X"00",X"78",X"18",X"30",X"0E",X"FC",
		X"07",X"FE",X"01",X"7F",X"00",X"79",X"00",X"79",X"00",X"79",X"00",X"7E",X"00",X"02",X"0F",X"28",
		X"00",X"68",X"00",X"78",X"00",X"FE",X"11",X"58",X"08",X"F8",X"04",X"78",X"02",X"30",X"03",X"FC",
		X"01",X"FE",X"01",X"7F",X"00",X"79",X"00",X"79",X"00",X"79",X"00",X"7E",X"00",X"02",X"07",X"7E",
		X"00",X"EC",X"00",X"CC",X"01",X"8C",X"01",X"C6",X"00",X"63",X"00",X"CE",X"01",X"02",X"07",X"7C",
		X"00",X"78",X"00",X"78",X"00",X"70",X"00",X"30",X"00",X"20",X"00",X"E0",X"00",X"02",X"07",X"7E",
		X"00",X"F8",X"00",X"E0",X"01",X"CC",X"01",X"86",X"00",X"C3",X"00",X"8E",X"03",X"02",X"0E",X"14",
		X"00",X"34",X"00",X"3C",X"00",X"FF",X"00",X"2C",X"00",X"7C",X"00",X"3C",X"00",X"18",X"00",X"7C",
		X"00",X"FE",X"00",X"3F",X"01",X"3D",X"02",X"3D",X"04",X"3D",X"00",X"02",X"0E",X"14",X"00",X"34",
		X"00",X"3C",X"00",X"FF",X"00",X"2C",X"00",X"7C",X"00",X"3C",X"00",X"18",X"00",X"FC",X"00",X"FE",
		X"03",X"3F",X"0E",X"3D",X"00",X"3D",X"00",X"3D",X"00",X"02",X"0E",X"14",X"00",X"34",X"00",X"3C",
		X"00",X"FF",X"00",X"2C",X"00",X"7C",X"00",X"3C",X"00",X"18",X"00",X"FC",X"01",X"FE",X"0F",X"3F",
		X"00",X"3D",X"00",X"3D",X"00",X"3D",X"00",X"02",X"0E",X"14",X"00",X"34",X"00",X"3C",X"00",X"FF",
		X"00",X"2C",X"00",X"7C",X"00",X"3C",X"00",X"18",X"0E",X"FC",X"03",X"7E",X"00",X"3F",X"00",X"3D",
		X"00",X"3D",X"00",X"3D",X"00",X"02",X"0E",X"14",X"00",X"34",X"00",X"3C",X"00",X"FF",X"00",X"2C",
		X"00",X"7C",X"00",X"3C",X"00",X"18",X"0E",X"FC",X"03",X"FE",X"00",X"3F",X"00",X"3D",X"00",X"3D",
		X"00",X"3D",X"00",X"02",X"0E",X"14",X"00",X"34",X"00",X"3C",X"00",X"FF",X"00",X"2C",X"00",X"7C",
		X"00",X"3C",X"08",X"18",X"06",X"FC",X"03",X"FE",X"00",X"3F",X"00",X"3D",X"00",X"3D",X"00",X"3D",
		X"00",X"02",X"0E",X"14",X"00",X"34",X"00",X"3C",X"00",X"FF",X"04",X"2C",X"02",X"7C",X"02",X"3C",
		X"01",X"98",X"01",X"FC",X"00",X"7E",X"00",X"3F",X"00",X"3D",X"00",X"3D",X"00",X"3D",X"00",X"01",
		X"05",X"7E",X"64",X"32",X"11",X"77",X"01",X"05",X"3E",X"38",X"18",X"10",X"70",X"01",X"05",X"7E",
		X"70",X"26",X"21",X"E7",X"01",X"1A",X"18",X"38",X"38",X"38",X"38",X"38",X"3A",X"3A",X"BE",X"B8",
		X"B8",X"F8",X"FB",X"3B",X"3B",X"3B",X"3F",X"3C",X"38",X"38",X"38",X"38",X"38",X"38",X"38",X"38",
		X"01",X"15",X"08",X"18",X"18",X"18",X"18",X"1A",X"1E",X"D8",X"58",X"78",X"78",X"19",X"19",X"1F",
		X"1E",X"18",X"18",X"18",X"18",X"18",X"18",X"01",X"0F",X"10",X"10",X"10",X"18",X"50",X"70",X"14",
		X"14",X"14",X"1C",X"10",X"10",X"10",X"10",X"10",X"03",X"1C",X"00",X"7E",X"00",X"80",X"FF",X"01",
		X"E0",X"FF",X"07",X"F0",X"FF",X"0F",X"F0",X"FF",X"0F",X"F8",X"FF",X"1F",X"F8",X"FF",X"1F",X"F8",
		X"FF",X"1F",X"F8",X"E7",X"1F",X"F0",X"C3",X"0F",X"F0",X"81",X"0F",X"E0",X"81",X"07",X"C0",X"81",
		X"03",X"80",X"C3",X"01",X"F0",X"FF",X"0F",X"E0",X"FF",X"07",X"E0",X"FF",X"07",X"F4",X"FF",X"2F",
		X"84",X"C3",X"21",X"04",X"81",X"20",X"04",X"81",X"20",X"06",X"81",X"60",X"F7",X"FF",X"EF",X"06",
		X"81",X"60",X"04",X"00",X"20",X"04",X"00",X"20",X"04",X"00",X"20",X"04",X"00",X"20",X"03",X"19",
		X"00",X"1E",X"00",X"80",X"7F",X"00",X"C0",X"FF",X"00",X"E0",X"FF",X"01",X"F0",X"FF",X"03",X"F0",
		X"FF",X"03",X"F8",X"F3",X"07",X"F8",X"E1",X"07",X"F8",X"C0",X"07",X"F0",X"C0",X"03",X"E0",X"C0",
		X"01",X"C0",X"E1",X"00",X"80",X"7F",X"00",X"F0",X"FF",X"03",X"E0",X"FF",X"01",X"E0",X"FF",X"01",
		X"F4",X"FF",X"0B",X"C4",X"E1",X"08",X"84",X"40",X"08",X"86",X"40",X"18",X"F7",X"FF",X"3B",X"86",
		X"40",X"18",X"04",X"00",X"08",X"04",X"00",X"08",X"04",X"00",X"08",X"02",X"13",X"E0",X"03",X"F8",
		X"0F",X"FC",X"1F",X"7C",X"1F",X"3E",X"3E",X"1E",X"3C",X"1E",X"3C",X"3C",X"1E",X"F8",X"0F",X"F0",
		X"07",X"FC",X"1F",X"F8",X"0F",X"FD",X"5F",X"39",X"4E",X"11",X"44",X"FD",X"5F",X"11",X"44",X"01",
		X"40",X"01",X"40",X"02",X"0F",X"C0",X"01",X"F0",X"07",X"F8",X"0F",X"78",X"0F",X"3C",X"1E",X"38",
		X"0E",X"70",X"07",X"E0",X"03",X"F8",X"0F",X"F0",X"07",X"3A",X"2E",X"12",X"24",X"FB",X"6F",X"02",
		X"20",X"02",X"20",X"02",X"0B",X"20",X"00",X"F8",X"00",X"FC",X"01",X"DE",X"03",X"8E",X"03",X"DC",
		X"01",X"F8",X"00",X"DC",X"01",X"89",X"04",X"FD",X"05",X"01",X"04",X"03",X"20",X"04",X"00",X"00",
		X"19",X"02",X"00",X"7A",X"01",X"00",X"FC",X"00",X"00",X"7E",X"05",X"00",X"FE",X"03",X"80",X"FC",
		X"03",X"40",X"FE",X"07",X"68",X"F9",X"03",X"3E",X"F0",X"FF",X"0F",X"A0",X"FF",X"03",X"80",X"FF",
		X"00",X"80",X"FF",X"00",X"C0",X"FF",X"00",X"E0",X"FF",X"00",X"E0",X"FF",X"01",X"70",X"FF",X"03",
		X"30",X"FE",X"07",X"30",X"FC",X"0F",X"30",X"FE",X"0F",X"30",X"FE",X"0F",X"30",X"F8",X"0F",X"20",
		X"F0",X"07",X"00",X"F0",X"07",X"00",X"F0",X"07",X"00",X"C0",X"07",X"00",X"80",X"07",X"00",X"00",
		X"07",X"00",X"00",X"03",X"00",X"40",X"03",X"00",X"80",X"03",X"00",X"00",X"0F",X"02",X"19",X"14",
		X"00",X"34",X"00",X"3C",X"00",X"FF",X"00",X"3C",X"00",X"2E",X"00",X"7E",X"00",X"3C",X"40",X"18",
		X"30",X"F8",X"1F",X"FC",X"07",X"FE",X"01",X"FE",X"01",X"F7",X"01",X"E3",X"03",X"C3",X"07",X"E3",
		X"0F",X"E2",X"1F",X"82",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"0E",X"00",X"0C",X"00",X"0E",X"00",
		X"3C",X"02",X"13",X"14",X"00",X"34",X"00",X"3C",X"00",X"FF",X"00",X"2E",X"00",X"7E",X"00",X"38",
		X"10",X"18",X"0C",X"FC",X"07",X"7E",X"00",X"7A",X"00",X"F2",X"01",X"F2",X"01",X"E0",X"03",X"E0",
		X"03",X"C0",X"01",X"80",X"01",X"C0",X"01",X"80",X"07",X"04",X"0B",X"A0",X"00",X"00",X"00",X"B0",
		X"01",X"00",X"00",X"B0",X"01",X"3C",X"00",X"F0",X"01",X"7E",X"00",X"F9",X"13",X"FF",X"00",X"FF",
		X"9F",X"FF",X"81",X"F8",X"C7",X"FF",X"9F",X"FC",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"00",
		X"00",X"FC",X"41",X"00",X"00",X"00",X"20",X"04",X"09",X"80",X"02",X"00",X"00",X"C0",X"06",X"00",
		X"00",X"C0",X"07",X"1C",X"00",X"C8",X"27",X"3E",X"00",X"F8",X"3F",X"7F",X"10",X"E0",X"0F",X"FF",
		X"13",X"F0",X"FF",X"FF",X"1F",X"F0",X"FF",X"FF",X"1F",X"00",X"00",X"7E",X"08",X"03",X"08",X"14",
		X"00",X"00",X"34",X"00",X"00",X"3C",X"F0",X"00",X"FF",X"F8",X"41",X"3C",X"FC",X"4F",X"FE",X"FF",
		X"7F",X"FE",X"FF",X"7F",X"00",X"E0",X"23",X"03",X"08",X"A0",X"00",X"00",X"A0",X"01",X"00",X"E0",
		X"C1",X"01",X"F8",X"E7",X"43",X"E0",X"F1",X"4F",X"F0",X"FF",X"7F",X"F0",X"FF",X"7F",X"00",X"C0",
		X"23",X"02",X"07",X"0A",X"00",X"1A",X"00",X"1E",X"00",X"7F",X"8E",X"1E",X"9F",X"FF",X"FF",X"00",
		X"40",X"02",X"16",X"01",X"04",X"08",X"1E",X"3C",X"0F",X"F8",X"4F",X"FC",X"07",X"FE",X"07",X"7F",
		X"0F",X"FE",X"3F",X"FC",X"7F",X"F0",X"3F",X"F9",X"39",X"F8",X"7F",X"D0",X"3F",X"FC",X"0F",X"FC",
		X"47",X"FE",X"07",X"FF",X"0D",X"E4",X"1F",X"C2",X"3F",X"C9",X"77",X"80",X"03",X"80",X"21",X"06",
		X"24",X"30",X"00",X"00",X"00",X"00",X"0C",X"F0",X"01",X"00",X"00",X"80",X"0F",X"F0",X"1F",X"00",
		X"00",X"F8",X"0F",X"E0",X"FF",X"FF",X"FF",X"FF",X"07",X"E0",X"FF",X"FF",X"FF",X"FF",X"07",X"E0",
		X"FF",X"FF",X"FF",X"FF",X"07",X"C0",X"FF",X"FF",X"FF",X"FF",X"03",X"C0",X"FF",X"FF",X"FF",X"FF",
		X"03",X"C0",X"FF",X"FF",X"FF",X"FF",X"03",X"80",X"FF",X"FF",X"FF",X"FF",X"01",X"80",X"FF",X"FF",
		X"FF",X"FF",X"01",X"80",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"FF",X"FF",X"FF",X"FF",X"03",X"C0",X"FF",X"FF",
		X"FF",X"FF",X"03",X"C0",X"FF",X"FF",X"FF",X"FF",X"03",X"C0",X"FF",X"FF",X"FF",X"FF",X"03",X"00",
		X"7C",X"00",X"00",X"3E",X"00",X"00",X"93",X"01",X"80",X"C9",X"00",X"80",X"10",X"02",X"40",X"08",
		X"01",X"40",X"11",X"05",X"A0",X"88",X"02",X"40",X"92",X"04",X"20",X"49",X"02",X"20",X"54",X"08",
		X"10",X"2A",X"04",X"20",X"38",X"08",X"10",X"1C",X"04",X"F0",X"EF",X"1F",X"F8",X"F7",X"0F",X"20",
		X"38",X"08",X"10",X"1C",X"04",X"20",X"54",X"08",X"10",X"2A",X"04",X"40",X"92",X"04",X"20",X"49",
		X"02",X"40",X"11",X"05",X"A0",X"88",X"02",X"80",X"10",X"02",X"40",X"08",X"01",X"00",X"93",X"01",
		X"80",X"C9",X"00",X"00",X"7C",X"00",X"00",X"3E",X"00",X"01",X"0F",X"18",X"3C",X"7E",X"FF",X"E7",
		X"E7",X"81",X"81",X"E7",X"E7",X"E7",X"E7",X"E7",X"FF",X"FF",X"CD",X"F5",X"0E",X"11",X"0B",X"20",
		X"1A",X"EE",X"FF",X"12",X"C2",X"EC",X"0E",X"CD",X"40",X"10",X"CD",X"E6",X"0F",X"C3",X"EC",X"0E",
		X"3A",X"0B",X"20",X"A7",X"CA",X"DE",X"0E",X"CD",X"40",X"10",X"CD",X"A0",X"13",X"CD",X"B7",X"0F",
		X"CD",X"B0",X"14",X"CD",X"29",X"15",X"CD",X"63",X"10",X"22",X"52",X"20",X"CD",X"60",X"12",X"21",
		X"00",X"00",X"22",X"33",X"20",X"2A",X"52",X"20",X"CD",X"2D",X"11",X"C3",X"EC",X"0E",X"2A",X"52",
		X"20",X"E5",X"CD",X"D0",X"10",X"CD",X"09",X"11",X"E1",X"CD",X"7B",X"10",X"CD",X"98",X"16",X"E1",
		X"D1",X"C1",X"F1",X"FB",X"C9",X"21",X"02",X"20",X"7E",X"A7",X"CA",X"FF",X"0E",X"35",X"C9",X"23",
		X"7E",X"A7",X"CA",X"0C",X"0F",X"35",X"2B",X"3A",X"05",X"20",X"77",X"C9",X"23",X"7E",X"A7",X"CA",
		X"18",X"0F",X"35",X"3E",X"00",X"D3",X"05",X"C9",X"2A",X"00",X"20",X"7E",X"A7",X"C2",X"2C",X"0F",
		X"3E",X"00",X"D3",X"05",X"3A",X"0A",X"20",X"A7",X"C0",X"D3",X"03",X"C9",X"F2",X"3B",X"0F",X"E6",
		X"7F",X"32",X"05",X"20",X"23",X"22",X"00",X"20",X"C3",X"1B",X"0F",X"32",X"03",X"20",X"23",X"3A",
		X"05",X"20",X"3D",X"32",X"02",X"20",X"3E",X"01",X"32",X"04",X"20",X"7E",X"23",X"22",X"00",X"20",
		X"E6",X"7F",X"07",X"4F",X"06",X"00",X"21",X"50",X"1D",X"09",X"7E",X"D3",X"05",X"23",X"7E",X"D3",
		X"06",X"C9",X"31",X"00",X"24",X"CD",X"49",X"12",X"AF",X"06",X"13",X"11",X"00",X"20",X"12",X"13",
		X"05",X"C2",X"6E",X"0F",X"3D",X"12",X"13",X"12",X"21",X"91",X"1A",X"22",X"06",X"20",X"21",X"7E",
		X"0F",X"E5",X"FB",X"D3",X"04",X"2A",X"06",X"20",X"7E",X"A7",X"CA",X"9F",X"0F",X"23",X"22",X"06",
		X"20",X"EB",X"21",X"51",X"19",X"07",X"4F",X"06",X"00",X"09",X"7E",X"23",X"66",X"6F",X"E9",X"CD",
		X"F3",X"12",X"CD",X"1A",X"17",X"CD",X"F6",X"16",X"CD",X"EB",X"14",X"3A",X"0A",X"20",X"A7",X"C8",
		X"CD",X"5A",X"15",X"CD",X"DD",X"16",X"C9",X"21",X"86",X"20",X"11",X"0B",X"00",X"19",X"E5",X"CD",
		X"D8",X"0F",X"E1",X"01",X"EF",X"00",X"FE",X"70",X"D2",X"CD",X"0F",X"06",X"10",X"7E",X"A1",X"B0",
		X"77",X"7D",X"FE",X"B2",X"C2",X"BA",X"0F",X"C9",X"7E",X"A7",X"F0",X"23",X"7E",X"23",X"86",X"77",
		X"23",X"7E",X"23",X"86",X"77",X"C9",X"21",X"4B",X"20",X"7E",X"A7",X"C0",X"47",X"21",X"09",X"20",
		X"35",X"C2",X"14",X"10",X"36",X"1E",X"3A",X"45",X"20",X"A7",X"C2",X"0E",X"10",X"21",X"08",X"20");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
