library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity GALAXIAN_1H is
  port (
    CLK         : in    std_logic;
    ADDR        : in    std_logic_vector(10 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end entity;

architecture prom of GALAXIAN_1H is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
    x"38",x"7C",x"C2",x"82",x"86",x"7C",x"38",x"00", -- 0x0000
    x"02",x"02",x"FE",x"FE",x"42",x"02",x"00",x"00", -- 0x0008
    x"62",x"F2",x"BA",x"9A",x"9E",x"CE",x"46",x"00", -- 0x0010
    x"8C",x"DE",x"F2",x"B2",x"92",x"86",x"04",x"00", -- 0x0018
    x"08",x"FE",x"FE",x"C8",x"68",x"38",x"18",x"00", -- 0x0020
    x"1C",x"BE",x"A2",x"A2",x"A2",x"E6",x"E4",x"00", -- 0x0028
    x"0C",x"9E",x"92",x"92",x"D2",x"7E",x"3C",x"00", -- 0x0030
    x"C0",x"E0",x"B0",x"9E",x"8E",x"C0",x"C0",x"00", -- 0x0038
    x"0C",x"6E",x"9A",x"9A",x"B2",x"F2",x"6C",x"00", -- 0x0040
    x"78",x"FC",x"96",x"92",x"92",x"F2",x"60",x"00", -- 0x0048
    x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00", -- 0x0050
    x"00",x"00",x"00",x"00",x"08",x"58",x"F0",x"F0", -- 0x0058
    x"00",x"00",x"00",x"02",x"07",x"07",x"06",x"00", -- 0x0060
    x"06",x"1E",x"3E",x"1A",x"19",x"3F",x"3F",x"7D", -- 0x0068
    x"37",x"36",x"32",x"76",x"74",x"1E",x"06",x"00", -- 0x0070
    x"00",x"07",x"02",x"3E",x"3E",x"02",x"07",x"00", -- 0x0078
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0080
    x"3E",x"7E",x"C8",x"88",x"C8",x"7E",x"3E",x"00", -- 0x0088
    x"6C",x"FE",x"92",x"92",x"92",x"FE",x"FE",x"00", -- 0x0090
    x"44",x"C6",x"82",x"82",x"C6",x"7C",x"38",x"00", -- 0x0098
    x"38",x"7C",x"C6",x"82",x"82",x"FE",x"FE",x"00", -- 0x00A0
    x"82",x"92",x"92",x"92",x"FE",x"FE",x"00",x"00", -- 0x00A8
    x"80",x"90",x"90",x"90",x"90",x"FE",x"FE",x"00", -- 0x00B0
    x"9E",x"9E",x"92",x"82",x"C6",x"7C",x"38",x"00", -- 0x00B8
    x"FE",x"FE",x"10",x"10",x"10",x"FE",x"FE",x"00", -- 0x00C0
    x"82",x"82",x"FE",x"FE",x"82",x"82",x"00",x"00", -- 0x00C8
    x"FC",x"FE",x"02",x"02",x"02",x"06",x"04",x"00", -- 0x00D0
    x"82",x"C6",x"6E",x"3C",x"18",x"FE",x"FE",x"00", -- 0x00D8
    x"02",x"02",x"02",x"02",x"FE",x"FE",x"00",x"00", -- 0x00E0
    x"FE",x"FE",x"70",x"38",x"70",x"FE",x"FE",x"00", -- 0x00E8
    x"FE",x"FE",x"1C",x"38",x"70",x"FE",x"FE",x"00", -- 0x00F0
    x"7C",x"FE",x"82",x"82",x"82",x"FE",x"7C",x"00", -- 0x00F8
    x"70",x"F8",x"88",x"88",x"88",x"FE",x"FE",x"00", -- 0x0100
    x"7A",x"FC",x"8E",x"8A",x"82",x"FE",x"7C",x"00", -- 0x0108
    x"72",x"F6",x"9E",x"8C",x"88",x"FE",x"FE",x"00", -- 0x0110
    x"0C",x"5E",x"D2",x"92",x"92",x"F6",x"64",x"00", -- 0x0118
    x"80",x"80",x"FE",x"FE",x"80",x"80",x"00",x"00", -- 0x0120
    x"FC",x"FE",x"02",x"02",x"02",x"FE",x"FC",x"00", -- 0x0128
    x"F0",x"F8",x"1C",x"0E",x"1C",x"F8",x"F0",x"00", -- 0x0130
    x"F8",x"FE",x"1C",x"38",x"1C",x"FE",x"F8",x"00", -- 0x0138
    x"C6",x"EE",x"7C",x"38",x"7C",x"EE",x"C6",x"00", -- 0x0140
    x"C0",x"F0",x"1E",x"1E",x"F0",x"C0",x"00",x"00", -- 0x0148
    x"C2",x"E2",x"F2",x"BA",x"9E",x"8E",x"86",x"00", -- 0x0150
    x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00", -- 0x0158
    x"02",x"02",x"07",x"02",x"00",x"00",x"00",x"00", -- 0x0160
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0168
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0170
    x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0178
    x"0F",x"0F",x"0F",x"07",x"07",x"07",x"03",x"01", -- 0x0180
    x"30",x"20",x"00",x"00",x"00",x"00",x"00",x"1C", -- 0x0188
    x"70",x"78",x"7C",x"7E",x"7F",x"7E",x"7E",x"3C", -- 0x0190
    x"00",x"00",x"00",x"00",x"00",x"40",x"40",x"20", -- 0x0198
    x"03",x"03",x"01",x"01",x"01",x"01",x"01",x"00", -- 0x01A0
    x"03",x"03",x"03",x"07",x"07",x"03",x"03",x"03", -- 0x01A8
    x"02",x"01",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01B0
    x"F8",x"FE",x"7F",x"7C",x"3C",x"1C",x"0E",x"06", -- 0x01B8
    x"00",x"80",x"C0",x"E0",x"E0",x"E0",x"F0",x"F0", -- 0x01C0
    x"FF",x"7F",x"1F",x"0F",x"93",x"F8",x"F0",x"58", -- 0x01C8
    x"00",x"01",x"01",x"03",x"03",x"03",x"00",x"00", -- 0x01D0
    x"FC",x"F0",x"F8",x"F8",x"F8",x"FC",x"7D",x"1C", -- 0x01D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FB",x"F1",x"F8", -- 0x01E0
    x"FF",x"FF",x"FE",x"FC",x"FE",x"FE",x"FF",x"FF", -- 0x01E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"0F", -- 0x01F0
    x"00",x"00",x"00",x"00",x"08",x"3C",x"7E",x"FF", -- 0x01F8
    x"00",x"00",x"00",x"02",x"06",x"0F",x"10",x"0F", -- 0x0200
    x"06",x"0E",x"1E",x"38",x"78",x"88",x"08",x"88", -- 0x0208
    x"06",x"02",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0210
    x"78",x"38",x"1E",x"0E",x"06",x"00",x"00",x"00", -- 0x0218
    x"01",x"02",x"06",x"0E",x"02",x"02",x"02",x"02", -- 0x0220
    x"00",x"80",x"C0",x"E0",x"80",x"80",x"80",x"80", -- 0x0228
    x"06",x"04",x"0C",x"0C",x"1C",x"3F",x"38",x"38", -- 0x0230
    x"C0",x"40",x"60",x"60",x"70",x"F8",x"38",x"38", -- 0x0238
    x"F8",x"B0",x"90",x"D0",x"E8",x"E4",x"97",x"10", -- 0x0240
    x"00",x"00",x"00",x"00",x"00",x"00",x"F0",x"E0", -- 0x0248
    x"09",x"08",x"0A",x"0C",x"0C",x"0E",x"0C",x"08", -- 0x0250
    x"40",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0258
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0260
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0268
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0270
    x"01",x"03",x"66",x"9C",x"9C",x"66",x"03",x"01", -- 0x0278
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0280
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0288
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0290
    x"3F",x"83",x"86",x"BC",x"BC",x"86",x"83",x"3F", -- 0x0298
    x"01",x"02",x"05",x"0B",x"17",x"2C",x"5C",x"9F", -- 0x02A0
    x"80",x"40",x"A0",x"D0",x"E8",x"34",x"3A",x"F9", -- 0x02A8
    x"9F",x"5C",x"2C",x"17",x"0B",x"05",x"02",x"01", -- 0x02B0
    x"F9",x"3A",x"34",x"E8",x"D0",x"A0",x"40",x"80", -- 0x02B8
    x"01",x"21",x"70",x"20",x"03",x"03",x"0F",x"CF", -- 0x02C0
    x"80",x"84",x"0E",x"04",x"C0",x"C0",x"F0",x"F3", -- 0x02C8
    x"CF",x"0F",x"03",x"03",x"20",x"70",x"21",x"01", -- 0x02D0
    x"F3",x"F0",x"C0",x"C0",x"04",x"0E",x"84",x"80", -- 0x02D8
    x"00",x"3E",x"7E",x"7F",x"7E",x"7E",x"7E",x"7E", -- 0x02E0
    x"00",x"80",x"C0",x"E0",x"70",x"B8",x"DC",x"EE", -- 0x02E8
    x"7E",x"7C",x"7C",x"0C",x"3C",x"7C",x"7F",x"7F", -- 0x02F0
    x"F6",x"FF",x"FE",x"EF",x"D6",x"EE",x"DE",x"DE", -- 0x02F8
    x"00",x"00",x"00",x"C0",x"F0",x"F8",x"7E",x"1F", -- 0x0300
    x"00",x"00",x"00",x"03",x"0F",x"1F",x"7E",x"F8", -- 0x0308
    x"1F",x"7E",x"F8",x"F0",x"C0",x"00",x"00",x"00", -- 0x0310
    x"F8",x"7E",x"1F",x"0F",x"03",x"00",x"00",x"00", -- 0x0318
    x"07",x"03",x"03",x"01",x"00",x"00",x"00",x"00", -- 0x0320
    x"00",x"00",x"00",x"00",x"01",x"03",x"03",x"07", -- 0x0328
    x"00",x"3F",x"3F",x"1D",x"1D",x"0D",x"0F",x"07", -- 0x0330
    x"07",x"0F",x"0D",x"1D",x"1D",x"3F",x"3F",x"00", -- 0x0338
    x"E0",x"FC",x"FF",x"3F",x"07",x"00",x"00",x"00", -- 0x0340
    x"00",x"00",x"00",x"07",x"3F",x"FF",x"FC",x"E0", -- 0x0348
    x"03",x"1F",x"FF",x"FE",x"F0",x"E0",x"E0",x"E0", -- 0x0350
    x"E0",x"E0",x"E0",x"F0",x"FE",x"FF",x"1F",x"03", -- 0x0358
    x"E3",x"E1",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0", -- 0x0360
    x"E0",x"F0",x"F8",x"FC",x"FE",x"FF",x"EF",x"E7", -- 0x0368
    x"07",x"07",x"07",x"07",x"07",x"07",x"87",x"C7", -- 0x0370
    x"E7",x"F7",x"FF",x"7F",x"3F",x"1F",x"0F",x"07", -- 0x0378
    x"00",x"00",x"00",x"02",x"05",x"00",x"03",x"0C", -- 0x0380
    x"00",x"00",x"00",x"10",x"50",x"68",x"88",x"C8", -- 0x0388
    x"03",x"0A",x"03",x"01",x"04",x"03",x"00",x"00", -- 0x0390
    x"F4",x"A0",x"C0",x"70",x"40",x"20",x"00",x"00", -- 0x0398
    x"00",x"00",x"00",x"00",x"02",x"0A",x"04",x"00", -- 0x03A0
    x"00",x"00",x"00",x"00",x"50",x"A0",x"00",x"20", -- 0x03A8
    x"00",x"09",x"01",x"02",x"00",x"00",x"00",x"00", -- 0x03B0
    x"38",x"10",x"00",x"40",x"20",x"00",x"00",x"00", -- 0x03B8
    x"00",x"02",x"01",x"01",x"01",x"40",x"13",x"01", -- 0x03C0
    x"00",x"00",x"00",x"04",x"0C",x"18",x"80",x"90", -- 0x03C8
    x"00",x"08",x"00",x"00",x"02",x"04",x"00",x"00", -- 0x03D0
    x"82",x"CC",x"00",x"10",x"98",x"84",x"00",x"00", -- 0x03D8
    x"08",x"04",x"00",x"02",x"8C",x"0E",x"07",x"0F", -- 0x03E0
    x"01",x"12",x"00",x"04",x"00",x"C0",x"C8",x"E0", -- 0x03E8
    x"07",x"03",x"21",x"00",x"80",x"21",x"48",x"81", -- 0x03F0
    x"C2",x"80",x"01",x"00",x"22",x"00",x"02",x"01", -- 0x03F8
    x"FF",x"FF",x"FF",x"FF",x"7F",x"7F",x"3F",x"1E", -- 0x0400
    x"8F",x"CF",x"9F",x"BF",x"3F",x"FF",x"FF",x"FF", -- 0x0408
    x"E0",x"F8",x"FE",x"FF",x"FF",x"FF",x"FE",x"E0", -- 0x0410
    x"E0",x"E0",x"C0",x"C0",x"80",x"80",x"00",x"00", -- 0x0418
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FC",x"F0", -- 0x0420
    x"00",x"80",x"F8",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0428
    x"00",x"00",x"00",x"00",x"E0",x"80",x"00",x"00", -- 0x0430
    x"FC",x"F8",x"F8",x"F0",x"E0",x"00",x"00",x"00", -- 0x0438
    x"00",x"00",x"00",x"80",x"E0",x"F0",x"F8",x"FC", -- 0x0440
    x"0F",x"1F",x"3F",x"3F",x"7F",x"7F",x"FF",x"FF", -- 0x0448
    x"00",x"00",x"00",x"00",x"01",x"01",x"04",x"0E", -- 0x0450
    x"3F",x"9F",x"9F",x"CF",x"CF",x"CF",x"E7",x"E7", -- 0x0458
    x"00",x"03",x"1F",x"7F",x"FF",x"FF",x"FF",x"7F", -- 0x0460
    x"FC",x"FC",x"FE",x"FE",x"FE",x"FF",x"FF",x"FF", -- 0x0468
    x"00",x"38",x"AF",x"CB",x"E5",x"F2",x"F9",x"F9", -- 0x0470
    x"BE",x"BF",x"5F",x"5F",x"5F",x"2F",x"2F",x"2F", -- 0x0478
    x"00",x"00",x"00",x"C0",x"F0",x"F8",x"7C",x"7E", -- 0x0480
    x"00",x"00",x"80",x"80",x"C0",x"C0",x"C0",x"00", -- 0x0488
    x"01",x"01",x"01",x"03",x"03",x"03",x"07",x"07", -- 0x0490
    x"07",x"0F",x"0F",x"0F",x"1F",x"1F",x"1F",x"1F", -- 0x0498
    x"1F",x"3F",x"3F",x"7F",x"7F",x"7F",x"FF",x"FF", -- 0x04A0
    x"FF",x"FF",x"FE",x"FE",x"FE",x"FE",x"FC",x"FC", -- 0x04A8
    x"0F",x"0F",x"0F",x"1F",x"1F",x"3F",x"3F",x"7F", -- 0x04B0
    x"7F",x"7E",x"FE",x"FE",x"FE",x"FC",x"FC",x"FC", -- 0x04B8
    x"00",x"00",x"00",x"00",x"01",x"01",x"03",x"03", -- 0x04C0
    x"07",x"07",x"0F",x"0F",x"1F",x"1F",x"3F",x"3F", -- 0x04C8
    x"07",x"07",x"0F",x"0F",x"1F",x"3F",x"3F",x"7F", -- 0x04D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FE", -- 0x04D8
    x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC", -- 0x04E0
    x"FC",x"FC",x"3C",x"18",x"08",x"00",x"00",x"00", -- 0x04E8
    x"E0",x"C0",x"80",x"80",x"00",x"00",x"00",x"00", -- 0x04F0
    x"FE",x"FE",x"FC",x"FC",x"F0",x"F0",x"F0",x"F0", -- 0x04F8
    x"7F",x"7F",x"FF",x"FF",x"FF",x"FF",x"FE",x"FE", -- 0x0500
    x"FC",x"FC",x"FC",x"FC",x"FC",x"FE",x"FE",x"FE", -- 0x0508
    x"FF",x"FF",x"FF",x"FF",x"C3",x"01",x"01",x"00", -- 0x0510
    x"33",x"3F",x"1F",x"00",x"00",x"00",x"00",x"00", -- 0x0518
    x"C0",x"80",x"80",x"00",x"00",x"00",x"00",x"00", -- 0x0520
    x"C0",x"40",x"40",x"40",x"60",x"60",x"40",x"C0", -- 0x0528
    x"00",x"00",x"80",x"80",x"80",x"C0",x"C0",x"C0", -- 0x0530
    x"F8",x"F0",x"F0",x"E0",x"E0",x"C0",x"80",x"80", -- 0x0538
    x"FF",x"F8",x"E0",x"C0",x"80",x"00",x"00",x"00", -- 0x0540
    x"E0",x"E0",x"E0",x"E0",x"F0",x"F0",x"FE",x"FF", -- 0x0548
    x"F8",x"F8",x"F8",x"F0",x"F0",x"F0",x"F0",x"E0", -- 0x0550
    x"E0",x"E0",x"40",x"00",x"00",x"00",x"00",x"00", -- 0x0558
    x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF", -- 0x0560
    x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00", -- 0x0568
    x"F0",x"F8",x"FC",x"FE",x"1F",x"0F",x"07",x"07", -- 0x0570
    x"07",x"07",x"0F",x"1F",x"FE",x"FC",x"F8",x"F0", -- 0x0578
    x"E1",x"E1",x"E1",x"E1",x"FF",x"FF",x"FF",x"FF", -- 0x0580
    x"1E",x"3F",x"7F",x"FF",x"F3",x"E1",x"E1",x"E1", -- 0x0588
    x"07",x"0F",x"9F",x"FF",x"FC",x"F8",x"F0",x"E0", -- 0x0590
    x"C0",x"C0",x"C0",x"C0",x"FF",x"FF",x"FF",x"FF", -- 0x0598
    x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF", -- 0x05A0
    x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05A8
    x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"01",x"07", -- 0x05B0
    x"1F",x"7F",x"FE",x"F8",x"FF",x"FF",x"FF",x"FF", -- 0x05B8
    x"FF",x"FF",x"FF",x"FF",x"1F",x"7F",x"FE",x"F8", -- 0x05C0
    x"E0",x"80",x"00",x"00",x"FF",x"FF",x"FF",x"FF", -- 0x05C8
    x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"FF", -- 0x05D0
    x"FF",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0", -- 0x05D8
    x"38",x"78",x"F8",x"F8",x"F0",x"E0",x"E0",x"E0", -- 0x05E0
    x"E0",x"E0",x"E0",x"F0",x"FF",x"FF",x"7F",x"3F", -- 0x05E8
    x"1C",x"1E",x"1F",x"1F",x"0F",x"07",x"07",x"07", -- 0x05F0
    x"07",x"07",x"07",x"0F",x"FF",x"FF",x"FE",x"FC", -- 0x05F8
    x"80",x"C0",x"E0",x"F0",x"F8",x"7C",x"3E",x"1F", -- 0x0600
    x"0F",x"07",x"03",x"03",x"FF",x"FF",x"FF",x"FF", -- 0x0608
    x"01",x"03",x"07",x"0F",x"1F",x"3E",x"7C",x"F8", -- 0x0610
    x"F0",x"E0",x"C0",x"C0",x"FF",x"FF",x"FF",x"FF", -- 0x0618
    x"00",x"00",x"00",x"00",x"81",x"87",x"00",x"00", -- 0x0620
    x"00",x"00",x"00",x"00",x"80",x"80",x"C0",x"00", -- 0x0628
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0630
    x"10",x"10",x"30",x"30",x"30",x"60",x"40",x"C0", -- 0x0638
    x"03",x"0F",x"1F",x"1B",x"39",x"70",x"73",x"37", -- 0x0640
    x"C0",x"C0",x"E8",x"FC",x"FC",x"9C",x"9C",x"EE", -- 0x0648
    x"3F",x"1F",x"07",x"1F",x"1E",x"0F",x"0F",x"01", -- 0x0650
    x"DE",x"DF",x"9F",x"A7",x"47",x"AF",x"FC",x"E0", -- 0x0658
    x"7F",x"7E",x"7E",x"7F",x"7F",x"7F",x"7E",x"78", -- 0x0660
    x"FE",x"EE",x"EE",x"F8",x"E0",x"80",x"00",x"00", -- 0x0668
    x"62",x"0E",x"3E",x"7E",x"7A",x"73",x"6B",x"59", -- 0x0670
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0678
    x"00",x"80",x"40",x"20",x"10",x"08",x"04",x"02", -- 0x0680
    x"00",x"10",x"08",x"08",x"1C",x"0C",x"00",x"00", -- 0x0688
    x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0690
    x"E0",x"E0",x"70",x"06",x"02",x"00",x"60",x"20", -- 0x0698
    x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"02", -- 0x06A0
    x"00",x"04",x"08",x"18",x"30",x"20",x"E0",x"40", -- 0x06A8
    x"00",x"00",x"71",x"12",x"11",x"16",x"04",x"04", -- 0x06B0
    x"00",x"00",x"80",x"00",x"00",x"00",x"00",x"70", -- 0x06B8
    x"31",x"08",x"00",x"00",x"00",x"00",x"01",x"01", -- 0x06C0
    x"C0",x"00",x"00",x"00",x"40",x"C0",x"78",x"00", -- 0x06C8
    x"01",x"06",x"0C",x"08",x"08",x"10",x"20",x"00", -- 0x06D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06D8
    x"00",x"00",x"00",x"00",x"00",x"0A",x"0F",x"03", -- 0x06E0
    x"38",x"1E",x"00",x"00",x"00",x"00",x"00",x"80", -- 0x06E8
    x"03",x"01",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06F0
    x"B0",x"30",x"30",x"1C",x"0C",x"04",x"02",x"00", -- 0x06F8
    x"00",x"80",x"40",x"30",x"08",x"05",x"07",x"03", -- 0x0700
    x"80",x"40",x"20",x"10",x"6C",x"90",x"0E",x"21", -- 0x0708
    x"01",x"01",x"03",x"06",x"04",x"04",x"1B",x"3A", -- 0x0710
    x"48",x"38",x"0E",x"1F",x"0F",x"07",x"01",x"D9", -- 0x0718
    x"00",x"00",x"00",x"00",x"00",x"06",x"04",x"09", -- 0x0720
    x"01",x"02",x"06",x"0C",x"38",x"70",x"58",x"AC", -- 0x0728
    x"D3",x"C6",x"87",x"6B",x"F4",x"A4",x"08",x"CC", -- 0x0730
    x"C8",x"D0",x"10",x"40",x"80",x"80",x"00",x"CF", -- 0x0738
    x"C5",x"02",x"00",x"06",x"02",x"01",x"00",x"02", -- 0x0740
    x"3F",x"8F",x"07",x"02",x"08",x"15",x"C7",x"F5", -- 0x0748
    x"02",x"06",x"0C",x"18",x"30",x"20",x"40",x"00", -- 0x0750
    x"74",x"22",x"01",x"00",x"02",x"04",x"08",x"10", -- 0x0758
    x"EF",x"EE",x"79",x"28",x"84",x"91",x"0B",x"15", -- 0x0760
    x"98",x"30",x"20",x"20",x"C0",x"00",x"40",x"F8", -- 0x0768
    x"94",x"C4",x"28",x"D0",x"30",x"00",x"00",x"00", -- 0x0770
    x"70",x"08",x"04",x"02",x"01",x"00",x"00",x"00", -- 0x0778
    x"00",x"80",x"60",x"10",x"0C",x"07",x"03",x"01", -- 0x0780
    x"20",x"20",x"10",x"10",x"08",x"9C",x"FF",x"FF", -- 0x0788
    x"10",x"0D",x"03",x"01",x"00",x"03",x"07",x"FF", -- 0x0790
    x"FF",x"FF",x"FB",x"FB",x"F7",x"E1",x"F0",x"E0", -- 0x0798
    x"00",x"00",x"40",x"41",x"42",x"46",x"DC",x"FD", -- 0x07A0
    x"00",x"02",x"04",x"18",x"20",x"60",x"C0",x"80", -- 0x07A8
    x"FF",x"FF",x"FF",x"FF",x"C7",x"03",x"07",x"00", -- 0x07B0
    x"80",x"04",x"18",x"20",x"C0",x"80",x"E0",x"FF", -- 0x07B8
    x"01",x"00",x"00",x"01",x"03",x"0F",x"18",x"60", -- 0x07C0
    x"80",x"F0",x"F0",x"F8",x"FC",x"7D",x"7F",x"FF", -- 0x07C8
    x"01",x"03",x"04",x"08",x"10",x"20",x"40",x"00", -- 0x07D0
    x"E7",x"83",x"01",x"01",x"00",x"00",x"00",x"00", -- 0x07D8
    x"0F",x"00",x"00",x"0B",x"0E",x"07",x"FF",x"FB", -- 0x07E0
    x"C0",x"00",x"40",x"C0",x"38",x"0C",x"80",x"80", -- 0x07E8
    x"F8",x"F8",x"DC",x"8C",x"86",x"82",x"82",x"80", -- 0x07F0
    x"C0",x"60",x"20",x"10",x"08",x"04",x"00",x"00"  -- 0x07F8
  );

begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
