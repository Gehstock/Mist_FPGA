library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity rom1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of rom1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"C3",X"18",X"00",X"00",X"00",X"E5",X"D5",X"C5",X"F5",X"C3",X"E8",X"0C",X"00",
		X"E5",X"D5",X"C5",X"F5",X"C3",X"B3",X"13",X"00",X"31",X"00",X"24",X"11",X"B0",X"03",X"CD",X"F2",
		X"04",X"21",X"43",X"23",X"36",X"01",X"11",X"40",X"22",X"21",X"7C",X"46",X"06",X"19",X"CD",X"41",
		X"0B",X"CD",X"D6",X"45",X"21",X"01",X"50",X"22",X"3F",X"23",X"DB",X"02",X"E6",X"04",X"C2",X"5A",
		X"47",X"CD",X"E8",X"45",X"CD",X"8C",X"04",X"C3",X"00",X"40",X"CD",X"EB",X"45",X"CD",X"2A",X"04",
		X"CD",X"DB",X"18",X"FE",X"03",X"CA",X"0E",X"46",X"FE",X"04",X"DA",X"E3",X"01",X"21",X"1C",X"21",
		X"36",X"FF",X"F5",X"21",X"00",X"07",X"11",X"04",X"22",X"06",X"0D",X"CD",X"41",X"0B",X"F1",X"FE",
		X"06",X"DA",X"7D",X"00",X"21",X"58",X"2A",X"22",X"06",X"22",X"22",X"08",X"22",X"FE",X"05",X"DA",
		X"85",X"00",X"CD",X"72",X"02",X"21",X"3C",X"20",X"36",X"06",X"CD",X"79",X"04",X"D3",X"06",X"21",
		X"1E",X"25",X"DA",X"98",X"00",X"21",X"1E",X"38",X"01",X"38",X"01",X"CD",X"DB",X"04",X"06",X"60",
		X"CD",X"81",X"04",X"11",X"DF",X"1C",X"21",X"1E",X"38",X"CD",X"79",X"04",X"D2",X"B5",X"00",X"11",
		X"CC",X"1C",X"21",X"1E",X"25",X"06",X"07",X"CD",X"22",X"08",X"06",X"60",X"CD",X"81",X"04",X"21",
		X"3C",X"20",X"35",X"C2",X"8A",X"00",X"21",X"42",X"23",X"36",X"FF",X"CD",X"AA",X"0C",X"CD",X"9F",
		X"0C",X"3E",X"02",X"CD",X"7E",X"06",X"3E",X"FF",X"CD",X"A0",X"06",X"3E",X"10",X"CD",X"95",X"06",
		X"21",X"3D",X"20",X"7E",X"A7",X"D3",X"06",X"C2",X"8B",X"05",X"3A",X"6F",X"20",X"A7",X"21",X"03",
		X"03",X"22",X"0C",X"20",X"CA",X"13",X"01",X"21",X"0A",X"21",X"7E",X"E6",X"40",X"CA",X"05",X"01",
		X"21",X"0C",X"20",X"36",X"05",X"21",X"0A",X"22",X"7E",X"E6",X"40",X"CA",X"13",X"01",X"21",X"0D",
		X"20",X"36",X"05",X"C3",X"5D",X"47",X"FE",X"5D",X"DA",X"3A",X"01",X"21",X"6F",X"20",X"36",X"00",
		X"3E",X"10",X"CD",X"89",X"06",X"3A",X"1D",X"20",X"FE",X"6D",X"D2",X"7C",X"02",X"FE",X"66",X"D2",
		X"8C",X"02",X"C3",X"6D",X"47",X"3E",X"08",X"CD",X"92",X"02",X"CD",X"37",X"02",X"21",X"1C",X"20",
		X"7E",X"A7",X"CA",X"61",X"01",X"36",X"00",X"2E",X"20",X"36",X"01",X"CD",X"79",X"04",X"21",X"33",
		X"23",X"DA",X"55",X"01",X"23",X"7E",X"32",X"02",X"23",X"CD",X"31",X"08",X"3E",X"01",X"CD",X"95",
		X"06",X"D3",X"06",X"CD",X"DB",X"18",X"FE",X"08",X"DA",X"7E",X"01",X"FE",X"0A",X"21",X"47",X"20",
		X"7E",X"D2",X"79",X"01",X"FE",X"02",X"C3",X"8E",X"01",X"FE",X"01",X"C3",X"8E",X"01",X"FE",X"06",
		X"21",X"47",X"20",X"7E",X"DA",X"8C",X"01",X"FE",X"03",X"C3",X"8E",X"01",X"FE",X"08",X"DA",X"AA",
		X"01",X"36",X"00",X"23",X"34",X"CD",X"53",X"05",X"06",X"02",X"AF",X"2A",X"14",X"20",X"11",X"E0",
		X"FF",X"77",X"19",X"22",X"14",X"20",X"05",X"C2",X"A1",X"01",X"CD",X"79",X"04",X"21",X"03",X"23",
		X"D2",X"CC",X"01",X"7E",X"FE",X"01",X"DA",X"E0",X"00",X"21",X"45",X"23",X"7E",X"A7",X"C2",X"E0",
		X"00",X"36",X"FF",X"2E",X"2F",X"34",X"CD",X"2A",X"04",X"C3",X"E0",X"00",X"2E",X"06",X"7E",X"FE",
		X"01",X"DA",X"E0",X"00",X"21",X"46",X"23",X"7E",X"A7",X"C2",X"E0",X"00",X"36",X"FF",X"2E",X"30",
		X"C3",X"C5",X"01",X"FE",X"02",X"DA",X"85",X"00",X"F5",X"21",X"1D",X"21",X"36",X"FF",X"21",X"B0",
		X"46",X"11",X"20",X"21",X"06",X"80",X"CD",X"41",X"0B",X"21",X"00",X"47",X"CD",X"22",X"04",X"21",
		X"10",X"01",X"22",X"1E",X"21",X"F1",X"FE",X"03",X"DA",X"85",X"00",X"CD",X"72",X"02",X"21",X"20",
		X"21",X"3E",X"04",X"77",X"2E",X"4E",X"77",X"2E",X"6C",X"77",X"2E",X"44",X"36",X"FC",X"2E",X"48",
		X"36",X"FC",X"C3",X"85",X"00",X"E5",X"06",X"08",X"C5",X"1A",X"77",X"13",X"01",X"20",X"00",X"09",
		X"C1",X"05",X"C2",X"28",X"02",X"E1",X"C9",X"21",X"02",X"20",X"7E",X"A7",X"CA",X"53",X"02",X"3A",
		X"04",X"20",X"21",X"0F",X"1C",X"3D",X"CA",X"50",X"02",X"11",X"16",X"00",X"19",X"C3",X"45",X"02",
		X"22",X"10",X"20",X"3A",X"02",X"21",X"A7",X"CA",X"63",X"02",X"3A",X"04",X"21",X"CD",X"F0",X"1A",
		X"22",X"0D",X"21",X"3A",X"02",X"22",X"A7",X"C8",X"3A",X"04",X"22",X"CD",X"F0",X"1A",X"22",X"0D",
		X"22",X"C9",X"21",X"6F",X"20",X"36",X"FF",X"3E",X"10",X"C3",X"7E",X"06",X"FE",X"7B",X"D2",X"9F",
		X"02",X"21",X"06",X"06",X"3E",X"04",X"CD",X"92",X"02",X"C3",X"3A",X"01",X"21",X"05",X"05",X"C3",
		X"84",X"02",X"22",X"0C",X"20",X"F5",X"3E",X"1C",X"CD",X"A0",X"06",X"F1",X"C3",X"95",X"06",X"3A",
		X"1C",X"20",X"A7",X"C2",X"81",X"02",X"21",X"42",X"23",X"36",X"00",X"3E",X"FF",X"CD",X"A0",X"06",
		X"CD",X"79",X"04",X"21",X"31",X"23",X"DA",X"BA",X"02",X"23",X"34",X"21",X"0D",X"25",X"01",X"03",
		X"D0",X"CD",X"DE",X"41",X"21",X"0D",X"C5",X"01",X"33",X"03",X"3E",X"01",X"CD",X"D2",X"08",X"21",
		X"0E",X"2B",X"11",X"15",X"47",X"06",X"0F",X"CD",X"22",X"08",X"CD",X"DB",X"42",X"CD",X"FD",X"05",
		X"CD",X"AA",X"41",X"CD",X"4C",X"04",X"21",X"01",X"00",X"22",X"6A",X"20",X"21",X"00",X"3B",X"06",
		X"0E",X"CD",X"CD",X"03",X"21",X"00",X"FF",X"22",X"6A",X"20",X"21",X"0E",X"3B",X"06",X"0B",X"CD",
		X"CD",X"03",X"21",X"6C",X"20",X"36",X"FF",X"21",X"FF",X"FF",X"22",X"6A",X"20",X"CD",X"79",X"04",
		X"21",X"1D",X"26",X"DA",X"19",X"03",X"21",X"1D",X"39",X"06",X"0E",X"CD",X"CD",X"03",X"CD",X"79",
		X"04",X"21",X"00",X"01",X"22",X"6A",X"20",X"06",X"09",X"21",X"0F",X"26",X"DA",X"3A",X"03",X"21",
		X"00",X"FF",X"22",X"6A",X"20",X"06",X"0A",X"21",X"0F",X"39",X"CD",X"CD",X"03",X"21",X"0E",X"2E",
		X"11",X"24",X"47",X"CD",X"25",X"02",X"21",X"0D",X"2E",X"01",X"30",X"01",X"3E",X"38",X"CD",X"DC",
		X"04",X"2A",X"12",X"20",X"22",X"01",X"23",X"CD",X"5E",X"04",X"3E",X"20",X"CD",X"9C",X"41",X"21",
		X"0C",X"2F",X"CD",X"79",X"04",X"11",X"03",X"23",X"DA",X"6E",X"03",X"11",X"06",X"23",X"CD",X"80",
		X"0C",X"CD",X"9A",X"41",X"CD",X"4C",X"04",X"CD",X"34",X"0C",X"CD",X"79",X"04",X"21",X"33",X"23",
		X"DA",X"84",X"03",X"23",X"22",X"6E",X"20",X"7E",X"C6",X"10",X"FE",X"A0",X"DA",X"91",X"03",X"3E",
		X"90",X"77",X"21",X"0F",X"2C",X"11",X"38",X"47",X"06",X"0D",X"CD",X"22",X"08",X"21",X"0F",X"31",
		X"22",X"28",X"23",X"2A",X"6E",X"20",X"22",X"26",X"23",X"06",X"01",X"CD",X"52",X"08",X"CD",X"9A",
		X"41",X"21",X"0B",X"CE",X"01",X"16",X"01",X"3E",X"01",X"CD",X"D2",X"08",X"21",X"0B",X"2F",X"11",
		X"45",X"47",X"06",X"09",X"CD",X"22",X"08",X"CD",X"AA",X"41",X"C3",X"4A",X"00",X"C5",X"E5",X"CD",
		X"F0",X"03",X"2A",X"6A",X"20",X"EB",X"E1",X"19",X"3A",X"6C",X"20",X"A7",X"C2",X"F6",X"03",X"11",
		X"12",X"20",X"CD",X"08",X"04",X"06",X"20",X"CD",X"81",X"04",X"C1",X"05",X"C2",X"CD",X"03",X"C9",
		X"01",X"01",X"28",X"C3",X"DE",X"41",X"CD",X"79",X"04",X"11",X"03",X"23",X"DA",X"02",X"04",X"11",
		X"06",X"23",X"CD",X"11",X"04",X"C3",X"E5",X"03",X"E5",X"CD",X"1A",X"04",X"CD",X"50",X"08",X"E1",
		X"C9",X"E5",X"CD",X"1A",X"04",X"CD",X"43",X"08",X"E1",X"C9",X"22",X"28",X"23",X"EB",X"22",X"26",
		X"23",X"C9",X"11",X"06",X"22",X"06",X"0E",X"C3",X"41",X"0B",X"21",X"2F",X"23",X"CD",X"79",X"04",
		X"DA",X"35",X"04",X"2E",X"30",X"7E",X"FE",X"02",X"D8",X"21",X"00",X"25",X"F5",X"11",X"4E",X"47",
		X"CD",X"25",X"02",X"F1",X"3D",X"FE",X"02",X"D8",X"24",X"C3",X"3C",X"04",X"21",X"01",X"24",X"01",
		X"1C",X"E0",X"CD",X"DE",X"41",X"21",X"01",X"C4",X"01",X"38",X"1B",X"C3",X"D0",X"08",X"21",X"02",
		X"23",X"11",X"05",X"23",X"3A",X"2A",X"23",X"5F",X"CD",X"81",X"08",X"13",X"23",X"CD",X"8F",X"08",
		X"21",X"00",X"23",X"11",X"03",X"00",X"C3",X"CA",X"0A",X"AF",X"3A",X"2C",X"23",X"A7",X"C0",X"37",
		X"C9",X"0E",X"FF",X"0D",X"C2",X"83",X"04",X"05",X"C2",X"81",X"04",X"C9",X"21",X"C9",X"04",X"11",
		X"2F",X"23",X"06",X"0C",X"CD",X"41",X"0B",X"DB",X"02",X"E6",X"03",X"06",X"03",X"80",X"21",X"2F",
		X"23",X"77",X"23",X"77",X"DB",X"02",X"E6",X"08",X"C8",X"21",X"04",X"23",X"36",X"90",X"2E",X"07",
		X"36",X"90",X"C3",X"BC",X"47",X"04",X"22",X"31",X"23",X"C9",X"05",X"23",X"1D",X"26",X"21",X"BA",
		X"04",X"11",X"26",X"23",X"06",X"04",X"C3",X"41",X"0B",X"05",X"05",X"01",X"01",X"10",X"10",X"00",
		X"40",X"00",X"40",X"D0",X"90",X"21",X"00",X"24",X"01",X"E0",X"20",X"AF",X"C5",X"E5",X"77",X"23",
		X"05",X"C2",X"DE",X"04",X"E1",X"11",X"20",X"00",X"19",X"C1",X"0D",X"C2",X"DC",X"04",X"C9",X"11",
		X"3F",X"02",X"21",X"00",X"20",X"C3",X"CA",X"0A",X"CD",X"EF",X"04",X"11",X"04",X"20",X"21",X"B3",
		X"1B",X"06",X"14",X"CD",X"41",X"0B",X"11",X"04",X"21",X"21",X"C6",X"1B",X"06",X"17",X"CD",X"41",
		X"0B",X"11",X"20",X"23",X"21",X"E7",X"1B",X"06",X"0A",X"CD",X"41",X"0B",X"21",X"72",X"20",X"22",
		X"70",X"20",X"21",X"2D",X"05",X"11",X"72",X"20",X"06",X"1B",X"C3",X"41",X"0B",X"03",X"01",X"07",
		X"01",X"07",X"05",X"07",X"01",X"03",X"05",X"07",X"01",X"03",X"01",X"07",X"05",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"0E",X"07",X"11",X"2A",X"23",X"06",X"03",
		X"C3",X"41",X"0B",X"21",X"12",X"20",X"7E",X"A7",X"C8",X"23",X"EB",X"21",X"0E",X"1C",X"0E",X"02",
		X"37",X"3E",X"99",X"CE",X"00",X"96",X"EB",X"86",X"27",X"77",X"EB",X"1B",X"2B",X"0D",X"C2",X"61",
		X"05",X"21",X"00",X"3B",X"22",X"28",X"23",X"21",X"12",X"20",X"22",X"26",X"23",X"06",X"02",X"CD",
		X"50",X"08",X"C3",X"BE",X"04",X"21",X"0B",X"07",X"C3",X"4B",X"05",X"CD",X"02",X"06",X"CD",X"B0",
		X"40",X"CD",X"FD",X"05",X"CD",X"95",X"02",X"3A",X"3B",X"23",X"A7",X"CA",X"07",X"06",X"CD",X"79",
		X"04",X"21",X"2F",X"23",X"D2",X"D0",X"05",X"7E",X"3D",X"77",X"C2",X"C7",X"05",X"CD",X"48",X"06",
		X"CD",X"11",X"07",X"CD",X"9A",X"41",X"21",X"30",X"23",X"7E",X"A7",X"CA",X"19",X"06",X"CD",X"08",
		X"46",X"CD",X"AC",X"06",X"C3",X"4A",X"00",X"23",X"7E",X"A7",X"CA",X"4A",X"00",X"C3",X"BE",X"05",
		X"23",X"7E",X"3D",X"77",X"C2",X"F4",X"05",X"CD",X"4E",X"06",X"CD",X"11",X"07",X"CD",X"9A",X"41",
		X"21",X"2F",X"23",X"7E",X"A7",X"CA",X"19",X"06",X"CD",X"9A",X"41",X"CD",X"D5",X"04",X"CD",X"C0",
		X"06",X"C3",X"4A",X"00",X"2B",X"7E",X"A7",X"CA",X"4A",X"00",X"C3",X"E8",X"05",X"3E",X"12",X"CD",
		X"89",X"06",X"3E",X"FF",X"C3",X"A0",X"06",X"21",X"2F",X"23",X"7E",X"3D",X"77",X"CA",X"16",X"06",
		X"CD",X"9A",X"41",X"C3",X"4A",X"00",X"CD",X"11",X"07",X"3E",X"02",X"CD",X"89",X"06",X"CD",X"9A",
		X"41",X"CD",X"4C",X"04",X"CD",X"8C",X"04",X"21",X"10",X"2D",X"CD",X"70",X"06",X"CD",X"9A",X"41",
		X"3A",X"0E",X"23",X"A7",X"C4",X"48",X"43",X"CD",X"D6",X"45",X"21",X"43",X"23",X"36",X"FF",X"21",
		X"00",X"00",X"22",X"45",X"23",X"C3",X"41",X"00",X"11",X"E3",X"06",X"C3",X"51",X"06",X"11",X"F6",
		X"06",X"D5",X"21",X"06",X"CD",X"01",X"14",X"01",X"CD",X"D0",X"08",X"21",X"03",X"CD",X"01",X"14",
		X"01",X"CD",X"D0",X"08",X"D1",X"21",X"06",X"2D",X"06",X"0A",X"CD",X"7B",X"41",X"21",X"03",X"2D",
		X"11",X"ED",X"06",X"06",X"09",X"C3",X"7B",X"41",X"21",X"10",X"2D",X"C3",X"70",X"06",X"C5",X"21",
		X"2D",X"23",X"46",X"B0",X"D3",X"05",X"77",X"C1",X"C9",X"C5",X"21",X"2D",X"23",X"46",X"2F",X"A0",
		X"D3",X"05",X"77",X"C1",X"C9",X"C5",X"21",X"2E",X"23",X"46",X"B0",X"D3",X"03",X"77",X"C1",X"C9",
		X"C5",X"21",X"2E",X"23",X"46",X"2F",X"A0",X"D3",X"03",X"77",X"C1",X"C9",X"21",X"0B",X"07",X"CD",
		X"CE",X"45",X"F3",X"3E",X"20",X"21",X"2D",X"23",X"46",X"B0",X"D3",X"05",X"77",X"C3",X"D5",X"06",
		X"CD",X"CB",X"45",X"F3",X"CD",X"DC",X"0E",X"D2",X"E1",X"06",X"3E",X"20",X"21",X"2D",X"23",X"46",
		X"2F",X"A0",X"D3",X"05",X"77",X"06",X"F0",X"0E",X"FF",X"0D",X"C2",X"D9",X"06",X"05",X"C2",X"D7",
		X"06",X"FB",X"C9",X"0F",X"0B",X"00",X"18",X"04",X"11",X"1B",X"1E",X"21",X"1F",X"06",X"00",X"0C",
		X"04",X"1B",X"0E",X"15",X"04",X"11",X"0F",X"0B",X"00",X"18",X"04",X"11",X"1B",X"1E",X"22",X"1F",
		X"05",X"05",X"B8",X"42",X"B8",X"42",X"48",X"9E",X"0A",X"9E",X"0A",X"08",X"39",X"FF",X"05",X"26",
		X"00",X"21",X"03",X"23",X"3A",X"2A",X"23",X"6F",X"2B",X"2B",X"22",X"09",X"23",X"06",X"03",X"11",
		X"3F",X"23",X"AF",X"1A",X"BE",X"DA",X"31",X"07",X"96",X"C0",X"23",X"13",X"05",X"C2",X"23",X"07",
		X"C9",X"06",X"03",X"2A",X"09",X"23",X"11",X"3F",X"23",X"7E",X"12",X"23",X"13",X"05",X"C2",X"39",
		X"07",X"CD",X"79",X"04",X"21",X"FF",X"00",X"DA",X"4D",X"07",X"21",X"FF",X"FF",X"22",X"0E",X"23",
		X"21",X"1D",X"2F",X"22",X"28",X"23",X"2A",X"09",X"23",X"22",X"26",X"23",X"C3",X"43",X"08",X"0F",
		X"0F",X"D2",X"93",X"07",X"CD",X"27",X"0B",X"7D",X"E6",X"1F",X"FE",X"0E",X"CA",X"7F",X"07",X"D6",
		X"02",X"21",X"B4",X"12",X"CA",X"7D",X"07",X"23",X"D6",X"03",X"C2",X"77",X"07",X"7E",X"C9",X"7C",
		X"FE",X"37",X"D2",X"8D",X"07",X"FE",X"2E",X"D2",X"90",X"07",X"3E",X"10",X"C9",X"3E",X"12",X"C9",
		X"3E",X"11",X"C9",X"CD",X"27",X"0B",X"7C",X"D6",X"25",X"21",X"BD",X"12",X"C3",X"74",X"07",X"21",
		X"8B",X"09",X"3E",X"18",X"CD",X"F2",X"07",X"21",X"B4",X"09",X"3E",X"FF",X"CD",X"F2",X"07",X"01",
		X"11",X"0A",X"21",X"F5",X"09",X"CD",X"DC",X"07",X"01",X"19",X"0A",X"21",X"FC",X"09",X"CD",X"DC",
		X"07",X"01",X"21",X"0A",X"21",X"03",X"0A",X"CD",X"DC",X"07",X"01",X"29",X"0A",X"21",X"0A",X"0A",
		X"CD",X"DC",X"07",X"01",X"6A",X"0A",X"21",X"31",X"0A",X"C3",X"DC",X"07",X"E5",X"7E",X"FE",X"FF",
		X"C2",X"E5",X"07",X"E1",X"C9",X"5F",X"23",X"56",X"EB",X"CD",X"10",X"08",X"E1",X"23",X"23",X"C3",
		X"DC",X"07",X"E5",X"47",X"7E",X"FE",X"FF",X"C2",X"FC",X"07",X"E1",X"C9",X"78",X"46",X"23",X"4E",
		X"23",X"5E",X"23",X"56",X"EB",X"CD",X"DC",X"04",X"E1",X"23",X"23",X"23",X"23",X"C3",X"F2",X"07",
		X"C5",X"16",X"08",X"D5",X"0A",X"77",X"11",X"20",X"00",X"19",X"03",X"D1",X"15",X"C2",X"13",X"08",
		X"C1",X"C9",X"D5",X"1A",X"CD",X"94",X"08",X"CD",X"AB",X"08",X"D1",X"13",X"05",X"C2",X"22",X"08",
		X"C9",X"CD",X"5E",X"04",X"21",X"2A",X"23",X"7E",X"3D",X"3D",X"2E",X"26",X"77",X"2E",X"2B",X"7E",
		X"2E",X"29",X"77",X"2A",X"26",X"23",X"7E",X"23",X"22",X"26",X"23",X"E6",X"0F",X"CD",X"71",X"08",
		X"06",X"02",X"C5",X"2A",X"26",X"23",X"7E",X"F5",X"E6",X"F0",X"0F",X"0F",X"0F",X"0F",X"CD",X"71",
		X"08",X"F1",X"E6",X"0F",X"CD",X"71",X"08",X"21",X"26",X"23",X"34",X"C1",X"05",X"C2",X"52",X"08",
		X"C9",X"C6",X"20",X"CD",X"94",X"08",X"2A",X"28",X"23",X"CD",X"AB",X"08",X"21",X"29",X"23",X"34",
		X"C9",X"06",X"03",X"AF",X"1A",X"8E",X"27",X"77",X"2B",X"1B",X"05",X"C2",X"84",X"08",X"C9",X"06",
		X"03",X"C3",X"41",X"0B",X"11",X"5C",X"1D",X"A7",X"C8",X"E5",X"21",X"00",X"00",X"C5",X"01",X"05",
		X"00",X"09",X"3D",X"C2",X"9E",X"08",X"19",X"EB",X"C1",X"E1",X"C9",X"C5",X"06",X"05",X"D3",X"06",
		X"C5",X"1A",X"07",X"77",X"13",X"01",X"20",X"00",X"09",X"C1",X"05",X"C2",X"AE",X"08",X"AF",X"77",
		X"01",X"20",X"00",X"09",X"77",X"09",X"77",X"09",X"C1",X"C9",X"21",X"00",X"C4",X"01",X"38",X"20",
		X"3E",X"FF",X"C5",X"E5",X"77",X"23",X"05",X"C2",X"D4",X"08",X"E1",X"11",X"80",X"00",X"19",X"C1",
		X"0D",X"C2",X"D2",X"08",X"C9",X"E5",X"7E",X"FE",X"FF",X"C2",X"EE",X"08",X"E1",X"C9",X"5F",X"23",
		X"56",X"23",X"46",X"EB",X"3A",X"39",X"20",X"A7",X"C2",X"05",X"09",X"CD",X"0B",X"09",X"E1",X"23",
		X"23",X"23",X"C3",X"E5",X"08",X"CD",X"1B",X"09",X"C3",X"FE",X"08",X"C5",X"E5",X"11",X"7B",X"09",
		X"CD",X"25",X"02",X"E1",X"23",X"C1",X"05",X"C2",X"0B",X"09",X"C9",X"C5",X"E5",X"11",X"83",X"09",
		X"CD",X"25",X"02",X"E1",X"24",X"C1",X"05",X"C2",X"1B",X"09",X"C9",X"05",X"26",X"08",X"11",X"26",
		X"08",X"08",X"29",X"05",X"11",X"29",X"05",X"0B",X"2C",X"02",X"11",X"2C",X"02",X"0B",X"2F",X"02",
		X"11",X"2F",X"02",X"0B",X"32",X"02",X"11",X"32",X"02",X"0B",X"35",X"02",X"11",X"35",X"02",X"0B",
		X"38",X"02",X"11",X"38",X"02",X"08",X"3B",X"05",X"11",X"3B",X"05",X"05",X"3E",X"08",X"11",X"3E",
		X"08",X"FF",X"03",X"28",X"08",X"03",X"35",X"07",X"06",X"2B",X"05",X"06",X"34",X"05",X"18",X"2B",
		X"05",X"18",X"34",X"05",X"1B",X"28",X"08",X"1B",X"34",X"08",X"FF",X"18",X"18",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"00",X"00",X"00",X"01",X"D0",X"01",X"25",X"01",
		X"40",X"04",X"28",X"01",X"40",X"04",X"34",X"01",X"28",X"07",X"2B",X"01",X"28",X"07",X"34",X"01",
		X"28",X"16",X"2B",X"01",X"28",X"16",X"34",X"01",X"40",X"19",X"28",X"01",X"40",X"19",X"34",X"01",
		X"D0",X"1C",X"25",X"FF",X"1A",X"02",X"62",X"24",X"08",X"02",X"65",X"27",X"08",X"02",X"71",X"27",
		X"05",X"02",X"68",X"2A",X"05",X"02",X"71",X"2A",X"08",X"02",X"6B",X"2D",X"02",X"02",X"6B",X"30",
		X"02",X"02",X"71",X"30",X"02",X"02",X"6B",X"33",X"02",X"02",X"71",X"33",X"08",X"02",X"6B",X"36",
		X"05",X"02",X"68",X"39",X"05",X"02",X"71",X"39",X"08",X"02",X"65",X"3C",X"08",X"02",X"71",X"3C",
		X"1A",X"02",X"62",X"3F",X"FF",X"01",X"24",X"04",X"27",X"07",X"2A",X"FF",X"01",X"3F",X"04",X"3C",
		X"07",X"39",X"FF",X"1C",X"24",X"19",X"27",X"16",X"2A",X"FF",X"1C",X"3F",X"19",X"3C",X"16",X"39",
		X"FF",X"00",X"00",X"00",X"F8",X"F8",X"18",X"18",X"18",X"18",X"18",X"18",X"F8",X"F8",X"00",X"00",
		X"00",X"00",X"00",X"00",X"1F",X"1F",X"18",X"18",X"18",X"18",X"18",X"18",X"1F",X"1F",X"00",X"00",
		X"00",X"0D",X"27",X"10",X"27",X"0D",X"2A",X"10",X"2A",X"0A",X"2D",X"13",X"2D",X"04",X"30",X"07",
		X"30",X"0A",X"30",X"0D",X"30",X"10",X"30",X"13",X"30",X"16",X"30",X"19",X"30",X"04",X"33",X"07",
		X"33",X"0A",X"33",X"0D",X"33",X"10",X"33",X"13",X"33",X"16",X"33",X"19",X"33",X"0A",X"36",X"13",
		X"36",X"0D",X"39",X"10",X"39",X"0D",X"3C",X"10",X"3C",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"08",X"00",X"18",X"02",X"30",X"04",X"F8",X"3F",X"30",X"04",X"18",X"02",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"20",X"00",X"20",X"00",X"70",X"00",
		X"A0",X"00",X"20",X"00",X"20",X"00",X"20",X"00",X"70",X"00",X"F8",X"00",X"AC",X"01",X"00",X"00",
		X"00",X"00",X"00",X"10",X"40",X"18",X"20",X"0C",X"FC",X"1F",X"20",X"0C",X"40",X"18",X"00",X"10",
		X"00",X"00",X"00",X"00",X"80",X"35",X"00",X"1F",X"00",X"0E",X"00",X"04",X"00",X"04",X"00",X"04",
		X"00",X"11",X"00",X"0E",X"00",X"04",X"00",X"04",X"00",X"04",X"AF",X"77",X"23",X"1B",X"BA",X"C2",
		X"CB",X"0A",X"BB",X"C2",X"CB",X"0A",X"C9",X"7D",X"E6",X"07",X"D3",X"02",X"CD",X"27",X"0B",X"01",
		X"0B",X"02",X"C9",X"CD",X"D7",X"0A",X"97",X"32",X"29",X"20",X"C5",X"E5",X"1A",X"D3",X"04",X"DB",
		X"03",X"F5",X"A6",X"CA",X"FE",X"0A",X"3E",X"01",X"32",X"29",X"20",X"22",X"2A",X"20",X"F1",X"B6",
		X"77",X"23",X"13",X"05",X"C2",X"EC",X"0A",X"97",X"D3",X"04",X"DB",X"03",X"F5",X"A6",X"CA",X"19",
		X"0B",X"3E",X"01",X"32",X"29",X"20",X"22",X"2A",X"20",X"F1",X"B6",X"77",X"E1",X"01",X"20",X"00",
		X"09",X"C1",X"0D",X"C2",X"EA",X"0A",X"C9",X"C5",X"06",X"03",X"7C",X"1F",X"67",X"7D",X"1F",X"6F",
		X"05",X"C2",X"2A",X"0B",X"7C",X"E6",X"3F",X"F6",X"20",X"67",X"C1",X"C9",X"06",X"06",X"11",X"23",
		X"20",X"7E",X"12",X"23",X"13",X"05",X"C2",X"41",X"0B",X"C9",X"CD",X"D7",X"0A",X"C5",X"E5",X"1A",
		X"D3",X"04",X"DB",X"03",X"AE",X"A6",X"77",X"23",X"13",X"05",X"C2",X"4F",X"0B",X"97",X"D3",X"04",
		X"DB",X"03",X"AE",X"A6",X"77",X"E1",X"01",X"20",X"00",X"09",X"C1",X"0D",X"C2",X"4D",X"0B",X"C9",
		X"CD",X"D7",X"0A",X"97",X"32",X"17",X"21",X"C5",X"E5",X"1A",X"D3",X"04",X"DB",X"03",X"F5",X"A6",
		X"CA",X"8B",X"0B",X"3E",X"01",X"32",X"17",X"21",X"22",X"18",X"21",X"F1",X"AE",X"77",X"23",X"13",
		X"05",X"C2",X"79",X"0B",X"97",X"D3",X"04",X"DB",X"03",X"F5",X"A6",X"CA",X"A6",X"0B",X"3E",X"01",
		X"32",X"17",X"21",X"22",X"18",X"21",X"F1",X"AE",X"77",X"E1",X"01",X"20",X"00",X"09",X"C1",X"0D",
		X"C2",X"77",X"0B",X"C9",X"CD",X"9F",X"07",X"21",X"2B",X"09",X"CD",X"E5",X"08",X"21",X"39",X"20",
		X"36",X"FF",X"21",X"62",X"09",X"CD",X"E5",X"08",X"21",X"3B",X"20",X"36",X"FF",X"E5",X"21",X"F2",
		X"1C",X"CD",X"EA",X"0B",X"E1",X"36",X"00",X"21",X"1B",X"1D",X"C3",X"EA",X"0B",X"AF",X"06",X"08",
		X"77",X"11",X"20",X"00",X"19",X"05",X"C2",X"E0",X"0B",X"C9",X"E5",X"7E",X"FE",X"FF",X"C2",X"F3",
		X"0B",X"E1",X"C9",X"5F",X"23",X"56",X"23",X"46",X"23",X"4E",X"EB",X"3A",X"3B",X"20",X"A7",X"CA",
		X"08",X"0C",X"CD",X"13",X"0C",X"C3",X"0B",X"0C",X"CD",X"1D",X"0C",X"E1",X"23",X"23",X"23",X"23",
		X"C3",X"EA",X"0B",X"71",X"11",X"80",X"00",X"19",X"05",X"C2",X"13",X"0C",X"C9",X"E5",X"71",X"11",
		X"80",X"00",X"19",X"71",X"E1",X"23",X"05",X"C2",X"1D",X"0C",X"C9",X"21",X"42",X"23",X"7E",X"A7",
		X"37",X"C8",X"3F",X"C9",X"CD",X"6A",X"42",X"21",X"1E",X"25",X"11",X"CC",X"1C",X"06",X"1A",X"CD",
		X"22",X"08",X"21",X"1D",X"26",X"11",X"03",X"23",X"CD",X"80",X"0C",X"21",X"1D",X"2F",X"11",X"3F",
		X"23",X"CD",X"80",X"0C",X"3A",X"3B",X"23",X"A7",X"CA",X"64",X"0C",X"21",X"1D",X"39",X"11",X"06",
		X"23",X"CD",X"80",X"0C",X"CD",X"A8",X"45",X"CD",X"9B",X"45",X"21",X"00",X"2A",X"11",X"E6",X"1C",
		X"06",X"04",X"CD",X"22",X"08",X"21",X"00",X"2E",X"01",X"01",X"30",X"3E",X"F8",X"C3",X"DF",X"41",
		X"CD",X"1A",X"04",X"C3",X"43",X"08",X"21",X"00",X"37",X"11",X"EA",X"1C",X"06",X"06",X"C3",X"22",
		X"08",X"3A",X"3D",X"23",X"C6",X"20",X"CD",X"94",X"08",X"21",X"00",X"3E",X"C3",X"AB",X"08",X"21",
		X"00",X"35",X"11",X"DD",X"1B",X"06",X"0A",X"C3",X"22",X"08",X"C3",X"DD",X"1F",X"11",X"B4",X"0A",
		X"CD",X"70",X"0B",X"CD",X"DB",X"18",X"FE",X"02",X"D8",X"FE",X"06",X"21",X"58",X"2A",X"D2",X"CF",
		X"0C",X"FE",X"04",X"21",X"28",X"D2",X"11",X"72",X"0A",X"DA",X"70",X"0B",X"21",X"B8",X"42",X"11",
		X"9E",X"0A",X"C3",X"70",X"0B",X"3A",X"44",X"23",X"A7",X"CA",X"CC",X"0E",X"C3",X"06",X"0D",X"CD",
		X"79",X"04",X"DB",X"01",X"D8",X"DB",X"00",X"C9",X"CD",X"39",X"17",X"21",X"91",X"22",X"35",X"CD",
		X"02",X"0E",X"DB",X"02",X"E6",X"10",X"C4",X"DE",X"0D",X"3A",X"51",X"22",X"A7",X"C2",X"B0",X"0D",
		X"CD",X"2B",X"0C",X"DA",X"D5",X"0C",X"21",X"00",X"20",X"34",X"7E",X"FE",X"03",X"D2",X"44",X"16",
		X"FE",X"02",X"D2",X"45",X"17",X"21",X"01",X"20",X"7E",X"A7",X"C2",X"C7",X"0E",X"23",X"7E",X"A7",
		X"C2",X"82",X"0E",X"2A",X"06",X"20",X"3A",X"04",X"20",X"CD",X"5F",X"07",X"32",X"0A",X"20",X"AF",
		X"47",X"3A",X"42",X"23",X"A7",X"CA",X"A3",X"0D",X"CD",X"D2",X"0E",X"E6",X"0F",X"A7",X"CA",X"76",
		X"12",X"21",X"03",X"20",X"36",X"FF",X"0F",X"DA",X"4F",X"0D",X"04",X"04",X"C3",X"46",X"0D",X"3E",
		X"01",X"80",X"23",X"23",X"77",X"2B",X"7E",X"47",X"23",X"BE",X"CA",X"50",X"12",X"C6",X"04",X"BE",
		X"CA",X"5E",X"12",X"D6",X"08",X"BE",X"CA",X"5E",X"12",X"2A",X"06",X"20",X"11",X"08",X"05",X"19",
		X"3A",X"05",X"20",X"FE",X"05",X"D2",X"64",X"12",X"FE",X"03",X"CA",X"70",X"12",X"11",X"0B",X"00",
		X"19",X"CD",X"27",X"0B",X"7E",X"A7",X"C2",X"76",X"12",X"2A",X"06",X"20",X"E5",X"21",X"28",X"13",
		X"3A",X"0A",X"20",X"E6",X"1F",X"3D",X"C2",X"9E",X"0D",X"5E",X"23",X"56",X"EB",X"E9",X"23",X"23",
		X"C3",X"95",X"0D",X"2A",X"70",X"20",X"7E",X"32",X"05",X"20",X"21",X"04",X"20",X"C3",X"56",X"0D",
		X"DB",X"01",X"E6",X"60",X"C4",X"D8",X"0D",X"CD",X"F2",X"0D",X"E6",X"10",X"06",X"01",X"21",X"40",
		X"22",X"C2",X"CD",X"0D",X"7E",X"A7",X"23",X"C2",X"CD",X"0D",X"2B",X"06",X"00",X"70",X"2A",X"4E",
		X"22",X"23",X"22",X"4E",X"22",X"C3",X"CC",X"0E",X"3E",X"01",X"32",X"56",X"22",X"C9",X"CD",X"E7",
		X"0D",X"CD",X"A8",X"45",X"C3",X"9B",X"45",X"06",X"19",X"21",X"7C",X"46",X"11",X"40",X"22",X"C3",
		X"41",X"0B",X"CD",X"03",X"46",X"DB",X"01",X"C8",X"3A",X"0F",X"23",X"A7",X"DB",X"00",X"C0",X"DB",
		X"01",X"C9",X"DB",X"02",X"E6",X"20",X"C8",X"21",X"90",X"20",X"7E",X"A7",X"C0",X"31",X"00",X"24",
		X"CD",X"4C",X"04",X"CD",X"BA",X"41",X"CD",X"02",X"06",X"21",X"51",X"22",X"77",X"21",X"0E",X"23",
		X"77",X"23",X"77",X"21",X"1C",X"21",X"36",X"00",X"3E",X"10",X"CD",X"89",X"06",X"21",X"00",X"FF",
		X"22",X"42",X"23",X"21",X"00",X"00",X"22",X"44",X"23",X"22",X"46",X"23",X"CD",X"8C",X"04",X"FB",
		X"CD",X"03",X"46",X"C2",X"4C",X"0E",X"CD",X"AC",X"06",X"C3",X"4F",X"0E",X"CD",X"C0",X"06",X"21",
		X"15",X"30",X"11",X"D9",X"1F",X"06",X"04",X"CD",X"22",X"08",X"CD",X"AA",X"41",X"D3",X"06",X"21",
		X"16",X"20",X"36",X"00",X"21",X"90",X"20",X"36",X"00",X"C3",X"19",X"06",X"11",X"C6",X"12",X"C3",
		X"90",X"12",X"3A",X"00",X"20",X"FE",X"03",X"CA",X"A3",X"1A",X"FE",X"02",X"CA",X"68",X"19",X"22",
		X"08",X"20",X"21",X"05",X"20",X"46",X"2B",X"7E",X"57",X"B8",X"C2",X"94",X"0E",X"2B",X"2B",X"36",
		X"00",X"C3",X"C7",X"0E",X"48",X"DA",X"BA",X"0F",X"07",X"07",X"07",X"07",X"B1",X"FE",X"71",X"36",
		X"08",X"CA",X"AD",X"0E",X"FE",X"81",X"36",X"01",X"CA",X"AD",X"0E",X"15",X"72",X"2B",X"2B",X"36",
		X"FF",X"CD",X"DC",X"0E",X"3A",X"09",X"20",X"DA",X"E6",X"0E",X"FE",X"80",X"D2",X"C7",X"0E",X"CD",
		X"89",X"13",X"21",X"01",X"20",X"36",X"01",X"21",X"2C",X"20",X"36",X"FF",X"F1",X"C1",X"D1",X"E1",
		X"FB",X"C9",X"DB",X"02",X"E6",X"40",X"C2",X"DF",X"0C",X"DB",X"01",X"C9",X"DB",X"02",X"E6",X"40",
		X"C2",X"79",X"04",X"37",X"3F",X"C9",X"FE",X"80",X"DA",X"C7",X"0E",X"C3",X"BF",X"0E",X"3A",X"70",
		X"22",X"A7",X"C4",X"0B",X"0F",X"3A",X"78",X"22",X"A7",X"C4",X"29",X"0F",X"3A",X"80",X"22",X"A7",
		X"C4",X"47",X"0F",X"3A",X"88",X"22",X"A7",X"C2",X"65",X"0F",X"C9",X"2A",X"73",X"22",X"7C",X"FE",
		X"30",X"DA",X"83",X"0F",X"7D",X"FE",X"E0",X"D2",X"83",X"0F",X"CD",X"AF",X"41",X"21",X"73",X"22",
		X"CD",X"CF",X"41",X"21",X"71",X"22",X"C3",X"5A",X"41",X"2A",X"7B",X"22",X"7C",X"FE",X"E0",X"D2",
		X"A5",X"0F",X"7D",X"FE",X"D0",X"D2",X"A5",X"0F",X"CD",X"AF",X"41",X"21",X"7B",X"22",X"CD",X"CF",
		X"41",X"21",X"79",X"22",X"C3",X"5A",X"41",X"2A",X"83",X"22",X"7C",X"FE",X"E0",X"D2",X"AC",X"0F",
		X"7D",X"FE",X"10",X"DA",X"AC",X"0F",X"CD",X"AF",X"41",X"21",X"83",X"22",X"CD",X"CF",X"41",X"21",
		X"81",X"22",X"C3",X"5A",X"41",X"2A",X"8B",X"22",X"7C",X"FE",X"30",X"DA",X"B3",X"0F",X"7D",X"FE",
		X"10",X"DA",X"B3",X"0F",X"CD",X"AF",X"41",X"21",X"8B",X"22",X"CD",X"CF",X"41",X"21",X"89",X"22",
		X"C3",X"5A",X"41",X"AF",X"32",X"70",X"22",X"3A",X"70",X"22",X"A7",X"C0",X"3A",X"78",X"22",X"A7",
		X"C0",X"3A",X"80",X"22",X"A7",X"C0",X"3A",X"88",X"22",X"A7",X"C0",X"32",X"90",X"22",X"32",X"92",
		X"22",X"32",X"3D",X"20",X"C9",X"AF",X"32",X"78",X"22",X"C3",X"87",X"0F",X"AF",X"32",X"80",X"22",
		X"C3",X"87",X"0F",X"AF",X"32",X"88",X"22",X"C3",X"87",X"0F",X"07",X"07",X"07",X"07",X"B1",X"FE",
		X"17",X"36",X"08",X"CA",X"AD",X"0E",X"FE",X"18",X"36",X"01",X"CA",X"AD",X"0E",X"14",X"C3",X"AC",
		X"0E",X"11",X"DE",X"12",X"C3",X"21",X"12",X"11",X"D8",X"12",X"C3",X"90",X"12",X"11",X"0E",X"13",
		X"C3",X"21",X"12",X"11",X"CC",X"12",X"C3",X"90",X"12",X"11",X"E4",X"12",X"C3",X"21",X"12",X"11",
		X"D2",X"12",X"C3",X"90",X"12",X"11",X"08",X"13",X"C3",X"21",X"12",X"11",X"EA",X"12",X"C3",X"21",
		X"12",X"11",X"F0",X"12",X"C3",X"21",X"12",X"11",X"FC",X"12",X"C3",X"21",X"12",X"11",X"02",X"13",
		X"C3",X"21",X"12",X"11",X"14",X"13",X"21",X"2F",X"20",X"06",X"0A",X"CD",X"47",X"12",X"E1",X"7C",
		X"FE",X"80",X"D2",X"33",X"10",X"FE",X"68",X"2A",X"31",X"20",X"D2",X"72",X"0E",X"2A",X"2F",X"20",
		X"C3",X"72",X"0E",X"FE",X"9C",X"D2",X"3E",X"10",X"2A",X"33",X"20",X"C3",X"72",X"0E",X"FE",X"B4",
		X"2A",X"37",X"20",X"D2",X"72",X"0E",X"2A",X"35",X"20",X"C3",X"72",X"0E",X"11",X"1E",X"13",X"C3",
		X"16",X"10",X"E1",X"7C",X"FE",X"38",X"D2",X"5F",X"10",X"21",X"70",X"2A",X"C3",X"72",X"0E",X"FE",
		X"50",X"21",X"70",X"5A",X"D2",X"72",X"0E",X"21",X"70",X"42",X"C3",X"72",X"0E",X"E1",X"7C",X"FE",
		X"80",X"D2",X"7A",X"10",X"21",X"70",X"72",X"C3",X"72",X"0E",X"FE",X"98",X"21",X"70",X"A2",X"D2",
		X"72",X"0E",X"21",X"70",X"8A",X"C3",X"72",X"0E",X"E1",X"7C",X"FE",X"C8",X"D2",X"95",X"10",X"21",
		X"70",X"BA",X"C3",X"72",X"0E",X"FE",X"E0",X"21",X"70",X"EA",X"D2",X"72",X"0E",X"21",X"70",X"D2",
		X"C3",X"72",X"0E",X"E1",X"7D",X"FE",X"B2",X"D2",X"B6",X"10",X"FE",X"39",X"DA",X"C4",X"10",X"E5",
		X"11",X"F6",X"12",X"C3",X"21",X"12",X"FE",X"C6",X"21",X"D0",X"8A",X"D2",X"72",X"0E",X"21",X"B8",
		X"8A",X"C3",X"72",X"0E",X"FE",X"22",X"21",X"28",X"8A",X"D2",X"72",X"0E",X"21",X"10",X"8A",X"C3",
		X"72",X"0E",X"21",X"2A",X"EA",X"22",X"17",X"20",X"E1",X"78",X"FE",X"03",X"CA",X"B1",X"11",X"7C",
		X"CD",X"0D",X"12",X"21",X"18",X"20",X"46",X"B8",X"D2",X"C7",X"0E",X"21",X"09",X"20",X"77",X"CD",
		X"DC",X"0E",X"3A",X"09",X"20",X"DA",X"82",X"11",X"FE",X"80",X"D2",X"C7",X"0E",X"CD",X"89",X"13",
		X"21",X"02",X"20",X"7E",X"A7",X"CA",X"0B",X"11",X"2B",X"36",X"01",X"3A",X"29",X"20",X"A7",X"C2",
		X"1D",X"11",X"21",X"2C",X"20",X"7E",X"A7",X"CA",X"C7",X"0E",X"C3",X"C0",X"14",X"2A",X"2A",X"20",
		X"22",X"1E",X"20",X"2A",X"06",X"21",X"CD",X"5C",X"11",X"D2",X"BF",X"1C",X"2A",X"06",X"22",X"CD",
		X"5C",X"11",X"D2",X"BF",X"1C",X"21",X"1C",X"20",X"36",X"FF",X"23",X"34",X"2A",X"2A",X"20",X"3E",
		X"1F",X"A5",X"6F",X"3A",X"05",X"20",X"0F",X"0F",X"DA",X"55",X"11",X"AF",X"77",X"11",X"20",X"00",
		X"19",X"77",X"C3",X"12",X"11",X"11",X"60",X"00",X"19",X"C3",X"4B",X"11",X"CD",X"27",X"0B",X"7D",
		X"E6",X"1F",X"47",X"3A",X"1E",X"20",X"E6",X"1F",X"B8",X"CA",X"73",X"11",X"3D",X"B8",X"CA",X"73",
		X"11",X"37",X"C9",X"3A",X"1F",X"20",X"BC",X"CA",X"7F",X"11",X"3D",X"BC",X"C2",X"71",X"11",X"37",
		X"3F",X"C9",X"FE",X"80",X"DA",X"C7",X"0E",X"C3",X"FD",X"10",X"21",X"42",X"D2",X"C3",X"D5",X"10",
		X"21",X"5A",X"BA",X"C3",X"D5",X"10",X"21",X"2A",X"5A",X"C3",X"D5",X"10",X"21",X"72",X"A2",X"C3",
		X"D5",X"10",X"21",X"BA",X"EA",X"C3",X"D5",X"10",X"C3",X"90",X"11",X"C3",X"8A",X"11",X"C3",X"D2",
		X"10",X"7C",X"CD",X"17",X"12",X"21",X"17",X"20",X"46",X"B8",X"DA",X"C7",X"0E",X"C3",X"EB",X"10",
		X"21",X"D2",X"12",X"22",X"19",X"20",X"E1",X"78",X"FE",X"01",X"CA",X"E0",X"11",X"7D",X"CD",X"17",
		X"12",X"21",X"1A",X"20",X"46",X"B8",X"DA",X"C7",X"0E",X"21",X"08",X"20",X"77",X"C3",X"EF",X"10",
		X"7D",X"CD",X"0D",X"12",X"21",X"19",X"20",X"46",X"B8",X"D2",X"C7",X"0E",X"C3",X"D9",X"11",X"21",
		X"BA",X"2A",X"C3",X"C3",X"11",X"21",X"A2",X"42",X"C3",X"C3",X"11",X"C3",X"F5",X"11",X"C3",X"C0",
		X"11",X"C3",X"F5",X"11",X"C3",X"F5",X"11",X"C3",X"EF",X"11",X"C3",X"C0",X"11",X"21",X"0B",X"20",
		X"46",X"3C",X"05",X"C2",X"11",X"12",X"C9",X"21",X"0B",X"20",X"46",X"3D",X"05",X"C2",X"1B",X"12",
		X"C9",X"21",X"2F",X"20",X"CD",X"45",X"12",X"E1",X"7D",X"FE",X"88",X"DA",X"34",X"12",X"2A",X"2F",
		X"20",X"C3",X"72",X"0E",X"FE",X"60",X"DA",X"3F",X"12",X"2A",X"31",X"20",X"C3",X"72",X"0E",X"2A",
		X"33",X"20",X"C3",X"72",X"0E",X"06",X"06",X"1A",X"77",X"23",X"13",X"05",X"C2",X"47",X"12",X"C9",
		X"2A",X"06",X"20",X"E5",X"21",X"04",X"20",X"46",X"21",X"4C",X"13",X"C3",X"90",X"0D",X"2A",X"06",
		X"20",X"C3",X"72",X"0E",X"11",X"00",X"0C",X"C2",X"80",X"0D",X"11",X"F5",X"FF",X"C3",X"80",X"0D",
		X"11",X"00",X"F5",X"C3",X"80",X"0D",X"21",X"03",X"20",X"36",X"00",X"21",X"04",X"20",X"46",X"23",
		X"70",X"C3",X"50",X"12",X"21",X"D0",X"EA",X"C3",X"7F",X"0E",X"21",X"D0",X"8A",X"C3",X"7F",X"0E",
		X"21",X"2F",X"20",X"CD",X"45",X"12",X"E1",X"7C",X"FE",X"80",X"D2",X"A3",X"12",X"2A",X"2F",X"20",
		X"C3",X"72",X"0E",X"FE",X"C0",X"D2",X"AE",X"12",X"2A",X"31",X"20",X"C3",X"72",X"0E",X"2A",X"33",
		X"20",X"C3",X"72",X"0E",X"23",X"47",X"8B",X"11",X"10",X"12",X"89",X"45",X"21",X"24",X"48",X"8C",
		X"0D",X"0E",X"0F",X"8A",X"46",X"22",X"D0",X"2A",X"D0",X"8A",X"D0",X"EA",X"B8",X"42",X"B8",X"8A",
		X"B8",X"D2",X"28",X"42",X"28",X"8A",X"28",X"D2",X"10",X"2A",X"10",X"8A",X"10",X"EA",X"D0",X"EA",
		X"70",X"EA",X"10",X"EA",X"B8",X"D2",X"70",X"D2",X"28",X"D2",X"A0",X"BA",X"70",X"BA",X"40",X"BA",
		X"A0",X"A2",X"70",X"A2",X"40",X"A2",X"A0",X"8A",X"70",X"8A",X"40",X"8A",X"A0",X"72",X"70",X"72",
		X"40",X"72",X"A0",X"5A",X"70",X"5A",X"40",X"5A",X"B8",X"42",X"70",X"42",X"28",X"42",X"D0",X"2A",
		X"70",X"2A",X"10",X"2A",X"A0",X"5A",X"A0",X"72",X"A0",X"8A",X"A0",X"A2",X"A0",X"BA",X"40",X"5A",
		X"40",X"72",X"40",X"8A",X"40",X"A2",X"40",X"BA",X"6C",X"0E",X"D1",X"0F",X"D7",X"0F",X"DD",X"0F",
		X"E3",X"0F",X"E9",X"0F",X"EF",X"0F",X"F5",X"0F",X"13",X"10",X"FB",X"0F",X"4C",X"10",X"0D",X"10",
		X"07",X"10",X"A3",X"10",X"01",X"10",X"52",X"10",X"6D",X"10",X"88",X"10",X"D2",X"10",X"C0",X"11",
		X"AE",X"11",X"0A",X"12",X"8A",X"11",X"EF",X"11",X"AB",X"11",X"07",X"12",X"90",X"11",X"F5",X"11",
		X"A8",X"11",X"04",X"12",X"01",X"12",X"FE",X"11",X"FB",X"11",X"96",X"11",X"9C",X"11",X"A2",X"11",
		X"2A",X"06",X"20",X"CD",X"A0",X"42",X"01",X"04",X"02",X"7B",X"C3",X"D2",X"08",X"2A",X"06",X"21",
		X"C3",X"73",X"13",X"2A",X"06",X"22",X"C3",X"73",X"13",X"2A",X"0E",X"20",X"EB",X"2A",X"06",X"20",
		X"CD",X"4A",X"0B",X"1E",X"FF",X"CD",X"70",X"13",X"2A",X"10",X"20",X"EB",X"2A",X"08",X"20",X"CD",
		X"E3",X"0A",X"2A",X"10",X"20",X"22",X"0E",X"20",X"2A",X"08",X"20",X"22",X"06",X"20",X"1E",X"05",
		X"C3",X"70",X"13",X"3A",X"92",X"22",X"A7",X"C4",X"EE",X"0E",X"DB",X"01",X"07",X"DA",X"04",X"14",
		X"21",X"3E",X"23",X"7E",X"A7",X"CA",X"E4",X"13",X"2B",X"7E",X"FE",X"09",X"D2",X"FC",X"13",X"3C",
		X"77",X"FE",X"09",X"D2",X"FC",X"13",X"3A",X"42",X"23",X"A7",X"C2",X"E0",X"13",X"CD",X"91",X"0C",
		X"AF",X"32",X"3E",X"23",X"3A",X"43",X"23",X"A7",X"CA",X"98",X"14",X"3A",X"42",X"23",X"A7",X"C2",
		X"98",X"14",X"3A",X"3D",X"23",X"A7",X"C2",X"09",X"14",X"C3",X"9B",X"40",X"3E",X"04",X"CD",X"7E",
		X"06",X"C3",X"DD",X"13",X"3E",X"01",X"C3",X"E1",X"13",X"3A",X"16",X"20",X"A7",X"C2",X"CC",X"0E",
		X"3E",X"01",X"32",X"16",X"20",X"31",X"00",X"24",X"FB",X"CD",X"BA",X"41",X"21",X"44",X"23",X"36",
		X"00",X"CD",X"D5",X"04",X"CD",X"F7",X"45",X"21",X"13",X"30",X"11",X"56",X"47",X"06",X"04",X"CD",
		X"22",X"08",X"3A",X"3D",X"23",X"3D",X"21",X"11",X"27",X"06",X"16",X"C2",X"75",X"14",X"11",X"F2",
		X"1B",X"CD",X"22",X"08",X"DB",X"01",X"E6",X"40",X"CA",X"32",X"14",X"CD",X"48",X"05",X"06",X"99",
		X"AF",X"32",X"3B",X"23",X"3A",X"3D",X"23",X"80",X"27",X"32",X"3D",X"23",X"3E",X"04",X"CD",X"89",
		X"06",X"CD",X"91",X"0C",X"21",X"43",X"23",X"36",X"00",X"C3",X"E1",X"47",X"11",X"06",X"00",X"CD",
		X"CA",X"0A",X"C3",X"4A",X"00",X"11",X"9D",X"1B",X"CD",X"22",X"08",X"DB",X"01",X"07",X"07",X"DA",
		X"4B",X"14",X"07",X"DA",X"89",X"14",X"C3",X"32",X"14",X"CD",X"48",X"05",X"21",X"3B",X"23",X"36",
		X"FF",X"06",X"98",X"3E",X"FF",X"C3",X"51",X"14",X"21",X"20",X"20",X"7E",X"A7",X"CA",X"A4",X"14",
		X"35",X"C3",X"A9",X"14",X"3E",X"01",X"CD",X"A0",X"06",X"21",X"2C",X"20",X"7E",X"A7",X"C2",X"C8",
		X"14",X"23",X"7E",X"A7",X"C2",X"FD",X"1A",X"23",X"7E",X"A7",X"C2",X"98",X"15",X"C3",X"CC",X"0E",
		X"21",X"2C",X"20",X"36",X"00",X"C3",X"CC",X"0E",X"21",X"01",X"20",X"7E",X"A7",X"CA",X"D4",X"14",
		X"35",X"C3",X"C0",X"14",X"CD",X"DC",X"0E",X"3A",X"09",X"20",X"DA",X"E8",X"14",X"FE",X"80",X"DA",
		X"C0",X"14",X"CD",X"89",X"13",X"C3",X"00",X"11",X"FE",X"80",X"D2",X"C0",X"14",X"C3",X"E2",X"14",
		X"21",X"3A",X"20",X"7E",X"A7",X"C2",X"DC",X"17",X"36",X"FF",X"3A",X"04",X"21",X"0F",X"0F",X"DA",
		X"1B",X"15",X"21",X"06",X"21",X"7E",X"26",X"20",X"46",X"B8",X"D2",X"16",X"15",X"3E",X"01",X"21",
		X"05",X"21",X"77",X"C3",X"6E",X"19",X"3E",X"05",X"C3",X"0F",X"15",X"21",X"07",X"21",X"7E",X"26",
		X"20",X"46",X"B8",X"3E",X"07",X"DA",X"0F",X"15",X"3E",X"03",X"C3",X"0F",X"15",X"C2",X"33",X"15",
		X"C3",X"BD",X"17",X"2A",X"06",X"21",X"CD",X"D4",X"1A",X"32",X"05",X"21",X"CD",X"E1",X"1A",X"C3",
		X"D3",X"17",X"21",X"0C",X"20",X"C3",X"10",X"12",X"21",X"0C",X"20",X"C3",X"1A",X"12",X"21",X"0D",
		X"20",X"C3",X"10",X"12",X"21",X"0D",X"20",X"C3",X"1A",X"12",X"21",X"14",X"21",X"36",X"07",X"C3",
		X"ED",X"18",X"21",X"14",X"21",X"36",X"03",X"21",X"BA",X"2A",X"C3",X"F0",X"18",X"21",X"14",X"21",
		X"36",X"07",X"C3",X"67",X"15",X"21",X"14",X"21",X"36",X"03",X"21",X"A2",X"42",X"C3",X"F0",X"18",
		X"21",X"14",X"21",X"36",X"07",X"C3",X"7A",X"15",X"C3",X"80",X"15",X"C3",X"E8",X"18",X"C3",X"80",
		X"15",X"2A",X"06",X"21",X"E5",X"C3",X"CF",X"18",X"21",X"46",X"20",X"7E",X"A7",X"C2",X"B6",X"15",
		X"2B",X"2B",X"34",X"7E",X"FE",X"F0",X"DA",X"B6",X"15",X"36",X"00",X"23",X"34",X"7E",X"FE",X"0A",
		X"DA",X"B6",X"15",X"23",X"36",X"FF",X"0E",X"03",X"3A",X"42",X"23",X"A7",X"CA",X"DC",X"15",X"CD",
		X"D2",X"0E",X"E6",X"10",X"A7",X"CA",X"13",X"16",X"21",X"48",X"20",X"7E",X"FE",X"18",X"D2",X"DC",
		X"15",X"3E",X"02",X"CD",X"95",X"06",X"21",X"47",X"20",X"34",X"0E",X"04",X"3A",X"46",X"20",X"A7",
		X"CA",X"E5",X"15",X"0E",X"02",X"21",X"0B",X"20",X"71",X"21",X"1C",X"21",X"7E",X"A7",X"C2",X"F7",
		X"15",X"23",X"7E",X"A7",X"CA",X"2A",X"16",X"CD",X"DC",X"0E",X"3A",X"09",X"22",X"DA",X"0B",X"16",
		X"FE",X"80",X"DA",X"2A",X"16",X"CD",X"00",X"17",X"C3",X"2A",X"16",X"FE",X"80",X"D2",X"2A",X"16",
		X"C3",X"05",X"16",X"3E",X"02",X"CD",X"A0",X"06",X"0E",X"03",X"C3",X"DC",X"15",X"21",X"2E",X"20",
		X"36",X"FF",X"21",X"00",X"20",X"36",X"00",X"C3",X"CC",X"0E",X"21",X"2E",X"20",X"36",X"00",X"C3",
		X"CC",X"0E",X"3A",X"17",X"21",X"A7",X"37",X"C8",X"2A",X"18",X"21",X"22",X"1E",X"20",X"2A",X"06",
		X"20",X"C3",X"5C",X"11",X"21",X"1C",X"21",X"7E",X"A7",X"C2",X"A8",X"19",X"23",X"7E",X"A7",X"CA",
		X"1D",X"16",X"CD",X"32",X"16",X"D2",X"BF",X"1C",X"2A",X"06",X"22",X"EB",X"2A",X"0F",X"22",X"19",
		X"EB",X"21",X"10",X"22",X"7E",X"07",X"D2",X"9D",X"16",X"2B",X"7E",X"07",X"23",X"23",X"7A",X"D2",
		X"73",X"16",X"7B",X"46",X"B8",X"DA",X"7B",X"16",X"C3",X"A9",X"16",X"CD",X"D6",X"16",X"CD",X"B0",
		X"16",X"CD",X"DC",X"0E",X"3A",X"09",X"22",X"DA",X"95",X"16",X"FE",X"80",X"D2",X"1D",X"16",X"CD",
		X"00",X"17",X"C3",X"1D",X"16",X"FE",X"80",X"DA",X"1D",X"16",X"C3",X"8F",X"16",X"A7",X"23",X"7A",
		X"C2",X"A4",X"16",X"7B",X"46",X"B8",X"D2",X"7B",X"16",X"EB",X"22",X"08",X"22",X"C3",X"81",X"16",
		X"21",X"10",X"22",X"7E",X"07",X"D2",X"C8",X"16",X"2B",X"7E",X"07",X"21",X"88",X"0A",X"D2",X"C4",
		X"16",X"21",X"9E",X"0A",X"22",X"0D",X"22",X"C9",X"0F",X"A7",X"21",X"B4",X"0A",X"C2",X"C4",X"16",
		X"21",X"72",X"0A",X"C3",X"C4",X"16",X"21",X"1F",X"21",X"34",X"7E",X"2B",X"BE",X"DA",X"E3",X"16",
		X"23",X"36",X"00",X"21",X"20",X"21",X"01",X"05",X"00",X"3D",X"CA",X"F1",X"16",X"09",X"C3",X"E9",
		X"16",X"11",X"0F",X"22",X"06",X"05",X"CD",X"41",X"0B",X"2A",X"12",X"22",X"22",X"08",X"22",X"C9",
		X"2A",X"0B",X"22",X"EB",X"2A",X"06",X"22",X"CD",X"70",X"0B",X"2A",X"0D",X"22",X"EB",X"2A",X"08",
		X"22",X"CD",X"70",X"0B",X"CD",X"DB",X"18",X"FE",X"04",X"DA",X"21",X"17",X"1E",X"FF",X"CD",X"83",
		X"13",X"2A",X"0D",X"22",X"22",X"0B",X"22",X"2A",X"08",X"22",X"22",X"06",X"22",X"CD",X"DB",X"18",
		X"FE",X"04",X"D8",X"1E",X"03",X"CD",X"83",X"13",X"C9",X"21",X"2C",X"20",X"36",X"00",X"23",X"36",
		X"00",X"23",X"36",X"00",X"C9",X"CD",X"39",X"17",X"CD",X"32",X"16",X"D2",X"BF",X"1C",X"21",X"02",
		X"21",X"7E",X"A7",X"C2",X"6B",X"19",X"2A",X"06",X"21",X"3A",X"04",X"21",X"CD",X"5F",X"07",X"FE",
		X"A0",X"C2",X"6C",X"17",X"3E",X"07",X"32",X"04",X"21",X"C3",X"6F",X"17",X"32",X"0A",X"21",X"21",
		X"15",X"21",X"7E",X"A7",X"CA",X"7B",X"17",X"35",X"C3",X"DC",X"17",X"21",X"14",X"21",X"36",X"00",
		X"21",X"0A",X"20",X"7E",X"26",X"21",X"BE",X"CA",X"F0",X"14",X"47",X"AF",X"32",X"3A",X"20",X"78",
		X"E6",X"1F",X"FE",X"0D",X"D2",X"A2",X"17",X"78",X"E6",X"E0",X"47",X"7E",X"E6",X"E0",X"B8",X"CA",
		X"E9",X"17",X"2E",X"1B",X"36",X"00",X"2E",X"0A",X"7E",X"E6",X"1F",X"FE",X"10",X"D2",X"54",X"1B",
		X"FE",X"0E",X"CA",X"22",X"18",X"3A",X"04",X"21",X"0F",X"0F",X"DA",X"33",X"15",X"2A",X"06",X"21",
		X"44",X"EB",X"3A",X"07",X"20",X"B8",X"3E",X"07",X"D2",X"CD",X"17",X"3E",X"03",X"32",X"05",X"21",
		X"CD",X"C5",X"1A",X"19",X"CD",X"27",X"0B",X"7E",X"A7",X"CA",X"5B",X"19",X"2A",X"06",X"21",X"E5",
		X"3A",X"0A",X"21",X"21",X"79",X"1B",X"C3",X"93",X"0D",X"7E",X"26",X"20",X"46",X"90",X"FE",X"02",
		X"CA",X"F8",X"17",X"FE",X"FE",X"C2",X"DC",X"17",X"21",X"0F",X"21",X"7E",X"A7",X"C2",X"DC",X"17",
		X"36",X"FF",X"3A",X"05",X"20",X"32",X"05",X"21",X"C3",X"6B",X"19",X"3A",X"04",X"21",X"FE",X"03",
		X"26",X"20",X"7E",X"C2",X"1D",X"18",X"E6",X"20",X"C0",X"2A",X"06",X"21",X"C9",X"E6",X"80",X"C3",
		X"18",X"18",X"26",X"20",X"7E",X"E6",X"20",X"CA",X"31",X"18",X"2A",X"06",X"21",X"E5",X"C3",X"ED",
		X"18",X"7E",X"FE",X"11",X"C2",X"B5",X"17",X"3A",X"06",X"21",X"FE",X"30",X"DA",X"B5",X"17",X"FE",
		X"C0",X"D2",X"B5",X"17",X"C3",X"2A",X"18",X"21",X"14",X"21",X"36",X"05",X"21",X"2A",X"EA",X"22",
		X"12",X"21",X"E1",X"3A",X"00",X"20",X"FE",X"03",X"D2",X"13",X"1A",X"3A",X"04",X"21",X"FE",X"03",
		X"CA",X"76",X"18",X"7C",X"CD",X"42",X"15",X"21",X"13",X"21",X"46",X"B8",X"D2",X"82",X"18",X"21",
		X"09",X"21",X"77",X"C3",X"87",X"19",X"7C",X"CD",X"48",X"15",X"21",X"12",X"21",X"46",X"B8",X"D2",
		X"6F",X"18",X"3A",X"14",X"21",X"A7",X"C2",X"53",X"19",X"21",X"06",X"21",X"7E",X"26",X"20",X"46",
		X"B8",X"3E",X"01",X"DA",X"53",X"19",X"3E",X"05",X"C3",X"53",X"19",X"21",X"14",X"21",X"36",X"01",
		X"C3",X"4C",X"18",X"21",X"14",X"21",X"36",X"05",X"21",X"42",X"D2",X"C3",X"4F",X"18",X"21",X"14",
		X"21",X"36",X"01",X"C3",X"A8",X"18",X"21",X"14",X"21",X"36",X"05",X"21",X"5A",X"BA",X"C3",X"4F",
		X"18",X"21",X"14",X"21",X"36",X"01",X"C3",X"BB",X"18",X"21",X"2A",X"5A",X"C3",X"4F",X"18",X"21",
		X"72",X"A2",X"C3",X"4F",X"18",X"21",X"BA",X"EA",X"C3",X"4F",X"18",X"CD",X"79",X"04",X"21",X"31",
		X"23",X"DA",X"E6",X"18",X"2E",X"32",X"7E",X"C9",X"21",X"14",X"21",X"36",X"03",X"21",X"D2",X"12",
		X"22",X"10",X"21",X"E1",X"3A",X"00",X"20",X"FE",X"03",X"D2",X"53",X"1A",X"3A",X"04",X"21",X"FE",
		X"01",X"CA",X"30",X"19",X"7D",X"CD",X"48",X"15",X"21",X"11",X"21",X"46",X"B8",X"DA",X"3C",X"19",
		X"21",X"08",X"21",X"77",X"CD",X"DC",X"0E",X"3A",X"09",X"21",X"DA",X"28",X"19",X"FE",X"80",X"D2",
		X"98",X"19",X"CD",X"2A",X"1B",X"C3",X"98",X"19",X"FE",X"80",X"DA",X"98",X"19",X"C3",X"22",X"19",
		X"7D",X"CD",X"42",X"15",X"21",X"10",X"21",X"46",X"B8",X"DA",X"10",X"19",X"21",X"07",X"21",X"3A",
		X"14",X"21",X"A7",X"C2",X"53",X"19",X"7C",X"21",X"07",X"20",X"46",X"B8",X"3E",X"07",X"DA",X"53",
		X"19",X"3E",X"03",X"32",X"05",X"21",X"21",X"14",X"21",X"36",X"00",X"2A",X"06",X"21",X"E5",X"3A",
		X"0A",X"21",X"21",X"28",X"13",X"C3",X"93",X"0D",X"22",X"08",X"21",X"21",X"05",X"21",X"46",X"2B",
		X"7E",X"57",X"B8",X"C2",X"82",X"19",X"2B",X"2B",X"36",X"00",X"21",X"15",X"21",X"36",X"06",X"C3",
		X"98",X"19",X"70",X"2B",X"2B",X"36",X"FF",X"CD",X"DC",X"0E",X"3A",X"09",X"21",X"DA",X"A0",X"19",
		X"FE",X"80",X"D2",X"98",X"19",X"CD",X"2A",X"1B",X"21",X"2D",X"20",X"36",X"FF",X"C3",X"CC",X"0E",
		X"FE",X"80",X"DA",X"98",X"19",X"C3",X"95",X"19",X"CD",X"32",X"16",X"D2",X"BF",X"1C",X"3A",X"02",
		X"22",X"A7",X"C2",X"A6",X"1A",X"2A",X"08",X"22",X"3A",X"04",X"22",X"CD",X"5F",X"07",X"32",X"0A",
		X"22",X"21",X"01",X"22",X"7E",X"A7",X"CA",X"CD",X"19",X"35",X"C3",X"FA",X"19",X"21",X"14",X"21",
		X"36",X"00",X"21",X"04",X"22",X"7E",X"0F",X"0F",X"DA",X"04",X"1A",X"2A",X"06",X"22",X"44",X"EB",
		X"3A",X"07",X"20",X"B8",X"3E",X"07",X"D2",X"EB",X"19",X"3E",X"03",X"32",X"05",X"22",X"CD",X"C5",
		X"1A",X"19",X"CD",X"27",X"0B",X"7E",X"A7",X"CA",X"99",X"1A",X"2A",X"06",X"22",X"E5",X"3A",X"0A",
		X"22",X"C3",X"E3",X"17",X"2A",X"06",X"22",X"CD",X"D4",X"1A",X"32",X"05",X"22",X"CD",X"E1",X"1A",
		X"C3",X"F1",X"19",X"3A",X"04",X"22",X"FE",X"03",X"CA",X"2E",X"1A",X"7C",X"CD",X"4E",X"15",X"21",
		X"13",X"21",X"46",X"B8",X"D2",X"3A",X"1A",X"21",X"09",X"22",X"77",X"C3",X"81",X"16",X"7C",X"CD",
		X"54",X"15",X"21",X"12",X"21",X"46",X"B8",X"D2",X"27",X"1A",X"3A",X"14",X"21",X"A7",X"C2",X"91",
		X"1A",X"21",X"06",X"22",X"7E",X"26",X"20",X"46",X"B8",X"3E",X"01",X"DA",X"91",X"1A",X"3E",X"05",
		X"C3",X"91",X"1A",X"3A",X"04",X"22",X"FE",X"01",X"CA",X"6E",X"1A",X"7D",X"CD",X"54",X"15",X"21",
		X"11",X"21",X"46",X"B8",X"DA",X"7A",X"1A",X"21",X"08",X"22",X"77",X"C3",X"81",X"16",X"7D",X"CD",
		X"4E",X"15",X"21",X"10",X"21",X"46",X"B8",X"DA",X"67",X"1A",X"21",X"07",X"22",X"3A",X"14",X"21",
		X"A7",X"C2",X"91",X"1A",X"7C",X"21",X"07",X"20",X"46",X"B8",X"3E",X"07",X"DA",X"91",X"1A",X"3E",
		X"03",X"32",X"05",X"22",X"21",X"14",X"21",X"36",X"00",X"2A",X"06",X"22",X"E5",X"3A",X"0A",X"22",
		X"C3",X"62",X"19",X"22",X"08",X"22",X"21",X"05",X"22",X"46",X"2B",X"7E",X"57",X"B8",X"C2",X"BD",
		X"1A",X"2B",X"2B",X"36",X"00",X"21",X"01",X"22",X"36",X"0A",X"C3",X"1D",X"16",X"70",X"2B",X"2B",
		X"36",X"FF",X"C3",X"81",X"16",X"EB",X"11",X"08",X"05",X"19",X"FE",X"03",X"11",X"00",X"0C",X"C0",
		X"11",X"00",X"F4",X"C9",X"45",X"EB",X"2A",X"06",X"20",X"7D",X"B8",X"3E",X"01",X"D0",X"3E",X"05",
		X"C9",X"EB",X"11",X"08",X"05",X"19",X"FE",X"01",X"11",X"F4",X"FF",X"C0",X"11",X"0C",X"00",X"C9",
		X"21",X"72",X"0A",X"3D",X"C8",X"11",X"16",X"00",X"19",X"3D",X"C3",X"F3",X"1A",X"21",X"01",X"21",
		X"7E",X"A7",X"CA",X"0E",X"1B",X"35",X"21",X"2D",X"20",X"36",X"00",X"C3",X"CC",X"0E",X"CD",X"DC",
		X"0E",X"3A",X"09",X"21",X"DA",X"22",X"1B",X"FE",X"80",X"DA",X"06",X"1B",X"CD",X"2A",X"1B",X"C3",
		X"06",X"1B",X"FE",X"80",X"D2",X"06",X"1B",X"C3",X"1C",X"1B",X"2A",X"0B",X"21",X"EB",X"2A",X"06",
		X"21",X"CD",X"70",X"0B",X"2A",X"0D",X"21",X"EB",X"2A",X"08",X"21",X"CD",X"70",X"0B",X"1E",X"FF",
		X"CD",X"7D",X"13",X"2A",X"0D",X"21",X"22",X"0B",X"21",X"2A",X"08",X"21",X"22",X"06",X"21",X"1E",
		X"03",X"C3",X"7D",X"13",X"0F",X"DA",X"91",X"15",X"0F",X"DA",X"B5",X"17",X"3A",X"04",X"21",X"FE",
		X"03",X"21",X"0A",X"20",X"7E",X"C2",X"B5",X"17",X"E6",X"20",X"CA",X"B5",X"17",X"21",X"14",X"21",
		X"36",X"05",X"2A",X"06",X"21",X"E5",X"C3",X"CF",X"18",X"47",X"18",X"E8",X"18",X"9B",X"18",X"5A",
		X"15",X"A3",X"18",X"62",X"15",X"AE",X"18",X"6D",X"15",X"B6",X"18",X"75",X"15",X"C1",X"18",X"80",
		X"15",X"88",X"15",X"8B",X"15",X"8E",X"15",X"C9",X"18",X"CF",X"18",X"D5",X"18",X"1B",X"21",X"1B",
		X"0E",X"11",X"1B",X"22",X"1B",X"0F",X"0B",X"00",X"18",X"04",X"11",X"12",X"1B",X"01",X"14",X"13",
		X"13",X"0E",X"0D",X"07",X"07",X"10",X"90",X"10",X"90",X"23",X"03",X"03",X"03",X"93",X"1C",X"93",
		X"1C",X"40",X"00",X"E0",X"33",X"00",X"07",X"07",X"D0",X"90",X"D0",X"90",X"21",X"B4",X"0A",X"B4",
		X"0A",X"03",X"00",X"80",X"BA",X"70",X"42",X"72",X"0A",X"70",X"42",X"72",X"0A",X"01",X"0E",X"0D",
		X"14",X"12",X"1B",X"24",X"20",X"20",X"20",X"1D",X"26",X"1D",X"29",X"1D",X"2F",X"05",X"23",X"1D",
		X"26",X"FF",X"1B",X"0E",X"0D",X"0B",X"18",X"1B",X"21",X"1B",X"0F",X"0B",X"00",X"18",X"04",X"11",
		X"12",X"1B",X"01",X"14",X"13",X"13",X"0E",X"0D",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"78",
		X"00",X"10",X"00",X"30",X"00",X"F8",X"00",X"F0",X"07",X"E0",X"3F",X"F0",X"07",X"F8",X"00",X"30",
		X"00",X"10",X"00",X"78",X"00",X"00",X"10",X"10",X"08",X"08",X"05",X"CC",X"03",X"F8",X"07",X"F0",
		X"03",X"A8",X"03",X"C0",X"01",X"80",X"09",X"40",X"07",X"00",X"02",X"00",X"01",X"00",X"01",X"00",
		X"01",X"80",X"03",X"80",X"03",X"80",X"03",X"C0",X"07",X"C8",X"27",X"E8",X"2F",X"F8",X"3E",X"48",
		X"24",X"04",X"00",X"08",X"04",X"50",X"08",X"E0",X"19",X"F0",X"0F",X"E0",X"07",X"E0",X"0A",X"C0",
		X"01",X"C8",X"00",X"70",X"01",X"20",X"00",X"00",X"1E",X"00",X"08",X"00",X"0C",X"00",X"1F",X"E0",
		X"0F",X"FC",X"07",X"E0",X"0F",X"00",X"1F",X"00",X"0C",X"00",X"08",X"00",X"1E",X"40",X"00",X"E0",
		X"02",X"90",X"01",X"80",X"03",X"C0",X"15",X"C0",X"0F",X"E0",X"1F",X"C0",X"33",X"A0",X"10",X"10",
		X"08",X"08",X"08",X"24",X"12",X"7C",X"1F",X"F4",X"17",X"E4",X"13",X"E0",X"03",X"C0",X"01",X"C0",
		X"01",X"C0",X"01",X"80",X"00",X"80",X"00",X"80",X"00",X"00",X"04",X"80",X"E0",X"00",X"13",X"80",
		X"03",X"50",X"07",X"E0",X"07",X"F0",X"0F",X"98",X"07",X"10",X"0A",X"20",X"10",X"00",X"20",X"21",
		X"42",X"23",X"36",X"00",X"21",X"3D",X"20",X"36",X"FF",X"C3",X"CC",X"0E",X"12",X"02",X"0E",X"11",
		X"04",X"1C",X"21",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"12",
		X"02",X"0E",X"11",X"04",X"1C",X"22",X"05",X"14",X"04",X"0B",X"02",X"11",X"04",X"03",X"08",X"13",
		X"1B",X"30",X"01",X"C4",X"38",X"06",X"04",X"C7",X"14",X"06",X"04",X"D3",X"14",X"06",X"07",X"CA",
		X"0E",X"06",X"07",X"D3",X"0E",X"06",X"16",X"CA",X"0E",X"06",X"16",X"D3",X"0E",X"06",X"19",X"C7",
		X"14",X"06",X"19",X"D3",X"14",X"06",X"1C",X"C4",X"38",X"06",X"FF",X"02",X"C4",X"1A",X"06",X"05",
		X"C7",X"09",X"06",X"10",X"C7",X"09",X"06",X"07",X"CA",X"07",X"06",X"10",X"CA",X"06",X"06",X"0A",
		X"CD",X"0A",X"06",X"0A",X"D0",X"04",X"06",X"10",X"D0",X"04",X"06",X"0A",X"D3",X"04",X"06",X"10",
		X"D3",X"04",X"06",X"0A",X"D6",X"0A",X"06",X"08",X"D9",X"06",X"06",X"10",X"D9",X"06",X"06",X"05",
		X"DC",X"09",X"06",X"10",X"DC",X"09",X"06",X"02",X"DF",X"1A",X"06",X"FF",X"1F",X"24",X"44",X"24",
		X"1F",X"7F",X"49",X"49",X"49",X"36",X"3E",X"41",X"41",X"41",X"22",X"7F",X"41",X"41",X"41",X"3E",
		X"7F",X"49",X"49",X"49",X"41",X"7F",X"48",X"48",X"48",X"40",X"3E",X"41",X"41",X"45",X"47",X"7F",
		X"08",X"08",X"08",X"7F",X"00",X"41",X"7F",X"41",X"00",X"02",X"01",X"01",X"01",X"7E",X"7F",X"08",
		X"14",X"22",X"41",X"7F",X"01",X"01",X"01",X"01",X"7F",X"20",X"18",X"20",X"7F",X"7F",X"10",X"08",
		X"04",X"7F",X"3E",X"41",X"41",X"41",X"3E",X"7F",X"48",X"48",X"48",X"30",X"3E",X"41",X"45",X"42",
		X"3D",X"7F",X"48",X"4C",X"4A",X"31",X"32",X"49",X"49",X"49",X"26",X"40",X"40",X"7F",X"40",X"40",
		X"7E",X"01",X"01",X"01",X"7E",X"7C",X"02",X"01",X"02",X"7C",X"7F",X"02",X"0C",X"02",X"7F",X"63",
		X"14",X"08",X"14",X"63",X"60",X"10",X"0F",X"10",X"60",X"43",X"45",X"49",X"51",X"61",X"00",X"00",
		X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"22",X"14",X"7F",
		X"14",X"22",X"08",X"14",X"22",X"41",X"00",X"00",X"41",X"22",X"14",X"08",X"3E",X"45",X"49",X"51",
		X"3E",X"00",X"21",X"7F",X"01",X"00",X"23",X"45",X"49",X"49",X"31",X"42",X"41",X"49",X"59",X"66",
		X"0C",X"14",X"24",X"7F",X"04",X"72",X"51",X"51",X"51",X"4E",X"1E",X"29",X"49",X"49",X"46",X"40",
		X"47",X"48",X"50",X"60",X"36",X"49",X"49",X"49",X"36",X"31",X"49",X"49",X"4A",X"3C",X"14",X"14",
		X"14",X"14",X"14",X"01",X"02",X"04",X"08",X"10",X"00",X"00",X"00",X"00",X"00",X"18",X"18",X"18",
		X"18",X"18",X"00",X"00",X"18",X"18",X"00",X"00",X"1F",X"14",X"16",X"09",X"00",X"1E",X"01",X"01",
		X"1E",X"00",X"1F",X"15",X"15",X"0A",X"00",X"00",X"1F",X"15",X"15",X"11",X"00",X"1F",X"08",X"04",
		X"1F",X"00",X"1F",X"11",X"11",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"40",X"0E",X"60",
		X"0C",X"10",X"10",X"00",X"03",X"80",X"07",X"00",X"0F",X"00",X"04",X"00",X"00",X"00",X"20",X"00",
		X"10",X"00",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"60",X"00",
		X"0A",X"00",X"1C",X"00",X"08",X"80",X"01",X"00",X"03",X"40",X"0B",X"80",X"5F",X"00",X"20",X"00",
		X"52",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"1F",X"00",X"16",X"00",X"A0",X"00",X"85",
		X"01",X"12",X"01",X"31",X"00",X"70",X"00",X"42",X"04",X"A4",X"08",X"0E",X"0C",X"0F",X"10",X"18",
		X"00",X"00",X"08",X"00",X"38",X"00",X"44",X"00",X"01",X"02",X"49",X"01",X"D0",X"01",X"54",X"02",
		X"08",X"00",X"84",X"00",X"60",X"00",X"31",X"00",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"18",X"80",X"00",X"40",X"C1",X"21",X"F2",X"03",X"18",X"0A",X"C8",X"18",X"02",X"3B",X"F4",X"46",
		X"24",X"10",X"4C",X"1B",X"40",X"49",X"10",X"00",X"B8",X"46",X"80",X"13",X"01",X"10",X"42",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"90",X"60",X"40",X"08",X"41",X"10",
		X"00",X"10",X"01",X"00",X"00",X"62",X"0D",X"00",X"08",X"F4",X"F8",X"11",X"00",X"38",X"B2",X"02",
		X"60",X"AB",X"C7",X"07",X"40",X"DB",X"DB",X"37",X"00",X"FD",X"3F",X"03",X"80",X"3D",X"FE",X"02",
		X"C1",X"8B",X"7F",X"07",X"E0",X"E7",X"F7",X"0F",X"E0",X"E9",X"FD",X"0F",X"E0",X"EC",X"AE",X"09",
		X"C0",X"DC",X"76",X"0D",X"80",X"8C",X"B9",X"05",X"80",X"2C",X"DF",X"03",X"C0",X"78",X"D3",X"03",
		X"20",X"59",X"EE",X"03",X"90",X"F9",X"FF",X"01",X"80",X"F1",X"C7",X"04",X"84",X"7B",X"17",X"10",
		X"80",X"F7",X"FB",X"02",X"00",X"2F",X"39",X"04",X"00",X"1E",X"1C",X"00",X"00",X"8C",X"01",X"10",
		X"00",X"80",X"00",X"00",X"00",X"80",X"00",X"41",X"10",X"00",X"04",X"C2",X"08",X"80",X"0C",X"00",
		X"1D",X"13",X"00",X"08",X"13",X"0E",X"1B",X"02",X"0E",X"11",X"0F",X"0E",X"11",X"00",X"13",X"08",
		X"0E",X"0D",X"1D",X"08",X"0D",X"12",X"04",X"11",X"13",X"1B",X"02",X"0E",X"08",X"0D",X"00",X"01",
		X"FF",X"00",X"00",X"67",X"1E",X"10",X"00",X"01",X"02",X"00",X"00",X"83",X"1E",X"10",X"00",X"FF",
		X"01",X"00",X"00",X"A1",X"1E",X"10",X"00",X"FF",X"FE",X"00",X"00",X"C0",X"1E",X"10",X"33",X"01",
		X"31",X"01",X"2D",X"01",X"2B",X"01",X"28",X"01",X"26",X"01",X"24",X"01",X"22",X"01",X"20",X"01",
		X"1E",X"01",X"1D",X"01",X"1B",X"01",X"19",X"01",X"00",X"13",X"08",X"0B",X"13",X"CD",X"DB",X"18",
		X"FE",X"03",X"21",X"D0",X"90",X"C2",X"AD",X"0C",X"2A",X"39",X"23",X"C3",X"AD",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"3A");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
