library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity spy_hunter_bg_bits_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of spy_hunter_bg_bits_1 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"FF",X"FF",X"FF",X"FF",X"57",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"D5",X"FF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"7F",X"FF",
		X"FF",X"FF",X"FF",X"3C",X"FF",X"FD",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"F7",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"7F",X"FF",X"FF",X"FF",X"FF",X"F5",X"FF",X"FD",X"DF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"FF",X"FF",X"FF",X"FF",X"DF",
		X"FF",X"FF",X"DD",X"FF",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",X"D7",X"DF",X"FF",X"F7",
		X"FF",X"FD",X"FD",X"FF",X"FD",X"FF",X"FF",X"FD",X"FF",X"FF",X"F5",X"FF",X"FF",X"7F",X"FF",X"FD",
		X"FD",X"FF",X"FF",X"7F",X"FF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"D7",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"FF",X"FF",X"FF",X"FF",X"DF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"FF",X"FF",
		X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"FF",X"FF",X"FF",X"FF",X"DF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"A5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"09",X"96",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"99",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"02",X"65",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"0A",X"69",X"99",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"26",X"66",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"98",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"56",X"68",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"56",X"9A",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"A6",X"80",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"66",X"9A",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"9A",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"10",
		X"00",X"00",X"00",X"00",X"10",X"41",X"00",X"04",X"00",X"04",X"00",X"41",X"00",X"04",X"44",X"11",
		X"41",X"10",X"51",X"00",X"11",X"01",X"15",X"45",X"10",X"11",X"44",X"45",X"05",X"85",X"51",X"55",
		X"44",X"41",X"11",X"44",X"55",X"54",X"55",X"55",X"45",X"14",X"45",X"15",X"51",X"59",X"55",X"55",
		X"11",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"91",X"59",X"59",X"55",X"55",X"59",X"55",
		X"45",X"55",X"55",X"55",X"59",X"55",X"55",X"65",X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"95",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"5D",X"5D",X"55",X"57",X"59",X"55",X"55",X"57",X"55",X"55",X"F7",X"75",
		X"55",X"57",X"57",X"55",X"57",X"77",X"DF",X"DF",X"55",X"75",X"75",X"77",X"DD",X"DF",X"F7",X"7F",
		X"77",X"5F",X"5F",X"7F",X"FF",X"FD",X"F7",X"FF",X"5D",X"F7",X"F7",X"DD",X"F7",X"FF",X"FF",X"FF",
		X"F7",X"7D",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"D7",X"7F",X"F7",X"FF",X"FF",X"FF",X"FF",
		X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7D",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"26",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"02",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"26",X"65",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"02",X"65",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"02",X"66",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"56",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"AA",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"AA",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"A8",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"56",X"A0",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"5A",X"A8",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"A8",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"10",
		X"00",X"00",X"00",X"00",X"10",X"41",X"00",X"04",X"00",X"04",X"00",X"41",X"00",X"04",X"44",X"11",
		X"41",X"10",X"51",X"00",X"11",X"01",X"15",X"45",X"10",X"11",X"44",X"45",X"05",X"85",X"51",X"55",
		X"44",X"41",X"11",X"44",X"55",X"54",X"55",X"55",X"45",X"14",X"45",X"15",X"51",X"59",X"55",X"55",
		X"11",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"91",X"59",X"59",X"55",X"55",X"59",X"55",
		X"45",X"55",X"55",X"55",X"59",X"55",X"55",X"65",X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"95",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"5D",X"5D",X"55",X"57",X"59",X"55",X"55",X"57",X"55",X"55",X"F7",X"75",
		X"55",X"57",X"57",X"55",X"57",X"77",X"DF",X"DF",X"55",X"75",X"75",X"77",X"DD",X"DF",X"F7",X"7F",
		X"77",X"5F",X"5F",X"7F",X"FF",X"FD",X"F7",X"FF",X"5D",X"F7",X"F7",X"DD",X"F7",X"FF",X"FF",X"FF",
		X"F7",X"7D",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"D7",X"7F",X"F7",X"FF",X"FF",X"FF",X"FF",
		X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7D",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"26",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"02",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"26",X"65",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"02",X"65",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"02",X"66",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"56",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"AA",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"AA",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"A8",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"56",X"A0",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"5A",X"A8",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"A8",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"10",
		X"00",X"00",X"00",X"00",X"10",X"41",X"00",X"04",X"00",X"04",X"00",X"41",X"00",X"04",X"44",X"11",
		X"41",X"10",X"51",X"00",X"11",X"01",X"15",X"45",X"10",X"11",X"44",X"45",X"05",X"85",X"51",X"55",
		X"44",X"41",X"11",X"44",X"55",X"54",X"55",X"55",X"45",X"14",X"45",X"15",X"51",X"59",X"55",X"55",
		X"11",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"91",X"59",X"59",X"55",X"55",X"59",X"55",
		X"45",X"55",X"55",X"55",X"59",X"55",X"55",X"65",X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"95",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"5D",X"5D",X"55",X"57",X"59",X"55",X"55",X"57",X"55",X"55",X"F7",X"75",
		X"55",X"57",X"57",X"55",X"57",X"77",X"DF",X"DF",X"55",X"75",X"75",X"77",X"DD",X"DF",X"F7",X"7F",
		X"77",X"5F",X"5F",X"7F",X"FF",X"FD",X"F7",X"FF",X"5D",X"F7",X"F7",X"DD",X"F7",X"FF",X"FF",X"FF",
		X"F7",X"7D",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"D7",X"7F",X"F7",X"FF",X"FF",X"FF",X"FF",
		X"66",X"7F",X"FF",X"FF",X"FF",X"DD",X"5A",X"AA",X"AE",X"BF",X"FF",X"FF",X"FF",X"FD",X"56",X"BA",
		X"AB",X"FF",X"FF",X"FF",X"FF",X"FD",X"56",X"AA",X"AA",X"FF",X"FF",X"FF",X"EF",X"D5",X"56",X"AA",
		X"AB",X"FF",X"FF",X"FF",X"BA",X"DD",X"56",X"BA",X"AF",X"FF",X"FF",X"FF",X"EF",X"F5",X"56",X"9A",
		X"AF",X"EF",X"FF",X"FF",X"FB",X"B6",X"56",X"6A",X"BF",X"FF",X"FF",X"FF",X"FE",X"FD",X"5A",X"AA",
		X"BF",X"EF",X"FF",X"FF",X"FF",X"F9",X"5A",X"AE",X"BF",X"FF",X"EF",X"FF",X"FF",X"BF",X"69",X"AA",
		X"BF",X"FF",X"FE",X"FF",X"FF",X"E5",X"5A",X"EA",X"BF",X"FF",X"FB",X"FF",X"FF",X"66",X"6A",X"AA",
		X"BF",X"FF",X"FE",X"FF",X"FE",X"55",X"A7",X"AA",X"BF",X"FF",X"FF",X"EF",X"BF",X"5A",X"AA",X"AA",
		X"BF",X"FF",X"FF",X"FE",X"7D",X"5A",X"6A",X"AA",X"AF",X"FF",X"FF",X"F9",X"99",X"66",X"AE",X"AA",
		X"AF",X"FF",X"FF",X"E9",X"65",X"5A",X"AA",X"AA",X"AF",X"FF",X"FF",X"EB",X"96",X"6A",X"BA",X"AA",
		X"AF",X"FF",X"FE",X"BA",X"A5",X"9A",X"AA",X"AA",X"AA",X"FF",X"FD",X"7A",X"A5",X"9B",X"AA",X"AA",
		X"AE",X"FF",X"F9",X"96",X"65",X"6A",X"AA",X"AA",X"AA",X"AF",X"DE",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AF",X"D5",X"9A",X"A6",X"6B",X"AA",X"AA",X"AA",X"AF",X"56",X"6A",X"AA",X"6A",X"AA",X"AA",
		X"AA",X"A6",X"65",X"A9",X"A6",X"6A",X"AA",X"AA",X"AA",X"A9",X"56",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"A9",X"96",X"AB",X"AA",X"AE",X"AA",X"AA",X"AA",X"AA",X"A6",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"A6",X"6A",X"EA",X"AA",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AB",X"AA",X"AE",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"BA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AE",X"66",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"95",X"BA",X"AA",X"AA",X"AA",X"AA",X"AA",X"BA",X"56",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"A9",X"56",X"AB",X"EA",X"6E",X"AA",X"AA",X"AB",X"A9",X"95",X"AA",X"A6",X"AB",X"AA",X"AA",
		X"AA",X"A5",X"55",X"6B",X"EA",X"AA",X"AA",X"AA",X"AA",X"97",X"FD",X"6A",X"99",X"AA",X"EA",X"AA",
		X"9A",X"97",X"FD",X"6B",X"A6",X"5A",X"AA",X"6A",X"AA",X"57",X"FD",X"AA",X"A5",X"6A",X"AA",X"AA",
		X"AA",X"7F",X"FF",X"6A",X"A5",X"6A",X"EA",X"AA",X"A9",X"7F",X"FF",X"DA",X"95",X"66",X"AA",X"9A",
		X"AB",X"FF",X"FD",X"D6",X"95",X"6A",X"BA",X"AA",X"A7",X"FF",X"FF",X"DA",X"95",X"5A",X"AA",X"AA",
		X"AF",X"FF",X"FF",X"56",X"5D",X"5A",X"AA",X"9A",X"AD",X"FF",X"FF",X"D6",X"5D",X"56",X"AA",X"AA",
		X"AB",X"FF",X"FF",X"D5",X"5D",X"5A",X"BA",X"9A",X"BF",X"FF",X"FF",X"F5",X"7F",X"56",X"AA",X"AA",
		X"BF",X"FF",X"FF",X"F6",X"7F",X"56",X"AE",X"AA",X"BF",X"FF",X"FF",X"F5",X"FF",X"D6",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FD",X"7F",X"56",X"6A",X"A9",X"FF",X"FF",X"FF",X"FF",X"FF",X"D6",X"AB",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"F7",X"D5",X"AA",X"A9",X"BF",X"FF",X"FF",X"FF",X"FF",X"D5",X"AA",X"AA",
		X"BF",X"FF",X"FF",X"FF",X"FF",X"F5",X"5A",X"AA",X"BF",X"FF",X"FF",X"FF",X"FF",X"F5",X"AA",X"EA",
		X"AF",X"FF",X"FF",X"FF",X"FF",X"D5",X"9A",X"AA",X"AB",X"FF",X"FF",X"FF",X"FF",X"F5",X"5A",X"AA",
		X"AB",X"FF",X"FF",X"FF",X"FF",X"75",X"5A",X"AE",X"AB",X"FF",X"FF",X"FF",X"FF",X"F5",X"56",X"AA",
		X"AA",X"FF",X"BF",X"FF",X"FF",X"F5",X"5A",X"6A",X"AA",X"FF",X"FF",X"FF",X"FF",X"FD",X"56",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"F7",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",
		X"FF",X"FF",X"F7",X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"D7",
		X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",
		X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",X"7F",X"FF",X"FF",X"FD",X"FD",X"FF",X"FF",X"FD",X"FF",
		X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",X"FD",X"F5",X"FF",X"FF",X"FF",X"DF",
		X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",X"DF",X"DF",X"FF",X"FD",X"FF",X"F7",X"FF",X"FD",X"FF",X"FF",
		X"FF",X"FD",X"FF",X"DF",X"FF",X"FD",X"F7",X"FF",X"FF",X"F7",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"F7",X"FF",X"FF",X"FF",X"FF",X"DF",X"7F",X"FF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"9A",X"AA",X"AA",X"AA",X"AA",X"9A",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"A9",X"AA",X"AA",X"AA",X"AA",X"9A",X"AA",X"AA",X"AA",X"AA",X"AA",X"69",X"AA",
		X"AA",X"AA",X"AA",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"6A",
		X"AA",X"A6",X"AA",X"AA",X"AA",X"A9",X"AA",X"AA",X"A6",X"AA",X"9A",X"AA",X"AA",X"9A",X"A6",X"66",
		X"A9",X"9A",X"65",X"A9",X"9A",X"AA",X"69",X"A9",X"55",X"55",X"6A",X"9A",X"A9",X"A6",X"56",X"59",
		X"95",X"56",X"59",X"AA",X"65",X"55",X"55",X"56",X"55",X"59",X"56",X"66",X"99",X"95",X"55",X"55",
		X"55",X"55",X"55",X"AA",X"56",X"56",X"55",X"55",X"55",X"55",X"56",X"66",X"55",X"55",X"65",X"55",
		X"55",X"55",X"55",X"95",X"59",X"59",X"55",X"65",X"55",X"95",X"59",X"59",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"DF",X"FF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",X"D7",X"FF",X"7F",
		X"F7",X"F7",X"F7",X"FD",X"F7",X"D7",X"FF",X"FF",X"FF",X"F7",X"FF",X"FD",X"FF",X"DF",X"7F",X"DF",
		X"FF",X"D7",X"FF",X"FD",X"FF",X"7F",X"FF",X"FF",X"FD",X"5F",X"FF",X"F7",X"FD",X"FF",X"FF",X"FF",
		X"FD",X"7F",X"FF",X"DF",X"F7",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",X"DF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"7F",X"FF",X"F7",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"F7",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"FF",X"FF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"DF",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FD",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"98",
		X"55",X"55",X"55",X"59",X"A6",X"9A",X"00",X"00",X"66",X"69",X"A6",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"A5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"09",X"96",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"99",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"02",X"65",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"0A",X"69",X"99",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"26",X"66",X"55",X"00",X"00",X"00",X"00",X"00",X"09",X"99",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"26",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"98",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"56",X"68",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"56",X"9A",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"A6",X"80",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"66",X"9A",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"9A",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"44",X"50",X"00",X"10",
		X"01",X"10",X"54",X"45",X"15",X"45",X"14",X"45",X"10",X"45",X"21",X"55",X"46",X"55",X"45",X"55",
		X"45",X"54",X"55",X"11",X"55",X"55",X"55",X"65",X"59",X"99",X"55",X"55",X"55",X"95",X"65",X"55",
		X"45",X"59",X"59",X"65",X"65",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",
		X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"59",X"59",X"55",X"55",X"59",X"55",
		X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"D5",X"55",X"D5",X"55",X"55",X"5F",X"55",X"77",X"5D",X"77",X"75",X"DD",
		X"D5",X"D7",X"DD",X"D5",X"F7",X"DF",X"DF",X"57",X"7F",X"7F",X"7F",X"DF",X"7F",X"7D",X"FD",X"DD",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"AA",X"AA",X"9A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"A9",X"AA",X"6A",X"AA",X"AA",X"AA",X"A9",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"6A",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"6A",X"AA",X"6A",X"AA",X"AA",X"AA",X"A9",X"A6",X"A6",X"9A",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"6A",X"AA",X"A6",X"AA",X"AA",X"6A",X"AA",X"99",X"99",X"66",X"6A",
		X"AA",X"AA",X"AA",X"A6",X"69",X"55",X"A9",X"9A",X"AA",X"6A",X"AA",X"AA",X"95",X"55",X"95",X"AA",
		X"AA",X"AA",X"AA",X"99",X"95",X"55",X"56",X"66",X"AA",X"A6",X"AA",X"AA",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"9A",X"A5",X"55",X"55",X"55",X"AA",X"AA",X"9A",X"69",X"55",X"55",X"59",X"55",
		X"AA",X"AA",X"AA",X"A6",X"55",X"55",X"55",X"55",X"9A",X"AA",X"AA",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"A5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"09",X"96",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"99",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"02",X"65",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"0A",X"69",X"99",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"26",X"66",X"55",
		X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",
		X"55",X"79",X"59",X"65",X"65",X"55",X"56",X"55",X"59",X"95",X"55",X"55",X"55",X"95",X"65",X"55",
		X"55",X"57",X"55",X"DD",X"55",X"55",X"55",X"65",X"55",X"55",X"ED",X"55",X"76",X"55",X"57",X"55",
		X"57",X"5F",X"57",X"75",X"D5",X"75",X"55",X"5D",X"5F",X"FD",X"FF",X"FF",X"55",X"5D",X"5D",X"55",
		X"FD",X"FF",X"FF",X"DD",X"FF",X"F5",X"F7",X"77",X"7F",X"DF",X"DF",X"FF",X"FD",X"FF",X"FF",X"FF",
		X"DF",X"FF",X"FF",X"F7",X"DF",X"DF",X"FF",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"98",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"56",X"68",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"56",X"9A",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"A6",X"80",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"66",X"9A",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"9A",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",X"FF",X"F7",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",X"7D",X"FD",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FD",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",X"F7",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"41",X"10",X"00",X"00",X"00",X"00",X"00",
		X"11",X"04",X"45",X"11",X"04",X"00",X"00",X"00",X"40",X"40",X"40",X"10",X"40",X"40",X"00",X"00",
		X"15",X"14",X"11",X"04",X"04",X"00",X"04",X"00",X"45",X"50",X"55",X"44",X"41",X"00",X"40",X"10",
		X"55",X"45",X"05",X"15",X"10",X"44",X"11",X"04",X"14",X"55",X"55",X"44",X"15",X"55",X"45",X"50",
		X"55",X"55",X"55",X"55",X"59",X"50",X"54",X"65",X"55",X"95",X"59",X"59",X"55",X"55",X"48",X"44",
		X"65",X"55",X"55",X"55",X"55",X"55",X"51",X"51",X"D5",X"55",X"55",X"55",X"55",X"59",X"55",X"54",
		X"75",X"79",X"59",X"65",X"65",X"55",X"56",X"55",X"5B",X"99",X"55",X"55",X"55",X"95",X"65",X"55",
		X"77",X"57",X"55",X"DD",X"55",X"55",X"55",X"65",X"FD",X"F5",X"ED",X"55",X"76",X"55",X"55",X"55",
		X"F7",X"7F",X"57",X"75",X"D5",X"75",X"55",X"55",X"FF",X"FD",X"FF",X"FF",X"77",X"5D",X"55",X"55",
		X"FF",X"FF",X"FF",X"DD",X"FF",X"F5",X"F5",X"75",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"5D",X"DD",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"FD",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"75",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"44",X"41",X"10",X"00",X"00",X"00",X"00",X"00",X"11",X"04",X"45",X"11",X"04",X"00",X"00",X"00",
		X"44",X"50",X"40",X"10",X"40",X"40",X"00",X"40",X"15",X"54",X"11",X"04",X"04",X"00",X"04",X"00",
		X"45",X"55",X"55",X"44",X"51",X"14",X"40",X"10",X"55",X"55",X"55",X"15",X"15",X"55",X"11",X"04",
		X"15",X"55",X"55",X"45",X"55",X"55",X"45",X"50",X"55",X"55",X"55",X"55",X"59",X"55",X"54",X"65",
		X"55",X"95",X"59",X"59",X"55",X"55",X"59",X"45",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"D5",X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"75",X"79",X"59",X"65",X"65",X"55",X"56",X"55",
		X"5B",X"99",X"55",X"55",X"55",X"95",X"65",X"55",X"77",X"57",X"55",X"DD",X"55",X"55",X"55",X"65",
		X"FD",X"F5",X"ED",X"55",X"76",X"55",X"55",X"55",X"F7",X"7F",X"57",X"75",X"D5",X"75",X"55",X"55",
		X"FF",X"FD",X"FF",X"FF",X"77",X"5D",X"55",X"55",X"FF",X"FF",X"FF",X"DD",X"FF",X"F5",X"F5",X"75",
		X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"5D",X"DD",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"FD",X"77",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"75",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"9A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A2",
		X"AA",X"AA",X"AA",X"A9",X"AA",X"6A",X"AA",X"AA",X"A9",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"6A",
		X"A9",X"AA",X"A9",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"9A",X"9A",X"6A",X"AA",X"AA",X"AA",
		X"9A",X"AA",X"A9",X"AA",X"AA",X"AA",X"AA",X"AA",X"A9",X"99",X"66",X"66",X"AA",X"A9",X"AA",X"AA",
		X"A6",X"6A",X"55",X"69",X"9A",X"AA",X"AA",X"AA",X"AA",X"56",X"55",X"56",X"AA",X"AA",X"A8",X"AA",
		X"99",X"95",X"55",X"56",X"66",X"AA",X"AA",X"AA",X"55",X"55",X"55",X"55",X"AA",X"AA",X"9A",X"AA",
		X"55",X"55",X"55",X"5A",X"A6",X"AA",X"AA",X"AA",X"55",X"65",X"55",X"55",X"69",X"A6",X"AA",X"AA",
		X"55",X"55",X"55",X"55",X"9A",X"AA",X"AA",X"AA",X"55",X"55",X"55",X"55",X"55",X"AA",X"AA",X"A6",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"41",X"10",X"00",X"00",X"00",X"00",X"00",
		X"11",X"04",X"45",X"11",X"04",X"00",X"00",X"00",X"44",X"50",X"40",X"10",X"40",X"40",X"00",X"40",
		X"15",X"54",X"11",X"04",X"04",X"00",X"04",X"00",X"45",X"55",X"55",X"44",X"51",X"14",X"40",X"10",
		X"55",X"55",X"55",X"15",X"15",X"55",X"11",X"04",X"15",X"55",X"55",X"45",X"55",X"55",X"45",X"50",
		X"55",X"55",X"55",X"55",X"59",X"55",X"54",X"65",X"55",X"95",X"59",X"59",X"55",X"55",X"59",X"45",
		X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"D5",X"55",X"55",X"55",X"55",X"59",X"55",X"55",
		X"75",X"79",X"59",X"65",X"65",X"55",X"56",X"55",X"5B",X"99",X"55",X"55",X"55",X"95",X"65",X"55",
		X"77",X"57",X"55",X"DD",X"55",X"55",X"55",X"65",X"FD",X"F5",X"ED",X"55",X"76",X"55",X"55",X"55",
		X"F7",X"7F",X"57",X"75",X"D5",X"75",X"55",X"55",X"FF",X"FD",X"FF",X"FF",X"77",X"5D",X"55",X"55",
		X"FF",X"FF",X"FF",X"DD",X"FF",X"F5",X"F5",X"75",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"5D",X"DD",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"FD",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"75",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F5",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",
		X"FD",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"FF",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"D7",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"5D",X"FD",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FD",X"FF",X"57",X"FF",X"FF",X"FF",X"FF",X"FF",X"F5",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FD",X"5F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"5F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"5D",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FD",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"DD",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F7",X"7D",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DD",X"F7",X"7D",X"DD",X"FF",X"FF",X"FF",X"FF",
		X"55",X"5F",X"7F",X"DF",X"7F",X"7F",X"FF",X"FF",X"55",X"57",X"DD",X"F7",X"F7",X"FF",X"F7",X"FF",
		X"56",X"55",X"55",X"77",X"5D",X"D7",X"7F",X"DF",X"55",X"55",X"55",X"D5",X"D5",X"55",X"DD",X"F7",
		X"55",X"55",X"55",X"75",X"55",X"75",X"75",X"5F",X"55",X"59",X"55",X"55",X"59",X"55",X"57",X"65",
		X"55",X"95",X"59",X"59",X"55",X"55",X"59",X"77",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"45",X"45",X"59",X"65",X"65",X"55",X"56",X"55",
		X"58",X"99",X"55",X"55",X"55",X"95",X"65",X"55",X"44",X"54",X"55",X"11",X"55",X"55",X"55",X"65",
		X"01",X"05",X"21",X"55",X"46",X"55",X"55",X"55",X"04",X"40",X"54",X"45",X"15",X"45",X"55",X"55",
		X"00",X"00",X"00",X"00",X"44",X"51",X"55",X"55",X"00",X"04",X"04",X"11",X"00",X"05",X"05",X"45",
		X"00",X"00",X"00",X"00",X"01",X"00",X"51",X"11",X"00",X"00",X"00",X"00",X"00",X"10",X"01",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"45",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"DD",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F7",X"7D",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DD",X"F7",X"7D",X"DD",X"FF",X"FF",X"FF",X"FF",
		X"55",X"5F",X"7F",X"DF",X"7F",X"7F",X"FF",X"FF",X"55",X"55",X"DD",X"F7",X"F7",X"FF",X"F7",X"FF",
		X"56",X"55",X"55",X"77",X"5D",X"D7",X"7F",X"DF",X"55",X"55",X"55",X"55",X"D5",X"55",X"DD",X"F7",
		X"55",X"55",X"55",X"55",X"55",X"75",X"75",X"5F",X"55",X"59",X"55",X"55",X"59",X"55",X"57",X"65",
		X"55",X"95",X"59",X"59",X"55",X"55",X"59",X"77",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"45",X"55",X"59",X"65",X"65",X"55",X"56",X"55",
		X"58",X"99",X"55",X"55",X"55",X"95",X"65",X"55",X"44",X"54",X"55",X"11",X"55",X"55",X"55",X"65",
		X"01",X"05",X"21",X"55",X"46",X"55",X"55",X"55",X"04",X"40",X"54",X"45",X"15",X"45",X"55",X"55",
		X"00",X"00",X"00",X"00",X"44",X"51",X"55",X"55",X"00",X"04",X"04",X"11",X"00",X"05",X"05",X"45",
		X"00",X"00",X"00",X"00",X"01",X"00",X"51",X"11",X"00",X"00",X"00",X"00",X"00",X"10",X"01",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"45",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"9A",X"9A",X"AA",X"AA",X"9A",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"AA",X"69",X"AA",X"AA",X"9A",
		X"AA",X"AA",X"AA",X"AA",X"A6",X"A9",X"AA",X"AA",X"AA",X"9A",X"A9",X"A9",X"5A",X"6A",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"A5",X"55",X"AA",X"AA",X"6A",X"A9",X"AA",X"66",X"55",X"55",X"56",X"9A",X"AA",
		X"9A",X"9A",X"A9",X"99",X"59",X"9A",X"AA",X"9A",X"55",X"56",X"56",X"55",X"55",X"56",X"99",X"AA",
		X"A5",X"65",X"55",X"55",X"55",X"55",X"69",X"6A",X"55",X"95",X"95",X"55",X"59",X"55",X"5A",X"55",
		X"59",X"55",X"55",X"55",X"55",X"59",X"65",X"56",X"95",X"55",X"56",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"65",X"55",X"95",X"59",X"59",X"55",X"55",X"55",X"55",
		X"59",X"99",X"55",X"55",X"55",X"95",X"65",X"55",X"54",X"54",X"55",X"11",X"55",X"55",X"55",X"65",
		X"01",X"05",X"21",X"55",X"46",X"55",X"55",X"55",X"44",X"40",X"54",X"45",X"15",X"45",X"55",X"55",
		X"00",X"00",X"00",X"00",X"44",X"51",X"55",X"55",X"01",X"04",X"04",X"11",X"00",X"05",X"05",X"45",
		X"00",X"00",X"00",X"00",X"01",X"00",X"51",X"11",X"00",X"00",X"00",X"00",X"00",X"10",X"01",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"45",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"7D",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"DD",X"F7",X"7D",X"DD",X"FF",X"FF",X"FF",X"FF",X"55",X"5F",X"7F",X"DF",X"7F",X"7F",X"FF",X"FF",
		X"55",X"55",X"DD",X"F7",X"F7",X"FF",X"F7",X"FF",X"56",X"55",X"55",X"77",X"5D",X"D7",X"7F",X"DF",
		X"55",X"55",X"55",X"55",X"D5",X"55",X"DD",X"F7",X"55",X"55",X"55",X"55",X"55",X"75",X"75",X"5F",
		X"55",X"59",X"55",X"55",X"59",X"55",X"57",X"65",X"55",X"95",X"59",X"59",X"55",X"55",X"59",X"77",
		X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",
		X"45",X"55",X"59",X"65",X"65",X"55",X"56",X"55",X"59",X"99",X"55",X"55",X"55",X"95",X"65",X"55",
		X"54",X"54",X"55",X"11",X"55",X"55",X"55",X"65",X"01",X"05",X"21",X"55",X"46",X"55",X"55",X"55",
		X"44",X"40",X"54",X"45",X"15",X"45",X"55",X"55",X"00",X"00",X"00",X"00",X"44",X"51",X"55",X"55",
		X"01",X"04",X"04",X"11",X"00",X"05",X"05",X"45",X"00",X"00",X"00",X"00",X"01",X"00",X"51",X"11",
		X"00",X"00",X"00",X"00",X"00",X"10",X"01",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"45",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"7D",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"D7",X"7D",X"DD",X"F7",X"FF",X"FF",X"FF",X"55",X"57",X"77",X"DF",X"7F",X"7F",X"FF",X"FF",
		X"55",X"55",X"D5",X"77",X"F7",X"FF",X"F7",X"FF",X"56",X"55",X"55",X"57",X"5D",X"D7",X"7F",X"DF",
		X"55",X"55",X"55",X"55",X"D5",X"55",X"DD",X"F7",X"55",X"55",X"55",X"55",X"55",X"75",X"75",X"5F",
		X"55",X"59",X"55",X"55",X"59",X"55",X"57",X"65",X"55",X"95",X"59",X"59",X"55",X"55",X"59",X"77",
		X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",
		X"55",X"55",X"59",X"65",X"65",X"55",X"56",X"55",X"59",X"99",X"55",X"55",X"55",X"95",X"65",X"55",
		X"14",X"54",X"55",X"55",X"55",X"55",X"55",X"65",X"45",X"05",X"21",X"55",X"56",X"55",X"55",X"55",
		X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",
		X"75",X"79",X"59",X"65",X"65",X"55",X"56",X"55",X"5B",X"99",X"55",X"55",X"55",X"95",X"65",X"55",
		X"57",X"57",X"55",X"DD",X"55",X"55",X"55",X"65",X"55",X"D5",X"ED",X"55",X"76",X"55",X"55",X"55",
		X"57",X"5F",X"57",X"75",X"D5",X"75",X"55",X"55",X"5F",X"FD",X"FF",X"FF",X"77",X"5D",X"55",X"55",
		X"FF",X"7F",X"FF",X"DD",X"FF",X"F5",X"F5",X"75",X"F7",X"FF",X"DF",X"FF",X"FD",X"FF",X"5D",X"DD",
		X"7F",X"FF",X"FF",X"FF",X"FF",X"DF",X"FD",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"75",
		X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"40",X"40",X"40",X"10",X"00",X"41",X"01",X"01",X"11",X"04",X"11",X"04",X"04",X"10",X"10",X"44",
		X"44",X"10",X"50",X"44",X"41",X"00",X"44",X"11",X"45",X"45",X"05",X"11",X"10",X"44",X"11",X"05",
		X"15",X"55",X"55",X"44",X"15",X"51",X"55",X"54",X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"65",
		X"55",X"95",X"59",X"59",X"55",X"55",X"59",X"55",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"55",X"59",X"59",X"65",X"65",X"55",X"56",X"55",
		X"59",X"99",X"55",X"55",X"55",X"95",X"65",X"55",X"75",X"55",X"55",X"DD",X"55",X"55",X"55",X"65",
		X"D7",X"75",X"ED",X"55",X"76",X"55",X"75",X"55",X"DD",X"D7",X"57",X"75",X"D5",X"75",X"D7",X"75",
		X"FD",X"75",X"F7",X"DF",X"77",X"5F",X"7D",X"DF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"55",X"57",X"77",X"DF",X"7F",X"7F",X"FF",X"FF",X"55",X"55",X"55",X"77",X"F7",X"FF",X"F7",X"FF",
		X"56",X"55",X"55",X"57",X"5D",X"D7",X"7F",X"FF",X"55",X"55",X"55",X"55",X"D5",X"55",X"DD",X"F7",
		X"55",X"55",X"55",X"55",X"55",X"75",X"75",X"5F",X"55",X"59",X"55",X"55",X"59",X"55",X"57",X"65",
		X"55",X"95",X"59",X"59",X"55",X"55",X"59",X"77",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"55",X"55",X"59",X"65",X"65",X"55",X"56",X"55",
		X"59",X"99",X"55",X"55",X"55",X"95",X"65",X"55",X"14",X"54",X"55",X"55",X"55",X"55",X"55",X"65",
		X"45",X"05",X"21",X"55",X"56",X"55",X"55",X"55",X"04",X"40",X"54",X"45",X"55",X"55",X"55",X"55",
		X"00",X"00",X"01",X"04",X"54",X"55",X"55",X"55",X"11",X"04",X"04",X"11",X"10",X"45",X"45",X"55",
		X"00",X"10",X"00",X"00",X"01",X"00",X"51",X"55",X"00",X"00",X"00",X"40",X"10",X"11",X"05",X"54",
		X"00",X"00",X"00",X"00",X"01",X"00",X"11",X"45",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"15",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"6A",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A9",X"9A",X"66",X"66",
		X"AA",X"AA",X"AA",X"99",X"9A",X"AA",X"A9",X"A9",X"AA",X"AA",X"AA",X"9A",X"A9",X"A6",X"56",X"99",
		X"AA",X"AA",X"59",X"AA",X"65",X"56",X"65",X"56",X"AA",X"A9",X"66",X"66",X"99",X"95",X"56",X"65",
		X"AA",X"9A",X"69",X"9A",X"56",X"66",X"95",X"55",X"AA",X"65",X"59",X"66",X"65",X"55",X"65",X"55",
		X"AA",X"96",X"66",X"55",X"59",X"5A",X"55",X"65",X"A9",X"95",X"59",X"59",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"57",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"5F",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"5D",X"DF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"7D",X"DF",X"7F",X"FF",X"FF",X"FF",X"FF",X"55",X"55",X"5D",X"DD",X"F7",X"FF",X"FF",X"FF",
		X"65",X"55",X"55",X"5F",X"7F",X"77",X"FF",X"FF",X"55",X"55",X"95",X"57",X"F7",X"FF",X"F7",X"FF",
		X"56",X"55",X"55",X"57",X"5D",X"D7",X"7F",X"FF",X"55",X"55",X"55",X"95",X"55",X"55",X"DD",X"F7",
		X"55",X"55",X"55",X"55",X"55",X"55",X"75",X"5F",X"55",X"59",X"55",X"55",X"59",X"55",X"57",X"65",
		X"55",X"95",X"59",X"59",X"55",X"55",X"59",X"77",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"15",X"55",X"55",X"55",X"59",X"55",X"55",X"51",X"55",X"59",X"65",X"65",X"55",X"56",X"55",
		X"05",X"51",X"45",X"55",X"55",X"95",X"65",X"55",X"04",X"44",X"55",X"15",X"55",X"55",X"55",X"65",
		X"00",X"05",X"21",X"55",X"56",X"55",X"55",X"55",X"00",X"40",X"54",X"45",X"55",X"55",X"55",X"55",
		X"00",X"00",X"01",X"04",X"54",X"55",X"55",X"55",X"00",X"00",X"04",X"11",X"10",X"45",X"45",X"55",
		X"00",X"00",X"00",X"00",X"01",X"00",X"51",X"55",X"00",X"00",X"00",X"40",X"10",X"11",X"05",X"54",
		X"00",X"00",X"00",X"00",X"01",X"00",X"11",X"45",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"15",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"41",X"10",X"04",X"00",X"00",X"00",X"00",
		X"11",X"04",X"45",X"11",X"04",X"04",X"00",X"00",X"44",X"50",X"44",X"10",X"50",X"41",X"01",X"01",
		X"15",X"15",X"11",X"44",X"05",X"10",X"10",X"44",X"55",X"55",X"55",X"44",X"41",X"41",X"44",X"11",
		X"55",X"55",X"55",X"55",X"14",X"54",X"51",X"05",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"54",
		X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"65",X"55",X"95",X"59",X"59",X"55",X"55",X"59",X"55",
		X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",
		X"75",X"59",X"59",X"65",X"65",X"55",X"56",X"55",X"59",X"99",X"55",X"55",X"55",X"95",X"65",X"55",
		X"75",X"57",X"55",X"DD",X"55",X"55",X"55",X"67",X"DF",X"75",X"ED",X"55",X"76",X"55",X"75",X"55",
		X"FD",X"DF",X"57",X"75",X"D5",X"75",X"D7",X"75",X"FF",X"FD",X"FD",X"FF",X"77",X"5D",X"FD",X"DF",
		X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",X"DF",X"7D",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"59",X"55",X"55",X"55",X"55",X"55",X"55",X"A5",X"55",X"55",X"55",X"55",X"59",X"55",X"55",
		X"A9",X"99",X"59",X"65",X"65",X"55",X"56",X"55",X"A9",X"59",X"55",X"55",X"55",X"95",X"65",X"55",
		X"A5",X"65",X"55",X"DD",X"55",X"55",X"55",X"65",X"A6",X"55",X"55",X"55",X"76",X"55",X"57",X"55",
		X"A9",X"55",X"57",X"75",X"D5",X"75",X"55",X"5D",X"95",X"55",X"55",X"FF",X"55",X"5D",X"5D",X"55",
		X"A5",X"55",X"FF",X"DD",X"FF",X"F5",X"F7",X"77",X"95",X"55",X"5D",X"FF",X"FD",X"FF",X"7F",X"FF",
		X"A5",X"55",X"57",X"77",X"DF",X"DF",X"FF",X"77",X"95",X"5F",X"7D",X"FF",X"FF",X"FF",X"F7",X"FF",
		X"95",X"77",X"DF",X"F7",X"F7",X"FF",X"FF",X"7F",X"55",X"DD",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"7F",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"57",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"59",X"55",X"55",X"59",X"55",X"57",X"65",X"55",X"95",X"59",X"59",X"55",X"55",X"59",X"77",
		X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",
		X"55",X"55",X"59",X"65",X"65",X"55",X"56",X"55",X"59",X"99",X"55",X"55",X"55",X"95",X"65",X"55",
		X"14",X"54",X"55",X"55",X"55",X"55",X"55",X"65",X"45",X"05",X"21",X"55",X"56",X"55",X"55",X"55",
		X"04",X"40",X"54",X"45",X"55",X"55",X"55",X"55",X"00",X"00",X"01",X"04",X"54",X"55",X"55",X"55",
		X"11",X"04",X"04",X"11",X"10",X"45",X"45",X"55",X"00",X"10",X"00",X"00",X"01",X"00",X"51",X"55",
		X"00",X"00",X"00",X"40",X"10",X"11",X"05",X"54",X"00",X"00",X"00",X"00",X"01",X"00",X"11",X"45",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"56",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"AA",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"AA",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"A8",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"56",X"A0",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"5A",X"A8",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"A8",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"DD",X"D5",X"55",X"55",X"55",X"55",X"55",X"55",
		X"65",X"57",X"55",X"55",X"55",X"55",X"55",X"55",X"FE",X"ED",X"55",X"D5",X"55",X"55",X"55",X"55",
		X"F7",X"F6",X"ED",X"55",X"55",X"55",X"55",X"55",X"FF",X"DF",X"F6",X"DD",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"F9",X"DD",X"55",X"55",X"55",X"FE",X"FF",X"BF",X"DF",X"95",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"F7",X"79",X"D5",X"55",X"55",X"FF",X"FF",X"FF",X"FF",X"D5",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"FF",
		X"FF",X"FF",X"FF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",X"DF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"69",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"A6",X"AA",X"AA",X"AA",X"AA",X"9A",X"A9",X"AA",X"AA",X"6A",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"A6",X"5A",X"AA",X"AA",X"AA",X"A9",X"AA",X"66",X"66",X"AA",X"A6",X"AA",X"AA",
		X"9A",X"9A",X"A9",X"99",X"59",X"9A",X"AA",X"AA",X"55",X"56",X"56",X"55",X"95",X"56",X"AA",X"AA",
		X"A5",X"65",X"65",X"96",X"55",X"AA",X"6A",X"AA",X"55",X"95",X"95",X"59",X"59",X"65",X"9A",X"AA",
		X"59",X"55",X"55",X"55",X"55",X"AA",X"A9",X"AA",X"95",X"55",X"56",X"55",X"65",X"99",X"6A",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"55",X"5A",X"66",X"55",X"55",X"55",X"55",X"55",X"59",X"6A",X"AA",
		X"55",X"55",X"55",X"55",X"59",X"95",X"66",X"5A",X"55",X"95",X"59",X"59",X"55",X"55",X"55",X"A6",
		X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"AA",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"56",X"AA",X"A0",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"5A",X"AA",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"08",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"D5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"DE",X"D9",X"55",X"55",X"55",X"55",X"55",X"55",X"FF",X"FD",X"95",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"F7",X"FB",X"B5",X"55",X"55",X"55",X"55",X"EF",X"FF",X"FD",X"DE",X"D5",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FB",X"55",X"55",X"55",X"FF",X"FF",X"EF",X"FF",X"FF",X"ED",X"D5",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"97",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"AA",X"55",X"55",X"55",X"55",X"55",X"59",X"59",X"A6",
		X"75",X"79",X"59",X"65",X"65",X"55",X"96",X"9A",X"5B",X"99",X"55",X"55",X"55",X"95",X"69",X"59",
		X"57",X"57",X"55",X"DD",X"55",X"55",X"55",X"65",X"55",X"D5",X"ED",X"55",X"76",X"55",X"55",X"99",
		X"57",X"5F",X"57",X"75",X"D5",X"75",X"55",X"55",X"5F",X"FD",X"FF",X"FF",X"77",X"5D",X"59",X"65",
		X"FF",X"7F",X"FF",X"DD",X"FF",X"F5",X"F5",X"55",X"F7",X"FF",X"DF",X"FF",X"FD",X"FF",X"5D",X"55",
		X"7F",X"FF",X"FF",X"FF",X"FF",X"DF",X"F5",X"57",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"DD",X"55",
		X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DD",X"57",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"D5",
		X"FF",X"FF",X"FF",X"E5",X"55",X"55",X"55",X"55",X"FF",X"FF",X"FF",X"F9",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FD",X"55",X"55",X"55",X"55",X"FF",X"FF",X"FF",X"FE",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"55",X"55",X"55",X"55",X"FF",X"FF",X"FF",X"FF",X"95",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"F5",X"55",X"55",X"55",X"FF",X"FF",X"FF",X"FF",X"F9",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"D5",X"55",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"E5",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"55",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F5",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AB",X"DA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AB",X"F6",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"FD",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"BF",X"D6",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AF",X"FD",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EF",X"DA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AF",X"F5",X"AA",X"AA",X"AA",X"AA",X"AF",X"6A",X"AA",X"FF",X"5A",X"AA",X"AA",
		X"AA",X"BD",X"6A",X"AA",X"AF",X"F5",X"55",X"55",X"AA",X"F5",X"AA",X"AA",X"AF",X"EF",X"FF",X"FE",
		X"2F",X"F6",X"AA",X"AA",X"AA",X"AF",X"FF",X"FE",X"BD",X"DA",X"AA",X"AA",X"AA",X"AA",X"AB",X"6A",
		X"A6",X"DA",X"AA",X"AA",X"AA",X"AA",X"AB",X"2A",X"AA",X"DA",X"AA",X"AA",X"AA",X"AA",X"AB",X"6A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"41",X"10",X"00",X"00",X"00",X"00",X"00",X"11",X"04",X"45",X"11",X"04",X"00",X"00",X"00",
		X"40",X"40",X"40",X"10",X"40",X"41",X"01",X"01",X"15",X"14",X"11",X"04",X"04",X"10",X"10",X"44",
		X"45",X"50",X"55",X"44",X"41",X"00",X"44",X"11",X"55",X"45",X"05",X"15",X"10",X"44",X"11",X"05",
		X"14",X"55",X"55",X"44",X"15",X"55",X"55",X"54",X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"65",
		X"55",X"95",X"59",X"59",X"55",X"55",X"59",X"55",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"75",X"59",X"59",X"65",X"65",X"55",X"56",X"55",
		X"59",X"99",X"55",X"55",X"55",X"95",X"65",X"55",X"75",X"57",X"55",X"DD",X"55",X"55",X"55",X"65",
		X"DF",X"75",X"ED",X"55",X"76",X"55",X"75",X"55",X"FD",X"DF",X"57",X"75",X"D5",X"75",X"D7",X"75",
		X"FF",X"FD",X"FF",X"FF",X"77",X"5F",X"FF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"41",X"10",X"00",X"00",X"00",X"00",X"00",X"11",X"04",X"45",X"11",X"04",X"00",X"00",X"00",
		X"40",X"40",X"40",X"10",X"40",X"41",X"01",X"01",X"15",X"14",X"11",X"04",X"04",X"10",X"10",X"44",
		X"45",X"50",X"55",X"44",X"41",X"00",X"44",X"11",X"55",X"45",X"05",X"15",X"10",X"44",X"11",X"05",
		X"14",X"55",X"55",X"44",X"15",X"55",X"55",X"54",X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"65",
		X"55",X"95",X"59",X"59",X"55",X"55",X"59",X"55",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"75",X"59",X"59",X"65",X"65",X"55",X"56",X"55",
		X"59",X"99",X"55",X"55",X"55",X"95",X"65",X"55",X"75",X"57",X"55",X"DD",X"55",X"55",X"55",X"65",
		X"DF",X"75",X"ED",X"55",X"76",X"55",X"75",X"55",X"FD",X"DF",X"57",X"75",X"D5",X"75",X"D7",X"75",
		X"FF",X"FD",X"FF",X"FF",X"77",X"5F",X"FF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"41",X"10",X"00",X"00",X"00",X"00",X"00",
		X"11",X"04",X"45",X"11",X"04",X"00",X"00",X"00",X"40",X"40",X"40",X"10",X"40",X"41",X"01",X"01",
		X"15",X"14",X"11",X"04",X"04",X"10",X"10",X"44",X"45",X"50",X"55",X"44",X"41",X"00",X"44",X"11",
		X"55",X"45",X"05",X"15",X"10",X"44",X"11",X"05",X"14",X"55",X"55",X"44",X"15",X"55",X"55",X"54",
		X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"65",X"55",X"95",X"59",X"59",X"55",X"55",X"59",X"55",
		X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",
		X"75",X"59",X"59",X"65",X"65",X"55",X"56",X"55",X"59",X"99",X"55",X"55",X"55",X"95",X"65",X"55",
		X"75",X"57",X"55",X"DD",X"55",X"55",X"55",X"67",X"DF",X"75",X"ED",X"55",X"76",X"55",X"75",X"57",
		X"FD",X"DF",X"57",X"75",X"D5",X"75",X"D7",X"77",X"FF",X"FD",X"FF",X"FF",X"77",X"5F",X"FF",X"DF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"FF",X"FF",X"FF",X"FF",X"F7",
		X"FF",X"FF",X"DF",X"FB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FD",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"D7",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FD",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"FF",X"7F",X"FF",
		X"FF",X"FF",X"DF",X"FF",X"F5",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"5F",X"FF",X"FF",
		X"FF",X"FD",X"7F",X"FF",X"FF",X"F5",X"55",X"55",X"FF",X"F5",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",
		X"F7",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"AA",X"DA",X"AA",X"AA",X"AA",X"AA",X"AB",X"6A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"41",X"10",X"00",X"00",X"00",X"00",X"00",
		X"11",X"04",X"45",X"11",X"04",X"00",X"00",X"00",X"40",X"40",X"40",X"10",X"40",X"41",X"01",X"01",
		X"15",X"14",X"11",X"04",X"04",X"10",X"10",X"44",X"45",X"50",X"55",X"44",X"41",X"00",X"44",X"11",
		X"55",X"45",X"05",X"15",X"10",X"44",X"11",X"05",X"14",X"55",X"55",X"44",X"15",X"55",X"55",X"54",
		X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"65",X"55",X"95",X"59",X"59",X"55",X"55",X"59",X"55",
		X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",
		X"75",X"59",X"59",X"65",X"65",X"55",X"56",X"55",X"59",X"99",X"55",X"55",X"55",X"95",X"65",X"55",
		X"75",X"57",X"55",X"DD",X"55",X"55",X"55",X"67",X"DF",X"75",X"ED",X"55",X"76",X"55",X"75",X"57",
		X"FD",X"DF",X"57",X"75",X"D5",X"75",X"D7",X"77",X"FF",X"FD",X"FF",X"FF",X"77",X"5F",X"FF",X"DF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FD",X"D5",X"55",X"55",X"55",X"55",X"59",X"AA",X"F7",X"5D",X"55",X"55",X"55",X"55",X"56",X"6A",
		X"DD",X"D5",X"55",X"55",X"55",X"55",X"99",X"9A",X"F7",X"55",X"D5",X"55",X"55",X"55",X"56",X"6A",
		X"7F",X"55",X"55",X"D5",X"55",X"55",X"56",X"AA",X"FD",X"DD",X"55",X"55",X"55",X"59",X"59",X"A6",
		X"F7",X"55",X"55",X"55",X"55",X"55",X"96",X"6A",X"DD",X"D5",X"55",X"55",X"55",X"55",X"59",X"AA",
		X"FF",X"57",X"55",X"55",X"55",X"55",X"56",X"A6",X"F7",X"55",X"5D",X"55",X"55",X"55",X"96",X"AA",
		X"DD",X"D5",X"55",X"55",X"55",X"55",X"59",X"9A",X"77",X"5D",X"55",X"55",X"55",X"55",X"56",X"6A",
		X"FD",X"D5",X"75",X"55",X"55",X"59",X"59",X"A6",X"F7",X"55",X"55",X"55",X"55",X"55",X"56",X"7A",
		X"DF",X"55",X"55",X"55",X"55",X"55",X"96",X"AA",X"FD",X"D7",X"55",X"55",X"55",X"55",X"59",X"A6",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"41",X"10",X"00",X"00",X"00",X"00",X"00",
		X"11",X"04",X"45",X"11",X"04",X"00",X"00",X"00",X"40",X"40",X"40",X"10",X"40",X"41",X"01",X"01",
		X"15",X"14",X"11",X"04",X"04",X"10",X"10",X"44",X"45",X"50",X"55",X"44",X"41",X"00",X"44",X"11",
		X"55",X"45",X"05",X"15",X"10",X"44",X"11",X"05",X"14",X"55",X"55",X"44",X"15",X"55",X"55",X"54",
		X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"65",X"55",X"95",X"59",X"59",X"55",X"55",X"59",X"55",
		X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",
		X"75",X"59",X"59",X"65",X"65",X"55",X"56",X"55",X"59",X"99",X"55",X"55",X"55",X"95",X"65",X"55",
		X"75",X"57",X"55",X"DD",X"55",X"55",X"55",X"67",X"DF",X"75",X"ED",X"55",X"76",X"55",X"75",X"55",
		X"FD",X"DF",X"57",X"75",X"D5",X"75",X"D7",X"75",X"FF",X"FD",X"FF",X"FF",X"77",X"5F",X"FF",X"DF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F7",X"55",X"55",X"D5",X"55",X"55",X"56",X"6A",X"7D",X"DD",X"55",X"55",X"55",X"55",X"59",X"9A",
		X"F7",X"55",X"55",X"55",X"55",X"56",X"66",X"AA",X"DF",X"55",X"D5",X"55",X"55",X"55",X"56",X"66",
		X"FD",X"DD",X"55",X"55",X"55",X"55",X"59",X"AA",X"F7",X"55",X"57",X"55",X"55",X"55",X"66",X"6A",
		X"DD",X"D5",X"55",X"55",X"55",X"65",X"59",X"AA",X"F7",X"57",X"55",X"55",X"55",X"55",X"56",X"6A",
		X"F7",X"55",X"55",X"55",X"55",X"55",X"96",X"9A",X"FD",X"D5",X"75",X"55",X"55",X"55",X"59",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5A",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FD",X"D5",X"55",X"55",X"55",X"55",X"A7",X"AA",
		X"FC",X"D5",X"55",X"55",X"55",X"55",X"A7",X"AA",X"A9",X"EA",X"AA",X"AA",X"AA",X"AA",X"A7",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"41",X"10",X"00",X"00",X"00",X"00",X"00",
		X"11",X"04",X"45",X"11",X"04",X"00",X"00",X"00",X"40",X"40",X"40",X"10",X"40",X"41",X"01",X"01",
		X"15",X"14",X"11",X"04",X"04",X"10",X"10",X"44",X"45",X"50",X"55",X"44",X"41",X"00",X"44",X"11",
		X"55",X"45",X"05",X"15",X"10",X"44",X"11",X"05",X"14",X"55",X"55",X"44",X"15",X"55",X"55",X"54",
		X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"65",X"55",X"95",X"59",X"59",X"55",X"55",X"59",X"55",
		X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",
		X"75",X"59",X"59",X"65",X"65",X"55",X"56",X"55",X"59",X"99",X"55",X"55",X"55",X"95",X"65",X"55",
		X"75",X"57",X"55",X"DD",X"55",X"55",X"55",X"67",X"DF",X"75",X"ED",X"55",X"76",X"55",X"75",X"55",
		X"FD",X"DF",X"57",X"75",X"D5",X"75",X"D7",X"75",X"FF",X"FD",X"FF",X"FF",X"77",X"5F",X"FF",X"DF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"95",X"55",X"55",X"55",X"55",X"AA",X"AA",X"AA",X"95",X"55",X"55",X"55",X"45",
		X"AA",X"9A",X"6A",X"65",X"55",X"55",X"65",X"65",X"AA",X"AA",X"A6",X"95",X"55",X"65",X"55",X"15",
		X"AA",X"AA",X"A9",X"55",X"55",X"55",X"55",X"55",X"AA",X"9A",X"66",X"55",X"55",X"55",X"D5",X"75",
		X"A9",X"A6",X"99",X"55",X"55",X"55",X"57",X"55",X"AA",X"A9",X"56",X"55",X"65",X"55",X"55",X"77",
		X"AA",X"A6",X"55",X"55",X"55",X"55",X"55",X"5D",X"A9",X"A9",X"55",X"55",X"55",X"59",X"77",X"55",
		X"AA",X"A5",X"95",X"55",X"55",X"55",X"55",X"75",X"9A",X"99",X"55",X"55",X"55",X"5D",X"75",X"DD",
		X"AA",X"95",X"55",X"55",X"55",X"55",X"57",X"77",X"AA",X"95",X"55",X"55",X"55",X"55",X"D5",X"DF",
		X"AA",X"65",X"95",X"55",X"56",X"55",X"57",X"77",X"AA",X"96",X"55",X"55",X"55",X"5D",X"75",X"FF",
		X"51",X"11",X"04",X"11",X"10",X"00",X"00",X"00",X"55",X"55",X"10",X"40",X"01",X"10",X"00",X"00",
		X"55",X"55",X"55",X"04",X"50",X"40",X"10",X"00",X"55",X"55",X"54",X"51",X"04",X"04",X"00",X"00",
		X"55",X"55",X"55",X"14",X"51",X"40",X"41",X"00",X"55",X"55",X"55",X"55",X"04",X"04",X"00",X"04",
		X"55",X"55",X"55",X"51",X"10",X"40",X"10",X"00",X"55",X"55",X"55",X"55",X"51",X"11",X"01",X"00",
		X"55",X"55",X"55",X"55",X"04",X"00",X"00",X"10",X"55",X"55",X"55",X"54",X"51",X"10",X"00",X"00",
		X"55",X"55",X"55",X"55",X"10",X"41",X"04",X"41",X"55",X"55",X"55",X"10",X"44",X"10",X"00",X"00",
		X"55",X"55",X"54",X"45",X"01",X"00",X"40",X"00",X"55",X"55",X"51",X"14",X"10",X"00",X"04",X"00",
		X"55",X"55",X"14",X"41",X"44",X"44",X"00",X"00",X"11",X"11",X"04",X"04",X"10",X"00",X"00",X"00",
		X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"41",X"10",X"00",X"00",X"00",X"00",X"00",
		X"11",X"04",X"45",X"11",X"04",X"00",X"00",X"00",X"40",X"40",X"40",X"10",X"40",X"41",X"01",X"01",
		X"15",X"14",X"11",X"04",X"04",X"10",X"10",X"44",X"45",X"50",X"55",X"44",X"41",X"00",X"44",X"11",
		X"55",X"45",X"05",X"15",X"10",X"44",X"11",X"05",X"14",X"55",X"55",X"44",X"15",X"55",X"55",X"54",
		X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"65",X"55",X"95",X"59",X"59",X"55",X"55",X"59",X"55",
		X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",
		X"75",X"59",X"59",X"65",X"65",X"55",X"56",X"55",X"59",X"99",X"55",X"55",X"55",X"95",X"65",X"55",
		X"75",X"57",X"55",X"DD",X"55",X"55",X"55",X"67",X"DF",X"75",X"ED",X"55",X"76",X"55",X"75",X"55",
		X"AA",X"65",X"55",X"55",X"55",X"55",X"57",X"7F",X"A9",X"95",X"55",X"55",X"55",X"55",X"75",X"DF",
		X"A6",X"66",X"55",X"55",X"55",X"55",X"57",X"77",X"A9",X"95",X"55",X"55",X"55",X"57",X"55",X"DF",
		X"AA",X"95",X"55",X"55",X"57",X"55",X"55",X"FD",X"9A",X"65",X"65",X"55",X"55",X"55",X"77",X"7F",
		X"A9",X"96",X"55",X"55",X"55",X"55",X"55",X"DF",X"AA",X"65",X"55",X"55",X"55",X"55",X"57",X"77",
		X"9A",X"95",X"55",X"55",X"55",X"55",X"D5",X"FF",X"AA",X"96",X"55",X"55",X"55",X"75",X"55",X"DF",
		X"A6",X"65",X"55",X"55",X"55",X"55",X"57",X"77",X"A9",X"95",X"55",X"55",X"55",X"55",X"75",X"DD",
		X"9A",X"65",X"65",X"55",X"55",X"5D",X"57",X"7F",X"A9",X"95",X"55",X"55",X"55",X"55",X"55",X"DF",
		X"AA",X"96",X"55",X"55",X"55",X"55",X"55",X"F7",X"9A",X"65",X"55",X"55",X"55",X"55",X"D7",X"7F",
		X"A9",X"95",X"55",X"55",X"57",X"55",X"55",X"DF",X"A6",X"65",X"55",X"55",X"55",X"55",X"77",X"7D",
		X"AA",X"99",X"95",X"55",X"55",X"55",X"55",X"DF",X"99",X"95",X"55",X"55",X"55",X"57",X"55",X"F7",
		X"AA",X"65",X"55",X"55",X"55",X"55",X"77",X"7F",X"A9",X"99",X"55",X"55",X"55",X"D5",X"55",X"DF",
		X"AA",X"65",X"59",X"55",X"55",X"55",X"57",X"77",X"A9",X"95",X"55",X"55",X"55",X"55",X"D5",X"DF",
		X"A6",X"96",X"55",X"55",X"55",X"55",X"55",X"DF",X"AA",X"65",X"55",X"55",X"55",X"5D",X"57",X"7F",
		X"A5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"DA",X"55",X"55",X"55",X"55",X"57",X"7F",
		X"AA",X"DA",X"55",X"55",X"55",X"55",X"57",X"3F",X"AA",X"DA",X"AA",X"AA",X"AA",X"AA",X"AB",X"6A",
		X"11",X"04",X"45",X"11",X"04",X"00",X"00",X"00",X"40",X"40",X"40",X"10",X"40",X"41",X"01",X"01",
		X"15",X"14",X"11",X"04",X"04",X"10",X"10",X"44",X"45",X"50",X"55",X"44",X"41",X"00",X"44",X"11",
		X"55",X"45",X"05",X"15",X"10",X"44",X"11",X"05",X"14",X"55",X"55",X"44",X"15",X"55",X"55",X"54",
		X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"65",X"55",X"95",X"59",X"59",X"55",X"55",X"59",X"55",
		X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",
		X"75",X"59",X"59",X"65",X"65",X"55",X"56",X"55",X"59",X"99",X"55",X"55",X"55",X"95",X"65",X"55",
		X"75",X"57",X"55",X"DD",X"55",X"55",X"55",X"67",X"DF",X"75",X"ED",X"55",X"76",X"55",X"75",X"55",
		X"FD",X"DF",X"57",X"75",X"D5",X"75",X"D7",X"75",X"FF",X"FD",X"FF",X"FF",X"77",X"5F",X"F7",X"DF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"F5",X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"F7",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"7F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"5F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"FF",
		X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",X"7F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"DF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"DF",X"FF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",X"DF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"D7",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",X"F5",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F5",X"5A",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"75",X"55",X"9F",
		X"FF",X"FF",X"DF",X"FF",X"7F",X"F5",X"56",X"A7",X"FF",X"FF",X"DF",X"FF",X"FF",X"D5",X"FE",X"7B",
		X"FF",X"FD",X"DF",X"FF",X"FF",X"D7",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"D5",X"FE",X"EF",
		X"FD",X"FF",X"FF",X"F7",X"FF",X"D7",X"FB",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",X"5F",X"FF",X"FF",
		X"FF",X"FF",X"F7",X"DF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"F5",X"FF",X"FF",X"7F",X"FF",X"FF",
		X"FF",X"FF",X"DF",X"FF",X"D5",X"FF",X"FF",X"FF",X"FF",X"DF",X"FF",X"FF",X"F7",X"DF",X"DF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"F5",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"F7",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"5F",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"56",X"AA",X"AA",X"AA",X"51",X"55",X"55",X"55",X"56",X"AA",X"AA",X"AA",
		X"59",X"59",X"55",X"55",X"59",X"A9",X"A6",X"AA",X"54",X"55",X"59",X"55",X"56",X"9A",X"AA",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"6A",X"AA",X"AA",X"5D",X"57",X"55",X"55",X"55",X"99",X"A6",X"AA",
		X"55",X"D5",X"55",X"55",X"55",X"66",X"9A",X"6A",X"DD",X"55",X"55",X"59",X"55",X"95",X"6A",X"AA",
		X"75",X"55",X"55",X"55",X"55",X"55",X"9A",X"AA",X"55",X"DD",X"65",X"55",X"55",X"55",X"6A",X"6A",
		X"5D",X"55",X"55",X"55",X"55",X"56",X"5A",X"AA",X"77",X"5D",X"75",X"55",X"55",X"55",X"66",X"A6",
		X"DD",X"D5",X"55",X"55",X"55",X"55",X"56",X"AA",X"F7",X"57",X"55",X"55",X"55",X"55",X"56",X"AA",
		X"DD",X"D5",X"55",X"95",X"55",X"56",X"59",X"AA",X"FF",X"5D",X"75",X"55",X"55",X"55",X"96",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"A5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"AA",X"DA",X"AA",X"AA",X"AA",X"AA",X"AB",X"6A",
		X"AA",X"DA",X"AA",X"AA",X"AA",X"AA",X"AB",X"2A",X"AA",X"DA",X"AA",X"AA",X"AA",X"AA",X"AB",X"6A",
		X"00",X"D0",X"00",X"00",X"00",X"00",X"03",X"40",X"00",X"D1",X"40",X"00",X"00",X"00",X"03",X"44",
		X"00",X"D4",X"00",X"00",X"00",X"00",X"03",X"50",X"00",X"D0",X"00",X"00",X"00",X"01",X"03",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"7F",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"5F",X"7D",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"F7",X"FF",X"FF",X"FF",
		X"FF",X"FD",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"7F",X"FF",X"DF",X"FF",
		X"FD",X"DF",X"5F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FD",X"FF",X"DF",X"7D",X"FF",X"FF",X"F7",X"FF",X"D7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",
		X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"D6",X"AF",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"D6",X"AF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"D7",X"AF",X"FF",X"FF",X"FF",X"F7",X"FD",X"FF",X"D5",X"5F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"D5",X"FF",X"FF",X"FF",X"7F",X"F7",X"FD",X"DF",X"D5",X"FF",
		X"FF",X"FD",X"FF",X"5F",X"F7",X"FF",X"D7",X"FF",X"FF",X"F5",X"FF",X"DF",X"FF",X"FF",X"5F",X"FF",
		X"FF",X"DD",X"FD",X"7F",X"FF",X"FF",X"5F",X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",X"F5",X"FF",X"FF",
		X"FF",X"FF",X"F5",X"FF",X"7F",X"FD",X"7F",X"FF",X"FF",X"FF",X"FF",X"57",X"FF",X"F5",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"F7",X"FD",X"57",X"FF",X"FF",X"FF",X"FF",X"FF",X"F5",X"DD",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"DF",X"FF",X"FF",X"FF",X"DD",X"FF",
		X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EA",X"FF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"6A",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"5D",X"FF",X"FF",X"77",X"FF",X"FF",X"FD",X"DF",X"77",
		X"FF",X"FF",X"FD",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",X"FF",X"FD",X"F7",X"FD",X"F7",X"77",X"7F",
		X"FF",X"FF",X"FF",X"F7",X"7F",X"F7",X"F5",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"DF",X"DF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"5F",X"FF",X"FD",X"FF",X"F7",X"FF",X"FF",X"F5",X"D7",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DA",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DA",X"BF",
		X"FF",X"7F",X"FF",X"FF",X"FF",X"7F",X"DA",X"BF",X"FD",X"7F",X"FF",X"F7",X"FF",X"FF",X"D5",X"7F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"57",X"7F",X"FF",X"DF",X"FF",X"DF",X"FF",X"7D",X"7D",X"FF",
		X"FF",X"FD",X"FF",X"FF",X"FF",X"FD",X"F7",X"FF",X"FF",X"FD",X"7F",X"7F",X"FD",X"FF",X"DF",X"FF",
		X"FF",X"FF",X"7D",X"7F",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"FD",X"5F",X"D7",X"D7",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"D7",X"55",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"D7",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"65",X"55",X"55",X"55",X"55",X"59",X"AA",X"AA",X"95",X"55",X"59",X"95",X"55",X"56",X"9A",
		X"A9",X"A5",X"55",X"55",X"55",X"55",X"59",X"AA",X"AA",X"99",X"55",X"55",X"95",X"55",X"56",X"6A",
		X"AA",X"55",X"55",X"59",X"65",X"55",X"59",X"AA",X"AA",X"99",X"55",X"55",X"55",X"55",X"56",X"9A",
		X"AA",X"A5",X"55",X"55",X"95",X"55",X"59",X"AA",X"AA",X"69",X"55",X"55",X"55",X"55",X"66",X"6A",
		X"AA",X"A6",X"55",X"55",X"95",X"55",X"59",X"AA",X"AA",X"A9",X"95",X"59",X"55",X"55",X"56",X"AA",
		X"AA",X"66",X"56",X"55",X"95",X"55",X"55",X"AA",X"AA",X"A9",X"55",X"65",X"55",X"55",X"55",X"6A",
		X"AA",X"A5",X"56",X"56",X"65",X"55",X"55",X"AA",X"AA",X"99",X"55",X"55",X"55",X"55",X"66",X"AA",
		X"AA",X"A9",X"55",X"55",X"95",X"55",X"99",X"AA",X"AA",X"A6",X"55",X"55",X"55",X"55",X"66",X"AA",
		X"AA",X"A9",X"55",X"59",X"55",X"55",X"5A",X"6A",X"AA",X"A6",X"55",X"55",X"55",X"55",X"56",X"AA",
		X"AA",X"A9",X"95",X"55",X"55",X"55",X"59",X"AA",X"AA",X"AA",X"65",X"56",X"55",X"55",X"56",X"AA",
		X"AA",X"A9",X"95",X"55",X"55",X"55",X"5A",X"9A",X"AA",X"AA",X"69",X"55",X"55",X"55",X"66",X"AA",
		X"AA",X"AA",X"95",X"55",X"55",X"59",X"9A",X"AA",X"AA",X"A9",X"A5",X"55",X"95",X"5A",X"69",X"AA",
		X"AA",X"AA",X"99",X"95",X"55",X"A6",X"AA",X"AA",X"AA",X"AA",X"A5",X"65",X"56",X"6A",X"9A",X"AA",
		X"AA",X"9A",X"A9",X"95",X"59",X"AA",X"AA",X"AA",X"AA",X"AA",X"9A",X"65",X"56",X"66",X"AA",X"AA",
		X"AA",X"AA",X"A9",X"99",X"59",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"6A",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"6A",X"A6",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"88",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"A5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"AA",X"DA",X"AA",X"AA",X"AA",X"AA",X"AB",X"6A",
		X"AA",X"DA",X"AA",X"AA",X"AA",X"AA",X"AB",X"2A",X"AA",X"DA",X"AA",X"AA",X"AA",X"AA",X"AB",X"6A",
		X"A0",X"D0",X"00",X"00",X"00",X"00",X"03",X"40",X"A0",X"D1",X"40",X"00",X"00",X"00",X"03",X"44",
		X"80",X"D4",X"00",X"00",X"00",X"00",X"03",X"50",X"80",X"D0",X"00",X"00",X"00",X"01",X"03",X"40",
		X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A8",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"AB",X"00",X"10",X"00",X"04",X"00",X"00",X"00",
		X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"10",X"00",X"01",X"00",X"00",X"00",X"00",
		X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A8",X"00",X"10",X"00",X"00",X"00",X"00",X"00",
		X"A0",X"00",X"00",X"00",X"00",X"40",X"01",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A0",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F6",X"AA",X"AA",X"00",X"00",X"00",X"00",X"40",X"B6",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"FA",X"AA",X"A6",X"10",X"00",X"00",X"00",X"00",X"EA",X"AA",X"AA",
		X"00",X"00",X"00",X"40",X"03",X"EA",X"AA",X"AA",X"00",X"00",X"00",X"00",X"03",X"6A",X"AA",X"AA",
		X"00",X"04",X"00",X"00",X"4D",X"6A",X"AA",X"AA",X"00",X"00",X"00",X"00",X"0E",X"6A",X"AA",X"AA",
		X"01",X"00",X"00",X"40",X"0B",X"5A",X"AA",X"AA",X"00",X"00",X"00",X"00",X"02",X"D6",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"D6",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"B6",X"AA",X"AA",
		X"03",X"00",X"00",X"00",X"70",X"26",X"AA",X"AA",X"07",X"00",X"00",X"01",X"70",X"36",X"AA",X"AA",
		X"07",X"00",X"00",X"14",X"70",X"BA",X"6A",X"AA",X"07",X"00",X"00",X"00",X"70",X"AA",X"AA",X"AA",
		X"A7",X"AA",X"AA",X"AA",X"7A",X"AA",X"AA",X"AA",X"A7",X"AA",X"AA",X"AA",X"7A",X"AA",X"AA",X"AA",
		X"A7",X"AA",X"AA",X"AA",X"7A",X"AA",X"AA",X"AA",X"BF",X"FF",X"FF",X"FF",X"FF",X"EA",X"AA",X"AA",
		X"BF",X"FF",X"FF",X"FF",X"FF",X"EA",X"AA",X"A6",X"95",X"55",X"55",X"55",X"55",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"9A",X"A6",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"A9",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"A6",X"AA",X"AA",X"AA",X"9A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"A9",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"1A",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"1A",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"1A",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"2A",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"01",X"6A",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"5A",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"1A",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"1A",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"2A",X"AA",X"6A",X"00",X"00",X"00",X"00",X"00",X"6A",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"5A",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"16",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"06",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"0A",X"AA",X"A6",
		X"00",X"00",X"00",X"00",X"00",X"2A",X"AA",X"A6",X"00",X"00",X"00",X"00",X"00",X"6A",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"6A",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"5A",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"1A",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"1A",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"2A",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"6A",X"A6",X"AA",
		X"00",X"00",X"00",X"00",X"01",X"6A",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"6A",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"6A",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"16",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"06",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"06",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"06",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"06",X"AA",X"AA");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
