library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity burnin_rubber_sound_prog is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of burnin_rubber_sound_prog is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"78",X"D8",X"A2",X"FF",X"9A",X"A2",X"72",X"A9",X"00",X"95",X"00",X"CA",X"D0",X"FB",X"20",X"1D",
		X"F0",X"AD",X"00",X"A0",X"A9",X"FF",X"8D",X"00",X"C0",X"58",X"4C",X"1A",X"F0",X"A2",X"0F",X"8E",
		X"00",X"40",X"8E",X"00",X"80",X"BD",X"50",X"F0",X"8D",X"00",X"20",X"8D",X"00",X"60",X"CA",X"10",
		X"EE",X"60",X"A2",X"0A",X"8E",X"00",X"40",X"BD",X"50",X"F0",X"8D",X"00",X"20",X"CA",X"10",X"F4",
		X"60",X"A2",X"0A",X"8E",X"00",X"80",X"BD",X"50",X"F0",X"8D",X"00",X"60",X"CA",X"10",X"F4",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"48",X"8A",X"48",X"98",X"48",X"AD",X"00",X"A0",X"30",X"37",X"A5",X"51",X"C9",X"01",X"F0",X"13",
		X"C9",X"05",X"F0",X"0F",X"AD",X"00",X"A0",X"85",X"51",X"85",X"6D",X"C9",X"14",X"90",X"0A",X"A9",
		X"00",X"85",X"51",X"68",X"A8",X"68",X"AA",X"68",X"40",X"A2",X"FF",X"9A",X"20",X"32",X"F0",X"A5",
		X"51",X"58",X"0A",X"AA",X"BD",X"2A",X"F1",X"85",X"4D",X"BD",X"2B",X"F1",X"85",X"4E",X"6C",X"4D",
		X"00",X"29",X"07",X"85",X"4A",X"A9",X"00",X"85",X"4C",X"A5",X"4A",X"48",X"20",X"FA",X"F0",X"AA",
		X"BD",X"06",X"F1",X"85",X"44",X"85",X"45",X"BD",X"09",X"F1",X"85",X"46",X"85",X"47",X"BD",X"0C",
		X"F1",X"85",X"48",X"85",X"49",X"BD",X"0F",X"F1",X"85",X"32",X"BD",X"12",X"F1",X"85",X"34",X"BD",
		X"15",X"F1",X"85",X"36",X"68",X"0A",X"AA",X"BD",X"18",X"F1",X"85",X"14",X"BD",X"19",X"F1",X"85",
		X"15",X"BD",X"1E",X"F1",X"85",X"16",X"BD",X"1F",X"F1",X"85",X"17",X"BD",X"24",X"F1",X"85",X"18",
		X"BD",X"25",X"F1",X"85",X"19",X"85",X"10",X"4C",X"83",X"F0",X"48",X"A2",X"49",X"A9",X"00",X"95",
		X"00",X"CA",X"D0",X"FB",X"68",X"60",X"0F",X"0A",X"0F",X"0F",X"0A",X"0F",X"0C",X"08",X"0C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"8B",X"F7",X"DA",X"F7",X"37",X"FC",X"A6",X"F7",
		X"65",X"F9",X"50",X"FC",X"C0",X"F7",X"EF",X"FA",X"68",X"FC",X"00",X"F0",X"52",X"F1",X"83",X"F1",
		X"83",X"F1",X"83",X"F1",X"52",X"F1",X"52",X"F1",X"52",X"F1",X"A4",X"F1",X"A4",X"F1",X"A4",X"F1",
		X"0F",X"F2",X"0F",X"F2",X"0F",X"F2",X"0F",X"F2",X"0F",X"F2",X"0F",X"F2",X"0F",X"F2",X"0F",X"F2",
		X"0F",X"F2",X"A5",X"6A",X"D0",X"27",X"A5",X"51",X"C9",X"01",X"D0",X"03",X"4C",X"63",X"F1",X"C9",
		X"05",X"D0",X"02",X"85",X"6A",X"0A",X"AA",X"BD",X"30",X"F2",X"85",X"53",X"85",X"5C",X"BD",X"31",
		X"F2",X"85",X"54",X"A9",X"00",X"85",X"59",X"85",X"5F",X"A9",X"08",X"85",X"62",X"4C",X"19",X"F0",
		X"4C",X"D2",X"F1",X"A5",X"10",X"F0",X"F9",X"A5",X"51",X"0A",X"AA",X"BD",X"30",X"F2",X"85",X"55",
		X"85",X"5D",X"BD",X"31",X"F2",X"85",X"56",X"A9",X"00",X"85",X"5A",X"85",X"60",X"A9",X"02",X"85",
		X"63",X"4C",X"19",X"F0",X"A5",X"6F",X"D0",X"20",X"A5",X"51",X"0A",X"AA",X"BD",X"30",X"F2",X"85",
		X"57",X"85",X"5E",X"BD",X"31",X"F2",X"85",X"58",X"A9",X"00",X"85",X"5B",X"85",X"61",X"A9",X"04",
		X"85",X"64",X"A5",X"51",X"C9",X"08",X"F0",X"03",X"4C",X"19",X"F0",X"A9",X"FF",X"85",X"6F",X"4C",
		X"19",X"F0",X"A9",X"00",X"85",X"6A",X"A2",X"04",X"BD",X"30",X"F2",X"85",X"65",X"BD",X"31",X"F2",
		X"85",X"66",X"A0",X"00",X"B1",X"65",X"C9",X"80",X"F0",X"15",X"8D",X"00",X"80",X"C8",X"B1",X"65",
		X"8D",X"00",X"60",X"C8",X"B1",X"65",X"85",X"67",X"20",X"02",X"F2",X"C8",X"4C",X"E4",X"F1",X"4C",
		X"19",X"F0",X"A9",X"F0",X"85",X"68",X"C6",X"68",X"D0",X"FC",X"C6",X"67",X"D0",X"F8",X"60",X"A5",
		X"6D",X"85",X"6E",X"0A",X"AA",X"BD",X"30",X"F2",X"85",X"53",X"85",X"5C",X"85",X"69",X"BD",X"31",
		X"F2",X"85",X"54",X"A9",X"00",X"85",X"59",X"85",X"5F",X"A9",X"01",X"85",X"62",X"4C",X"19",X"F0",
		X"83",X"F0",X"58",X"F2",X"89",X"F2",X"ED",X"F2",X"87",X"F3",X"B5",X"F3",X"E6",X"F3",X"17",X"F4",
		X"30",X"F4",X"61",X"F4",X"71",X"F4",X"96",X"F4",X"AF",X"F4",X"C8",X"F4",X"E1",X"F4",X"FA",X"F4",
		X"13",X"F5",X"23",X"F5",X"33",X"F5",X"43",X"F5",X"00",X"00",X"01",X"01",X"00",X"01",X"07",X"F7",
		X"01",X"08",X"0C",X"01",X"06",X"1F",X"20",X"08",X"0B",X"01",X"06",X"1C",X"10",X"08",X"0C",X"01",
		X"06",X"1F",X"20",X"08",X"0B",X"01",X"06",X"1C",X"20",X"08",X"09",X"01",X"06",X"16",X"30",X"06",
		X"1A",X"10",X"06",X"00",X"01",X"08",X"00",X"01",X"80",X"07",X"F0",X"01",X"03",X"00",X"01",X"02",
		X"B3",X"08",X"09",X"0F",X"08",X"02",X"59",X"08",X"09",X"0E",X"08",X"02",X"B3",X"08",X"09",X"0D",
		X"08",X"02",X"59",X"08",X"09",X"0C",X"08",X"02",X"B3",X"08",X"09",X"0B",X"08",X"02",X"59",X"08",
		X"09",X"0A",X"08",X"02",X"B3",X"08",X"09",X"09",X"08",X"02",X"59",X"08",X"09",X"08",X"08",X"02",
		X"B3",X"08",X"09",X"07",X"08",X"02",X"59",X"08",X"09",X"06",X"08",X"02",X"B3",X"08",X"09",X"05",
		X"08",X"02",X"59",X"08",X"09",X"04",X"08",X"02",X"B3",X"08",X"09",X"03",X"08",X"02",X"59",X"08",
		X"09",X"02",X"08",X"02",X"B3",X"08",X"09",X"00",X"01",X"02",X"00",X"01",X"80",X"09",X"0B",X"01",
		X"03",X"00",X"01",X"02",X"5F",X"04",X"02",X"3C",X"04",X"02",X"5C",X"04",X"02",X"3A",X"04",X"02",
		X"5A",X"04",X"02",X"39",X"04",X"02",X"58",X"04",X"02",X"37",X"04",X"02",X"57",X"04",X"02",X"35",
		X"04",X"02",X"54",X"04",X"02",X"33",X"04",X"02",X"53",X"04",X"02",X"31",X"04",X"02",X"51",X"04",
		X"02",X"2E",X"04",X"02",X"4F",X"04",X"02",X"2D",X"04",X"02",X"4D",X"04",X"02",X"2B",X"04",X"02",
		X"4B",X"04",X"02",X"29",X"04",X"02",X"49",X"04",X"02",X"27",X"04",X"02",X"47",X"04",X"02",X"26",
		X"04",X"02",X"45",X"04",X"02",X"24",X"04",X"02",X"44",X"04",X"02",X"22",X"04",X"02",X"42",X"04",
		X"02",X"20",X"04",X"02",X"40",X"04",X"02",X"2E",X"04",X"02",X"3E",X"04",X"02",X"28",X"04",X"02",
		X"3C",X"04",X"02",X"1A",X"04",X"02",X"3A",X"04",X"02",X"18",X"04",X"02",X"38",X"04",X"02",X"16",
		X"04",X"02",X"36",X"04",X"02",X"14",X"04",X"02",X"34",X"04",X"02",X"12",X"04",X"02",X"30",X"04",
		X"02",X"0E",X"04",X"02",X"00",X"01",X"80",X"09",X"0B",X"01",X"02",X"00",X"01",X"02",X"2A",X"05",
		X"02",X"8E",X"05",X"02",X"25",X"05",X"02",X"7E",X"05",X"02",X"21",X"05",X"02",X"20",X"05",X"02",
		X"1D",X"05",X"02",X"64",X"05",X"02",X"1C",X"05",X"02",X"5E",X"05",X"02",X"1F",X"05",X"02",X"6A",
		X"05",X"02",X"00",X"06",X"80",X"07",X"F7",X"01",X"08",X"0A",X"01",X"06",X"10",X"20",X"08",X"0C",
		X"01",X"06",X"1F",X"20",X"08",X"0B",X"01",X"06",X"1C",X"10",X"08",X"0C",X"01",X"06",X"1F",X"20",
		X"08",X"0B",X"01",X"06",X"1C",X"20",X"08",X"09",X"01",X"06",X"16",X"30",X"06",X"1A",X"10",X"06",
		X"00",X"01",X"08",X"00",X"01",X"80",X"00",X"00",X"01",X"01",X"00",X"01",X"06",X"1F",X"01",X"08",
		X"0A",X"05",X"06",X"14",X"01",X"08",X"0C",X"05",X"06",X"18",X"01",X"08",X"0D",X"05",X"06",X"10",
		X"01",X"08",X"0C",X"10",X"08",X"0A",X"05",X"08",X"08",X"05",X"08",X"06",X"05",X"08",X"04",X"05",
		X"08",X"02",X"05",X"06",X"00",X"01",X"80",X"08",X"0B",X"01",X"06",X"1F",X"0A",X"08",X"0A",X"02",
		X"06",X"1C",X"02",X"08",X"0B",X"02",X"06",X"18",X"02",X"08",X"07",X"02",X"08",X"00",X"01",X"80",
		X"0A",X"0D",X"01",X"05",X"00",X"01",X"04",X"77",X"0A",X"04",X"3B",X"0A",X"04",X"77",X"0A",X"04",
		X"3B",X"0A",X"04",X"77",X"0A",X"04",X"3B",X"0A",X"04",X"77",X"0A",X"04",X"3B",X"0A",X"04",X"77",
		X"0A",X"04",X"3B",X"0A",X"04",X"77",X"0A",X"04",X"3B",X"0A",X"0A",X"00",X"01",X"04",X"00",X"01",
		X"80",X"05",X"00",X"01",X"04",X"2F",X"01",X"0A",X"0F",X"0F",X"0A",X"00",X"01",X"04",X"00",X"01",
		X"80",X"05",X"00",X"01",X"0A",X"0D",X"01",X"04",X"7F",X"04",X"04",X"5F",X"04",X"04",X"78",X"04",
		X"04",X"58",X"04",X"04",X"70",X"04",X"04",X"50",X"04",X"04",X"68",X"04",X"04",X"48",X"04",X"0A",
		X"00",X"01",X"04",X"00",X"01",X"80",X"00",X"FF",X"01",X"01",X"08",X"01",X"08",X"0A",X"02",X"00",
		X"FF",X"01",X"01",X"07",X"01",X"08",X"09",X"02",X"00",X"BF",X"01",X"01",X"07",X"01",X"81",X"00",
		X"6F",X"01",X"01",X"08",X"01",X"08",X"0A",X"02",X"00",X"6F",X"01",X"01",X"07",X"01",X"08",X"09",
		X"02",X"00",X"2F",X"01",X"01",X"07",X"01",X"81",X"00",X"BF",X"01",X"01",X"07",X"01",X"08",X"0A",
		X"02",X"00",X"BF",X"01",X"01",X"06",X"01",X"08",X"09",X"02",X"00",X"7F",X"01",X"01",X"06",X"01",
		X"81",X"00",X"1F",X"01",X"01",X"07",X"01",X"08",X"0A",X"01",X"00",X"1F",X"01",X"01",X"06",X"01",
		X"08",X"0A",X"01",X"00",X"CF",X"01",X"01",X"05",X"01",X"81",X"00",X"6F",X"01",X"01",X"06",X"01",
		X"08",X"0A",X"01",X"00",X"6F",X"01",X"01",X"05",X"01",X"08",X"0A",X"01",X"00",X"2F",X"01",X"01",
		X"05",X"01",X"81",X"00",X"BF",X"01",X"01",X"05",X"01",X"08",X"0A",X"01",X"00",X"BF",X"01",X"01",
		X"04",X"01",X"81",X"00",X"2F",X"01",X"01",X"05",X"01",X"08",X"0A",X"01",X"00",X"2F",X"01",X"01",
		X"04",X"01",X"81",X"00",X"1F",X"01",X"01",X"05",X"01",X"08",X"0A",X"01",X"00",X"1F",X"01",X"01",
		X"04",X"01",X"81",X"00",X"00",X"01",X"01",X"00",X"01",X"08",X"00",X"01",X"81",X"4C",X"83",X"F0",
		X"48",X"8A",X"48",X"98",X"48",X"A5",X"10",X"F0",X"F4",X"A5",X"11",X"29",X"07",X"E6",X"11",X"0A",
		X"AA",X"BD",X"7E",X"F5",X"85",X"12",X"BD",X"7F",X"F5",X"85",X"13",X"A9",X"07",X"8D",X"00",X"80",
		X"A5",X"62",X"05",X"63",X"05",X"64",X"49",X"FF",X"8D",X"00",X"60",X"6C",X"12",X"00",X"67",X"F6",
		X"67",X"F6",X"67",X"F6",X"10",X"F7",X"8E",X"F5",X"E9",X"F5",X"20",X"F6",X"83",X"F0",X"A5",X"5C",
		X"F0",X"23",X"A5",X"59",X"D0",X"1D",X"A4",X"5F",X"B1",X"53",X"C9",X"80",X"F0",X"21",X"C9",X"81",
		X"F0",X"16",X"8D",X"00",X"80",X"C8",X"B1",X"53",X"8D",X"00",X"60",X"C8",X"B1",X"53",X"85",X"59",
		X"C8",X"84",X"5F",X"C6",X"59",X"4C",X"83",X"F0",X"A9",X"00",X"85",X"5F",X"4C",X"83",X"F0",X"A5",
		X"51",X"C9",X"01",X"F0",X"0F",X"C9",X"05",X"F0",X"0B",X"A9",X"00",X"85",X"6A",X"A5",X"6E",X"85",
		X"6D",X"4C",X"0F",X"F2",X"A9",X"08",X"8D",X"00",X"80",X"A9",X"00",X"8D",X"00",X"60",X"85",X"5C",
		X"85",X"6A",X"85",X"51",X"85",X"62",X"4C",X"83",X"F0",X"A5",X"5D",X"F0",X"1F",X"A5",X"5A",X"D0",
		X"19",X"A4",X"60",X"B1",X"55",X"C9",X"80",X"F0",X"16",X"8D",X"00",X"80",X"C8",X"B1",X"55",X"8D",
		X"00",X"60",X"C8",X"B1",X"55",X"85",X"5A",X"C8",X"84",X"60",X"C6",X"5A",X"4C",X"83",X"F0",X"A9",
		X"09",X"8D",X"00",X"80",X"A9",X"00",X"8D",X"00",X"60",X"85",X"5D",X"85",X"63",X"4C",X"83",X"F0",
		X"A5",X"5E",X"F0",X"1F",X"A5",X"5B",X"D0",X"19",X"A4",X"61",X"B1",X"57",X"C9",X"80",X"F0",X"16",
		X"8D",X"00",X"80",X"C8",X"B1",X"57",X"8D",X"00",X"60",X"C8",X"B1",X"57",X"85",X"5B",X"C8",X"84",
		X"61",X"C6",X"5B",X"4C",X"83",X"F0",X"A9",X"00",X"85",X"6F",X"85",X"5E",X"85",X"64",X"4C",X"83",
		X"F0",X"20",X"FA",X"F0",X"20",X"32",X"F0",X"E6",X"4C",X"4C",X"A9",X"F0",X"20",X"FA",X"F0",X"20",
		X"32",X"F0",X"A9",X"01",X"4C",X"A1",X"F0",X"B5",X"1A",X"D0",X"75",X"A1",X"14",X"C9",X"FE",X"F0",
		X"E0",X"C9",X"FF",X"F0",X"E7",X"20",X"64",X"F7",X"48",X"29",X"0F",X"A8",X"B9",X"6B",X"F7",X"95",
		X"26",X"B9",X"7B",X"F7",X"95",X"27",X"68",X"85",X"4B",X"4A",X"4A",X"4A",X"4A",X"A8",X"D0",X"0A",
		X"95",X"26",X"95",X"27",X"95",X"2C",X"95",X"2D",X"F0",X"29",X"56",X"27",X"76",X"26",X"88",X"D0",
		X"F9",X"18",X"A5",X"4B",X"75",X"32",X"48",X"29",X"0F",X"A8",X"B9",X"6B",X"F7",X"95",X"2C",X"B9",
		X"7B",X"F7",X"95",X"2D",X"68",X"4A",X"4A",X"4A",X"4A",X"A8",X"56",X"2D",X"76",X"2C",X"88",X"D0",
		X"F9",X"B5",X"44",X"95",X"45",X"A1",X"14",X"20",X"64",X"F7",X"95",X"1A",X"95",X"20",X"A0",X"02",
		X"56",X"20",X"88",X"D0",X"FB",X"B5",X"20",X"95",X"21",X"D6",X"1A",X"D6",X"21",X"4C",X"83",X"F0",
		X"D6",X"1A",X"D6",X"21",X"D0",X"0A",X"B5",X"20",X"95",X"21",X"B5",X"45",X"F0",X"02",X"D6",X"45",
		X"B5",X"3E",X"29",X"01",X"D0",X"0D",X"F6",X"3E",X"B5",X"26",X"95",X"38",X"B5",X"27",X"95",X"39",
		X"4C",X"83",X"F0",X"F6",X"3E",X"B5",X"2C",X"95",X"38",X"B5",X"2D",X"95",X"39",X"4C",X"83",X"F0",
		X"A2",X"05",X"8E",X"00",X"40",X"B5",X"38",X"8D",X"00",X"20",X"CA",X"10",X"F5",X"A5",X"4C",X"29",
		X"01",X"D0",X"0C",X"A9",X"07",X"8D",X"00",X"40",X"A9",X"F8",X"8D",X"00",X"20",X"D0",X"0A",X"A9",
		X"07",X"8D",X"00",X"40",X"A9",X"DC",X"8D",X"00",X"20",X"A9",X"08",X"8D",X"00",X"40",X"A5",X"45",
		X"8D",X"00",X"20",X"A9",X"09",X"8D",X"00",X"40",X"A5",X"47",X"8D",X"00",X"20",X"A9",X"0A",X"8D",
		X"00",X"40",X"A5",X"49",X"8D",X"00",X"20",X"A9",X"06",X"8D",X"00",X"40",X"A9",X"02",X"8D",X"00",
		X"20",X"4C",X"83",X"F0",X"F6",X"14",X"D0",X"02",X"F6",X"15",X"60",X"65",X"23",X"F3",X"D5",X"C6",
		X"C7",X"D6",X"F2",X"1B",X"51",X"91",X"DD",X"32",X"91",X"F9",X"6A",X"16",X"15",X"13",X"12",X"11",
		X"10",X"0F",X"0E",X"0E",X"0D",X"0C",X"0B",X"0B",X"0A",X"09",X"09",X"47",X"20",X"47",X"10",X"47",
		X"10",X"47",X"60",X"49",X"20",X"47",X"20",X"49",X"20",X"47",X"20",X"47",X"10",X"47",X"10",X"47",
		X"40",X"47",X"40",X"00",X"40",X"FF",X"44",X"20",X"44",X"10",X"44",X"10",X"44",X"60",X"45",X"20",
		X"44",X"20",X"45",X"20",X"44",X"20",X"44",X"10",X"44",X"10",X"44",X"40",X"44",X"40",X"00",X"40",
		X"40",X"20",X"40",X"10",X"40",X"10",X"40",X"60",X"40",X"20",X"40",X"20",X"40",X"20",X"40",X"20",
		X"40",X"10",X"40",X"10",X"40",X"40",X"40",X"40",X"00",X"40",X"44",X"18",X"44",X"18",X"40",X"18",
		X"40",X"18",X"42",X"18",X"42",X"18",X"45",X"30",X"44",X"18",X"44",X"18",X"40",X"18",X"40",X"18",
		X"42",X"18",X"42",X"18",X"37",X"30",X"44",X"18",X"44",X"18",X"40",X"18",X"40",X"18",X"42",X"18",
		X"42",X"18",X"44",X"18",X"45",X"18",X"47",X"18",X"47",X"18",X"50",X"18",X"47",X"18",X"44",X"18",
		X"47",X"18",X"50",X"30",X"50",X"18",X"49",X"30",X"45",X"18",X"4B",X"18",X"47",X"30",X"44",X"18",
		X"49",X"18",X"45",X"30",X"42",X"18",X"47",X"18",X"44",X"30",X"40",X"18",X"40",X"18",X"44",X"18",
		X"47",X"18",X"47",X"18",X"42",X"18",X"45",X"18",X"49",X"18",X"49",X"18",X"47",X"18",X"4B",X"18",
		X"52",X"18",X"54",X"18",X"50",X"30",X"00",X"30",X"50",X"24",X"4B",X"0C",X"45",X"30",X"4B",X"24",
		X"49",X"0C",X"44",X"30",X"44",X"24",X"45",X"0C",X"47",X"30",X"30",X"0C",X"32",X"0C",X"34",X"0C",
		X"35",X"0C",X"37",X"0C",X"39",X"0C",X"3B",X"0C",X"40",X"0C",X"45",X"24",X"47",X"0C",X"49",X"30",
		X"32",X"0C",X"34",X"0C",X"35",X"0C",X"37",X"0C",X"39",X"0C",X"3B",X"0C",X"30",X"0C",X"32",X"0C",
		X"44",X"18",X"44",X"18",X"45",X"18",X"45",X"18",X"47",X"18",X"47",X"18",X"40",X"30",X"44",X"18",
		X"40",X"18",X"42",X"18",X"45",X"18",X"44",X"18",X"42",X"18",X"40",X"30",X"44",X"18",X"44",X"0C",
		X"44",X"0C",X"40",X"18",X"40",X"0C",X"40",X"0C",X"45",X"18",X"44",X"18",X"42",X"30",X"44",X"18",
		X"44",X"0C",X"44",X"0C",X"40",X"18",X"40",X"0C",X"40",X"0C",X"44",X"18",X"42",X"18",X"40",X"30",
		X"44",X"18",X"44",X"0C",X"44",X"0C",X"40",X"18",X"40",X"0C",X"40",X"0C",X"42",X"0C",X"44",X"0C",
		X"45",X"0C",X"47",X"0C",X"4B",X"30",X"44",X"18",X"44",X"0C",X"44",X"0C",X"40",X"18",X"40",X"0C",
		X"40",X"0C",X"45",X"18",X"44",X"18",X"42",X"30",X"44",X"18",X"44",X"0C",X"44",X"0C",X"40",X"18",
		X"40",X"0C",X"40",X"0C",X"3B",X"0C",X"39",X"0C",X"3B",X"0C",X"40",X"0C",X"42",X"30",X"44",X"18",
		X"44",X"0C",X"44",X"0C",X"40",X"18",X"40",X"0C",X"40",X"0C",X"42",X"0C",X"44",X"0C",X"45",X"0C",
		X"47",X"0C",X"49",X"30",X"4B",X"18",X"4B",X"0C",X"4B",X"0C",X"47",X"18",X"47",X"0C",X"47",X"0C",
		X"50",X"0C",X"4B",X"0C",X"49",X"0C",X"4B",X"0C",X"50",X"30",X"50",X"18",X"49",X"18",X"45",X"18",
		X"47",X"18",X"4B",X"18",X"47",X"18",X"44",X"18",X"45",X"18",X"49",X"18",X"45",X"18",X"42",X"18",
		X"44",X"18",X"47",X"18",X"44",X"18",X"40",X"30",X"50",X"30",X"49",X"18",X"45",X"18",X"4B",X"18",
		X"4B",X"18",X"47",X"18",X"44",X"18",X"49",X"30",X"45",X"18",X"42",X"18",X"47",X"18",X"47",X"18",
		X"44",X"18",X"40",X"18",X"FE",X"40",X"18",X"40",X"18",X"39",X"18",X"39",X"18",X"3B",X"18",X"3B",
		X"18",X"42",X"30",X"40",X"18",X"40",X"18",X"39",X"18",X"39",X"18",X"3B",X"18",X"3B",X"18",X"34",
		X"30",X"40",X"18",X"40",X"18",X"39",X"18",X"39",X"18",X"3B",X"18",X"3B",X"18",X"40",X"18",X"42",
		X"18",X"44",X"18",X"44",X"18",X"49",X"18",X"44",X"18",X"40",X"18",X"44",X"18",X"49",X"30",X"49",
		X"18",X"45",X"30",X"42",X"18",X"47",X"18",X"44",X"30",X"40",X"18",X"45",X"18",X"42",X"30",X"3B",
		X"18",X"44",X"18",X"40",X"30",X"39",X"18",X"39",X"18",X"40",X"18",X"44",X"18",X"44",X"18",X"3B",
		X"18",X"42",X"18",X"45",X"18",X"45",X"18",X"44",X"18",X"47",X"18",X"4B",X"18",X"50",X"18",X"49",
		X"30",X"00",X"30",X"49",X"24",X"47",X"0C",X"42",X"30",X"47",X"24",X"45",X"0C",X"40",X"30",X"40",
		X"24",X"42",X"0C",X"44",X"30",X"29",X"0C",X"2B",X"0C",X"30",X"0C",X"32",X"0C",X"34",X"0C",X"35",
		X"0C",X"37",X"0C",X"39",X"0C",X"42",X"24",X"44",X"0C",X"45",X"30",X"2B",X"0C",X"30",X"0C",X"32",
		X"0C",X"34",X"0C",X"35",X"0C",X"37",X"0C",X"39",X"0C",X"3B",X"0C",X"40",X"18",X"40",X"18",X"42",
		X"18",X"42",X"18",X"44",X"18",X"44",X"18",X"39",X"30",X"40",X"18",X"39",X"18",X"3B",X"18",X"42",
		X"18",X"40",X"18",X"3B",X"18",X"39",X"30",X"40",X"18",X"40",X"0C",X"40",X"0C",X"39",X"18",X"39",
		X"0C",X"39",X"0C",X"42",X"18",X"40",X"18",X"3B",X"30",X"3B",X"18",X"3B",X"0C",X"3B",X"0C",X"39",
		X"18",X"39",X"0C",X"39",X"0C",X"40",X"18",X"3B",X"18",X"39",X"30",X"40",X"18",X"40",X"0C",X"40",
		X"0C",X"39",X"18",X"39",X"0C",X"39",X"0C",X"3B",X"0C",X"40",X"0C",X"42",X"0C",X"44",X"0C",X"47",
		X"30",X"40",X"18",X"40",X"0C",X"40",X"0C",X"39",X"18",X"39",X"0C",X"39",X"0C",X"42",X"18",X"40",
		X"18",X"3B",X"30",X"40",X"18",X"40",X"0C",X"40",X"0C",X"39",X"18",X"39",X"0C",X"39",X"0C",X"37",
		X"0C",X"35",X"0C",X"37",X"0C",X"39",X"0C",X"3B",X"30",X"40",X"18",X"40",X"0C",X"40",X"0C",X"39",
		X"18",X"39",X"0C",X"39",X"0C",X"3B",X"0C",X"40",X"0C",X"42",X"0C",X"44",X"0C",X"45",X"30",X"47",
		X"18",X"47",X"0C",X"47",X"0C",X"44",X"18",X"44",X"0C",X"44",X"0C",X"49",X"0C",X"47",X"0C",X"45",
		X"0C",X"47",X"0C",X"49",X"30",X"49",X"18",X"45",X"18",X"42",X"18",X"44",X"18",X"47",X"18",X"44",
		X"18",X"40",X"18",X"42",X"18",X"45",X"18",X"42",X"18",X"3B",X"18",X"40",X"18",X"44",X"18",X"40",
		X"18",X"39",X"30",X"49",X"30",X"45",X"18",X"42",X"18",X"47",X"18",X"47",X"18",X"44",X"18",X"40",
		X"18",X"45",X"30",X"42",X"18",X"3B",X"18",X"44",X"18",X"44",X"18",X"40",X"18",X"39",X"18",X"34",
		X"24",X"34",X"0C",X"30",X"30",X"32",X"24",X"32",X"0C",X"35",X"30",X"34",X"24",X"34",X"0C",X"30",
		X"30",X"32",X"24",X"32",X"0C",X"27",X"30",X"34",X"24",X"34",X"0C",X"30",X"30",X"32",X"24",X"32",
		X"0C",X"35",X"30",X"30",X"18",X"34",X"18",X"32",X"18",X"35",X"18",X"34",X"24",X"30",X"0C",X"34",
		X"30",X"40",X"24",X"39",X"0C",X"39",X"30",X"3B",X"24",X"37",X"0C",X"37",X"30",X"39",X"24",X"35",
		X"0C",X"32",X"30",X"37",X"24",X"34",X"0C",X"34",X"30",X"30",X"30",X"34",X"18",X"34",X"18",X"32",
		X"30",X"35",X"18",X"35",X"18",X"34",X"30",X"30",X"18",X"32",X"18",X"30",X"30",X"00",X"30",X"40",
		X"24",X"3B",X"0C",X"35",X"30",X"3B",X"24",X"39",X"0C",X"34",X"30",X"34",X"24",X"35",X"0C",X"40",
		X"30",X"00",X"60",X"35",X"24",X"37",X"0C",X"42",X"30",X"00",X"60",X"34",X"18",X"34",X"18",X"32",
		X"18",X"32",X"18",X"30",X"18",X"30",X"18",X"30",X"30",X"34",X"24",X"34",X"0C",X"30",X"30",X"32",
		X"24",X"32",X"0C",X"35",X"30",X"34",X"24",X"34",X"0C",X"30",X"30",X"30",X"24",X"32",X"0C",X"35",
		X"30",X"35",X"24",X"35",X"0C",X"32",X"30",X"30",X"24",X"30",X"0C",X"34",X"30",X"34",X"24",X"34",
		X"0C",X"30",X"30",X"32",X"24",X"32",X"0C",X"37",X"30",X"54",X"18",X"54",X"0C",X"54",X"0C",X"50",
		X"18",X"50",X"0C",X"50",X"0C",X"55",X"18",X"54",X"18",X"52",X"30",X"54",X"18",X"54",X"0C",X"54",
		X"0C",X"50",X"18",X"50",X"0C",X"50",X"0C",X"4B",X"0C",X"49",X"0C",X"4B",X"0C",X"50",X"0C",X"52",
		X"30",X"54",X"18",X"54",X"0C",X"54",X"0C",X"50",X"18",X"50",X"0C",X"50",X"0C",X"52",X"0C",X"54",
		X"0C",X"55",X"0C",X"57",X"0C",X"59",X"30",X"5B",X"18",X"5B",X"0C",X"5B",X"0C",X"57",X"18",X"57",
		X"0C",X"57",X"0C",X"60",X"0C",X"5B",X"0C",X"59",X"0C",X"5B",X"0C",X"60",X"30",X"60",X"18",X"59",
		X"18",X"55",X"18",X"57",X"18",X"5B",X"18",X"57",X"18",X"54",X"18",X"55",X"18",X"59",X"18",X"55",
		X"18",X"52",X"18",X"54",X"18",X"57",X"18",X"54",X"18",X"50",X"30",X"60",X"30",X"59",X"18",X"55",
		X"18",X"5B",X"18",X"5B",X"18",X"57",X"18",X"54",X"18",X"59",X"30",X"55",X"18",X"52",X"18",X"57",
		X"18",X"57",X"18",X"54",X"18",X"50",X"18",X"47",X"60",X"49",X"18",X"47",X"18",X"45",X"18",X"47",
		X"78",X"44",X"18",X"45",X"18",X"49",X"18",X"47",X"18",X"45",X"18",X"47",X"C0",X"00",X"60",X"FF",
		X"44",X"60",X"45",X"18",X"44",X"18",X"42",X"18",X"44",X"78",X"40",X"18",X"42",X"18",X"45",X"18",
		X"44",X"18",X"42",X"18",X"44",X"C0",X"00",X"60",X"40",X"60",X"40",X"60",X"40",X"60",X"40",X"60",
		X"40",X"30",X"40",X"30",X"40",X"78",X"00",X"60",X"78",X"D8",X"A2",X"FF",X"9A",X"AD",X"00",X"A0",
		X"A9",X"00",X"8D",X"00",X"C0",X"A0",X"00",X"A2",X"00",X"B9",X"00",X"F0",X"95",X"00",X"C8",X"E8",
		X"D0",X"F7",X"B9",X"00",X"F0",X"9D",X"00",X"01",X"C8",X"E8",X"D0",X"F6",X"B5",X"00",X"D9",X"00",
		X"F0",X"D0",X"4E",X"C8",X"E8",X"D0",X"F5",X"BD",X"00",X"01",X"D9",X"00",X"F0",X"D0",X"42",X"C8",
		X"E8",X"D0",X"F4",X"C8",X"C0",X"40",X"D0",X"CF",X"A2",X"00",X"BD",X"D9",X"FC",X"8D",X"00",X"40",
		X"E8",X"BD",X"D9",X"FC",X"8D",X"00",X"20",X"E8",X"E0",X"18",X"D0",X"EE",X"A2",X"00",X"A0",X"00",
		X"88",X"D0",X"FD",X"CA",X"D0",X"FA",X"4C",X"00",X"F0",X"00",X"66",X"01",X"01",X"02",X"1C",X"03",
		X"01",X"04",X"EF",X"05",X"00",X"07",X"F8",X"08",X"10",X"09",X"10",X"0A",X"10",X"0C",X"30",X"0D",
		X"09",X"A0",X"00",X"B9",X"12",X"FD",X"8D",X"00",X"40",X"C8",X"B9",X"12",X"FD",X"8D",X"00",X"20",
		X"C8",X"C0",X"18",X"D0",X"EE",X"A2",X"A0",X"A0",X"00",X"88",X"D0",X"FD",X"CA",X"D0",X"FA",X"4C",
		X"F1",X"FC",X"00",X"CC",X"01",X"02",X"02",X"A4",X"03",X"02",X"04",X"7E",X"05",X"02",X"07",X"38",
		X"08",X"10",X"09",X"10",X"0A",X"10",X"0C",X"30",X"0D",X"09",X"20",X"42",X"55",X"52",X"4E",X"49",
		X"4E",X"22",X"20",X"52",X"55",X"42",X"42",X"45",X"52",X"20",X"53",X"6F",X"75",X"6E",X"64",X"20",
		X"50",X"72",X"6F",X"67",X"72",X"61",X"6D",X"20",X"20",X"43",X"6F",X"70",X"79",X"72",X"69",X"67",
		X"68",X"74",X"20",X"31",X"39",X"38",X"32",X"20",X"28",X"63",X"29",X"20",X"44",X"41",X"54",X"41",
		X"20",X"45",X"41",X"53",X"54",X"20",X"63",X"6F",X"72",X"70",X"2E",X"20",X"20",X"70",X"72",X"6F",
		X"67",X"72",X"61",X"6D",X"65",X"64",X"20",X"62",X"79",X"20",X"54",X"2E",X"4B",X"69",X"74",X"61",
		X"7A",X"61",X"77",X"61",X"20",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"50",X"F5",X"78",X"FC",X"60",X"F0");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
