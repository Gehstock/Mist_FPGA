library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity bwidow_vec_rom4 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of bwidow_vec_rom4 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"08",X"5E",X"3A",X"40",X"3C",X"5D",X"06",X"5B",X"05",X"5A",X"23",X"44",X"20",X"46",X"02",X"58",
		X"22",X"44",X"3F",X"45",X"01",X"44",X"24",X"5C",X"25",X"42",X"13",X"41",X"00",X"C0",X"02",X"43",
		X"3D",X"46",X"25",X"43",X"1A",X"58",X"3C",X"42",X"3C",X"41",X"06",X"5B",X"3B",X"42",X"3B",X"5F",
		X"03",X"58",X"03",X"59",X"24",X"43",X"22",X"45",X"1F",X"58",X"23",X"43",X"22",X"45",X"02",X"45",
		X"23",X"59",X"24",X"40",X"15",X"46",X"00",X"C0",X"03",X"42",X"21",X"46",X"24",X"42",X"18",X"5A",
		X"3D",X"44",X"3C",X"42",X"04",X"59",X"3C",X"44",X"3B",X"41",X"00",X"58",X"00",X"58",X"25",X"41",
		X"24",X"44",X"1C",X"59",X"24",X"42",X"23",X"44",X"03",X"42",X"21",X"5A",X"24",X"5E",X"18",X"4A",
		X"00",X"C0",X"04",X"41",X"23",X"45",X"24",X"40",X"17",X"5E",X"3E",X"45",X"3D",X"43",X"01",X"58",
		X"3E",X"45",X"3C",X"43",X"1D",X"59",X"1D",X"58",X"25",X"5F",X"25",X"42",X"1A",X"5B",X"24",X"41",
		X"24",X"42",X"04",X"41",X"3D",X"5A",X"25",X"5D",X"1C",X"4C",X"00",X"C0",X"04",X"41",X"24",X"42",
		X"25",X"5E",X"16",X"42",X"21",X"45",X"3E",X"44",X"1E",X"58",X"20",X"46",X"3D",X"44",X"1B",X"5A",
		X"1A",X"5B",X"24",X"5D",X"26",X"40",X"18",X"5E",X"24",X"5E",X"25",X"41",X"02",X"5F",X"3E",X"5C",
		X"22",X"5B",X"01",X"4D",X"00",X"C0",X"03",X"5E",X"26",X"43",X"23",X"5B",X"18",X"46",X"22",X"44",
		X"21",X"44",X"1B",X"5A",X"22",X"45",X"3F",X"45",X"18",X"5D",X"19",X"5D",X"23",X"5C",X"25",X"5E",
		X"18",X"41",X"23",X"5D",X"25",X"5E",X"03",X"5E",X"3B",X"5D",X"20",X"5C",X"06",X"4B",X"00",X"C0",
		X"02",X"5D",X"26",X"5F",X"22",X"5C",X"1A",X"48",X"24",X"43",X"22",X"44",X"19",X"5C",X"24",X"44",
		X"21",X"45",X"18",X"40",X"18",X"40",X"21",X"5B",X"24",X"5C",X"19",X"44",X"22",X"5C",X"24",X"5D",
		X"02",X"5D",X"3A",X"5F",X"3E",X"5C",X"0A",X"48",X"00",X"C0",X"1F",X"5C",X"27",X"5D",X"20",X"5C",
		X"1E",X"49",X"25",X"42",X"23",X"43",X"18",X"5F",X"25",X"42",X"23",X"44",X"19",X"43",X"18",X"43",
		X"3F",X"5B",X"22",X"5B",X"1B",X"46",X"21",X"5C",X"22",X"5C",X"01",X"5C",X"3A",X"43",X"3D",X"5B",
		X"0C",X"44",X"00",X"C0",X"1F",X"5C",X"24",X"5C",X"3E",X"5B",X"02",X"4A",X"25",X"5F",X"24",X"42",
		X"18",X"42",X"26",X"40",X"24",X"43",X"1A",X"45",X"1B",X"46",X"3D",X"5C",X"20",X"5A",X"1E",X"48",
		X"3E",X"5C",X"21",X"5B",X"1F",X"5E",X"3C",X"42",X"3B",X"5E",X"0D",X"5F",X"00",X"C0",X"1E",X"5D",
		X"21",X"5A",X"3D",X"5D",X"06",X"48",X"24",X"5E",X"24",X"5F",X"1A",X"45",X"25",X"5E",X"25",X"41",
		X"1D",X"48",X"1D",X"47",X"3C",X"5D",X"3E",X"5B",X"01",X"48",X"3D",X"5D",X"3E",X"5B",X"1E",X"5D",
		X"3D",X"45",X"3C",X"40",X"0B",X"5A",X"00",X"C0",X"1D",X"5E",X"3F",X"5A",X"3C",X"5E",X"08",X"46",
		X"23",X"5C",X"24",X"5E",X"1C",X"47",X"24",X"5C",X"25",X"5F",X"00",X"48",X"00",X"48",X"3B",X"5F",
		X"3C",X"5C",X"04",X"47",X"3C",X"5E",X"3D",X"5C",X"1D",X"5E",X"3F",X"46",X"3C",X"42",X"08",X"56",
		X"00",X"C0",X"1C",X"41",X"3D",X"59",X"3C",X"40",X"09",X"42",X"22",X"5B",X"23",X"5D",X"1F",X"48",
		X"22",X"5B",X"24",X"5D",X"03",X"47",X"03",X"48",X"3B",X"41",X"3B",X"5E",X"06",X"45",X"3C",X"5F",
		X"3C",X"5E",X"1C",X"5F",X"21",X"46",X"3D",X"43",X"04",X"54",X"00",X"C0",X"1C",X"41",X"3C",X"5C",
		X"3B",X"42",X"0A",X"5E",X"3F",X"5B",X"22",X"5C",X"02",X"48",X"20",X"5A",X"23",X"5C",X"05",X"46",
		X"06",X"45",X"3C",X"43",X"3A",X"40",X"08",X"42",X"3C",X"42",X"3B",X"5F",X"1C",X"41",X"24",X"44",
		X"3E",X"45",X"1F",X"53",X"00",X"C0",X"1D",X"42",X"3A",X"5F",X"3D",X"43",X"08",X"5A",X"3E",X"5C",
		X"3F",X"5C",X"05",X"46",X"3E",X"5B",X"21",X"5B",X"08",X"43",X"07",X"43",X"3D",X"44",X"3B",X"42",
		X"08",X"5F",X"3D",X"43",X"3B",X"42",X"1B",X"42",X"27",X"43",X"20",X"44",X"1A",X"55",X"00",X"C0",
		X"1E",X"43",X"36",X"57",X"3F",X"5C",X"27",X"5E",X"26",X"4C",X"26",X"54",X"27",X"42",X"3F",X"44",
		X"36",X"49",X"1E",X"5D",X"00",X"C0",X"1F",X"44",X"34",X"5D",X"3D",X"5B",X"26",X"5B",X"2A",X"49",
		X"3F",X"53",X"29",X"5F",X"21",X"44",X"3A",X"4C",X"1D",X"5E",X"00",X"C0",X"1F",X"44",X"34",X"40",
		X"3D",X"5E",X"23",X"5A",X"2D",X"44",X"3C",X"53",X"26",X"5D",X"22",X"43",X"20",X"4E",X"1C",X"5F",
		X"00",X"C0",X"02",X"43",X"34",X"46",X"3C",X"5F",X"21",X"59",X"2D",X"5F",X"37",X"56",X"25",X"5A",
		X"23",X"43",X"25",X"4E",X"1C",X"5F",X"00",X"C0",X"03",X"42",X"37",X"4A",X"3C",X"41",X"3E",X"59",
		X"2C",X"5A",X"34",X"5A",X"22",X"59",X"24",X"41",X"29",X"4A",X"1D",X"42",X"00",X"C0",X"04",X"41",
		X"3B",X"4C",X"3D",X"43",X"3B",X"5A",X"29",X"56",X"33",X"41",X"3F",X"57",X"24",X"5F",X"2C",X"46",
		X"1E",X"43",X"00",X"C0",X"04",X"41",X"20",X"4C",X"3E",X"43",X"3A",X"5D",X"24",X"53",X"33",X"44",
		X"3D",X"5A",X"23",X"5E",X"2C",X"40",X"01",X"44",X"00",X"C0",X"03",X"5E",X"26",X"4C",X"3F",X"44",
		X"37",X"5F",X"21",X"53",X"36",X"49",X"3A",X"5B",X"23",X"5D",X"2C",X"5B",X"01",X"44",X"00",X"C0",
		X"02",X"5D",X"2A",X"49",X"21",X"44",X"39",X"42",X"3A",X"54",X"3A",X"4C",X"39",X"5E",X"21",X"5C",
		X"2A",X"57",X"02",X"43",X"00",X"C0",X"1F",X"5C",X"2E",X"45",X"23",X"43",X"3A",X"45",X"36",X"57",
		X"3F",X"4D",X"39",X"41",X"3F",X"5C",X"26",X"54",X"03",X"42",X"00",X"C0",X"1F",X"5C",X"2E",X"40",
		X"23",X"42",X"3D",X"46",X"33",X"5C",X"24",X"4D",X"3A",X"43",X"3E",X"5D",X"20",X"54",X"04",X"5F",
		X"00",X"C0",X"1E",X"5D",X"2C",X"5A",X"24",X"41",X"3F",X"49",X"33",X"5F",X"29",X"4A",X"3B",X"46",
		X"3B",X"5D",X"3D",X"54",X"04",X"5F",X"00",X"C0",X"1D",X"5E",X"29",X"56",X"24",X"5F",X"22",X"47",
		X"34",X"46",X"2C",X"46",X"3E",X"47",X"3C",X"5F",X"37",X"56",X"03",X"5E",X"00",X"C0",X"1C",X"41",
		X"23",X"52",X"25",X"5D",X"25",X"46",X"37",X"4A",X"2D",X"41",X"21",X"47",X"3C",X"41",X"34",X"5A",
		X"02",X"5D",X"00",X"C0",X"1C",X"41",X"20",X"52",X"22",X"5D",X"26",X"43",X"3C",X"4D",X"2D",X"5C",
		X"23",X"46",X"3D",X"42",X"32",X"40",X"01",X"5C",X"00",X"C0",X"1D",X"42",X"3A",X"54",X"21",X"5C",
		X"27",X"41",X"21",X"4D",X"2A",X"57",X"26",X"45",X"3D",X"45",X"32",X"43",X"01",X"5C",X"00",X"C0",
		X"1E",X"43",X"34",X"5A",X"3F",X"5C",X"27",X"5E",X"28",X"49",X"28",X"57",X"27",X"42",X"3F",X"44",
		X"34",X"46",X"1E",X"5D",X"00",X"C0",X"1F",X"44",X"33",X"5F",X"3D",X"5E",X"26",X"5A",X"2B",X"45",
		X"24",X"55",X"27",X"5F",X"21",X"44",X"37",X"4A",X"1D",X"5E",X"00",X"C0",X"1F",X"44",X"35",X"44",
		X"3C",X"5E",X"24",X"5B",X"2C",X"5F",X"3F",X"54",X"27",X"5C",X"22",X"44",X"3C",X"4D",X"1C",X"5F",
		X"00",X"C0",X"02",X"43",X"36",X"49",X"3C",X"5F",X"21",X"59",X"2B",X"5C",X"3B",X"55",X"24",X"5A",
		X"24",X"43",X"21",X"4F",X"1C",X"5F",X"00",X"C0",X"03",X"42",X"3A",X"4C",X"3C",X"41",X"3E",X"59",
		X"29",X"58",X"37",X"58",X"22",X"59",X"24",X"41",X"26",X"4C",X"1D",X"42",X"00",X"C0",X"04",X"41",
		X"3F",X"4D",X"3C",X"43",X"3C",X"5A",X"25",X"55",X"35",X"5C",X"3F",X"59",X"24",X"5F",X"2A",X"49",
		X"1E",X"43",X"00",X"C0",X"04",X"41",X"24",X"4B",X"3E",X"44",X"39",X"5C",X"21",X"54",X"34",X"41",
		X"3C",X"59",X"24",X"5E",X"2B",X"44",X"01",X"44",X"00",X"C0",X"03",X"5E",X"29",X"4A",X"3F",X"44",
		X"39",X"5F",X"3C",X"55",X"35",X"45",X"3A",X"5C",X"23",X"5C",X"2D",X"5F",X"01",X"44",X"00",X"C0",
		X"02",X"5D",X"2C",X"46",X"21",X"44",X"39",X"42",X"38",X"57",X"38",X"49",X"39",X"5E",X"21",X"5C",
		X"2C",X"5A",X"02",X"43",X"00",X"C0",X"1F",X"5C",X"2F",X"41",X"23",X"44",X"3A",X"44",X"35",X"5B",
		X"3C",X"4B",X"39",X"41",X"3F",X"5C",X"29",X"56",X"03",X"42",X"00",X"C0",X"1F",X"5C",X"2D",X"5C",
		X"24",X"42",X"3C",X"47",X"34",X"5F",X"3F",X"4C",X"3B",X"44",X"3E",X"5C",X"24",X"55",X"04",X"5F",
		X"00",X"C0",X"1E",X"5D",X"2A",X"57",X"24",X"41",X"3F",X"47",X"35",X"44",X"25",X"4B",X"3A",X"46",
		X"3E",X"5D",X"3F",X"53",X"04",X"5F",X"00",X"C0",X"1D",X"5E",X"26",X"54",X"24",X"5F",X"22",X"47",
		X"37",X"48",X"29",X"48",X"3E",X"47",X"3C",X"5F",X"3A",X"54",X"03",X"5E",X"00",X"C0",X"1C",X"41",
		X"21",X"51",X"22",X"5D",X"26",X"46",X"3B",X"4B",X"2B",X"44",X"21",X"47",X"3C",X"41",X"36",X"57",
		X"02",X"5D",X"00",X"C0",X"1C",X"41",X"3C",X"53",X"22",X"5C",X"25",X"44",X"21",X"4C",X"2C",X"41",
		X"24",X"45",X"3C",X"42",X"33",X"5C",X"01",X"5C",X"00",X"C0",X"1D",X"42",X"37",X"56",X"21",X"5C",
		X"27",X"41",X"24",X"4B",X"2B",X"5B",X"26",X"46",X"3D",X"42",X"31",X"41",X"01",X"5C",X"00",X"C0",
		X"1E",X"43",X"33",X"5D",X"3E",X"5C",X"26",X"5D",X"2B",X"47",X"2B",X"59",X"26",X"43",X"3E",X"44",
		X"33",X"43",X"1E",X"5D",X"00",X"C0",X"1F",X"44",X"33",X"42",X"3D",X"5D",X"24",X"5B",X"2D",X"42",
		X"27",X"55",X"27",X"41",X"20",X"44",X"35",X"48",X"1D",X"5E",X"00",X"C0",X"FE",X"00",X"1F",X"44",
		X"36",X"47",X"3C",X"5E",X"22",X"5A",X"2D",X"5D",X"23",X"53",X"26",X"5E",X"22",X"44",X"39",X"4C",
		X"1C",X"5F",X"00",X"C0",X"02",X"43",X"38",X"4B",X"3C",X"40",X"3F",X"59",X"2B",X"59",X"3E",X"53",
		X"25",X"5C",X"23",X"43",X"3E",X"4F",X"1C",X"5F",X"00",X"C0",X"03",X"42",X"3D",X"4D",X"3C",X"42",
		X"3D",X"5A",X"27",X"55",X"39",X"55",X"23",X"5A",X"24",X"42",X"23",X"4D",X"1D",X"42",X"00",X"C0",
		X"04",X"41",X"22",X"4D",X"3D",X"43",X"3B",X"5C",X"22",X"53",X"35",X"59",X"21",X"59",X"24",X"40",
		X"28",X"4B",X"1E",X"43",X"00",X"C0",X"04",X"41",X"27",X"4A",X"3E",X"44",X"3A",X"5E",X"3D",X"53",
		X"33",X"5D",X"3E",X"5A",X"24",X"5E",X"2A",X"47",X"01",X"44",X"00",X"C0",X"03",X"5E",X"2B",X"48",
		X"20",X"44",X"39",X"41",X"39",X"55",X"33",X"42",X"3C",X"5B",X"23",X"5D",X"2D",X"42",X"01",X"44",
		X"00",X"C0",X"02",X"5D",X"2D",X"43",X"22",X"44",X"3A",X"43",X"35",X"59",X"35",X"47",X"3A",X"5D",
		X"22",X"5C",X"2D",X"5D",X"02",X"43",X"00",X"C0",X"1F",X"5C",X"2F",X"5E",X"23",X"43",X"3C",X"45",
		X"33",X"5E",X"39",X"4B",X"39",X"5F",X"20",X"5C",X"2B",X"58",X"03",X"42",X"00",X"C0",X"1F",X"5C",
		X"2C",X"59",X"24",X"42",X"3E",X"46",X"33",X"43",X"3D",X"4D",X"3A",X"42",X"3E",X"5C",X"27",X"56",
		X"04",X"5F",X"00",X"C0",X"1E",X"5D",X"28",X"55",X"24",X"40",X"21",X"47",X"35",X"47",X"22",X"4D",
		X"3B",X"44",X"3D",X"5D",X"22",X"53",X"04",X"5F",X"00",X"C0",X"1D",X"5E",X"23",X"53",X"24",X"5E",
		X"23",X"46",X"39",X"4B",X"27",X"4B",X"3D",X"46",X"3C",X"5E",X"3D",X"53",X"03",X"5E",X"00",X"C0",
		X"1C",X"41",X"3E",X"51",X"23",X"5D",X"25",X"44",X"3E",X"4D",X"2B",X"47",X"3F",X"47",X"3C",X"40",
		X"38",X"55",X"02",X"5D",X"00",X"C0",X"1C",X"41",X"39",X"54",X"22",X"5C",X"26",X"42",X"23",X"4D",
		X"2D",X"43",X"22",X"46",X"3C",X"42",X"34",X"59",X"01",X"5C",X"00",X"C0",X"1D",X"42",X"35",X"58",
		X"20",X"5C",X"27",X"5F",X"27",X"4B",X"2D",X"5E",X"24",X"45",X"3D",X"43",X"31",X"5E",X"01",X"5C",
		X"00",X"C0",X"A0",X"A7",X"60",X"A7",X"39",X"BB",X"8B",X"BB",X"E3",X"BB",X"39",X"BC",X"AE",X"BC",
		X"4D",X"BD",X"00",X"60",X"3F",X"5F",X"C4",X"60",X"24",X"40",X"22",X"5F",X"21",X"5E",X"20",X"5F",
		X"3B",X"5E",X"3B",X"42",X"20",X"41",X"21",X"42",X"22",X"41",X"87",X"60",X"3D",X"40",X"3D",X"5F",
		X"3F",X"5F",X"39",X"40",X"3C",X"43",X"20",X"42",X"C4",X"60",X"29",X"45",X"29",X"40",X"22",X"5F",
		X"22",X"41",X"29",X"40",X"29",X"5B",X"87",X"60",X"20",X"5E",X"3C",X"5D",X"35",X"40",X"00",X"60",
		X"3B",X"4F",X"C4",X"60",X"37",X"BD",X"C4",X"60",X"24",X"44",X"23",X"41",X"00",X"60",X"3F",X"5E",
		X"C4",X"60",X"3F",X"40",X"3B",X"5D",X"00",X"60",X"D6",X"1F",X"F8",X"3F",X"C2",X"60",X"3F",X"41",
		X"3F",X"5F",X"3F",X"40",X"3E",X"43",X"3F",X"40",X"3F",X"5F",X"00",X"60",X"22",X"5E",X"C2",X"60",
		X"21",X"5F",X"21",X"40",X"00",X"60",X"33",X"4C",X"C2",X"60",X"21",X"40",X"21",X"5E",X"23",X"40",
		X"21",X"42",X"3B",X"40",X"00",X"60",X"25",X"40",X"87",X"60",X"2F",X"40",X"C2",X"60",X"21",X"5E",
		X"23",X"40",X"21",X"42",X"3B",X"40",X"00",X"60",X"25",X"40",X"87",X"60",X"2E",X"40",X"00",X"60",
		X"FC",X"1F",X"D8",X"3F",X"00",X"C0",X"00",X"60",X"20",X"4C",X"C4",X"60",X"21",X"43",X"22",X"43",
		X"22",X"40",X"00",X"60",X"3F",X"5E",X"C4",X"60",X"3F",X"40",X"3D",X"5C",X"37",X"BD",X"00",X"60",
		X"EC",X"1F",X"28",X"20",X"C4",X"60",X"3C",X"43",X"38",X"44",X"3D",X"40",X"3D",X"5F",X"3E",X"5E",
		X"3E",X"42",X"3D",X"41",X"3D",X"40",X"38",X"5C",X"3C",X"5D",X"87",X"60",X"2F",X"43",X"25",X"5E",
		X"25",X"42",X"2F",X"5D",X"00",X"60",X"34",X"5A",X"C2",X"60",X"21",X"41",X"20",X"41",X"3F",X"41",
		X"3E",X"40",X"3F",X"5F",X"00",X"60",X"36",X"40",X"C2",X"60",X"3F",X"41",X"3E",X"40",X"3F",X"5F",
		X"20",X"5F",X"21",X"5F",X"00",X"60",X"34",X"46",X"87",X"60",X"20",X"5E",X"28",X"5C",X"24",X"40",
		X"24",X"42",X"00",X"60",X"28",X"40",X"87",X"60",X"24",X"5E",X"24",X"40",X"28",X"44",X"20",X"42",
		X"00",X"60",X"F8",X"1F",X"E0",X"3F",X"C4",X"60",X"21",X"5E",X"20",X"5F",X"3B",X"5E",X"3B",X"42",
		X"20",X"41",X"21",X"42",X"22",X"41",X"24",X"40",X"22",X"5F",X"00",X"60",X"3E",X"59",X"C2",X"60",
		X"3F",X"40",X"3F",X"5F",X"3F",X"40",X"3D",X"42",X"3E",X"5F",X"00",X"60",X"22",X"5F",X"C2",X"60",
		X"21",X"5F",X"22",X"40",X"00",X"C0",X"00",X"60",X"20",X"4C",X"C4",X"60",X"20",X"43",X"22",X"43",
		X"22",X"41",X"00",X"60",X"3F",X"5D",X"C4",X"60",X"3E",X"5F",X"3F",X"5D",X"37",X"BD",X"00",X"60",
		X"20",X"5A",X"C4",X"60",X"23",X"43",X"25",X"40",X"28",X"5C",X"24",X"5D",X"87",X"60",X"34",X"45",
		X"3B",X"40",X"3D",X"5E",X"3D",X"42",X"3B",X"40",X"34",X"5B",X"C4",X"60",X"24",X"43",X"28",X"44",
		X"25",X"40",X"23",X"5D",X"00",X"60",X"25",X"57",X"C2",X"60",X"20",X"41",X"21",X"41",X"22",X"40",
		X"21",X"5E",X"3F",X"5F",X"00",X"60",X"33",X"41",X"C2",X"60",X"20",X"41",X"3F",X"41",X"3E",X"40",
		X"3F",X"5E",X"21",X"5F",X"00",X"60",X"23",X"41",X"87",X"60",X"3C",X"5E",X"3D",X"40",X"3D",X"41",
		X"3B",X"44",X"20",X"42",X"00",X"60",X"00",X"00",X"50",X"20",X"87",X"60",X"20",X"5E",X"3B",X"5C",
		X"3D",X"5F",X"3D",X"40",X"3C",X"42",X"C4",X"60",X"20",X"5E",X"3B",X"5E",X"3B",X"42",X"20",X"42",
		X"22",X"42",X"26",X"40",X"22",X"5E",X"00",X"60",X"20",X"59",X"C2",X"60",X"3E",X"5F",X"3D",X"41",
		X"3D",X"5F",X"3E",X"41",X"00",X"60",X"23",X"5E",X"C2",X"60",X"24",X"40",X"00",X"60",X"3E",X"4C",
		X"00",X"C0",X"00",X"60",X"20",X"4F",X"C4",X"60",X"20",X"44",X"21",X"43",X"00",X"60",X"21",X"5E",
		X"C4",X"60",X"3F",X"5E",X"3F",X"5D",X"23",X"40",X"27",X"5D",X"25",X"5D",X"26",X"5A",X"21",X"5D",
		X"22",X"41",X"00",X"60",X"3E",X"5F",X"C4",X"60",X"20",X"5E",X"3B",X"59",X"32",X"5A",X"3A",X"40",
		X"32",X"46",X"3B",X"47",X"20",X"42",X"3E",X"41",X"00",X"60",X"22",X"5F",X"C4",X"60",X"21",X"43",
		X"26",X"46",X"25",X"43",X"27",X"43",X"23",X"40",X"00",X"60",X"20",X"5D",X"87",X"60",X"3E",X"41",
		X"3E",X"40",X"3B",X"5E",X"39",X"5A",X"3E",X"5D",X"20",X"5D",X"23",X"5E",X"23",X"5E",X"22",X"40",
		X"25",X"41",X"00",X"60",X"2A",X"40",X"87",X"60",X"25",X"5F",X"22",X"40",X"23",X"42",X"23",X"42",
		X"20",X"43",X"3E",X"43",X"39",X"46",X"3B",X"42",X"3E",X"40",X"3E",X"5F",X"00",X"60",X"23",X"53",
		X"C2",X"60",X"21",X"41",X"22",X"40",X"21",X"5F",X"20",X"5E",X"3E",X"5F",X"3F",X"41",X"00",X"60",
		X"38",X"40",X"C2",X"60",X"3F",X"5F",X"3E",X"41",X"20",X"42",X"21",X"41",X"22",X"40",X"21",X"5F",
		X"C4",X"60",X"22",X"42",X"22",X"40",X"22",X"5E",X"21",X"5F",X"20",X"5D",X"3C",X"5E",X"3C",X"42",
		X"20",X"43",X"21",X"41",X"00",X"60",X"3F",X"57",X"C2",X"60",X"23",X"41",X"22",X"40",X"23",X"5F",
		X"20",X"5F",X"3D",X"5E",X"3E",X"40",X"3D",X"42",X"20",X"41",X"00",X"60",X"21",X"5E",X"C4",X"60",
		X"21",X"41",X"21",X"40",X"21",X"5F",X"21",X"41",X"21",X"40",X"21",X"5F",X"00",X"60",X"21",X"5F",
		X"3E",X"5F",X"3C",X"40",X"3E",X"41",X"00",X"60",X"24",X"4D",X"00",X"C0",X"00",X"60",X"26",X"00",
		X"00",X"20",X"C4",X"60",X"3F",X"48",X"00",X"60",X"22",X"5E",X"C4",X"60",X"3F",X"5A",X"21",X"40",
		X"24",X"5F",X"24",X"5D",X"2A",X"52",X"21",X"5E",X"24",X"42",X"00",X"60",X"3C",X"5E",X"C4",X"60",
		X"20",X"5D",X"3C",X"59",X"35",X"59",X"3C",X"5E",X"3E",X"40",X"3C",X"42",X"35",X"47",X"3C",X"47",
		X"20",X"43",X"3C",X"42",X"00",X"60",X"24",X"5E",X"C4",X"60",X"21",X"42",X"2A",X"4E",X"24",X"43",
		X"24",X"41",X"21",X"40",X"00",X"60",X"3F",X"5F",X"87",X"60",X"21",X"5F",X"21",X"41",X"00",X"60",
		X"3F",X"5C",X"87",X"60",X"3E",X"42",X"3E",X"40",X"3D",X"5E",X"3B",X"57",X"3E",X"5B",X"20",X"5C",
		X"23",X"5C",X"22",X"40",X"27",X"44",X"00",X"60",X"24",X"40",X"87",X"60",X"27",X"5C",X"22",X"40",
		X"23",X"44",X"20",X"44",X"3E",X"45",X"3B",X"49",X"3D",X"42",X"3E",X"40",X"3E",X"5E",X"00",X"60",
		X"DC",X"1F",X"04",X"20",X"C2",X"60",X"20",X"42",X"21",X"41",X"21",X"40",X"21",X"5F",X"20",X"5E",
		X"3F",X"5F",X"00",X"60",X"22",X"5F",X"C5",X"60",X"22",X"42",X"20",X"43",X"3D",X"43",X"3E",X"40",
		X"3E",X"5E",X"00",X"60",X"3E",X"40",X"C5",X"60",X"3E",X"42",X"3E",X"40",X"3D",X"5D",X"20",X"5D",
		X"22",X"5E",X"00",X"60",X"22",X"41",X"C2",X"60",X"3F",X"41",X"20",X"42",X"21",X"41",X"21",X"40",
		X"21",X"5F",X"20",X"5E",X"C4",X"60",X"21",X"44",X"21",X"41",X"21",X"5F",X"21",X"5C",X"20",X"5D",
		X"3E",X"5D",X"3E",X"43",X"20",X"43",X"00",X"60",X"21",X"5A",X"C2",X"60",X"22",X"40",X"24",X"5B",
		X"20",X"5F",X"3E",X"40",X"3E",X"41",X"3E",X"40",X"3E",X"5F",X"3E",X"40",X"20",X"41",X"24",X"45",
		X"00",X"60",X"3E",X"5A",X"C4",X"60",X"3F",X"41",X"21",X"42",X"22",X"40",X"21",X"5F",X"21",X"41",
		X"22",X"40",X"21",X"5E",X"3F",X"5F",X"00",X"60",X"20",X"00",X"FA",X"3F",X"00",X"C0",X"25",X"40",
		X"26",X"5E",X"27",X"5C",X"23",X"5E",X"24",X"5B",X"20",X"5E",X"3D",X"5D",X"39",X"5C",X"3B",X"5E",
		X"3B",X"5F",X"36",X"40",X"3B",X"41",X"3B",X"42",X"39",X"44",X"3D",X"43",X"20",X"42",X"24",X"45",
		X"23",X"42",X"27",X"44",X"26",X"42",X"25",X"40",X"00",X"C0",X"00",X"60",X"02",X"00",X"D0",X"3F",
		X"C4",X"60",X"36",X"5C",X"DA",X"1F",X"16",X"20",X"3F",X"40",X"26",X"00",X"E2",X"3F",X"21",X"43",
		X"2A",X"44",X"24",X"5D",X"00",X"60",X"3C",X"43",X"C4",X"60",X"3F",X"41",X"37",X"44",X"DA",X"1F",
		X"EA",X"3F",X"3F",X"40",X"2C",X"00",X"12",X"20",X"23",X"42",X"27",X"5D",X"20",X"5E",X"22",X"5C",
		X"00",X"60",X"3E",X"46",X"C4",X"60",X"20",X"41",X"21",X"42",X"3C",X"45",X"E4",X"1F",X"DE",X"3F",
		X"3F",X"40",X"24",X"00",X"24",X"20",X"23",X"40",X"25",X"5A",X"3D",X"5D",X"00",X"60",X"23",X"43",
		X"C4",X"60",X"23",X"43",X"2A",X"45",X"29",X"42",X"2A",X"40",X"29",X"5E",X"2A",X"5B",X"26",X"5A",
		X"00",X"60",X"3D",X"43",X"C4",X"60",X"25",X"46",X"23",X"40",X"DC",X"1F",X"24",X"20",X"3F",X"40",
		X"1C",X"00",X"DE",X"3F",X"3C",X"5B",X"21",X"5E",X"20",X"5F",X"00",X"60",X"3E",X"5A",X"C4",X"60",
		X"22",X"44",X"20",X"42",X"27",X"43",X"23",X"5E",X"D4",X"1F",X"12",X"20",X"3F",X"40",X"26",X"00",
		X"EA",X"3F",X"37",X"5C",X"3F",X"5F",X"3C",X"5D",X"00",X"60",X"24",X"43",X"C4",X"60",X"2A",X"5C",
		X"21",X"5D",X"DA",X"1F",X"E2",X"3F",X"3F",X"40",X"26",X"00",X"16",X"20",X"36",X"44",X"00",X"60",
		X"FE",X"1F",X"D0",X"3F",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"48",X"24",X"44",X"24",X"5C",X"20",X"58",X"18",X"44",X"28",X"40",X"04",X"5C",X"00",X"C0",
		X"20",X"4C",X"26",X"40",X"22",X"5E",X"20",X"5E",X"3E",X"5E",X"3A",X"40",X"06",X"40",X"22",X"5E",
		X"20",X"5E",X"3E",X"5E",X"3A",X"40",X"52",X"FE",X"20",X"4C",X"28",X"40",X"18",X"54",X"95",X"FE",
		X"20",X"4C",X"24",X"40",X"24",X"5C",X"20",X"5C",X"3C",X"5C",X"3C",X"40",X"52",X"FE",X"28",X"40",
		X"18",X"40",X"20",X"4C",X"28",X"40",X"1E",X"5A",X"3A",X"40",X"0C",X"5A",X"00",X"C0",X"20",X"4C",
		X"28",X"40",X"20",X"5C",X"1C",X"5C",X"24",X"40",X"20",X"5C",X"51",X"FE",X"20",X"4C",X"00",X"5A",
		X"28",X"40",X"00",X"46",X"AE",X"FE",X"28",X"40",X"18",X"4C",X"28",X"40",X"1C",X"40",X"20",X"54",
		X"08",X"40",X"00",X"C0",X"00",X"44",X"24",X"5C",X"24",X"40",X"73",X"FE",X"20",X"4C",X"06",X"40",
		X"3A",X"5A",X"26",X"5A",X"06",X"40",X"00",X"C0",X"00",X"4C",X"20",X"54",X"95",X"FE",X"20",X"4C",
		X"24",X"5C",X"24",X"44",X"AE",X"FE",X"20",X"4C",X"28",X"54",X"73",X"FE",X"20",X"4C",X"28",X"40",
		X"20",X"54",X"38",X"40",X"0C",X"40",X"00",X"C0",X"20",X"4C",X"28",X"40",X"20",X"5A",X"38",X"40",
		X"25",X"FE",X"20",X"4C",X"28",X"40",X"20",X"58",X"3C",X"5C",X"3C",X"40",X"04",X"44",X"24",X"5C",
		X"96",X"FE",X"20",X"4C",X"28",X"40",X"20",X"5A",X"38",X"40",X"02",X"40",X"26",X"5A",X"96",X"FE",
		X"28",X"40",X"20",X"46",X"38",X"40",X"20",X"46",X"28",X"40",X"74",X"FE",X"00",X"4C",X"35",X"FE",
		X"00",X"4C",X"20",X"54",X"28",X"40",X"20",X"4C",X"04",X"54",X"00",X"C0",X"00",X"4C",X"24",X"54",
		X"24",X"4C",X"74",X"FE",X"00",X"4C",X"20",X"54",X"24",X"44",X"24",X"5C",X"73",X"FE",X"28",X"4C",
		X"18",X"40",X"28",X"54",X"AF",X"FE",X"04",X"40",X"20",X"48",X"3C",X"44",X"08",X"40",X"3C",X"5C",
		X"08",X"58",X"00",X"C0",X"00",X"4C",X"28",X"40",X"38",X"54",X"95",X"FE",X"04",X"4C",X"37",X"FE",
		X"00",X"4C",X"28",X"40",X"20",X"5A",X"38",X"40",X"20",X"5A",X"28",X"40",X"04",X"40",X"00",X"C0",
		X"00",X"4C",X"28",X"40",X"20",X"54",X"38",X"40",X"00",X"46",X"28",X"40",X"04",X"5A",X"00",X"C0",
		X"00",X"4C",X"20",X"5A",X"28",X"40",X"00",X"46",X"AE",X"FE",X"00",X"46",X"28",X"40",X"20",X"5A",
		X"38",X"40",X"20",X"4C",X"0C",X"54",X"00",X"C0",X"00",X"4C",X"28",X"40",X"20",X"54",X"04",X"40",
		X"00",X"C0",X"20",X"4C",X"99",X"FE",X"08",X"46",X"38",X"40",X"20",X"46",X"AD",X"FE",X"A9",X"FF",
		X"95",X"FE",X"05",X"00",X"02",X"00",X"21",X"43",X"3E",X"42",X"23",X"40",X"05",X"00",X"02",X"20",
		X"FB",X"1F",X"02",X"20",X"23",X"40",X"3E",X"5E",X"21",X"5D",X"03",X"00",X"FA",X"3F",X"FD",X"1F",
		X"FA",X"3F",X"FB",X"1F",X"0E",X"00",X"04",X"40",X"00",X"C0",X"00",X"42",X"20",X"48",X"22",X"42",
		X"24",X"40",X"22",X"5E",X"20",X"58",X"3E",X"5E",X"3C",X"40",X"3E",X"42",X"06",X"42",X"3C",X"40",
		X"20",X"44",X"24",X"40",X"06",X"58",X"00",X"C0",X"00",X"46",X"28",X"46",X"20",X"54",X"38",X"46",
		X"0C",X"5A",X"00",X"C0",X"52",X"BE",X"4E",X"BE",X"8E",X"BE",X"90",X"BE",X"98",X"BE",X"A0",X"BE",
		X"68",X"BE",X"A5",X"BE",X"AC",X"BE",X"B1",X"BE",X"B3",X"BE",X"00",X"BE",X"08",X"BE",X"14",X"BE",
		X"18",X"BE",X"1F",X"BE",X"21",X"BE",X"27",X"BE",X"2E",X"BE",X"33",X"BE",X"3A",X"BE",X"3E",X"BE",
		X"44",X"BE",X"47",X"BE",X"4B",X"BE",X"4E",X"BE",X"54",X"BE",X"59",X"BE",X"61",X"BE",X"68",X"BE",
		X"6E",X"BE",X"70",X"BE",X"76",X"BE",X"7A",X"BE",X"7F",X"BE",X"83",X"BE",X"8A",X"BE",X"B9",X"BE",
		X"B8",X"BE",X"B7",X"BE",X"CD",X"BE",X"DC",X"BE",X"00",X"C0",X"40",X"80",X"00",X"71",X"00",X"C0",
		X"0D",X"BF",X"5E",X"1E",X"3E",X"1E",X"00",X"00",X"84",X"23",X"48",X"03",X"00",X"20",X"00",X"00",
		X"7C",X"3C",X"B8",X"1C",X"00",X"20",X"00",X"C0",X"5E",X"1E",X"3E",X"1E",X"48",X"03",X"48",X"23",
		X"C4",X"1F",X"3C",X"20",X"F4",X"1C",X"F4",X"3C",X"78",X"00",X"88",X"3F",X"D0",X"02",X"D0",X"22",
		X"4C",X"1F",X"B4",X"20",X"6C",X"1D",X"6C",X"3D",X"F0",X"00",X"10",X"3F",X"58",X"02",X"58",X"22",
		X"D4",X"1E",X"2C",X"21",X"E4",X"1D",X"E4",X"3D",X"68",X"01",X"98",X"3E",X"E0",X"01",X"E0",X"21",
		X"5C",X"1E",X"A4",X"21",X"5C",X"1E",X"5C",X"3E",X"E0",X"01",X"20",X"3E",X"68",X"01",X"68",X"21",
		X"E4",X"1D",X"1C",X"22",X"D4",X"1E",X"D4",X"3E",X"58",X"02",X"A8",X"3D",X"F0",X"00",X"F0",X"20",
		X"6C",X"1D",X"94",X"22",X"4C",X"1F",X"4C",X"3F",X"D0",X"02",X"30",X"3D",X"78",X"00",X"78",X"20",
		X"F4",X"1C",X"0C",X"23",X"C4",X"1F",X"C4",X"3F",X"48",X"03",X"B8",X"3C",X"01",X"1E",X"00",X"00",
		X"14",X"71",X"E2",X"FE",X"10",X"00",X"00",X"1F",X"00",X"C0",X"00",X"00",X"00",X"E1",X"5A",X"BF",
		X"00",X"00",X"00",X"C1",X"5A",X"BF",X"00",X"00",X"00",X"A1",X"5A",X"BF",X"00",X"00",X"00",X"81",
		X"5A",X"BF",X"00",X"00",X"00",X"61",X"5A",X"BF",X"00",X"00",X"00",X"41",X"00",X"C0",X"17",X"60",
		X"00",X"00",X"40",X"40",X"10",X"00",X"C0",X"1E",X"00",X"00",X"00",X"21",X"00",X"C0",X"B8",X"1C",
		X"00",X"20",X"40",X"80",X"00",X"C0",X"00",X"00",X"84",X"23",X"40",X"80",X"00",X"C0",X"C7",X"60",
		X"40",X"80",X"1C",X"FF",X"99",X"BF",X"00",X"70",X"C0",X"00",X"00",X"00",X"99",X"BF",X"25",X"40",
		X"99",X"BF",X"40",X"1F",X"00",X"00",X"99",X"BF",X"25",X"40",X"99",X"BF",X"00",X"00",X"00",X"01",
		X"99",X"BF",X"20",X"45",X"99",X"BF",X"00",X"00",X"00",X"1F",X"99",X"BF",X"20",X"45",X"40",X"80",
		X"00",X"C0",X"87",X"60",X"40",X"80",X"40",X"80",X"00",X"C0",X"00",X"00",X"84",X"23",X"00",X"5F",
		X"00",X"00",X"7C",X"3C",X"00",X"C0",X"40",X"80",X"00",X"71",X"87",X"60",X"20",X"00",X"3E",X"1E",
		X"00",X"C0",X"04",X"4C",X"20",X"5B",X"04",X"5F",X"38",X"40",X"01",X"5F",X"26",X"40",X"FB",X"1F",
		X"00",X"20",X"3A",X"40",X"FB",X"1F",X"00",X"20",X"26",X"40",X"05",X"40",X"00",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
