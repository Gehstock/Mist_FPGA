library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_PGM is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_PGM is
	type rom is array(0 to  24575) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"F3",X"C3",X"69",X"00",X"FF",X"FF",X"FF",X"C3",X"3E",X"09",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C3",X"1F",X"0A",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"2B",X"0A",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C3",X"3E",X"0A",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C3",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"12",X"0F",X"AF",X"21",X"00",X"A8",X"06",X"08",X"77",
		X"23",X"10",X"FC",X"3E",X"9B",X"32",X"03",X"98",X"3A",X"02",X"98",X"E6",X"01",X"CA",X"3F",X"08",
		X"21",X"00",X"88",X"11",X"00",X"8C",X"FD",X"21",X"8D",X"00",X"C3",X"48",X"01",X"FD",X"21",X"94",
		X"00",X"C3",X"25",X"02",X"21",X"9A",X"00",X"C3",X"58",X"02",X"52",X"41",X"4D",X"20",X"31",X"47",
		X"48",X"4A",X"4B",X"00",X"21",X"00",X"80",X"11",X"00",X"88",X"FD",X"21",X"B1",X"00",X"C3",X"48",
		X"01",X"21",X"B7",X"00",X"C3",X"58",X"02",X"32",X"43",X"20",X"52",X"4F",X"4D",X"20",X"20",X"20",
		X"00",X"21",X"00",X"00",X"DD",X"21",X"CB",X"00",X"C3",X"30",X"01",X"21",X"D1",X"00",X"C3",X"58",
		X"02",X"32",X"45",X"00",X"21",X"00",X"10",X"DD",X"21",X"DE",X"00",X"C3",X"30",X"01",X"21",X"E4",
		X"00",X"C3",X"58",X"02",X"32",X"46",X"00",X"21",X"00",X"20",X"DD",X"21",X"F1",X"00",X"C3",X"30",
		X"01",X"21",X"F7",X"00",X"C3",X"58",X"02",X"32",X"48",X"00",X"21",X"00",X"30",X"DD",X"21",X"04",
		X"01",X"C3",X"30",X"01",X"21",X"0A",X"01",X"C3",X"58",X"02",X"32",X"4A",X"00",X"21",X"00",X"40",
		X"DD",X"21",X"17",X"01",X"C3",X"30",X"01",X"21",X"1D",X"01",X"C3",X"58",X"02",X"32",X"4C",X"00",
		X"21",X"26",X"01",X"C3",X"58",X"02",X"20",X"20",X"20",X"20",X"20",X"20",X"00",X"C3",X"B6",X"17",
		X"01",X"00",X"10",X"AF",X"86",X"23",X"0D",X"C2",X"34",X"01",X"08",X"3A",X"00",X"70",X"08",X"10",
		X"F3",X"FE",X"FF",X"C2",X"79",X"02",X"DD",X"E9",X"DD",X"21",X"4F",X"01",X"C3",X"8F",X"01",X"44",
		X"4D",X"36",X"00",X"23",X"7D",X"BB",X"C2",X"51",X"01",X"08",X"3A",X"00",X"B0",X"08",X"7C",X"BA",
		X"C2",X"51",X"01",X"69",X"60",X"01",X"55",X"00",X"DD",X"21",X"6F",X"01",X"C3",X"A0",X"01",X"01",
		X"AA",X"55",X"DD",X"21",X"79",X"01",X"C3",X"E2",X"01",X"01",X"FF",X"AA",X"DD",X"21",X"83",X"01",
		X"C3",X"A0",X"01",X"01",X"00",X"FF",X"DD",X"21",X"8D",X"01",X"C3",X"E2",X"01",X"FD",X"E9",X"06",
		X"00",X"70",X"7E",X"B8",X"C2",X"7F",X"02",X"08",X"3A",X"00",X"B0",X"08",X"10",X"F3",X"DD",X"E9",
		X"08",X"3A",X"00",X"B0",X"08",X"7C",X"D9",X"67",X"D9",X"7D",X"D9",X"6F",X"D9",X"7B",X"D9",X"5F",
		X"D9",X"7A",X"D9",X"57",X"D9",X"7E",X"A8",X"C2",X"7F",X"02",X"71",X"7E",X"A9",X"C2",X"7F",X"02",
		X"23",X"7D",X"BB",X"C2",X"B5",X"01",X"08",X"3A",X"00",X"B0",X"08",X"7C",X"BA",X"C2",X"B5",X"01",
		X"D9",X"7C",X"D9",X"67",X"D9",X"7D",X"D9",X"6F",X"D9",X"7B",X"D9",X"5F",X"D9",X"7A",X"D9",X"57",
		X"DD",X"E9",X"08",X"3A",X"00",X"B0",X"08",X"7C",X"D9",X"67",X"D9",X"7D",X"D9",X"6F",X"D9",X"7B",
		X"D9",X"5F",X"D9",X"7A",X"D9",X"57",X"D9",X"EB",X"2B",X"7E",X"A8",X"C2",X"7F",X"02",X"71",X"7E",
		X"A9",X"C2",X"7F",X"02",X"08",X"3A",X"00",X"B0",X"08",X"7D",X"BB",X"C2",X"F8",X"01",X"7C",X"BA",
		X"C2",X"F8",X"01",X"D9",X"7C",X"D9",X"67",X"D9",X"7D",X"D9",X"6F",X"D9",X"7B",X"D9",X"5F",X"D9",
		X"7A",X"D9",X"57",X"DD",X"E9",X"21",X"00",X"88",X"11",X"00",X"8C",X"06",X"10",X"DD",X"21",X"34",
		X"02",X"C3",X"45",X"02",X"21",X"00",X"90",X"11",X"00",X"94",X"06",X"00",X"DD",X"21",X"43",X"02",
		X"C3",X"45",X"02",X"FD",X"E9",X"70",X"23",X"7D",X"BB",X"C2",X"45",X"02",X"08",X"3A",X"00",X"B0",
		X"08",X"7C",X"BA",X"C2",X"45",X"02",X"DD",X"E9",X"EB",X"21",X"6E",X"8B",X"1A",X"B7",X"CA",X"76",
		X"02",X"D6",X"30",X"F2",X"68",X"02",X"3E",X"10",X"77",X"08",X"3A",X"00",X"B0",X"08",X"01",X"E0",
		X"FF",X"09",X"13",X"C3",X"5C",X"02",X"EB",X"23",X"E9",X"3A",X"00",X"B0",X"C3",X"79",X"02",X"3A",
		X"00",X"B0",X"C3",X"7F",X"02",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3A",X"9F",X"86",X"B7",X"C4",X"1F",X"4C",X"3A",X"8F",X"86",X"B7",X"28",X"16",X"3A",X"90",X"86",
		X"3C",X"3C",X"32",X"90",X"86",X"21",X"04",X"90",X"06",X"03",X"77",X"23",X"23",X"10",X"FB",X"AF",
		X"32",X"8F",X"86",X"3A",X"86",X"86",X"B7",X"CA",X"9B",X"04",X"FE",X"FF",X"28",X"0B",X"FE",X"FE",
		X"28",X"2F",X"FE",X"FD",X"28",X"40",X"C3",X"9B",X"04",X"AF",X"32",X"86",X"86",X"21",X"87",X"86",
		X"34",X"3A",X"87",X"86",X"21",X"07",X"90",X"06",X"07",X"CD",X"8B",X"04",X"21",X"35",X"90",X"06",
		X"01",X"CD",X"8B",X"04",X"3A",X"87",X"86",X"21",X"1B",X"90",X"06",X"07",X"CD",X"8B",X"04",X"18",
		X"3A",X"AF",X"32",X"86",X"86",X"21",X"87",X"86",X"34",X"3A",X"87",X"86",X"21",X"07",X"90",X"06",
		X"0C",X"CD",X"92",X"04",X"18",X"25",X"AF",X"32",X"86",X"86",X"21",X"87",X"86",X"34",X"3A",X"87",
		X"86",X"21",X"05",X"90",X"06",X"1C",X"CD",X"8B",X"04",X"18",X"10",X"77",X"23",X"23",X"3C",X"10",
		X"FA",X"C9",X"77",X"23",X"23",X"23",X"23",X"3C",X"10",X"F8",X"C9",X"3A",X"8C",X"86",X"CB",X"4F",
		X"C8",X"3A",X"3D",X"86",X"47",X"3A",X"3E",X"86",X"80",X"47",X"3A",X"3F",X"86",X"80",X"47",X"3A",
		X"40",X"86",X"80",X"B7",X"C8",X"F5",X"21",X"8D",X"86",X"34",X"CB",X"46",X"CA",X"CE",X"04",X"11",
		X"3C",X"80",X"01",X"00",X"80",X"21",X"8E",X"86",X"36",X"00",X"CB",X"FE",X"18",X"10",X"F1",X"3D",
		X"B7",X"C8",X"F5",X"11",X"3E",X"80",X"01",X"01",X"80",X"21",X"8E",X"86",X"CB",X"BE",X"0A",X"E6",
		X"1C",X"CA",X"FD",X"07",X"21",X"8E",X"86",X"34",X"FE",X"04",X"CA",X"FF",X"04",X"FE",X"08",X"CA",
		X"C7",X"05",X"FE",X"10",X"CA",X"91",X"06",X"FE",X"18",X"CA",X"47",X"07",X"C3",X"FD",X"07",X"D5",
		X"EB",X"5E",X"23",X"56",X"EB",X"D1",X"7E",X"FE",X"2E",X"38",X"18",X"FE",X"30",X"30",X"14",X"0A",
		X"E6",X"E3",X"02",X"D5",X"11",X"20",X"00",X"19",X"7E",X"FE",X"B0",X"38",X"25",X"36",X"10",X"D1",
		X"C3",X"FD",X"07",X"D5",X"11",X"20",X"00",X"19",X"D1",X"7E",X"FE",X"2E",X"38",X"18",X"FE",X"30",
		X"30",X"14",X"0A",X"E6",X"E3",X"02",X"D5",X"11",X"E0",X"FF",X"19",X"7E",X"FE",X"B0",X"38",X"02",
		X"36",X"10",X"D1",X"C3",X"FD",X"07",X"0A",X"3C",X"E6",X"03",X"FE",X"03",X"20",X"02",X"3E",X"00",
		X"67",X"0A",X"E6",X"FC",X"B4",X"02",X"E6",X"03",X"B7",X"C2",X"7F",X"05",X"D5",X"EB",X"5E",X"23",
		X"56",X"21",X"E0",X"FF",X"19",X"7E",X"FE",X"50",X"38",X"0E",X"FE",X"A0",X"30",X"0A",X"D1",X"0A",
		X"E6",X"E3",X"CB",X"E7",X"02",X"C3",X"E1",X"06",X"EB",X"E1",X"73",X"23",X"72",X"2B",X"EB",X"1A",
		X"6F",X"13",X"1A",X"67",X"0A",X"E6",X"03",X"C5",X"E5",X"26",X"00",X"6F",X"0A",X"E6",X"60",X"28",
		X"17",X"CB",X"6F",X"28",X"0E",X"CB",X"77",X"28",X"05",X"01",X"32",X"08",X"18",X"0D",X"01",X"0E",
		X"08",X"18",X"08",X"01",X"1A",X"08",X"18",X"03",X"01",X"26",X"08",X"09",X"7E",X"E1",X"77",X"C1",
		X"C5",X"F5",X"0A",X"E6",X"03",X"FE",X"02",X"C1",X"20",X"02",X"06",X"11",X"05",X"78",X"01",X"20",
		X"00",X"09",X"77",X"C1",X"C3",X"FE",X"07",X"D5",X"EB",X"5E",X"23",X"56",X"EB",X"D1",X"7E",X"FE",
		X"2E",X"38",X"18",X"FE",X"30",X"30",X"14",X"0A",X"E6",X"E3",X"02",X"D5",X"11",X"E0",X"FF",X"19",
		X"7E",X"FE",X"B0",X"38",X"25",X"36",X"10",X"D1",X"C3",X"FD",X"07",X"D5",X"11",X"E0",X"FF",X"19",
		X"D1",X"7E",X"FE",X"2E",X"38",X"18",X"FE",X"30",X"30",X"14",X"0A",X"E6",X"E3",X"02",X"D5",X"11",
		X"20",X"00",X"19",X"7E",X"FE",X"B0",X"38",X"02",X"36",X"10",X"D1",X"C3",X"FD",X"07",X"0A",X"3C",
		X"E6",X"03",X"FE",X"03",X"20",X"02",X"3E",X"00",X"67",X"0A",X"E6",X"FC",X"B4",X"02",X"E6",X"03",
		X"B7",X"C2",X"49",X"06",X"D5",X"EB",X"5E",X"23",X"56",X"21",X"20",X"00",X"19",X"7E",X"FE",X"50",
		X"38",X"10",X"FE",X"A0",X"30",X"0C",X"D1",X"0A",X"E6",X"E3",X"CB",X"DF",X"CB",X"E7",X"02",X"C3",
		X"97",X"07",X"EB",X"E1",X"73",X"23",X"72",X"2B",X"EB",X"1A",X"6F",X"13",X"1A",X"67",X"0A",X"E6",
		X"03",X"C5",X"E5",X"26",X"00",X"6F",X"0A",X"E6",X"60",X"28",X"17",X"CB",X"6F",X"28",X"0E",X"CB",
		X"77",X"28",X"05",X"01",X"35",X"08",X"18",X"0D",X"01",X"11",X"08",X"18",X"08",X"01",X"1D",X"08",
		X"18",X"03",X"01",X"29",X"08",X"09",X"7E",X"E1",X"77",X"C1",X"C5",X"F5",X"0A",X"E6",X"03",X"FE",
		X"02",X"C1",X"20",X"02",X"06",X"0F",X"04",X"78",X"01",X"E0",X"FF",X"09",X"77",X"C1",X"C3",X"FE",
		X"07",X"D5",X"EB",X"5E",X"23",X"56",X"EB",X"D1",X"7E",X"FE",X"2E",X"38",X"14",X"FE",X"30",X"30",
		X"10",X"0A",X"E6",X"E3",X"02",X"2B",X"7E",X"FE",X"B0",X"DA",X"FD",X"07",X"36",X"10",X"C3",X"FD",
		X"07",X"2B",X"7E",X"FE",X"2E",X"38",X"14",X"FE",X"30",X"30",X"10",X"0A",X"E6",X"E3",X"02",X"23",
		X"7E",X"FE",X"B0",X"DA",X"FD",X"07",X"36",X"10",X"C3",X"FD",X"07",X"0A",X"3C",X"E6",X"03",X"FE",
		X"03",X"20",X"02",X"3E",X"00",X"67",X"0A",X"E6",X"FC",X"B4",X"02",X"E6",X"03",X"B7",X"C2",X"02",
		X"07",X"D5",X"EB",X"5E",X"23",X"56",X"13",X"EB",X"7E",X"FE",X"50",X"38",X"0E",X"FE",X"A0",X"30",
		X"0A",X"D1",X"0A",X"E6",X"E3",X"CB",X"DF",X"02",X"C3",X"24",X"06",X"EB",X"E1",X"73",X"23",X"72",
		X"2B",X"EB",X"1A",X"6F",X"13",X"1A",X"67",X"0A",X"E6",X"03",X"C5",X"E5",X"26",X"00",X"6F",X"0A",
		X"E6",X"60",X"28",X"17",X"CB",X"6F",X"28",X"0E",X"CB",X"77",X"28",X"05",X"01",X"38",X"08",X"18",
		X"0D",X"01",X"14",X"08",X"18",X"08",X"01",X"20",X"08",X"18",X"03",X"01",X"2C",X"08",X"09",X"7E",
		X"E1",X"77",X"C1",X"C5",X"F5",X"0A",X"E6",X"03",X"FE",X"02",X"C1",X"20",X"02",X"06",X"11",X"05",
		X"78",X"2B",X"77",X"C1",X"C3",X"FE",X"07",X"D5",X"EB",X"5E",X"23",X"56",X"EB",X"D1",X"7E",X"FE",
		X"2E",X"38",X"14",X"FE",X"30",X"30",X"10",X"0A",X"E6",X"E3",X"02",X"23",X"7E",X"FE",X"B0",X"DA",
		X"FD",X"07",X"36",X"10",X"C3",X"FD",X"07",X"23",X"7E",X"FE",X"2E",X"38",X"14",X"FE",X"30",X"30",
		X"10",X"0A",X"E6",X"E3",X"02",X"2B",X"7E",X"FE",X"B0",X"DA",X"FD",X"07",X"36",X"10",X"C3",X"FD",
		X"07",X"0A",X"3C",X"E6",X"03",X"FE",X"03",X"20",X"02",X"3E",X"00",X"67",X"0A",X"E6",X"FC",X"B4",
		X"02",X"E6",X"03",X"B7",X"C2",X"B8",X"07",X"D5",X"EB",X"5E",X"23",X"56",X"1B",X"EB",X"7E",X"FE",
		X"50",X"38",X"0E",X"FE",X"A0",X"30",X"0A",X"D1",X"0A",X"E6",X"E3",X"CB",X"D7",X"02",X"C3",X"5C",
		X"05",X"EB",X"E1",X"73",X"23",X"72",X"2B",X"EB",X"1A",X"6F",X"13",X"1A",X"67",X"0A",X"E6",X"03",
		X"C5",X"E5",X"26",X"00",X"6F",X"0A",X"E6",X"60",X"28",X"17",X"CB",X"6F",X"28",X"0E",X"CB",X"77",
		X"28",X"05",X"01",X"3B",X"08",X"18",X"0D",X"01",X"17",X"08",X"18",X"08",X"01",X"23",X"08",X"18",
		X"03",X"01",X"2F",X"08",X"09",X"7E",X"E1",X"77",X"C1",X"C5",X"F5",X"0A",X"E6",X"03",X"FE",X"02",
		X"C1",X"20",X"02",X"06",X"0F",X"04",X"78",X"23",X"77",X"C1",X"C3",X"FE",X"07",X"13",X"F1",X"3D",
		X"B7",X"C8",X"3D",X"B7",X"C8",X"F5",X"13",X"13",X"13",X"03",X"03",X"C3",X"DE",X"04",X"FE",X"FC",
		X"FF",X"F8",X"F6",X"FA",X"F4",X"F2",X"F5",X"EE",X"EC",X"F0",X"EA",X"E8",X"EB",X"E4",X"E2",X"E6",
		X"E0",X"DE",X"E1",X"DA",X"D8",X"DC",X"D6",X"D4",X"D7",X"D0",X"CE",X"D2",X"CC",X"CA",X"CD",X"C6",
		X"C4",X"C7",X"C2",X"C0",X"C3",X"BC",X"BA",X"BE",X"B8",X"B6",X"B9",X"B2",X"B0",X"B4",X"DC",X"31",
		X"80",X"80",X"F5",X"3A",X"00",X"B0",X"F1",X"CD",X"C1",X"09",X"F5",X"3A",X"00",X"B0",X"F1",X"D7",
		X"00",X"E7",X"04",X"04",X"01",X"E7",X"04",X"08",X"02",X"E7",X"04",X"0C",X"03",X"E7",X"04",X"10",
		X"04",X"3E",X"9B",X"32",X"03",X"98",X"3E",X"88",X"32",X"03",X"A0",X"F5",X"3A",X"00",X"B0",X"F1",
		X"3E",X"10",X"32",X"02",X"98",X"3E",X"00",X"32",X"02",X"98",X"CF",X"68",X"40",X"50",X"4F",X"52",
		X"54",X"20",X"41",X"00",X"21",X"50",X"40",X"CD",X"FE",X"08",X"3A",X"00",X"98",X"CD",X"E6",X"08",
		X"CF",X"68",X"60",X"50",X"4F",X"52",X"54",X"20",X"42",X"00",X"21",X"70",X"40",X"CD",X"FE",X"08",
		X"3A",X"01",X"98",X"CD",X"E6",X"08",X"CF",X"68",X"80",X"50",X"4F",X"52",X"54",X"20",X"43",X"00",
		X"21",X"90",X"40",X"CD",X"FE",X"08",X"3A",X"02",X"98",X"CD",X"E6",X"08",X"CF",X"40",X"A8",X"37",
		X"20",X"36",X"20",X"35",X"20",X"34",X"20",X"33",X"20",X"32",X"20",X"31",X"20",X"30",X"00",X"CF",
		X"50",X"B0",X"42",X"49",X"54",X"20",X"4E",X"55",X"4D",X"42",X"45",X"52",X"53",X"00",X"2E",X"00",
		X"2D",X"20",X"FD",X"C3",X"6B",X"08",X"06",X"08",X"07",X"F5",X"E6",X"01",X"F6",X"30",X"CD",X"A9",
		X"09",X"AF",X"CD",X"A9",X"09",X"F5",X"3A",X"00",X"B0",X"F1",X"F1",X"10",X"EB",X"C9",X"F5",X"AF",
		X"C3",X"03",X"09",X"94",X"3D",X"67",X"CB",X"3C",X"CB",X"3C",X"CB",X"3C",X"CB",X"3C",X"CB",X"1D",
		X"CB",X"3C",X"CB",X"1D",X"CB",X"3C",X"CB",X"1D",X"D5",X"11",X"00",X"88",X"19",X"D1",X"F1",X"C9",
		X"D5",X"11",X"00",X"88",X"B7",X"ED",X"52",X"CB",X"25",X"CB",X"14",X"CB",X"25",X"CB",X"14",X"CB",
		X"25",X"CB",X"14",X"7C",X"2F",X"67",X"CB",X"24",X"CB",X"24",X"CB",X"24",X"D1",X"C9",X"E3",X"F5",
		X"C5",X"D5",X"56",X"23",X"5E",X"23",X"EB",X"CD",X"FE",X"08",X"1A",X"13",X"B7",X"CA",X"56",X"09",
		X"CD",X"A9",X"09",X"C3",X"4A",X"09",X"EB",X"D1",X"C1",X"F1",X"E3",X"C9",X"0E",X"03",X"C3",X"68",
		X"09",X"0E",X"00",X"C3",X"68",X"09",X"0E",X"01",X"F5",X"C5",X"D5",X"E5",X"CD",X"FE",X"08",X"78",
		X"3D",X"20",X"02",X"CB",X"81",X"1A",X"CB",X"40",X"20",X"05",X"07",X"07",X"07",X"07",X"1B",X"13",
		X"E6",X"0F",X"C2",X"94",X"09",X"CB",X"41",X"CA",X"96",X"09",X"3E",X"20",X"CB",X"49",X"C2",X"A2",
		X"09",X"C3",X"9F",X"09",X"CB",X"81",X"C6",X"30",X"FE",X"3A",X"DA",X"9F",X"09",X"C6",X"07",X"CD",
		X"A9",X"09",X"10",X"CB",X"E1",X"D1",X"C1",X"F1",X"C9",X"C5",X"D6",X"30",X"F2",X"B1",X"09",X"3E",
		X"10",X"77",X"01",X"E0",X"FF",X"09",X"7C",X"FE",X"88",X"30",X"04",X"01",X"00",X"04",X"09",X"C1",
		X"C9",X"F5",X"C5",X"E5",X"D5",X"3E",X"00",X"32",X"86",X"86",X"06",X"14",X"21",X"6B",X"86",X"36",
		X"00",X"23",X"10",X"FB",X"21",X"00",X"88",X"0E",X"04",X"3E",X"10",X"CD",X"F7",X"09",X"21",X"00",
		X"90",X"0E",X"01",X"CD",X"F6",X"09",X"3E",X"00",X"32",X"03",X"A8",X"32",X"05",X"A8",X"32",X"04",
		X"A8",X"D1",X"E1",X"C1",X"F1",X"C9",X"AF",X"06",X"00",X"77",X"23",X"10",X"FC",X"0D",X"20",X"F9",
		X"C9",X"F5",X"C5",X"D5",X"E5",X"50",X"E5",X"CD",X"FE",X"08",X"3E",X"20",X"CD",X"A9",X"09",X"10",
		X"F9",X"E1",X"7D",X"C6",X"08",X"6F",X"42",X"0D",X"20",X"EC",X"E1",X"D1",X"C1",X"F1",X"C9",X"E1",
		X"7E",X"23",X"E5",X"11",X"00",X"00",X"06",X"20",X"C3",X"48",X"0A",X"E1",X"7E",X"23",X"E5",X"47",
		X"0F",X"0F",X"E6",X"3E",X"4F",X"78",X"06",X"00",X"21",X"01",X"90",X"09",X"77",X"C9",X"E1",X"46",
		X"23",X"5E",X"16",X"00",X"23",X"7E",X"23",X"E5",X"21",X"01",X"90",X"19",X"19",X"77",X"23",X"23",
		X"10",X"FB",X"C9",X"21",X"01",X"90",X"19",X"19",X"77",X"23",X"23",X"10",X"FB",X"C9",X"77",X"3C",
		X"23",X"77",X"3C",X"11",X"1F",X"00",X"19",X"77",X"3C",X"23",X"77",X"C9",X"DF",X"FC",X"CF",X"10",
		X"F8",X"3B",X"31",X"39",X"38",X"32",X"20",X"20",X"54",X"41",X"47",X"4F",X"20",X"45",X"4C",X"45",
		X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",X"43",X"00",X"C9",X"AF",X"32",
		X"65",X"86",X"3A",X"CA",X"81",X"B7",X"28",X"1E",X"DF",X"F2",X"CF",X"80",X"E8",X"20",X"43",X"52",
		X"45",X"44",X"49",X"54",X"53",X"5B",X"20",X"20",X"20",X"00",X"21",X"E8",X"C8",X"11",X"CA",X"81",
		X"06",X"02",X"CD",X"66",X"09",X"C9",X"DF",X"F6",X"CF",X"80",X"E8",X"49",X"4E",X"53",X"45",X"52",
		X"54",X"20",X"43",X"4F",X"49",X"4E",X"00",X"C9",X"3A",X"66",X"86",X"B7",X"C0",X"AF",X"32",X"64",
		X"86",X"DF",X"0B",X"CF",X"10",X"00",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"31",X"00",X"21",
		X"08",X"10",X"11",X"07",X"82",X"06",X"06",X"CD",X"66",X"09",X"CF",X"70",X"00",X"48",X"49",X"47",
		X"48",X"00",X"21",X"08",X"68",X"11",X"CB",X"81",X"06",X"06",X"CD",X"66",X"09",X"3A",X"67",X"86",
		X"FE",X"02",X"C0",X"CF",X"B0",X"00",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"32",X"00",X"21",
		X"08",X"C0",X"11",X"0A",X"82",X"06",X"06",X"CD",X"66",X"09",X"C9",X"DF",X"F9",X"CF",X"10",X"18",
		X"20",X"20",X"20",X"20",X"20",X"20",X"00",X"CF",X"C0",X"18",X"20",X"20",X"20",X"20",X"20",X"20",
		X"00",X"3A",X"33",X"86",X"B7",X"28",X"0F",X"3D",X"28",X"0C",X"FE",X"05",X"38",X"02",X"3E",X"05",
		X"21",X"18",X"18",X"CD",X"56",X"0B",X"3A",X"47",X"86",X"B7",X"C8",X"3D",X"C8",X"FE",X"05",X"38",
		X"02",X"3E",X"05",X"21",X"18",X"C8",X"E5",X"CD",X"FE",X"08",X"36",X"2C",X"E1",X"3D",X"C8",X"08",
		X"7C",X"C6",X"08",X"67",X"08",X"18",X"EF",X"C9",X"3A",X"CA",X"81",X"B7",X"C8",X"21",X"A8",X"00",
		X"01",X"05",X"20",X"CD",X"01",X"0A",X"E7",X"07",X"15",X"05",X"3A",X"CA",X"81",X"FE",X"01",X"20",
		X"41",X"CF",X"18",X"A8",X"50",X"55",X"53",X"48",X"20",X"31",X"20",X"50",X"4C",X"41",X"59",X"45",
		X"52",X"20",X"53",X"54",X"41",X"52",X"54",X"20",X"42",X"55",X"54",X"54",X"4F",X"4E",X"00",X"CF",
		X"68",X"B8",X"5B",X"20",X"4F",X"52",X"20",X"5B",X"00",X"CF",X"30",X"C8",X"49",X"4E",X"53",X"45",
		X"52",X"54",X"20",X"41",X"4E",X"4F",X"54",X"48",X"45",X"52",X"20",X"43",X"4F",X"49",X"4E",X"00",
		X"18",X"34",X"CF",X"48",X"A8",X"50",X"55",X"53",X"48",X"20",X"31",X"20",X"50",X"4C",X"41",X"59",
		X"45",X"52",X"00",X"CF",X"68",X"B8",X"5B",X"20",X"4F",X"52",X"20",X"5B",X"00",X"CF",X"28",X"C8",
		X"32",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"53",X"54",X"41",X"52",X"54",X"20",X"42",
		X"55",X"54",X"54",X"4F",X"4E",X"00",X"06",X"05",X"C5",X"E7",X"07",X"15",X"01",X"3E",X"02",X"CD",
		X"7B",X"18",X"E7",X"07",X"15",X"02",X"3E",X"02",X"CD",X"7B",X"18",X"E7",X"07",X"15",X"03",X"3E",
		X"02",X"CD",X"7B",X"18",X"E7",X"07",X"15",X"04",X"3E",X"02",X"CD",X"7B",X"18",X"E7",X"07",X"15",
		X"05",X"3E",X"02",X"CD",X"7B",X"18",X"E7",X"07",X"15",X"06",X"3E",X"02",X"CD",X"7B",X"18",X"E7",
		X"07",X"15",X"07",X"3E",X"02",X"CD",X"7B",X"18",X"E7",X"07",X"15",X"00",X"3E",X"02",X"CD",X"7B",
		X"18",X"C1",X"10",X"B4",X"C9",X"F5",X"3A",X"66",X"86",X"B7",X"28",X"09",X"3A",X"01",X"98",X"E6",
		X"02",X"28",X"02",X"F1",X"C9",X"F1",X"F3",X"32",X"00",X"A0",X"AF",X"32",X"01",X"A0",X"E3",X"E3",
		X"3E",X"08",X"32",X"01",X"A0",X"FB",X"C9",X"D5",X"E5",X"ED",X"5B",X"5F",X"86",X"21",X"AA",X"AA",
		X"19",X"29",X"19",X"29",X"19",X"29",X"19",X"29",X"29",X"19",X"29",X"29",X"19",X"29",X"29",X"19",
		X"29",X"19",X"29",X"29",X"19",X"29",X"19",X"29",X"19",X"11",X"2F",X"6A",X"19",X"22",X"5F",X"86",
		X"7C",X"E1",X"D1",X"C9",X"FD",X"E1",X"DD",X"21",X"4A",X"83",X"DD",X"CB",X"00",X"C6",X"DD",X"CB",
		X"00",X"CE",X"CD",X"B2",X"0D",X"31",X"44",X"81",X"FD",X"E9",X"FD",X"E1",X"DD",X"21",X"EE",X"82",
		X"DD",X"CB",X"00",X"C6",X"DD",X"CB",X"00",X"CE",X"CD",X"B2",X"0D",X"31",X"6C",X"81",X"DD",X"21",
		X"67",X"82",X"DD",X"CB",X"00",X"C6",X"CD",X"9B",X"0D",X"CD",X"C6",X"0D",X"FD",X"E9",X"FD",X"E1",
		X"DD",X"21",X"1C",X"83",X"DD",X"CB",X"00",X"C6",X"DD",X"CB",X"00",X"CE",X"CD",X"B2",X"0D",X"31",
		X"94",X"81",X"DD",X"21",X"76",X"82",X"DD",X"CB",X"00",X"C6",X"CD",X"9B",X"0D",X"CD",X"C6",X"0D",
		X"FD",X"E9",X"D9",X"21",X"E2",X"0E",X"CD",X"80",X"0D",X"D9",X"D0",X"CD",X"9B",X"0D",X"CD",X"C6",
		X"0D",X"37",X"C9",X"D9",X"21",X"F0",X"0E",X"CD",X"80",X"0D",X"D9",X"D0",X"CD",X"9B",X"0D",X"CD",
		X"C6",X"0D",X"37",X"C9",X"FD",X"E1",X"CD",X"68",X"0D",X"30",X"14",X"DD",X"CB",X"00",X"C6",X"DD",
		X"CB",X"00",X"CE",X"CD",X"B2",X"0D",X"CD",X"5B",X"0E",X"CD",X"03",X"0D",X"37",X"FD",X"E9",X"C3",
		X"12",X"0E",X"FD",X"E1",X"CD",X"70",X"0D",X"30",X"F6",X"DD",X"CB",X"00",X"C6",X"DD",X"CB",X"00",
		X"CE",X"CD",X"B2",X"0D",X"CD",X"5B",X"0E",X"CD",X"03",X"0D",X"37",X"FD",X"E9",X"C3",X"12",X"0E",
		X"E1",X"D9",X"21",X"00",X"0F",X"CD",X"80",X"0D",X"D9",X"D2",X"67",X"0D",X"DD",X"22",X"B6",X"81",
		X"CD",X"B2",X"0D",X"CD",X"5B",X"0E",X"37",X"E9",X"E1",X"D9",X"21",X"D0",X"0E",X"C3",X"55",X"0D",
		X"E1",X"D9",X"21",X"D0",X"0E",X"C3",X"55",X"0D",X"E1",X"D9",X"21",X"E0",X"0E",X"C3",X"55",X"0D",
		X"E5",X"D1",X"7E",X"23",X"66",X"6F",X"B4",X"C8",X"7E",X"B7",X"28",X"06",X"13",X"13",X"D5",X"E1",
		X"18",X"F0",X"E5",X"DD",X"E1",X"DD",X"CB",X"00",X"C6",X"37",X"C9",X"D9",X"DD",X"E5",X"E1",X"DD",
		X"2A",X"B6",X"81",X"DD",X"75",X"01",X"DD",X"74",X"02",X"DD",X"CB",X"00",X"DE",X"E5",X"DD",X"E1",
		X"D9",X"C9",X"D9",X"DD",X"CB",X"00",X"CE",X"DD",X"E5",X"E1",X"22",X"B6",X"81",X"AF",X"06",X"0F",
		X"23",X"77",X"10",X"FC",X"D9",X"C9",X"D9",X"DD",X"E5",X"E1",X"22",X"B4",X"81",X"AF",X"06",X"0E",
		X"23",X"77",X"10",X"FC",X"D9",X"C9",X"21",X"00",X"00",X"39",X"31",X"1C",X"81",X"FD",X"E5",X"FD",
		X"2A",X"B6",X"81",X"FD",X"22",X"BA",X"81",X"FD",X"75",X"0E",X"FD",X"74",X"0F",X"C9",X"21",X"00",
		X"00",X"39",X"31",X"1C",X"81",X"DD",X"2A",X"B6",X"81",X"DD",X"75",X"0E",X"DD",X"74",X"0F",X"2A",
		X"BA",X"81",X"7C",X"B5",X"28",X"0C",X"DD",X"2A",X"BA",X"81",X"21",X"00",X"00",X"22",X"BA",X"81",
		X"18",X"04",X"DD",X"2A",X"B6",X"81",X"CD",X"2B",X"0E",X"DD",X"CB",X"00",X"46",X"28",X"F7",X"DD",
		X"22",X"B6",X"81",X"DD",X"66",X"0F",X"DD",X"6E",X"0E",X"F9",X"C9",X"D9",X"01",X"2E",X"00",X"DD",
		X"09",X"DD",X"E5",X"E1",X"01",X"2A",X"86",X"B7",X"ED",X"42",X"38",X"04",X"DD",X"21",X"EE",X"82",
		X"D9",X"C9",X"DD",X"2A",X"B6",X"81",X"DD",X"77",X"03",X"DD",X"CB",X"00",X"EE",X"CD",X"EE",X"0D",
		X"DD",X"2A",X"B6",X"81",X"DD",X"CB",X"00",X"6E",X"20",X"F3",X"C9",X"D9",X"D1",X"01",X"2E",X"00",
		X"DD",X"E5",X"E1",X"09",X"F9",X"D5",X"D9",X"C9",X"CD",X"78",X"0E",X"D9",X"2A",X"B6",X"81",X"06",
		X"10",X"AF",X"77",X"23",X"10",X"FC",X"D9",X"C9",X"DD",X"2A",X"B6",X"81",X"DD",X"CB",X"00",X"5E",
		X"C8",X"DD",X"CB",X"00",X"9E",X"D9",X"DD",X"6E",X"01",X"DD",X"66",X"02",X"06",X"0F",X"AF",X"77",
		X"23",X"10",X"FC",X"DD",X"77",X"01",X"DD",X"77",X"01",X"D9",X"C9",X"CD",X"00",X"10",X"DD",X"21",
		X"EE",X"82",X"AF",X"DD",X"77",X"00",X"DD",X"21",X"1C",X"83",X"AF",X"DD",X"77",X"00",X"DD",X"21",
		X"78",X"83",X"DD",X"77",X"00",X"CD",X"2B",X"0E",X"30",X"02",X"18",X"F6",X"DD",X"21",X"0D",X"82",
		X"11",X"0F",X"00",X"06",X"0F",X"DD",X"77",X"00",X"DD",X"19",X"10",X"F9",X"CD",X"06",X"10",X"C9",
		X"E8",X"84",X"16",X"85",X"44",X"85",X"00",X"00",X"72",X"85",X"A0",X"85",X"CE",X"85",X"00",X"00",
		X"00",X"00",X"0D",X"82",X"1C",X"82",X"2B",X"82",X"3A",X"82",X"49",X"82",X"58",X"82",X"00",X"00",
		X"85",X"82",X"94",X"82",X"A3",X"82",X"B2",X"82",X"C1",X"82",X"D0",X"82",X"DF",X"82",X"00",X"00",
		X"78",X"83",X"A6",X"83",X"D4",X"83",X"02",X"84",X"30",X"84",X"5E",X"84",X"8C",X"84",X"BA",X"84",
		X"00",X"00",X"F5",X"3A",X"00",X"B0",X"AF",X"32",X"01",X"A8",X"3C",X"32",X"01",X"A8",X"3A",X"BE",
		X"81",X"CB",X"0F",X"32",X"BE",X"81",X"DA",X"DA",X"0F",X"3A",X"BF",X"81",X"B7",X"C2",X"D8",X"0F",
		X"3C",X"32",X"BF",X"81",X"ED",X"73",X"B8",X"81",X"31",X"F4",X"80",X"08",X"F5",X"C5",X"D5",X"E5",
		X"DD",X"E5",X"FD",X"E5",X"D9",X"C5",X"D5",X"E5",X"21",X"0D",X"82",X"11",X"40",X"90",X"06",X"08",
		X"C5",X"CB",X"46",X"CC",X"C9",X"11",X"01",X"06",X"00",X"09",X"7E",X"12",X"23",X"13",X"7E",X"12",
		X"23",X"13",X"7E",X"12",X"23",X"23",X"23",X"23",X"13",X"7E",X"12",X"23",X"23",X"23",X"13",X"C1",
		X"10",X"DE",X"21",X"85",X"82",X"11",X"61",X"90",X"06",X"07",X"C5",X"E5",X"DD",X"E1",X"01",X"06",
		X"00",X"09",X"7E",X"C6",X"08",X"12",X"01",X"06",X"00",X"09",X"13",X"13",X"7E",X"2F",X"C6",X"F1",
		X"12",X"13",X"13",X"23",X"23",X"23",X"C1",X"10",X"E1",X"CD",X"00",X"04",X"CD",X"48",X"14",X"21",
		X"EE",X"82",X"06",X"11",X"C5",X"46",X"CB",X"40",X"C4",X"0C",X"10",X"CB",X"58",X"C4",X"5B",X"10",
		X"11",X"2E",X"00",X"19",X"C1",X"10",X"ED",X"CD",X"1A",X"11",X"CD",X"96",X"11",X"CD",X"E8",X"11",
		X"CD",X"EE",X"12",X"E1",X"D1",X"C1",X"D9",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"F1",X"08",
		X"ED",X"7B",X"B8",X"81",X"AF",X"32",X"BF",X"81",X"F1",X"C9",X"ED",X"73",X"BC",X"81",X"31",X"B4",
		X"81",X"C5",X"D5",X"E5",X"DD",X"E5",X"08",X"D9",X"F5",X"C5",X"D5",X"E5",X"CD",X"EE",X"12",X"E1",
		X"D1",X"C1",X"F1",X"D9",X"08",X"DD",X"E1",X"E1",X"D1",X"C1",X"ED",X"7B",X"BC",X"81",X"F1",X"C9",
		X"3E",X"FF",X"32",X"BE",X"81",X"C9",X"3E",X"55",X"32",X"BE",X"81",X"C9",X"E5",X"CB",X"48",X"CA",
		X"58",X"10",X"23",X"5E",X"23",X"56",X"D5",X"FD",X"E1",X"23",X"CB",X"68",X"28",X"05",X"35",X"20",
		X"02",X"CB",X"A8",X"23",X"CB",X"60",X"28",X"2C",X"35",X"20",X"29",X"CB",X"F8",X"23",X"5E",X"23",
		X"56",X"13",X"13",X"13",X"13",X"13",X"1A",X"B7",X"C2",X"4C",X"10",X"13",X"1A",X"B7",X"C2",X"45",
		X"10",X"CB",X"A0",X"CB",X"B8",X"EB",X"23",X"7E",X"23",X"66",X"6F",X"EB",X"72",X"2B",X"73",X"13",
		X"13",X"1A",X"2B",X"77",X"CB",X"50",X"28",X"00",X"E1",X"70",X"C9",X"CB",X"48",X"C8",X"E5",X"DD",
		X"E1",X"E5",X"FD",X"CB",X"00",X"66",X"28",X"17",X"DD",X"7E",X"08",X"C6",X"08",X"67",X"DD",X"7E",
		X"0A",X"C6",X"08",X"6F",X"CD",X"FE",X"08",X"FD",X"7E",X"0E",X"77",X"FD",X"CB",X"00",X"A6",X"E1",
		X"CB",X"78",X"28",X"14",X"CB",X"BE",X"DD",X"66",X"06",X"DD",X"6E",X"05",X"23",X"23",X"23",X"7E",
		X"FD",X"77",X"07",X"23",X"7E",X"FD",X"77",X"08",X"FD",X"CB",X"00",X"4E",X"28",X"09",X"FD",X"35",
		X"01",X"20",X"04",X"FD",X"CB",X"00",X"8E",X"FD",X"CB",X"00",X"56",X"28",X"09",X"FD",X"35",X"02",
		X"20",X"04",X"FD",X"CB",X"00",X"96",X"CB",X"50",X"28",X"49",X"DD",X"7E",X"07",X"FD",X"77",X"05",
		X"DD",X"7E",X"08",X"FD",X"77",X"06",X"DD",X"7E",X"09",X"FD",X"77",X"0B",X"DD",X"7E",X"0A",X"FD",
		X"77",X"0C",X"FD",X"E5",X"E1",X"23",X"23",X"23",X"5E",X"23",X"56",X"23",X"4E",X"23",X"46",X"EB",
		X"09",X"EB",X"DD",X"72",X"08",X"DD",X"73",X"07",X"2B",X"73",X"23",X"72",X"23",X"23",X"23",X"5E",
		X"23",X"56",X"23",X"4E",X"23",X"46",X"EB",X"09",X"EB",X"DD",X"72",X"0A",X"DD",X"73",X"09",X"2B",
		X"73",X"23",X"72",X"DD",X"7E",X"08",X"C6",X"08",X"67",X"DD",X"7E",X"0A",X"C6",X"08",X"6F",X"CD",
		X"FE",X"08",X"7E",X"FD",X"77",X"0D",X"DD",X"E5",X"E1",X"C9",X"DD",X"21",X"E8",X"84",X"06",X"07",
		X"DD",X"CB",X"00",X"46",X"C4",X"2F",X"11",X"11",X"2E",X"00",X"DD",X"19",X"10",X"F2",X"C9",X"DD",
		X"7E",X"0D",X"FE",X"FF",X"C8",X"DD",X"66",X"02",X"DD",X"6E",X"01",X"E5",X"FD",X"E1",X"FD",X"7E",
		X"0D",X"D9",X"FE",X"50",X"38",X"4E",X"DD",X"36",X"0D",X"FF",X"FE",X"A0",X"38",X"46",X"01",X"01",
		X"02",X"DD",X"CB",X"0C",X"76",X"28",X"05",X"CD",X"8B",X"1B",X"18",X"03",X"CD",X"03",X"1C",X"DD",
		X"7E",X"08",X"C6",X"08",X"67",X"DD",X"7E",X"0A",X"C6",X"08",X"6F",X"CD",X"FE",X"08",X"36",X"2E",
		X"EB",X"21",X"6B",X"86",X"CD",X"67",X"0C",X"E6",X"03",X"20",X"01",X"3C",X"CD",X"45",X"0C",X"06",
		X"09",X"4E",X"23",X"7E",X"23",X"B1",X"20",X"07",X"2B",X"2B",X"73",X"23",X"72",X"18",X"05",X"10",
		X"F0",X"EB",X"36",X"10",X"D9",X"C9",X"21",X"6A",X"86",X"35",X"7E",X"B7",X"C0",X"36",X"05",X"21",
		X"6B",X"86",X"06",X"0A",X"5E",X"23",X"56",X"23",X"7A",X"B3",X"28",X"1A",X"1A",X"FE",X"2E",X"38",
		X"0A",X"FE",X"37",X"28",X"06",X"30",X"04",X"3C",X"12",X"18",X"0B",X"3E",X"10",X"12",X"2B",X"2B",
		X"36",X"00",X"23",X"36",X"00",X"23",X"10",X"DC",X"C9",X"AF",X"E5",X"DD",X"E1",X"DD",X"77",X"06",
		X"DD",X"77",X"0C",X"C9",X"7A",X"2F",X"57",X"7B",X"2F",X"5F",X"13",X"C9",X"78",X"2F",X"47",X"79",
		X"2F",X"4F",X"03",X"C9",X"00",X"00",X"00",X"00",X"DD",X"21",X"EE",X"82",X"FD",X"21",X"78",X"83",
		X"3E",X"08",X"6F",X"DD",X"4E",X"0A",X"CD",X"0B",X"12",X"DD",X"21",X"1C",X"83",X"FD",X"21",X"78",
		X"83",X"3E",X"08",X"6F",X"DD",X"4E",X"0A",X"CD",X"0B",X"12",X"C9",X"D9",X"3E",X"08",X"6F",X"DD",
		X"4E",X"08",X"06",X"08",X"FD",X"7E",X"00",X"E6",X"41",X"EE",X"41",X"20",X"3B",X"FD",X"56",X"06",
		X"FD",X"5E",X"05",X"1A",X"67",X"13",X"1A",X"D9",X"85",X"1F",X"67",X"FD",X"7E",X"0A",X"91",X"30",
		X"02",X"ED",X"44",X"BC",X"D9",X"30",X"21",X"7C",X"85",X"1F",X"67",X"FD",X"7E",X"08",X"91",X"30",
		X"02",X"ED",X"44",X"BC",X"30",X"12",X"DD",X"7E",X"0D",X"FD",X"B6",X"0C",X"DD",X"77",X"0D",X"FD",
		X"7E",X"0D",X"DD",X"B6",X"0C",X"FD",X"77",X"0D",X"11",X"2E",X"00",X"FD",X"19",X"10",X"B5",X"DD",
		X"21",X"E8",X"84",X"CD",X"86",X"12",X"DD",X"21",X"16",X"85",X"CD",X"86",X"12",X"DD",X"21",X"44",
		X"85",X"CD",X"86",X"12",X"DD",X"21",X"72",X"85",X"CD",X"86",X"12",X"DD",X"21",X"A0",X"85",X"CD",
		X"86",X"12",X"DD",X"21",X"CE",X"85",X"DD",X"7E",X"00",X"E6",X"41",X"EE",X"41",X"C0",X"FD",X"21",
		X"EE",X"82",X"3E",X"02",X"6F",X"DD",X"4E",X"0A",X"D9",X"3E",X"02",X"6F",X"DD",X"4E",X"08",X"06",
		X"0B",X"FD",X"7E",X"00",X"E6",X"41",X"EE",X"41",X"20",X"3B",X"FD",X"56",X"06",X"FD",X"5E",X"05",
		X"1A",X"67",X"13",X"1A",X"D9",X"85",X"1F",X"67",X"FD",X"7E",X"0A",X"91",X"30",X"02",X"ED",X"44",
		X"BC",X"D9",X"30",X"21",X"7C",X"85",X"1F",X"67",X"FD",X"7E",X"08",X"91",X"30",X"02",X"ED",X"44",
		X"BC",X"30",X"12",X"DD",X"7E",X"0D",X"FD",X"B6",X"0C",X"DD",X"77",X"0D",X"FD",X"7E",X"0D",X"DD",
		X"B6",X"0C",X"FD",X"77",X"0D",X"11",X"2E",X"00",X"FD",X"19",X"10",X"B5",X"D9",X"C9",X"21",X"C0",
		X"81",X"7E",X"23",X"46",X"A8",X"4F",X"3A",X"00",X"98",X"2F",X"77",X"2B",X"70",X"A1",X"E6",X"C0",
		X"23",X"23",X"CB",X"7F",X"28",X"01",X"34",X"23",X"CB",X"77",X"28",X"01",X"34",X"CD",X"3B",X"13",
		X"CD",X"A2",X"13",X"C9",X"3A",X"CA",X"81",X"C6",X"99",X"27",X"32",X"CA",X"81",X"C9",X"47",X"B7",
		X"C8",X"3E",X"FF",X"32",X"65",X"86",X"3A",X"CA",X"81",X"FE",X"99",X"C8",X"80",X"27",X"30",X"02",
		X"3E",X"99",X"32",X"CA",X"81",X"3E",X"05",X"CD",X"45",X"0C",X"C9",X"D9",X"11",X"C2",X"81",X"3A",
		X"C4",X"81",X"4F",X"21",X"E7",X"13",X"CD",X"60",X"13",X"79",X"32",X"C4",X"81",X"11",X"C3",X"81",
		X"3A",X"C5",X"81",X"4F",X"21",X"17",X"14",X"CD",X"60",X"13",X"79",X"32",X"C5",X"81",X"D9",X"C9",
		X"3A",X"02",X"98",X"2F",X"E6",X"06",X"CB",X"3F",X"47",X"28",X"08",X"D5",X"11",X"0C",X"00",X"19",
		X"10",X"FD",X"D1",X"1A",X"B7",X"C8",X"09",X"AF",X"86",X"08",X"79",X"FE",X"0B",X"20",X"0A",X"D5",
		X"11",X"0C",X"00",X"AF",X"ED",X"52",X"0E",X"FF",X"D1",X"0C",X"23",X"08",X"EB",X"35",X"CD",X"98",
		X"13",X"EB",X"20",X"E4",X"CD",X"1E",X"13",X"C9",X"F5",X"3A",X"C6",X"81",X"3C",X"32",X"C6",X"81",
		X"F1",X"C9",X"3A",X"C9",X"81",X"B7",X"28",X"25",X"3A",X"C8",X"81",X"B7",X"28",X"05",X"3D",X"32",
		X"C8",X"81",X"C9",X"3A",X"C7",X"81",X"B7",X"28",X"0E",X"3E",X"00",X"32",X"02",X"A8",X"32",X"C7",
		X"81",X"3E",X"0C",X"32",X"C8",X"81",X"C9",X"3E",X"00",X"32",X"C9",X"81",X"C9",X"3A",X"C6",X"81",
		X"B7",X"C8",X"3D",X"32",X"C6",X"81",X"3E",X"FF",X"32",X"C9",X"81",X"32",X"C7",X"81",X"32",X"02",
		X"A8",X"3E",X"04",X"32",X"C8",X"81",X"C9",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",
		X"04",X"04",X"04",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"01",X"00",X"00",X"01",X"00",X"00",X"01",X"00",X"00",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"C9",X"DD",X"21",X"2A",X"86",X"21",X"00",X"98",X"CD",
		X"95",X"14",X"DD",X"23",X"23",X"CD",X"95",X"14",X"DD",X"23",X"23",X"CD",X"95",X"14",X"3A",X"69",
		X"86",X"FE",X"02",X"C0",X"3A",X"02",X"98",X"E6",X"08",X"C0",X"3A",X"2D",X"86",X"E6",X"C0",X"6F",
		X"3A",X"2E",X"86",X"E6",X"3C",X"B5",X"32",X"2D",X"86",X"3A",X"2E",X"86",X"CB",X"3F",X"CB",X"3F",
		X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"E6",X"03",X"6F",X"3A",X"2D",X"86",X"E6",X"FC",
		X"B5",X"32",X"2D",X"86",X"C9",X"DD",X"7E",X"00",X"DD",X"46",X"03",X"A8",X"57",X"7E",X"2F",X"4F",
		X"7A",X"A1",X"DD",X"77",X"06",X"DD",X"70",X"00",X"DD",X"71",X"03",X"C9",X"06",X"FF",X"DD",X"7E",
		X"08",X"C6",X"04",X"67",X"DD",X"7E",X"0A",X"6F",X"E5",X"CD",X"FE",X"08",X"7E",X"FE",X"5B",X"38",
		X"06",X"FE",X"A0",X"30",X"02",X"CB",X"80",X"E1",X"E5",X"7C",X"C6",X"06",X"67",X"CD",X"FE",X"08",
		X"7E",X"FE",X"5B",X"38",X"06",X"FE",X"A0",X"30",X"02",X"CB",X"88",X"E1",X"7D",X"C6",X"10",X"6F",
		X"E5",X"CD",X"FE",X"08",X"7E",X"FE",X"5B",X"38",X"06",X"FE",X"A0",X"30",X"02",X"CB",X"A8",X"E1",
		X"7C",X"C6",X"06",X"67",X"CD",X"FE",X"08",X"7E",X"FE",X"5B",X"38",X"06",X"FE",X"A0",X"30",X"02",
		X"CB",X"A0",X"DD",X"7E",X"08",X"67",X"DD",X"7E",X"0A",X"C6",X"04",X"6F",X"E5",X"CD",X"FE",X"08",
		X"7E",X"FE",X"5B",X"38",X"06",X"FE",X"A0",X"30",X"02",X"CB",X"B8",X"E1",X"E5",X"7C",X"C6",X"10",
		X"67",X"CD",X"FE",X"08",X"7E",X"FE",X"5B",X"38",X"06",X"FE",X"A0",X"30",X"02",X"CB",X"90",X"E1",
		X"7D",X"C6",X"06",X"6F",X"E5",X"CD",X"FE",X"08",X"7E",X"FE",X"5B",X"38",X"06",X"FE",X"A0",X"30",
		X"02",X"CB",X"B0",X"E1",X"7C",X"C6",X"10",X"67",X"CD",X"FE",X"08",X"7E",X"FE",X"5B",X"38",X"06",
		X"FE",X"A0",X"30",X"02",X"CB",X"98",X"C9",X"DD",X"7E",X"08",X"C6",X"08",X"67",X"DD",X"7E",X"0A",
		X"C6",X"08",X"6F",X"CD",X"FE",X"08",X"7E",X"DD",X"77",X"0D",X"C9",X"AF",X"32",X"68",X"86",X"21",
		X"F8",X"00",X"01",X"01",X"1F",X"CD",X"01",X"0A",X"11",X"3C",X"80",X"3A",X"3D",X"86",X"4F",X"3A",
		X"3E",X"86",X"81",X"4F",X"3A",X"3F",X"86",X"81",X"4F",X"3A",X"40",X"86",X"81",X"B7",X"CA",X"FA",
		X"15",X"47",X"C5",X"21",X"58",X"16",X"CD",X"67",X"0C",X"E6",X"03",X"CB",X"27",X"06",X"00",X"4F",
		X"09",X"7E",X"12",X"13",X"23",X"7E",X"12",X"13",X"C1",X"10",X"E7",X"21",X"00",X"80",X"3A",X"3D",
		X"86",X"B7",X"28",X"06",X"47",X"0E",X"40",X"CD",X"E5",X"15",X"3A",X"3E",X"86",X"B7",X"28",X"06",
		X"47",X"0E",X"20",X"CD",X"E5",X"15",X"3A",X"3F",X"86",X"B7",X"28",X"06",X"47",X"0E",X"00",X"CD",
		X"E5",X"15",X"3A",X"40",X"86",X"B7",X"28",X"06",X"47",X"0E",X"60",X"CD",X"E5",X"15",X"2B",X"CB",
		X"FE",X"CD",X"FA",X"15",X"C9",X"E5",X"CD",X"67",X"0C",X"E6",X"03",X"11",X"54",X"16",X"26",X"00",
		X"6F",X"19",X"7E",X"B1",X"E1",X"77",X"23",X"10",X"EC",X"C9",X"3A",X"41",X"86",X"B7",X"C0",X"3E",
		X"60",X"32",X"90",X"86",X"21",X"04",X"90",X"06",X"03",X"77",X"23",X"23",X"10",X"FB",X"21",X"00",
		X"00",X"01",X"04",X"1F",X"CD",X"01",X"0A",X"3E",X"93",X"21",X"04",X"88",X"11",X"20",X"00",X"06",
		X"20",X"77",X"19",X"10",X"FC",X"11",X"60",X"16",X"21",X"04",X"89",X"CD",X"46",X"16",X"21",X"03",
		X"89",X"CD",X"46",X"16",X"21",X"02",X"89",X"CD",X"46",X"16",X"3E",X"FF",X"32",X"03",X"A8",X"DF",
		X"11",X"DF",X"18",X"DF",X"25",X"C9",X"06",X"06",X"C5",X"1A",X"77",X"01",X"20",X"00",X"09",X"13",
		X"C1",X"10",X"F5",X"C9",X"04",X"0A",X"12",X"19",X"AC",X"8B",X"2C",X"88",X"B9",X"8B",X"39",X"88",
		X"89",X"8B",X"85",X"87",X"81",X"83",X"88",X"8A",X"84",X"86",X"80",X"82",X"10",X"7F",X"7E",X"7D",
		X"7C",X"10",X"21",X"AC",X"16",X"3A",X"38",X"86",X"BE",X"28",X"14",X"38",X"0C",X"3E",X"FF",X"BE",
		X"28",X"07",X"11",X"06",X"00",X"19",X"C3",X"75",X"16",X"11",X"06",X"00",X"B7",X"ED",X"52",X"23",
		X"7E",X"32",X"3D",X"86",X"23",X"7E",X"32",X"3E",X"86",X"23",X"7E",X"32",X"3F",X"86",X"23",X"7E",
		X"32",X"40",X"86",X"23",X"7E",X"32",X"42",X"86",X"32",X"43",X"86",X"C9",X"01",X"10",X"0A",X"00",
		X"00",X"02",X"02",X"10",X"10",X"00",X"00",X"04",X"03",X"0A",X"0A",X"1E",X"00",X"05",X"04",X"10",
		X"00",X"00",X"28",X"06",X"05",X"14",X"14",X"00",X"00",X"07",X"06",X"10",X"10",X"10",X"00",X"08",
		X"07",X"10",X"10",X"10",X"0C",X"0A",X"08",X"3C",X"00",X"00",X"00",X"0C",X"09",X"00",X"3C",X"00",
		X"00",X"0E",X"0A",X"00",X"00",X"3C",X"00",X"10",X"0B",X"00",X"00",X"00",X"3C",X"12",X"0C",X"20",
		X"1C",X"00",X"00",X"14",X"0D",X"20",X"00",X"1C",X"00",X"16",X"0E",X"10",X"10",X"10",X"0C",X"18",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3E",X"02",X"32",X"8C",X"86",X"21",X"52",X"17",X"06",
		X"00",X"3A",X"38",X"86",X"F5",X"4F",X"09",X"7E",X"32",X"38",X"86",X"CF",X"60",X"F8",X"4C",X"45",
		X"56",X"45",X"4C",X"20",X"00",X"21",X"F8",X"90",X"11",X"38",X"86",X"06",X"02",X"CD",X"66",X"09",
		X"CF",X"18",X"F8",X"41",X"49",X"52",X"20",X"00",X"3A",X"67",X"86",X"FE",X"02",X"20",X"08",X"CF",
		X"A8",X"F8",X"41",X"49",X"52",X"20",X"00",X"F1",X"32",X"38",X"86",X"CD",X"48",X"3A",X"CD",X"86",
		X"59",X"C9",X"00",X"01",X"02",X"03",X"04",X"05",X"06",X"07",X"08",X"09",X"10",X"11",X"12",X"13",
		X"14",X"15",X"16",X"17",X"18",X"19",X"20",X"21",X"22",X"23",X"24",X"25",X"26",X"27",X"28",X"29",
		X"30",X"31",X"32",X"33",X"34",X"35",X"36",X"37",X"38",X"39",X"40",X"41",X"42",X"43",X"44",X"45",
		X"46",X"47",X"48",X"49",X"50",X"51",X"52",X"53",X"54",X"55",X"56",X"57",X"58",X"59",X"60",X"61",
		X"62",X"63",X"64",X"65",X"66",X"67",X"68",X"69",X"70",X"71",X"72",X"73",X"74",X"75",X"76",X"77",
		X"78",X"79",X"80",X"81",X"82",X"83",X"84",X"85",X"86",X"87",X"88",X"89",X"90",X"91",X"92",X"93",
		X"94",X"95",X"96",X"97",X"98",X"99",X"3E",X"00",X"32",X"01",X"A8",X"32",X"02",X"A8",X"32",X"03",
		X"A8",X"32",X"04",X"A8",X"32",X"07",X"A8",X"32",X"06",X"A8",X"3E",X"9B",X"32",X"03",X"98",X"3E",
		X"88",X"32",X"03",X"A0",X"31",X"1C",X"81",X"21",X"1C",X"81",X"0E",X"08",X"CD",X"F6",X"09",X"3E",
		X"FF",X"32",X"C0",X"81",X"32",X"C1",X"81",X"21",X"A6",X"18",X"11",X"CB",X"81",X"01",X"3C",X"00",
		X"ED",X"B0",X"31",X"1C",X"81",X"21",X"00",X"90",X"0E",X"01",X"CD",X"F6",X"09",X"CD",X"53",X"18",
		X"CD",X"E2",X"18",X"3E",X"01",X"CD",X"70",X"18",X"CD",X"7B",X"1C",X"3E",X"01",X"CD",X"70",X"18",
		X"CD",X"16",X"18",X"C3",X"FD",X"17",X"3E",X"FF",X"32",X"66",X"86",X"3E",X"01",X"32",X"38",X"86",
		X"AF",X"32",X"7F",X"86",X"32",X"80",X"86",X"32",X"81",X"86",X"32",X"AB",X"86",X"3E",X"02",X"32",
		X"67",X"86",X"21",X"33",X"86",X"CD",X"AA",X"29",X"CD",X"72",X"16",X"21",X"47",X"86",X"CD",X"AA",
		X"29",X"CD",X"72",X"16",X"CD",X"D5",X"29",X"3E",X"00",X"32",X"33",X"86",X"32",X"47",X"86",X"CD",
		X"45",X"0C",X"C9",X"E1",X"22",X"61",X"86",X"32",X"63",X"86",X"CD",X"9B",X"0E",X"CD",X"94",X"0C",
		X"AF",X"32",X"BF",X"81",X"3E",X"FF",X"32",X"01",X"A8",X"2A",X"61",X"86",X"3A",X"63",X"86",X"E9",
		X"F5",X"3E",X"1E",X"CD",X"7B",X"18",X"F1",X"3D",X"20",X"F6",X"C9",X"F5",X"D5",X"E5",X"C5",X"DD",
		X"2A",X"B6",X"81",X"DD",X"CB",X"00",X"EE",X"DD",X"36",X"03",X"01",X"CD",X"67",X"0C",X"CD",X"0B",
		X"28",X"3A",X"65",X"86",X"B7",X"C4",X"8E",X"0A",X"DD",X"CB",X"00",X"6E",X"20",X"ED",X"C1",X"E1",
		X"D1",X"F1",X"3D",X"20",X"D6",X"C9",X"01",X"04",X"80",X"4A",X"4D",X"48",X"01",X"01",X"00",X"52",
		X"41",X"51",X"00",X"39",X"10",X"55",X"52",X"4C",X"00",X"28",X"70",X"4D",X"53",X"20",X"00",X"18",
		X"30",X"45",X"4C",X"50",X"00",X"17",X"70",X"4A",X"49",X"4D",X"00",X"16",X"40",X"42",X"49",X"4C",
		X"00",X"15",X"90",X"44",X"41",X"4E",X"00",X"14",X"10",X"41",X"50",X"48",X"00",X"12",X"00",X"4F",
		X"42",X"45",X"CD",X"C1",X"09",X"CD",X"69",X"1D",X"CD",X"6C",X"0A",X"CD",X"8E",X"0A",X"CF",X"28",
		X"00",X"20",X"54",X"41",X"47",X"4F",X"20",X"50",X"52",X"4F",X"55",X"44",X"4C",X"59",X"20",X"50",
		X"52",X"45",X"53",X"45",X"4E",X"54",X"53",X"00",X"CF",X"60",X"18",X"43",X"41",X"4C",X"49",X"50",
		X"53",X"4F",X"00",X"E7",X"06",X"07",X"05",X"E7",X"06",X"0D",X"02",X"E7",X"07",X"13",X"07",X"DF",
		X"30",X"CF",X"40",X"30",X"20",X"54",X"4F",X"50",X"20",X"31",X"30",X"20",X"53",X"43",X"4F",X"52",
		X"45",X"53",X"20",X"00",X"11",X"CB",X"81",X"21",X"40",X"38",X"3E",X"01",X"08",X"D5",X"EB",X"7E",
		X"23",X"B6",X"23",X"B6",X"EB",X"D1",X"C8",X"E5",X"D5",X"08",X"32",X"00",X"80",X"08",X"06",X"02",
		X"11",X"00",X"80",X"CD",X"66",X"09",X"01",X"00",X"20",X"09",X"D1",X"06",X"06",X"CD",X"66",X"09",
		X"13",X"13",X"13",X"01",X"00",X"30",X"09",X"CD",X"FE",X"08",X"06",X"03",X"3E",X"20",X"CD",X"A9",
		X"09",X"10",X"F9",X"06",X"03",X"1A",X"13",X"CD",X"A9",X"09",X"10",X"F9",X"E1",X"01",X"10",X"00",
		X"09",X"08",X"C6",X"01",X"27",X"FE",X"11",X"DA",X"3C",X"19",X"06",X"05",X"C5",X"DF",X"19",X"3E",
		X"02",X"CD",X"7B",X"18",X"DF",X"1A",X"3E",X"02",X"CD",X"7B",X"18",X"DF",X"1B",X"3E",X"02",X"CD",
		X"7B",X"18",X"DF",X"1C",X"3E",X"02",X"CD",X"7B",X"18",X"DF",X"1D",X"3E",X"02",X"CD",X"7B",X"18",
		X"DF",X"1E",X"3E",X"02",X"CD",X"7B",X"18",X"DF",X"1F",X"3E",X"02",X"CD",X"7B",X"18",X"DF",X"18",
		X"3E",X"02",X"CD",X"7B",X"18",X"C1",X"10",X"C4",X"C9",X"0E",X"0A",X"11",X"CB",X"81",X"E5",X"D5",
		X"06",X"03",X"1A",X"BE",X"38",X"11",X"20",X"04",X"13",X"23",X"10",X"F6",X"D1",X"21",X"06",X"00",
		X"19",X"EB",X"E1",X"0D",X"20",X"E8",X"C9",X"D1",X"D5",X"0D",X"28",X"16",X"06",X"00",X"21",X"00",
		X"00",X"09",X"29",X"09",X"29",X"E5",X"19",X"2B",X"54",X"5D",X"01",X"06",X"00",X"09",X"EB",X"C1",
		X"ED",X"B8",X"D1",X"E1",X"01",X"03",X"00",X"ED",X"B0",X"D5",X"CD",X"C1",X"09",X"CD",X"88",X"29",
		X"CD",X"C8",X"0A",X"DF",X"1A",X"3A",X"8A",X"86",X"FE",X"01",X"20",X"1E",X"CF",X"20",X"28",X"43",
		X"4F",X"4E",X"47",X"52",X"41",X"54",X"55",X"4C",X"41",X"54",X"49",X"4F",X"4E",X"53",X"20",X"50",
		X"4C",X"41",X"59",X"45",X"52",X"20",X"31",X"00",X"18",X"1C",X"CF",X"20",X"28",X"43",X"4F",X"4E",
		X"47",X"52",X"41",X"54",X"55",X"4C",X"41",X"54",X"49",X"4F",X"4E",X"53",X"20",X"50",X"4C",X"41",
		X"59",X"45",X"52",X"20",X"32",X"00",X"E7",X"16",X"00",X"04",X"DF",X"4E",X"CF",X"38",X"38",X"59",
		X"4F",X"55",X"20",X"48",X"41",X"56",X"45",X"20",X"4D",X"41",X"44",X"45",X"20",X"54",X"48",X"45",
		X"00",X"CF",X"60",X"48",X"43",X"41",X"4C",X"49",X"50",X"53",X"4F",X"00",X"CF",X"50",X"58",X"48",
		X"41",X"4C",X"4C",X"20",X"4F",X"46",X"20",X"46",X"41",X"4D",X"45",X"00",X"E7",X"03",X"0F",X"05",
		X"CF",X"28",X"78",X"45",X"4E",X"54",X"45",X"52",X"20",X"59",X"4F",X"55",X"52",X"20",X"49",X"4E",
		X"49",X"54",X"49",X"41",X"4C",X"53",X"20",X"5B",X"00",X"CF",X"70",X"88",X"5B",X"5B",X"5B",X"00",
		X"E7",X"03",X"16",X"07",X"CF",X"20",X"B0",X"4D",X"4F",X"56",X"45",X"20",X"53",X"54",X"49",X"43",
		X"4B",X"20",X"4C",X"45",X"46",X"54",X"20",X"4F",X"52",X"20",X"52",X"49",X"47",X"48",X"54",X"00",
		X"CF",X"30",X"C0",X"54",X"4F",X"20",X"43",X"48",X"41",X"4E",X"47",X"45",X"20",X"54",X"48",X"45",
		X"20",X"4C",X"45",X"54",X"54",X"45",X"52",X"00",X"CF",X"20",X"D0",X"50",X"55",X"4C",X"4C",X"20",
		X"53",X"54",X"49",X"43",X"4B",X"20",X"44",X"4F",X"57",X"4E",X"20",X"54",X"4F",X"20",X"45",X"4E",
		X"54",X"45",X"52",X"00",X"E1",X"E5",X"06",X"03",X"36",X"20",X"23",X"10",X"FB",X"21",X"88",X"70",
		X"CD",X"FE",X"08",X"D1",X"06",X"03",X"0E",X"41",X"3E",X"C8",X"32",X"61",X"86",X"CD",X"4C",X"1B",
		X"20",X"FB",X"79",X"E5",X"CD",X"A9",X"09",X"C5",X"D5",X"3E",X"09",X"CD",X"7B",X"18",X"D1",X"C1",
		X"E1",X"3A",X"61",X"86",X"3D",X"32",X"61",X"86",X"C8",X"CD",X"4C",X"1B",X"20",X"05",X"CD",X"5C",
		X"1B",X"18",X"DA",X"79",X"12",X"13",X"CD",X"A9",X"09",X"10",X"CD",X"C9",X"3A",X"8A",X"86",X"FE",
		X"02",X"3A",X"2E",X"86",X"28",X"03",X"3A",X"2D",X"86",X"E6",X"08",X"C9",X"F5",X"D5",X"3A",X"8A",
		X"86",X"FE",X"02",X"3A",X"2E",X"86",X"28",X"03",X"3A",X"2D",X"86",X"57",X"79",X"CB",X"62",X"28",
		X"0A",X"C6",X"01",X"FE",X"5B",X"38",X"10",X"3E",X"40",X"18",X"0C",X"CB",X"6A",X"28",X"08",X"D6",
		X"01",X"FE",X"40",X"30",X"02",X"3E",X"5A",X"4F",X"D1",X"F1",X"C9",X"3A",X"66",X"86",X"B7",X"C0",
		X"3E",X"FF",X"32",X"64",X"86",X"21",X"07",X"82",X"1E",X"04",X"23",X"23",X"23",X"CB",X"38",X"08",
		X"04",X"2B",X"1D",X"10",X"FC",X"08",X"30",X"08",X"CB",X"21",X"CB",X"21",X"CB",X"21",X"CB",X"21",
		X"79",X"86",X"27",X"77",X"30",X"08",X"2B",X"1D",X"28",X"04",X"0E",X"01",X"18",X"F2",X"CD",X"FB",
		X"1B",X"EB",X"2A",X"3A",X"86",X"7A",X"BC",X"D8",X"7B",X"BD",X"D8",X"3A",X"33",X"86",X"C6",X"01",
		X"27",X"32",X"33",X"86",X"3E",X"0F",X"CD",X"45",X"0C",X"CD",X"E0",X"1B",X"CD",X"1B",X"0B",X"C9",
		X"2A",X"3A",X"86",X"1E",X"30",X"16",X"00",X"06",X"04",X"CB",X"23",X"CB",X"12",X"10",X"FA",X"7D",
		X"83",X"27",X"6F",X"7C",X"8A",X"27",X"67",X"22",X"3A",X"86",X"C9",X"21",X"07",X"82",X"7E",X"23",
		X"6E",X"67",X"C9",X"3A",X"66",X"86",X"B7",X"C0",X"3E",X"FF",X"32",X"64",X"86",X"21",X"0A",X"82",
		X"1E",X"04",X"23",X"23",X"23",X"CB",X"38",X"08",X"04",X"2B",X"1D",X"10",X"FC",X"08",X"30",X"08",
		X"CB",X"21",X"CB",X"21",X"CB",X"21",X"CB",X"21",X"79",X"86",X"27",X"77",X"30",X"08",X"2B",X"1D",
		X"28",X"04",X"0E",X"01",X"18",X"F2",X"CD",X"73",X"1C",X"EB",X"2A",X"4E",X"86",X"7A",X"BC",X"D8",
		X"7B",X"BD",X"D8",X"3A",X"47",X"86",X"C6",X"01",X"27",X"32",X"47",X"86",X"3E",X"0F",X"CD",X"45",
		X"0C",X"CD",X"58",X"1C",X"CD",X"1B",X"0B",X"C9",X"2A",X"4E",X"86",X"1E",X"30",X"16",X"00",X"06",
		X"04",X"CB",X"23",X"CB",X"12",X"10",X"FA",X"7D",X"83",X"27",X"6F",X"7C",X"8A",X"27",X"67",X"22",
		X"4E",X"86",X"C9",X"21",X"0A",X"82",X"7E",X"23",X"6E",X"67",X"C9",X"CD",X"C1",X"09",X"3E",X"00",
		X"32",X"07",X"A8",X"32",X"06",X"A8",X"3E",X"01",X"32",X"69",X"86",X"AF",X"32",X"38",X"86",X"CD",
		X"B0",X"4B",X"CD",X"69",X"1D",X"CD",X"6C",X"0A",X"CD",X"8E",X"0A",X"E7",X"02",X"00",X"02",X"CF",
		X"28",X"00",X"20",X"54",X"41",X"47",X"4F",X"20",X"50",X"52",X"4F",X"55",X"44",X"4C",X"59",X"20",
		X"50",X"52",X"45",X"53",X"45",X"4E",X"54",X"53",X"00",X"CF",X"28",X"08",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"00",X"DF",X"AF",X"CF",X"10",X"A8",X"45",X"58",X"54",X"52",X"41",X"20",X"4D",X"41",
		X"4E",X"20",X"45",X"56",X"45",X"52",X"59",X"20",X"33",X"30",X"30",X"30",X"30",X"20",X"50",X"4F",
		X"49",X"4E",X"54",X"53",X"00",X"3E",X"01",X"CD",X"70",X"18",X"CF",X"10",X"C8",X"50",X"4C",X"41",
		X"59",X"20",X"20",X"31",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"4F",X"52",X"20",X"54",
		X"45",X"41",X"4D",X"5B",X"50",X"4C",X"41",X"59",X"20",X"00",X"06",X"08",X"C5",X"DF",X"C9",X"3E",
		X"02",X"CD",X"7B",X"18",X"DF",X"CA",X"3E",X"02",X"CD",X"7B",X"18",X"DF",X"CB",X"3E",X"02",X"CD",
		X"7B",X"18",X"DF",X"CC",X"3E",X"02",X"CD",X"7B",X"18",X"DF",X"CD",X"3E",X"02",X"CD",X"7B",X"18",
		X"DF",X"CE",X"3E",X"02",X"CD",X"7B",X"18",X"DF",X"CF",X"3E",X"02",X"CD",X"7B",X"18",X"DF",X"C8",
		X"3E",X"02",X"CD",X"7B",X"18",X"C1",X"10",X"C4",X"3E",X"02",X"CD",X"70",X"18",X"21",X"A8",X"10",
		X"01",X"08",X"1C",X"CD",X"01",X"0A",X"C3",X"68",X"0B",X"3A",X"2D",X"86",X"CB",X"57",X"C8",X"3A",
		X"2D",X"86",X"CB",X"4F",X"C8",X"CB",X"47",X"C8",X"21",X"81",X"88",X"11",X"20",X"00",X"3A",X"82",
		X"86",X"E6",X"0F",X"CD",X"DD",X"1D",X"3A",X"82",X"86",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",
		X"3F",X"CD",X"DD",X"1D",X"3A",X"83",X"86",X"E6",X"0F",X"CD",X"DD",X"1D",X"3A",X"83",X"86",X"CB",
		X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CD",X"DD",X"1D",X"21",X"01",X"8B",X"11",X"20",X"00",
		X"3A",X"84",X"86",X"E6",X"0F",X"CD",X"DD",X"1D",X"3A",X"84",X"86",X"CB",X"3F",X"CB",X"3F",X"CB",
		X"3F",X"CB",X"3F",X"CD",X"DD",X"1D",X"3A",X"85",X"86",X"E6",X"0F",X"CD",X"DD",X"1D",X"3A",X"85",
		X"86",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CD",X"DD",X"1D",X"C9",X"01",X"E6",X"1D",
		X"81",X"4F",X"0A",X"77",X"19",X"C9",X"00",X"01",X"02",X"03",X"04",X"05",X"06",X"07",X"08",X"09",
		X"11",X"12",X"13",X"14",X"15",X"16",X"17",X"18",X"CD",X"50",X"0D",X"D2",X"12",X"0E",X"CD",X"F2",
		X"0C",X"D2",X"61",X"1F",X"FD",X"2A",X"B6",X"81",X"FD",X"66",X"02",X"FD",X"6E",X"01",X"E5",X"DD",
		X"E1",X"CD",X"BD",X"1F",X"FD",X"CB",X"00",X"F6",X"FD",X"CB",X"0C",X"D6",X"FD",X"CB",X"00",X"D6",
		X"FD",X"36",X"0D",X"00",X"DD",X"E5",X"CD",X"EE",X"0D",X"FD",X"E1",X"DD",X"7E",X"0D",X"B7",X"C2",
		X"36",X"1F",X"CD",X"3C",X"1E",X"FD",X"E5",X"CD",X"EE",X"0D",X"18",X"ED",X"DD",X"7E",X"0B",X"E6",
		X"07",X"4F",X"5F",X"DD",X"36",X"0B",X"00",X"DD",X"CB",X"0B",X"FE",X"FD",X"CB",X"00",X"4E",X"20",
		X"2A",X"CD",X"67",X"0C",X"E6",X"0F",X"CB",X"D7",X"FD",X"77",X"01",X"FD",X"CB",X"00",X"CE",X"C5",
		X"CD",X"15",X"1F",X"21",X"05",X"1F",X"06",X"00",X"09",X"5E",X"C1",X"CD",X"67",X"0C",X"FE",X"64",
		X"38",X"09",X"E6",X"07",X"28",X"F5",X"FE",X"04",X"28",X"F1",X"5F",X"CD",X"AC",X"14",X"16",X"00",
		X"CB",X"23",X"21",X"02",X"20",X"19",X"19",X"19",X"11",X"00",X"00",X"FD",X"36",X"04",X"00",X"FD",
		X"36",X"03",X"00",X"FD",X"36",X"0A",X"00",X"FD",X"36",X"09",X"00",X"78",X"A6",X"BE",X"28",X"0D",
		X"78",X"23",X"23",X"A6",X"BE",X"28",X"06",X"78",X"23",X"23",X"A6",X"BE",X"C0",X"23",X"7E",X"B9",
		X"20",X"04",X"DD",X"CB",X"0B",X"BE",X"5F",X"DD",X"7E",X"0B",X"E6",X"F8",X"B3",X"DD",X"77",X"0B",
		X"CB",X"23",X"CB",X"23",X"21",X"42",X"20",X"19",X"7E",X"FD",X"77",X"03",X"23",X"7E",X"FD",X"77",
		X"04",X"23",X"7E",X"FD",X"77",X"09",X"23",X"7E",X"FD",X"77",X"0A",X"DD",X"CB",X"0B",X"7E",X"C8",
		X"DD",X"CB",X"0B",X"BE",X"DD",X"4E",X"0B",X"06",X"00",X"21",X"32",X"20",X"09",X"09",X"7E",X"23",
		X"66",X"6F",X"DD",X"CB",X"00",X"A6",X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",X"36",X"04",X"01",
		X"DD",X"CB",X"00",X"E6",X"C9",X"00",X"06",X"04",X"05",X"02",X"00",X"03",X"00",X"00",X"07",X"00",
		X"00",X"01",X"00",X"00",X"00",X"0E",X"00",X"3A",X"73",X"82",X"FD",X"BE",X"0C",X"38",X"04",X"CB",
		X"C9",X"18",X"04",X"28",X"02",X"CB",X"D9",X"3A",X"6D",X"82",X"FD",X"BE",X"06",X"38",X"03",X"CB",
		X"D1",X"C9",X"C8",X"CB",X"C1",X"C9",X"CB",X"77",X"28",X"08",X"01",X"02",X"02",X"CD",X"8B",X"1B",
		X"18",X"0A",X"CB",X"7F",X"28",X"06",X"01",X"02",X"02",X"CD",X"03",X"1C",X"3E",X"05",X"CD",X"45",
		X"0C",X"CD",X"69",X"1F",X"21",X"43",X"86",X"35",X"2B",X"7E",X"B7",X"28",X"04",X"35",X"C3",X"04",
		X"1E",X"CD",X"68",X"0E",X"CD",X"EE",X"0D",X"18",X"FB",X"AF",X"DD",X"77",X"0D",X"FD",X"77",X"04",
		X"FD",X"77",X"03",X"FD",X"77",X"0A",X"FD",X"77",X"09",X"DD",X"CB",X"0C",X"96",X"DD",X"CB",X"00",
		X"A6",X"DD",X"CB",X"00",X"B6",X"21",X"4A",X"21",X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",X"36",
		X"04",X"01",X"DD",X"CB",X"00",X"E6",X"CD",X"EE",X"0D",X"DD",X"CB",X"00",X"66",X"20",X"F7",X"DD",
		X"36",X"0A",X"00",X"DD",X"36",X"08",X"00",X"DD",X"66",X"02",X"DD",X"6E",X"01",X"E5",X"FD",X"E1",
		X"FD",X"36",X"06",X"00",X"FD",X"36",X"0C",X"00",X"DD",X"CB",X"00",X"96",X"C9",X"CD",X"67",X"0C",
		X"CB",X"6F",X"28",X"1F",X"FD",X"36",X"08",X"02",X"FD",X"36",X"0A",X"C8",X"21",X"7F",X"20",X"FD",
		X"75",X"05",X"FD",X"74",X"06",X"FD",X"36",X"04",X"01",X"FD",X"CB",X"00",X"E6",X"3E",X"02",X"FD",
		X"77",X"0B",X"C9",X"FD",X"36",X"08",X"EE",X"FD",X"36",X"0A",X"C8",X"21",X"62",X"20",X"FD",X"75",
		X"05",X"FD",X"74",X"06",X"FD",X"36",X"04",X"01",X"FD",X"CB",X"00",X"E6",X"3E",X"06",X"FD",X"77",
		X"0B",X"C9",X"03",X"00",X"03",X"00",X"03",X"00",X"0F",X"01",X"0C",X"02",X"03",X"00",X"0C",X"02",
		X"0C",X"02",X"0C",X"02",X"3C",X"03",X"30",X"04",X"0C",X"02",X"30",X"04",X"30",X"04",X"30",X"04",
		X"F0",X"05",X"C0",X"06",X"30",X"04",X"C0",X"06",X"C0",X"06",X"C0",X"06",X"C3",X"07",X"03",X"00",
		X"C0",X"06",X"9C",X"20",X"F3",X"20",X"7F",X"20",X"2D",X"21",X"B9",X"20",X"10",X"21",X"62",X"20",
		X"D6",X"20",X"00",X"00",X"00",X"FE",X"00",X"03",X"00",X"FE",X"00",X"03",X"00",X"00",X"00",X"03",
		X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"FD",X"00",X"02",X"00",X"FD",X"00",X"00",X"00",X"FD",
		X"00",X"FE",X"00",X"00",X"01",X"00",X"00",X"0C",X"0C",X"05",X"59",X"07",X"0C",X"0C",X"04",X"5A",
		X"07",X"0C",X"0C",X"05",X"5B",X"07",X"0C",X"0C",X"04",X"5A",X"07",X"00",X"01",X"67",X"20",X"00",
		X"00",X"01",X"00",X"00",X"0C",X"0C",X"04",X"5C",X"07",X"0C",X"0C",X"03",X"5D",X"07",X"0C",X"0C",
		X"05",X"5E",X"07",X"0C",X"0C",X"03",X"5D",X"07",X"00",X"01",X"84",X"20",X"00",X"00",X"01",X"00",
		X"00",X"0C",X"0C",X"04",X"5F",X"07",X"0C",X"0C",X"03",X"60",X"07",X"0C",X"0C",X"05",X"61",X"07",
		X"0C",X"0C",X"03",X"60",X"07",X"00",X"01",X"A1",X"20",X"00",X"00",X"01",X"00",X"00",X"0C",X"0C",
		X"04",X"62",X"07",X"0C",X"0C",X"03",X"63",X"07",X"0C",X"0C",X"05",X"64",X"07",X"0C",X"0C",X"03",
		X"63",X"07",X"00",X"01",X"BE",X"20",X"00",X"00",X"01",X"00",X"00",X"0C",X"0C",X"05",X"5F",X"07",
		X"0C",X"0C",X"04",X"60",X"07",X"0C",X"0C",X"05",X"61",X"07",X"0C",X"0C",X"04",X"60",X"07",X"00",
		X"01",X"DB",X"20",X"00",X"00",X"01",X"00",X"00",X"0C",X"0C",X"04",X"62",X"07",X"0C",X"0C",X"03",
		X"63",X"07",X"0C",X"0C",X"05",X"64",X"07",X"0C",X"0C",X"03",X"63",X"07",X"00",X"01",X"F8",X"20",
		X"00",X"00",X"01",X"00",X"00",X"0C",X"0C",X"04",X"65",X"07",X"0C",X"0C",X"03",X"66",X"07",X"0C",
		X"0C",X"05",X"67",X"07",X"0C",X"0C",X"03",X"66",X"07",X"00",X"01",X"15",X"21",X"00",X"00",X"01",
		X"00",X"00",X"0C",X"0C",X"04",X"68",X"07",X"0C",X"0C",X"03",X"69",X"07",X"0C",X"0C",X"05",X"6A",
		X"07",X"0C",X"0C",X"03",X"69",X"07",X"00",X"01",X"32",X"21",X"00",X"00",X"01",X"00",X"00",X"01",
		X"00",X"01",X"CA",X"00",X"01",X"00",X"01",X"CA",X"01",X"01",X"00",X"01",X"CA",X"02",X"01",X"00",
		X"01",X"CA",X"03",X"01",X"00",X"01",X"CA",X"04",X"01",X"00",X"01",X"CA",X"05",X"01",X"00",X"01",
		X"CA",X"06",X"01",X"00",X"01",X"CA",X"07",X"01",X"00",X"01",X"C5",X"00",X"01",X"00",X"01",X"C5",
		X"01",X"01",X"00",X"01",X"C5",X"02",X"01",X"00",X"01",X"C5",X"03",X"01",X"00",X"01",X"C5",X"04",
		X"01",X"00",X"01",X"C5",X"05",X"01",X"00",X"01",X"C5",X"06",X"01",X"00",X"01",X"C5",X"07",X"01",
		X"00",X"01",X"C6",X"00",X"01",X"00",X"01",X"C6",X"01",X"01",X"00",X"01",X"C6",X"02",X"01",X"00",
		X"01",X"C6",X"03",X"01",X"00",X"01",X"C6",X"04",X"01",X"00",X"01",X"C6",X"05",X"01",X"00",X"01",
		X"C6",X"06",X"01",X"00",X"01",X"C6",X"07",X"01",X"00",X"01",X"C7",X"00",X"01",X"00",X"01",X"C7",
		X"01",X"01",X"00",X"01",X"C7",X"02",X"01",X"00",X"01",X"C7",X"03",X"01",X"00",X"01",X"C7",X"04",
		X"01",X"00",X"01",X"C7",X"05",X"01",X"00",X"01",X"C7",X"06",X"01",X"00",X"01",X"C7",X"07",X"01",
		X"00",X"01",X"C8",X"00",X"01",X"00",X"01",X"C8",X"01",X"01",X"00",X"01",X"C8",X"02",X"01",X"00",
		X"01",X"C8",X"03",X"01",X"00",X"01",X"C8",X"04",X"01",X"00",X"01",X"C8",X"05",X"01",X"00",X"01",
		X"C8",X"06",X"01",X"00",X"01",X"C8",X"07",X"01",X"00",X"01",X"C9",X"00",X"01",X"00",X"01",X"C9",
		X"01",X"01",X"00",X"01",X"C9",X"02",X"01",X"00",X"01",X"C9",X"03",X"01",X"00",X"01",X"C9",X"04",
		X"01",X"00",X"01",X"C9",X"05",X"01",X"00",X"01",X"C9",X"06",X"01",X"00",X"01",X"C9",X"07",X"00",
		X"00",X"00",X"00",X"CD",X"50",X"0D",X"D2",X"12",X"0E",X"CD",X"F2",X"0C",X"D2",X"CD",X"23",X"3E",
		X"1E",X"CD",X"42",X"0E",X"DD",X"66",X"02",X"DD",X"6E",X"01",X"E5",X"FD",X"E1",X"CD",X"D5",X"23",
		X"DD",X"CB",X"00",X"F6",X"DD",X"CB",X"0C",X"D6",X"DD",X"CB",X"00",X"D6",X"DD",X"36",X"0D",X"00",
		X"FD",X"E5",X"FD",X"E1",X"DD",X"7E",X"0D",X"B7",X"C2",X"AC",X"23",X"FD",X"CB",X"00",X"56",X"20",
		X"13",X"CD",X"67",X"0C",X"E6",X"0F",X"CB",X"CF",X"FD",X"77",X"02",X"FD",X"CB",X"00",X"D6",X"3E",
		X"0A",X"CD",X"45",X"0C",X"CD",X"9E",X"22",X"FD",X"E5",X"CD",X"EE",X"0D",X"18",X"D4",X"DD",X"7E",
		X"0B",X"E6",X"07",X"4F",X"5F",X"DD",X"36",X"0B",X"00",X"DD",X"CB",X"0B",X"FE",X"FD",X"CB",X"00",
		X"4E",X"20",X"2A",X"CD",X"67",X"0C",X"E6",X"0F",X"CB",X"D7",X"FD",X"77",X"01",X"FD",X"CB",X"00",
		X"CE",X"C5",X"CD",X"83",X"23",X"21",X"73",X"23",X"06",X"00",X"09",X"5E",X"C1",X"CD",X"67",X"0C",
		X"FE",X"C8",X"38",X"09",X"E6",X"07",X"28",X"F5",X"FE",X"04",X"28",X"F1",X"5F",X"CD",X"AC",X"14",
		X"16",X"00",X"CB",X"23",X"21",X"18",X"24",X"19",X"19",X"19",X"11",X"00",X"00",X"FD",X"36",X"04",
		X"00",X"FD",X"36",X"03",X"00",X"FD",X"36",X"0A",X"00",X"FD",X"36",X"09",X"00",X"78",X"A6",X"BE",
		X"28",X"0D",X"78",X"23",X"23",X"A6",X"BE",X"28",X"06",X"78",X"23",X"23",X"A6",X"BE",X"C0",X"23",
		X"7E",X"B9",X"20",X"04",X"DD",X"CB",X"0B",X"BE",X"5F",X"DD",X"7E",X"0B",X"E6",X"F8",X"B3",X"DD",
		X"77",X"0B",X"CB",X"23",X"CB",X"23",X"3A",X"2C",X"86",X"CB",X"5F",X"28",X"05",X"21",X"58",X"24",
		X"18",X"03",X"21",X"78",X"24",X"19",X"7E",X"FD",X"77",X"03",X"23",X"7E",X"FD",X"77",X"04",X"23",
		X"7E",X"FD",X"77",X"09",X"23",X"7E",X"FD",X"77",X"0A",X"DD",X"CB",X"0B",X"7E",X"C8",X"DD",X"CB",
		X"0B",X"BE",X"DD",X"4E",X"0B",X"06",X"00",X"21",X"48",X"24",X"09",X"09",X"7E",X"23",X"66",X"6F",
		X"DD",X"CB",X"00",X"A6",X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",X"36",X"04",X"01",X"DD",X"CB",
		X"00",X"E6",X"C9",X"00",X"06",X"04",X"05",X"02",X"00",X"03",X"00",X"00",X"07",X"00",X"00",X"01",
		X"00",X"00",X"00",X"DD",X"E5",X"DD",X"2A",X"A8",X"86",X"DD",X"7E",X"0A",X"FD",X"BE",X"0C",X"38",
		X"04",X"CB",X"C9",X"18",X"04",X"28",X"02",X"CB",X"D9",X"DD",X"7E",X"08",X"FD",X"BE",X"06",X"38",
		X"05",X"CB",X"D1",X"DD",X"E1",X"C9",X"C8",X"CB",X"C1",X"DD",X"E1",X"C9",X"CB",X"77",X"28",X"08",
		X"01",X"01",X"02",X"CD",X"8B",X"1B",X"18",X"0A",X"CB",X"7F",X"28",X"06",X"01",X"01",X"02",X"CD",
		X"03",X"1C",X"3E",X"05",X"CD",X"45",X"0C",X"CD",X"69",X"1F",X"C3",X"4F",X"22",X"CD",X"68",X"0E",
		X"CD",X"EE",X"0D",X"18",X"FB",X"3E",X"0A",X"CD",X"45",X"0C",X"21",X"08",X"24",X"3A",X"38",X"86",
		X"E6",X"07",X"CB",X"27",X"16",X"00",X"5F",X"19",X"5E",X"23",X"56",X"DD",X"73",X"08",X"DD",X"72",
		X"0A",X"21",X"B5",X"24",X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",X"36",X"04",X"01",X"DD",X"CB",
		X"00",X"E6",X"3E",X"02",X"DD",X"77",X"0B",X"C9",X"51",X"E0",X"DB",X"DF",X"A1",X"E2",X"DB",X"E2",
		X"D5",X"68",X"85",X"A1",X"95",X"E6",X"D5",X"E6",X"03",X"00",X"03",X"00",X"03",X"00",X"0F",X"01",
		X"0C",X"02",X"03",X"00",X"0C",X"02",X"0C",X"02",X"0C",X"02",X"3C",X"03",X"30",X"04",X"0C",X"02",
		X"30",X"04",X"30",X"04",X"30",X"04",X"F0",X"05",X"C0",X"06",X"30",X"04",X"C0",X"06",X"C0",X"06",
		X"C0",X"06",X"C3",X"07",X"03",X"00",X"C0",X"06",X"D2",X"24",X"D2",X"24",X"B5",X"24",X"EF",X"24",
		X"EF",X"24",X"EF",X"24",X"98",X"24",X"D2",X"24",X"00",X"00",X"C0",X"FE",X"A0",X"01",X"C0",X"FE",
		X"00",X"01",X"00",X"00",X"00",X"01",X"7F",X"01",X"00",X"00",X"7F",X"01",X"00",X"FE",X"7F",X"01",
		X"00",X"FE",X"00",X"00",X"A0",X"FE",X"C0",X"FE",X"00",X"00",X"C0",X"FD",X"A0",X"01",X"C0",X"FD",
		X"C0",X"01",X"00",X"00",X"00",X"01",X"7F",X"02",X"00",X"00",X"7F",X"02",X"00",X"FE",X"7F",X"02",
		X"00",X"FD",X"00",X"00",X"A0",X"FE",X"C0",X"FD",X"00",X"00",X"01",X"00",X"00",X"0C",X"0C",X"06",
		X"6B",X"03",X"0C",X"0C",X"06",X"6C",X"03",X"0C",X"0C",X"06",X"6D",X"03",X"0C",X"0C",X"06",X"6C",
		X"03",X"00",X"01",X"9D",X"24",X"00",X"00",X"01",X"00",X"00",X"0C",X"0C",X"06",X"6B",X"03",X"0C",
		X"0C",X"06",X"6C",X"03",X"0C",X"0C",X"06",X"6D",X"03",X"0C",X"0C",X"06",X"6C",X"03",X"00",X"01",
		X"BA",X"24",X"00",X"00",X"01",X"00",X"00",X"0C",X"0C",X"06",X"6B",X"03",X"0C",X"0C",X"06",X"6C",
		X"03",X"0C",X"0C",X"06",X"6D",X"03",X"0C",X"0C",X"06",X"6C",X"03",X"00",X"01",X"D7",X"24",X"00",
		X"00",X"01",X"00",X"00",X"0C",X"0C",X"06",X"6B",X"03",X"0C",X"0C",X"06",X"6C",X"03",X"0C",X"0C",
		X"06",X"6D",X"03",X"0C",X"0C",X"06",X"6C",X"03",X"00",X"01",X"F4",X"24",X"C9",X"CD",X"50",X"0D",
		X"D2",X"12",X"0E",X"CD",X"F2",X"0C",X"D2",X"76",X"26",X"FD",X"2A",X"B6",X"81",X"FD",X"66",X"02",
		X"FD",X"6E",X"01",X"E5",X"DD",X"E1",X"CD",X"7E",X"26",X"FD",X"CB",X"00",X"F6",X"FD",X"CB",X"0C",
		X"D6",X"FD",X"CB",X"00",X"D6",X"FD",X"36",X"0D",X"00",X"DD",X"E5",X"CD",X"EE",X"0D",X"FD",X"E1",
		X"DD",X"7E",X"0D",X"B7",X"C2",X"4B",X"26",X"CD",X"51",X"25",X"FD",X"E5",X"CD",X"EE",X"0D",X"18",
		X"ED",X"DD",X"7E",X"0B",X"E6",X"07",X"4F",X"5F",X"DD",X"36",X"0B",X"00",X"DD",X"CB",X"0B",X"FE",
		X"FD",X"CB",X"00",X"4E",X"20",X"2A",X"CD",X"67",X"0C",X"E6",X"0F",X"CB",X"D7",X"FD",X"77",X"01",
		X"FD",X"CB",X"00",X"CE",X"C5",X"CD",X"2A",X"26",X"21",X"1A",X"26",X"06",X"00",X"09",X"5E",X"C1",
		X"CD",X"67",X"0C",X"FE",X"64",X"38",X"09",X"E6",X"07",X"28",X"F5",X"FE",X"04",X"28",X"F1",X"5F",
		X"CD",X"AC",X"14",X"16",X"00",X"CB",X"23",X"21",X"C3",X"26",X"19",X"19",X"19",X"11",X"00",X"00",
		X"FD",X"36",X"04",X"00",X"FD",X"36",X"03",X"00",X"FD",X"36",X"0A",X"00",X"FD",X"36",X"09",X"00",
		X"78",X"A6",X"BE",X"28",X"0D",X"78",X"23",X"23",X"A6",X"BE",X"28",X"06",X"78",X"23",X"23",X"A6",
		X"BE",X"C0",X"23",X"7E",X"B9",X"20",X"04",X"DD",X"CB",X"0B",X"BE",X"5F",X"DD",X"7E",X"0B",X"E6",
		X"F8",X"B3",X"DD",X"77",X"0B",X"CB",X"23",X"CB",X"23",X"21",X"03",X"27",X"19",X"7E",X"FD",X"77",
		X"03",X"23",X"7E",X"FD",X"77",X"04",X"23",X"7E",X"FD",X"77",X"09",X"23",X"7E",X"FD",X"77",X"0A",
		X"DD",X"CB",X"0B",X"7E",X"C8",X"DD",X"CB",X"0B",X"BE",X"DD",X"4E",X"0B",X"06",X"00",X"21",X"F3",
		X"26",X"09",X"09",X"7E",X"23",X"66",X"6F",X"DD",X"CB",X"00",X"A6",X"DD",X"75",X"05",X"DD",X"74",
		X"06",X"DD",X"36",X"04",X"01",X"DD",X"CB",X"00",X"E6",X"C9",X"00",X"06",X"04",X"05",X"02",X"00",
		X"03",X"00",X"00",X"07",X"00",X"00",X"01",X"00",X"00",X"00",X"0E",X"00",X"3A",X"73",X"82",X"FD",
		X"BE",X"0C",X"38",X"04",X"CB",X"C9",X"18",X"04",X"28",X"02",X"CB",X"D9",X"3A",X"6D",X"82",X"FD",
		X"BE",X"06",X"38",X"03",X"CB",X"D1",X"C9",X"C8",X"CB",X"C1",X"C9",X"CB",X"77",X"28",X"08",X"01",
		X"02",X"02",X"CD",X"8B",X"1B",X"18",X"0A",X"CB",X"7F",X"28",X"06",X"01",X"02",X"02",X"CD",X"03",
		X"1C",X"3E",X"05",X"CD",X"45",X"0C",X"CD",X"69",X"1F",X"21",X"43",X"86",X"35",X"2B",X"7E",X"B7",
		X"28",X"04",X"35",X"C3",X"19",X"25",X"CD",X"68",X"0E",X"CD",X"EE",X"0D",X"18",X"FB",X"CD",X"67",
		X"0C",X"CB",X"6F",X"28",X"1F",X"FD",X"36",X"08",X"02",X"FD",X"36",X"0A",X"C8",X"21",X"40",X"27",
		X"FD",X"75",X"05",X"FD",X"74",X"06",X"FD",X"36",X"04",X"01",X"FD",X"CB",X"00",X"E6",X"3E",X"02",
		X"FD",X"77",X"0B",X"C9",X"FD",X"36",X"08",X"EE",X"FD",X"36",X"0A",X"C8",X"21",X"23",X"27",X"FD",
		X"75",X"05",X"FD",X"74",X"06",X"FD",X"36",X"04",X"01",X"FD",X"CB",X"00",X"E6",X"3E",X"06",X"FD",
		X"77",X"0B",X"C9",X"03",X"00",X"03",X"00",X"03",X"00",X"0F",X"01",X"0C",X"02",X"03",X"00",X"0C",
		X"02",X"0C",X"02",X"0C",X"02",X"3C",X"03",X"30",X"04",X"0C",X"02",X"30",X"04",X"30",X"04",X"30",
		X"04",X"F0",X"05",X"C0",X"06",X"30",X"04",X"C0",X"06",X"C0",X"06",X"C0",X"06",X"C3",X"07",X"03",
		X"00",X"C0",X"06",X"5D",X"27",X"B4",X"27",X"40",X"27",X"EE",X"27",X"7A",X"27",X"D1",X"27",X"23",
		X"27",X"97",X"27",X"00",X"00",X"00",X"FD",X"00",X"03",X"00",X"FD",X"00",X"03",X"00",X"00",X"00",
		X"03",X"00",X"03",X"00",X"00",X"00",X"03",X"00",X"FD",X"00",X"03",X"00",X"FD",X"00",X"00",X"00",
		X"FD",X"00",X"FD",X"00",X"00",X"01",X"00",X"00",X"0C",X"0C",X"05",X"6E",X"07",X"0C",X"0C",X"04",
		X"6F",X"07",X"0C",X"0C",X"05",X"70",X"07",X"0C",X"0C",X"04",X"6F",X"07",X"00",X"01",X"28",X"27",
		X"00",X"00",X"01",X"00",X"00",X"0C",X"0C",X"04",X"71",X"07",X"0C",X"0C",X"03",X"72",X"07",X"0C",
		X"0C",X"05",X"73",X"07",X"0C",X"0C",X"03",X"72",X"07",X"00",X"01",X"45",X"27",X"00",X"00",X"01",
		X"00",X"00",X"0C",X"0C",X"04",X"74",X"07",X"0C",X"0C",X"03",X"75",X"07",X"0C",X"0C",X"05",X"76",
		X"07",X"0C",X"0C",X"03",X"75",X"07",X"00",X"01",X"62",X"27",X"00",X"00",X"01",X"00",X"00",X"0C",
		X"0C",X"04",X"7D",X"07",X"0C",X"0C",X"03",X"7E",X"07",X"0C",X"0C",X"05",X"7F",X"07",X"0C",X"0C",
		X"03",X"1A",X"07",X"00",X"01",X"7F",X"27",X"00",X"00",X"01",X"00",X"00",X"0C",X"0C",X"05",X"74",
		X"07",X"0C",X"0C",X"04",X"75",X"07",X"0C",X"0C",X"05",X"76",X"07",X"0C",X"0C",X"04",X"75",X"07",
		X"00",X"01",X"9C",X"27",X"00",X"00",X"01",X"00",X"00",X"0C",X"0C",X"04",X"77",X"07",X"0C",X"0C",
		X"03",X"78",X"07",X"0C",X"0C",X"05",X"79",X"07",X"0C",X"0C",X"03",X"78",X"07",X"00",X"01",X"B9",
		X"27",X"00",X"00",X"01",X"00",X"00",X"0C",X"0C",X"04",X"7A",X"07",X"0C",X"0C",X"03",X"7B",X"07",
		X"0C",X"0C",X"05",X"7C",X"07",X"0C",X"0C",X"03",X"7B",X"07",X"00",X"01",X"D6",X"27",X"00",X"00",
		X"01",X"00",X"00",X"0C",X"0C",X"04",X"7D",X"07",X"0C",X"0C",X"03",X"7E",X"07",X"0C",X"0C",X"05",
		X"7F",X"07",X"0C",X"0C",X"03",X"7E",X"07",X"00",X"01",X"F3",X"27",X"3A",X"CA",X"81",X"B7",X"C8",
		X"FE",X"01",X"28",X"07",X"3A",X"30",X"86",X"CB",X"47",X"20",X"08",X"3A",X"32",X"86",X"CB",X"47",
		X"20",X"19",X"C9",X"AF",X"32",X"8C",X"86",X"CD",X"14",X"13",X"3E",X"02",X"32",X"67",X"86",X"21",
		X"47",X"86",X"CD",X"AA",X"29",X"CD",X"72",X"16",X"C3",X"47",X"28",X"AF",X"32",X"8C",X"86",X"AF",
		X"32",X"47",X"86",X"3C",X"32",X"67",X"86",X"3E",X"11",X"CD",X"45",X"0C",X"3E",X"01",X"CD",X"42",
		X"0E",X"3E",X"12",X"CD",X"45",X"0C",X"3E",X"01",X"CD",X"42",X"0E",X"CD",X"14",X"13",X"21",X"33",
		X"86",X"CD",X"AA",X"29",X"CD",X"72",X"16",X"CD",X"53",X"18",X"21",X"00",X"00",X"22",X"07",X"82",
		X"22",X"09",X"82",X"22",X"0B",X"82",X"22",X"C2",X"81",X"21",X"00",X"03",X"22",X"3A",X"86",X"21",
		X"00",X"03",X"22",X"4E",X"86",X"AF",X"32",X"66",X"86",X"3E",X"01",X"32",X"69",X"86",X"AF",X"32",
		X"7F",X"86",X"32",X"80",X"86",X"32",X"81",X"86",X"CD",X"88",X"29",X"CD",X"D5",X"29",X"3E",X"0A",
		X"CD",X"42",X"0E",X"CD",X"9B",X"0E",X"AF",X"CD",X"45",X"0C",X"3A",X"33",X"86",X"21",X"47",X"86",
		X"B6",X"20",X"E5",X"CD",X"ED",X"28",X"2A",X"80",X"86",X"ED",X"4B",X"82",X"86",X"09",X"22",X"82",
		X"86",X"2A",X"84",X"86",X"23",X"3A",X"67",X"86",X"FE",X"02",X"20",X"01",X"23",X"22",X"84",X"86",
		X"3E",X"01",X"32",X"8A",X"86",X"21",X"07",X"82",X"CD",X"C9",X"19",X"3E",X"02",X"32",X"8A",X"86",
		X"21",X"0A",X"82",X"CD",X"C9",X"19",X"AF",X"32",X"8A",X"86",X"C3",X"FD",X"17",X"3E",X"05",X"CD",
		X"42",X"0E",X"3E",X"00",X"32",X"3C",X"86",X"CF",X"28",X"68",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"00",X"CF",X"28",X"78",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"00",X"3A",X"67",X"86",X"FE",X"01",
		X"20",X"1C",X"CF",X"28",X"68",X"20",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"31",X"20",
		X"47",X"41",X"4D",X"45",X"20",X"4F",X"56",X"45",X"52",X"20",X"20",X"00",X"18",X"1D",X"CF",X"18",
		X"68",X"50",X"4C",X"41",X"59",X"45",X"52",X"53",X"20",X"31",X"20",X"41",X"4E",X"44",X"20",X"32",
		X"20",X"47",X"41",X"4D",X"45",X"20",X"4F",X"56",X"45",X"52",X"00",X"06",X"19",X"3E",X"FD",X"32",
		X"86",X"86",X"3E",X"03",X"CD",X"42",X"0E",X"10",X"F4",X"C9",X"3A",X"01",X"98",X"2F",X"E6",X"01",
		X"28",X"03",X"36",X"05",X"C9",X"36",X"03",X"C9",X"18",X"17",X"3A",X"69",X"86",X"FE",X"02",X"20",
		X"10",X"3A",X"02",X"98",X"E6",X"08",X"20",X"09",X"3E",X"FF",X"32",X"07",X"A8",X"32",X"06",X"A8",
		X"C9",X"3E",X"00",X"32",X"07",X"A8",X"32",X"06",X"A8",X"C9",X"CD",X"7A",X"29",X"23",X"36",X"00",
		X"23",X"36",X"00",X"23",X"36",X"0F",X"23",X"36",X"0F",X"23",X"36",X"01",X"23",X"36",X"02",X"21",
		X"3C",X"86",X"36",X"00",X"21",X"50",X"86",X"36",X"00",X"3E",X"00",X"32",X"8A",X"86",X"32",X"41",
		X"86",X"32",X"55",X"86",X"C9",X"3E",X"FF",X"32",X"A4",X"86",X"32",X"AA",X"86",X"AF",X"32",X"64",
		X"86",X"32",X"68",X"86",X"32",X"AB",X"86",X"3E",X"05",X"32",X"6A",X"86",X"CD",X"19",X"2B",X"CD",
		X"6B",X"15",X"CD",X"5A",X"4B",X"CD",X"07",X"17",X"3E",X"01",X"CD",X"42",X"0E",X"DD",X"21",X"EE",
		X"82",X"DD",X"7E",X"00",X"B7",X"20",X"F1",X"3A",X"33",X"86",X"FE",X"00",X"28",X"0A",X"FD",X"21",
		X"27",X"2D",X"CD",X"D6",X"0D",X"CD",X"C4",X"39",X"3A",X"67",X"86",X"FE",X"01",X"28",X"11",X"3A",
		X"47",X"86",X"FE",X"00",X"28",X"0A",X"FD",X"21",X"5D",X"2F",X"CD",X"D6",X"0D",X"CD",X"FA",X"39",
		X"FD",X"21",X"8E",X"39",X"CD",X"D6",X"0D",X"FD",X"21",X"9B",X"5D",X"CD",X"D6",X"0D",X"CD",X"1B",
		X"0B",X"3A",X"66",X"86",X"B7",X"28",X"44",X"CF",X"00",X"00",X"20",X"20",X"20",X"47",X"45",X"54",
		X"20",X"54",X"48",X"45",X"20",X"54",X"52",X"45",X"41",X"53",X"55",X"52",X"45",X"20",X"41",X"4E",
		X"44",X"20",X"42",X"52",X"49",X"4E",X"47",X"20",X"00",X"CF",X"00",X"08",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"49",X"54",X"20",X"54",X"4F",X"20",X"54",X"48",X"45",X"20",X"42",X"4F",
		X"41",X"54",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"00",X"3E",X"01",X"32",X"AB",X"86",
		X"CD",X"C8",X"0A",X"DD",X"21",X"EE",X"82",X"DD",X"7E",X"00",X"DD",X"21",X"1C",X"83",X"DD",X"B6",
		X"00",X"20",X"09",X"3E",X"00",X"32",X"8C",X"86",X"CD",X"16",X"5A",X"C9",X"3A",X"66",X"86",X"B7",
		X"C4",X"0B",X"28",X"3A",X"64",X"86",X"B7",X"C4",X"C8",X"0A",X"3A",X"68",X"86",X"FE",X"02",X"CA",
		X"D5",X"37",X"DD",X"21",X"EE",X"82",X"DD",X"7E",X"00",X"FE",X"00",X"20",X"19",X"3A",X"33",X"86",
		X"FE",X"00",X"28",X"12",X"3E",X"0A",X"CD",X"42",X"0E",X"FD",X"21",X"27",X"2D",X"CD",X"D6",X"0D",
		X"CD",X"C4",X"39",X"CD",X"1B",X"0B",X"3A",X"67",X"86",X"FE",X"01",X"28",X"24",X"DD",X"21",X"1C",
		X"83",X"DD",X"7E",X"00",X"FE",X"00",X"20",X"19",X"3A",X"47",X"86",X"FE",X"00",X"28",X"12",X"3E",
		X"0A",X"CD",X"42",X"0E",X"FD",X"21",X"5D",X"2F",X"CD",X"D6",X"0D",X"CD",X"FA",X"39",X"CD",X"1B",
		X"0B",X"3E",X"01",X"CD",X"42",X"0E",X"C3",X"8B",X"2A",X"3A",X"33",X"86",X"B7",X"20",X"04",X"32",
		X"AA",X"86",X"C9",X"3A",X"47",X"86",X"B7",X"C0",X"32",X"AA",X"86",X"C9",X"3A",X"8E",X"86",X"FE",
		X"19",X"D0",X"AF",X"32",X"A4",X"86",X"21",X"C0",X"2B",X"3A",X"38",X"86",X"BE",X"28",X"14",X"38",
		X"0C",X"3E",X"FF",X"BE",X"28",X"07",X"11",X"0B",X"00",X"19",X"C3",X"39",X"2B",X"11",X"0B",X"00",
		X"B7",X"ED",X"52",X"23",X"E5",X"7E",X"B7",X"28",X"14",X"47",X"C5",X"21",X"42",X"86",X"7E",X"B7",
		X"28",X"08",X"35",X"FD",X"21",X"F8",X"1D",X"CD",X"D6",X"0D",X"C1",X"10",X"ED",X"E1",X"23",X"E5",
		X"7E",X"B7",X"28",X"14",X"47",X"C5",X"21",X"42",X"86",X"7E",X"B7",X"28",X"08",X"35",X"FD",X"21",
		X"43",X"22",X"CD",X"D6",X"0D",X"C1",X"10",X"ED",X"E1",X"23",X"E5",X"7E",X"B7",X"28",X"14",X"47",
		X"C5",X"21",X"42",X"86",X"7E",X"B7",X"28",X"08",X"35",X"FD",X"21",X"0D",X"25",X"CD",X"D6",X"0D",
		X"C1",X"10",X"ED",X"E1",X"23",X"E5",X"7E",X"B7",X"28",X"14",X"47",X"C5",X"21",X"42",X"86",X"7E",
		X"B7",X"28",X"08",X"35",X"FD",X"21",X"B9",X"5A",X"CD",X"D6",X"0D",X"C1",X"10",X"ED",X"E1",X"C9",
		X"01",X"01",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"01",X"00",X"02",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"02",X"00",X"02",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"02",X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"01",X"00",X"04",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"03",X"00",X"03",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"03",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"01",X"00",
		X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"06",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0A",X"02",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"06",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",
		X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"06",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"12",X"06",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"13",X"01",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"14",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"01",X"00",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"16",X"01",X"00",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"17",X"01",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"01",X"00",
		X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"01",X"00",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"1A",X"01",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1B",X"01",
		X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"00",X"00",X"05",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"1D",X"01",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1E",
		X"01",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"01",X"00",X"04",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"01",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CF",X"10",X"00",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"00",X"CF",X"28",X"08",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"00",X"CD",
		X"AA",X"0C",X"3A",X"AB",X"86",X"B7",X"28",X"05",X"3E",X"5A",X"CD",X"42",X"0E",X"DD",X"21",X"EE",
		X"82",X"FD",X"21",X"67",X"82",X"21",X"34",X"86",X"36",X"00",X"21",X"35",X"86",X"36",X"00",X"CD",
		X"77",X"2E",X"DD",X"CB",X"00",X"D6",X"AF",X"DD",X"77",X"0D",X"DD",X"CB",X"0C",X"C6",X"DD",X"CB",
		X"00",X"F6",X"3E",X"05",X"FD",X"77",X"01",X"FD",X"CB",X"00",X"CE",X"CD",X"CC",X"2E",X"3E",X"01",
		X"CD",X"42",X"0E",X"3A",X"A4",X"86",X"B7",X"C4",X"2C",X"2B",X"FD",X"21",X"67",X"82",X"CD",X"93",
		X"31",X"DD",X"7E",X"08",X"FE",X"08",X"30",X"04",X"3E",X"E7",X"18",X"06",X"FE",X"E8",X"38",X"0A",
		X"3E",X"09",X"DD",X"77",X"08",X"3E",X"06",X"CD",X"45",X"0C",X"21",X"92",X"86",X"3A",X"91",X"86",
		X"B6",X"23",X"B6",X"23",X"B6",X"CA",X"24",X"2E",X"CD",X"86",X"59",X"21",X"89",X"86",X"7E",X"B7",
		X"28",X"01",X"35",X"DD",X"7E",X"0D",X"CB",X"57",X"C2",X"24",X"2E",X"CB",X"7F",X"C2",X"20",X"2E",
		X"FD",X"7E",X"0D",X"FE",X"A0",X"D2",X"24",X"2E",X"01",X"00",X"00",X"11",X"00",X"00",X"3A",X"66",
		X"86",X"B7",X"28",X"2F",X"3A",X"A6",X"86",X"FD",X"CB",X"00",X"56",X"20",X"49",X"3E",X"14",X"FD",
		X"77",X"02",X"FD",X"CB",X"00",X"D6",X"CD",X"67",X"0C",X"E6",X"3C",X"32",X"A6",X"86",X"18",X"36",
		X"AF",X"32",X"AA",X"86",X"3A",X"33",X"86",X"B7",X"28",X"06",X"C6",X"99",X"27",X"32",X"33",X"86",
		X"C3",X"78",X"32",X"3A",X"2F",X"86",X"E6",X"01",X"20",X"07",X"3A",X"2D",X"86",X"E6",X"3C",X"20",
		X"12",X"FD",X"36",X"04",X"00",X"FD",X"36",X"03",X"00",X"FD",X"36",X"0A",X"00",X"FD",X"36",X"09",
		X"00",X"18",X"09",X"3A",X"2D",X"86",X"E6",X"3C",X"67",X"CD",X"BF",X"31",X"3A",X"66",X"86",X"B7",
		X"28",X"05",X"CD",X"67",X"0C",X"18",X"03",X"3A",X"2F",X"86",X"E6",X"01",X"C4",X"99",X"2E",X"3E",
		X"01",X"CD",X"42",X"0E",X"C3",X"A3",X"2D",X"DD",X"36",X"08",X"91",X"DD",X"36",X"07",X"00",X"DD",
		X"36",X"0A",X"08",X"DD",X"36",X"09",X"00",X"21",X"B7",X"34",X"DD",X"75",X"05",X"DD",X"74",X"06",
		X"DD",X"36",X"04",X"01",X"DD",X"CB",X"00",X"E6",X"C9",X"3A",X"66",X"86",X"B7",X"20",X"06",X"3A",
		X"2D",X"86",X"E6",X"3C",X"C8",X"DD",X"CB",X"0C",X"4E",X"C0",X"3A",X"34",X"86",X"FE",X"03",X"C8",
		X"D0",X"3A",X"89",X"86",X"B7",X"C0",X"3E",X"03",X"32",X"89",X"86",X"FD",X"E5",X"FD",X"21",X"C5",
		X"35",X"CD",X"D6",X"0D",X"FD",X"E1",X"3E",X"04",X"CD",X"45",X"0C",X"C9",X"CD",X"86",X"59",X"3A",
		X"66",X"86",X"B7",X"28",X"05",X"CD",X"67",X"0C",X"18",X"03",X"3A",X"2D",X"86",X"E6",X"3C",X"06",
		X"01",X"C5",X"06",X"FF",X"26",X"04",X"CD",X"C4",X"31",X"CD",X"86",X"59",X"3E",X"01",X"CD",X"42",
		X"0E",X"FD",X"21",X"67",X"82",X"C1",X"10",X"E9",X"06",X"01",X"C5",X"06",X"FF",X"26",X"24",X"CD",
		X"C4",X"31",X"3E",X"01",X"CD",X"42",X"0E",X"CD",X"86",X"59",X"FD",X"21",X"67",X"82",X"C1",X"10",
		X"E9",X"06",X"06",X"C5",X"06",X"FF",X"26",X"20",X"CD",X"C4",X"31",X"3E",X"01",X"CD",X"42",X"0E",
		X"CD",X"86",X"59",X"FD",X"21",X"67",X"82",X"C1",X"10",X"E9",X"06",X"06",X"C5",X"06",X"FF",X"26",
		X"28",X"CD",X"C4",X"31",X"3E",X"01",X"CD",X"42",X"0E",X"CD",X"86",X"59",X"FD",X"21",X"67",X"82",
		X"C1",X"10",X"E9",X"06",X"0A",X"C5",X"06",X"FF",X"26",X"08",X"CD",X"C4",X"31",X"3E",X"01",X"CD",
		X"42",X"0E",X"CD",X"86",X"59",X"FD",X"21",X"67",X"82",X"C1",X"10",X"E9",X"C9",X"CF",X"10",X"00",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"00",X"CF",X"28",X"08",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"00",X"CD",X"CE",X"0C",X"3A",X"AB",X"86",X"B7",X"28",X"05",X"3E",X"5A",
		X"CD",X"42",X"0E",X"DD",X"21",X"1C",X"83",X"FD",X"21",X"76",X"82",X"21",X"48",X"86",X"36",X"00",
		X"21",X"49",X"86",X"36",X"00",X"CD",X"AD",X"30",X"DD",X"CB",X"00",X"D6",X"AF",X"DD",X"77",X"0D",
		X"DD",X"CB",X"0C",X"DE",X"DD",X"CB",X"00",X"F6",X"3E",X"05",X"FD",X"77",X"01",X"FD",X"CB",X"00",
		X"CE",X"CD",X"CF",X"30",X"3E",X"01",X"CD",X"42",X"0E",X"3A",X"A4",X"86",X"B7",X"C4",X"2C",X"2B",
		X"FD",X"21",X"76",X"82",X"CD",X"93",X"31",X"DD",X"7E",X"08",X"FE",X"08",X"30",X"04",X"3E",X"E7",
		X"18",X"06",X"FE",X"E8",X"38",X"0A",X"3E",X"09",X"DD",X"77",X"08",X"3E",X"06",X"CD",X"45",X"0C",
		X"21",X"96",X"86",X"3A",X"95",X"86",X"B6",X"23",X"B6",X"23",X"B6",X"CA",X"5A",X"30",X"CD",X"86",
		X"59",X"21",X"89",X"86",X"7E",X"B7",X"28",X"01",X"35",X"DD",X"7E",X"0D",X"CB",X"57",X"C2",X"5A",
		X"30",X"CB",X"77",X"C2",X"56",X"30",X"FD",X"7E",X"0D",X"FE",X"A0",X"D2",X"5A",X"30",X"01",X"00",
		X"00",X"11",X"00",X"00",X"3A",X"66",X"86",X"B7",X"28",X"2F",X"3A",X"A6",X"86",X"FD",X"CB",X"00",
		X"56",X"20",X"4B",X"3E",X"14",X"FD",X"77",X"02",X"FD",X"CB",X"00",X"D6",X"CD",X"67",X"0C",X"E6",
		X"3C",X"32",X"A6",X"86",X"18",X"38",X"AF",X"32",X"AA",X"86",X"3A",X"47",X"86",X"B7",X"28",X"06",
		X"C6",X"99",X"27",X"32",X"47",X"86",X"C3",X"78",X"32",X"3A",X"2D",X"86",X"E6",X"01",X"20",X"07",
		X"3A",X"2E",X"86",X"E6",X"3C",X"20",X"12",X"FD",X"36",X"04",X"00",X"FD",X"36",X"03",X"00",X"FD",
		X"36",X"0A",X"00",X"FD",X"36",X"09",X"00",X"18",X"09",X"3A",X"2E",X"86",X"E6",X"3C",X"67",X"CD",
		X"BF",X"31",X"3A",X"66",X"86",X"B7",X"28",X"05",X"CD",X"67",X"0C",X"18",X"03",X"3A",X"2D",X"86",
		X"E6",X"01",X"C4",X"60",X"31",X"3E",X"01",X"CD",X"42",X"0E",X"C3",X"D9",X"2F",X"DD",X"36",X"08",
		X"B9",X"DD",X"36",X"07",X"00",X"DD",X"36",X"0A",X"0A",X"DD",X"36",X"09",X"00",X"21",X"AD",X"35",
		X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",X"36",X"04",X"01",X"DD",X"CB",X"00",X"E6",X"C9",X"CD",
		X"86",X"59",X"3A",X"66",X"86",X"B7",X"28",X"05",X"CD",X"67",X"0C",X"18",X"03",X"3A",X"2E",X"86",
		X"E6",X"3C",X"06",X"01",X"C5",X"06",X"FF",X"26",X"04",X"CD",X"C4",X"31",X"CD",X"86",X"59",X"3E",
		X"01",X"CD",X"42",X"0E",X"FD",X"21",X"76",X"82",X"C1",X"10",X"E9",X"06",X"01",X"C5",X"06",X"FF",
		X"26",X"24",X"CD",X"C4",X"31",X"3E",X"01",X"CD",X"42",X"0E",X"CD",X"86",X"59",X"FD",X"21",X"76",
		X"82",X"C1",X"10",X"E9",X"06",X"06",X"C5",X"06",X"FF",X"26",X"20",X"CD",X"C4",X"31",X"3E",X"01",
		X"CD",X"42",X"0E",X"CD",X"86",X"59",X"FD",X"21",X"76",X"82",X"C1",X"10",X"E9",X"06",X"06",X"C5",
		X"06",X"FF",X"26",X"28",X"CD",X"C4",X"31",X"3E",X"01",X"CD",X"42",X"0E",X"CD",X"86",X"59",X"FD",
		X"21",X"76",X"82",X"C1",X"10",X"E9",X"06",X"0A",X"C5",X"06",X"FF",X"26",X"08",X"CD",X"C4",X"31",
		X"3E",X"01",X"CD",X"42",X"0E",X"CD",X"86",X"59",X"FD",X"21",X"76",X"82",X"C1",X"10",X"E9",X"C9",
		X"3A",X"66",X"86",X"B7",X"20",X"06",X"3A",X"2E",X"86",X"E6",X"3C",X"C8",X"DD",X"CB",X"0C",X"4E",
		X"C0",X"3A",X"48",X"86",X"FE",X"03",X"C8",X"D0",X"3A",X"89",X"86",X"B7",X"C0",X"3E",X"03",X"32",
		X"89",X"86",X"FD",X"E5",X"FD",X"21",X"D2",X"36",X"CD",X"D6",X"0D",X"FD",X"E1",X"3E",X"04",X"CD",
		X"45",X"0C",X"C9",X"DD",X"CB",X"0C",X"4E",X"C8",X"DD",X"7E",X"0A",X"FE",X"38",X"D0",X"DD",X"7E",
		X"08",X"FE",X"78",X"D8",X"FE",X"90",X"D0",X"3E",X"0E",X"CD",X"45",X"0C",X"3E",X"10",X"32",X"C5",
		X"89",X"32",X"C6",X"89",X"3E",X"02",X"32",X"68",X"86",X"3E",X"01",X"32",X"41",X"86",X"C9",X"E5",
		X"CD",X"AC",X"14",X"E1",X"FD",X"36",X"04",X"00",X"FD",X"36",X"03",X"00",X"FD",X"36",X"0A",X"00",
		X"FD",X"36",X"09",X"00",X"DD",X"7E",X"0B",X"E6",X"0F",X"4F",X"DD",X"36",X"0B",X"00",X"DD",X"CB",
		X"0B",X"FE",X"7C",X"1F",X"1F",X"E6",X"0F",X"C8",X"16",X"00",X"5F",X"CB",X"23",X"21",X"2F",X"33",
		X"19",X"19",X"19",X"11",X"00",X"00",X"78",X"A6",X"BE",X"28",X"0D",X"78",X"23",X"23",X"A6",X"BE",
		X"28",X"06",X"78",X"23",X"23",X"A6",X"BE",X"C0",X"23",X"7E",X"1C",X"1F",X"30",X"FC",X"7B",X"B9",
		X"20",X"04",X"DD",X"CB",X"0B",X"BE",X"DD",X"7E",X"0B",X"E6",X"F0",X"B3",X"DD",X"77",X"0B",X"1D",
		X"DD",X"CB",X"0C",X"4E",X"28",X"05",X"21",X"AF",X"33",X"18",X"03",X"21",X"8F",X"33",X"19",X"19",
		X"19",X"19",X"7E",X"FD",X"77",X"03",X"23",X"7E",X"FD",X"77",X"04",X"23",X"7E",X"FD",X"77",X"09",
		X"23",X"7E",X"FD",X"77",X"0A",X"DD",X"CB",X"0B",X"7E",X"C8",X"DD",X"CB",X"0B",X"BE",X"DD",X"4E",
		X"0B",X"06",X"00",X"21",X"0B",X"33",X"DD",X"CB",X"0C",X"46",X"20",X"03",X"21",X"1D",X"33",X"09",
		X"09",X"7E",X"23",X"66",X"6F",X"DD",X"CB",X"00",X"A6",X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",
		X"36",X"04",X"01",X"DD",X"CB",X"00",X"E6",X"C9",X"3E",X"02",X"32",X"41",X"86",X"DD",X"CB",X"0C",
		X"86",X"3E",X"05",X"CD",X"45",X"0C",X"AF",X"FD",X"77",X"03",X"FD",X"77",X"04",X"FD",X"77",X"09",
		X"FD",X"77",X"0A",X"DD",X"CB",X"00",X"B6",X"DD",X"CB",X"00",X"A6",X"21",X"4A",X"21",X"DD",X"75",
		X"05",X"DD",X"74",X"06",X"DD",X"36",X"04",X"01",X"DD",X"CB",X"00",X"E6",X"DD",X"CB",X"00",X"66",
		X"28",X"05",X"CD",X"EE",X"0D",X"18",X"F5",X"AF",X"DD",X"77",X"08",X"DD",X"77",X"0A",X"CD",X"68",
		X"0E",X"CD",X"EE",X"0D",X"18",X"FB",X"00",X"00",X"01",X"00",X"00",X"01",X"00",X"03",X"1B",X"02",
		X"01",X"00",X"03",X"9B",X"03",X"01",X"00",X"03",X"1A",X"04",X"01",X"00",X"03",X"9A",X"05",X"01",
		X"00",X"03",X"19",X"06",X"01",X"00",X"03",X"99",X"07",X"01",X"00",X"03",X"17",X"02",X"01",X"00",
		X"03",X"97",X"03",X"01",X"00",X"03",X"16",X"04",X"01",X"00",X"03",X"96",X"05",X"01",X"00",X"03",
		X"12",X"06",X"01",X"00",X"03",X"92",X"07",X"00",X"00",X"00",X"00",X"B7",X"34",X"60",X"34",X"7D",
		X"34",X"CF",X"33",X"43",X"34",X"09",X"34",X"26",X"34",X"EC",X"33",X"9A",X"34",X"AD",X"35",X"56",
		X"35",X"73",X"35",X"C5",X"34",X"39",X"35",X"FF",X"34",X"1C",X"35",X"E2",X"34",X"90",X"35",X"3C",
		X"08",X"30",X"10",X"0C",X"04",X"03",X"01",X"03",X"01",X"03",X"01",X"30",X"10",X"30",X"10",X"30",
		X"10",X"3C",X"08",X"30",X"10",X"0C",X"04",X"0C",X"04",X"0C",X"04",X"0C",X"04",X"0F",X"02",X"0C",
		X"04",X"03",X"01",X"3C",X"08",X"30",X"10",X"0C",X"04",X"F0",X"20",X"C0",X"40",X"30",X"10",X"C0",
		X"40",X"C0",X"40",X"C0",X"40",X"C3",X"80",X"03",X"01",X"C0",X"40",X"F0",X"20",X"C0",X"40",X"30",
		X"10",X"3C",X"08",X"30",X"10",X"0C",X"04",X"F0",X"20",X"C0",X"40",X"30",X"10",X"F0",X"20",X"C0",
		X"40",X"30",X"10",X"3C",X"08",X"30",X"10",X"0C",X"04",X"F0",X"20",X"C0",X"40",X"30",X"10",X"00",
		X"00",X"80",X"FD",X"80",X"02",X"80",X"FD",X"80",X"02",X"00",X"00",X"80",X"02",X"80",X"02",X"00",
		X"00",X"80",X"02",X"80",X"FD",X"80",X"02",X"80",X"FD",X"00",X"00",X"80",X"FD",X"80",X"FD",X"00",
		X"00",X"D0",X"FE",X"00",X"01",X"00",X"FF",X"00",X"02",X"00",X"00",X"00",X"03",X"00",X"03",X"00",
		X"00",X"00",X"03",X"00",X"FD",X"00",X"03",X"00",X"FE",X"00",X"00",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"01",X"00",X"00",X"06",X"06",X"03",X"40",X"07",X"06",X"06",X"03",X"41",X"07",X"06",X"06",
		X"03",X"42",X"07",X"06",X"06",X"03",X"41",X"07",X"00",X"01",X"D4",X"33",X"00",X"00",X"01",X"00",
		X"00",X"06",X"06",X"03",X"43",X"07",X"06",X"06",X"03",X"45",X"07",X"06",X"06",X"03",X"46",X"07",
		X"06",X"06",X"03",X"45",X"07",X"00",X"01",X"F1",X"33",X"00",X"00",X"01",X"00",X"00",X"06",X"06",
		X"03",X"47",X"07",X"06",X"06",X"03",X"48",X"07",X"06",X"06",X"03",X"49",X"07",X"06",X"06",X"03",
		X"48",X"07",X"00",X"01",X"0E",X"34",X"00",X"00",X"01",X"00",X"00",X"06",X"06",X"03",X"53",X"07",
		X"06",X"06",X"03",X"54",X"07",X"06",X"06",X"03",X"55",X"07",X"06",X"06",X"03",X"54",X"07",X"00",
		X"01",X"2B",X"34",X"00",X"00",X"01",X"00",X"00",X"06",X"06",X"03",X"56",X"07",X"06",X"06",X"03",
		X"57",X"07",X"06",X"06",X"03",X"58",X"07",X"06",X"06",X"03",X"57",X"07",X"00",X"01",X"48",X"34",
		X"00",X"00",X"01",X"00",X"00",X"06",X"06",X"03",X"4A",X"07",X"06",X"06",X"03",X"4B",X"07",X"06",
		X"06",X"03",X"4C",X"07",X"06",X"06",X"03",X"4B",X"07",X"00",X"01",X"65",X"34",X"00",X"00",X"01",
		X"00",X"00",X"06",X"06",X"03",X"4D",X"07",X"06",X"06",X"03",X"4E",X"07",X"06",X"06",X"03",X"4F",
		X"07",X"06",X"06",X"03",X"4E",X"07",X"00",X"01",X"82",X"34",X"00",X"00",X"01",X"00",X"00",X"06",
		X"06",X"03",X"50",X"07",X"06",X"06",X"03",X"51",X"07",X"06",X"06",X"03",X"52",X"07",X"06",X"06",
		X"03",X"51",X"07",X"00",X"01",X"9F",X"34",X"00",X"00",X"01",X"00",X"00",X"06",X"04",X"01",X"4A",
		X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"06",X"06",X"03",X"40",X"02",X"06",
		X"06",X"03",X"41",X"02",X"06",X"06",X"03",X"42",X"02",X"06",X"06",X"03",X"41",X"02",X"00",X"01",
		X"CA",X"34",X"00",X"00",X"01",X"00",X"00",X"06",X"06",X"03",X"43",X"02",X"06",X"06",X"03",X"45",
		X"02",X"06",X"06",X"03",X"46",X"02",X"06",X"06",X"03",X"45",X"02",X"00",X"01",X"E7",X"34",X"00",
		X"00",X"01",X"00",X"00",X"06",X"06",X"03",X"47",X"02",X"06",X"06",X"03",X"48",X"02",X"06",X"06",
		X"03",X"49",X"02",X"06",X"06",X"03",X"48",X"02",X"00",X"01",X"04",X"35",X"00",X"00",X"01",X"00",
		X"00",X"06",X"06",X"03",X"53",X"02",X"06",X"06",X"03",X"54",X"02",X"06",X"06",X"03",X"55",X"02",
		X"06",X"06",X"03",X"54",X"02",X"00",X"01",X"21",X"35",X"00",X"00",X"01",X"00",X"00",X"06",X"06",
		X"03",X"56",X"02",X"06",X"06",X"03",X"57",X"02",X"06",X"06",X"03",X"58",X"02",X"06",X"06",X"03",
		X"57",X"02",X"00",X"01",X"3E",X"35",X"00",X"00",X"01",X"00",X"00",X"06",X"06",X"03",X"4A",X"02",
		X"06",X"06",X"03",X"4B",X"02",X"06",X"06",X"03",X"4C",X"02",X"06",X"06",X"03",X"4B",X"02",X"00",
		X"01",X"5B",X"35",X"00",X"00",X"01",X"00",X"00",X"06",X"06",X"03",X"4D",X"02",X"06",X"06",X"03",
		X"4E",X"02",X"06",X"06",X"03",X"4F",X"02",X"06",X"06",X"03",X"4E",X"02",X"00",X"01",X"78",X"35",
		X"00",X"00",X"01",X"00",X"00",X"06",X"06",X"03",X"50",X"02",X"06",X"06",X"03",X"51",X"02",X"06",
		X"06",X"03",X"52",X"02",X"06",X"06",X"03",X"51",X"02",X"00",X"01",X"95",X"35",X"00",X"00",X"01",
		X"00",X"00",X"06",X"04",X"01",X"4A",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",
		X"04",X"04",X"00",X"00",X"00",X"CD",X"14",X"0D",X"D2",X"1B",X"36",X"DD",X"E5",X"FD",X"E1",X"DD",
		X"2A",X"B6",X"81",X"21",X"34",X"86",X"34",X"CD",X"27",X"36",X"CD",X"55",X"36",X"DD",X"CB",X"0C",
		X"F6",X"21",X"BB",X"35",X"DD",X"75",X"05",X"DD",X"74",X"06",X"3E",X"0F",X"DD",X"77",X"03",X"DD",
		X"CB",X"00",X"EE",X"DD",X"36",X"0D",X"00",X"DD",X"CB",X"00",X"D6",X"DD",X"CB",X"00",X"F6",X"FD",
		X"E5",X"CD",X"EE",X"0D",X"FD",X"E1",X"DD",X"7E",X"0D",X"CB",X"87",X"B7",X"20",X"0D",X"DD",X"CB",
		X"00",X"6E",X"28",X"07",X"FD",X"E5",X"CD",X"EE",X"0D",X"18",X"E9",X"21",X"34",X"86",X"35",X"CD",
		X"68",X"0E",X"CD",X"EE",X"0D",X"18",X"FB",X"FD",X"E5",X"FD",X"21",X"EE",X"82",X"FD",X"46",X"08",
		X"05",X"05",X"CD",X"67",X"0C",X"E6",X"07",X"FE",X"06",X"30",X"F7",X"80",X"DD",X"77",X"08",X"FD",
		X"46",X"0A",X"05",X"05",X"05",X"CD",X"67",X"0C",X"E6",X"07",X"FE",X"06",X"30",X"F7",X"80",X"DD",
		X"77",X"0A",X"FD",X"E1",X"C9",X"3A",X"66",X"86",X"B7",X"28",X"05",X"CD",X"67",X"0C",X"18",X"03",
		X"3A",X"2D",X"86",X"E6",X"3C",X"C8",X"CB",X"3F",X"CB",X"3F",X"5F",X"16",X"00",X"21",X"88",X"36",
		X"19",X"19",X"19",X"19",X"5E",X"23",X"56",X"23",X"4E",X"23",X"46",X"FD",X"73",X"03",X"FD",X"72",
		X"04",X"FD",X"71",X"09",X"FD",X"70",X"0A",X"C9",X"EE",X"FA",X"EE",X"FA",X"00",X"00",X"5E",X"F9",
		X"00",X"00",X"A2",X"06",X"A2",X"06",X"00",X"00",X"A2",X"06",X"00",X"00",X"12",X"05",X"EE",X"FA",
		X"12",X"05",X"12",X"05",X"EE",X"FA",X"EE",X"FA",X"5E",X"F9",X"00",X"00",X"EE",X"FA",X"EE",X"FA",
		X"EE",X"FA",X"12",X"05",X"12",X"05",X"EE",X"FA",X"12",X"05",X"12",X"05",X"EE",X"FA",X"EE",X"FA",
		X"5E",X"F9",X"00",X"00",X"EE",X"FA",X"EE",X"FA",X"00",X"00",X"01",X"00",X"00",X"04",X"04",X"00",
		X"00",X"00",X"CD",X"32",X"0D",X"D2",X"28",X"37",X"DD",X"E5",X"FD",X"E1",X"DD",X"2A",X"B6",X"81",
		X"21",X"48",X"86",X"34",X"CD",X"34",X"37",X"CD",X"62",X"37",X"DD",X"CB",X"0C",X"FE",X"21",X"C8",
		X"36",X"DD",X"75",X"05",X"DD",X"74",X"06",X"3E",X"0F",X"DD",X"77",X"03",X"DD",X"CB",X"00",X"EE",
		X"DD",X"36",X"0D",X"00",X"DD",X"CB",X"00",X"D6",X"DD",X"CB",X"00",X"F6",X"FD",X"E5",X"CD",X"EE",
		X"0D",X"FD",X"E1",X"DD",X"7E",X"0D",X"CB",X"9F",X"B7",X"20",X"0D",X"DD",X"CB",X"00",X"6E",X"28",
		X"07",X"FD",X"E5",X"CD",X"EE",X"0D",X"18",X"E9",X"21",X"48",X"86",X"35",X"CD",X"68",X"0E",X"CD",
		X"EE",X"0D",X"18",X"FB",X"FD",X"E5",X"FD",X"21",X"1C",X"83",X"FD",X"46",X"08",X"05",X"05",X"CD",
		X"67",X"0C",X"E6",X"07",X"FE",X"06",X"30",X"F7",X"80",X"DD",X"77",X"08",X"FD",X"46",X"0A",X"05",
		X"05",X"05",X"CD",X"67",X"0C",X"E6",X"07",X"FE",X"06",X"30",X"F7",X"80",X"DD",X"77",X"0A",X"FD",
		X"E1",X"C9",X"3A",X"66",X"86",X"B7",X"28",X"05",X"CD",X"67",X"0C",X"18",X"03",X"3A",X"2E",X"86",
		X"E6",X"3C",X"C8",X"CB",X"3F",X"CB",X"3F",X"5F",X"16",X"00",X"21",X"95",X"37",X"19",X"19",X"19",
		X"19",X"5E",X"23",X"56",X"23",X"4E",X"23",X"46",X"FD",X"73",X"03",X"FD",X"72",X"04",X"FD",X"71",
		X"09",X"FD",X"70",X"0A",X"C9",X"EE",X"FA",X"EE",X"FA",X"00",X"00",X"5E",X"F9",X"00",X"00",X"A2",
		X"06",X"A2",X"06",X"00",X"00",X"A2",X"06",X"00",X"00",X"12",X"05",X"EE",X"FA",X"12",X"05",X"12",
		X"05",X"EE",X"FA",X"EE",X"FA",X"5E",X"F9",X"00",X"00",X"EE",X"FA",X"EE",X"FA",X"EE",X"FA",X"12",
		X"05",X"12",X"05",X"EE",X"FA",X"12",X"05",X"12",X"05",X"EE",X"FA",X"EE",X"FA",X"5E",X"F9",X"00",
		X"00",X"EE",X"FA",X"EE",X"FA",X"AF",X"32",X"8C",X"86",X"CD",X"9B",X"0E",X"3E",X"00",X"CD",X"45",
		X"0C",X"3E",X"01",X"CD",X"42",X"0E",X"3E",X"10",X"CD",X"45",X"0C",X"3E",X"01",X"CD",X"42",X"0E",
		X"21",X"38",X"86",X"34",X"CD",X"72",X"16",X"3E",X"00",X"32",X"68",X"86",X"CD",X"C8",X"0A",X"CD",
		X"1B",X"0B",X"21",X"78",X"18",X"01",X"08",X"1A",X"CD",X"01",X"0A",X"3A",X"67",X"86",X"FE",X"02",
		X"CA",X"A4",X"38",X"CF",X"40",X"88",X"59",X"4F",X"55",X"52",X"20",X"4F",X"4C",X"44",X"20",X"53",
		X"43",X"4F",X"52",X"45",X"00",X"21",X"88",X"B0",X"11",X"07",X"82",X"06",X"06",X"CD",X"66",X"09",
		X"CF",X"40",X"98",X"59",X"4F",X"55",X"52",X"20",X"41",X"49",X"52",X"20",X"42",X"4F",X"4E",X"55",
		X"53",X"00",X"21",X"93",X"88",X"CD",X"A7",X"3A",X"3A",X"94",X"86",X"4F",X"06",X"03",X"CD",X"8B",
		X"1B",X"3E",X"01",X"CD",X"42",X"0E",X"3A",X"93",X"86",X"4F",X"06",X"02",X"CD",X"8B",X"1B",X"3E",
		X"01",X"CD",X"42",X"0E",X"3A",X"92",X"86",X"4F",X"06",X"01",X"CD",X"8B",X"1B",X"3E",X"01",X"CD",
		X"42",X"0E",X"3A",X"91",X"86",X"4F",X"06",X"00",X"CD",X"8B",X"1B",X"3E",X"01",X"CD",X"42",X"0E",
		X"CF",X"20",X"A8",X"59",X"4F",X"55",X"52",X"20",X"43",X"55",X"52",X"52",X"45",X"4E",X"54",X"20",
		X"53",X"43",X"4F",X"52",X"45",X"00",X"21",X"A8",X"B0",X"11",X"07",X"82",X"06",X"06",X"CD",X"66",
		X"09",X"C3",X"7B",X"39",X"3A",X"94",X"86",X"4F",X"06",X"03",X"CD",X"8B",X"1B",X"3E",X"01",X"CD",
		X"42",X"0E",X"3A",X"93",X"86",X"4F",X"06",X"02",X"CD",X"8B",X"1B",X"3E",X"01",X"CD",X"42",X"0E",
		X"3A",X"92",X"86",X"4F",X"06",X"01",X"CD",X"8B",X"1B",X"3E",X"01",X"CD",X"42",X"0E",X"3A",X"91",
		X"86",X"4F",X"06",X"00",X"CD",X"8B",X"1B",X"3E",X"01",X"CD",X"42",X"0E",X"3A",X"98",X"86",X"4F",
		X"06",X"03",X"CD",X"03",X"1C",X"3E",X"01",X"CD",X"42",X"0E",X"3A",X"97",X"86",X"4F",X"06",X"02",
		X"CD",X"03",X"1C",X"3E",X"01",X"CD",X"42",X"0E",X"3A",X"96",X"86",X"4F",X"06",X"01",X"CD",X"03",
		X"1C",X"3E",X"01",X"CD",X"42",X"0E",X"3A",X"95",X"86",X"4F",X"06",X"00",X"CD",X"03",X"1C",X"3E",
		X"01",X"CD",X"42",X"0E",X"CF",X"30",X"98",X"20",X"42",X"55",X"44",X"44",X"59",X"20",X"53",X"59",
		X"53",X"54",X"45",X"4D",X"20",X"42",X"4F",X"4E",X"55",X"53",X"20",X"00",X"3A",X"AA",X"86",X"B7",
		X"20",X"19",X"CF",X"30",X"A8",X"30",X"30",X"30",X"20",X"20",X"46",X"4F",X"52",X"20",X"45",X"41",
		X"43",X"48",X"20",X"44",X"49",X"56",X"45",X"52",X"00",X"18",X"30",X"CF",X"30",X"A8",X"32",X"30",
		X"30",X"30",X"20",X"20",X"46",X"4F",X"52",X"20",X"45",X"41",X"43",X"48",X"20",X"44",X"49",X"56",
		X"45",X"52",X"00",X"0E",X"02",X"06",X"03",X"CD",X"8B",X"1B",X"3E",X"01",X"CD",X"42",X"0E",X"0E",
		X"02",X"06",X"03",X"CD",X"03",X"1C",X"3E",X"01",X"CD",X"42",X"0E",X"3E",X"04",X"CD",X"42",X"0E",
		X"CD",X"C8",X"0A",X"3E",X"32",X"CD",X"42",X"0E",X"CD",X"9B",X"0E",X"C3",X"D5",X"29",X"CD",X"50",
		X"0D",X"D2",X"12",X"0E",X"DD",X"E5",X"DD",X"21",X"EE",X"82",X"DD",X"7E",X"00",X"B7",X"28",X"03",
		X"CD",X"57",X"3A",X"3A",X"67",X"86",X"FE",X"01",X"28",X"0D",X"DD",X"21",X"1C",X"83",X"DD",X"7E",
		X"00",X"B7",X"28",X"03",X"CD",X"BE",X"3A",X"DD",X"E1",X"CD",X"EE",X"0D",X"3E",X"01",X"CD",X"42",
		X"0E",X"C3",X"94",X"39",X"3A",X"38",X"86",X"FE",X"0A",X"38",X"02",X"3E",X"0A",X"CB",X"27",X"21",
		X"2E",X"3A",X"06",X"00",X"4F",X"09",X"56",X"23",X"5E",X"3A",X"2C",X"86",X"CB",X"5F",X"28",X"0A",
		X"1C",X"1C",X"3E",X"09",X"BB",X"30",X"03",X"1E",X"00",X"14",X"7A",X"32",X"94",X"86",X"7B",X"32",
		X"93",X"86",X"AF",X"32",X"92",X"86",X"32",X"91",X"86",X"C9",X"3A",X"38",X"86",X"FE",X"0A",X"38",
		X"02",X"3E",X"0A",X"CB",X"27",X"21",X"2E",X"3A",X"06",X"00",X"4F",X"09",X"56",X"23",X"5E",X"3A",
		X"2C",X"86",X"CB",X"5F",X"28",X"0A",X"1C",X"1C",X"3E",X"09",X"BB",X"30",X"03",X"1E",X"00",X"14",
		X"7A",X"32",X"98",X"86",X"7B",X"32",X"97",X"86",X"AF",X"32",X"96",X"86",X"32",X"95",X"86",X"C9",
		X"00",X"08",X"00",X"08",X"00",X"09",X"00",X"09",X"01",X"00",X"01",X"00",X"01",X"01",X"01",X"01",
		X"01",X"02",X"01",X"02",X"01",X"04",X"01",X"04",X"AF",X"32",X"91",X"86",X"32",X"95",X"86",X"32",
		X"92",X"86",X"32",X"96",X"86",X"18",X"49",X"3A",X"91",X"86",X"3D",X"32",X"91",X"86",X"FE",X"FF",
		X"20",X"3E",X"3E",X"09",X"32",X"91",X"86",X"3A",X"92",X"86",X"3D",X"32",X"92",X"86",X"FE",X"FF",
		X"20",X"2E",X"3E",X"09",X"32",X"92",X"86",X"3A",X"93",X"86",X"3D",X"32",X"93",X"86",X"FE",X"FF",
		X"20",X"1E",X"3E",X"09",X"32",X"93",X"86",X"3A",X"94",X"86",X"3D",X"32",X"94",X"86",X"FE",X"FF",
		X"20",X"0E",X"3E",X"00",X"32",X"91",X"86",X"32",X"92",X"86",X"32",X"93",X"86",X"32",X"94",X"86",
		X"21",X"7F",X"88",X"11",X"40",X"02",X"19",X"11",X"20",X"00",X"3A",X"91",X"86",X"77",X"19",X"3A",
		X"92",X"86",X"77",X"19",X"3A",X"93",X"86",X"77",X"19",X"3A",X"94",X"86",X"77",X"C9",X"3A",X"95",
		X"86",X"3D",X"32",X"95",X"86",X"FE",X"FF",X"20",X"3E",X"3E",X"09",X"32",X"95",X"86",X"3A",X"96",
		X"86",X"3D",X"32",X"96",X"86",X"FE",X"FF",X"20",X"2E",X"3E",X"09",X"32",X"96",X"86",X"3A",X"97",
		X"86",X"3D",X"32",X"97",X"86",X"FE",X"FF",X"20",X"1E",X"3E",X"09",X"32",X"97",X"86",X"3A",X"98",
		X"86",X"3D",X"32",X"98",X"86",X"FE",X"FF",X"20",X"0E",X"3E",X"00",X"32",X"95",X"86",X"32",X"96",
		X"86",X"32",X"97",X"86",X"32",X"98",X"86",X"21",X"7F",X"88",X"11",X"20",X"00",X"3A",X"95",X"86",
		X"77",X"19",X"3A",X"96",X"86",X"77",X"19",X"3A",X"97",X"86",X"77",X"19",X"3A",X"98",X"86",X"77",
		X"C9",X"17",X"46",X"56",X"5A",X"3E",X"1A",X"48",X"9A",X"41",X"DA",X"44",X"86",X"4C",X"C6",X"4F",
		X"06",X"53",X"34",X"3B",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"5F",X"60",X"60",X"60",X"60",X"60",X"62",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"63",X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"5E",X"10",X"10",X"10",X"10",X"10",
		X"61",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"5F",X"60",
		X"60",X"5C",X"60",X"60",X"60",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"63",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"5E",X"60",X"60",X"5D",X"60",X"60",X"60",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"60",X"10",X"60",X"60",X"60",X"60",X"60",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"5F",X"60",X"60",X"60",X"60",X"60",X"5C",X"60",X"60",X"60",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",
		X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"5E",X"60",X"60",X"60",X"60",X"60",X"61",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"5F",X"60",X"60",X"62",X"10",X"10",
		X"62",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"63",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"5E",X"10",
		X"10",X"5E",X"60",X"60",X"61",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"5F",X"60",X"60",X"60",X"60",X"60",X"62",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",
		X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"5E",X"60",X"60",X"60",X"60",X"60",X"61",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",
		X"8F",X"9F",X"9E",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",
		X"8F",X"9C",X"9D",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"10",X"10",X"8F",X"8F",X"8F",
		X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"10",X"10",X"8F",X"8F",X"8F",X"8F",X"9C",X"9E",
		X"9F",X"9D",X"9E",X"9F",X"9D",X"10",X"10",X"9C",X"9F",X"9C",X"9D",X"9E",X"9F",X"9C",X"9E",X"9D",
		X"9F",X"9C",X"10",X"10",X"9F",X"9D",X"9C",X"8F",X"10",X"10",X"10",X"8D",X"10",X"10",X"8F",X"10",
		X"10",X"8E",X"10",X"10",X"8F",X"10",X"10",X"10",X"8D",X"10",X"10",X"8D",X"10",X"10",X"8F",X"10",
		X"10",X"8F",X"10",X"10",X"10",X"8E",X"10",X"10",X"8E",X"10",X"10",X"8D",X"10",X"10",X"90",X"10",
		X"10",X"10",X"90",X"10",X"10",X"8E",X"10",X"10",X"8E",X"10",X"10",X"8F",X"10",X"10",X"10",X"8E",
		X"10",X"10",X"8D",X"10",X"10",X"90",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"8D",
		X"10",X"10",X"90",X"10",X"10",X"8F",X"10",X"10",X"10",X"8F",X"10",X"10",X"8F",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"8F",X"10",X"10",X"10",X"10",X"10",X"8F",
		X"10",X"10",X"10",X"8E",X"10",X"10",X"8E",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"8E",X"10",X"10",X"10",X"10",X"10",X"8F",X"10",X"10",X"10",X"8F",X"10",X"10",
		X"8F",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"8D",X"10",X"10",
		X"10",X"10",X"10",X"8F",X"10",X"10",X"10",X"8E",X"10",X"10",X"8E",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"8E",X"10",X"10",X"10",X"10",X"10",X"8F",X"10",X"10",
		X"10",X"8D",X"10",X"10",X"8F",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"8F",X"10",X"10",X"10",X"10",X"10",X"8F",X"10",X"10",X"10",X"8F",X"10",X"10",X"8E",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"8E",X"10",X"10",X"10",X"10",
		X"10",X"8F",X"10",X"10",X"10",X"90",X"10",X"10",X"8F",X"10",X"10",X"10",X"10",X"10",X"91",X"10",
		X"10",X"10",X"10",X"10",X"10",X"90",X"10",X"10",X"10",X"10",X"10",X"8F",X"10",X"10",X"10",X"10",
		X"10",X"10",X"8D",X"10",X"10",X"10",X"10",X"10",X"8E",X"10",X"10",X"10",X"91",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"8F",X"10",X"10",X"10",X"10",X"10",X"10",X"8E",X"10",X"10",X"10",
		X"10",X"10",X"8F",X"10",X"10",X"10",X"8E",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"8F",
		X"10",X"10",X"10",X"10",X"10",X"10",X"8F",X"10",X"10",X"10",X"10",X"10",X"8E",X"10",X"10",X"10",
		X"8F",X"10",X"10",X"10",X"10",X"10",X"91",X"10",X"10",X"8F",X"10",X"10",X"10",X"10",X"10",X"10",
		X"90",X"10",X"10",X"10",X"10",X"10",X"8F",X"10",X"10",X"10",X"8E",X"10",X"10",X"10",X"10",X"10",
		X"8E",X"10",X"10",X"8F",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"8E",X"10",X"10",X"10",X"8F",X"10",X"10",X"10",X"10",X"10",X"8F",X"10",X"10",X"8F",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"8F",X"10",X"10",X"10",X"8E",X"10",
		X"10",X"10",X"10",X"10",X"8D",X"10",X"10",X"8F",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"8E",X"10",X"10",X"10",X"8F",X"10",X"10",X"10",X"10",X"10",X"8F",X"10",
		X"10",X"8F",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"8F",X"10",
		X"10",X"10",X"8E",X"10",X"10",X"10",X"10",X"10",X"8E",X"10",X"10",X"8F",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"8E",X"10",X"10",X"10",X"8F",X"10",X"10",X"10",
		X"10",X"10",X"8F",X"10",X"10",X"8F",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"8F",X"10",X"10",X"10",X"90",X"10",X"10",X"10",X"10",X"10",X"8E",X"10",X"10",X"8F",
		X"10",X"10",X"10",X"10",X"10",X"91",X"10",X"10",X"10",X"10",X"10",X"10",X"8E",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"90",X"10",X"10",X"8F",X"10",X"10",X"10",X"10",X"10",X"9F",
		X"10",X"10",X"10",X"10",X"10",X"10",X"8D",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"8F",X"10",X"10",X"10",X"10",X"10",X"8E",X"10",X"10",X"10",X"10",X"10",X"10",
		X"8F",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"8F",X"10",X"10",
		X"10",X"10",X"10",X"8D",X"10",X"10",X"10",X"10",X"10",X"10",X"8E",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"8F",X"10",X"10",X"91",X"10",X"10",X"8E",X"10",X"10",
		X"10",X"10",X"10",X"10",X"8F",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"8F",X"10",X"10",X"8F",X"10",X"10",X"8F",X"10",X"10",X"10",X"10",X"10",X"10",X"8D",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"8F",X"9C",X"98",X"8F",X"9A",
		X"98",X"8F",X"98",X"10",X"10",X"9B",X"99",X"98",X"8F",X"9B",X"98",X"9A",X"8F",X"9B",X"9A",X"8F",
		X"10",X"10",X"8F",X"99",X"9B",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"10",X"10",X"8F",
		X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"10",X"10",X"8F",X"8F",X"8F",X"8F",
		X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"99",X"98",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",
		X"8F",X"8F",X"8F",X"8F",X"9A",X"9B",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",
		X"8F",X"72",X"71",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",
		X"8F",X"71",X"73",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"10",X"10",X"8F",X"8F",X"8F",
		X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"10",X"10",X"8F",X"8F",X"8F",X"69",X"71",X"72",
		X"70",X"72",X"70",X"72",X"70",X"10",X"10",X"73",X"71",X"70",X"73",X"73",X"70",X"72",X"71",X"73",
		X"72",X"71",X"10",X"10",X"73",X"73",X"71",X"6B",X"64",X"10",X"10",X"10",X"10",X"64",X"10",X"10",
		X"10",X"65",X"10",X"10",X"10",X"10",X"10",X"10",X"65",X"10",X"10",X"64",X"10",X"10",X"64",X"10",
		X"10",X"6B",X"65",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"64",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"65",X"10",X"10",X"67",X"10",X"10",X"69",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"64",
		X"10",X"10",X"10",X"10",X"10",X"6B",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"65",X"67",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"68",
		X"10",X"10",X"64",X"66",X"65",X"66",X"10",X"10",X"65",X"64",X"10",X"10",X"64",X"10",X"10",X"10",
		X"66",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"6A",X"10",X"10",X"10",X"10",X"10",X"65",
		X"10",X"10",X"10",X"10",X"10",X"10",X"66",X"10",X"10",X"10",X"64",X"10",X"10",X"10",X"10",X"10",
		X"67",X"10",X"10",X"69",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"65",X"10",X"10",X"10",X"65",X"10",X"10",X"64",X"10",X"10",X"64",X"10",X"10",X"6A",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"66",X"64",X"10",
		X"10",X"10",X"10",X"10",X"65",X"10",X"10",X"6B",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"64",X"66",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"68",X"10",X"10",X"10",X"66",X"65",X"67",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"66",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"6A",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"65",X"67",X"64",X"66",X"10",X"10",X"10",X"67",X"10",X"10",X"66",
		X"10",X"10",X"10",X"10",X"10",X"69",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"64",X"10",X"10",X"10",X"10",X"10",X"6B",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"65",X"10",X"10",X"10",X"10",X"10",X"69",X"10",X"10",X"10",X"10",X"10",X"67",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"6A",X"10",X"10",X"66",X"65",X"66",X"64",X"10",X"10",X"10",X"10",X"10",X"10",
		X"66",X"64",X"10",X"10",X"67",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"68",X"10",X"10",
		X"10",X"10",X"10",X"65",X"10",X"10",X"65",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"64",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"6B",X"10",X"10",X"10",X"10",X"10",X"65",X"10",X"10",
		X"66",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"65",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"68",X"10",X"10",X"10",X"10",X"10",X"66",X"10",X"10",X"64",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"66",X"10",X"10",X"6B",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"67",X"65",X"66",X"64",X"67",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"64",X"10",X"10",X"6A",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"65",X"10",X"10",X"10",X"10",X"10",X"65",X"10",X"10",X"6B",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"65",
		X"64",X"10",X"10",X"66",X"10",X"10",X"10",X"10",X"10",X"68",X"10",X"10",X"10",X"10",X"10",X"64",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"64",X"10",X"10",
		X"10",X"10",X"10",X"6A",X"10",X"10",X"10",X"10",X"10",X"65",X"10",X"10",X"67",X"66",X"65",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"65",X"10",X"10",X"10",X"10",X"10",X"69",X"10",X"10",
		X"10",X"10",X"10",X"65",X"10",X"10",X"65",X"64",X"66",X"10",X"10",X"64",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"66",X"10",X"10",X"6A",X"10",X"10",X"10",X"10",X"10",X"65",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"66",X"10",X"10",X"64",X"10",X"10",X"10",X"10",X"10",X"65",X"10",
		X"10",X"68",X"10",X"10",X"10",X"10",X"10",X"66",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"65",
		X"10",X"10",X"66",X"10",X"10",X"10",X"10",X"10",X"66",X"10",X"10",X"69",X"6C",X"6F",X"6E",X"6D",
		X"6E",X"6F",X"6D",X"10",X"10",X"6C",X"6F",X"6C",X"6D",X"6E",X"6F",X"6C",X"6E",X"6D",X"6F",X"6C",
		X"10",X"10",X"6C",X"6C",X"6E",X"6A",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"10",X"10",X"8F",
		X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"10",X"10",X"8F",X"8F",X"8F",X"8F",
		X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"6D",X"6F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",
		X"8F",X"8F",X"8F",X"8F",X"6C",X"6E",X"8F",X"8F",X"8F",X"8F",X"5F",X"60",X"60",X"60",X"60",X"60",
		X"5C",X"60",X"60",X"5C",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"5C",X"60",X"60",
		X"5C",X"60",X"60",X"60",X"63",X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"63",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"63",X"10",X"10",X"69",X"5E",X"5C",
		X"60",X"60",X"5C",X"60",X"61",X"10",X"10",X"5E",X"60",X"5C",X"60",X"60",X"60",X"60",X"60",X"60",
		X"5C",X"61",X"10",X"10",X"5E",X"60",X"60",X"60",X"10",X"63",X"10",X"10",X"63",X"10",X"10",X"10",
		X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",
		X"10",X"6B",X"5F",X"61",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"69",X"63",X"10",X"10",X"10",
		X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"63",X"10",
		X"10",X"10",X"10",X"10",X"10",X"6B",X"63",X"10",X"10",X"10",X"5E",X"60",X"60",X"60",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"68",
		X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"63",
		X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"6A",X"63",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"63",X"10",X"10",X"63",X"10",X"10",X"10",
		X"10",X"10",X"10",X"69",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"63",
		X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"60",X"60",X"60",X"5E",X"60",
		X"10",X"10",X"10",X"60",X"60",X"60",X"60",X"5C",X"60",X"61",X"10",X"10",X"10",X"63",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"6B",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"68",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",
		X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"6A",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"69",X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"63",
		X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"6B",
		X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"5F",X"60",X"5D",
		X"60",X"60",X"60",X"10",X"10",X"10",X"60",X"60",X"60",X"60",X"10",X"10",X"10",X"10",X"10",X"63",
		X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"6A",X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"63",X"10",X"10",
		X"5F",X"61",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"68",X"10",X"10",
		X"10",X"10",X"10",X"63",X"10",X"10",X"5F",X"61",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"6B",X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",
		X"63",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",
		X"10",X"68",X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"63",X"10",X"10",X"10",X"63",X"10",
		X"10",X"10",X"63",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"6B",X"10",X"10",X"10",X"10",
		X"10",X"63",X"10",X"10",X"5E",X"60",X"60",X"60",X"61",X"10",X"10",X"10",X"63",X"10",X"10",X"10",
		X"5E",X"60",X"60",X"60",X"60",X"60",X"10",X"10",X"10",X"10",X"5F",X"61",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"6B",
		X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"68",X"10",X"10",X"10",X"10",X"63",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"6A",X"63",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"60",X"5C",X"60",
		X"10",X"10",X"10",X"5F",X"61",X"10",X"10",X"10",X"10",X"10",X"10",X"60",X"60",X"60",X"63",X"10",
		X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"63",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"6A",X"5E",X"62",X"10",X"10",X"63",X"10",X"10",X"10",
		X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"68",X"10",X"63",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",
		X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"69",X"5F",X"5D",X"60",X"60",
		X"5D",X"60",X"62",X"10",X"10",X"5F",X"5D",X"60",X"60",X"60",X"60",X"5D",X"60",X"60",X"60",X"62",
		X"10",X"10",X"5F",X"60",X"60",X"60",X"63",X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"63",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"63",X"10",X"10",X"68",
		X"5E",X"60",X"60",X"60",X"60",X"60",X"5D",X"60",X"60",X"5D",X"60",X"60",X"60",X"60",X"60",X"60",
		X"60",X"60",X"60",X"5D",X"60",X"60",X"5D",X"60",X"60",X"60",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",
		X"8F",X"9F",X"9E",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",
		X"8F",X"9C",X"9D",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"10",X"10",X"8F",X"8F",X"8F",
		X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"10",X"10",X"8F",X"8F",X"8F",X"8F",X"9C",X"9E",
		X"9F",X"9D",X"9E",X"9F",X"9D",X"10",X"10",X"9C",X"9F",X"9C",X"9D",X"9E",X"9F",X"9C",X"9E",X"9D",
		X"9F",X"9C",X"10",X"10",X"9F",X"9D",X"9C",X"8F",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"8F",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"8D",X"10",X"10",X"10",X"10",
		X"10",X"8F",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"8D",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"90",X"10",X"10",X"10",X"10",X"10",X"8F",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"8E",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"8F",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"90",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"8F",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"8F",X"10",X"10",X"10",X"10",X"10",X"91",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"8F",X"10",X"10",X"10",X"10",X"10",X"8D",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"8F",X"10",X"10",
		X"10",X"10",X"69",X"8E",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"8F",X"10",X"10",X"10",X"10",X"6B",X"8E",X"10",X"10",
		X"10",X"10",X"10",X"10",X"91",X"10",X"10",X"10",X"10",X"10",X"10",X"91",X"10",X"10",X"10",X"10",
		X"10",X"8F",X"10",X"10",X"10",X"10",X"69",X"8F",X"10",X"10",X"10",X"10",X"10",X"10",X"8D",X"10",
		X"10",X"10",X"10",X"10",X"68",X"8D",X"10",X"10",X"10",X"10",X"10",X"8F",X"10",X"10",X"10",X"10",
		X"6B",X"8E",X"10",X"10",X"10",X"10",X"10",X"68",X"8E",X"10",X"10",X"10",X"10",X"10",X"69",X"8F",
		X"10",X"10",X"10",X"10",X"10",X"8F",X"10",X"10",X"10",X"10",X"10",X"8D",X"10",X"10",X"10",X"10",
		X"10",X"69",X"8F",X"10",X"10",X"10",X"10",X"10",X"6B",X"8D",X"10",X"10",X"10",X"10",X"10",X"8F",
		X"10",X"10",X"10",X"10",X"10",X"8E",X"10",X"10",X"10",X"10",X"10",X"6A",X"8E",X"10",X"10",X"10",
		X"10",X"10",X"10",X"8E",X"10",X"10",X"10",X"10",X"10",X"8F",X"10",X"10",X"10",X"10",X"10",X"8F",
		X"10",X"10",X"10",X"10",X"10",X"6B",X"8D",X"10",X"10",X"10",X"10",X"10",X"10",X"90",X"10",X"10",
		X"10",X"10",X"10",X"8F",X"10",X"10",X"10",X"10",X"10",X"8E",X"10",X"10",X"10",X"10",X"10",X"68",
		X"8F",X"10",X"10",X"10",X"91",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"8F",X"10",X"10",
		X"10",X"10",X"10",X"8D",X"10",X"10",X"10",X"10",X"10",X"10",X"8E",X"10",X"10",X"10",X"8D",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"69",X"8F",X"10",X"10",X"10",X"10",X"10",X"8D",X"10",X"10",
		X"10",X"10",X"10",X"10",X"90",X"10",X"10",X"10",X"8E",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"68",X"8F",X"10",X"10",X"10",X"10",X"6B",X"8E",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"8D",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"8F",X"10",X"10",X"10",X"10",
		X"69",X"8E",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"90",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"8F",X"10",X"10",X"10",X"10",X"68",X"8F",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"6A",X"8F",
		X"10",X"10",X"10",X"10",X"6B",X"8D",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"6B",X"8F",X"10",X"10",X"10",X"10",X"10",X"90",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"8F",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"8F",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"8F",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"91",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"8F",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"8F",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"8F",X"9C",X"98",X"99",X"9A",
		X"98",X"8F",X"98",X"10",X"10",X"9B",X"99",X"98",X"8F",X"9B",X"98",X"9A",X"8F",X"9B",X"9A",X"8F",
		X"10",X"10",X"8F",X"99",X"9B",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"10",X"10",X"8F",
		X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"10",X"10",X"8F",X"8F",X"8F",X"8F",
		X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"99",X"98",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",
		X"8F",X"8F",X"8F",X"8F",X"9A",X"9B",X"8F",X"8F",X"8F",X"8F",X"CD",X"0E",X"16",X"3A",X"67",X"86",
		X"FE",X"01",X"28",X"35",X"3A",X"47",X"86",X"B7",X"28",X"2F",X"3A",X"33",X"86",X"B7",X"20",X"11",
		X"CF",X"50",X"08",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"32",X"20",X"55",X"50",X"00",X"18",
		X"27",X"CF",X"38",X"08",X"50",X"4C",X"41",X"59",X"45",X"52",X"53",X"20",X"31",X"20",X"41",X"4E",
		X"44",X"20",X"32",X"20",X"55",X"50",X"00",X"18",X"0F",X"CF",X"50",X"08",X"50",X"4C",X"41",X"59",
		X"45",X"52",X"20",X"31",X"20",X"55",X"50",X"00",X"3A",X"41",X"86",X"FE",X"02",X"CA",X"52",X"4C",
		X"3E",X"00",X"32",X"BE",X"81",X"CD",X"6B",X"4C",X"CD",X"D5",X"4B",X"3E",X"FE",X"32",X"9D",X"86",
		X"3E",X"FF",X"32",X"9F",X"86",X"3A",X"9D",X"86",X"B7",X"20",X"F5",X"AF",X"32",X"9F",X"86",X"3E",
		X"55",X"32",X"BE",X"81",X"C9",X"21",X"22",X"3B",X"3A",X"38",X"86",X"B7",X"CB",X"DF",X"28",X"02",
		X"E6",X"07",X"CB",X"27",X"06",X"00",X"4F",X"09",X"5E",X"23",X"56",X"EB",X"11",X"1F",X"8C",X"22",
		X"A2",X"86",X"ED",X"53",X"A0",X"86",X"3A",X"38",X"86",X"E6",X"03",X"FE",X"01",X"28",X"0C",X"FE",
		X"02",X"28",X"0D",X"FE",X"03",X"28",X"0E",X"FE",X"00",X"28",X"0F",X"E7",X"1A",X"05",X"00",X"C9",
		X"E7",X"1A",X"05",X"01",X"C9",X"E7",X"1A",X"05",X"02",X"C9",X"E7",X"1A",X"05",X"03",X"C9",X"AF",
		X"32",X"9F",X"86",X"3A",X"9D",X"86",X"3D",X"3D",X"32",X"9D",X"86",X"21",X"0A",X"90",X"06",X"1A",
		X"77",X"23",X"23",X"10",X"FB",X"E6",X"07",X"C0",X"ED",X"5B",X"A2",X"86",X"2A",X"A0",X"86",X"01",
		X"C6",X"FF",X"09",X"EB",X"06",X"00",X"0E",X"1A",X"ED",X"B0",X"22",X"A2",X"86",X"ED",X"53",X"A0",
		X"86",X"C9",X"AF",X"32",X"9F",X"86",X"32",X"9D",X"86",X"CD",X"D5",X"4B",X"06",X"20",X"C5",X"CD",
		X"38",X"4C",X"C1",X"10",X"F9",X"3E",X"32",X"CD",X"42",X"0E",X"C9",X"3A",X"41",X"86",X"B7",X"C0",
		X"3E",X"01",X"32",X"8F",X"86",X"3A",X"90",X"86",X"E6",X"6F",X"FE",X"07",X"28",X"F2",X"3A",X"90",
		X"86",X"B7",X"20",X"EC",X"C9",X"72",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"72",X"71",X"8F",
		X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"71",X"73",X"8F",
		X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"10",X"10",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",
		X"8F",X"8F",X"8F",X"8F",X"10",X"10",X"8F",X"8F",X"8F",X"69",X"71",X"72",X"70",X"72",X"70",X"72",
		X"70",X"10",X"10",X"73",X"71",X"70",X"73",X"73",X"70",X"72",X"8D",X"73",X"72",X"71",X"10",X"10",
		X"73",X"73",X"73",X"6B",X"64",X"10",X"10",X"10",X"10",X"64",X"10",X"10",X"10",X"65",X"10",X"10",
		X"10",X"10",X"10",X"10",X"8E",X"10",X"10",X"64",X"10",X"10",X"10",X"10",X"10",X"6B",X"65",X"10",
		X"10",X"10",X"10",X"65",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"8F",X"10",
		X"10",X"65",X"10",X"10",X"10",X"10",X"10",X"69",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"8D",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"6B",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"8F",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"68",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"65",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"90",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"6A",X"10",X"10",X"10",X"10",X"10",X"64",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"91",X"10",X"10",X"10",X"69",
		X"10",X"10",X"64",X"66",X"65",X"66",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"8D",X"64",X"10",X"10",X"6A",X"10",X"10",X"10",X"10",X"10",X"65",
		X"66",X"10",X"10",X"60",X"60",X"62",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"8E",
		X"62",X"10",X"10",X"6B",X"10",X"10",X"10",X"10",X"10",X"65",X"10",X"10",X"10",X"10",X"10",X"63",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"68",X"8F",X"63",X"10",X"10",X"68",X"10",X"10",
		X"10",X"10",X"10",X"66",X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"90",X"63",X"10",X"10",X"6A",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"63",X"10",
		X"10",X"69",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"5E",X"62",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"6B",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"60",X"5C",X"60",X"10",
		X"10",X"10",X"10",X"10",X"10",X"69",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"91",X"10",
		X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"6A",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"8D",X"10",X"10",X"10",X"63",X"10",X"10",X"10",
		X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"68",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"8E",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"6B",X"10",X"10",X"10",X"10",X"10",X"10",X"60",X"60",X"8D",X"60",X"60",X"60",
		X"61",X"10",X"10",X"10",X"5F",X"5D",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"8F",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"63",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"6B",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"8E",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"6A",X"10",X"10",X"10",X"10",X"68",X"8E",X"8D",X"8F",X"90",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"6B",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"60",X"5D",X"60",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"68",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"6A",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"69",X"10",X"10",X"10",X"10",X"10",X"64",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"6A",X"10",X"10",X"10",X"10",X"10",X"65",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"68",X"10",X"10",
		X"10",X"10",X"10",X"66",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"65",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"66",X"10",X"10",X"69",X"6C",X"6F",X"6E",X"6D",X"6E",X"6F",X"6D",X"10",
		X"10",X"6C",X"6F",X"6C",X"6D",X"6E",X"6F",X"6C",X"6E",X"6D",X"6F",X"6C",X"10",X"10",X"6C",X"6C",
		X"6E",X"6A",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"10",X"10",X"8F",X"8F",X"8F",X"8F",X"8F",
		X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"10",X"10",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",
		X"8F",X"8F",X"8F",X"6D",X"6F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",
		X"6C",X"6E",X"8F",X"8F",X"8F",X"8F",X"5F",X"60",X"60",X"60",X"60",X"60",X"5C",X"60",X"60",X"5C",
		X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"5C",X"60",X"60",X"5C",X"60",X"60",X"60",
		X"63",X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"63",X"10",X"10",X"63",X"10",X"10",X"69",X"5E",X"5C",X"60",X"60",X"5C",X"60",
		X"61",X"10",X"10",X"5E",X"60",X"5C",X"60",X"60",X"60",X"60",X"60",X"5C",X"60",X"61",X"10",X"10",
		X"5E",X"60",X"60",X"60",X"10",X"63",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"63",
		X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"6B",X"5F",X"61",
		X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"63",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"69",X"63",X"10",X"10",X"10",X"63",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"6B",X"63",X"10",X"10",X"10",X"5E",X"60",X"60",X"60",X"60",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"68",X"63",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"6A",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"69",
		X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"5E",X"60",X"60",X"60",X"60",X"60",X"60",X"5E",X"60",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"6B",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"91",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"68",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"69",X"8E",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"6A",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"6B",
		X"8D",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"91",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"69",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"6A",X"8E",X"10",X"10",X"10",X"10",X"63",
		X"10",X"10",X"8E",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"6B",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"69",X"8F",X"10",X"10",X"10",X"5F",X"5D",X"60",X"60",X"8F",X"10",X"10",X"10",
		X"10",X"5E",X"60",X"60",X"60",X"60",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"6A",X"8E",X"10",
		X"10",X"10",X"63",X"10",X"10",X"10",X"8E",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"6A",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"90",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"8D",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"68",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"8F",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"6B",X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"8D",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"68",X"10",X"10",
		X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"90",X"10",
		X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"6B",X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",
		X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"5E",X"60",X"60",X"60",
		X"60",X"60",X"10",X"10",X"10",X"10",X"5F",X"61",X"10",X"10",X"63",X"10",X"10",X"63",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"6B",X"10",X"10",X"10",X"10",
		X"63",X"10",X"10",X"10",X"63",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"68",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"63",X"10",
		X"10",X"63",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"6A",
		X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"5E",X"60",X"5C",X"61",X"10",X"10",X"10",X"5F",
		X"61",X"10",X"10",X"10",X"10",X"10",X"10",X"60",X"60",X"60",X"10",X"10",X"10",X"10",X"63",X"10",
		X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"6A",X"5E",X"62",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"63",X"10",
		X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"68",X"10",X"63",
		X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"63",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"69",X"5F",X"5D",X"60",X"60",X"5D",X"60",X"62",X"10",
		X"10",X"5F",X"5D",X"60",X"60",X"60",X"60",X"5D",X"60",X"60",X"60",X"62",X"10",X"10",X"5F",X"60",
		X"60",X"60",X"63",X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"63",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"63",X"10",X"10",X"68",X"5E",X"60",X"60",X"60",
		X"60",X"60",X"5D",X"60",X"60",X"5D",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"5D",
		X"60",X"60",X"5D",X"60",X"60",X"60",X"5F",X"60",X"60",X"60",X"60",X"60",X"5C",X"60",X"60",X"5C",
		X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"5C",X"60",X"60",X"60",
		X"63",X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"63",X"10",X"10",X"63",X"10",X"10",X"69",X"5E",X"5C",X"60",X"60",X"5C",X"60",
		X"61",X"10",X"10",X"5E",X"60",X"5C",X"60",X"60",X"60",X"60",X"5C",X"60",X"60",X"61",X"10",X"10",
		X"5E",X"60",X"60",X"60",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"63",
		X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"6B",X"10",X"10",
		X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"63",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"69",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"6B",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"68",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"6A",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"69",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"69",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"6B",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"68",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"6A",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"69",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"6B",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"91",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"91",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"6B",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"8E",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"90",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"6A",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"90",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"68",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"6B",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"91",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"68",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"90",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"6B",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"68",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"6B",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"68",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"6A",
		X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"60",X"60",X"60",X"10",X"10",X"10",X"10",X"63",X"10",
		X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"6A",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"63",X"10",
		X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"68",X"10",X"10",
		X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"63",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"69",X"5F",X"5D",X"60",X"60",X"5D",X"60",X"62",X"10",
		X"10",X"5F",X"5D",X"60",X"60",X"60",X"60",X"5D",X"60",X"60",X"60",X"62",X"10",X"10",X"5F",X"60",
		X"60",X"60",X"63",X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"63",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"63",X"10",X"10",X"68",X"5E",X"60",X"60",X"60",
		X"60",X"60",X"5D",X"60",X"60",X"5D",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"5D",
		X"60",X"60",X"5D",X"60",X"60",X"60",X"5F",X"60",X"60",X"60",X"60",X"60",X"5C",X"60",X"60",X"5C",
		X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"5C",X"60",X"60",X"5C",X"60",X"60",X"60",
		X"63",X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"63",X"10",X"10",X"63",X"10",X"10",X"69",X"5E",X"5C",X"60",X"60",X"60",X"60",
		X"61",X"10",X"10",X"5E",X"60",X"60",X"5C",X"60",X"60",X"60",X"60",X"60",X"60",X"61",X"10",X"10",
		X"5E",X"60",X"60",X"60",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"6B",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"69",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"6B",X"10",X"10",X"10",X"10",X"91",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"63",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"68",X"10",X"10",X"10",X"10",
		X"90",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"91",X"10",X"10",X"6A",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"91",X"10",X"10",X"10",X"10",X"10",X"90",X"10",X"10",X"69",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"90",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"69",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"91",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"6B",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"90",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"68",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"6A",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"91",X"10",
		X"10",X"69",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"90",X"10",X"10",X"6B",X"10",X"10",X"10",X"10",
		X"10",X"91",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"6B",X"10",X"10",X"10",X"10",X"10",X"90",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"6A",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"68",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"6B",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"91",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"91",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"68",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"90",X"10",X"10",X"10",X"10",X"91",X"10",X"10",X"90",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"6B",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"90",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"68",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"6B",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"68",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"6A",
		X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"68",X"10",X"10",X"10",X"10",X"63",X"10",
		X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"6A",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"63",X"10",
		X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"68",X"10",X"10",
		X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"10",X"10",X"63",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"69",X"5F",X"5D",X"60",X"60",X"5D",X"60",X"62",X"10",
		X"10",X"5F",X"5D",X"60",X"60",X"60",X"60",X"5D",X"60",X"60",X"60",X"62",X"10",X"10",X"5F",X"60",
		X"60",X"60",X"63",X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"63",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"63",X"10",X"10",X"63",X"10",X"10",X"68",X"5E",X"60",X"60",X"60",
		X"60",X"60",X"5D",X"60",X"60",X"5D",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"5D",
		X"60",X"60",X"5D",X"60",X"60",X"60",X"3A",X"8C",X"86",X"B7",X"C8",X"DD",X"7E",X"08",X"C6",X"08",
		X"67",X"DD",X"7E",X"0A",X"C6",X"08",X"6F",X"CD",X"FE",X"08",X"E5",X"3A",X"3D",X"86",X"4F",X"3A",
		X"3E",X"86",X"81",X"4F",X"3A",X"3F",X"86",X"81",X"4F",X"3A",X"40",X"86",X"81",X"B7",X"20",X"02",
		X"E1",X"C9",X"47",X"21",X"00",X"80",X"11",X"3C",X"80",X"7E",X"E6",X"1C",X"CA",X"0F",X"5A",X"7E",
		X"E6",X"03",X"FE",X"02",X"C2",X"0F",X"5A",X"D5",X"D9",X"D1",X"E1",X"E5",X"7D",X"E6",X"1F",X"4F",
		X"1A",X"E6",X"1F",X"B9",X"30",X"04",X"06",X"10",X"18",X"02",X"06",X"18",X"13",X"1A",X"1B",X"BC",
		X"38",X"0E",X"28",X"02",X"18",X"0E",X"1A",X"E6",X"E0",X"4F",X"7D",X"E6",X"E0",X"B9",X"38",X"04",
		X"0E",X"08",X"18",X"02",X"0E",X"04",X"CD",X"67",X"0C",X"FE",X"32",X"30",X"03",X"D9",X"18",X"0F",
		X"CB",X"4F",X"28",X"03",X"78",X"18",X"01",X"79",X"D9",X"4F",X"7E",X"E6",X"E3",X"B1",X"77",X"23",
		X"13",X"13",X"10",X"A5",X"E1",X"C9",X"3A",X"3D",X"86",X"4F",X"3A",X"3E",X"86",X"81",X"4F",X"3A",
		X"3F",X"86",X"81",X"4F",X"3A",X"40",X"86",X"81",X"47",X"C5",X"3A",X"3D",X"86",X"B7",X"28",X"1A",
		X"AF",X"32",X"3D",X"86",X"11",X"00",X"80",X"21",X"3D",X"86",X"1A",X"E6",X"60",X"FE",X"40",X"20",
		X"06",X"1A",X"E6",X"1C",X"28",X"01",X"34",X"13",X"10",X"F0",X"C1",X"C5",X"3A",X"3E",X"86",X"B7",
		X"28",X"1A",X"AF",X"32",X"3E",X"86",X"11",X"00",X"80",X"21",X"3E",X"86",X"1A",X"E6",X"60",X"FE",
		X"20",X"20",X"06",X"1A",X"E6",X"1C",X"28",X"01",X"34",X"13",X"10",X"F0",X"C1",X"C5",X"3A",X"3F",
		X"86",X"B7",X"28",X"1B",X"47",X"AF",X"32",X"3F",X"86",X"11",X"00",X"80",X"21",X"3F",X"86",X"1A",
		X"E6",X"60",X"FE",X"00",X"20",X"06",X"1A",X"E6",X"1C",X"28",X"01",X"34",X"13",X"10",X"F0",X"C1",
		X"3A",X"40",X"86",X"B7",X"28",X"1B",X"47",X"AF",X"32",X"40",X"86",X"11",X"00",X"80",X"21",X"40",
		X"86",X"1A",X"E6",X"60",X"FE",X"60",X"20",X"06",X"1A",X"E6",X"1C",X"28",X"01",X"34",X"13",X"10",
		X"F0",X"21",X"43",X"86",X"7E",X"32",X"42",X"86",X"C9",X"CD",X"50",X"0D",X"D2",X"12",X"0E",X"CD",
		X"F2",X"0C",X"D2",X"26",X"5C",X"FD",X"2A",X"B6",X"81",X"FD",X"66",X"02",X"FD",X"6E",X"01",X"E5",
		X"DD",X"E1",X"CD",X"82",X"5C",X"FD",X"CB",X"00",X"F6",X"FD",X"CB",X"0C",X"D6",X"FD",X"CB",X"00",
		X"D6",X"FD",X"36",X"0D",X"00",X"DD",X"E5",X"CD",X"EE",X"0D",X"FD",X"E1",X"DD",X"7E",X"0D",X"B7",
		X"C2",X"F7",X"5B",X"CD",X"FD",X"5A",X"FD",X"E5",X"CD",X"EE",X"0D",X"18",X"ED",X"DD",X"7E",X"0B",
		X"E6",X"07",X"4F",X"5F",X"DD",X"36",X"0B",X"00",X"DD",X"CB",X"0B",X"FE",X"FD",X"CB",X"00",X"4E",
		X"20",X"2A",X"CD",X"67",X"0C",X"E6",X"0C",X"CB",X"D7",X"FD",X"77",X"01",X"FD",X"CB",X"00",X"CE",
		X"C5",X"CD",X"D6",X"5B",X"21",X"C6",X"5B",X"06",X"00",X"09",X"5E",X"C1",X"CD",X"67",X"0C",X"FE",
		X"64",X"38",X"09",X"E6",X"07",X"28",X"F5",X"FE",X"04",X"28",X"F1",X"5F",X"CD",X"AC",X"14",X"16",
		X"00",X"CB",X"23",X"21",X"C7",X"5C",X"19",X"19",X"19",X"11",X"00",X"00",X"FD",X"36",X"04",X"00",
		X"FD",X"36",X"03",X"00",X"FD",X"36",X"0A",X"00",X"FD",X"36",X"09",X"00",X"78",X"A6",X"BE",X"28",
		X"0D",X"78",X"23",X"23",X"A6",X"BE",X"28",X"06",X"78",X"23",X"23",X"A6",X"BE",X"C0",X"23",X"7E",
		X"B9",X"20",X"04",X"DD",X"CB",X"0B",X"BE",X"5F",X"DD",X"7E",X"0B",X"E6",X"F8",X"B3",X"DD",X"77",
		X"0B",X"CB",X"23",X"CB",X"23",X"21",X"07",X"5D",X"19",X"7E",X"FD",X"77",X"03",X"23",X"7E",X"FD",
		X"77",X"04",X"23",X"7E",X"FD",X"77",X"09",X"23",X"7E",X"FD",X"77",X"0A",X"DD",X"CB",X"0B",X"7E",
		X"C8",X"DD",X"CB",X"0B",X"BE",X"DD",X"4E",X"0B",X"06",X"00",X"21",X"F7",X"5C",X"09",X"09",X"7E",
		X"23",X"66",X"6F",X"DD",X"CB",X"00",X"A6",X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",X"36",X"04",
		X"01",X"DD",X"CB",X"00",X"E6",X"C9",X"00",X"06",X"04",X"05",X"02",X"00",X"03",X"00",X"00",X"07",
		X"00",X"00",X"01",X"00",X"00",X"00",X"0E",X"00",X"3A",X"73",X"82",X"FD",X"BE",X"0C",X"38",X"04",
		X"CB",X"C9",X"18",X"04",X"28",X"02",X"CB",X"D9",X"3A",X"6D",X"82",X"FD",X"BE",X"06",X"38",X"03",
		X"CB",X"D1",X"C9",X"C8",X"CB",X"C1",X"C9",X"CB",X"77",X"28",X"08",X"01",X"02",X"02",X"CD",X"8B",
		X"1B",X"18",X"0A",X"CB",X"7F",X"28",X"06",X"01",X"02",X"02",X"CD",X"03",X"1C",X"3E",X"05",X"CD",
		X"45",X"0C",X"CD",X"2E",X"5C",X"21",X"43",X"86",X"7E",X"B7",X"28",X"0A",X"35",X"2B",X"7E",X"B7",
		X"28",X"04",X"35",X"C3",X"C5",X"5A",X"CD",X"68",X"0E",X"CD",X"EE",X"0D",X"18",X"FB",X"AF",X"DD",
		X"77",X"0D",X"FD",X"77",X"04",X"FD",X"77",X"03",X"FD",X"77",X"0A",X"FD",X"77",X"09",X"DD",X"CB",
		X"0C",X"96",X"DD",X"CB",X"00",X"A6",X"DD",X"CB",X"00",X"B6",X"21",X"4A",X"21",X"DD",X"75",X"05",
		X"DD",X"74",X"06",X"DD",X"36",X"04",X"01",X"DD",X"CB",X"00",X"E6",X"CD",X"EE",X"0D",X"DD",X"CB",
		X"00",X"66",X"20",X"F7",X"DD",X"36",X"0A",X"00",X"DD",X"36",X"08",X"00",X"DD",X"66",X"02",X"DD",
		X"6E",X"01",X"E5",X"FD",X"E1",X"FD",X"36",X"06",X"00",X"FD",X"36",X"0C",X"00",X"DD",X"CB",X"00",
		X"96",X"C9",X"CD",X"67",X"0C",X"CB",X"6F",X"28",X"1F",X"FD",X"36",X"08",X"02",X"FD",X"36",X"0A",
		X"C8",X"21",X"27",X"5D",X"FD",X"75",X"05",X"FD",X"74",X"06",X"FD",X"36",X"04",X"01",X"FD",X"CB",
		X"00",X"E6",X"3E",X"02",X"FD",X"77",X"0B",X"C9",X"FD",X"36",X"08",X"EE",X"FD",X"36",X"0A",X"C8",
		X"21",X"44",X"5D",X"FD",X"75",X"05",X"FD",X"74",X"06",X"FD",X"36",X"04",X"01",X"FD",X"CB",X"00",
		X"E6",X"3E",X"06",X"FD",X"77",X"0B",X"C9",X"03",X"00",X"03",X"00",X"03",X"00",X"0F",X"01",X"0C",
		X"02",X"03",X"00",X"0C",X"02",X"0C",X"02",X"0C",X"02",X"3C",X"03",X"30",X"04",X"0C",X"02",X"30",
		X"04",X"30",X"04",X"30",X"04",X"F0",X"05",X"C0",X"06",X"30",X"04",X"C0",X"06",X"C0",X"06",X"C0",
		X"06",X"C3",X"07",X"03",X"00",X"C0",X"06",X"61",X"5D",X"27",X"5D",X"27",X"5D",X"27",X"5D",X"7E",
		X"5D",X"44",X"5D",X"44",X"5D",X"44",X"5D",X"00",X"00",X"00",X"FE",X"00",X"03",X"00",X"FE",X"00",
		X"03",X"00",X"00",X"00",X"03",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"FD",X"00",X"02",X"00",
		X"FD",X"00",X"00",X"00",X"FD",X"00",X"FE",X"00",X"00",X"01",X"00",X"00",X"0C",X"0C",X"05",X"80",
		X"01",X"0C",X"0C",X"05",X"81",X"01",X"0C",X"0C",X"05",X"82",X"01",X"0C",X"0C",X"05",X"81",X"01",
		X"00",X"01",X"2C",X"5D",X"00",X"00",X"01",X"00",X"00",X"0C",X"0C",X"04",X"83",X"01",X"0C",X"0C",
		X"03",X"85",X"01",X"0C",X"0C",X"05",X"86",X"01",X"0C",X"0C",X"03",X"85",X"01",X"00",X"01",X"49",
		X"5D",X"00",X"00",X"01",X"00",X"00",X"0C",X"0C",X"04",X"87",X"01",X"0C",X"0C",X"03",X"88",X"01",
		X"0C",X"0C",X"05",X"89",X"01",X"0C",X"0C",X"03",X"88",X"01",X"00",X"01",X"66",X"5D",X"00",X"00",
		X"01",X"00",X"00",X"0C",X"0C",X"04",X"8A",X"01",X"0C",X"0C",X"03",X"8B",X"01",X"0C",X"0C",X"05",
		X"8C",X"01",X"0C",X"0C",X"03",X"8B",X"01",X"00",X"01",X"83",X"5D",X"CD",X"50",X"0D",X"D2",X"12",
		X"0E",X"CD",X"F2",X"0C",X"D2",X"8F",X"5E",X"FD",X"2A",X"B6",X"81",X"FD",X"22",X"A8",X"86",X"FD",
		X"66",X"02",X"FD",X"6E",X"01",X"E5",X"DD",X"E1",X"CD",X"97",X"5E",X"FD",X"CB",X"00",X"F6",X"FD",
		X"CB",X"00",X"D6",X"FD",X"36",X"0D",X"00",X"DD",X"E5",X"CD",X"EE",X"0D",X"FD",X"E1",X"DD",X"7E",
		X"0D",X"CB",X"47",X"20",X"15",X"CB",X"5F",X"20",X"63",X"DD",X"7E",X"0D",X"CB",X"87",X"CB",X"9F",
		X"DD",X"77",X"0D",X"FD",X"E5",X"CD",X"EE",X"0D",X"18",X"E2",X"3A",X"EE",X"82",X"B7",X"28",X"E9",
		X"21",X"FA",X"82",X"CB",X"CE",X"01",X"03",X"02",X"CD",X"8B",X"1B",X"3E",X"13",X"CD",X"45",X"0C",
		X"FD",X"E5",X"DD",X"E5",X"FD",X"21",X"43",X"22",X"CD",X"D6",X"0D",X"FD",X"21",X"43",X"22",X"CD",
		X"D6",X"0D",X"DD",X"E1",X"3E",X"5A",X"32",X"C4",X"89",X"3E",X"5B",X"32",X"C5",X"89",X"32",X"C6",
		X"89",X"FD",X"E1",X"3A",X"EE",X"82",X"B7",X"28",X"B0",X"3A",X"F6",X"82",X"DD",X"77",X"08",X"3A",
		X"F8",X"82",X"DD",X"77",X"0A",X"FD",X"E5",X"CD",X"EE",X"0D",X"18",X"E5",X"3A",X"1C",X"83",X"B7",
		X"28",X"97",X"21",X"28",X"83",X"CB",X"CE",X"01",X"03",X"02",X"CD",X"03",X"1C",X"3E",X"13",X"CD",
		X"45",X"0C",X"FD",X"E5",X"DD",X"E5",X"FD",X"21",X"43",X"22",X"CD",X"D6",X"0D",X"FD",X"21",X"43",
		X"22",X"CD",X"D6",X"0D",X"DD",X"E1",X"3E",X"5A",X"32",X"C4",X"89",X"3E",X"5B",X"32",X"C5",X"89",
		X"32",X"C6",X"89",X"FD",X"E1",X"3A",X"1C",X"83",X"B7",X"CA",X"D9",X"5D",X"3A",X"24",X"83",X"DD",
		X"77",X"08",X"3A",X"26",X"83",X"DD",X"77",X"0A",X"FD",X"E5",X"CD",X"EE",X"0D",X"18",X"E4",X"CD",
		X"68",X"0E",X"CD",X"EE",X"0D",X"18",X"FB",X"AF",X"DD",X"77",X"04",X"DD",X"77",X"03",X"DD",X"77",
		X"0A",X"DD",X"77",X"09",X"21",X"DB",X"5E",X"3A",X"38",X"86",X"E6",X"07",X"CB",X"27",X"16",X"00",
		X"5F",X"19",X"5E",X"23",X"56",X"FD",X"73",X"08",X"FD",X"72",X"0A",X"21",X"EB",X"5E",X"3A",X"38",
		X"86",X"E6",X"03",X"CB",X"27",X"16",X"00",X"5F",X"19",X"5E",X"23",X"56",X"FD",X"73",X"05",X"FD",
		X"72",X"06",X"FD",X"36",X"04",X"01",X"FD",X"CB",X"00",X"E6",X"C9",X"51",X"E0",X"DB",X"DF",X"A1",
		X"E2",X"DB",X"E2",X"D5",X"68",X"85",X"A1",X"95",X"E6",X"D5",X"E6",X"F3",X"5E",X"24",X"5F",X"55",
		X"5F",X"86",X"5F",X"00",X"00",X"01",X"00",X"00",X"14",X"14",X"03",X"C0",X"00",X"14",X"14",X"03",
		X"C0",X"01",X"14",X"14",X"03",X"C0",X"02",X"14",X"14",X"03",X"C0",X"03",X"14",X"14",X"03",X"C0",
		X"04",X"14",X"14",X"03",X"C0",X"05",X"14",X"14",X"03",X"C0",X"06",X"14",X"14",X"03",X"C0",X"07",
		X"00",X"01",X"F8",X"5E",X"00",X"00",X"01",X"00",X"00",X"14",X"14",X"03",X"C1",X"00",X"14",X"14",
		X"03",X"C1",X"01",X"14",X"14",X"03",X"C1",X"02",X"14",X"14",X"03",X"C1",X"03",X"14",X"14",X"03",
		X"C1",X"04",X"14",X"14",X"03",X"C1",X"05",X"14",X"14",X"03",X"C1",X"06",X"14",X"14",X"03",X"C1",
		X"07",X"00",X"01",X"29",X"5F",X"00",X"00",X"01",X"00",X"00",X"14",X"14",X"03",X"C2",X"00",X"14",
		X"14",X"03",X"C2",X"01",X"14",X"14",X"03",X"C2",X"02",X"14",X"14",X"03",X"C2",X"03",X"14",X"14",
		X"03",X"C2",X"04",X"14",X"14",X"03",X"C2",X"05",X"14",X"14",X"03",X"C2",X"06",X"14",X"14",X"03",
		X"C2",X"07",X"00",X"01",X"5A",X"5F",X"00",X"00",X"01",X"00",X"00",X"14",X"14",X"03",X"C3",X"00",
		X"14",X"14",X"03",X"C3",X"01",X"14",X"14",X"03",X"C3",X"02",X"14",X"14",X"03",X"C3",X"03",X"14",
		X"14",X"03",X"C3",X"04",X"14",X"14",X"03",X"C3",X"05",X"14",X"14",X"03",X"C3",X"06",X"14",X"14",
		X"03",X"C3",X"07",X"00",X"01",X"8B",X"5F",X"00",X"00",X"00",X"00",X"D7",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
