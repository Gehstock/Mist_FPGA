library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity romh is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of romh is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"AF",X"D3",X"03",X"C3",X"17",X"00",X"F5",X"C5",X"D5",X"E5",X"C3",X"9A",X"0E",X"00",
		X"F5",X"C5",X"D5",X"E5",X"C3",X"B0",X"0E",X"DB",X"02",X"E6",X"10",X"CA",X"62",X"0F",X"06",X"01",
		X"11",X"00",X"00",X"21",X"00",X"20",X"D3",X"04",X"70",X"7E",X"A8",X"CA",X"3D",X"00",X"4F",X"7D",
		X"E6",X"01",X"79",X"C2",X"3B",X"00",X"B2",X"57",X"C3",X"3D",X"00",X"B3",X"5F",X"23",X"7C",X"FE",
		X"40",X"C2",X"26",X"00",X"D3",X"04",X"2B",X"7C",X"FE",X"1F",X"CA",X"7A",X"00",X"7E",X"A8",X"CA",
		X"61",X"00",X"4F",X"7D",X"E6",X"01",X"79",X"C2",X"5F",X"00",X"B2",X"57",X"C3",X"61",X"00",X"B3",
		X"5F",X"78",X"2F",X"77",X"AE",X"CA",X"44",X"00",X"4F",X"7D",X"E6",X"01",X"79",X"C2",X"75",X"00",
		X"B2",X"57",X"C3",X"77",X"00",X"B3",X"5F",X"C3",X"44",X"00",X"D3",X"04",X"23",X"7C",X"FE",X"40",
		X"CA",X"9D",X"00",X"78",X"2F",X"AE",X"CA",X"98",X"00",X"4F",X"7D",X"E6",X"01",X"79",X"C2",X"96",
		X"00",X"B2",X"57",X"C3",X"98",X"00",X"B3",X"5F",X"AF",X"77",X"C3",X"7A",X"00",X"78",X"07",X"47",
		X"D2",X"23",X"00",X"7A",X"B3",X"CA",X"CC",X"00",X"EB",X"F9",X"11",X"00",X"20",X"06",X"00",X"21",
		X"00",X"00",X"39",X"0E",X"10",X"AF",X"29",X"DA",X"BB",X"00",X"2F",X"12",X"13",X"3E",X"08",X"12",
		X"13",X"0D",X"C2",X"B5",X"00",X"05",X"C2",X"AF",X"00",X"C3",X"1A",X"01",X"31",X"00",X"24",X"21",
		X"00",X"00",X"11",X"00",X"00",X"0E",X"04",X"AF",X"86",X"D3",X"04",X"23",X"47",X"79",X"BC",X"78",
		X"C2",X"D8",X"00",X"E5",X"21",X"1F",X"01",X"19",X"BE",X"3E",X"40",X"CA",X"F7",X"00",X"21",X"00",
		X"20",X"34",X"21",X"28",X"01",X"19",X"7E",X"21",X"29",X"20",X"19",X"77",X"E1",X"13",X"0C",X"0C",
		X"0C",X"0C",X"3E",X"24",X"B9",X"C2",X"D7",X"00",X"21",X"29",X"20",X"3A",X"00",X"20",X"A7",X"CA",
		X"00",X"00",X"11",X"08",X"30",X"3E",X"08",X"CD",X"30",X"01",X"D3",X"04",X"C3",X"1A",X"01",X"00",
		X"CA",X"40",X"19",X"47",X"E8",X"B8",X"00",X"BC",X"48",X"48",X"47",X"47",X"46",X"46",X"45",X"44",
		X"F5",X"7E",X"23",X"A7",X"FA",X"31",X"01",X"D6",X"30",X"F2",X"4D",X"01",X"47",X"13",X"7B",X"E6",
		X"1F",X"C2",X"46",X"01",X"14",X"14",X"04",X"C2",X"3D",X"01",X"C3",X"31",X"01",X"E5",X"D5",X"3C",
		X"FE",X"0B",X"FA",X"57",X"01",X"D6",X"06",X"21",X"71",X"01",X"01",X"0A",X"00",X"09",X"3D",X"C2",
		X"5D",X"01",X"EB",X"01",X"20",X"00",X"3E",X"0A",X"F5",X"1A",X"13",X"77",X"09",X"F1",X"3D",X"C2",
		X"68",X"01",X"D1",X"E1",X"13",X"F1",X"3D",X"C2",X"30",X"01",X"C9",X"3C",X"7E",X"66",X"66",X"66",
		X"66",X"66",X"66",X"7E",X"3C",X"18",X"1C",X"18",X"18",X"18",X"18",X"18",X"18",X"3C",X"3C",X"3C",
		X"7E",X"66",X"60",X"7C",X"3E",X"06",X"06",X"7E",X"7E",X"3C",X"7E",X"66",X"60",X"38",X"78",X"60",
		X"66",X"7E",X"3C",X"66",X"66",X"66",X"66",X"7E",X"7E",X"60",X"60",X"60",X"60",X"3E",X"3E",X"06",
		X"06",X"3E",X"7E",X"60",X"66",X"7E",X"3C",X"3C",X"3E",X"06",X"06",X"3E",X"7E",X"66",X"66",X"7E",
		X"3C",X"7E",X"7E",X"60",X"70",X"30",X"38",X"18",X"1C",X"0C",X"0C",X"3C",X"7E",X"66",X"66",X"3C",
		X"7E",X"66",X"66",X"7E",X"3C",X"3C",X"7E",X"66",X"66",X"7E",X"7C",X"60",X"60",X"7C",X"3C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"3C",X"7E",X"66",X"66",X"66",X"7E",
		X"7E",X"66",X"66",X"3E",X"7E",X"66",X"66",X"3E",X"7E",X"66",X"66",X"7E",X"3E",X"3C",X"7E",X"66",
		X"06",X"06",X"06",X"06",X"66",X"7E",X"3C",X"3E",X"7E",X"66",X"66",X"66",X"66",X"66",X"66",X"7E",
		X"3E",X"7E",X"7E",X"06",X"06",X"3E",X"3E",X"06",X"06",X"7E",X"7E",X"7E",X"7E",X"06",X"06",X"3E",
		X"3E",X"06",X"06",X"06",X"06",X"3C",X"7E",X"66",X"06",X"06",X"76",X"76",X"66",X"7E",X"3C",X"66",
		X"66",X"66",X"66",X"7E",X"7E",X"66",X"66",X"66",X"66",X"3C",X"3C",X"18",X"18",X"18",X"18",X"18",
		X"18",X"3C",X"3C",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"66",X"7E",X"3C",X"66",X"66",X"76",
		X"3E",X"1E",X"1E",X"3E",X"76",X"66",X"66",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"7E",
		X"7E",X"C3",X"C3",X"E7",X"E7",X"FF",X"FF",X"DB",X"C3",X"C3",X"C3",X"66",X"66",X"6E",X"6E",X"7E",
		X"7E",X"76",X"76",X"66",X"66",X"3C",X"7E",X"66",X"66",X"66",X"66",X"66",X"66",X"7E",X"3C",X"3E",
		X"7E",X"66",X"66",X"7E",X"3E",X"06",X"06",X"06",X"06",X"3C",X"7E",X"66",X"66",X"66",X"66",X"66",
		X"66",X"7E",X"5C",X"3E",X"7E",X"66",X"66",X"7E",X"3E",X"76",X"66",X"66",X"66",X"3C",X"7E",X"66",
		X"06",X"3E",X"7C",X"60",X"66",X"7E",X"3C",X"7E",X"7E",X"18",X"18",X"18",X"18",X"18",X"18",X"18",
		X"18",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"7E",X"3C",X"66",X"66",X"66",X"66",X"66",
		X"7E",X"3C",X"3C",X"18",X"18",X"C3",X"C3",X"C3",X"DB",X"FF",X"FF",X"E7",X"E7",X"C3",X"C3",X"66",
		X"66",X"7E",X"3C",X"18",X"18",X"3C",X"7E",X"66",X"66",X"66",X"66",X"7E",X"3C",X"18",X"18",X"18",
		X"18",X"18",X"18",X"7E",X"7E",X"60",X"70",X"38",X"1C",X"0E",X"06",X"7E",X"7E",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"00",X"00",X"C0",X"C0",X"10",X"38",X"38",X"38",X"38",X"38",X"38",X"38",X"38",
		X"7C",X"47",X"03",X"51",X"03",X"79",X"03",X"6F",X"03",X"8D",X"03",X"5B",X"03",X"83",X"03",X"65",
		X"03",X"97",X"03",X"A1",X"03",X"AB",X"03",X"29",X"03",X"33",X"03",X"3D",X"03",X"1F",X"03",X"89",
		X"0E",X"89",X"0E",X"89",X"0E",X"89",X"0E",X"89",X"0E",X"81",X"0D",X"81",X"0D",X"81",X"0D",X"81",
		X"0D",X"81",X"0D",X"2B",X"0C",X"2B",X"0C",X"8D",X"0C",X"8D",X"0C",X"C1",X"0C",X"E9",X"0C",X"17",
		X"0D",X"3D",X"0D",X"57",X"0D",X"71",X"0D",X"28",X"0B",X"7E",X"0B",X"CB",X"0B",X"F3",X"0B",X"13",
		X"0C",X"C1",X"03",X"D6",X"05",X"B5",X"07",X"ED",X"08",X"FD",X"09",X"02",X"04",X"11",X"06",X"D9",
		X"07",X"0D",X"09",X"1B",X"0A",X"43",X"04",X"4C",X"06",X"FD",X"07",X"2D",X"09",X"39",X"0A",X"84",
		X"04",X"87",X"06",X"21",X"08",X"4D",X"09",X"57",X"0A",X"C5",X"04",X"C2",X"06",X"45",X"08",X"6D",
		X"09",X"75",X"0A",X"06",X"05",X"FD",X"06",X"69",X"08",X"8D",X"09",X"93",X"0A",X"47",X"05",X"38",
		X"07",X"8D",X"08",X"AD",X"09",X"B1",X"0A",X"88",X"05",X"73",X"07",X"B1",X"08",X"CD",X"09",X"CF",
		X"0A",X"A2",X"05",X"89",X"07",X"C5",X"08",X"DD",X"09",X"D6",X"0A",X"BC",X"05",X"9F",X"07",X"D9",
		X"08",X"ED",X"09",X"DD",X"0A",X"CD",X"09",X"DD",X"09",X"ED",X"09",X"CF",X"0A",X"D6",X"0A",X"DD",
		X"0A",X"03",X"15",X"00",X"05",X"00",X"80",X"0D",X"00",X"80",X"0D",X"00",X"80",X"0F",X"00",X"C8",
		X"9F",X"00",X"F8",X"FF",X"00",X"C0",X"17",X"00",X"C0",X"3F",X"00",X"C0",X"7F",X"00",X"C0",X"1F",
		X"00",X"80",X"1F",X"00",X"00",X"07",X"00",X"80",X"0F",X"00",X"F8",X"3F",X"00",X"FC",X"7F",X"00",
		X"CE",X"FF",X"01",X"C6",X"FF",X"03",X"C6",X"1F",X"17",X"C6",X"1F",X"0E",X"C6",X"1F",X"14",X"FA",
		X"3F",X"20",X"03",X"15",X"00",X"05",X"00",X"80",X"0D",X"00",X"80",X"0D",X"00",X"80",X"0F",X"00",
		X"C8",X"9F",X"00",X"F8",X"FF",X"00",X"C0",X"17",X"00",X"C0",X"3F",X"00",X"C0",X"7F",X"00",X"C0",
		X"1F",X"00",X"80",X"1F",X"00",X"00",X"07",X"00",X"80",X"0F",X"00",X"F8",X"3F",X"00",X"FC",X"7F",
		X"00",X"CE",X"FF",X"01",X"C6",X"FF",X"07",X"C6",X"1F",X"1E",X"C6",X"1F",X"70",X"C6",X"1F",X"00",
		X"FA",X"3F",X"00",X"03",X"15",X"00",X"05",X"00",X"80",X"0D",X"00",X"80",X"0D",X"00",X"80",X"0F",
		X"00",X"C8",X"9F",X"00",X"F8",X"FF",X"00",X"C0",X"17",X"00",X"C0",X"3F",X"00",X"C0",X"7F",X"00",
		X"C0",X"1F",X"00",X"80",X"1F",X"00",X"00",X"07",X"00",X"80",X"0F",X"00",X"F8",X"3F",X"00",X"FC",
		X"FF",X"01",X"CE",X"FF",X"0F",X"C6",X"1F",X"7F",X"C6",X"1F",X"00",X"C6",X"1F",X"00",X"C6",X"1F",
		X"00",X"FA",X"3F",X"00",X"03",X"15",X"00",X"05",X"00",X"80",X"0D",X"00",X"80",X"0D",X"00",X"80",
		X"0F",X"00",X"C8",X"9F",X"00",X"F8",X"FF",X"00",X"C0",X"17",X"00",X"C0",X"3F",X"00",X"C0",X"7F",
		X"00",X"C0",X"1F",X"00",X"80",X"1F",X"00",X"00",X"07",X"08",X"80",X"0F",X"F0",X"F8",X"FF",X"1F",
		X"FC",X"FF",X"0F",X"CE",X"FF",X"00",X"C6",X"1F",X"00",X"C6",X"1F",X"00",X"C6",X"1F",X"00",X"C6",
		X"1F",X"00",X"FA",X"3F",X"00",X"03",X"15",X"00",X"05",X"00",X"80",X"0D",X"00",X"80",X"0D",X"00",
		X"80",X"0F",X"00",X"C8",X"9F",X"00",X"F8",X"FF",X"00",X"C0",X"17",X"00",X"C0",X"3F",X"00",X"C0",
		X"7F",X"00",X"C0",X"1F",X"00",X"80",X"1F",X"C0",X"00",X"07",X"38",X"80",X"0F",X"0C",X"F8",X"FF",
		X"0F",X"FC",X"FF",X"03",X"CE",X"FF",X"00",X"C6",X"1F",X"00",X"C6",X"1F",X"00",X"C6",X"1F",X"00",
		X"C6",X"1F",X"00",X"FA",X"3F",X"00",X"03",X"15",X"00",X"05",X"00",X"80",X"0D",X"00",X"80",X"0D",
		X"00",X"80",X"0F",X"00",X"C8",X"9F",X"00",X"F8",X"FF",X"00",X"C0",X"17",X"00",X"C0",X"3F",X"00",
		X"C0",X"7F",X"00",X"C0",X"1F",X"C0",X"80",X"1F",X"70",X"00",X"07",X"3C",X"80",X"0F",X"0F",X"F8",
		X"FF",X"03",X"FC",X"FF",X"01",X"CE",X"FF",X"00",X"C6",X"1F",X"00",X"C6",X"1F",X"00",X"C6",X"1F",
		X"00",X"C6",X"1F",X"00",X"FA",X"3F",X"00",X"03",X"15",X"00",X"05",X"00",X"80",X"0D",X"00",X"80",
		X"0D",X"00",X"80",X"0F",X"00",X"C8",X"9F",X"00",X"F8",X"FF",X"00",X"C0",X"17",X"80",X"C0",X"3F",
		X"50",X"C0",X"7F",X"60",X"C0",X"1F",X"30",X"80",X"1F",X"38",X"00",X"07",X"1C",X"80",X"0F",X"0E",
		X"F8",X"FF",X"07",X"FC",X"FF",X"03",X"CE",X"FF",X"01",X"C6",X"1F",X"00",X"C6",X"1F",X"00",X"C6",
		X"1F",X"00",X"C6",X"1F",X"00",X"FA",X"3F",X"00",X"02",X"0C",X"F0",X"3F",X"F0",X"3F",X"E0",X"3D",
		X"C0",X"79",X"C0",X"71",X"C0",X"E1",X"C0",X"E1",X"E0",X"60",X"70",X"70",X"34",X"34",X"38",X"38",
		X"F0",X"F0",X"02",X"0C",X"F0",X"3F",X"E0",X"3F",X"C0",X"1F",X"C0",X"1F",X"C0",X"1F",X"00",X"1F",
		X"00",X"1E",X"00",X"1C",X"00",X"0C",X"00",X"0D",X"00",X"0E",X"00",X"3C",X"02",X"0C",X"F0",X"3F",
		X"F0",X"3F",X"E0",X"1F",X"C0",X"0F",X"80",X"1F",X"00",X"3E",X"C0",X"7D",X"E0",X"78",X"70",X"30",
		X"34",X"34",X"38",X"38",X"F0",X"F0",X"03",X"13",X"40",X"01",X"00",X"60",X"03",X"00",X"E0",X"03",
		X"00",X"F4",X"17",X"00",X"FC",X"1F",X"00",X"E0",X"02",X"00",X"E0",X"0F",X"00",X"E0",X"03",X"00",
		X"E0",X"03",X"00",X"C0",X"01",X"00",X"E0",X"03",X"00",X"FC",X"0F",X"00",X"FE",X"3F",X"00",X"F3",
		X"7F",X"00",X"F3",X"E3",X"02",X"F3",X"C3",X"01",X"F1",X"83",X"02",X"FE",X"03",X"04",X"FC",X"07",
		X"00",X"03",X"13",X"40",X"01",X"00",X"60",X"03",X"00",X"E0",X"03",X"00",X"F4",X"17",X"00",X"FC",
		X"1F",X"00",X"E0",X"02",X"00",X"E0",X"0F",X"00",X"E0",X"03",X"00",X"E0",X"03",X"00",X"C0",X"01",
		X"00",X"E0",X"03",X"00",X"FC",X"0F",X"00",X"FE",X"1F",X"00",X"F3",X"7F",X"00",X"F3",X"E3",X"01",
		X"F3",X"03",X"07",X"F1",X"03",X"00",X"FE",X"03",X"00",X"FC",X"07",X"00",X"03",X"13",X"40",X"01",
		X"00",X"60",X"03",X"00",X"E0",X"03",X"00",X"F4",X"17",X"00",X"FC",X"1F",X"00",X"E0",X"02",X"00",
		X"E0",X"0F",X"00",X"E0",X"03",X"00",X"E0",X"03",X"00",X"C0",X"01",X"00",X"E0",X"03",X"00",X"FC",
		X"1F",X"00",X"FE",X"FF",X"00",X"F3",X"FF",X"07",X"F3",X"03",X"00",X"F3",X"03",X"00",X"F1",X"03",
		X"00",X"FE",X"03",X"00",X"FC",X"07",X"00",X"03",X"13",X"40",X"01",X"00",X"60",X"03",X"00",X"E0",
		X"03",X"00",X"F4",X"17",X"00",X"FC",X"1F",X"00",X"E0",X"02",X"00",X"E0",X"0F",X"00",X"E0",X"03",
		X"00",X"E0",X"03",X"00",X"C0",X"01",X"01",X"E0",X"03",X"1E",X"FC",X"FF",X"03",X"FE",X"FF",X"03",
		X"F3",X"0F",X"00",X"F3",X"03",X"00",X"F3",X"03",X"00",X"F1",X"03",X"00",X"FE",X"03",X"00",X"FC",
		X"07",X"00",X"03",X"13",X"40",X"01",X"00",X"60",X"03",X"00",X"E0",X"03",X"00",X"F4",X"17",X"00",
		X"FC",X"1F",X"00",X"E0",X"02",X"00",X"E0",X"0F",X"00",X"E0",X"03",X"00",X"E0",X"03",X"0C",X"C0",
		X"81",X"03",X"E0",X"C3",X"00",X"FC",X"FF",X"00",X"FE",X"3F",X"00",X"F3",X"0F",X"00",X"F3",X"03",
		X"00",X"F3",X"03",X"00",X"F1",X"03",X"00",X"FE",X"03",X"00",X"FC",X"07",X"00",X"03",X"13",X"40",
		X"01",X"00",X"60",X"03",X"00",X"E0",X"03",X"00",X"F4",X"17",X"00",X"FC",X"1F",X"00",X"E0",X"02",
		X"00",X"E0",X"0F",X"00",X"E0",X"03",X"00",X"E0",X"03",X"06",X"C0",X"C1",X"03",X"E0",X"F3",X"00",
		X"FC",X"3F",X"00",X"FE",X"1F",X"00",X"F3",X"0F",X"00",X"F3",X"03",X"00",X"F3",X"03",X"00",X"F1",
		X"03",X"00",X"FE",X"03",X"00",X"FC",X"07",X"00",X"03",X"13",X"40",X"01",X"00",X"60",X"03",X"00",
		X"E0",X"03",X"00",X"F4",X"17",X"00",X"FC",X"1F",X"00",X"E0",X"02",X"04",X"E0",X"8F",X"06",X"E0",
		X"03",X"03",X"E0",X"83",X"03",X"C0",X"C1",X"01",X"E0",X"E3",X"00",X"FC",X"7F",X"00",X"FE",X"3F",
		X"00",X"F3",X"1F",X"00",X"F3",X"03",X"00",X"F3",X"03",X"00",X"F1",X"03",X"00",X"FE",X"03",X"00",
		X"FC",X"07",X"00",X"02",X"0A",X"F8",X"07",X"70",X"0F",X"70",X"0E",X"70",X"1C",X"30",X"1C",X"38",
		X"0C",X"1C",X"0E",X"0C",X"06",X"0E",X"07",X"3C",X"1E",X"02",X"0A",X"FC",X"03",X"F8",X"03",X"F0",
		X"03",X"F0",X"03",X"C0",X"03",X"C0",X"03",X"80",X"03",X"80",X"01",X"C0",X"01",X"80",X"07",X"02",
		X"0A",X"FC",X"03",X"F8",X"01",X"F0",X"00",X"E0",X"01",X"C8",X"03",X"9C",X"07",X"0E",X"07",X"06",
		X"03",X"87",X"03",X"1E",X"0F",X"02",X"11",X"50",X"00",X"D8",X"00",X"F8",X"00",X"FE",X"03",X"B8",
		X"00",X"F8",X"01",X"F8",X"00",X"60",X"00",X"F0",X"00",X"FC",X"03",X"FE",X"07",X"FF",X"06",X"F9",
		X"0C",X"F9",X"18",X"F9",X"20",X"FE",X"01",X"FE",X"01",X"02",X"11",X"50",X"00",X"D8",X"00",X"F8",
		X"00",X"FE",X"03",X"B8",X"00",X"F8",X"01",X"F8",X"00",X"60",X"00",X"F0",X"00",X"FC",X"03",X"FE",
		X"0F",X"FF",X"3C",X"F9",X"60",X"F9",X"00",X"F9",X"00",X"FE",X"01",X"FE",X"01",X"02",X"11",X"50");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
