library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity cpu2_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of cpu2_rom is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"E8",X"ED",X"08",X"86",X"00",X"A7",X"42",X"39",X"30",X"88",X"10",X"33",X"44",X"8C",X"53",
		X"B0",X"25",X"B8",X"39",X"96",X"AF",X"26",X"05",X"96",X"38",X"27",X"05",X"39",X"96",X"39",X"26",
		X"FB",X"DC",X"1A",X"10",X"83",X"04",X"80",X"25",X"F3",X"10",X"83",X"05",X"81",X"24",X"ED",X"DC",
		X"1C",X"10",X"83",X"06",X"00",X"25",X"E5",X"10",X"83",X"07",X"01",X"24",X"DF",X"96",X"AF",X"26",
		X"04",X"0C",X"38",X"20",X"02",X"0C",X"39",X"8E",X"53",X"50",X"CE",X"51",X"BC",X"A6",X"84",X"26",
		X"3C",X"6A",X"84",X"7C",X"52",X"34",X"86",X"0A",X"A7",X"03",X"B6",X"52",X"41",X"8B",X"40",X"2B",
		X"16",X"CC",X"FC",X"80",X"A7",X"43",X"E7",X"C4",X"CC",X"FF",X"18",X"ED",X"06",X"CC",X"00",X"00",
		X"ED",X"08",X"86",X"40",X"A7",X"42",X"39",X"CC",X"04",X"80",X"A7",X"43",X"E7",X"C4",X"CC",X"00",
		X"E8",X"ED",X"06",X"CC",X"00",X"00",X"ED",X"08",X"86",X"C0",X"A7",X"42",X"39",X"30",X"88",X"10",
		X"33",X"44",X"8C",X"53",X"B0",X"25",X"B6",X"39",X"CC",X"37",X"D1",X"DD",X"D0",X"39",X"96",X"D0",
		X"8B",X"59",X"97",X"D0",X"98",X"D1",X"97",X"D1",X"39",X"0F",X"DC",X"8E",X"52",X"F0",X"CE",X"51",
		X"A4",X"B6",X"57",X"DD",X"27",X"02",X"0A",X"DC",X"B6",X"54",X"60",X"26",X"0B",X"B6",X"52",X"34",
		X"27",X"06",X"86",X"0C",X"97",X"34",X"20",X"04",X"86",X"06",X"97",X"34",X"A6",X"84",X"27",X"1D",
		X"CC",X"A0",X"ED",X"34",X"06",X"A6",X"84",X"4C",X"27",X"0A",X"4C",X"26",X"75",X"6A",X"0E",X"26",
		X"02",X"6C",X"84",X"39",X"A6",X"03",X"10",X"8E",X"F5",X"98",X"48",X"6E",X"B6",X"30",X"88",X"10",
		X"33",X"44",X"0A",X"34",X"10",X"26",X"FF",X"D4",X"B6",X"54",X"40",X"10",X"26",X"04",X"9E",X"39",
		X"A6",X"43",X"E6",X"0C",X"F3",X"57",X"C0",X"A7",X"43",X"E7",X"0C",X"A6",X"C4",X"E6",X"0D",X"F3",
		X"57",X"C2",X"A7",X"C4",X"E7",X"0D",X"39",X"0A",X"E8",X"26",X"2E",X"CC",X"06",X"09",X"BD",X"8F",
		X"0C",X"C6",X"04",X"BD",X"A5",X"AB",X"20",X"21",X"0A",X"D5",X"26",X"1D",X"7C",X"57",X"DE",X"86",
		X"06",X"D6",X"DD",X"CB",X"05",X"BD",X"8F",X"0C",X"D6",X"DD",X"0C",X"DD",X"96",X"DD",X"81",X"03",
		X"25",X"04",X"C6",X"02",X"D7",X"DD",X"BD",X"A5",X"AB",X"7A",X"52",X"34",X"4F",X"A7",X"84",X"A7",
		X"43",X"39",X"81",X"78",X"24",X"36",X"8D",X"A8",X"6A",X"84",X"26",X"12",X"A6",X"03",X"10",X"8E",
		X"F5",X"AE",X"A6",X"A6",X"27",X"E6",X"4C",X"27",X"BF",X"4C",X"27",X"AB",X"20",X"DB",X"86",X"5B",
		X"E6",X"03",X"C0",X"06",X"27",X"05",X"5A",X"27",X"02",X"86",X"AF",X"97",X"F6",X"A6",X"84",X"46",
		X"46",X"84",X"07",X"9B",X"F6",X"A7",X"41",X"86",X"40",X"A7",X"42",X"39",X"E6",X"03",X"C1",X"08",
		X"22",X"33",X"27",X"09",X"C1",X"06",X"24",X"12",X"7C",X"57",X"DC",X"0C",X"EC",X"86",X"18",X"A7",
		X"84",X"BD",X"92",X"1A",X"CC",X"06",X"04",X"7E",X"8F",X"0C",X"86",X"10",X"A7",X"84",X"C1",X"06",
		X"26",X"0A",X"7C",X"57",X"DB",X"0C",X"EB",X"BD",X"92",X"0A",X"20",X"03",X"BD",X"92",X"12",X"CC",
		X"06",X"01",X"7E",X"8F",X"0C",X"86",X"18",X"A7",X"84",X"BD",X"92",X"58",X"C1",X"09",X"26",X"05",
		X"7C",X"57",X"D7",X"20",X"03",X"7C",X"57",X"D8",X"7C",X"57",X"D0",X"F6",X"57",X"D0",X"86",X"07",
		X"7E",X"8F",X"0C",X"96",X"DC",X"27",X"04",X"6F",X"0A",X"20",X"03",X"BD",X"A6",X"CE",X"A6",X"0B",
		X"27",X"04",X"6A",X"0B",X"20",X"5E",X"A6",X"0A",X"26",X"04",X"E6",X"02",X"20",X"12",X"6A",X"0A",
		X"26",X"09",X"B6",X"52",X"41",X"80",X"80",X"A7",X"02",X"20",X"05",X"BD",X"A5",X"DE",X"E7",X"02",
		X"E0",X"01",X"27",X"2D",X"D7",X"F6",X"A6",X"04",X"AB",X"05",X"44",X"69",X"05",X"44",X"69",X"05",
		X"44",X"69",X"05",X"44",X"69",X"05",X"E6",X"05",X"C4",X"0F",X"E7",X"05",X"D6",X"F6",X"2A",X"01",
		X"40",X"AB",X"01",X"A7",X"01",X"A0",X"02",X"8B",X"01",X"81",X"02",X"22",X"04",X"A6",X"02",X"A7",
		X"01",X"E6",X"01",X"BD",X"A6",X"21",X"CC",X"00",X"C4",X"BD",X"A6",X"6F",X"DC",X"3A",X"ED",X"06",
		X"DC",X"3C",X"ED",X"08",X"A6",X"43",X"E6",X"0C",X"E3",X"06",X"F3",X"57",X"C0",X"A7",X"43",X"E7",
		X"0C",X"A6",X"C4",X"E6",X"0D",X"E3",X"08",X"F3",X"57",X"C2",X"A7",X"C4",X"E7",X"0D",X"10",X"8E",
		X"F5",X"DA",X"B6",X"57",X"D6",X"48",X"10",X"AE",X"A6",X"A6",X"01",X"8B",X"08",X"44",X"44",X"44",
		X"44",X"A6",X"A6",X"A7",X"41",X"5F",X"A6",X"01",X"2A",X"02",X"C6",X"40",X"D7",X"F6",X"10",X"8E",
		X"F5",X"B9",X"B6",X"57",X"C7",X"44",X"44",X"44",X"44",X"84",X"07",X"A6",X"A6",X"9B",X"F6",X"A7",
		X"42",X"7E",X"A5",X"72",X"BD",X"A6",X"CE",X"A6",X"43",X"80",X"80",X"8B",X"34",X"81",X"68",X"22",
		X"4A",X"A6",X"C4",X"80",X"78",X"8B",X"34",X"81",X"68",X"22",X"40",X"A6",X"02",X"E6",X"04",X"26",
		X"1A",X"6A",X"04",X"CC",X"80",X"78",X"BD",X"A5",X"E0",X"E7",X"02",X"BD",X"A0",X"9E",X"84",X"01",
		X"8B",X"58",X"85",X"01",X"27",X"01",X"40",X"AB",X"02",X"A7",X"02",X"A0",X"01",X"27",X"1C",X"C6",
		X"08",X"81",X"80",X"25",X"01",X"50",X"EB",X"01",X"E7",X"01",X"BD",X"A6",X"21",X"CC",X"01",X"10",
		X"BD",X"A6",X"6F",X"DC",X"3A",X"ED",X"06",X"DC",X"3C",X"ED",X"08",X"A6",X"43",X"E6",X"0C",X"E3",
		X"06",X"F3",X"57",X"C0",X"A7",X"43",X"E7",X"0C",X"A6",X"C4",X"E6",X"0D",X"E3",X"08",X"F3",X"57",
		X"C2",X"A7",X"C4",X"E7",X"0D",X"B6",X"57",X"C7",X"44",X"84",X"03",X"8B",X"32",X"A7",X"41",X"7E",
		X"A5",X"83",X"B6",X"57",X"C7",X"84",X"03",X"26",X"03",X"BD",X"A6",X"CE",X"6A",X"05",X"26",X"02",
		X"8D",X"41",X"A6",X"43",X"E6",X"0C",X"F3",X"57",X"C0",X"A7",X"43",X"E7",X"0C",X"EC",X"06",X"A3",
		X"08",X"ED",X"06",X"A6",X"C4",X"E6",X"0D",X"E3",X"06",X"F3",X"57",X"C2",X"A7",X"C4",X"E7",X"0D",
		X"BD",X"A3",X"56",X"7E",X"A5",X"83",X"A6",X"04",X"46",X"24",X"17",X"46",X"24",X"06",X"86",X"20",
		X"A0",X"05",X"20",X"02",X"A6",X"05",X"47",X"47",X"10",X"8E",X"F5",X"C1",X"31",X"A6",X"A6",X"A4",
		X"A7",X"41",X"39",X"A6",X"04",X"48",X"10",X"8E",X"F5",X"CA",X"6E",X"B6",X"6C",X"04",X"86",X"20",
		X"A7",X"05",X"EC",X"06",X"47",X"56",X"47",X"56",X"47",X"56",X"47",X"56",X"ED",X"08",X"39",X"6C",
		X"04",X"86",X"0C",X"A7",X"05",X"CC",X"00",X"00",X"ED",X"08",X"39",X"6F",X"04",X"86",X"20",X"A7",
		X"05",X"CC",X"00",X"00",X"ED",X"08",X"39",X"B6",X"57",X"C7",X"84",X"03",X"26",X"03",X"BD",X"A6",
		X"CE",X"A6",X"04",X"27",X"11",X"4A",X"26",X"3E",X"A6",X"0A",X"AB",X"01",X"A7",X"01",X"6A",X"05",
		X"26",X"21",X"6C",X"04",X"20",X"1D",X"6A",X"05",X"26",X"2C",X"6C",X"04",X"BD",X"A0",X"9E",X"84",
		X"3F",X"8B",X"70",X"A7",X"05",X"A6",X"43",X"2B",X"06",X"86",X"FC",X"A7",X"0A",X"20",X"04",X"86",
		X"04",X"A7",X"0A",X"E6",X"01",X"BD",X"A6",X"21",X"CC",X"01",X"80",X"BD",X"A6",X"6F",X"DC",X"3A",
		X"ED",X"06",X"DC",X"3C",X"ED",X"08",X"A6",X"43",X"E6",X"0C",X"E3",X"06",X"F3",X"57",X"C0",X"A7",
		X"43",X"E7",X"0C",X"A6",X"C4",X"E6",X"0D",X"E3",X"08",X"F3",X"57",X"C2",X"A7",X"C4",X"E7",X"0D",
		X"6A",X"0B",X"26",X"04",X"86",X"2F",X"A7",X"0B",X"A6",X"0B",X"44",X"44",X"44",X"8B",X"2C",X"A7",
		X"41",X"7E",X"A5",X"83",X"B6",X"57",X"C7",X"84",X"03",X"26",X"03",X"BD",X"A6",X"CE",X"8D",X"03",
		X"7E",X"A5",X"83",X"A6",X"04",X"27",X"05",X"4A",X"27",X"0E",X"20",X"2E",X"6A",X"02",X"26",X"2A",
		X"6C",X"04",X"86",X"40",X"A7",X"05",X"20",X"42",X"6A",X"05",X"27",X"05",X"BD",X"A1",X"00",X"20",
		X"39",X"6C",X"04",X"CC",X"00",X"00",X"ED",X"0A",X"A6",X"43",X"2A",X"07",X"CC",X"FF",X"F6",X"ED",
		X"08",X"20",X"27",X"CC",X"00",X"0A",X"ED",X"08",X"20",X"20",X"EC",X"06",X"E3",X"08",X"ED",X"06",
		X"A6",X"43",X"E6",X"0C",X"E3",X"06",X"F3",X"57",X"C0",X"A7",X"43",X"E7",X"0C",X"A6",X"C4",X"E6",
		X"0D",X"E3",X"0A",X"F3",X"57",X"C2",X"A7",X"C4",X"E7",X"0D",X"A6",X"04",X"27",X"33",X"4A",X"26",
		X"07",X"A6",X"05",X"84",X"01",X"27",X"03",X"39",X"6A",X"05",X"A6",X"04",X"4A",X"27",X"0A",X"A6",
		X"06",X"2B",X"10",X"10",X"8E",X"F5",X"D6",X"20",X"0E",X"A6",X"43",X"2B",X"06",X"10",X"8E",X"F5",
		X"D6",X"20",X"04",X"10",X"8E",X"F5",X"D2",X"A6",X"05",X"46",X"46",X"84",X"03",X"A6",X"A6",X"A7",
		X"41",X"39",X"B6",X"57",X"C7",X"84",X"03",X"26",X"03",X"BD",X"A6",X"CE",X"6A",X"04",X"26",X"1E",
		X"BD",X"A0",X"9E",X"AB",X"01",X"A7",X"01",X"E6",X"01",X"BD",X"A6",X"21",X"CC",X"01",X"50",X"BD",
		X"A6",X"6F",X"DC",X"3A",X"ED",X"06",X"DC",X"3C",X"ED",X"08",X"A6",X"05",X"A7",X"04",X"A6",X"43",
		X"E6",X"0C",X"E3",X"06",X"F3",X"57",X"C0",X"A7",X"43",X"E7",X"0C",X"A6",X"C4",X"E6",X"0D",X"E3",
		X"08",X"F3",X"57",X"C2",X"A7",X"C4",X"E7",X"0D",X"B6",X"57",X"C7",X"44",X"84",X"03",X"8B",X"20",
		X"A7",X"41",X"86",X"40",X"A7",X"42",X"7E",X"A5",X"83",X"B6",X"57",X"C7",X"84",X"07",X"26",X"03",
		X"BD",X"A6",X"CE",X"B6",X"57",X"C7",X"44",X"84",X"03",X"8B",X"28",X"A7",X"41",X"20",X"26",X"C6",
		X"3E",X"D7",X"F6",X"20",X"04",X"C6",X"36",X"D7",X"F6",X"B6",X"57",X"C7",X"44",X"84",X"01",X"9B",
		X"F6",X"A7",X"41",X"20",X"10",X"10",X"8E",X"F6",X"4E",X"B6",X"57",X"C7",X"44",X"44",X"44",X"84",
		X"03",X"A6",X"A6",X"A7",X"41",X"A6",X"43",X"E6",X"0C",X"E3",X"06",X"F3",X"57",X"C0",X"A7",X"43",
		X"E7",X"0C",X"A6",X"C4",X"E6",X"0D",X"E3",X"08",X"F3",X"57",X"C2",X"A7",X"C4",X"E7",X"0D",X"7E",
		X"A5",X"83",X"A6",X"43",X"8B",X"04",X"81",X"08",X"25",X"1D",X"A6",X"C4",X"8B",X"10",X"81",X"10",
		X"25",X"15",X"39",X"A6",X"43",X"8B",X"04",X"81",X"08",X"25",X"09",X"A6",X"C4",X"8B",X"10",X"81",
		X"10",X"25",X"01",X"39",X"7A",X"52",X"34",X"4F",X"A7",X"84",X"A7",X"43",X"39",X"7A",X"54",X"40",
		X"27",X"01",X"39",X"4F",X"B7",X"51",X"FB",X"B7",X"51",X"FF",X"39",X"10",X"8E",X"F6",X"52",X"58",
		X"58",X"31",X"A5",X"EC",X"A1",X"B7",X"51",X"F9",X"F7",X"51",X"FA",X"EC",X"A4",X"B7",X"51",X"FD",
		X"F7",X"51",X"FE",X"CC",X"18",X"28",X"B7",X"51",X"FB",X"F7",X"51",X"FF",X"CC",X"13",X"13",X"B7",
		X"51",X"F8",X"F7",X"51",X"FC",X"86",X"60",X"B7",X"54",X"40",X"BD",X"92",X"8F",X"39",X"DC",X"ED",
		X"34",X"10",X"CB",X"08",X"D7",X"F6",X"5F",X"A0",X"43",X"24",X"03",X"C6",X"02",X"40",X"DD",X"F7",
		X"C6",X"01",X"A6",X"C4",X"8B",X"08",X"90",X"F6",X"24",X"02",X"5F",X"40",X"DA",X"F8",X"D7",X"F8",
		X"5A",X"C1",X"02",X"D6",X"F7",X"24",X"02",X"1E",X"89",X"54",X"54",X"54",X"54",X"D7",X"F6",X"84",
		X"F0",X"9B",X"F6",X"8E",X"F6",X"EA",X"E6",X"86",X"96",X"F8",X"8E",X"F6",X"66",X"EB",X"86",X"35",
		X"90",X"34",X"10",X"D7",X"F6",X"C4",X"3F",X"26",X"15",X"0F",X"3B",X"0F",X"3D",X"08",X"F6",X"59",
		X"08",X"F6",X"59",X"8E",X"F7",X"EA",X"EC",X"85",X"D7",X"3A",X"97",X"3C",X"35",X"90",X"0F",X"3A",
		X"0F",X"3C",X"8E",X"F7",X"6A",X"30",X"85",X"A6",X"84",X"E6",X"88",X"40",X"08",X"F6",X"25",X"0B",
		X"08",X"F6",X"24",X"15",X"1E",X"89",X"50",X"03",X"3A",X"20",X"0E",X"1E",X"89",X"40",X"03",X"3C",
		X"08",X"F6",X"25",X"05",X"1E",X"89",X"40",X"03",X"3A",X"D7",X"3B",X"97",X"3D",X"35",X"90",X"DD",
		X"D6",X"DC",X"3A",X"2A",X"04",X"4F",X"5F",X"93",X"3A",X"DD",X"F6",X"0D",X"F6",X"27",X"04",X"DC",
		X"D6",X"20",X"10",X"0F",X"F9",X"96",X"F7",X"D6",X"D7",X"3D",X"97",X"FA",X"96",X"F7",X"D6",X"D6",
		X"3D",X"D3",X"F9",X"DD",X"F6",X"0D",X"3A",X"2A",X"04",X"4F",X"5F",X"93",X"F6",X"DD",X"3A",X"DC",
		X"3C",X"2A",X"04",X"4F",X"5F",X"93",X"3C",X"DD",X"F6",X"0D",X"F6",X"27",X"04",X"DC",X"D6",X"20",
		X"10",X"0F",X"F9",X"96",X"F7",X"D6",X"D7",X"3D",X"97",X"FA",X"96",X"F7",X"D6",X"D6",X"3D",X"D3",
		X"F9",X"DD",X"F6",X"0D",X"3C",X"2A",X"04",X"4F",X"5F",X"93",X"F6",X"DD",X"3C",X"39",X"96",X"A7",
		X"10",X"27",X"00",X"72",X"96",X"9C",X"10",X"26",X"00",X"6C",X"B6",X"57",X"C7",X"44",X"44",X"44",
		X"44",X"84",X"0F",X"97",X"F6",X"A6",X"0F",X"84",X"0F",X"91",X"F6",X"10",X"26",X"00",X"57",X"D6",
		X"9D",X"DB",X"9D",X"D7",X"F6",X"A6",X"43",X"80",X"80",X"9B",X"9D",X"91",X"F6",X"24",X"0A",X"A6",
		X"C4",X"80",X"78",X"9B",X"9D",X"91",X"F6",X"25",X"3D",X"BD",X"A5",X"DE",X"D7",X"CB",X"CB",X"80",
		X"D7",X"F6",X"B6",X"52",X"41",X"90",X"F6",X"9B",X"A2",X"D6",X"A2",X"DB",X"A2",X"D7",X"F6",X"91",
		X"F6",X"25",X"23",X"10",X"8E",X"51",X"D4",X"10",X"9F",X"5C",X"10",X"8E",X"53",X"B0",X"86",X"06",
		X"97",X"32",X"A6",X"A4",X"10",X"27",X"00",X"0F",X"31",X"A8",X"10",X"CC",X"00",X"04",X"D3",X"5C",
		X"DD",X"5C",X"0A",X"32",X"26",X"EC",X"39",X"96",X"9B",X"97",X"9C",X"86",X"FF",X"A7",X"A4",X"D6",
		X"CB",X"BD",X"A6",X"21",X"CC",X"01",X"90",X"BD",X"A6",X"6F",X"DC",X"3A",X"ED",X"24",X"DC",X"3C",
		X"ED",X"26",X"CC",X"00",X"00",X"ED",X"28",X"A7",X"23",X"10",X"9E",X"5C",X"A6",X"43",X"A7",X"23",
		X"A6",X"C4",X"A7",X"A4",X"CC",X"1F",X"40",X"ED",X"21",X"7E",X"92",X"06",X"8E",X"53",X"B0",X"CE",
		X"51",X"D4",X"A6",X"84",X"27",X"2E",X"4C",X"27",X"05",X"4C",X"27",X"28",X"20",X"31",X"A6",X"43",
		X"E6",X"08",X"E3",X"04",X"F3",X"57",X"C0",X"A7",X"43",X"E7",X"08",X"8B",X"03",X"81",X"07",X"25",
		X"1E",X"A6",X"C4",X"E6",X"09",X"E3",X"06",X"F3",X"57",X"C2",X"A7",X"C4",X"E7",X"09",X"8B",X"03",
		X"81",X"07",X"25",X"0B",X"30",X"88",X"10",X"33",X"44",X"8C",X"54",X"40",X"25",X"C4",X"39",X"4F",
		X"A7",X"84",X"A7",X"43",X"20",X"EE",X"8E",X"BD",X"5E",X"C6",X"06",X"A6",X"80",X"AB",X"80",X"5A",
		X"26",X"FB",X"81",X"1B",X"27",X"0A",X"B6",X"57",X"C8",X"88",X"01",X"B7",X"57",X"C8",X"20",X"0F",
		X"B6",X"B5",X"62",X"81",X"1B",X"27",X"08",X"B6",X"57",X"C8",X"88",X"01",X"B7",X"57",X"C8",X"B6",
		X"55",X"20",X"26",X"52",X"8E",X"F7",X"FF",X"0F",X"F7",X"EC",X"84",X"83",X"00",X"07",X"93",X"1A",
		X"84",X"07",X"26",X"16",X"D7",X"F8",X"EC",X"02",X"93",X"1C",X"84",X"07",X"26",X"0C",X"D7",X"F9",
		X"96",X"F7",X"CE",X"44",X"24",X"A6",X"C6",X"27",X"0B",X"39",X"0C",X"F7",X"30",X"04",X"8C",X"F8",
		X"1F",X"25",X"D6",X"39",X"CE",X"55",X"20",X"DC",X"F8",X"B7",X"52",X"33",X"F7",X"52",X"30",X"CC",
		X"FF",X"40",X"FD",X"52",X"31",X"EC",X"84",X"ED",X"43",X"EC",X"02",X"ED",X"45",X"96",X"F7",X"A7",
		X"41",X"6F",X"42",X"6A",X"C4",X"39",X"8E",X"55",X"20",X"CE",X"52",X"30",X"A6",X"84",X"4C",X"26",
		X"66",X"EC",X"03",X"83",X"00",X"07",X"93",X"1A",X"84",X"07",X"26",X"48",X"D7",X"F6",X"EC",X"05",
		X"93",X"1C",X"84",X"07",X"26",X"3E",X"E7",X"C4",X"96",X"F6",X"A7",X"43",X"A6",X"02",X"81",X"02",
		X"27",X"1C",X"A6",X"84",X"4C",X"26",X"16",X"E6",X"02",X"27",X"12",X"A6",X"07",X"27",X"0E",X"6A",
		X"07",X"44",X"44",X"84",X"07",X"10",X"8E",X"F7",X"EF",X"A6",X"A6",X"A7",X"41",X"39",X"A6",X"07",
		X"27",X"12",X"6A",X"07",X"A6",X"07",X"44",X"44",X"44",X"84",X"07",X"10",X"8E",X"F7",X"F7",X"A6",
		X"A6",X"A7",X"41",X"39",X"A6",X"02",X"27",X"0A",X"10",X"8E",X"44",X"24",X"A6",X"01",X"C6",X"FF",
		X"E7",X"A6",X"6F",X"43",X"6F",X"84",X"39",X"81",X"78",X"24",X"19",X"6A",X"84",X"27",X"E5",X"A6",
		X"84",X"44",X"44",X"44",X"10",X"8E",X"F8",X"1F",X"A6",X"A6",X"A7",X"41",X"86",X"40",X"A7",X"42",
		X"7E",X"A8",X"51",X"39",X"86",X"28",X"A7",X"84",X"C6",X"03",X"BD",X"A5",X"AB",X"CC",X"06",X"08",
		X"BD",X"8F",X"0C",X"7E",X"A8",X"51",X"FC",X"52",X"35",X"10",X"83",X"FF",X"FF",X"26",X"1A",X"8E",
		X"C2",X"4D",X"C6",X"1B",X"A6",X"80",X"AB",X"80",X"5A",X"26",X"FB",X"81",X"34",X"27",X"0A",X"86",
		X"01",X"B7",X"57",X"C8",X"7F",X"57",X"D0",X"20",X"11",X"B6",X"83",X"61",X"81",X"1B",X"27",X"0A",
		X"CC",X"00",X"52",X"BD",X"8F",X"0C",X"5C",X"BD",X"8F",X"0C",X"B6",X"57",X"C7",X"84",X"03",X"26",
		X"2C",X"FC",X"57",X"C0",X"58",X"49",X"58",X"49",X"58",X"49",X"58",X"49",X"DD",X"F6",X"58",X"49",
		X"D3",X"F6",X"40",X"8B",X"80",X"97",X"ED",X"FC",X"57",X"C2",X"58",X"49",X"58",X"49",X"58",X"49",
		X"58",X"49",X"DD",X"F6",X"58",X"49",X"D3",X"F6",X"40",X"8B",X"78",X"97",X"EE",X"39",X"CE",X"F8",
		X"35",X"8E",X"55",X"30",X"86",X"18",X"97",X"F6",X"86",X"FF",X"97",X"F7",X"8D",X"1C",X"4F",X"F6",
		X"57",X"D4",X"26",X"04",X"0F",X"2E",X"86",X"FF",X"97",X"F7",X"CE",X"F8",X"DD",X"B6",X"57",X"D6",
		X"48",X"EE",X"C6",X"8E",X"56",X"B0",X"86",X"08",X"97",X"F6",X"EC",X"C4",X"ED",X"04",X"EC",X"42",
		X"ED",X"06",X"EC",X"44",X"ED",X"08",X"A6",X"46",X"A7",X"01",X"96",X"F7",X"A7",X"02",X"CC",X"00",
		X"00",X"ED",X"0C",X"6F",X"0A",X"30",X"88",X"10",X"33",X"47",X"0A",X"F6",X"26",X"DC",X"8E",X"BD",
		X"5E",X"C6",X"06",X"A6",X"80",X"AB",X"80",X"5A",X"26",X"FB",X"81",X"1B",X"27",X"0A",X"86",X"01",
		X"B7",X"57",X"C8",X"7F",X"57",X"D0",X"20",X"20",X"B6",X"A7",X"E4",X"81",X"1B",X"27",X"0A",X"B6",
		X"57",X"C8",X"88",X"01",X"B7",X"57",X"C8",X"20",X"0F",X"B6",X"B5",X"62",X"81",X"1B",X"27",X"08",
		X"B6",X"57",X"C8",X"88",X"01",X"B7",X"57",X"C8",X"39",X"8E",X"55",X"30",X"86",X"20",X"97",X"7A",
		X"A6",X"02",X"27",X"18",X"EC",X"04",X"93",X"1A",X"84",X"07",X"26",X"0D",X"EC",X"06",X"93",X"1C",
		X"84",X"07",X"26",X"05",X"BD",X"AA",X"BB",X"20",X"03",X"BD",X"AA",X"07",X"0A",X"7A",X"10",X"27",
		X"00",X"F4",X"30",X"88",X"10",X"20",X"D9",X"A6",X"0A",X"26",X"03",X"BD",X"AA",X"44",X"6A",X"0A",
		X"A6",X"0B",X"10",X"8E",X"FB",X"94",X"E6",X"08",X"59",X"24",X"04",X"10",X"8E",X"FB",X"B8",X"31",
		X"A6",X"E6",X"0C",X"EB",X"21",X"E7",X"0C",X"C6",X"00",X"E9",X"A4",X"1D",X"E3",X"04",X"84",X"07",
		X"ED",X"04",X"E6",X"0D",X"EB",X"23",X"E7",X"0D",X"C6",X"00",X"E9",X"22",X"1D",X"E3",X"06",X"84",
		X"07",X"ED",X"06",X"39",X"A6",X"08",X"2B",X"5F",X"10",X"8E",X"FA",X"41",X"48",X"10",X"AE",X"A6",
		X"A6",X"09",X"6C",X"09",X"A6",X"A6",X"81",X"FF",X"27",X"1D",X"81",X"FE",X"27",X"3F",X"81",X"FD",
		X"27",X"27",X"81",X"FC",X"27",X"2D",X"1F",X"89",X"84",X"0F",X"48",X"48",X"48",X"48",X"A7",X"0A",
		X"C4",X"F0",X"54",X"54",X"E7",X"0B",X"39",X"86",X"01",X"A7",X"09",X"A6",X"A4",X"20",X"E7",X"A6",
		X"08",X"8B",X"80",X"A7",X"08",X"6C",X"09",X"20",X"BB",X"A6",X"08",X"8B",X"08",X"A7",X"08",X"6F",
		X"09",X"20",X"B1",X"A6",X"08",X"80",X"08",X"A7",X"08",X"6F",X"09",X"20",X"A7",X"A6",X"08",X"8B",
		X"80",X"A7",X"08",X"6A",X"09",X"6A",X"09",X"10",X"8E",X"FA",X"41",X"48",X"10",X"AE",X"A6",X"A6",
		X"09",X"81",X"FF",X"27",X"CA",X"6A",X"09",X"A6",X"A6",X"20",X"AB",X"CE",X"54",X"A0",X"86",X"08",
		X"97",X"F6",X"A6",X"C4",X"27",X"0C",X"0A",X"F6",X"27",X"05",X"33",X"C8",X"10",X"20",X"F3",X"7E",
		X"AA",X"07",X"6A",X"C4",X"EC",X"04",X"ED",X"44",X"EC",X"06",X"ED",X"46",X"EC",X"08",X"ED",X"48",
		X"EC",X"0A",X"ED",X"4A",X"EC",X"0C",X"ED",X"4C",X"A6",X"01",X"27",X"02",X"0C",X"DA",X"A7",X"41",
		X"4F",X"A7",X"42",X"A7",X"02",X"39",X"8E",X"54",X"A0",X"CE",X"52",X"10",X"A6",X"84",X"10",X"27",
		X"00",X"A1",X"4C",X"10",X"26",X"00",X"A9",X"BD",X"AA",X"07",X"EC",X"04",X"93",X"1A",X"84",X"07",
		X"26",X"36",X"D7",X"F6",X"EC",X"06",X"93",X"1C",X"84",X"07",X"26",X"2C",X"E7",X"C4",X"96",X"F6",
		X"A7",X"43",X"BD",X"AC",X"4E",X"A6",X"02",X"10",X"8E",X"F8",X"24",X"E6",X"01",X"27",X"02",X"8B",
		X"04",X"A6",X"A6",X"A7",X"41",X"10",X"8E",X"F8",X"2C",X"B6",X"57",X"C7",X"44",X"44",X"44",X"44",
		X"84",X"03",X"A6",X"A6",X"A7",X"42",X"20",X"5B",X"10",X"8E",X"55",X"30",X"86",X"20",X"97",X"F6",
		X"6D",X"22",X"27",X"0B",X"0A",X"F6",X"27",X"05",X"31",X"A8",X"10",X"20",X"F3",X"20",X"44",X"6A",
		X"22",X"EC",X"04",X"ED",X"24",X"EC",X"06",X"ED",X"26",X"EC",X"08",X"ED",X"28",X"EC",X"0A",X"ED",
		X"2A",X"EC",X"0C",X"ED",X"2C",X"A6",X"01",X"27",X"02",X"0A",X"DA",X"A7",X"21",X"4F",X"A7",X"84",
		X"A7",X"23",X"A6",X"02",X"27",X"1D",X"81",X"03",X"24",X"19",X"10",X"8E",X"54",X"10",X"86",X"03",
		X"A7",X"7F",X"A6",X"A4",X"81",X"FE",X"27",X"09",X"31",X"A8",X"10",X"6A",X"7F",X"26",X"F3",X"20",
		X"02",X"6F",X"A4",X"30",X"88",X"10",X"33",X"44",X"8C",X"55",X"20",X"10",X"25",X"FF",X"4D",X"39",
		X"81",X"78",X"24",X"46",X"6A",X"84",X"27",X"28",X"A6",X"84",X"44",X"44",X"44",X"10",X"8E",X"F8",
		X"30",X"A6",X"A6",X"A7",X"41",X"86",X"40",X"A7",X"42",X"EC",X"04",X"93",X"1A",X"84",X"07",X"26",
		X"0F",X"E7",X"43",X"EC",X"06",X"93",X"1C",X"84",X"07",X"26",X"05",X"E7",X"C4",X"7E",X"AB",X"A3",
		X"A6",X"01",X"26",X"08",X"CC",X"06",X"02",X"BD",X"8F",X"0C",X"20",X"06",X"CC",X"06",X"04",X"BD",
		X"8F",X"0C",X"4F",X"A7",X"43",X"A7",X"84",X"7E",X"AB",X"A3",X"BD",X"92",X"16",X"86",X"28",X"A7",
		X"84",X"A6",X"01",X"27",X"24",X"0A",X"DA",X"0C",X"2E",X"96",X"2E",X"81",X"08",X"26",X"1A",X"B6",
		X"54",X"60",X"4A",X"2B",X"06",X"B6",X"54",X"6D",X"26",X"01",X"39",X"CC",X"06",X"09",X"BD",X"8F",
		X"0C",X"C6",X"04",X"BD",X"A5",X"AB",X"7A",X"57",X"D4",X"A6",X"02",X"27",X"87",X"81",X"03",X"24",
		X"83",X"10",X"8E",X"54",X"10",X"86",X"03",X"97",X"F6",X"A6",X"A4",X"81",X"FE",X"27",X"0A",X"31",
		X"A8",X"10",X"0A",X"F6",X"26",X"F3",X"7E",X"AB",X"B4",X"6F",X"A4",X"7E",X"AB",X"B4",X"A6",X"02",
		X"26",X"68",X"B6",X"57",X"C9",X"81",X"07",X"26",X"60",X"A6",X"01",X"26",X"49",X"96",X"A7",X"26",
		X"58",X"B6",X"57",X"C7",X"49",X"49",X"49",X"49",X"84",X"0F",X"97",X"F6",X"A6",X"0F",X"84",X"0F",
		X"91",X"F6",X"26",X"45",X"D6",X"9D",X"DB",X"9D",X"D7",X"F6",X"A6",X"43",X"80",X"80",X"9B",X"9D",
		X"91",X"F6",X"22",X"0A",X"A6",X"C4",X"80",X"78",X"9B",X"9D",X"91",X"F6",X"23",X"2B",X"BD",X"A5",
		X"DE",X"CB",X"80",X"D7",X"F6",X"B6",X"52",X"41",X"90",X"F6",X"9B",X"A2",X"D6",X"A2",X"DB",X"A2",
		X"D7",X"F6",X"91",X"F6",X"25",X"13",X"10",X"8E",X"54",X"10",X"86",X"03",X"97",X"F6",X"A6",X"A4",
		X"27",X"18",X"31",X"A8",X"10",X"0A",X"F6",X"26",X"F5",X"39",X"6A",X"0E",X"27",X"01",X"39",X"81",
		X"02",X"25",X"0B",X"81",X"03",X"26",X"0E",X"6F",X"02",X"39",X"86",X"FE",X"A7",X"A4",X"6C",X"02",
		X"86",X"08",X"A7",X"0E",X"39",X"10",X"8E",X"51",X"EC",X"10",X"9F",X"CE",X"10",X"8E",X"54",X"10",
		X"86",X"03",X"97",X"F6",X"A6",X"A4",X"81",X"FE",X"27",X"0F",X"31",X"A8",X"10",X"CC",X"00",X"04",
		X"D3",X"CE",X"DD",X"CE",X"0A",X"F6",X"26",X"EC",X"39",X"6C",X"A4",X"34",X"20",X"10",X"9E",X"CE",
		X"CC",X"1F",X"40",X"ED",X"21",X"A6",X"C4",X"E6",X"43",X"A7",X"A4",X"E7",X"23",X"35",X"20",X"BD",
		X"A5",X"DE",X"BD",X"A6",X"21",X"CC",X"01",X"90",X"BD",X"A6",X"6F",X"DC",X"3A",X"ED",X"24",X"DC",
		X"3C",X"ED",X"26",X"CC",X"00",X"00",X"ED",X"28",X"6C",X"02",X"86",X"10",X"A7",X"0E",X"7E",X"92",
		X"06",X"8E",X"52",X"40",X"CE",X"51",X"78",X"CC",X"78",X"08",X"ED",X"C4",X"CC",X"40",X"80",X"ED",
		X"42",X"86",X"FF",X"A7",X"84",X"86",X"C0",X"A7",X"01",X"A7",X"02",X"5F",X"E7",X"0F",X"30",X"88",
		X"10",X"5C",X"C1",X"2F",X"25",X"F6",X"39",X"8E",X"52",X"40",X"CE",X"51",X"78",X"A6",X"84",X"4C",
		X"10",X"26",X"00",X"5E",X"BD",X"85",X"2E",X"84",X"0F",X"81",X"00",X"27",X"25",X"10",X"8E",X"FB",
		X"FC",X"31",X"A6",X"A6",X"A4",X"A7",X"02",X"A0",X"01",X"27",X"17",X"C6",X"03",X"81",X"80",X"25",
		X"01",X"50",X"EB",X"01",X"E7",X"01",X"E0",X"02",X"CB",X"02",X"C1",X"05",X"22",X"04",X"A6",X"02",
		X"A7",X"01",X"10",X"8E",X"FB",X"DC",X"A6",X"01",X"8B",X"04",X"1F",X"89",X"44",X"44",X"44",X"A6",
		X"A6",X"A7",X"41",X"86",X"00",X"59",X"24",X"02",X"86",X"40",X"A7",X"42",X"E6",X"01",X"BD",X"A6",
		X"21",X"CC",X"00",X"00",X"93",X"3A",X"FD",X"57",X"C0",X"CC",X"00",X"00",X"93",X"3C",X"FD",X"57",
		X"C2",X"39",X"81",X"78",X"24",X"35",X"6A",X"84",X"10",X"27",X"00",X"7A",X"A6",X"84",X"44",X"44",
		X"48",X"10",X"8E",X"FC",X"07",X"10",X"AE",X"A6",X"C6",X"40",X"A6",X"A0",X"B7",X"51",X"79",X"F7",
		X"51",X"7A",X"A6",X"A0",X"B7",X"51",X"7D",X"F7",X"51",X"7E",X"A6",X"A0",X"B7",X"51",X"81",X"F7",
		X"51",X"82",X"A6",X"A4",X"B7",X"51",X"85",X"F7",X"51",X"86",X"39",X"BD",X"91",X"EF",X"BD",X"92",
		X"5D",X"C6",X"78",X"F7",X"51",X"7B",X"F7",X"51",X"83",X"CB",X"10",X"F7",X"51",X"7F",X"F7",X"51",
		X"87",X"C6",X"70",X"F7",X"51",X"78",X"F7",X"51",X"7C",X"CB",X"10",X"F7",X"51",X"80",X"F7",X"51",
		X"84",X"86",X"34",X"A7",X"84",X"7F",X"51",X"8B",X"7F",X"51",X"8F",X"7F",X"51",X"93",X"7F",X"52",
		X"80",X"7F",X"52",X"90",X"7F",X"52",X"A0",X"7F",X"52",X"B8",X"7F",X"52",X"C8",X"7F",X"51",X"9C",
		X"7F",X"51",X"A0",X"7E",X"AD",X"C2",X"7F",X"51",X"7B",X"7F",X"51",X"7F",X"7F",X"51",X"83",X"7F",
		X"51",X"87",X"6C",X"84",X"0C",X"CC",X"96",X"CC",X"81",X"50",X"25",X"02",X"6F",X"84",X"39",X"B6",
		X"52",X"40",X"4C",X"10",X"26",X"01",X"31",X"BD",X"85",X"2E",X"48",X"48",X"48",X"79",X"57",X"BF",
		X"48",X"79",X"57",X"BE",X"96",X"EF",X"26",X"0F",X"B6",X"57",X"BE",X"84",X"07",X"81",X"01",X"26",
		X"60",X"86",X"0C",X"97",X"EF",X"20",X"09",X"4A",X"97",X"EF",X"27",X"04",X"81",X"06",X"26",X"51",
		X"8E",X"52",X"50",X"CE",X"51",X"7C",X"A6",X"84",X"26",X"3D",X"BD",X"92",X"02",X"4F",X"5F",X"B3",
		X"57",X"C0",X"58",X"49",X"58",X"49",X"ED",X"03",X"8B",X"80",X"ED",X"07",X"A7",X"43",X"4F",X"5F",
		X"B3",X"57",X"C2",X"58",X"49",X"58",X"49",X"ED",X"05",X"8B",X"78",X"ED",X"09",X"A7",X"C4",X"6A",
		X"84",X"B6",X"52",X"41",X"5F",X"ED",X"01",X"8B",X"04",X"84",X"F8",X"44",X"44",X"10",X"8E",X"FC",
		X"55",X"EC",X"A6",X"ED",X"41",X"20",X"0A",X"30",X"88",X"10",X"33",X"44",X"8C",X"52",X"B0",X"25",
		X"B5",X"B6",X"57",X"BF",X"84",X"07",X"81",X"01",X"26",X"49",X"8E",X"52",X"C0",X"CE",X"51",X"98",
		X"5F",X"A6",X"10",X"4A",X"81",X"FF",X"59",X"A6",X"84",X"4A",X"81",X"FF",X"59",X"A6",X"18",X"48",
		X"59",X"A6",X"08",X"48",X"59",X"10",X"8E",X"FC",X"95",X"A6",X"A5",X"27",X"26",X"2A",X"04",X"30",
		X"10",X"33",X"5C",X"BD",X"92",X"3E",X"6F",X"88",X"20",X"6A",X"84",X"86",X"80",X"A7",X"43",X"CC",
		X"78",X"FF",X"ED",X"C4",X"B6",X"52",X"41",X"A7",X"01",X"6C",X"4A",X"6F",X"09",X"A6",X"08",X"26",
		X"02",X"6F",X"0A",X"8E",X"52",X"50",X"CE",X"51",X"7C",X"A6",X"84",X"27",X"29",X"4C",X"26",X"32",
		X"EC",X"03",X"E3",X"07",X"F3",X"57",X"C0",X"ED",X"07",X"8B",X"03",X"81",X"07",X"25",X"43",X"80",
		X"03",X"A7",X"43",X"EC",X"05",X"E3",X"09",X"F3",X"57",X"C2",X"ED",X"09",X"8B",X"03",X"81",X"07",
		X"25",X"30",X"80",X"03",X"A7",X"C4",X"30",X"88",X"10",X"33",X"44",X"8C",X"52",X"B0",X"26",X"C9",
		X"20",X"26",X"81",X"78",X"23",X"0E",X"86",X"0C",X"A7",X"84",X"CC",X"1E",X"48",X"ED",X"41",X"BD",
		X"91",X"FE",X"20",X"E2",X"6A",X"84",X"27",X"0A",X"A6",X"84",X"85",X"03",X"26",X"D8",X"6C",X"42",
		X"20",X"D4",X"6F",X"84",X"6F",X"43",X"20",X"CE",X"8E",X"52",X"C8",X"CE",X"51",X"A0",X"A6",X"84",
		X"27",X"56",X"10",X"AE",X"05",X"A6",X"23",X"10",X"8C",X"52",X"00",X"26",X"02",X"8B",X"08",X"A7",
		X"43",X"8B",X"08",X"81",X"10",X"23",X"3B",X"A6",X"A4",X"10",X"8C",X"52",X"00",X"26",X"02",X"8B",
		X"08",X"A7",X"C4",X"4A",X"81",X"EF",X"24",X"2A",X"A6",X"18",X"26",X"2C",X"6A",X"01",X"26",X"12",
		X"10",X"8C",X"52",X"30",X"26",X"1C",X"86",X"02",X"B7",X"55",X"22",X"86",X"20",X"B7",X"55",X"27",
		X"20",X"10",X"A6",X"01",X"80",X"30",X"23",X"10",X"44",X"25",X"01",X"40",X"AB",X"43",X"A7",X"43",
		X"20",X"06",X"6F",X"84",X"6F",X"43",X"6A",X"04",X"30",X"10",X"33",X"5C",X"8C",X"52",X"B8",X"27",
		X"9D",X"8E",X"52",X"C0",X"CE",X"51",X"98",X"A6",X"84",X"10",X"27",X"00",X"B8",X"4C",X"10",X"26",
		X"00",X"DE",X"E6",X"08",X"26",X"2D",X"A6",X"43",X"A8",X"C4",X"E6",X"43",X"C0",X"50",X"C1",X"60",
		X"24",X"36",X"E6",X"C4",X"C0",X"48",X"C1",X"60",X"24",X"2E",X"84",X"3F",X"97",X"F6",X"4F",X"E6",
		X"43",X"58",X"46",X"E6",X"C4",X"CB",X"08",X"58",X"46",X"88",X"80",X"2B",X"02",X"88",X"40",X"9A",
		X"F6",X"20",X"15",X"10",X"AE",X"0D",X"A6",X"23",X"E6",X"A4",X"10",X"8C",X"52",X"00",X"26",X"03",
		X"C3",X"08",X"08",X"BD",X"A5",X"E0",X"1F",X"98",X"6A",X"88",X"20",X"26",X"03",X"6C",X"88",X"20",
		X"E6",X"88",X"20",X"50",X"59",X"59",X"59",X"C4",X"07",X"A0",X"01",X"2A",X"01",X"50",X"EB",X"01",
		X"E7",X"01",X"BD",X"A6",X"21",X"CC",X"02",X"20",X"BD",X"A6",X"6F",X"DC",X"3A",X"ED",X"04",X"DC",
		X"3C",X"ED",X"06",X"A6",X"43",X"E6",X"02",X"E3",X"04",X"F3",X"57",X"C0",X"A7",X"43",X"E7",X"02",
		X"8B",X"F9",X"81",X"02",X"23",X"3B",X"A6",X"C4",X"E6",X"03",X"E3",X"06",X"F3",X"57",X"C2",X"A7",
		X"C4",X"E7",X"03",X"8B",X"02",X"81",X"02",X"23",X"28",X"A6",X"84",X"2A",X"18",X"10",X"8E",X"FC",
		X"A5",X"A6",X"0A",X"27",X"03",X"31",X"A8",X"20",X"A6",X"01",X"8B",X"08",X"84",X"F0",X"44",X"44",
		X"44",X"EC",X"A6",X"ED",X"41",X"30",X"10",X"33",X"5C",X"8C",X"52",X"B0",X"10",X"27",X"FF",X"37",
		X"39",X"6F",X"08",X"6F",X"4B",X"10",X"AE",X"0B",X"6A",X"0C",X"10",X"8C",X"55",X"20",X"26",X"0A",
		X"86",X"02",X"B7",X"55",X"22",X"86",X"20",X"B7",X"55",X"27",X"6F",X"84",X"6F",X"43",X"20",X"D5",
		X"81",X"78",X"23",X"0A",X"6F",X"08",X"6F",X"4B",X"6A",X"0C",X"86",X"11",X"A7",X"84",X"6A",X"84",
		X"27",X"E8",X"A6",X"84",X"85",X"03",X"26",X"BD",X"10",X"8E",X"F4",X"D3",X"44",X"44",X"A6",X"A6",
		X"A7",X"41",X"7E",X"B0",X"83",X"B6",X"52",X"40",X"4C",X"27",X"01",X"39",X"8E",X"52",X"50",X"A6",
		X"84",X"4C",X"26",X"79",X"A6",X"01",X"8B",X"04",X"84",X"78",X"44",X"44",X"CE",X"FC",X"E5",X"EC",
		X"C6",X"DD",X"F6",X"48",X"58",X"DD",X"F8",X"CE",X"52",X"F0",X"10",X"8E",X"51",X"A4",X"86",X"0C",
		X"F6",X"52",X"34",X"FA",X"54",X"60",X"26",X"01",X"44",X"97",X"FA",X"A6",X"C4",X"4C",X"26",X"2A",
		X"A6",X"07",X"A0",X"23",X"9B",X"F6",X"91",X"F8",X"22",X"20",X"A6",X"09",X"A0",X"A4",X"9B",X"F7",
		X"91",X"F9",X"22",X"16",X"86",X"78",X"11",X"83",X"53",X"50",X"25",X"4A",X"F6",X"54",X"60",X"27",
		X"38",X"F6",X"54",X"6D",X"2A",X"40",X"A7",X"84",X"20",X"23",X"31",X"24",X"33",X"C8",X"10",X"0A",
		X"FA",X"26",X"C8",X"B6",X"54",X"60",X"4C",X"26",X"14",X"A6",X"07",X"B0",X"52",X"03",X"81",X"10",
		X"22",X"0B",X"86",X"78",X"E6",X"09",X"F0",X"52",X"00",X"C1",X"10",X"23",X"D9",X"30",X"88",X"10",
		X"8C",X"52",X"B0",X"10",X"26",X"FF",X"78",X"20",X"13",X"E6",X"43",X"C0",X"07",X"27",X"07",X"5A",
		X"26",X"C4",X"6A",X"41",X"26",X"C0",X"A7",X"C4",X"60",X"84",X"20",X"E1",X"8E",X"52",X"C8",X"A6",
		X"84",X"AA",X"18",X"27",X"0A",X"30",X"10",X"A6",X"84",X"AA",X"18",X"10",X"26",X"00",X"E4",X"4F",
		X"5F",X"B3",X"57",X"C2",X"58",X"49",X"58",X"49",X"58",X"49",X"58",X"49",X"DD",X"F6",X"58",X"49",
		X"D3",X"F6",X"8B",X"88",X"97",X"F8",X"4F",X"5F",X"B3",X"57",X"C0",X"58",X"49",X"58",X"49",X"58",
		X"49",X"58",X"49",X"DD",X"F6",X"58",X"49",X"D3",X"F6",X"8B",X"90",X"97",X"F9",X"0F",X"FB",X"CE",
		X"53",X"50",X"B6",X"52",X"34",X"27",X"72",X"10",X"8E",X"51",X"BC",X"86",X"06",X"97",X"FA",X"A6",
		X"C4",X"4C",X"26",X"5C",X"11",X"83",X"54",X"A0",X"24",X"06",X"A6",X"43",X"81",X"07",X"27",X"50",
		X"DC",X"F8",X"E0",X"23",X"C1",X"20",X"22",X"48",X"A0",X"A4",X"81",X"20",X"22",X"42",X"86",X"F3",
		X"8C",X"52",X"C8",X"27",X"02",X"86",X"13",X"11",X"A3",X"86",X"27",X"34",X"11",X"83",X"55",X"20",
		X"26",X"0D",X"A6",X"42",X"26",X"2A",X"6C",X"42",X"86",X"20",X"A7",X"47",X"BD",X"92",X"94",X"6A",
		X"84",X"86",X"50",X"D6",X"FB",X"ED",X"01",X"EF",X"03",X"10",X"AF",X"05",X"E6",X"07",X"CB",X"02",
		X"58",X"58",X"4F",X"C3",X"51",X"79",X"1F",X"01",X"CC",X"FE",X"06",X"ED",X"84",X"7E",X"92",X"1E",
		X"31",X"24",X"33",X"C8",X"10",X"0A",X"FA",X"26",X"96",X"11",X"83",X"54",X"70",X"27",X"34",X"22",
		X"0E",X"CE",X"54",X"A0",X"10",X"8E",X"52",X"10",X"0C",X"FB",X"86",X"09",X"7E",X"B2",X"0D",X"CE",
		X"54",X"60",X"A6",X"C4",X"4C",X"26",X"1C",X"10",X"8E",X"52",X"00",X"DC",X"F8",X"E0",X"23",X"C0",
		X"08",X"C1",X"20",X"22",X"0E",X"0C",X"FA",X"0F",X"FB",X"A0",X"A4",X"80",X"08",X"81",X"20",X"10",
		X"23",X"FF",X"7B",X"8E",X"52",X"C0",X"CE",X"51",X"98",X"A6",X"84",X"A4",X"08",X"4C",X"26",X"2E",
		X"A6",X"98",X"0B",X"4C",X"26",X"28",X"A6",X"43",X"E6",X"C4",X"EE",X"0D",X"11",X"83",X"52",X"00",
		X"26",X"03",X"83",X"08",X"08",X"A0",X"43",X"2A",X"01",X"40",X"97",X"F6",X"E0",X"C4",X"2A",X"01",
		X"50",X"DB",X"F6",X"C1",X"08",X"22",X"07",X"86",X"78",X"A7",X"84",X"A7",X"98",X"0B",X"30",X"10",
		X"CE",X"51",X"94",X"8C",X"52",X"B0",X"27",X"C1",X"39",X"B6",X"57",X"C6",X"8E",X"FD",X"3D",X"48",
		X"6E",X"96",X"7C",X"57",X"C6",X"86",X"20",X"B7",X"57",X"CE",X"BD",X"B5",X"CF",X"BD",X"90",X"35",
		X"CC",X"00",X"29",X"BD",X"8F",X"0C",X"8E",X"FD",X"43",X"B6",X"57",X"C9",X"48",X"6E",X"96",X"7A",
		X"57",X"CE",X"26",X"03",X"7C",X"57",X"C6",X"39",X"B6",X"57",X"30",X"84",X"08",X"27",X"11",X"7F",
		X"57",X"C6",X"7C",X"57",X"C9",X"B6",X"57",X"C9",X"81",X"06",X"25",X"03",X"7F",X"57",X"C9",X"39",
		X"8E",X"FD",X"4F",X"B6",X"57",X"C9",X"48",X"6E",X"96",X"CC",X"00",X"02",X"B7",X"3A",X"00",X"B7",
		X"38",X"00",X"D7",X"8C",X"7E",X"81",X"42",X"39",X"CC",X"00",X"2A",X"BD",X"8F",X"0C",X"5C",X"BD",
		X"8F",X"0C",X"5C",X"BD",X"8F",X"0C",X"CE",X"FD",X"5B",X"E6",X"C0",X"8E",X"40",X"A4",X"86",X"02",
		X"97",X"F9",X"86",X"04",X"97",X"F8",X"86",X"05",X"97",X"F7",X"86",X"05",X"97",X"F6",X"86",X"0A",
		X"E7",X"89",X"08",X"00",X"A7",X"80",X"0A",X"F6",X"26",X"F6",X"30",X"88",X"1B",X"0A",X"F7",X"26",
		X"E9",X"30",X"88",X"20",X"E6",X"C0",X"0A",X"F8",X"26",X"DC",X"8E",X"40",X"AA",X"0A",X"F9",X"26",
		X"D1",X"8E",X"51",X"78",X"CC",X"02",X"04",X"DD",X"F6",X"CC",X"98",X"D0",X"A7",X"84",X"A7",X"04",
		X"8B",X"10",X"A7",X"08",X"A7",X"0C",X"E7",X"03",X"E7",X"0B",X"C0",X"10",X"E7",X"07",X"E7",X"0F",
		X"30",X"88",X"10",X"83",X"10",X"20",X"0A",X"F7",X"26",X"E2",X"86",X"04",X"97",X"F7",X"CC",X"C8",
		X"D0",X"0A",X"F6",X"26",X"D7",X"86",X"08",X"97",X"F6",X"8E",X"51",X"78",X"86",X"FD",X"33",X"5F",
		X"E6",X"C0",X"ED",X"01",X"ED",X"05",X"ED",X"09",X"ED",X"0D",X"30",X"88",X"10",X"0A",X"F6",X"26",
		X"EF",X"39",X"CC",X"00",X"2D",X"BD",X"8F",X"0C",X"5C",X"C1",X"38",X"23",X"F8",X"39",X"8E",X"40",
		X"85",X"B6",X"57",X"32",X"8D",X"12",X"8E",X"42",X"45",X"B6",X"57",X"31",X"8D",X"0A",X"8E",X"41",
		X"72",X"B6",X"57",X"30",X"C6",X"05",X"20",X"02",X"C6",X"06",X"D7",X"F6",X"44",X"1F",X"A9",X"C4",
		X"01",X"CB",X"30",X"E7",X"81",X"0A",X"F6",X"26",X"F3",X"39",X"0F",X"83",X"0F",X"84",X"86",X"01",
		X"97",X"82",X"CC",X"00",X"39",X"7E",X"8F",X"0C",X"8E",X"44",X"83",X"CE",X"30",X"02",X"0D",X"82",
		X"26",X"04",X"30",X"01",X"33",X"5F",X"6A",X"84",X"A6",X"84",X"84",X"1F",X"27",X"09",X"81",X"04",
		X"26",X"04",X"86",X"01",X"A7",X"C4",X"39",X"A7",X"C4",X"6D",X"84",X"26",X"F9",X"0A",X"82",X"10",
		X"2B",X"FE",X"CC",X"86",X"32",X"B7",X"41",X"69",X"39",X"CC",X"00",X"3C",X"BD",X"8F",X"0C",X"5C",
		X"C1",X"45",X"23",X"F8",X"CC",X"00",X"4E",X"BD",X"8F",X"0C",X"5C",X"C1",X"51",X"23",X"F8",X"39",
		X"B6",X"28",X"60",X"85",X"0F",X"27",X"53",X"81",X"10",X"25",X"54",X"CC",X"01",X"3B",X"BD",X"8F",
		X"0C",X"CC",X"00",X"3D",X"BD",X"8F",X"0C",X"5C",X"BD",X"8F",X"0C",X"C6",X"4E",X"BD",X"8F",X"0C",
		X"5C",X"BD",X"8F",X"0C",X"5C",X"BD",X"8F",X"0C",X"5C",X"BD",X"8F",X"0C",X"CE",X"BC",X"0C",X"8E",
		X"42",X"66",X"B6",X"28",X"60",X"43",X"84",X"0F",X"48",X"EC",X"C6",X"C3",X"30",X"30",X"E7",X"89",
		X"FE",X"E0",X"A7",X"81",X"B6",X"28",X"60",X"43",X"84",X"F0",X"44",X"44",X"44",X"EC",X"C6",X"C3",
		X"30",X"30",X"A7",X"84",X"E7",X"89",X"FE",X"E0",X"20",X"37",X"CC",X"00",X"3A",X"20",X"03",X"CC",
		X"00",X"3B",X"BD",X"8F",X"0C",X"CC",X"01",X"3D",X"BD",X"8F",X"0C",X"5C",X"BD",X"8F",X"0C",X"C6",
		X"4E",X"BD",X"8F",X"0C",X"5C",X"BD",X"8F",X"0C",X"5C",X"BD",X"8F",X"0C",X"5C",X"BD",X"8F",X"0C",
		X"86",X"20",X"8E",X"42",X"66",X"A7",X"84",X"A7",X"02",X"A7",X"89",X"FE",X"E0",X"A7",X"89",X"FE",
		X"E2",X"8E",X"41",X"CE",X"B6",X"30",X"00",X"43",X"84",X"18",X"44",X"44",X"44",X"8B",X"31",X"A7",
		X"84",X"8B",X"04",X"A7",X"02",X"B6",X"30",X"00",X"48",X"CC",X"4E",X"20",X"24",X"03",X"CC",X"46",
		X"46",X"A7",X"88",X"E6",X"E7",X"88",X"C6",X"B6",X"30",X"00",X"43",X"84",X"03",X"26",X"03",X"86",
		X"02",X"44",X"49",X"8B",X"30",X"A7",X"08",X"B6",X"30",X"00",X"C6",X"45",X"84",X"04",X"27",X"02",
		X"5A",X"4F",X"7E",X"8F",X"0C",X"8E",X"BD",X"5E",X"C6",X"06",X"A6",X"80",X"AB",X"80",X"5A",X"26",
		X"FB",X"81",X"1B",X"27",X"08",X"CC",X"00",X"52",X"BD",X"8F",X"0C",X"D7",X"00",X"86",X"1B",X"97",
		X"E7",X"CC",X"00",X"01",X"DD",X"D8",X"CC",X"00",X"46",X"BD",X"8F",X"0C",X"5C",X"7E",X"8F",X"0C",
		X"DC",X"D8",X"83",X"00",X"01",X"DD",X"D8",X"27",X"0E",X"10",X"83",X"01",X"E0",X"24",X"07",X"B6",
		X"57",X"30",X"84",X"10",X"26",X"01",X"39",X"CC",X"02",X"00",X"DD",X"D8",X"96",X"E7",X"4C",X"81",
		X"1B",X"23",X"01",X"4F",X"97",X"E7",X"84",X"0F",X"81",X"0A",X"25",X"02",X"8B",X"07",X"8B",X"30",
		X"B7",X"41",X"69",X"96",X"E7",X"44",X"44",X"44",X"44",X"81",X"0A",X"25",X"02",X"8B",X"07",X"8B",
		X"30",X"B7",X"41",X"89",X"BD",X"91",X"EF",X"96",X"E7",X"48",X"8E",X"FD",X"05",X"6E",X"96",X"4F",
		X"B7",X"57",X"C8",X"B7",X"30",X"05",X"B7",X"30",X"04",X"97",X"02",X"B7",X"3E",X"00",X"97",X"00",
		X"B7",X"3C",X"00",X"86",X"0E",X"B7",X"45",X"06",X"B7",X"28",X"00",X"8E",X"40",X"00",X"CC",X"20",
		X"0F",X"B7",X"20",X"00",X"E7",X"89",X"08",X"00",X"A7",X"80",X"8C",X"44",X"00",X"25",X"F2",X"30",
		X"88",X"40",X"A7",X"84",X"E7",X"89",X"08",X"00",X"A7",X"01",X"E7",X"89",X"08",X"01",X"A7",X"88",
		X"1E",X"E7",X"89",X"08",X"1E",X"A7",X"88",X"1F",X"E7",X"89",X"08",X"1F",X"30",X"88",X"20",X"8C",
		X"47",X"C0",X"25",X"DE",X"39",X"10",X"CE",X"57",X"FF",X"8D",X"A4",X"C6",X"4D",X"BD",X"83",X"C8",
		X"C6",X"48",X"BD",X"83",X"C8",X"BD",X"B7",X"79",X"20",X"FE",X"10",X"CE",X"57",X"FF",X"8D",X"8F",
		X"C6",X"4D",X"BD",X"83",X"C8",X"C6",X"4B",X"BD",X"83",X"C8",X"BD",X"B7",X"79",X"20",X"FE",X"10",
		X"CE",X"57",X"FF",X"BD",X"B5",X"CF",X"C6",X"4D",X"BD",X"83",X"C8",X"C6",X"49",X"BD",X"83",X"C8",
		X"C6",X"4C",X"BD",X"83",X"C8",X"BD",X"B7",X"79",X"20",X"FE",X"7F",X"30",X"00",X"B6",X"7F",X"FF",
		X"81",X"55",X"26",X"03",X"7E",X"60",X"00",X"B7",X"20",X"00",X"4F",X"B7",X"3A",X"00",X"B7",X"38",
		X"00",X"B7",X"57",X"FF",X"8E",X"40",X"00",X"B7",X"20",X"00",X"A7",X"84",X"A1",X"80",X"26",X"95",
		X"8C",X"57",X"FF",X"25",X"F2",X"8B",X"55",X"81",X"54",X"26",X"E9",X"4C",X"81",X"FF",X"26",X"01",
		X"4F",X"B7",X"20",X"00",X"A7",X"82",X"A1",X"84",X"10",X"26",X"FF",X"79",X"8C",X"40",X"00",X"22",
		X"EA",X"4F",X"A7",X"80",X"8C",X"57",X"FF",X"25",X"F8",X"86",X"10",X"BA",X"57",X"FF",X"B7",X"57",
		X"FF",X"10",X"8E",X"00",X"00",X"B7",X"20",X"00",X"3D",X"31",X"3F",X"26",X"F8",X"B6",X"57",X"FF",
		X"85",X"10",X"10",X"26",X"FF",X"79",X"48",X"10",X"25",X"FF",X"5F",X"44",X"44",X"10",X"25",X"FF",
		X"6E",X"B7",X"20",X"00",X"10",X"CE",X"57",X"FF",X"BD",X"B5",X"CF",X"B7",X"20",X"00",X"C6",X"4D",
		X"BD",X"83",X"C8",X"C6",X"49",X"BD",X"83",X"C8",X"C6",X"4A",X"BD",X"83",X"C8",X"B7",X"20",X"00",
		X"10",X"8E",X"00",X"00",X"CE",X"FD",X"73",X"8E",X"20",X"00",X"4F",X"5F",X"B7",X"20",X"00",X"EB",
		X"A2",X"89",X"00",X"30",X"1F",X"26",X"F5",X"10",X"A3",X"C3",X"34",X"01",X"11",X"83",X"FD",X"6B",
		X"26",X"E5",X"C6",X"22",X"E7",X"7D",X"BD",X"83",X"C8",X"6C",X"7D",X"E6",X"7D",X"C1",X"27",X"25",
		X"F5",X"8E",X"42",X"6B",X"6F",X"7F",X"35",X"01",X"27",X"2F",X"C6",X"07",X"86",X"42",X"A7",X"84",
		X"E7",X"89",X"08",X"00",X"86",X"41",X"A7",X"88",X"E0",X"E7",X"89",X"07",X"E0",X"86",X"44",X"A7",
		X"88",X"C0",X"E7",X"89",X"07",X"C0",X"E7",X"89",X"08",X"C0",X"E7",X"89",X"08",X"A0",X"E7",X"89",
		X"08",X"80",X"E7",X"89",X"08",X"60",X"B7",X"57",X"FA",X"30",X"02",X"8C",X"42",X"73",X"26",X"C6",
		X"8D",X"07",X"6D",X"7B",X"26",X"FE",X"7E",X"80",X"00",X"86",X"02",X"8E",X"00",X"00",X"B7",X"20",
		X"00",X"30",X"1F",X"26",X"F9",X"4A",X"26",X"F6",X"39",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E0",X"00",X"C0",X"04",X"A0",X"06",X"80",X"0C",X"02",X"03",X"05",X"07",X"01",X"01",X"01",X"02",
		X"01",X"03",X"01",X"04",X"01",X"05",X"01",X"06",X"01",X"07",X"02",X"01",X"02",X"03",X"02",X"05",
		X"03",X"01",X"03",X"02",X"03",X"04",X"04",X"01",X"04",X"03",X"00",X"00",X"00",X"02",X"00",X"47",
		X"53",X"58",X"00",X"01",X"75",X"58",X"4A",X"53",X"00",X"01",X"50",X"43",X"42",X"52",X"00",X"01",
		X"25",X"52",X"47",X"42",X"00",X"01",X"00",X"43",X"52",X"54",X"B2",X"F9",X"8C",X"F3",X"8E",X"3B",
		X"85",X"25",X"69",X"B7",X"83",X"C8",X"83",X"E5",X"00",X"00",X"84",X"05",X"84",X"12",X"84",X"38",
		X"84",X"45",X"84",X"9F",X"94",X"23",X"84",X"B3",X"8F",X"ED",X"84",X"C0",X"84",X"E7",X"BD",X"1A",
		X"BD",X"22",X"BD",X"2A",X"BD",X"36",X"BD",X"40",X"BD",X"4D",X"BD",X"5B",X"BD",X"6B",X"BD",X"82",
		X"BD",X"89",X"BD",X"90",X"BD",X"97",X"BD",X"9E",X"BD",X"A5",X"BD",X"BA",X"BD",X"CD",X"BD",X"E3",
		X"BD",X"FA",X"BE",X"11",X"BE",X"28",X"BE",X"3F",X"BE",X"56",X"BE",X"6D",X"BE",X"84",X"BE",X"9B",
		X"BE",X"A8",X"BE",X"B1",X"BE",X"BA",X"BE",X"C5",X"BE",X"CD",X"BE",X"D9",X"BE",X"E5",X"BE",X"EF",
		X"BF",X"00",X"BF",X"11",X"BF",X"1E",X"BF",X"2B",X"BF",X"38",X"BF",X"45",X"BF",X"52",X"BF",X"6A",
		X"BF",X"82",X"BF",X"92",X"BF",X"A2",X"BF",X"B1",X"BF",X"C0",X"BF",X"CB",X"BF",X"E8",X"C0",X"05",
		X"C0",X"22",X"C0",X"3F",X"C0",X"5C",X"C0",X"79",X"C0",X"88",X"C0",X"97",X"C0",X"A6",X"C0",X"B5",
		X"C0",X"C4",X"C0",X"D6",X"C0",X"E4",X"C0",X"F2",X"C1",X"04",X"C1",X"0D",X"C1",X"16",X"C1",X"26",
		X"C1",X"3E",X"C1",X"56",X"C1",X"68",X"C1",X"72",X"C1",X"7E",X"C1",X"8A",X"C1",X"9A",X"C1",X"A8",
		X"C1",X"B5",X"C1",X"C2",X"C1",X"CF",X"C1",X"DC",X"C1",X"E9",X"C1",X"FC",X"C2",X"04",X"C2",X"0C",
		X"C2",X"14",X"C2",X"1C",X"C2",X"3C",X"C2",X"5C",X"C2",X"6B",X"47",X"40",X"0F",X"10",X"12",X"1D",
		X"19",X"40",X"45",X"00",X"0F",X"11",X"12",X"1D",X"19",X"40",X"46",X"60",X"0F",X"16",X"17",X"12",
		X"1B",X"13",X"18",X"1A",X"15",X"40",X"45",X"5F",X"0F",X"13",X"1A",X"15",X"14",X"17",X"1C",X"40",
		X"45",X"5F",X"0F",X"46",X"52",X"45",X"45",X"20",X"50",X"4C",X"41",X"59",X"40",X"45",X"7F",X"0F",
		X"49",X"4E",X"56",X"41",X"4C",X"49",X"44",X"49",X"54",X"59",X"40",X"42",X"BC",X"0E",X"5C",X"4B",
		X"4F",X"4E",X"41",X"4D",X"49",X"20",X"31",X"39",X"38",X"34",X"40",X"43",X"0E",X"0E",X"1B",X"13",
		X"18",X"1A",X"15",X"20",X"1A",X"23",X"29",X"26",X"17",X"29",X"25",X"20",X"1C",X"23",X"24",X"27",
		X"15",X"40",X"42",X"F0",X"0A",X"31",X"53",X"54",X"40",X"42",X"F2",X"0B",X"32",X"4E",X"44",X"40",
		X"42",X"F4",X"0C",X"33",X"52",X"44",X"40",X"42",X"F6",X"0D",X"34",X"54",X"48",X"40",X"42",X"F8",
		X"0E",X"35",X"54",X"48",X"40",X"43",X"10",X"0E",X"50",X"55",X"53",X"48",X"20",X"53",X"54",X"41",
		X"52",X"54",X"20",X"42",X"55",X"54",X"54",X"4F",X"4E",X"40",X"42",X"F2",X"0E",X"4F",X"4E",X"45",
		X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"4F",X"4E",X"4C",X"59",X"40",X"43",X"12",X"0E",
		X"4F",X"4E",X"45",X"20",X"4F",X"52",X"20",X"54",X"57",X"4F",X"20",X"50",X"4C",X"41",X"59",X"45",
		X"52",X"53",X"40",X"43",X"35",X"0E",X"31",X"53",X"54",X"20",X"42",X"4F",X"4E",X"55",X"53",X"20",
		X"31",X"30",X"30",X"30",X"30",X"20",X"50",X"54",X"53",X"40",X"43",X"37",X"0E",X"41",X"4E",X"44",
		X"20",X"45",X"56",X"45",X"52",X"59",X"20",X"35",X"30",X"30",X"30",X"30",X"20",X"50",X"54",X"53",
		X"40",X"43",X"35",X"0E",X"31",X"53",X"54",X"20",X"42",X"4F",X"4E",X"55",X"53",X"20",X"32",X"30",
		X"30",X"30",X"30",X"20",X"50",X"54",X"53",X"40",X"43",X"37",X"0E",X"41",X"4E",X"44",X"20",X"45",
		X"56",X"45",X"52",X"59",X"20",X"36",X"30",X"30",X"30",X"30",X"20",X"50",X"54",X"53",X"40",X"43",
		X"35",X"0E",X"31",X"53",X"54",X"20",X"42",X"4F",X"4E",X"55",X"53",X"20",X"33",X"30",X"30",X"30",
		X"30",X"20",X"50",X"54",X"53",X"40",X"43",X"37",X"0E",X"41",X"4E",X"44",X"20",X"45",X"56",X"45",
		X"52",X"59",X"20",X"37",X"30",X"30",X"30",X"30",X"20",X"50",X"54",X"53",X"40",X"43",X"35",X"0E",
		X"31",X"53",X"54",X"20",X"42",X"4F",X"4E",X"55",X"53",X"20",X"34",X"30",X"30",X"30",X"30",X"20",
		X"50",X"54",X"53",X"40",X"43",X"37",X"0E",X"41",X"4E",X"44",X"20",X"45",X"56",X"45",X"52",X"59",
		X"20",X"38",X"30",X"30",X"30",X"30",X"20",X"50",X"54",X"53",X"40",X"42",X"91",X"0E",X"47",X"41",
		X"4D",X"45",X"20",X"4F",X"56",X"45",X"52",X"40",X"47",X"BF",X"0F",X"1B",X"1C",X"23",X"25",X"15",
		X"40",X"41",X"68",X"3D",X"E8",X"E9",X"4E",X"EB",X"EC",X"40",X"41",X"69",X"3D",X"F8",X"F9",X"FA",
		X"FB",X"FC",X"FD",X"FE",X"40",X"41",X"6A",X"3D",X"D8",X"D9",X"DA",X"DB",X"40",X"41",X"6B",X"3D",
		X"D0",X"D1",X"D2",X"D3",X"D4",X"D5",X"D6",X"D7",X"40",X"41",X"6C",X"3D",X"E0",X"E1",X"E2",X"E3",
		X"E4",X"E5",X"E6",X"E7",X"40",X"41",X"6D",X"3D",X"F0",X"F1",X"F2",X"F3",X"F4",X"F5",X"40",X"42",
		X"BA",X"0B",X"60",X"61",X"62",X"63",X"64",X"65",X"66",X"67",X"68",X"69",X"6A",X"6B",X"6C",X"40",
		X"42",X"BB",X"0B",X"70",X"71",X"72",X"73",X"74",X"75",X"76",X"77",X"78",X"79",X"7A",X"7B",X"7C",
		X"40",X"43",X"28",X"0F",X"52",X"41",X"4D",X"20",X"20",X"20",X"20",X"4F",X"4B",X"40",X"43",X"2B",
		X"0F",X"52",X"4F",X"4D",X"31",X"20",X"20",X"20",X"4F",X"4B",X"40",X"43",X"2D",X"0F",X"52",X"4F",
		X"4D",X"32",X"20",X"20",X"20",X"4F",X"4B",X"40",X"43",X"2F",X"0F",X"52",X"4F",X"4D",X"33",X"20",
		X"20",X"20",X"4F",X"4B",X"40",X"43",X"31",X"0F",X"52",X"4F",X"4D",X"34",X"20",X"20",X"20",X"4F",
		X"4B",X"40",X"43",X"34",X"1A",X"31",X"45",X"B9",X"B9",X"B2",X"B9",X"B9",X"B9",X"B9",X"B9",X"C2",
		X"B9",X"B9",X"B9",X"E5",X"B9",X"F6",X"B9",X"B9",X"B9",X"40",X"43",X"35",X"1A",X"52",X"76",X"48",
		X"77",X"58",X"59",X"6F",X"7E",X"7F",X"C0",X"D0",X"E2",X"F3",X"F4",X"F5",X"D6",X"E6",X"CA",X"BB",
		X"CF",X"40",X"46",X"BE",X"0E",X"5C",X"4B",X"4F",X"4E",X"41",X"4D",X"49",X"20",X"31",X"39",X"38",
		X"34",X"40",X"42",X"C2",X"0F",X"43",X"4F",X"4C",X"4F",X"52",X"20",X"20",X"20",X"54",X"45",X"53",
		X"54",X"40",X"43",X"63",X"0F",X"56",X"52",X"41",X"4D",X"20",X"20",X"43",X"4F",X"4C",X"4F",X"52",
		X"40",X"43",X"71",X"0F",X"4F",X"42",X"4A",X"20",X"20",X"20",X"43",X"4F",X"4C",X"4F",X"52",X"40",
		X"42",X"62",X"0F",X"49",X"4F",X"20",X"54",X"45",X"53",X"54",X"40",X"43",X"85",X"0F",X"31",X"50",
		X"20",X"4C",X"45",X"46",X"54",X"20",X"20",X"20",X"30",X"20",X"20",X"20",X"32",X"50",X"20",X"4C",
		X"45",X"46",X"54",X"20",X"20",X"20",X"30",X"40",X"43",X"87",X"0F",X"31",X"50",X"20",X"52",X"49",
		X"47",X"48",X"54",X"20",X"20",X"30",X"20",X"20",X"20",X"32",X"50",X"20",X"52",X"49",X"47",X"48");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
