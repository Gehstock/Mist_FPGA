library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity gravitar_vec_rom1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of gravitar_vec_rom1 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"FF",X"80",X"00",X"C0",X"00",X"00",X"40",X"80",X"60",X"00",X"60",X"80",X"40",X"1F",
		X"60",X"80",X"60",X"1F",X"A0",X"9F",X"00",X"00",X"60",X"80",X"00",X"C0",X"40",X"01",X"C0",X"80",
		X"C0",X"00",X"40",X"9F",X"40",X"00",X"60",X"80",X"00",X"00",X"40",X"80",X"A0",X"1F",X"60",X"80",
		X"00",X"C0",X"80",X"1F",X"80",X"80",X"40",X"1F",X"80",X"9F",X"00",X"00",X"FF",X"80",X"00",X"C0",
		X"C0",X"00",X"60",X"80",X"E0",X"00",X"A0",X"9F",X"00",X"00",X"40",X"80",X"A0",X"1F",X"C0",X"80",
		X"60",X"1E",X"40",X"9F",X"80",X"1F",X"C0",X"80",X"00",X"C0",X"40",X"01",X"A0",X"80",X"E0",X"00",
		X"60",X"9F",X"A0",X"1F",X"FF",X"80",X"00",X"C0",X"40",X"1F",X"FF",X"80",X"00",X"C0",X"C0",X"00",
		X"FF",X"80",X"00",X"C0",X"80",X"1F",X"FF",X"80",X"00",X"C0",X"E0",X"1E",X"FF",X"80",X"00",X"C0",
		X"00",X"00",X"FF",X"80",X"E0",X"00",X"00",X"00",X"40",X"00",X"40",X"9F",X"80",X"00",X"40",X"80",
		X"A0",X"00",X"80",X"9F",X"00",X"00",X"FF",X"80",X"00",X"C0",X"00",X"00",X"FF",X"80",X"E0",X"00",
		X"01",X"1F",X"60",X"01",X"FF",X"80",X"00",X"00",X"01",X"9F",X"00",X"C0",X"00",X"00",X"A0",X"80",
		X"20",X"01",X"60",X"9F",X"00",X"00",X"80",X"80",X"FF",X"00",X"80",X"80",X"00",X"C0",X"01",X"1F",
		X"C0",X"80",X"00",X"00",X"40",X"80",X"00",X"C0",X"FF",X"00",X"80",X"00",X"FF",X"80",X"E0",X"01",
		X"00",X"00",X"60",X"1F",X"C0",X"9F",X"A0",X"00",X"C0",X"9F",X"00",X"00",X"80",X"9F",X"40",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"80",X"00",X"C0",X"00",X"00",X"80",X"80",X"80",X"00",X"40",X"80",
		X"40",X"1F",X"40",X"80",X"20",X"02",X"00",X"00",X"A0",X"1F",X"C0",X"9F",X"60",X"00",X"C0",X"9F",
		X"00",X"00",X"80",X"9F",X"40",X"00",X"00",X"00",X"00",X"00",X"FF",X"80",X"00",X"C0",X"20",X"00",
		X"20",X"80",X"00",X"00",X"60",X"80",X"60",X"00",X"40",X"80",X"A0",X"1F",X"40",X"80",X"00",X"02",
		X"00",X"00",X"00",X"00",X"01",X"9F",X"40",X"00",X"00",X"00",X"00",X"00",X"FF",X"80",X"00",X"C0",
		X"C0",X"1F",X"40",X"80",X"00",X"00",X"80",X"80",X"40",X"00",X"40",X"80",X"00",X"02",X"00",X"00",
		X"00",X"00",X"01",X"9F",X"40",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",X"C0",X"1F",X"40",X"80",
		X"00",X"C0",X"C0",X"00",X"40",X"80",X"40",X"1F",X"40",X"80",X"A0",X"1F",X"80",X"80",X"00",X"C0",
		X"80",X"00",X"20",X"80",X"00",X"00",X"40",X"80",X"80",X"1F",X"A0",X"80",X"60",X"02",X"00",X"00",
		X"00",X"00",X"80",X"9F",X"60",X"1F",X"C0",X"9F",X"A0",X"00",X"C0",X"9F",X"40",X"00",X"40",X"80",
		X"00",X"00",X"C0",X"80",X"00",X"C0",X"80",X"00",X"20",X"80",X"00",X"00",X"40",X"80",X"80",X"1F",
		X"20",X"80",X"80",X"00",X"80",X"80",X"E0",X"01",X"00",X"00",X"00",X"00",X"80",X"9F",X"80",X"1F",
		X"C0",X"9F",X"80",X"00",X"C0",X"9F",X"40",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",X"C0",X"1F",
		X"40",X"80",X"00",X"C0",X"A0",X"1F",X"40",X"80",X"00",X"00",X"60",X"80",X"A0",X"00",X"60",X"80",
		X"00",X"C0",X"00",X"00",X"80",X"80",X"60",X"00",X"40",X"80",X"A0",X"1F",X"40",X"80",X"A0",X"01",
		X"00",X"00",X"60",X"1F",X"C0",X"9F",X"A0",X"00",X"C0",X"9F",X"00",X"00",X"80",X"9F",X"40",X"00",
		X"40",X"80",X"00",X"00",X"C0",X"80",X"00",X"C0",X"60",X"00",X"40",X"80",X"A0",X"1F",X"40",X"80",
		X"00",X"00",X"60",X"80",X"80",X"1F",X"20",X"80",X"20",X"02",X"00",X"00",X"A0",X"1F",X"C0",X"9F",
		X"60",X"00",X"C0",X"9F",X"00",X"00",X"80",X"9F",X"40",X"00",X"00",X"00",X"00",X"00",X"FF",X"80",
		X"00",X"C0",X"00",X"00",X"40",X"80",X"40",X"00",X"40",X"80",X"80",X"00",X"40",X"80",X"80",X"1F",
		X"40",X"80",X"E0",X"01",X"00",X"00",X"00",X"00",X"01",X"9F",X"40",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"80",X"00",X"C0",X"A0",X"1F",X"40",X"80",X"00",X"00",X"40",X"80",X"80",X"00",X"40",X"80",
		X"80",X"1F",X"40",X"80",X"40",X"02",X"00",X"00",X"00",X"00",X"01",X"9F",X"40",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"80",X"00",X"C0",X"20",X"00",X"40",X"80",X"00",X"00",X"40",X"80",X"C0",X"00",
		X"40",X"80",X"40",X"1F",X"40",X"80",X"20",X"02",X"00",X"00",X"00",X"00",X"01",X"9F",X"40",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"80",X"00",X"C0",X"40",X"00",X"40",X"80",X"00",X"00",X"40",X"80",
		X"C0",X"1F",X"80",X"80",X"20",X"02",X"00",X"00",X"80",X"1F",X"C0",X"9F",X"80",X"00",X"C0",X"9F",
		X"00",X"00",X"80",X"9F",X"40",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",X"C0",X"1F",X"40",X"80",
		X"00",X"C0",X"40",X"00",X"60",X"80",X"00",X"00",X"A0",X"80",X"00",X"C0",X"A0",X"00",X"40",X"80",
		X"60",X"1F",X"40",X"80",X"00",X"00",X"40",X"80",X"80",X"1F",X"40",X"80",X"60",X"02",X"00",X"00",
		X"00",X"00",X"01",X"9F",X"40",X"00",X"40",X"80",X"00",X"00",X"C0",X"80",X"00",X"C0",X"00",X"00",
		X"C0",X"80",X"40",X"00",X"40",X"80",X"A0",X"1E",X"00",X"00",X"00",X"00",X"60",X"9F",X"A0",X"00",
		X"A0",X"80",X"00",X"00",X"80",X"9F",X"80",X"00",X"80",X"9F",X"00",X"C0",X"A0",X"1F",X"60",X"80",
		X"40",X"00",X"60",X"80",X"C0",X"1F",X"40",X"80",X"40",X"1F",X"00",X"00",X"C0",X"1F",X"C0",X"9F",
		X"00",X"00",X"40",X"80",X"80",X"03",X"00",X"00",X"00",X"00",X"C0",X"9F",X"40",X"1F",X"40",X"9F",
		X"00",X"C0",X"A0",X"1F",X"60",X"80",X"A0",X"1F",X"A0",X"9F",X"C0",X"1F",X"00",X"00",X"00",X"00",
		X"60",X"80",X"A0",X"00",X"A0",X"80",X"80",X"00",X"80",X"9F",X"80",X"00",X"80",X"80",X"20",X"03",
		X"00",X"00",X"A0",X"1F",X"A0",X"9F",X"A0",X"1F",X"60",X"80",X"00",X"00",X"80",X"9F",X"80",X"1F",
		X"80",X"9F",X"00",X"C0",X"00",X"00",X"A0",X"80",X"A0",X"1F",X"60",X"80",X"00",X"03",X"00",X"00",
		X"00",X"00",X"80",X"9F",X"80",X"00",X"80",X"9F",X"00",X"C0",X"00",X"00",X"FF",X"80",X"00",X"03",
		X"01",X"1F",X"00",X"00",X"60",X"80",X"80",X"00",X"80",X"80",X"80",X"00",X"80",X"9F",X"00",X"00",
		X"A0",X"9F",X"80",X"00",X"FF",X"80",X"00",X"C0",X"00",X"00",X"FF",X"80",X"01",X"1F",X"01",X"9F",
		X"60",X"1F",X"A0",X"80",X"60",X"00",X"60",X"80",X"00",X"00",X"A0",X"9F",X"60",X"00",X"60",X"80",
		X"E0",X"03",X"00",X"00",X"00",X"00",X"A0",X"9F",X"80",X"01",X"60",X"9F",X"00",X"C0",X"40",X"00",
		X"40",X"80",X"00",X"00",X"80",X"80",X"40",X"00",X"40",X"80",X"60",X"00",X"A0",X"9F",X"80",X"00",
		X"60",X"80",X"40",X"00",X"C0",X"9F",X"40",X"00",X"40",X"80",X"20",X"01",X"00",X"00",X"40",X"00",
		X"C0",X"9F",X"40",X"00",X"40",X"80",X"00",X"00",X"60",X"9F",X"60",X"00",X"A0",X"9F",X"00",X"C0",
		X"00",X"00",X"C0",X"80",X"40",X"00",X"40",X"80",X"80",X"00",X"80",X"9F",X"00",X"00",X"E0",X"9F",
		X"60",X"00",X"A0",X"9F",X"00",X"C0",X"00",X"00",X"FF",X"80",X"40",X"1F",X"40",X"9F",X"40",X"1F",
		X"C0",X"80",X"00",X"C0",X"20",X"1F",X"FF",X"80",X"80",X"01",X"00",X"00",X"E0",X"00",X"A0",X"9F",
		X"00",X"00",X"60",X"80",X"00",X"C0",X"00",X"00",X"FF",X"80",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"A0",X"9F",X"A0",X"00",X"60",X"9F",X"E0",X"00",X"00",X"00",X"00",X"00",X"FF",X"80",X"00",X"C0",
		X"00",X"00",X"A0",X"80",X"60",X"00",X"60",X"80",X"80",X"01",X"00",X"00",X"01",X"1F",X"01",X"9F",
		X"80",X"01",X"00",X"00",X"00",X"00",X"FF",X"80",X"00",X"C0",X"A0",X"00",X"60",X"80",X"00",X"00",
		X"60",X"80",X"40",X"00",X"40",X"80",X"A0",X"00",X"00",X"00",X"40",X"00",X"A0",X"9F",X"00",X"00",
		X"C0",X"9F",X"C0",X"1F",X"A0",X"9F",X"80",X"00",X"00",X"00",X"00",X"00",X"FF",X"80",X"00",X"C0",
		X"00",X"00",X"80",X"80",X"A0",X"00",X"80",X"9F",X"80",X"00",X"00",X"00",X"00",X"00",X"FF",X"80",
		X"01",X"1F",X"00",X"00",X"20",X"1F",X"60",X"9F",X"A0",X"1F",X"60",X"80",X"00",X"00",X"40",X"80",
		X"00",X"C0",X"40",X"00",X"60",X"80",X"00",X"00",X"A0",X"80",X"FF",X"00",X"00",X"00",X"80",X"1F",
		X"C0",X"9F",X"80",X"00",X"A0",X"9F",X"00",X"00",X"A0",X"9F",X"FF",X"00",X"00",X"00",X"C0",X"1F",
		X"40",X"80",X"C0",X"1F",X"C0",X"9F",X"80",X"1F",X"FF",X"80",X"00",X"C0",X"80",X"00",X"A0",X"80",
		X"A0",X"00",X"60",X"80",X"E0",X"00",X"01",X"9F",X"00",X"00",X"FF",X"80",X"00",X"C0",X"80",X"1E",
		X"FF",X"80",X"FF",X"00",X"00",X"00",X"80",X"00",X"A0",X"9F",X"00",X"00",X"60",X"80",X"00",X"C0",
		X"C0",X"1F",X"FF",X"80",X"C0",X"00",X"00",X"00",X"00",X"00",X"C0",X"9F",X"80",X"00",X"40",X"9F",
		X"80",X"00",X"00",X"00",X"00",X"00",X"FF",X"80",X"00",X"C0",X"80",X"1F",X"80",X"80",X"00",X"00",
		X"80",X"80",X"80",X"01",X"00",X"00",X"00",X"00",X"20",X"9F",X"C0",X"1F",X"E0",X"9F",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"80",X"00",X"C0",X"80",X"00",X"60",X"80",X"00",X"00",X"A0",X"80",
		X"40",X"01",X"00",X"00",X"00",X"00",X"20",X"9F",X"C0",X"1F",X"E0",X"9F",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"80",X"00",X"C0",X"80",X"00",X"60",X"80",X"00",X"00",X"A0",X"80",X"C0",X"00",
		X"40",X"9F",X"00",X"00",X"C0",X"9F",X"80",X"00",X"00",X"00",X"00",X"00",X"FF",X"80",X"00",X"C0",
		X"80",X"1F",X"40",X"80",X"A0",X"1F",X"40",X"80",X"40",X"1F",X"80",X"80",X"00",X"C0",X"00",X"00",
		X"80",X"80",X"40",X"00",X"40",X"80",X"00",X"00",X"40",X"80",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"01",X"9F",X"80",X"00",X"80",X"80",X"00",X"00",X"80",X"80",X"00",X"C0",X"00",X"00",X"C0",X"80",
		X"E0",X"00",X"40",X"9F",X"80",X"00",X"00",X"00",X"00",X"00",X"FF",X"80",X"00",X"C0",X"01",X"1F",
		X"FF",X"C0",X"00",X"02",X"00",X"00",X"01",X"1F",X"01",X"DF",X"00",X"C0",X"01",X"1F",X"FF",X"C0",
		X"80",X"01",X"00",X"00",X"80",X"00",X"80",X"DF",X"80",X"00",X"80",X"C0",X"80",X"01",X"00",X"00",
		X"01",X"1F",X"01",X"DF",X"00",X"03",X"FF",X"00",X"80",X"00",X"80",X"DF",X"00",X"C0",X"01",X"1F",
		X"FF",X"C0",X"80",X"01",X"00",X"00",X"FF",X"00",X"01",X"DF",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"FF",X"C0",X"80",X"01",X"00",X"00",X"01",X"1F",X"01",X"DF",X"00",X"02",X"00",X"00",X"01",X"1F",
		X"FF",X"C0",X"00",X"C0",X"00",X"00",X"FF",X"C0",X"FF",X"00",X"00",X"00",X"00",X"00",X"80",X"DF",
		X"80",X"00",X"80",X"DF",X"00",X"03",X"00",X"00",X"FF",X"00",X"FF",X"C0",X"00",X"C0",X"00",X"00",
		X"FF",X"C0",X"FF",X"00",X"00",X"00",X"00",X"00",X"01",X"DF",X"80",X"03",X"00",X"00",X"01",X"1F",
		X"FF",X"C0",X"00",X"02",X"00",X"00",X"01",X"1F",X"01",X"DF",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"FF",X"C0",X"00",X"C0",X"00",X"00",X"FF",X"C0",X"FF",X"00",X"00",X"00",X"00",X"00",X"01",X"DF",
		X"80",X"02",X"00",X"00",X"01",X"1F",X"FF",X"C0",X"80",X"01",X"00",X"00",X"80",X"00",X"80",X"DF",
		X"00",X"00",X"80",X"C0",X"FF",X"00",X"00",X"00",X"00",X"00",X"01",X"DF",X"FF",X"00",X"00",X"00",
		X"FF",X"00",X"FF",X"C0",X"00",X"C0",X"00",X"00",X"FF",X"C0",X"80",X"01",X"00",X"00",X"80",X"1F",
		X"80",X"DF",X"00",X"00",X"80",X"DF",X"80",X"01",X"00",X"00",X"00",X"00",X"FF",X"C0",X"80",X"01",
		X"00",X"00",X"00",X"00",X"01",X"DF",X"80",X"00",X"00",X"00",X"00",X"00",X"FF",X"C0",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"01",X"DF",X"00",X"C0",X"FF",X"00",X"FF",X"C0",X"80",X"00",X"01",X"1F",
		X"FF",X"00",X"FF",X"C0",X"80",X"00",X"00",X"00",X"80",X"1F",X"80",X"DF",X"00",X"00",X"80",X"DF",
		X"80",X"00",X"FF",X"00",X"FF",X"00",X"01",X"DF",X"80",X"00",X"00",X"00",X"01",X"1F",X"FF",X"C0",
		X"80",X"01",X"00",X"00",X"80",X"00",X"80",X"DF",X"00",X"00",X"80",X"DF",X"00",X"C0",X"FF",X"00",
		X"FF",X"C0",X"80",X"00",X"01",X"1F",X"80",X"00",X"80",X"C0",X"80",X"00",X"80",X"DF",X"80",X"01",
		X"00",X"00",X"01",X"1F",X"FF",X"C0",X"00",X"C0",X"FF",X"00",X"FF",X"C0",X"FF",X"00",X"01",X"DF",
		X"00",X"C0",X"01",X"1F",X"FF",X"80",X"00",X"C0",X"FF",X"00",X"FF",X"80",X"00",X"C0",X"00",X"00",
		X"FF",X"80",X"00",X"00",X"01",X"1F",X"FF",X"00",X"FF",X"80",X"FF",X"00",X"01",X"1F",X"FF",X"00",
		X"FF",X"80",X"00",X"C0",X"00",X"00",X"FF",X"80",X"FF",X"00",X"01",X"1F",X"FF",X"00",X"FF",X"80",
		X"FF",X"00",X"01",X"9F",X"00",X"C0",X"00",X"00",X"FF",X"80",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"01",X"9F",X"FF",X"00",X"FF",X"80",X"00",X"C0",X"00",X"00",X"FF",X"80",X"FF",X"00",X"01",X"9F",
		X"FF",X"01",X"00",X"00",X"01",X"1F",X"FF",X"80",X"00",X"C0",X"00",X"00",X"FF",X"80",X"FF",X"00",
		X"00",X"00",X"01",X"1F",X"01",X"9F",X"FF",X"01",X"00",X"00",X"00",X"00",X"FF",X"80",X"00",X"C0",
		X"FF",X"00",X"FF",X"80",X"00",X"00",X"01",X"1F",X"FF",X"00",X"FF",X"80",X"00",X"00",X"01",X"9F",
		X"00",X"C0",X"00",X"00",X"FF",X"80",X"FF",X"00",X"01",X"9F",X"00",X"00",X"FF",X"80",X"00",X"C0",
		X"00",X"00",X"FF",X"80",X"00",X"00",X"01",X"1F",X"FF",X"00",X"FF",X"80",X"00",X"00",X"01",X"9F",
		X"00",X"C0",X"01",X"1F",X"FF",X"80",X"FF",X"00",X"01",X"1F",X"FF",X"00",X"FF",X"80",X"00",X"00",
		X"01",X"9F",X"FF",X"00",X"FF",X"80",X"01",X"1F",X"01",X"1E",X"FF",X"00",X"FF",X"80",X"FF",X"01",
		X"FF",X"80",X"00",X"C0",X"01",X"1F",X"FF",X"80",X"FF",X"03",X"01",X"1F",X"FF",X"00",X"FF",X"80",
		X"00",X"00",X"01",X"9F",X"FF",X"00",X"FF",X"80",X"00",X"00",X"01",X"1F",X"FF",X"01",X"FF",X"80",
		X"00",X"C0",X"00",X"00",X"FF",X"80",X"FF",X"00",X"00",X"00",X"FF",X"00",X"01",X"9F",X"00",X"00",
		X"FF",X"80",X"00",X"03",X"00",X"00",X"FF",X"00",X"01",X"9F",X"FF",X"01",X"00",X"00",X"00",X"00",
		X"FF",X"80",X"00",X"C0",X"FF",X"00",X"FF",X"80",X"00",X"00",X"01",X"9F",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"80",X"00",X"03",X"01",X"1F",X"00",X"00",X"FF",X"80",X"FF",X"00",X"01",X"9F",
		X"FF",X"00",X"FF",X"80",X"FF",X"00",X"01",X"9F",X"00",X"C0",X"FF",X"00",X"FF",X"80",X"FF",X"01");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
