library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity travusa_chr_bit2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of travusa_chr_bit2 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"04",X"3C",X"00",X"24",X"18",X"3F",X"00",
		X"80",X"40",X"F3",X"0C",X"30",X"C0",X"38",X"04",X"3F",X"00",X"3F",X"06",X"0C",X"06",X"3F",X"00",
		X"80",X"40",X"F3",X"0C",X"30",X"C0",X"00",X"A0",X"3F",X"00",X"01",X"00",X"12",X"21",X"21",X"1E",
		X"00",X"01",X"FF",X"41",X"00",X"19",X"24",X"24",X"61",X"91",X"89",X"47",X"00",X"19",X"24",X"24",
		X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"6C",X"82",X"82",X"82",X"82",X"6C",X"00",X"00",
		X"6C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"92",X"92",X"92",X"92",X"60",X"00",X"00",
		X"6C",X"92",X"92",X"92",X"92",X"00",X"00",X"00",X"6C",X"10",X"10",X"10",X"10",X"0C",X"00",X"00",
		X"60",X"92",X"92",X"92",X"92",X"0C",X"00",X"00",X"60",X"92",X"92",X"92",X"92",X"6C",X"00",X"00",
		X"6C",X"02",X"02",X"02",X"02",X"00",X"00",X"00",X"6C",X"92",X"92",X"92",X"92",X"6C",X"00",X"00",
		X"6C",X"92",X"92",X"92",X"92",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"41",
		X"00",X"3F",X"7F",X"77",X"6F",X"7B",X"73",X"77",X"00",X"FC",X"FE",X"EE",X"F6",X"9E",X"0E",X"6E",
		X"76",X"70",X"79",X"6F",X"77",X"7F",X"3F",X"00",X"EE",X"CE",X"DE",X"F6",X"EE",X"FE",X"FC",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",
		X"FF",X"FF",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"C0",X"C0",X"C0",X"00",X"80",X"80",X"80",X"FC",
		X"FF",X"FF",X"FF",X"82",X"82",X"7F",X"7F",X"FF",X"FC",X"FC",X"FC",X"40",X"40",X"C0",X"80",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5F",X"5F",X"00",X"00",X"00",
		X"00",X"00",X"03",X"03",X"00",X"03",X"03",X"00",X"00",X"14",X"3E",X"14",X"28",X"7C",X"28",X"00",
		X"00",X"24",X"76",X"52",X"FF",X"4A",X"6E",X"24",X"00",X"42",X"A4",X"48",X"10",X"24",X"4A",X"84",
		X"00",X"50",X"20",X"56",X"49",X"59",X"76",X"20",X"00",X"00",X"00",X"03",X"07",X"00",X"00",X"00",
		X"1F",X"9F",X"91",X"81",X"81",X"81",X"FF",X"7E",X"46",X"CF",X"89",X"99",X"99",X"91",X"F3",X"62",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"30",X"70",X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"08",X"08",X"00",
		X"00",X"00",X"00",X"00",X"60",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"3E",X"41",X"41",X"41",X"7F",X"7F",X"3E",X"00",X"00",X"00",X"7F",X"7F",X"7F",X"01",X"00",
		X"00",X"46",X"4F",X"4F",X"49",X"79",X"79",X"71",X"00",X"36",X"7F",X"7F",X"49",X"49",X"41",X"22",
		X"00",X"20",X"7F",X"7F",X"7F",X"21",X"22",X"3C",X"00",X"31",X"79",X"79",X"49",X"4F",X"4F",X"4F",
		X"00",X"31",X"79",X"79",X"49",X"4F",X"4F",X"3E",X"00",X"03",X"0F",X"7F",X"7D",X"71",X"01",X"03",
		X"00",X"36",X"79",X"79",X"49",X"4F",X"4F",X"36",X"00",X"3E",X"79",X"79",X"49",X"4F",X"4F",X"46",
		X"00",X"00",X"00",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"12",X"32",X"00",X"00",X"00",
		X"7C",X"08",X"00",X"06",X"09",X"09",X"7F",X"00",X"00",X"14",X"14",X"14",X"14",X"14",X"14",X"14",
		X"40",X"00",X"24",X"54",X"54",X"48",X"00",X"48",X"00",X"02",X"07",X"0D",X"59",X"01",X"03",X"02",
		X"00",X"63",X"36",X"1C",X"08",X"1C",X"36",X"63",X"00",X"7E",X"7F",X"7F",X"11",X"11",X"11",X"7E",
		X"00",X"36",X"49",X"49",X"49",X"7F",X"7F",X"7F",X"00",X"22",X"41",X"41",X"41",X"7F",X"7F",X"3E",
		X"00",X"3E",X"7F",X"7F",X"41",X"41",X"41",X"7F",X"00",X"49",X"49",X"49",X"49",X"7F",X"7F",X"7F",
		X"00",X"09",X"09",X"09",X"09",X"7F",X"7F",X"7F",X"00",X"3A",X"7B",X"7B",X"49",X"49",X"41",X"3E",
		X"00",X"7F",X"08",X"08",X"08",X"7F",X"7F",X"7F",X"00",X"00",X"00",X"7F",X"7F",X"7F",X"00",X"00",
		X"00",X"00",X"00",X"3F",X"7F",X"7F",X"40",X"40",X"00",X"61",X"72",X"7C",X"18",X"0F",X"0F",X"7F",
		X"00",X"40",X"40",X"40",X"40",X"7F",X"7F",X"7F",X"00",X"7E",X"7F",X"01",X"7F",X"7F",X"01",X"7F",
		X"00",X"7E",X"7F",X"7F",X"01",X"01",X"01",X"7F",X"00",X"3E",X"41",X"41",X"41",X"7F",X"7F",X"3E",
		X"00",X"0E",X"11",X"11",X"11",X"7F",X"7F",X"7F",X"00",X"7E",X"71",X"41",X"41",X"7F",X"7F",X"3E",
		X"00",X"76",X"79",X"79",X"09",X"0F",X"0F",X"7F",X"00",X"32",X"79",X"79",X"49",X"4F",X"4F",X"26",
		X"00",X"01",X"01",X"7F",X"7F",X"7F",X"01",X"01",X"00",X"3F",X"40",X"40",X"40",X"7F",X"7F",X"3F",
		X"00",X"0F",X"10",X"20",X"60",X"7F",X"3F",X"1F",X"00",X"3F",X"40",X"7F",X"7F",X"40",X"7F",X"3F",
		X"00",X"61",X"72",X"7C",X"1C",X"3F",X"67",X"43",X"00",X"07",X"08",X"70",X"78",X"7F",X"0F",X"07",
		X"00",X"43",X"47",X"4F",X"5D",X"79",X"71",X"61",X"A2",X"A2",X"A2",X"A2",X"A2",X"9C",X"41",X"3E",
		X"00",X"7E",X"7E",X"7E",X"7E",X"7E",X"00",X"00",X"00",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"04",X"00",X"09",X"40",X"00",X"24",X"46",X"00",X"00",X"02",X"80",X"48",X"00",X"00",X"44",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",X"3F",X"3F",
		X"80",X"C0",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"C0",X"00",X"60",X"40",X"80",X"70",X"4C",X"64",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"E0",X"A8",X"01",X"82",X"00",X"20",X"04",
		X"9D",X"73",X"84",X"94",X"64",X"89",X"20",X"12",X"DD",X"A5",X"B0",X"C6",X"09",X"5A",X"22",X"85",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F5",X"A5",X"3A",X"9C",X"A5",X"5E",X"E0",X"04",
		X"B8",X"E4",X"28",X"7C",X"D6",X"8F",X"6A",X"79",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",
		X"01",X"C4",X"E0",X"F8",X"FE",X"FF",X"FF",X"FF",X"00",X"80",X"02",X"50",X"44",X"84",X"E0",X"F8",
		X"AE",X"49",X"BD",X"26",X"6A",X"B9",X"0E",X"6F",X"40",X"00",X"80",X"C0",X"70",X"C0",X"40",X"70",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C8",X"90",X"3C",X"E6",X"2C",X"79",X"C4",X"16",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"40",X"80",X"C0",X"00",X"50",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"FF",X"FF",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"FF",X"FF",X"FF",X"FF",X"F8",X"F8",X"F8",X"F8",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"1F",X"1F",X"1F",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"E7",X"C3",X"C3",X"E7",X"FF",X"FF",X"FF",X"FF",X"F9",X"F4",X"F0",X"F9",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"03",X"0F",X"1F",X"7C",X"F8",X"E0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E0",X"83",X"07",X"1F",X"7F",X"FF",X"FF",X"FF",
		X"03",X"0F",X"1F",X"7C",X"F8",X"E0",X"83",X"07",X"00",X"00",X"00",X"00",X"00",X"03",X"0F",X"1F",
		X"7C",X"F8",X"E0",X"83",X"07",X"1F",X"7F",X"FF",X"1F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"1F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"1F",X"7C",X"F8",X"E0",X"83",X"07",X"1F",X"7F",X"00",X"00",X"00",X"03",X"0F",X"1F",X"7C",X"F8",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"83",X"07",X"1F",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"30",X"60",X"98",X"D0",X"3F",X"7B",X"51",X"10",X"F8",X"E0",X"83",X"07",X"1F",X"7F",X"FF",X"FF",
		X"00",X"03",X"0F",X"1F",X"7C",X"F8",X"E0",X"83",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0F",
		X"0F",X"1F",X"7C",X"F8",X"E0",X"83",X"07",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E7",X"2A",X"9F",X"D5",X"D0",X"82",X"1C",X"02",
		X"01",X"03",X"02",X"00",X"03",X"0F",X"1F",X"7C",X"3F",X"1C",X"86",X"C7",X"E7",X"F3",X"F8",X"FC",
		X"FF",X"FF",X"9F",X"0F",X"0F",X"9F",X"FF",X"FF",X"00",X"80",X"40",X"40",X"80",X"00",X"00",X"00",
		X"00",X"40",X"60",X"00",X"10",X"08",X"06",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"E0",X"78",X"1F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"0A",X"5F",X"79",X"0B",X"1E",X"04",X"17",X"03",X"00",X"01",X"03",X"00",X"00",X"00",X"00",
		X"DB",X"85",X"48",X"20",X"10",X"06",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"1F",X"7E",X"FE",X"FF",
		X"00",X"00",X"80",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"07",X"1F",X"7F",X"07",X"1F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",
		X"00",X"03",X"07",X"1F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"03",X"07",X"1F",X"7F",X"FF",X"1F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"F8",X"E0",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"40",X"40",X"40",X"40",X"40",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"04",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"C8",X"E8",X"E8",X"D8",X"B0",X"60",X"E0",X"C0",
		X"97",X"9C",X"9E",X"9B",X"8B",X"8D",X"87",X"C3",X"30",X"30",X"10",X"18",X"18",X"08",X"C8",X"68",
		X"F8",X"FC",X"FC",X"F2",X"BC",X"BE",X"B5",X"BF",X"A0",X"60",X"E0",X"E0",X"E0",X"60",X"60",X"30",
		X"DF",X"EE",X"CF",X"C7",X"EE",X"FC",X"FC",X"F8",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",
		X"0D",X"09",X"09",X"08",X"0D",X"0C",X"06",X"07",X"BF",X"DF",X"FD",X"DD",X"7B",X"7F",X"FF",X"F7",
		X"00",X"03",X"0C",X"B0",X"00",X"00",X"00",X"00",X"1E",X"7C",X"C0",X"00",X"00",X"00",X"C0",X"00",
		X"FF",X"FF",X"EF",X"01",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"C6",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"DE",X"FF",X"98",X"20",X"00",X"00",X"40",X"DB",X"3F",X"07",
		X"00",X"00",X"00",X"00",X"80",X"40",X"BC",X"FF",X"00",X"05",X"00",X"00",X"00",X"00",X"82",X"00",
		X"00",X"00",X"00",X"80",X"E0",X"F0",X"F8",X"FC",X"80",X"60",X"1C",X"04",X"07",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"E0",X"30",X"18",X"00",X"80",X"E0",X"E0",X"F0",X"FC",X"FE",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"E0",X"FC",X"3F",X"07",X"00",X"00",X"00",X"00",X"00",X"80",X"FF",X"FF",X"7F",X"03",X"00",
		X"00",X"00",X"00",X"E0",X"FC",X"F8",X"E0",X"00",X"E0",X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"80",X"E0",X"F8",X"FE",X"C0",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"80",X"F8",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"0F",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3E",X"3E",X"3E",X"3E",X"3D",X"30",X"06",X"FA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A8",X"80",X"80",X"06",X"1E",X"3E",X"3E",X"3E",X"3E",X"3E",X"3E",X"3E",X"3E",X"3E",X"3E",X"3E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"FC",
		X"00",X"00",X"00",X"00",X"F0",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FE",X"FF",X"FF",X"FF",X"01",
		X"00",X"00",X"00",X"00",X"80",X"E0",X"F0",X"FC",X"80",X"E0",X"F8",X"FE",X"7F",X"1F",X"07",X"01",
		X"FF",X"FF",X"1F",X"03",X"00",X"00",X"E0",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"80",X"C0",X"F0",X"F8",X"7E",X"3F",X"0F",X"80",X"C0",X"E0",X"70",X"38",X"1C",X"0E",X"87",
		X"00",X"00",X"00",X"00",X"80",X"C0",X"F0",X"F8",X"E0",X"F0",X"FC",X"7E",X"1F",X"0F",X"03",X"81",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"FC",X"FF",X"00",X"80",X"E0",X"F8",X"FE",X"7F",X"1F",X"07",
		X"80",X"FF",X"FF",X"FF",X"7F",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"1F",X"00",X"00",X"00",X"E0",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"3F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",
		X"FF",X"FF",X"F0",X"00",X"00",X"00",X"0F",X"FF",X"0F",X"FF",X"FF",X"FF",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"FF",X"FF",X"FF",X"F0",X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"FF",X"FF",
		X"00",X"00",X"07",X"3F",X"FF",X"FF",X"F8",X"C0",X"00",X"00",X"00",X"00",X"01",X"0F",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"3F",X"FF",X"FF",X"F8",X"C0",X"00",X"00",X"00",
		X"00",X"01",X"0F",X"FF",X"FF",X"FE",X"F0",X"00",X"00",X"00",X"00",X"00",X"07",X"3F",X"FF",X"FF",
		X"FF",X"C0",X"00",X"00",X"00",X"3F",X"FF",X"FF",X"FF",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"E0",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"0F",X"FF",X"FF",X"FF",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"3F",X"FF",X"FF",X"F8",X"C0",
		X"FE",X"F0",X"00",X"00",X"01",X"0F",X"FF",X"FF",X"FE",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"FF",X"FF",X"F8",X"C0",X"00",X"00",X"00",X"00",X"0F",X"7F",X"FF",X"FF",X"F0",X"80",X"00",
		X"FF",X"FF",X"FC",X"E0",X"00",X"00",X"03",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"FE",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"3F",X"07",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"FC",X"7E",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"C0",X"E0",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"0F",X"07",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"F8",X"00",X"00",X"00",X"00",X"E0",X"FC",X"FF",X"FF",
		X"00",X"C0",X"F8",X"FF",X"FF",X"FF",X"FF",X"F9",X"FF",X"FF",X"7F",X"1F",X"0F",X"07",X"03",X"81",
		X"C7",X"E1",X"F0",X"F8",X"FC",X"7E",X"3F",X"1F",X"0F",X"07",X"03",X"81",X"C0",X"E0",X"F0",X"F8",
		X"FC",X"7E",X"3F",X"1F",X"0F",X"07",X"03",X"01",X"3C",X"3C",X"3C",X"3C",X"3C",X"3E",X"3F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"F0",X"FC",X"E0",X"F0",X"F8",X"FC",X"FE",X"7F",X"3F",X"9F",
		X"CF",X"E7",X"F3",X"F9",X"FC",X"7E",X"3F",X"1F",X"C0",X"E0",X"F0",X"F8",X"FC",X"7E",X"3F",X"1F",
		X"3C",X"3E",X"3F",X"3F",X"3F",X"3F",X"3F",X"3D",X"3F",X"3F",X"3F",X"3D",X"3C",X"3C",X"3C",X"3C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"F0",X"F8",X"FC",X"FE",X"7F",X"3F",X"9F",
		X"FF",X"FF",X"FF",X"FB",X"FC",X"7E",X"3F",X"1F",X"00",X"00",X"00",X"00",X"C0",X"F0",X"FC",X"FF",
		X"00",X"E0",X"FC",X"FF",X"FF",X"7F",X"3F",X"1F",X"FF",X"FF",X"7F",X"8F",X"C1",X"E0",X"F0",X"F8",
		X"FF",X"7F",X"3F",X"1F",X"0F",X"07",X"03",X"81",X"1F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"7F",X"07",X"00",X"00",X"00",X"00",X"C1",X"FF",X"FF",X"BF",X"3F",X"00",X"00",X"00",
		X"80",X"FE",X"FF",X"FF",X"FF",X"03",X"00",X"00",X"F8",X"7C",X"7C",X"3E",X"3E",X"1F",X"1F",X"0F",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"F0",X"F0",X"F0",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"00",X"40",X"7E",X"40",X"00",X"5E",X"72",X"00",X"00",X"78",X"48",X"7E",X"00",X"7E",X"42",X"7E",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FE",X"D4",X"FA",X"A0",X"51",X"A2",X"08",X"FF",X"DF",X"16",X"AF",X"4D",X"1A",X"05",X"50",
		X"FF",X"7E",X"AE",X"54",X"29",X"88",X"22",X"49",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"CF",X"40",X"50",X"50",X"70",X"40",X"3F",X"00",X"00",X"00",X"02",X"03",X"40",X"40",X"FF",X"DF",
		X"00",X"00",X"43",X"C3",X"03",X"03",X"FF",X"FB",X"F2",X"06",X"0E",X"18",X"00",X"02",X"FC",X"00",
		X"5A",X"48",X"7E",X"7E",X"40",X"7E",X"7E",X"64",X"7E",X"7E",X"7E",X"7E",X"00",X"00",X"18",X"18",
		X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"6E",X"BB",X"77",X"DD",X"DD",X"77",X"BB",X"6E",
		X"FF",X"FF",X"D7",X"BD",X"D7",X"4B",X"81",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"F0",X"FF",X"F0",X"E1",X"ED",X"CC",X"0E",X"0F",X"07",
		X"F4",X"E6",X"EF",X"EF",X"CF",X"87",X"B1",X"BC",X"A7",X"B7",X"E7",X"EF",X"EF",X"EF",X"FF",X"FF",
		X"FF",X"F9",X"C1",X"F1",X"FC",X"F4",X"F6",X"F6",X"F9",X"F5",X"FD",X"E9",X"EB",X"A3",X"23",X"23",
		X"A2",X"DA",X"C8",X"89",X"01",X"01",X"1B",X"FF",X"07",X"07",X"CF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"9F",X"9F",X"8B",X"CA",X"C2",X"C0",X"C0",X"E9",X"FF",X"FF",X"CF",X"1F",X"7F",X"FD",X"FB",X"D3",
		X"FD",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"D2",X"99",X"1C",X"14",X"40",X"C0",X"F0",X"FF",
		X"EF",X"EF",X"C3",X"CB",X"9B",X"F9",X"FD",X"FD",X"FF",X"FF",X"DE",X"FF",X"FF",X"EF",X"FB",X"FF",
		X"FF",X"FB",X"7F",X"FF",X"FB",X"DF",X"FF",X"FF",X"BF",X"F5",X"FF",X"EF",X"FF",X"FA",X"BF",X"FF",
		X"00",X"00",X"00",X"00",X"87",X"80",X"83",X"87",X"00",X"00",X"00",X"00",X"FF",X"00",X"55",X"D5",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"9C",X"F6",X"00",X"00",X"00",X"00",X"FF",X"00",X"B9",X"EF",
		X"00",X"00",X"00",X"00",X"E0",X"30",X"90",X"D0",X"87",X"82",X"81",X"85",X"87",X"83",X"87",X"83",
		X"90",X"D0",X"90",X"90",X"D0",X"10",X"D0",X"D0",X"86",X"87",X"83",X"80",X"C0",X"60",X"30",X"1F",
		X"FE",X"FB",X"D3",X"02",X"00",X"00",X"00",X"FF",X"FB",X"FF",X"29",X"00",X"00",X"00",X"00",X"FF",
		X"7F",X"EB",X"D9",X"41",X"00",X"00",X"00",X"FF",X"D0",X"D0",X"90",X"00",X"00",X"00",X"00",X"E0",
		X"FF",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"3F",X"60",X"C1",X"83",X"87",X"86",X"84",X"80",X"FC",X"06",X"83",X"C1",X"E1",X"61",X"21",X"01",
		X"FF",X"1F",X"83",X"38",X"FC",X"F9",X"E3",X"DF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"9F",X"8F",
		X"FB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"B6",X"67",X"AA",X"75",X"56",X"EA",X"97",X"67",X"E5",X"22",X"54",X"DE",X"BB",X"FD",X"FF",
		X"B5",X"6D",X"C2",X"4E",X"D5",X"BF",X"FF",X"FF",X"6D",X"B7",X"4E",X"A8",X"B5",X"53",X"EF",X"FF",
		X"00",X"FF",X"CF",X"A7",X"08",X"15",X"42",X"E8",X"00",X"FF",X"FF",X"FF",X"00",X"4D",X"84",X"53",
		X"3C",X"BF",X"BF",X"BF",X"16",X"2D",X"91",X"66",X"00",X"FF",X"C0",X"FF",X"FF",X"FF",X"E0",X"FF",
		X"00",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"00",X"FF",X"03",X"FB",X"FB",X"FB",X"03",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F8",X"F8",X"18",X"18",X"18",X"18",X"18",X"00",X"00",X"7E",X"66",X"72",X"7A",
		X"7E",X"7E",X"40",X"7E",X"7E",X"72",X"5E",X"70",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C0",X"FF",X"EF",X"E8",X"EE",X"EE",X"EE",X"FE",
		X"C1",X"FC",X"BE",X"BE",X"BE",X"8E",X"FE",X"FF",X"C0",X"FF",X"EF",X"E1",X"FC",X"FE",X"8F",X"FF",
		X"C1",X"FC",X"BE",X"BE",X"BE",X"BE",X"CF",X"FF",X"8F",X"EF",X"EF",X"EF",X"EF",X"EF",X"E0",X"FF",
		X"E3",X"FB",X"BB",X"39",X"39",X"39",X"BB",X"FF",X"81",X"FC",X"8E",X"BE",X"BE",X"BE",X"BE",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"E0",X"00",X"00",X"00",X"01",X"0F",X"FF",
		X"00",X"0F",X"7F",X"F0",X"80",X"00",X"00",X"00",X"00",X"07",X"3F",X"F8",X"C0",X"00",X"00",X"07",
		X"FF",X"FF",X"FF",X"F6",X"C0",X"40",X"00",X"00",X"FF",X"FA",X"C0",X"00",X"00",X"00",X"01",X"0F",
		X"80",X"00",X"00",X"00",X"07",X"3F",X"F8",X"C0",X"00",X"00",X"0F",X"FF",X"F0",X"00",X"00",X"00",
		X"0F",X"FF",X"F0",X"00",X"00",X"00",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"F2",X"40",X"00",X"00",
		X"FF",X"FF",X"FA",X"40",X"00",X"00",X"00",X"00",X"F7",X"A0",X"00",X"00",X"00",X"00",X"0F",X"FF",
		X"00",X"00",X"00",X"00",X"0F",X"FF",X"F0",X"00",X"00",X"00",X"0F",X"FF",X"F0",X"00",X"00",X"00",
		X"0F",X"FF",X"F0",X"00",X"00",X"00",X"0F",X"FF",X"00",X"00",X"50",X"FB",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"80",X"E1",X"FF",X"FF",X"3F",X"00",X"00",X"00",X"00",X"80",X"E9",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"B5",X"00",X"FC",X"FE",X"07",X"03",X"01",X"00",X"00",
		X"00",X"00",X"00",X"03",X"17",X"FF",X"FF",X"FF",X"00",X"07",X"6F",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"F8",X"C0",X"00",X"00",X"07",X"3F",X"F8",X"C0",X"00",X"01",X"0F",X"FE",X"F0",X"00",X"00",X"00",
		X"3F",X"F8",X"C0",X"00",X"00",X"00",X"02",X"1F",X"00",X"00",X"00",X"00",X"05",X"6F",X"FF",X"FF",
		X"00",X"03",X"17",X"7F",X"FF",X"FF",X"FF",X"FF",X"FE",X"F0",X"00",X"00",X"01",X"0F",X"FE",X"F0",
		X"00",X"00",X"07",X"7F",X"F8",X"80",X"00",X"00",X"0F",X"FF",X"F0",X"00",X"00",X"00",X"00",X"07",
		X"F0",X"00",X"00",X"00",X"00",X"06",X"6F",X"FF",X"00",X"00",X"00",X"02",X"AF",X"FF",X"FF",X"FF",
		X"00",X"06",X"5F",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"00",X"00",X"0F",X"FF",X"F0",X"00",
		X"00",X"00",X"0F",X"FF",X"F0",X"00",X"00",X"00",X"0F",X"FF",X"F0",X"00",X"00",X"00",X"00",X"05",
		X"F0",X"00",X"00",X"00",X"00",X"02",X"CF",X"FF",X"00",X"00",X"00",X"00",X"16",X"DF",X"FF",X"FF",
		X"00",X"00",X"00",X"5D",X"FB",X"FF",X"FF",X"FF",X"01",X"00",X"4A",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"C0",X"00",X"00",X"00",X"3F",X"FF",X"C0",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"FC",X"FE",X"07",X"03",X"01",X"C0",X"C0",X"C8",X"F8",X"F6",X"FF",X"FF",X"FF",
		X"03",X"00",X"00",X"00",X"80",X"E8",X"FD",X"F9",X"FF",X"1F",X"00",X"00",X"00",X"00",X"40",X"ED",
		X"80",X"FF",X"7F",X"00",X"00",X"00",X"00",X"80",X"78",X"F4",X"F6",X"7E",X"7F",X"77",X"77",X"7F",
		X"0E",X"07",X"01",X"00",X"80",X"C0",X"F0",X"FC",X"01",X"80",X"E0",X"78",X"1E",X"07",X"01",X"00",
		X"FF",X"3F",X"03",X"00",X"00",X"C0",X"FC",X"3F",X"C0",X"E0",X"F0",X"E8",X"FC",X"FA",X"FF",X"FF",
		X"E0",X"70",X"1C",X"0E",X"03",X"01",X"00",X"C0",X"7E",X"3F",X"0F",X"07",X"81",X"C0",X"70",X"38",
		X"C0",X"E0",X"F0",X"E8",X"FC",X"FA",X"FD",X"FF",X"C3",X"61",X"30",X"18",X"0C",X"06",X"03",X"C1",
		X"00",X"80",X"E0",X"F0",X"F4",X"FE",X"FE",X"FF",X"C3",X"61",X"30",X"18",X"0C",X"06",X"03",X"81",
		X"C0",X"F0",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"0E",X"03",X"01",X"80",X"C0",X"E0",X"F8",X"FC",
		X"07",X"81",X"C0",X"70",X"38",X"0E",X"07",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"4A",X"EF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"60",X"F5",X"FF",X"FF",X"FF",
		X"1F",X"03",X"00",X"00",X"00",X"A0",X"F4",X"FF",X"80",X"E0",X"78",X"1E",X"07",X"01",X"00",X"00",
		X"7F",X"1F",X"0F",X"03",X"81",X"E0",X"70",X"1C",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"FE",X"FF",X"01",X"00",X"00",X"0F",X"00",X"00",X"00",X"F0",X"FF",X"0F",X"00",
		X"00",X"00",X"01",X"03",X"07",X"06",X"04",X"00",X"00",X"00",X"80",X"C0",X"E0",X"60",X"20",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"69",X"D6",X"F4",X"E0",X"F0",X"D4",X"80",
		X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"26",X"42",X"40",X"00",X"00",X"00",X"00",X"00",
		X"08",X"04",X"04",X"00",X"10",X"08",X"00",X"00",X"00",X"00",X"08",X"D0",X"68",X"E8",X"D0",X"D4",
		X"00",X"00",X"01",X"02",X"07",X"02",X"01",X"01",X"6C",X"F8",X"F2",X"FA",X"F4",X"71",X"7B",X"7A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",
		X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",
		X"44",X"CC",X"41",X"2F",X"77",X"23",X"63",X"FA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7A",X"7E",X"D8",X"7B",X"87",X"5A",X"B9",X"12",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"04",X"08",X"61",X"20",X"08",X"04",X"03",X"80",X"C0",X"72",X"3B",X"3B",X"72",X"C0",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"0F",X"1F",X"3F",X"3F",X"7F",X"7F",X"00",X"00",X"10",X"1C",X"38",X"1C",X"10",X"00",
		X"7F",X"7F",X"3F",X"3F",X"1F",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",X"20",X"18",X"00",X"00",
		X"00",X"10",X"1C",X"18",X"0C",X"10",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"69",X"69",X"69",X"69",X"69",X"69",X"69",X"69",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"BF",X"FF",X"FF",X"EF",X"FF",X"7F",X"FF",X"F7",X"FF",X"DF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"BB",X"FF",X"FF",X"F7",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"03",X"0F",X"1F",X"3F",X"3F",X"7F",X"7F",X"FF",X"C0",X"F0",X"F8",X"FC",X"FC",X"FE",X"FE",X"FF",
		X"FF",X"7F",X"7F",X"3F",X"3F",X"1F",X"0F",X"03",X"FF",X"FE",X"FE",X"FC",X"FC",X"F8",X"F0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"7F",X"00",X"0E",X"06",X"06",X"06",X"06",X"BE",X"BE",
		X"FF",X"F4",X"F4",X"F4",X"F4",X"F4",X"F4",X"F4",X"FF",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",
		X"F4",X"F4",X"F4",X"F4",X"F4",X"F4",X"F4",X"FF",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"FF",
		X"F4",X"F4",X"F4",X"F4",X"F4",X"F4",X"F4",X"F4",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",
		X"0C",X"17",X"29",X"5F",X"7D",X"3F",X"1F",X"0C",X"0C",X"17",X"21",X"41",X"41",X"21",X"17",X"0C",
		X"00",X"00",X"00",X"60",X"7F",X"7F",X"60",X"00",X"00",X"00",X"00",X"06",X"BE",X"BE",X"06",X"00",
		X"00",X"00",X"3E",X"7F",X"71",X"71",X"7F",X"7F",X"00",X"00",X"3E",X"BE",X"80",X"80",X"BE",X"BE",
		X"00",X"01",X"03",X"06",X"0C",X"18",X"30",X"60",X"80",X"C0",X"60",X"30",X"18",X"0C",X"06",X"03",
		X"C0",X"F8",X"08",X"09",X"0B",X"0B",X"0B",X"0B",X"01",X"07",X"04",X"F4",X"F4",X"04",X"F4",X"F4",
		X"00",X"1C",X"3C",X"7C",X"70",X"61",X"73",X"7F",X"00",X"3C",X"7E",X"FF",X"E7",X"C3",X"87",X"9F",
		X"BF",X"9E",X"00",X"3F",X"7F",X"7F",X"60",X"60",X"1E",X"1C",X"00",X"FF",X"FF",X"FF",X"C0",X"C0",
		X"00",X"FF",X"00",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"00",X"FF",X"00",X"FF",X"00",X"00",
		X"FF",X"91",X"00",X"6E",X"6E",X"00",X"91",X"FF",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",
		X"FD",X"A5",X"95",X"FD",X"A5",X"95",X"FD",X"C5",X"B7",X"FF",X"97",X"87",X"FF",X"87",X"CF",X"87",
		X"AD",X"C5",X"FD",X"F5",X"85",X"FD",X"B5",X"85",X"FF",X"87",X"AF",X"C7",X"FF",X"C7",X"BF",X"87",
		X"FD",X"95",X"05",X"6D",X"05",X"05",X"FD",X"55",X"05",X"FD",X"4D",X"45",X"15",X"95",X"FD",X"05",
		X"55",X"05",X"05",X"FD",X"3D",X"0D",X"E5",X"0D",X"05",X"CD",X"9D",X"05",X"05",X"FD",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",X"97",X"87",X"FF",X"07",X"FF",X"87",
		X"FD",X"AD",X"AD",X"FD",X"FD",X"55",X"55",X"05",X"B7",X"CF",X"FF",X"C7",X"BF",X"87",X"BF",X"87",
		X"3D",X"FD",X"05",X"05",X"FD",X"95",X"05",X"6D",X"05",X"05",X"FD",X"75",X"75",X"05",X"8D",X"FD",
		X"05",X"05",X"FD",X"8D",X"05",X"75",X"05",X"05",X"05",X"05",X"FD",X"F5",X"F5",X"05",X"05",X"FD",
		X"FF",X"81",X"00",X"7E",X"7E",X"00",X"81",X"FF",X"7F",X"3F",X"9F",X"CF",X"E7",X"FF",X"A7",X"CF",
		X"FF",X"9E",X"0E",X"6E",X"6E",X"60",X"70",X"FF",X"97",X"FF",X"97",X"87",X"FF",X"47",X"17",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"08",X"08",X"0B",X"0B",X"08",X"08",X"08",X"08",X"04",X"04",X"74",X"74",X"04",X"04",X"04",X"04",
		X"08",X"08",X"08",X"0F",X"00",X"00",X"00",X"00",X"04",X"04",X"04",X"FC",X"00",X"00",X"00",X"00",
		X"70",X"7F",X"3F",X"0F",X"00",X"1C",X"3C",X"7C",X"C0",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",
		X"70",X"60",X"60",X"70",X"7F",X"3F",X"1F",X"00",X"C3",X"C3",X"C3",X"07",X"FF",X"FE",X"FC",X"00",
		X"00",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"00",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"00",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",
		X"00",X"04",X"07",X"1D",X"7D",X"1D",X"07",X"04",X"00",X"0E",X"7C",X"B0",X"A0",X"B0",X"7C",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"7D",X"7D",X"7D",X"00",X"00",X"00",X"00",X"00",X"8E",X"8E",X"8E",
		X"00",X"00",X"3C",X"7C",X"71",X"71",X"7D",X"3C",X"00",X"00",X"3C",X"BE",X"8E",X"8E",X"3E",X"3C",
		X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"00",X"00",X"7D",X"7D",X"00",X"00",X"7D",X"7D",X"00",X"00",X"BC",X"BE",X"0E",X"0E",X"BE",X"BC",
		X"00",X"00",X"3C",X"7C",X"70",X"70",X"7D",X"3D",X"00",X"00",X"3C",X"3E",X"0E",X"0E",X"BE",X"BC",
		X"00",X"00",X"60",X"60",X"7D",X"7D",X"60",X"60",X"00",X"00",X"00",X"00",X"BE",X"BE",X"00",X"00",
		X"00",X"00",X"3D",X"7D",X"71",X"71",X"7D",X"3D",X"00",X"00",X"BE",X"BE",X"80",X"80",X"BE",X"BE",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"00",X"00",X"39",X"79",X"71",X"70",X"7D",X"3D",X"00",X"00",X"BE",X"BE",X"8E",X"0E",X"BE",X"BC",
		X"00",X"00",X"7D",X"7D",X"01",X"0D",X"7D",X"7D",X"00",X"00",X"BE",X"BE",X"B0",X"80",X"BE",X"BE",
		X"00",X"00",X"3D",X"7D",X"70",X"70",X"7D",X"3D",X"00",X"00",X"BC",X"BE",X"0E",X"0E",X"BE",X"BC",
		X"69",X"69",X"69",X"69",X"69",X"68",X"69",X"6B",X"22",X"14",X"48",X"80",X"40",X"32",X"00",X"00",
		X"6B",X"69",X"68",X"69",X"69",X"69",X"69",X"69",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"23",X"77",X"5D",X"EB",X"B7",X"7E",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"BE",X"CD",X"FF",X"7F",X"77",X"23",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"7F",X"7F",X"7F",X"7E",X"79",X"77",X"77",X"00",X"FF",X"FF",X"80",X"7F",X"FF",X"FF",X"FE",
		X"6F",X"5F",X"5F",X"5F",X"3F",X"3F",X"3F",X"3F",X"FC",X"F8",X"F0",X"E2",X"FE",X"FC",X"F8",X"F0",
		X"00",X"FF",X"FF",X"03",X"FC",X"43",X"7E",X"01",X"00",X"FE",X"FE",X"FE",X"FE",X"1E",X"E6",X"38",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",
		X"3F",X"3F",X"3F",X"3F",X"5F",X"5F",X"5F",X"6F",X"C3",X"FE",X"FC",X"E0",X"F0",X"FC",X"FE",X"FE",
		X"6F",X"77",X"79",X"7E",X"7F",X"7F",X"7F",X"00",X"FF",X"FF",X"FF",X"3F",X"C0",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"18",X"10",X"02",X"06",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"0C",
		X"01",X"FE",X"C3",X"F8",X"07",X"FF",X"FF",X"00",X"32",X"CE",X"3E",X"FE",X"FE",X"FE",X"FE",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"FF",X"FB",X"00",X"00",X"7B",X"03",X"83",X"FF",
		X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"40",X"00",X"00",X"00",X"23",X"3F",X"9F",X"8F",X"0D",X"02",X"05",X"02",X"01",X"C2",X"E0",X"F0",
		X"C7",X"E0",X"F0",X"60",X"21",X"03",X"E7",X"FF",X"F1",X"52",X"11",X"00",X"81",X"80",X"C2",X"E0",
		X"EF",X"EF",X"E7",X"E2",X"F0",X"F9",X"FF",X"CF",X"F0",X"E1",X"E2",X"40",X"00",X"00",X"C3",X"E0",
		X"E3",X"7F",X"3F",X"3E",X"00",X"4A",X"92",X"35",X"E2",X"C2",X"81",X"0A",X"53",X"A4",X"04",X"49",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"FF",X"F1",X"60",X"6E",X"6E",X"00",X"81",X"FF",
		X"FF",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FF",X"8F",X"07",X"77",X"77",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"36",X"3C",X"18",X"10",X"00",X"00",X"00",X"00",
		X"FE",X"FE",X"7E",X"7E",X"3E",X"3C",X"10",X"00",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",
		X"1F",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"FF",X"FF",X"7F",X"3F",X"1F",X"07",X"00",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"8C",X"84",X"FC",X"00",X"00",X"00",X"00",X"0F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"20",X"00",X"40",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"81",X"01",X"22",
		X"80",X"C0",X"E0",X"F0",X"F0",X"F8",X"FC",X"FC",X"FF",X"FF",X"3F",X"1F",X"0F",X"07",X"03",X"01",
		X"7F",X"7E",X"7C",X"7E",X"3E",X"3F",X"3F",X"1F",X"00",X"80",X"80",X"C0",X"C0",X"E0",X"F0",X"F8",
		X"1F",X"1F",X"1F",X"0F",X"0F",X"0F",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"80",X"FE",X"03",X"00",X"00",X"00",X"00",X"E0",X"3F",X"00",X"00",
		X"00",X"00",X"00",X"F8",X"0F",X"00",X"00",X"00",X"00",X"80",X"FE",X"03",X"00",X"00",X"00",X"00",
		X"22",X"23",X"A3",X"A1",X"3F",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"F0",X"FC",X"FE",X"FF",
		X"FF",X"FF",X"3F",X"00",X"0F",X"3F",X"3F",X"7F",X"FF",X"0F",X"00",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"03",X"00",X"00",X"07",X"0F",X"1F",X"1F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"FC",X"FC",X"BC",X"8C",X"CC",X"8C",X"0C",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"03",X"00",
		X"00",X"80",X"FF",X"FF",X"3F",X"00",X"00",X"00",X"80",X"C0",X"E1",X"01",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"03",X"00",X"00",X"00",X"00",X"00",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"F0",X"00",X"00",X"00",X"00",X"00",X"C0",X"FE",
		X"8F",X"80",X"C0",X"C0",X"C0",X"F0",X"FF",X"FF",X"1F",X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"7F",X"7F",X"7F",X"7F",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"18",X"FE",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"C0",X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"07",X"07",X"06",X"04",X"80",X"80",
		X"70",X"18",X"0C",X"06",X"03",X"01",X"C1",X"FF",X"60",X"C0",X"80",X"80",X"80",X"F0",X"FF",X"FF",
		X"20",X"20",X"22",X"23",X"23",X"23",X"23",X"23",X"00",X"00",X"00",X"00",X"C0",X"E0",X"E0",X"F0",
		X"FE",X"FC",X"00",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"C7",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",
		X"F9",X"FF",X"FF",X"FF",X"FF",X"1F",X"00",X"00",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"5B",X"BD",X"D5",X"F3",X"FB",X"FB",X"7E",
		X"04",X"2C",X"36",X"3F",X"0F",X"AF",X"7F",X"FF",X"FF",X"FF",X"7F",X"7F",X"FF",X"FF",X"DF",X"DF",
		X"00",X"8B",X"8B",X"EE",X"EF",X"F7",X"F7",X"FB",X"5F",X"3F",X"5F",X"3F",X"0F",X"1A",X"00",X"00",
		X"FB",X"FB",X"F1",X"F8",X"F8",X"F8",X"FC",X"BC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"BF",X"BF",X"3F",X"7E",X"6E",X"ED",X"FF",X"9C",X"B8",X"F8",X"78",X"79",X"FB",X"FB",X"F7",
		X"DF",X"9E",X"1E",X"3C",X"31",X"40",X"00",X"00",X"D6",X"F5",X"E0",X"C6",X"84",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",X"FF",X"FF",X"FF",X"E0",X"80",X"00",X"00",X"00",
		X"F0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"40",X"50",X"40",X"58",X"50",X"40",X"50",X"FF",X"00",X"3F",X"7F",X"FF",X"3F",X"7F",X"3D",
		X"40",X"5F",X"50",X"40",X"58",X"50",X"40",X"48",X"71",X"B2",X"23",X"60",X"60",X"20",X"20",X"20",
		X"50",X"56",X"40",X"40",X"53",X"50",X"40",X"48",X"E0",X"60",X"20",X"20",X"60",X"3F",X"7F",X"3F",
		X"50",X"56",X"44",X"40",X"40",X"50",X"40",X"7F",X"7F",X"3F",X"3F",X"3F",X"7F",X"FF",X"00",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"F8",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"F0",X"F0",X"F8",X"F8",X"FC",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"FF",X"FF",X"FF",X"FF",X"0F",X"E0",X"FE",X"FF",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FE",X"FC",X"FD",X"F9",X"FB",X"F3",X"F7",
		X"00",X"80",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"80",X"F8",X"FF",X"FF",X"FF",
		X"03",X"03",X"03",X"03",X"03",X"03",X"77",X"07",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FC",X"F9",
		X"07",X"77",X"77",X"07",X"07",X"77",X"77",X"07",X"F1",X"F1",X"E1",X"E1",X"E0",X"E1",X"E1",X"F1",
		X"F1",X"F9",X"FC",X"FE",X"00",X"67",X"FF",X"F7",X"FF",X"FF",X"FF",X"00",X"00",X"69",X"F7",X"BF",
		X"FF",X"FF",X"95",X"FF",X"FF",X"4E",X"F7",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"0F",
		X"0F",X"0F",X"1F",X"1F",X"00",X"1F",X"1F",X"0F",X"78",X"D0",X"F0",X"60",X"80",X"E0",X"FC",X"FE",
		X"3C",X"3C",X"3C",X"3C",X"3C",X"3F",X"3F",X"3F",X"EF",X"FF",X"DF",X"FD",X"FF",X"BB",X"49",X"00",
		X"03",X"07",X"3F",X"7D",X"FF",X"FD",X"EE",X"F8",X"17",X"1F",X"0F",X"1D",X"0F",X"0F",X"1B",X"0F",
		X"0F",X"0F",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FB",X"FC",X"D1",X"E7",X"4D",X"D7",X"9F",X"AF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"00",X"00",X"38",X"FE",X"FF",X"FF",
		X"03",X"07",X"07",X"07",X"0F",X"0F",X"0E",X"0E",X"FF",X"FF",X"C7",X"83",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"C0",X"C0",X"E0",X"F0",X"F8",X"7C",X"3C",X"00",X"00",X"00",X"00",X"00",X"70",X"F8",X"F8",
		X"0E",X"0E",X"0F",X"07",X"07",X"07",X"03",X"03",X"00",X"00",X"00",X"00",X"80",X"CC",X"FE",X"FE",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FE",X"FC",X"38",X"00",X"00",X"00",X"00",
		X"1C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"F8",X"70",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"7E",X"7F",X"60",X"7F",X"71",X"7E",X"6E",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F9",
		X"62",X"7F",X"7F",X"60",X"7F",X"6F",X"60",X"7F",X"E3",X"EF",X"CF",X"9F",X"BE",X"04",X"60",X"73",
		X"AF",X"AF",X"A7",X"E7",X"80",X"07",X"8F",X"8F",X"80",X"80",X"80",X"80",X"00",X"00",X"80",X"C0",
		X"C7",X"E0",X"F0",X"60",X"21",X"03",X"E7",X"FF",X"E0",X"40",X"00",X"00",X"80",X"80",X"C0",X"E0",
		X"7F",X"60",X"7E",X"62",X"7E",X"7F",X"60",X"7F",X"7F",X"FF",X"E7",X"81",X"81",X"84",X"C7",X"C3",
		X"65",X"7C",X"7F",X"6E",X"62",X"7F",X"7F",X"7F",X"E0",X"E0",X"F0",X"FC",X"FF",X"FF",X"FF",X"FF",
		X"EF",X"EF",X"E7",X"E2",X"F0",X"F9",X"FF",X"CF",X"F0",X"E0",X"E0",X"40",X"00",X"00",X"C0",X"E0",
		X"E3",X"7F",X"3F",X"3E",X"80",X"8B",X"CB",X"DB",X"E0",X"C0",X"80",X"00",X"C0",X"C0",X"C0",X"C0",
		X"0F",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"FC",X"04",X"04",X"04",X"04",X"04",X"04",X"04",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",
		X"00",X"1C",X"3C",X"7C",X"70",X"61",X"73",X"7F",X"00",X"3C",X"7E",X"FF",X"E7",X"C3",X"87",X"9F",
		X"3F",X"1E",X"00",X"3F",X"7F",X"7F",X"60",X"60",X"1E",X"1C",X"00",X"FF",X"FF",X"FF",X"C0",X"C0",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"0F",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"FC",
		X"70",X"7F",X"3F",X"0F",X"00",X"1C",X"3C",X"7C",X"C0",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",
		X"70",X"60",X"60",X"70",X"7F",X"3F",X"1F",X"00",X"C3",X"C3",X"C3",X"07",X"FF",X"FE",X"FC",X"00",
		X"00",X"38",X"30",X"20",X"20",X"20",X"36",X"20",X"00",X"9F",X"3F",X"7F",X"1F",X"3F",X"DF",X"1B",
		X"20",X"20",X"36",X"24",X"20",X"20",X"30",X"38",X"1D",X"3C",X"1E",X"1F",X"1F",X"3F",X"7F",X"1F",
		X"00",X"FF",X"FE",X"DF",X"DF",X"CF",X"CF",X"E7",X"00",X"FC",X"FC",X"FC",X"7C",X"7C",X"7C",X"3C",
		X"E7",X"E2",X"30",X"10",X"88",X"C0",X"E0",X"80",X"3C",X"3C",X"1C",X"1C",X"0C",X"0C",X"0C",X"0C",
		X"30",X"20",X"20",X"20",X"38",X"30",X"20",X"20",X"1F",X"3F",X"1C",X"3B",X"1F",X"1F",X"3F",X"1F",
		X"20",X"38",X"30",X"20",X"20",X"20",X"3F",X"00",X"3F",X"3F",X"1F",X"1F",X"1F",X"3F",X"FF",X"00",
		X"00",X"30",X"F8",X"F0",X"F1",X"E3",X"E6",X"CE",X"0C",X"0C",X"1C",X"1C",X"3C",X"3C",X"7C",X"7C",
		X"DE",X"BE",X"FE",X"7E",X"FF",X"FB",X"FF",X"00",X"7C",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"00",
		X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FE",X"02",X"FA",X"EA",X"CA",X"8A",X"0A",X"0A",
		X"FB",X"FB",X"2B",X"0B",X"EB",X"EB",X"EB",X"EB",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"F0",X"F8",X"1F",X"0F",X"07",X"03",X"00",X"00",X"00",X"00",
		X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"80",X"E0",X"FF",X"FF",X"FF",X"FF",
		X"EB",X"EB",X"EB",X"EA",X"08",X"F8",X"FB",X"FE",X"8A",X"8A",X"9A",X"0A",X"0A",X"1A",X"3A",X"0A",
		X"FC",X"FC",X"FE",X"FC",X"FC",X"FF",X"00",X"FF",X"0A",X"1A",X"0A",X"0A",X"1A",X"FA",X"02",X"FE",
		X"60",X"7E",X"7E",X"60",X"7E",X"60",X"7C",X"6A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"62",X"3E",X"1F",X"00",X"7F",X"6F",X"60",X"7F",X"00",X"00",X"00",X"80",X"E0",X"F0",X"B4",X"BE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"02",X"08",X"5A",
		X"7F",X"60",X"7E",X"62",X"7E",X"7F",X"70",X"7F",X"BF",X"3D",X"3D",X"3D",X"3D",X"39",X"B8",X"F0",
		X"64",X"7E",X"7F",X"6A",X"62",X"7F",X"7F",X"73",X"E0",X"E0",X"C0",X"C0",X"80",X"80",X"80",X"80",
		X"43",X"61",X"72",X"D1",X"C2",X"01",X"01",X"00",X"FE",X"FE",X"BE",X"2C",X"2E",X"3E",X"14",X"3A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"32",X"0E",X"1E",X"14",X"0E",X"04",X"02",X"0A",
		X"60",X"01",X"00",X"01",X"20",X"71",X"78",X"79",X"BF",X"70",X"A0",X"6F",X"A0",X"7F",X"B1",X"6E",
		X"38",X"09",X"08",X"01",X"00",X"01",X"00",X"01",X"AE",X"60",X"B1",X"7F",X"A0",X"7F",X"AF",X"60",
		X"E5",X"E7",X"F7",X"F7",X"FD",X"FF",X"E6",X"E6",X"8E",X"1E",X"9E",X"9E",X"CE",X"4E",X"DE",X"8E",
		X"FF",X"F7",X"FD",X"E7",X"E7",X"EF",X"F7",X"EE",X"1E",X"9E",X"1E",X"8E",X"9E",X"4E",X"8E",X"9E",
		X"00",X"01",X"00",X"01",X"10",X"31",X"70",X"79",X"AF",X"7F",X"A0",X"7E",X"A0",X"60",X"BF",X"70",
		X"38",X"11",X"00",X"01",X"20",X"61",X"70",X"79",X"AD",X"60",X"B8",X"7F",X"AE",X"60",X"B1",X"7F",
		X"E7",X"F7",X"F7",X"F7",X"EF",X"FF",X"F7",X"E7",X"DE",X"CE",X"6E",X"AE",X"CE",X"4E",X"8E",X"9E",
		X"F6",X"F7",X"F7",X"CF",X"DF",X"D7",X"EF",X"E6",X"9E",X"CE",X"AE",X"CE",X"6E",X"CE",X"8E",X"CE",
		X"00",X"3A",X"3A",X"00",X"3A",X"3A",X"00",X"32",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"3E",X"3E",X"00",X"22",X"22",X"3E",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"04",X"18",X"38",X"38",X"38",X"3C",X"00",X"00",X"00",X"20",X"B0",X"90",X"90",X"00",
		X"2C",X"04",X"04",X"00",X"08",X"1C",X"1C",X"38",X"40",X"40",X"00",X"40",X"60",X"68",X"48",X"18",
		X"00",X"2A",X"2A",X"3E",X"3E",X"00",X"3E",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3E",X"3E",X"00",X"22",X"22",X"3E",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3B",X"37",X"37",X"AF",X"8E",X"4C",X"59",X"3A",X"38",X"28",X"28",X"18",X"08",X"C0",X"80",X"60",
		X"AB",X"7A",X"02",X"02",X"00",X"00",X"00",X"00",X"10",X"90",X"F0",X"60",X"00",X"00",X"00",X"00",
		X"00",X"00",X"1F",X"1F",X"1C",X"1F",X"10",X"10",X"00",X"00",X"EF",X"EF",X"2F",X"AF",X"2F",X"3F",
		X"10",X"1F",X"1C",X"18",X"10",X"16",X"17",X"18",X"0F",X"EF",X"2F",X"3E",X"1D",X"4F",X"7F",X"1F",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"00",X"00",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"F8",X"86",X"71",X"FD",X"E2",X"F8",X"FD",X"9D",X"F8",X"78",X"78",X"20",X"B0",X"B0",X"30",X"20",
		X"1F",X"18",X"14",X"17",X"10",X"10",X"18",X"1D",X"EF",X"6F",X"2E",X"AD",X"3F",X"3E",X"0F",X"EF",
		X"14",X"14",X"17",X"10",X"10",X"18",X"00",X"00",X"2F",X"2F",X"AF",X"3F",X"3F",X"7F",X"00",X"00",
		X"8D",X"87",X"C7",X"FF",X"3B",X"8E",X"71",X"87",X"A0",X"A0",X"80",X"C8",X"F8",X"F8",X"F8",X"F8",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"00",X"00",
		X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"EF",X"FF",X"FD",X"FF",X"FF",X"FF",X"F7",X"7F",X"FF",X"FE",
		X"FF",X"FB",X"FF",X"FD",X"DF",X"FF",X"7D",X"FF",X"FF",X"FB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"BF",X"FF",X"FF",X"DF",
		X"FF",X"FF",X"FF",X"FF",X"BE",X"8F",X"E7",X"63",X"FF",X"FF",X"F7",X"FF",X"FD",X"FF",X"DF",X"FF",
		X"63",X"F7",X"96",X"7F",X"FD",X"FB",X"FF",X"EF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FA",X"FF",X"FB",X"FD",X"FD",X"FF",X"FB",X"FD",X"AF",X"4F",X"A7",X"D7",X"A3",X"D3",X"E9",X"D1",
		X"FD",X"FC",X"FC",X"FC",X"FE",X"FF",X"FF",X"FF",X"81",X"01",X"13",X"03",X"07",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"F1",X"E0",X"DA",X"D5",X"EA",X"7D",X"6A",X"2D",X"B6",X"BD",X"DE",X"DE",
		X"FD",X"EF",X"C1",X"C1",X"D9",X"80",X"A2",X"A2",X"C8",X"86",X"3D",X"5D",X"B0",X"C0",X"BE",X"FF",
		X"00",X"00",X"00",X"02",X"05",X"28",X"20",X"29",X"00",X"00",X"00",X"40",X"A0",X"10",X"08",X"10",
		X"23",X"2B",X"61",X"30",X"39",X"1C",X"0F",X"02",X"00",X"90",X"88",X"00",X"80",X"00",X"E0",X"00",
		X"AA",X"A2",X"84",X"D8",X"C1",X"E2",X"FF",X"FB",X"9B",X"D2",X"E0",X"39",X"9D",X"3D",X"87",X"C7",
		X"7F",X"3F",X"BF",X"3F",X"9F",X"5F",X"9F",X"4F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"02",X"03",X"03",X"01",X"00",X"02",X"01",X"62",X"94",X"AD",X"A5",X"91",X"CB",X"0A",X"0B",
		X"05",X"04",X"04",X"0E",X"0E",X"18",X"03",X"1D",X"40",X"82",X"C7",X"77",X"6F",X"AF",X"1F",X"9F",
		X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"03",X"05",X"38",X"6F",X"2F",X"6B",X"51",X"F6",X"EE",
		X"02",X"0E",X"0B",X"03",X"1D",X"03",X"1B",X"1F",X"E5",X"7A",X"98",X"30",X"61",X"53",X"E7",X"A7",
		X"90",X"56",X"AA",X"33",X"CB",X"DA",X"96",X"0C",X"9F",X"7C",X"E0",X"80",X"00",X"00",X"00",X"05",
		X"2C",X"B8",X"98",X"98",X"50",X"31",X"91",X"13",X"0D",X"1B",X"39",X"3F",X"6F",X"5D",X"7B",X"37",
		X"AC",X"C2",X"40",X"30",X"60",X"9E",X"D0",X"04",X"B4",X"00",X"C0",X"00",X"00",X"00",X"02",X"17",
		X"70",X"28",X"80",X"58",X"D0",X"21",X"A3",X"03",X"1F",X"CF",X"6F",X"3F",X"3E",X"84",X"E0",X"F3",
		X"E7",X"E5",X"A2",X"24",X"44",X"60",X"AA",X"68",X"7F",X"2B",X"7F",X"2D",X"3F",X"95",X"1D",X"0F",
		X"55",X"F4",X"96",X"2A",X"A3",X"75",X"2E",X"6D",X"07",X"00",X"84",X"44",X"31",X"8A",X"C1",X"78",
		X"A7",X"07",X"23",X"F1",X"00",X"10",X"80",X"58",X"FF",X"FF",X"E7",X"81",X"01",X"04",X"07",X"03",
		X"20",X"86",X"08",X"61",X"16",X"34",X"8D",X"40",X"00",X"00",X"00",X"00",X"88",X"65",X"00",X"59",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"9F",X"9F",X"8F",X"00",X"80",X"E0",X"FC",X"FF",X"FF",X"FF",X"FF",
		X"C7",X"C3",X"80",X"40",X"80",X"C0",X"80",X"80",X"FF",X"FF",X"FF",X"1F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"06",X"07",X"03",X"01",X"00",X"00",
		X"FF",X"00",X"FF",X"EE",X"FE",X"DC",X"EE",X"FE",X"FF",X"00",X"FF",X"EE",X"FE",X"DC",X"EE",X"FE",
		X"07",X"1C",X"21",X"43",X"47",X"87",X"8F",X"8F",X"DB",X"35",X"DA",X"EA",X"ED",X"F5",X"F5",X"F5");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
