library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity prog is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of prog is
	type rom is array(0 to  24575) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"3E",X"00",X"32",X"84",X"7D",X"C3",X"66",X"02",X"3A",X"07",X"60",X"0F",X"D0",X"33",X"33",X"C9",
		X"3A",X"00",X"62",X"0F",X"D8",X"33",X"33",X"C9",X"21",X"09",X"60",X"35",X"C8",X"33",X"33",X"C9",
		X"21",X"08",X"60",X"35",X"28",X"F2",X"E1",X"C9",X"87",X"E1",X"5F",X"16",X"00",X"C3",X"32",X"00",
		X"18",X"12",X"19",X"5E",X"23",X"56",X"EB",X"E9",X"C3",X"36",X"57",X"06",X"0A",X"C3",X"2B",X"57",
		X"19",X"10",X"FA",X"C9",X"21",X"27",X"62",X"46",X"0F",X"10",X"FD",X"D8",X"E1",X"C9",X"11",X"08",
		X"69",X"01",X"28",X"00",X"ED",X"B0",X"C9",X"3A",X"18",X"60",X"21",X"1A",X"60",X"86",X"21",X"19",
		X"60",X"86",X"32",X"18",X"60",X"C9",X"F5",X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",X"AF",X"32",
		X"84",X"7D",X"3A",X"00",X"7D",X"E6",X"01",X"C2",X"03",X"80",X"21",X"38",X"01",X"CD",X"41",X"01",
		X"3A",X"07",X"60",X"A7",X"C2",X"B5",X"00",X"3A",X"26",X"60",X"A7",X"C2",X"98",X"00",X"3A",X"0E",
		X"60",X"A7",X"3A",X"80",X"7C",X"C2",X"9B",X"00",X"3A",X"00",X"7C",X"47",X"E6",X"0F",X"4F",X"3A",
		X"11",X"60",X"2F",X"A0",X"E6",X"10",X"17",X"17",X"17",X"B1",X"60",X"6F",X"22",X"10",X"60",X"78",
		X"CB",X"77",X"C2",X"00",X"00",X"21",X"1A",X"60",X"35",X"CD",X"57",X"00",X"CD",X"7B",X"01",X"CD",
		X"E0",X"00",X"21",X"D2",X"00",X"E5",X"3A",X"05",X"60",X"EF",X"C3",X"01",X"3C",X"07",X"B2",X"08",
		X"FE",X"06",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"3E",X"01",X"32",X"84",X"7D",X"F1",X"C9",
		X"21",X"80",X"60",X"11",X"00",X"7D",X"3A",X"07",X"60",X"A7",X"C0",X"06",X"07",X"7E",X"A7",X"CA",
		X"F5",X"00",X"35",X"3E",X"01",X"12",X"1C",X"2C",X"10",X"F3",X"CD",X"31",X"38",X"7E",X"A7",X"C2",
		X"08",X"01",X"2D",X"2D",X"7E",X"C3",X"0B",X"01",X"35",X"2D",X"7E",X"32",X"00",X"7C",X"21",X"88",
		X"60",X"AF",X"BE",X"CA",X"18",X"01",X"35",X"3C",X"CD",X"2F",X"0C",X"C9",X"06",X"08",X"AF",X"21",
		X"00",X"7D",X"11",X"80",X"60",X"77",X"12",X"2C",X"1C",X"10",X"FA",X"06",X"05",X"12",X"1C",X"10",
		X"FC",X"32",X"80",X"7D",X"CD",X"8D",X"2E",X"C9",X"53",X"00",X"69",X"80",X"41",X"00",X"70",X"80",
		X"81",X"AF",X"32",X"85",X"7D",X"7E",X"32",X"08",X"78",X"23",X"7E",X"32",X"00",X"78",X"23",X"7E",
		X"32",X"00",X"78",X"23",X"7E",X"32",X"01",X"78",X"23",X"7E",X"32",X"01",X"78",X"23",X"7E",X"32",
		X"02",X"78",X"23",X"7E",X"32",X"02",X"78",X"23",X"7E",X"32",X"03",X"78",X"23",X"7E",X"32",X"03",
		X"78",X"3E",X"01",X"32",X"85",X"7D",X"AF",X"32",X"85",X"7D",X"C9",X"3A",X"00",X"7D",X"CB",X"7F",
		X"21",X"03",X"60",X"C2",X"89",X"01",X"36",X"01",X"C9",X"7E",X"A7",X"C8",X"E5",X"3A",X"05",X"60",
		X"FE",X"03",X"CA",X"9D",X"01",X"CD",X"1C",X"01",X"3E",X"03",X"32",X"85",X"60",X"E1",X"36",X"00",
		X"2B",X"34",X"11",X"24",X"60",X"1A",X"96",X"C0",X"77",X"13",X"2B",X"EB",X"1A",X"FE",X"90",X"D0",
		X"86",X"27",X"12",X"11",X"00",X"04",X"CD",X"9F",X"30",X"C9",X"00",X"37",X"00",X"AA",X"AA",X"AA",
		X"00",X"18",X"01",X"CD",X"74",X"08",X"21",X"BA",X"01",X"11",X"B2",X"60",X"01",X"09",X"00",X"ED",
		X"B0",X"3E",X"01",X"32",X"07",X"60",X"32",X"29",X"62",X"32",X"28",X"62",X"CD",X"B8",X"06",X"CD",
		X"07",X"02",X"3E",X"01",X"32",X"82",X"7D",X"32",X"05",X"60",X"32",X"27",X"62",X"AF",X"32",X"0A",
		X"60",X"CD",X"53",X"0A",X"11",X"04",X"03",X"CD",X"9F",X"30",X"11",X"02",X"02",X"CD",X"9F",X"30",
		X"11",X"00",X"02",X"CD",X"9F",X"30",X"C9",X"3A",X"80",X"7D",X"4F",X"21",X"20",X"60",X"E6",X"03",
		X"C6",X"03",X"77",X"23",X"79",X"0F",X"0F",X"E6",X"03",X"47",X"3E",X"10",X"CA",X"26",X"02",X"3E",
		X"0A",X"C6",X"05",X"27",X"10",X"FB",X"77",X"23",X"79",X"01",X"01",X"01",X"11",X"02",X"01",X"E6",
		X"70",X"17",X"17",X"17",X"17",X"CA",X"47",X"02",X"DA",X"41",X"02",X"3C",X"4F",X"5A",X"C3",X"47",
		X"02",X"C6",X"02",X"47",X"57",X"87",X"5F",X"72",X"23",X"73",X"23",X"70",X"23",X"71",X"23",X"3A",
		X"80",X"7D",X"07",X"3E",X"01",X"DA",X"59",X"02",X"3D",X"77",X"21",X"65",X"35",X"11",X"00",X"61",
		X"01",X"AA",X"00",X"ED",X"B0",X"C9",X"06",X"10",X"21",X"00",X"60",X"AF",X"4F",X"77",X"23",X"0D",
		X"20",X"FB",X"10",X"F8",X"06",X"04",X"21",X"00",X"70",X"4F",X"77",X"23",X"0D",X"20",X"FB",X"10",
		X"F8",X"06",X"04",X"3E",X"10",X"21",X"00",X"74",X"0E",X"00",X"77",X"23",X"0D",X"20",X"FB",X"10",
		X"F7",X"21",X"C0",X"60",X"06",X"40",X"3E",X"FF",X"77",X"23",X"10",X"FC",X"3E",X"C0",X"32",X"B0",
		X"60",X"32",X"B1",X"60",X"AF",X"32",X"83",X"7D",X"32",X"86",X"7D",X"32",X"87",X"7D",X"3C",X"32",
		X"82",X"7D",X"C3",X"12",X"12",X"CD",X"1C",X"01",X"3E",X"01",X"32",X"84",X"7D",X"26",X"60",X"3A",
		X"B1",X"60",X"6F",X"7E",X"87",X"30",X"1C",X"CD",X"15",X"03",X"CD",X"50",X"03",X"21",X"19",X"60",
		X"34",X"21",X"83",X"63",X"3A",X"1A",X"60",X"BE",X"28",X"E3",X"77",X"CD",X"7F",X"03",X"CD",X"A2",
		X"03",X"18",X"DA",X"E6",X"1F",X"5F",X"16",X"00",X"36",X"FF",X"2C",X"4E",X"36",X"FF",X"2C",X"7D",
		X"FE",X"C0",X"30",X"02",X"3E",X"C0",X"32",X"B1",X"60",X"79",X"21",X"BD",X"02",X"E5",X"21",X"07",
		X"03",X"19",X"5E",X"23",X"56",X"EB",X"E9",X"1C",X"05",X"9B",X"05",X"C6",X"05",X"E9",X"05",X"11",
		X"06",X"2A",X"06",X"B8",X"06",X"3A",X"1A",X"60",X"47",X"E6",X"0F",X"C0",X"CF",X"3A",X"0D",X"60",
		X"CD",X"47",X"03",X"11",X"E0",X"FF",X"CB",X"60",X"28",X"14",X"3E",X"10",X"77",X"19",X"77",X"19",
		X"77",X"3A",X"0F",X"60",X"A7",X"C8",X"3A",X"0D",X"60",X"EE",X"01",X"CD",X"47",X"03",X"3C",X"77",
		X"19",X"36",X"25",X"19",X"36",X"20",X"C9",X"21",X"40",X"77",X"A7",X"C8",X"21",X"E0",X"74",X"C9",
		X"3A",X"2D",X"62",X"A7",X"C0",X"21",X"B3",X"60",X"3A",X"0D",X"60",X"A7",X"28",X"03",X"21",X"B6",
		X"60",X"7E",X"E6",X"F0",X"47",X"23",X"7E",X"E6",X"0F",X"B0",X"0F",X"0F",X"0F",X"0F",X"21",X"21",
		X"60",X"BE",X"D8",X"3E",X"01",X"32",X"2D",X"62",X"21",X"28",X"62",X"34",X"C3",X"B8",X"06",X"21",
		X"84",X"63",X"7E",X"34",X"A7",X"C0",X"21",X"81",X"63",X"7E",X"47",X"34",X"E6",X"07",X"C0",X"78",
		X"0F",X"0F",X"0F",X"47",X"CD",X"5B",X"56",X"80",X"FE",X"03",X"38",X"02",X"3E",X"05",X"32",X"80",
		X"63",X"C9",X"3E",X"03",X"F7",X"D7",X"3A",X"50",X"63",X"0F",X"D8",X"21",X"B8",X"62",X"35",X"C0",
		X"36",X"04",X"3A",X"B9",X"62",X"0F",X"D0",X"21",X"29",X"6A",X"06",X"40",X"DD",X"21",X"A0",X"66",
		X"0F",X"D2",X"E4",X"03",X"DD",X"36",X"09",X"02",X"DD",X"36",X"0A",X"02",X"04",X"04",X"CD",X"F2",
		X"03",X"21",X"BA",X"62",X"35",X"C0",X"3E",X"01",X"32",X"B9",X"62",X"32",X"A0",X"63",X"3E",X"10",
		X"32",X"BA",X"62",X"C9",X"DD",X"36",X"09",X"02",X"DD",X"36",X"0A",X"00",X"CD",X"F2",X"03",X"C3",
		X"DE",X"03",X"70",X"3A",X"19",X"60",X"0F",X"D8",X"04",X"70",X"C9",X"C9",X"38",X"95",X"00",X"48",
		X"A1",X"43",X"0B",X"87",X"A1",X"43",X"0B",X"97",X"99",X"6C",X"07",X"9D",X"A9",X"08",X"07",X"9D",
		X"AF",X"CD",X"36",X"0B",X"3C",X"32",X"86",X"7D",X"11",X"12",X"38",X"CD",X"A7",X"0D",X"3E",X"10",
		X"32",X"57",X"76",X"32",X"B7",X"75",X"21",X"D0",X"27",X"11",X"30",X"69",X"01",X"08",X"00",X"ED",
		X"B0",X"21",X"D8",X"27",X"11",X"0C",X"6A",X"01",X"10",X"00",X"ED",X"B0",X"21",X"5C",X"38",X"CD",
		X"4E",X"00",X"3A",X"19",X"69",X"F6",X"80",X"32",X"1D",X"69",X"3A",X"21",X"69",X"F6",X"80",X"32",
		X"25",X"69",X"21",X"08",X"69",X"11",X"04",X"00",X"01",X"54",X"0A",X"CD",X"3D",X"00",X"21",X"E8",
		X"27",X"11",X"1C",X"6A",X"01",X"08",X"00",X"ED",X"B0",X"21",X"0B",X"69",X"11",X"04",X"00",X"01",
		X"A0",X"0A",X"CD",X"3D",X"00",X"3E",X"3F",X"32",X"8E",X"63",X"AF",X"32",X"AF",X"62",X"21",X"CB",
		X"0B",X"11",X"00",X"69",X"01",X"08",X"00",X"ED",X"B0",X"3E",X"40",X"32",X"09",X"60",X"21",X"85",
		X"63",X"34",X"22",X"C0",X"63",X"C9",X"21",X"AF",X"62",X"34",X"7E",X"CB",X"47",X"C0",X"E6",X"07",
		X"FE",X"06",X"F5",X"21",X"19",X"6A",X"28",X"04",X"7E",X"EE",X"0E",X"77",X"2B",X"35",X"F1",X"21",
		X"15",X"6A",X"28",X"04",X"7E",X"EE",X"0E",X"77",X"2B",X"35",X"7E",X"FE",X"9E",X"D0",X"21",X"00",
		X"69",X"11",X"04",X"00",X"01",X"FF",X"0C",X"CD",X"3D",X"00",X"3A",X"08",X"69",X"FE",X"37",X"D0",
		X"3E",X"30",X"C3",X"8B",X"04",X"21",X"AF",X"62",X"35",X"7E",X"11",X"82",X"39",X"FE",X"80",X"28",
		X"12",X"11",X"5A",X"39",X"FE",X"50",X"28",X"0B",X"11",X"5C",X"38",X"FE",X"30",X"28",X"04",X"A7",
		X"28",X"0F",X"C9",X"EB",X"D5",X"CD",X"4E",X"00",X"21",X"83",X"60",X"36",X"03",X"D1",X"1A",X"A7",
		X"C0",X"21",X"85",X"63",X"34",X"C9",X"AF",X"32",X"85",X"63",X"21",X"09",X"60",X"34",X"23",X"36",
		X"0A",X"C9",X"00",X"00",X"06",X"03",X"77",X"19",X"3D",X"10",X"FB",X"C9",X"4F",X"CF",X"CD",X"5F",
		X"05",X"C3",X"B9",X"11",X"4F",X"21",X"29",X"35",X"06",X"00",X"09",X"A7",X"06",X"03",X"1A",X"8E",
		X"27",X"12",X"13",X"23",X"10",X"F8",X"D5",X"1B",X"3A",X"0D",X"60",X"CD",X"6B",X"05",X"D1",X"1B",
		X"21",X"BA",X"60",X"06",X"03",X"1A",X"BE",X"D8",X"C2",X"50",X"05",X"1B",X"2B",X"10",X"F6",X"C9",
		X"CD",X"5F",X"05",X"21",X"B8",X"60",X"1A",X"77",X"13",X"23",X"10",X"FA",X"C3",X"DA",X"05",X"11",
		X"B2",X"60",X"3A",X"0D",X"60",X"A7",X"C8",X"11",X"B5",X"60",X"C9",X"DD",X"21",X"81",X"77",X"A7",
		X"28",X"0A",X"DD",X"21",X"21",X"75",X"18",X"04",X"DD",X"21",X"41",X"76",X"EB",X"11",X"E0",X"FF",
		X"01",X"04",X"03",X"7E",X"0F",X"0F",X"0F",X"0F",X"CD",X"93",X"05",X"7E",X"CD",X"93",X"05",X"2B",
		X"10",X"F1",X"C9",X"E6",X"0F",X"DD",X"77",X"00",X"DD",X"19",X"C9",X"FE",X"03",X"D2",X"BD",X"05",
		X"F5",X"21",X"B2",X"60",X"A7",X"CA",X"AB",X"05",X"21",X"B5",X"60",X"FE",X"02",X"C2",X"B3",X"05",
		X"21",X"B8",X"60",X"AF",X"77",X"23",X"77",X"23",X"77",X"F1",X"C3",X"C6",X"05",X"3D",X"F5",X"CD",
		X"9B",X"05",X"F1",X"C8",X"18",X"F7",X"FE",X"03",X"CA",X"E0",X"05",X"11",X"B4",X"60",X"A7",X"CA",
		X"D5",X"05",X"11",X"B7",X"60",X"FE",X"02",X"C2",X"6B",X"05",X"11",X"BA",X"60",X"C3",X"78",X"05",
		X"3D",X"F5",X"CD",X"C6",X"05",X"F1",X"C8",X"18",X"F7",X"21",X"4B",X"36",X"87",X"F5",X"E6",X"7F",
		X"5F",X"16",X"00",X"19",X"5E",X"23",X"56",X"EB",X"5E",X"23",X"56",X"23",X"01",X"E0",X"FF",X"EB",
		X"1A",X"FE",X"3F",X"CA",X"26",X"00",X"77",X"F1",X"30",X"02",X"36",X"10",X"F5",X"13",X"09",X"18",
		X"EF",X"CD",X"28",X"0D",X"0F",X"D0",X"3E",X"05",X"CD",X"E9",X"05",X"21",X"01",X"60",X"11",X"E0",
		X"FF",X"DD",X"21",X"BF",X"74",X"06",X"01",X"C3",X"83",X"05",X"A7",X"CA",X"91",X"06",X"3A",X"8C",
		X"63",X"A7",X"C2",X"A8",X"06",X"3A",X"B8",X"63",X"A7",X"C0",X"3A",X"B0",X"62",X"01",X"0A",X"00",
		X"04",X"91",X"C2",X"40",X"06",X"78",X"07",X"07",X"07",X"07",X"32",X"8C",X"63",X"21",X"44",X"38",
		X"11",X"63",X"74",X"3E",X"08",X"DD",X"21",X"1D",X"00",X"01",X"03",X"00",X"ED",X"B0",X"DD",X"19",
		X"DD",X"E5",X"D1",X"3D",X"C2",X"55",X"06",X"CD",X"32",X"07",X"4F",X"E6",X"0F",X"47",X"79",X"0F",
		X"0F",X"0F",X"0F",X"E6",X"0F",X"C2",X"89",X"06",X"3E",X"05",X"32",X"89",X"60",X"3E",X"70",X"32",
		X"C4",X"74",X"32",X"E4",X"74",X"80",X"47",X"3E",X"10",X"32",X"24",X"75",X"78",X"32",X"04",X"75",
		X"C9",X"3A",X"8C",X"63",X"47",X"E6",X"0F",X"C5",X"CD",X"1C",X"05",X"C1",X"78",X"0F",X"0F",X"0F",
		X"0F",X"E6",X"0F",X"C6",X"0A",X"C3",X"1C",X"05",X"D6",X"01",X"20",X"05",X"21",X"B8",X"63",X"36",
		X"01",X"27",X"32",X"8C",X"63",X"C3",X"6A",X"06",X"4F",X"CF",X"06",X"06",X"11",X"E0",X"FF",X"21",
		X"E2",X"74",X"36",X"10",X"19",X"10",X"FB",X"3A",X"28",X"62",X"91",X"CA",X"D7",X"06",X"47",X"21",
		X"E2",X"74",X"36",X"FF",X"19",X"10",X"FB",X"21",X"03",X"75",X"00",X"00",X"21",X"E3",X"74",X"00",
		X"00",X"3A",X"29",X"62",X"FE",X"64",X"38",X"05",X"3E",X"63",X"32",X"29",X"62",X"01",X"0A",X"FF",
		X"04",X"91",X"D2",X"F0",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C9",X"3A",X"0A",
		X"60",X"EF",X"86",X"09",X"AB",X"09",X"D6",X"09",X"FE",X"09",X"1B",X"0A",X"37",X"0A",X"63",X"0A",
		X"76",X"0A",X"FD",X"26",X"2F",X"26",X"70",X"0C",X"47",X"12",X"7A",X"19",X"7C",X"12",X"F2",X"12",
		X"44",X"13",X"8F",X"13",X"A1",X"13",X"AA",X"13",X"BB",X"13",X"1E",X"14",X"86",X"14",X"15",X"16",
		X"6B",X"19",X"3A",X"29",X"62",X"32",X"84",X"74",X"3A",X"8C",X"63",X"C9",X"21",X"0A",X"60",X"3A",
		X"01",X"60",X"A7",X"C2",X"5C",X"07",X"7E",X"EF",X"79",X"07",X"63",X"07",X"47",X"12",X"77",X"19",
		X"7C",X"12",X"C3",X"07",X"CB",X"07",X"4B",X"08",X"00",X"00",X"00",X"00",X"36",X"00",X"21",X"05",
		X"60",X"34",X"C9",X"E7",X"AF",X"32",X"92",X"63",X"32",X"A0",X"63",X"3E",X"02",X"32",X"27",X"62",
		X"CD",X"D6",X"5F",X"32",X"28",X"62",X"C3",X"92",X"0C",X"21",X"86",X"7D",X"36",X"00",X"23",X"36",
		X"00",X"11",X"1B",X"03",X"CD",X"9F",X"30",X"1C",X"CD",X"9F",X"30",X"CD",X"65",X"09",X"21",X"09",
		X"60",X"36",X"02",X"23",X"34",X"CD",X"74",X"08",X"CD",X"53",X"0A",X"3A",X"0F",X"60",X"FE",X"01",
		X"CC",X"EE",X"09",X"ED",X"5B",X"22",X"60",X"21",X"6C",X"75",X"CD",X"AD",X"07",X"73",X"23",X"23",
		X"72",X"7A",X"D6",X"0A",X"C2",X"BC",X"07",X"77",X"3C",X"32",X"8E",X"75",X"11",X"01",X"02",X"21",
		X"8C",X"76",X"C9",X"CD",X"74",X"08",X"21",X"0A",X"60",X"34",X"C9",X"3A",X"8A",X"63",X"FE",X"00",
		X"C2",X"2D",X"08",X"3E",X"60",X"32",X"8A",X"63",X"0E",X"5F",X"FE",X"00",X"CA",X"3B",X"08",X"21",
		X"86",X"7D",X"36",X"00",X"79",X"CB",X"07",X"30",X"02",X"36",X"01",X"23",X"36",X"00",X"CB",X"07",
		X"30",X"02",X"36",X"01",X"32",X"8B",X"63",X"3E",X"01",X"32",X"80",X"7C",X"C3",X"52",X"0C",X"1A",
		X"77",X"23",X"13",X"10",X"FA",X"C9",X"CD",X"FF",X"07",X"D5",X"11",X"1D",X"00",X"19",X"D1",X"0D",
		X"C2",X"6A",X"0C",X"11",X"1E",X"03",X"CD",X"9F",X"30",X"21",X"FC",X"03",X"11",X"00",X"69",X"06",
		X"14",X"7E",X"12",X"23",X"13",X"10",X"FA",X"C9",X"00",X"00",X"00",X"00",X"00",X"3A",X"8B",X"63",
		X"4F",X"3A",X"8A",X"63",X"3D",X"32",X"8A",X"63",X"C3",X"DA",X"07",X"21",X"09",X"60",X"36",X"02",
		X"23",X"34",X"21",X"8A",X"63",X"36",X"00",X"23",X"36",X"00",X"C9",X"E7",X"CD",X"89",X"0C",X"36",
		X"00",X"C9",X"21",X"00",X"74",X"0E",X"04",X"06",X"00",X"3E",X"10",X"77",X"23",X"10",X"FC",X"0D",
		X"C2",X"57",X"08",X"21",X"00",X"69",X"0E",X"02",X"06",X"C0",X"AF",X"77",X"23",X"10",X"FC",X"0D",
		X"C2",X"68",X"08",X"C9",X"21",X"03",X"74",X"0E",X"20",X"06",X"1D",X"3E",X"10",X"11",X"03",X"00",
		X"77",X"23",X"10",X"FC",X"19",X"0D",X"C2",X"79",X"08",X"21",X"22",X"75",X"11",X"20",X"00",X"0E",
		X"02",X"3E",X"10",X"06",X"0E",X"77",X"19",X"10",X"FC",X"21",X"23",X"75",X"0D",X"C2",X"93",X"08",
		X"21",X"00",X"69",X"06",X"00",X"3E",X"00",X"77",X"23",X"10",X"FC",X"06",X"80",X"77",X"23",X"10",
		X"FC",X"C9",X"3A",X"0A",X"60",X"EF",X"BA",X"08",X"F8",X"08",X"CD",X"74",X"08",X"AF",X"32",X"07",
		X"60",X"11",X"0C",X"03",X"CD",X"9F",X"30",X"21",X"0A",X"60",X"34",X"CD",X"65",X"09",X"AF",X"21",
		X"86",X"7D",X"77",X"2C",X"77",X"06",X"04",X"1E",X"09",X"3A",X"01",X"60",X"FE",X"01",X"CA",X"E4",
		X"08",X"06",X"0C",X"1C",X"3A",X"1A",X"60",X"E6",X"07",X"C2",X"F3",X"08",X"7B",X"CD",X"E9",X"05",
		X"CD",X"16",X"06",X"3A",X"00",X"7D",X"A0",X"C9",X"CD",X"D5",X"08",X"FE",X"04",X"CA",X"06",X"09",
		X"FE",X"08",X"CA",X"19",X"09",X"C9",X"CD",X"77",X"09",X"21",X"48",X"60",X"06",X"08",X"AF",X"77",
		X"2C",X"10",X"FC",X"21",X"00",X"00",X"C3",X"38",X"09",X"CD",X"77",X"09",X"CD",X"77",X"09",X"11",
		X"48",X"60",X"3A",X"20",X"60",X"12",X"1C",X"21",X"5E",X"09",X"01",X"07",X"00",X"ED",X"B0",X"11",
		X"01",X"01",X"CD",X"9F",X"30",X"21",X"00",X"01",X"22",X"0E",X"60",X"CD",X"74",X"08",X"11",X"40",
		X"60",X"3A",X"20",X"60",X"12",X"1C",X"21",X"5E",X"09",X"01",X"07",X"00",X"ED",X"B0",X"11",X"00",
		X"01",X"CD",X"9F",X"30",X"AF",X"32",X"0A",X"60",X"3E",X"03",X"32",X"05",X"60",X"C9",X"01",X"65",
		X"3A",X"01",X"00",X"00",X"00",X"11",X"00",X"04",X"CD",X"9F",X"30",X"11",X"14",X"03",X"06",X"06",
		X"CD",X"9F",X"30",X"1C",X"10",X"FA",X"C9",X"21",X"01",X"60",X"3E",X"99",X"86",X"27",X"77",X"11",
		X"00",X"04",X"CD",X"9F",X"30",X"C9",X"CD",X"52",X"08",X"CD",X"1C",X"01",X"11",X"82",X"7D",X"3E",
		X"01",X"12",X"21",X"0A",X"60",X"3A",X"0E",X"60",X"A7",X"C2",X"9F",X"09",X"36",X"01",X"C9",X"3A",
		X"26",X"60",X"3D",X"CA",X"A8",X"09",X"AF",X"12",X"36",X"03",X"C9",X"21",X"40",X"60",X"11",X"28",
		X"62",X"01",X"08",X"00",X"ED",X"B0",X"2A",X"2A",X"62",X"7E",X"32",X"27",X"62",X"3A",X"0F",X"60",
		X"A7",X"21",X"09",X"60",X"11",X"0A",X"60",X"CA",X"D0",X"09",X"36",X"78",X"EB",X"36",X"02",X"C9",
		X"36",X"01",X"EB",X"36",X"05",X"C9",X"AF",X"32",X"86",X"7D",X"32",X"87",X"7D",X"11",X"02",X"03",
		X"CD",X"9F",X"30",X"11",X"01",X"02",X"CD",X"9F",X"30",X"3E",X"05",X"32",X"0A",X"60",X"3E",X"02",
		X"32",X"E0",X"74",X"3E",X"25",X"32",X"C0",X"74",X"3E",X"20",X"32",X"A0",X"74",X"C9",X"21",X"48",
		X"60",X"11",X"28",X"62",X"01",X"08",X"00",X"ED",X"B0",X"2A",X"2A",X"62",X"7E",X"32",X"27",X"62",
		X"3E",X"78",X"32",X"09",X"60",X"3E",X"04",X"32",X"0A",X"60",X"C9",X"AF",X"32",X"86",X"7D",X"32",
		X"87",X"7D",X"11",X"03",X"03",X"CD",X"9F",X"30",X"11",X"01",X"02",X"CD",X"9F",X"30",X"CD",X"EE",
		X"09",X"3E",X"05",X"32",X"0A",X"60",X"C9",X"11",X"04",X"03",X"CD",X"9F",X"30",X"11",X"02",X"02",
		X"CD",X"9F",X"30",X"11",X"00",X"02",X"CD",X"9F",X"30",X"11",X"00",X"06",X"CD",X"9F",X"30",X"21",
		X"0A",X"60",X"34",X"3E",X"01",X"32",X"40",X"77",X"3E",X"25",X"32",X"20",X"77",X"3E",X"20",X"32",
		X"00",X"77",X"C9",X"DF",X"CD",X"74",X"08",X"21",X"09",X"60",X"36",X"01",X"2C",X"34",X"11",X"2C",
		X"62",X"1A",X"A7",X"C3",X"01",X"19",X"3A",X"85",X"63",X"EF",X"10",X"04",X"8A",X"0A",X"69",X"30",
		X"96",X"04",X"D5",X"04",X"31",X"0B",X"69",X"30",X"06",X"05",X"21",X"AF",X"62",X"34",X"CB",X"46",
		X"C0",X"E5",X"21",X"03",X"69",X"11",X"04",X"00",X"01",X"FF",X"0E",X"CD",X"3D",X"00",X"E1",X"7E",
		X"E6",X"0F",X"F5",X"CC",X"4A",X"30",X"3A",X"0B",X"69",X"FE",X"70",X"30",X"07",X"AF",X"32",X"0C",
		X"6A",X"32",X"10",X"6A",X"F1",X"E6",X"07",X"FE",X"06",X"20",X"2D",X"3A",X"15",X"6A",X"EE",X"0F",
		X"32",X"15",X"6A",X"CB",X"47",X"3E",X"C6",X"28",X"02",X"3E",X"10",X"32",X"88",X"75",X"32",X"68",
		X"76",X"3A",X"19",X"6A",X"EE",X"0F",X"32",X"19",X"6A",X"DD",X"21",X"1C",X"6A",X"DD",X"7E",X"01",
		X"EE",X"80",X"DD",X"77",X"01",X"DD",X"77",X"05",X"3A",X"0B",X"69",X"FE",X"40",X"D0",X"AF",X"32",
		X"0C",X"6A",X"32",X"10",X"6A",X"32",X"AF",X"62",X"3E",X"19",X"32",X"15",X"6A",X"32",X"19",X"6A",
		X"21",X"63",X"76",X"CD",X"26",X"18",X"3E",X"10",X"32",X"88",X"75",X"32",X"68",X"76",X"AF",X"32",
		X"1C",X"6A",X"32",X"20",X"6A",X"32",X"30",X"69",X"32",X"34",X"69",X"21",X"70",X"77",X"11",X"8A",
		X"0B",X"CD",X"65",X"0B",X"21",X"BB",X"0B",X"06",X"04",X"CD",X"42",X"0B",X"3E",X"20",X"C3",X"8B",
		X"04",X"3E",X"40",X"C3",X"8B",X"04",X"32",X"87",X"7D",X"21",X"8A",X"60",X"36",X"08",X"23",X"36",
		X"03",X"C9",X"DD",X"21",X"4C",X"69",X"11",X"08",X"00",X"7E",X"DD",X"77",X"00",X"23",X"7E",X"DD",
		X"77",X"01",X"23",X"7E",X"DD",X"77",X"02",X"23",X"7E",X"DD",X"77",X"03",X"23",X"DD",X"19",X"11",
		X"04",X"00",X"10",X"E5",X"C9",X"01",X"E0",X"FF",X"22",X"B9",X"63",X"1A",X"13",X"3C",X"28",X"0C",
		X"3C",X"28",X"0F",X"3D",X"3D",X"FE",X"AA",X"C8",X"77",X"09",X"18",X"EF",X"2A",X"B9",X"63",X"23",
		X"18",X"E6",X"C5",X"01",X"20",X"00",X"09",X"C1",X"18",X"E1",X"17",X"15",X"24",X"10",X"10",X"10",
		X"10",X"1B",X"15",X"29",X"10",X"16",X"22",X"1F",X"1D",X"10",X"10",X"10",X"10",X"1D",X"11",X"22",
		X"19",X"1F",X"2B",X"FF",X"FF",X"10",X"10",X"10",X"10",X"10",X"23",X"11",X"26",X"15",X"10",X"29",
		X"1F",X"25",X"22",X"10",X"20",X"11",X"20",X"11",X"10",X"38",X"AA",X"78",X"69",X"07",X"C8",X"88",
		X"05",X"07",X"C8",X"48",X"5F",X"0D",X"80",X"A8",X"16",X"00",X"80",X"7F",X"2D",X"08",X"CE",X"7F",
		X"2D",X"88",X"E0",X"32",X"03",X"7D",X"32",X"83",X"60",X"C9",X"32",X"80",X"60",X"3A",X"15",X"62",
		X"A7",X"3E",X"01",X"28",X"01",X"AF",X"32",X"07",X"7D",X"C9",X"F5",X"32",X"07",X"62",X"E6",X"7F",
		X"FE",X"08",X"CC",X"8F",X"1D",X"F1",X"C9",X"32",X"15",X"62",X"CD",X"8F",X"1D",X"C9",X"3E",X"03",
		X"32",X"82",X"60",X"AF",X"32",X"8C",X"60",X"7E",X"E6",X"80",X"C9",X"00",X"00",X"3E",X"29",X"32",
		X"8F",X"60",X"3E",X"20",X"32",X"09",X"60",X"21",X"4C",X"69",X"36",X"00",X"21",X"54",X"69",X"36",
		X"00",X"E1",X"C9",X"AF",X"32",X"8C",X"60",X"3E",X"01",X"32",X"82",X"60",X"C3",X"AC",X"50",X"32",
		X"80",X"7D",X"3A",X"8C",X"60",X"32",X"81",X"7D",X"C9",X"CD",X"1C",X"01",X"06",X"28",X"21",X"58",
		X"69",X"36",X"00",X"23",X"10",X"FB",X"C9",X"00",X"D2",X"E6",X"16",X"AF",X"32",X"89",X"60",X"C3",
		X"EE",X"16",X"21",X"8A",X"74",X"11",X"0A",X"3D",X"0E",X"14",X"06",X"06",X"CD",X"FF",X"07",X"D5",
		X"11",X"1A",X"00",X"19",X"D1",X"0D",X"20",X"F2",X"0E",X"05",X"06",X"03",X"C3",X"06",X"08",X"00",
		X"3A",X"85",X"63",X"EF",X"78",X"0C",X"91",X"0C",X"DF",X"21",X"09",X"60",X"36",X"20",X"21",X"85",
		X"63",X"34",X"CD",X"1C",X"01",X"CD",X"74",X"08",X"C9",X"AF",X"32",X"80",X"7C",X"21",X"0A",X"60",
		X"C9",X"DF",X"CD",X"74",X"08",X"AF",X"32",X"8C",X"63",X"11",X"01",X"05",X"CD",X"9F",X"30",X"21",
		X"86",X"7D",X"36",X"00",X"23",X"36",X"01",X"3A",X"27",X"62",X"3D",X"CA",X"D4",X"0C",X"3D",X"CA",
		X"DF",X"0C",X"3D",X"CA",X"F2",X"0C",X"00",X"00",X"00",X"21",X"86",X"7D",X"36",X"01",X"3E",X"03",
		X"32",X"89",X"60",X"11",X"40",X"3C",X"CD",X"A7",X"0D",X"3A",X"27",X"62",X"FE",X"03",X"00",X"00",
		X"00",X"C3",X"A0",X"3F",X"11",X"86",X"3B",X"3E",X"02",X"32",X"89",X"60",X"C3",X"E7",X"0C",X"11",
		X"C6",X"3A",X"3E",X"01",X"32",X"89",X"60",X"21",X"86",X"7D",X"36",X"01",X"23",X"36",X"00",X"C3",
		X"C6",X"0C",X"00",X"00",X"00",X"3E",X"04",X"32",X"89",X"60",X"11",X"BE",X"3F",X"C3",X"C6",X"0C",
		X"31",X"44",X"57",X"10",X"7A",X"92",X"99",X"A7",X"30",X"43",X"56",X"10",X"79",X"91",X"98",X"A6",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CD",X"89",X"0C",X"3A",X"07",X"60",X"C9",X"00",
		X"DD",X"77",X"07",X"3A",X"27",X"62",X"FE",X"02",X"3E",X"02",X"C0",X"3E",X"04",X"C9",X"00",X"00",
		X"00",X"00",X"00",X"21",X"87",X"76",X"CD",X"4C",X"0D",X"21",X"47",X"75",X"06",X"04",X"36",X"FD",
		X"23",X"10",X"FB",X"11",X"1C",X"00",X"19",X"06",X"04",X"36",X"FC",X"23",X"10",X"FB",X"C9",X"CD",
		X"56",X"0F",X"CD",X"41",X"24",X"21",X"09",X"60",X"36",X"40",X"23",X"34",X"21",X"5C",X"38",X"CD",
		X"C0",X"57",X"11",X"00",X"69",X"01",X"08",X"00",X"ED",X"B0",X"3A",X"27",X"62",X"FE",X"03",X"28",
		X"0A",X"0F",X"0F",X"D8",X"21",X"0B",X"69",X"0E",X"00",X"FF",X"C9",X"21",X"08",X"69",X"0E",X"54",
		X"FF",X"11",X"04",X"00",X"01",X"54",X"02",X"21",X"00",X"69",X"CD",X"3D",X"00",X"01",X"F8",X"0C",
		X"21",X"03",X"69",X"CD",X"3D",X"00",X"C9",X"1A",X"32",X"B3",X"63",X"CD",X"15",X"0F",X"13",X"1A",
		X"67",X"44",X"13",X"1A",X"6F",X"4D",X"D5",X"CD",X"F0",X"2F",X"D1",X"22",X"AB",X"63",X"78",X"E6",
		X"07",X"32",X"B4",X"63",X"79",X"E6",X"07",X"32",X"AF",X"63",X"13",X"1A",X"67",X"90",X"D2",X"D3",
		X"0D",X"ED",X"44",X"32",X"B1",X"63",X"13",X"1A",X"6F",X"91",X"32",X"B2",X"63",X"1A",X"E6",X"07",
		X"32",X"B0",X"63",X"D5",X"CD",X"F0",X"2F",X"D1",X"22",X"AD",X"63",X"3A",X"B3",X"63",X"FE",X"05",
		X"D2",X"46",X"0E",X"3A",X"B2",X"63",X"D6",X"08",X"47",X"3A",X"AF",X"63",X"80",X"32",X"B2",X"63",
		X"2A",X"AB",X"63",X"3A",X"B3",X"63",X"3D",X"28",X"19",X"3D",X"28",X"12",X"3D",X"28",X"0B",X"3D",
		X"28",X"04",X"3E",X"C2",X"18",X"0E",X"3E",X"B7",X"18",X"0A",X"3E",X"C0",X"18",X"06",X"3E",X"C4",
		X"18",X"02",X"3E",X"C6",X"77",X"32",X"B5",X"63",X"3A",X"B2",X"63",X"D6",X"08",X"32",X"B2",X"63",
		X"38",X"07",X"2C",X"3A",X"B5",X"63",X"77",X"18",X"EF",X"C3",X"0A",X"0F",X"00",X"00",X"30",X"01",
		X"3C",X"77",X"13",X"C3",X"A7",X"0D",X"FE",X"08",X"D2",X"91",X"0E",X"D6",X"05",X"28",X"07",X"3D",
		X"28",X"08",X"3E",X"F2",X"18",X"06",X"3E",X"E1",X"18",X"02",X"3E",X"E4",X"2A",X"AB",X"63",X"77",
		X"3C",X"32",X"B5",X"63",X"01",X"20",X"00",X"09",X"3A",X"B1",X"63",X"D6",X"10",X"38",X"12",X"32",
		X"B1",X"63",X"3A",X"B5",X"63",X"77",X"01",X"20",X"00",X"09",X"3A",X"B1",X"63",X"D6",X"08",X"18",
		X"EC",X"3A",X"B3",X"63",X"FE",X"08",X"3A",X"B5",X"63",X"30",X"02",X"3C",X"77",X"13",X"C3",X"A7",
		X"0D",X"FE",X"0C",X"D2",X"C1",X"0E",X"D6",X"08",X"28",X"0A",X"3D",X"28",X"0B",X"3D",X"28",X"0C",
		X"3E",X"AF",X"18",X"0A",X"3E",X"F1",X"18",X"06",X"3E",X"E0",X"18",X"02",X"3E",X"B5",X"32",X"B5",
		X"63",X"2A",X"AB",X"63",X"77",X"01",X"20",X"00",X"09",X"3A",X"B1",X"63",X"D6",X"08",X"C3",X"6D",
		X"0E",X"FE",X"0C",X"20",X"2A",X"3E",X"D0",X"2A",X"AB",X"63",X"77",X"32",X"B5",X"63",X"01",X"20",
		X"00",X"09",X"3A",X"B1",X"63",X"D6",X"08",X"32",X"B1",X"63",X"38",X"0B",X"3A",X"B5",X"63",X"3C",
		X"FE",X"D8",X"CA",X"8D",X"0E",X"18",X"E3",X"2A",X"AB",X"63",X"2C",X"3E",X"D4",X"18",X"DB",X"FE",
		X"0D",X"28",X"0F",X"FE",X"0E",X"28",X"03",X"C3",X"43",X"0F",X"3E",X"CA",X"2A",X"AB",X"63",X"C3",
		X"24",X"0E",X"3E",X"AE",X"2A",X"AB",X"63",X"C3",X"24",X"0E",X"3A",X"B3",X"63",X"FE",X"03",X"3A",
		X"B5",X"63",X"C3",X"3E",X"0E",X"FE",X"AA",X"C0",X"3A",X"27",X"62",X"FE",X"04",X"28",X"0B",X"FE",
		X"02",X"28",X"16",X"CD",X"BC",X"59",X"00",X"33",X"33",X"C9",X"0E",X"F7",X"06",X"0D",X"13",X"1A",
		X"6F",X"13",X"1A",X"67",X"71",X"10",X"F7",X"18",X"EE",X"0E",X"C3",X"18",X"EF",X"0E",X"F0",X"06",
		X"04",X"18",X"EB",X"FE",X"0F",X"28",X"0A",X"FE",X"10",X"3E",X"E7",X"CA",X"AE",X"0E",X"C3",X"A7",
		X"0D",X"3E",X"F8",X"18",X"F6",X"0F",X"06",X"27",X"21",X"00",X"62",X"AF",X"77",X"2C",X"10",X"FC",
		X"0E",X"11",X"16",X"80",X"21",X"80",X"62",X"42",X"77",X"23",X"10",X"FC",X"0D",X"20",X"F8",X"21",
		X"9C",X"3D",X"11",X"80",X"62",X"01",X"40",X"00",X"ED",X"B0",X"3A",X"29",X"62",X"47",X"A7",X"17",
		X"A7",X"17",X"A7",X"17",X"80",X"80",X"C6",X"28",X"FE",X"51",X"38",X"02",X"3E",X"50",X"21",X"B0",
		X"62",X"06",X"03",X"77",X"2C",X"10",X"FC",X"87",X"47",X"3E",X"DC",X"90",X"FE",X"28",X"30",X"02",
		X"3E",X"28",X"77",X"2C",X"77",X"21",X"09",X"62",X"36",X"04",X"2C",X"36",X"08",X"3A",X"27",X"62",
		X"4F",X"21",X"34",X"6A",X"36",X"00",X"2C",X"36",X"96",X"2C",X"36",X"00",X"2C",X"36",X"40",X"C3",
		X"CB",X"0F",X"32",X"25",X"62",X"21",X"8D",X"60",X"36",X"03",X"C9",X"79",X"EF",X"00",X"00",X"D7",
		X"0F",X"1F",X"10",X"87",X"10",X"4F",X"11",X"CD",X"89",X"48",X"CD",X"E9",X"48",X"CD",X"55",X"48",
		X"00",X"00",X"CD",X"50",X"4D",X"11",X"07",X"64",X"0E",X"1C",X"06",X"05",X"CD",X"2A",X"12",X"00",
		X"00",X"00",X"00",X"00",X"00",X"18",X"09",X"00",X"32",X"AF",X"62",X"AF",X"32",X"8C",X"60",X"C9",
		X"21",X"0C",X"3E",X"CD",X"A6",X"11",X"21",X"1B",X"10",X"11",X"07",X"67",X"01",X"1C",X"08",X"CD",
		X"2A",X"12",X"11",X"07",X"68",X"06",X"02",X"C3",X"3E",X"55",X"C9",X"00",X"00",X"02",X"02",X"21",
		X"EC",X"3D",X"11",X"07",X"64",X"01",X"1C",X"05",X"CD",X"2A",X"12",X"CD",X"86",X"11",X"21",X"18",
		X"3E",X"11",X"A7",X"65",X"01",X"0C",X"06",X"CD",X"2A",X"12",X"DD",X"21",X"A0",X"65",X"21",X"B8",
		X"69",X"11",X"10",X"00",X"06",X"06",X"CD",X"D3",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"21",
		X"04",X"3E",X"11",X"FC",X"69",X"01",X"04",X"00",X"ED",X"B0",X"21",X"1C",X"3E",X"11",X"44",X"69",
		X"01",X"08",X"00",X"ED",X"B0",X"21",X"7C",X"10",X"CD",X"A6",X"11",X"21",X"3C",X"3E",X"11",X"0C",
		X"6A",X"01",X"14",X"00",X"ED",X"B0",X"3E",X"01",X"C3",X"FB",X"53",X"C9",X"2B",X"63",X"6B",X"63",
		X"8B",X"A3",X"A3",X"6B",X"9B",X"18",X"C9",X"21",X"EC",X"3D",X"11",X"07",X"64",X"01",X"1C",X"05",
		X"CD",X"2A",X"12",X"CD",X"86",X"11",X"21",X"00",X"66",X"11",X"10",X"00",X"3E",X"01",X"06",X"06",
		X"77",X"19",X"10",X"FC",X"21",X"35",X"5E",X"11",X"A3",X"65",X"01",X"0E",X"06",X"CD",X"EC",X"11",
		X"21",X"41",X"5E",X"11",X"A7",X"65",X"01",X"0C",X"06",X"CD",X"2A",X"12",X"DD",X"21",X"A0",X"65",
		X"21",X"B8",X"69",X"06",X"06",X"11",X"10",X"00",X"CD",X"D3",X"11",X"21",X"A0",X"65",X"06",X"06",
		X"36",X"01",X"19",X"10",X"FB",X"21",X"2B",X"5E",X"CD",X"A6",X"11",X"21",X"23",X"5E",X"11",X"0C",
		X"6A",X"01",X"08",X"00",X"ED",X"B0",X"00",X"00",X"00",X"DD",X"21",X"00",X"64",X"DD",X"36",X"00",
		X"01",X"DD",X"36",X"16",X"4B",X"DD",X"36",X"0E",X"A0",X"DD",X"36",X"05",X"38",X"DD",X"36",X"0F",
		X"40",X"DD",X"36",X"20",X"01",X"DD",X"36",X"36",X"4B",X"DD",X"36",X"2E",X"D8",X"DD",X"36",X"25",
		X"60",X"DD",X"36",X"2F",X"40",X"C9",X"11",X"F7",X"39",X"E5",X"21",X"8A",X"60",X"36",X"0E",X"23",
		X"36",X"03",X"E1",X"C9",X"3A",X"27",X"62",X"FE",X"03",X"C8",X"21",X"8A",X"60",X"36",X"07",X"23",
		X"36",X"03",X"C9",X"11",X"20",X"00",X"3A",X"29",X"62",X"FE",X"03",X"06",X"08",X"D8",X"C3",X"CA",
		X"5F",X"16",X"00",X"3A",X"29",X"62",X"FE",X"03",X"3E",X"08",X"D8",X"C3",X"D0",X"5F",X"00",X"CD",
		X"10",X"4F",X"CD",X"D0",X"51",X"CD",X"54",X"52",X"21",X"5C",X"3E",X"11",X"0C",X"6A",X"01",X"0C",
		X"00",X"ED",X"B0",X"CD",X"A6",X"11",X"DD",X"21",X"A0",X"64",X"DD",X"36",X"00",X"01",X"DD",X"36",
		X"20",X"01",X"21",X"50",X"69",X"06",X"02",X"11",X"20",X"00",X"CD",X"D3",X"11",X"C9",X"3F",X"0C",
		X"08",X"08",X"73",X"50",X"8D",X"50",X"CD",X"48",X"3A",X"11",X"07",X"65",X"01",X"0C",X"0A",X"CD",
		X"2A",X"12",X"DD",X"21",X"00",X"65",X"21",X"58",X"69",X"06",X"0A",X"11",X"10",X"00",X"CD",X"D3",
		X"11",X"C9",X"3B",X"0F",X"04",X"01",X"11",X"83",X"66",X"01",X"0E",X"05",X"CD",X"EC",X"11",X"21",
		X"08",X"3E",X"11",X"87",X"66",X"01",X"0C",X"02",X"C9",X"79",X"FE",X"15",X"30",X"05",X"81",X"81",
		X"C3",X"24",X"05",X"21",X"A0",X"59",X"FE",X"15",X"CA",X"2B",X"05",X"23",X"23",X"23",X"C3",X"2B",
		X"05",X"00",X"00",X"DD",X"7E",X"03",X"77",X"2C",X"DD",X"7E",X"07",X"77",X"2C",X"DD",X"7E",X"08",
		X"77",X"2C",X"DD",X"7E",X"05",X"77",X"2C",X"DD",X"19",X"10",X"E8",X"C9",X"7E",X"12",X"23",X"1C",
		X"1C",X"7E",X"12",X"23",X"7B",X"81",X"5F",X"10",X"F3",X"C9",X"3A",X"05",X"62",X"FE",X"48",X"C2",
		X"A6",X"1D",X"3A",X"03",X"62",X"FE",X"A0",X"D2",X"A6",X"1D",X"3E",X"A0",X"32",X"03",X"62",X"C3",
		X"A6",X"1D",X"3A",X"00",X"7D",X"E6",X"01",X"C2",X"00",X"80",X"31",X"00",X"6C",X"C3",X"B5",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E5",X"C5",X"06",X"04",X"7E",X"12",
		X"23",X"1C",X"10",X"FA",X"C1",X"E1",X"7B",X"81",X"5F",X"10",X"EF",X"C9",X"3A",X"27",X"62",X"FE",
		X"04",X"36",X"0A",X"C0",X"36",X"08",X"C9",X"DF",X"CD",X"31",X"4F",X"DD",X"21",X"00",X"62",X"21",
		X"4C",X"69",X"DD",X"36",X"00",X"01",X"DD",X"71",X"03",X"71",X"2C",X"DD",X"36",X"07",X"05",X"36",
		X"05",X"2C",X"DD",X"36",X"08",X"07",X"36",X"07",X"2C",X"DD",X"70",X"05",X"70",X"DD",X"36",X"0F",
		X"01",X"CD",X"95",X"40",X"34",X"11",X"01",X"06",X"CD",X"9F",X"30",X"C9",X"CD",X"BD",X"1D",X"3A",
		X"9D",X"63",X"EF",X"8B",X"12",X"AC",X"12",X"DE",X"12",X"00",X"00",X"DF",X"21",X"4D",X"69",X"CD",
		X"7C",X"47",X"21",X"9D",X"63",X"34",X"7A",X"32",X"9E",X"63",X"3E",X"08",X"32",X"09",X"60",X"AF",
		X"32",X"8C",X"60",X"32",X"89",X"60",X"3E",X"03",X"32",X"88",X"60",X"C9",X"DF",X"3E",X"08",X"32",
		X"09",X"60",X"21",X"9E",X"63",X"35",X"CA",X"CB",X"12",X"21",X"4D",X"69",X"3E",X"18",X"AE",X"77",
		X"21",X"55",X"69",X"3E",X"18",X"AE",X"77",X"00",X"00",X"00",X"C9",X"21",X"4D",X"69",X"00",X"00",
		X"00",X"00",X"00",X"00",X"21",X"9D",X"63",X"34",X"3E",X"56",X"32",X"09",X"60",X"C9",X"DF",X"CD",
		X"92",X"4E",X"21",X"0A",X"60",X"3A",X"0E",X"60",X"A7",X"CA",X"ED",X"12",X"34",X"34",X"2B",X"36",
		X"01",X"C9",X"CD",X"8E",X"59",X"AF",X"32",X"2C",X"62",X"21",X"28",X"62",X"35",X"7E",X"11",X"40",
		X"60",X"01",X"08",X"00",X"ED",X"B0",X"A7",X"C2",X"34",X"13",X"3E",X"01",X"21",X"B2",X"60",X"CD",
		X"CA",X"13",X"21",X"D4",X"76",X"3A",X"0F",X"60",X"A7",X"28",X"07",X"11",X"02",X"03",X"CD",X"9F",
		X"30",X"2B",X"CD",X"26",X"18",X"11",X"00",X"03",X"CD",X"9F",X"30",X"21",X"09",X"60",X"36",X"C0",
		X"23",X"36",X"10",X"C9",X"0E",X"0A",X"3A",X"0F",X"60",X"A7",X"CA",X"3F",X"13",X"0E",X"17",X"79",
		X"32",X"0A",X"60",X"C9",X"CD",X"1C",X"01",X"AF",X"32",X"2C",X"62",X"21",X"28",X"62",X"35",X"7E",
		X"11",X"48",X"60",X"01",X"08",X"00",X"ED",X"B0",X"A7",X"C2",X"7F",X"13",X"3E",X"03",X"21",X"B5",
		X"60",X"CD",X"CA",X"13",X"11",X"03",X"03",X"CD",X"9F",X"30",X"11",X"00",X"03",X"CD",X"9F",X"30",
		X"21",X"D3",X"76",X"CD",X"26",X"18",X"21",X"09",X"60",X"36",X"C0",X"23",X"36",X"11",X"C9",X"0E",
		X"17",X"3A",X"40",X"60",X"A7",X"C2",X"8A",X"13",X"0E",X"0A",X"79",X"32",X"0A",X"60",X"C9",X"DF",
		X"0E",X"17",X"3A",X"48",X"60",X"34",X"A7",X"C2",X"9C",X"13",X"0E",X"14",X"79",X"32",X"0A",X"60",
		X"C9",X"DF",X"0E",X"17",X"3A",X"40",X"60",X"C3",X"95",X"13",X"3A",X"26",X"60",X"32",X"82",X"7D",
		X"AF",X"32",X"0A",X"60",X"21",X"01",X"01",X"22",X"0D",X"60",X"C9",X"AF",X"32",X"0D",X"60",X"32",
		X"0E",X"60",X"32",X"0A",X"60",X"3C",X"32",X"82",X"7D",X"C9",X"11",X"C6",X"61",X"12",X"CF",X"13",
		X"01",X"03",X"00",X"ED",X"B0",X"06",X"03",X"21",X"B1",X"61",X"1B",X"1A",X"0F",X"0F",X"0F",X"0F",
		X"E6",X"0F",X"77",X"23",X"1A",X"E6",X"0F",X"77",X"23",X"10",X"EF",X"06",X"0E",X"36",X"10",X"23",
		X"10",X"FB",X"36",X"3F",X"06",X"05",X"21",X"A5",X"61",X"11",X"C7",X"61",X"1A",X"96",X"23",X"13",
		X"1A",X"9E",X"23",X"13",X"1A",X"9E",X"D8",X"C5",X"06",X"19",X"4E",X"1A",X"77",X"79",X"12",X"2B",
		X"1B",X"10",X"F7",X"01",X"F5",X"FF",X"09",X"EB",X"09",X"EB",X"C1",X"10",X"DF",X"C9",X"CD",X"16",
		X"06",X"DF",X"CD",X"74",X"08",X"3E",X"00",X"32",X"0E",X"60",X"32",X"0D",X"60",X"21",X"1C",X"61",
		X"11",X"22",X"00",X"06",X"05",X"3E",X"01",X"BE",X"CA",X"59",X"14",X"19",X"10",X"F9",X"21",X"1C",
		X"61",X"06",X"05",X"3E",X"03",X"BE",X"CA",X"4F",X"14",X"19",X"10",X"F9",X"C3",X"75",X"14",X"3E",
		X"01",X"32",X"0E",X"60",X"32",X"0D",X"60",X"3E",X"00",X"21",X"26",X"60",X"B6",X"32",X"82",X"7D",
		X"3E",X"00",X"32",X"09",X"60",X"21",X"0A",X"60",X"34",X"11",X"0D",X"03",X"06",X"0C",X"CD",X"9F",
		X"30",X"13",X"10",X"FA",X"C9",X"3E",X"01",X"32",X"82",X"7D",X"32",X"05",X"60",X"32",X"07",X"60",
		X"3E",X"00",X"32",X"0A",X"60",X"C9",X"CD",X"16",X"06",X"21",X"09",X"60",X"7E",X"A7",X"C2",X"DC",
		X"14",X"32",X"86",X"7D",X"32",X"87",X"7D",X"36",X"01",X"21",X"30",X"60",X"36",X"0A",X"23",X"36",
		X"00",X"23",X"36",X"03",X"23",X"36",X"3C",X"23",X"36",X"3E",X"23",X"36",X"00",X"21",X"E8",X"75",
		X"22",X"36",X"60",X"21",X"1C",X"61",X"3A",X"0E",X"60",X"07",X"3C",X"4F",X"11",X"22",X"00",X"06",
		X"04",X"7E",X"B9",X"CA",X"C9",X"14",X"19",X"10",X"F8",X"22",X"38",X"60",X"11",X"F3",X"FF",X"19",
		X"22",X"3A",X"60",X"06",X"00",X"3A",X"35",X"60",X"4F",X"CD",X"FA",X"15",X"21",X"34",X"60",X"35",
		X"C2",X"FC",X"14",X"36",X"3E",X"2B",X"35",X"CA",X"C6",X"15",X"7E",X"06",X"FF",X"04",X"D6",X"0A",
		X"D2",X"ED",X"14",X"C6",X"0A",X"32",X"52",X"75",X"78",X"32",X"72",X"75",X"21",X"30",X"60",X"46",
		X"36",X"0A",X"3A",X"10",X"60",X"CB",X"7F",X"C2",X"46",X"15",X"E6",X"03",X"C2",X"14",X"15",X"3C",
		X"77",X"C3",X"8A",X"15",X"05",X"CA",X"1D",X"15",X"78",X"77",X"C3",X"8A",X"15",X"CB",X"4F",X"C2",
		X"39",X"15",X"3A",X"35",X"60",X"3C",X"FE",X"1E",X"C2",X"2D",X"15",X"3E",X"00",X"32",X"35",X"60",
		X"4F",X"06",X"00",X"CD",X"FA",X"15",X"C3",X"8A",X"15",X"3A",X"35",X"60",X"D6",X"01",X"F2",X"2D",
		X"15",X"3E",X"1D",X"C3",X"2D",X"15",X"3A",X"35",X"60",X"FE",X"1C",X"CA",X"6D",X"15",X"FE",X"1D",
		X"CA",X"C6",X"15",X"2A",X"36",X"60",X"01",X"68",X"74",X"A7",X"ED",X"42",X"CA",X"8A",X"15",X"09",
		X"C6",X"11",X"77",X"01",X"E0",X"FF",X"09",X"22",X"36",X"60",X"C3",X"8A",X"15",X"2A",X"36",X"60",
		X"01",X"20",X"00",X"09",X"A7",X"01",X"08",X"76",X"ED",X"42",X"C2",X"86",X"15",X"21",X"E8",X"75",
		X"3E",X"10",X"77",X"C3",X"67",X"15",X"09",X"C3",X"80",X"15",X"21",X"32",X"60",X"35",X"C2",X"F9",
		X"15",X"3A",X"31",X"60",X"A7",X"C2",X"B8",X"15",X"3E",X"01",X"32",X"31",X"60",X"11",X"BF",X"01",
		X"FD",X"2A",X"38",X"60",X"FD",X"6E",X"04",X"FD",X"66",X"05",X"E5",X"DD",X"E1",X"CD",X"7C",X"05",
		X"3E",X"10",X"32",X"32",X"60",X"C3",X"F9",X"15",X"AF",X"32",X"31",X"60",X"ED",X"5B",X"38",X"60",
		X"13",X"13",X"13",X"C3",X"A0",X"15",X"ED",X"5B",X"38",X"60",X"AF",X"12",X"21",X"09",X"60",X"36",
		X"80",X"23",X"35",X"06",X"0C",X"21",X"E8",X"75",X"FD",X"2A",X"3A",X"60",X"11",X"E0",X"FF",X"7E",
		X"FD",X"77",X"00",X"FD",X"23",X"19",X"10",X"F7",X"06",X"05",X"11",X"14",X"03",X"CD",X"9F",X"30",
		X"13",X"10",X"FA",X"11",X"1A",X"03",X"CD",X"9F",X"30",X"C9",X"D5",X"E5",X"CB",X"21",X"21",X"0F",
		X"36",X"09",X"EB",X"21",X"74",X"69",X"1A",X"13",X"77",X"23",X"36",X"60",X"23",X"36",X"04",X"23",
		X"1A",X"77",X"E1",X"D1",X"C9",X"3A",X"27",X"62",X"FE",X"03",X"CA",X"41",X"16",X"CD",X"BD",X"30",
		X"21",X"58",X"69",X"06",X"14",X"36",X"00",X"23",X"10",X"FB",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"3A",X"88",X"63",X"EF",X"A3",X"16",X"BB",X"16",X"57",X"17",X"8E",X"17",X"8E",
		X"17",X"CD",X"BD",X"1D",X"3A",X"88",X"63",X"EF",X"B6",X"17",X"69",X"30",X"39",X"18",X"6F",X"18",
		X"80",X"18",X"C6",X"18",X"45",X"5E",X"00",X"3A",X"27",X"62",X"FE",X"04",X"C2",X"2F",X"20",X"7D",
		X"FE",X"60",X"D2",X"2F",X"20",X"C3",X"BA",X"21",X"DA",X"B4",X"2A",X"3A",X"03",X"62",X"67",X"3A",
		X"05",X"62",X"C6",X"04",X"6F",X"CD",X"F0",X"2F",X"7E",X"FE",X"D0",X"D2",X"B4",X"2A",X"AF",X"32",
		X"8C",X"6A",X"C3",X"AC",X"2A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"CD",X"08",X"17",X"3A",X"08",X"69",X"C6",X"14",X"32",X"34",X"6A",X"00",X"3E",
		X"FF",X"21",X"08",X"69",X"4F",X"FF",X"21",X"88",X"63",X"34",X"C9",X"AF",X"CD",X"0F",X"58",X"3A",
		X"A3",X"63",X"4F",X"3A",X"34",X"6A",X"FE",X"08",X"DA",X"E1",X"16",X"CB",X"79",X"CA",X"D5",X"16",
		X"3E",X"01",X"32",X"A0",X"62",X"CD",X"02",X"26",X"3A",X"A3",X"63",X"4F",X"CD",X"CC",X"1D",X"FF",
		X"C9",X"FE",X"08",X"C3",X"48",X"0C",X"CB",X"79",X"CA",X"D0",X"16",X"C3",X"D5",X"16",X"21",X"88",
		X"63",X"34",X"C9",X"00",X"3E",X"66",X"32",X"0C",X"69",X"AF",X"32",X"24",X"69",X"32",X"2C",X"69",
		X"32",X"AF",X"62",X"21",X"88",X"63",X"34",X"C9",X"CD",X"1C",X"01",X"3E",X"00",X"32",X"38",X"6A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"05",X"69",X"36",X"2D",X"21",X"C4",
		X"75",X"11",X"20",X"00",X"3E",X"10",X"CD",X"14",X"05",X"21",X"8A",X"60",X"CD",X"B0",X"1F",X"36",
		X"03",X"C9",X"CD",X"6F",X"30",X"3A",X"13",X"69",X"FE",X"2C",X"D0",X"AF",X"32",X"00",X"69",X"32",
		X"04",X"69",X"32",X"0C",X"69",X"3E",X"6B",X"32",X"24",X"69",X"3D",X"32",X"2C",X"69",X"21",X"21",
		X"6A",X"34",X"21",X"88",X"63",X"34",X"C9",X"CD",X"6F",X"30",X"CD",X"6C",X"17",X"23",X"13",X"CD",
		X"83",X"17",X"3E",X"40",X"32",X"09",X"60",X"CD",X"0B",X"18",X"34",X"C9",X"11",X"03",X"00",X"21",
		X"2F",X"69",X"06",X"0A",X"A7",X"7E",X"ED",X"52",X"FE",X"19",X"D2",X"7F",X"17",X"36",X"00",X"2B",
		X"10",X"F2",X"C9",X"06",X"0A",X"7E",X"A7",X"C2",X"26",X"00",X"19",X"10",X"F8",X"C9",X"DF",X"2A",
		X"2A",X"62",X"23",X"7E",X"FE",X"7F",X"C2",X"9D",X"17",X"21",X"75",X"3A",X"7E",X"22",X"2A",X"62",
		X"32",X"27",X"62",X"11",X"00",X"05",X"CD",X"9F",X"30",X"AF",X"32",X"88",X"63",X"21",X"09",X"60",
		X"36",X"30",X"23",X"C3",X"3C",X"12",X"00",X"CD",X"39",X"0C",X"21",X"8A",X"60",X"36",X"0E",X"23",
		X"36",X"03",X"18",X"50",X"21",X"00",X"62",X"11",X"E0",X"64",X"01",X"20",X"00",X"ED",X"B0",X"FD",
		X"21",X"E0",X"64",X"3E",X"0F",X"FD",X"86",X"05",X"FD",X"77",X"05",X"C9",X"3A",X"27",X"62",X"FE",
		X"03",X"DD",X"21",X"00",X"66",X"C8",X"DD",X"21",X"90",X"65",X"C9",X"00",X"3A",X"27",X"62",X"FE",
		X"03",X"3A",X"10",X"69",X"C2",X"00",X"00",X"AF",X"32",X"00",X"69",X"32",X"04",X"69",X"32",X"20",
		X"69",X"32",X"24",X"69",X"32",X"28",X"69",X"32",X"2C",X"69",X"C9",X"3E",X"40",X"32",X"38",X"6A",
		X"21",X"88",X"63",X"C9",X"3E",X"20",X"32",X"09",X"60",X"3E",X"80",X"32",X"90",X"63",X"21",X"88",
		X"63",X"34",X"22",X"C0",X"63",X"C9",X"11",X"DB",X"FF",X"0E",X"0E",X"3E",X"10",X"06",X"05",X"77",
		X"23",X"10",X"FC",X"19",X"0D",X"C2",X"2D",X"18",X"C9",X"21",X"90",X"63",X"34",X"CA",X"65",X"18",
		X"7E",X"C3",X"33",X"1A",X"11",X"CF",X"39",X"CB",X"66",X"20",X"03",X"CD",X"16",X"11",X"EB",X"CD",
		X"4E",X"00",X"21",X"08",X"69",X"0E",X"00",X"FF",X"21",X"0B",X"69",X"0E",X"08",X"FF",X"C9",X"00",
		X"00",X"00",X"00",X"00",X"00",X"3E",X"20",X"32",X"09",X"60",X"21",X"88",X"63",X"34",X"C9",X"DF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"03",X"32",X"8C",X"60",X"21",X"88",X"63",X"34",X"C9",
		X"21",X"0B",X"69",X"0E",X"02",X"FF",X"CD",X"24",X"19",X"3A",X"1B",X"69",X"FE",X"C8",X"D4",X"06",
		X"19",X"FE",X"D6",X"D8",X"3E",X"20",X"32",X"15",X"69",X"00",X"00",X"00",X"00",X"00",X"00",X"21",
		X"C6",X"76",X"CD",X"26",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"04",X"00",X"01",X"28",
		X"02",X"21",X"03",X"69",X"CD",X"3D",X"00",X"3E",X"00",X"CD",X"F8",X"0F",X"3E",X"03",X"32",X"82",
		X"60",X"21",X"88",X"63",X"34",X"C9",X"CD",X"24",X"19",X"35",X"7E",X"FE",X"C0",X"D0",X"21",X"15",
		X"69",X"7E",X"EE",X"01",X"F6",X"20",X"77",X"CD",X"13",X"19",X"C3",X"3D",X"19",X"32",X"28",X"6A",
		X"32",X"40",X"63",X"3A",X"07",X"62",X"E6",X"7F",X"FE",X"04",X"C0",X"3E",X"0A",X"32",X"0F",X"62",
		X"C9",X"3A",X"27",X"62",X"FE",X"04",X"20",X"04",X"79",X"C6",X"10",X"4F",X"79",X"E6",X"7F",X"12",
		X"C9",X"C0",X"36",X"0A",X"C9",X"00",X"F5",X"3E",X"90",X"32",X"4D",X"69",X"3E",X"F4",X"32",X"55",
		X"69",X"F1",X"C9",X"21",X"8A",X"60",X"36",X"0C",X"3A",X"29",X"62",X"0F",X"38",X"02",X"36",X"0D",
		X"23",X"36",X"03",X"C9",X"3A",X"37",X"6A",X"C6",X"02",X"FE",X"F2",X"30",X"07",X"32",X"37",X"6A",
		X"21",X"AF",X"62",X"C9",X"3E",X"F1",X"32",X"35",X"6A",X"18",X"F5",X"00",X"00",X"2A",X"2A",X"62",
		X"23",X"7E",X"FE",X"7F",X"C2",X"4B",X"19",X"21",X"75",X"3A",X"7E",X"22",X"2A",X"62",X"00",X"00",
		X"00",X"21",X"29",X"62",X"34",X"11",X"00",X"05",X"CD",X"9F",X"30",X"AF",X"32",X"2E",X"62",X"00",
		X"00",X"00",X"21",X"88",X"63",X"34",X"C3",X"C7",X"1F",X"00",X"00",X"CD",X"52",X"08",X"3A",X"0E",
		X"60",X"C6",X"12",X"32",X"0A",X"60",X"C9",X"CD",X"EE",X"21",X"CD",X"BD",X"1D",X"CD",X"8C",X"1E",
		X"CD",X"C3",X"1A",X"CD",X"72",X"1F",X"CD",X"8F",X"2C",X"CD",X"03",X"2C",X"CD",X"3A",X"4D",X"CD",
		X"04",X"2E",X"CD",X"EA",X"24",X"CD",X"DB",X"2D",X"CD",X"D4",X"2E",X"CD",X"07",X"22",X"00",X"00",
		X"00",X"CD",X"85",X"2A",X"CD",X"46",X"1F",X"CD",X"FA",X"26",X"CD",X"F2",X"25",X"CD",X"DA",X"19",
		X"CD",X"FB",X"03",X"CD",X"08",X"28",X"CD",X"1D",X"28",X"CD",X"57",X"1E",X"CD",X"07",X"1A",X"CD",
		X"CB",X"2F",X"CD",X"F2",X"4E",X"CD",X"49",X"58",X"A7",X"C0",X"CD",X"1C",X"01",X"21",X"86",X"60",
		X"36",X"03",X"CD",X"B2",X"59",X"34",X"2B",X"36",X"40",X"C9",X"3A",X"94",X"6A",X"A7",X"C0",X"C3",
		X"B9",X"55",X"BE",X"CA",X"ED",X"19",X"2C",X"2C",X"2C",X"2C",X"10",X"F6",X"C9",X"3A",X"05",X"62",
		X"2C",X"2C",X"2C",X"BE",X"C0",X"2D",X"2D",X"CB",X"5E",X"C0",X"2D",X"22",X"43",X"63",X"AF",X"32",
		X"42",X"63",X"3C",X"32",X"40",X"63",X"C9",X"3A",X"86",X"63",X"EF",X"1E",X"1A",X"15",X"1A",X"1F",
		X"1A",X"2A",X"1A",X"00",X"00",X"AF",X"32",X"87",X"63",X"3E",X"02",X"32",X"86",X"63",X"C9",X"21",
		X"87",X"63",X"35",X"C0",X"3E",X"03",X"32",X"86",X"63",X"C9",X"3A",X"16",X"62",X"A7",X"C0",X"E1",
		X"C3",X"D2",X"19",X"FE",X"E0",X"F5",X"CC",X"40",X"1A",X"F1",X"E6",X"0F",X"C0",X"C3",X"44",X"18",
		X"3E",X"10",X"11",X"20",X"00",X"21",X"27",X"76",X"CD",X"14",X"05",X"21",X"A7",X"75",X"CD",X"14",
		X"05",X"21",X"48",X"77",X"11",X"CA",X"FF",X"0E",X"16",X"3E",X"10",X"06",X"16",X"77",X"23",X"10",
		X"FC",X"19",X"0D",X"20",X"F6",X"CD",X"76",X"1A",X"CD",X"BD",X"30",X"06",X"1C",X"21",X"58",X"69",
		X"36",X"00",X"23",X"10",X"FB",X"C9",X"DD",X"21",X"4C",X"69",X"DD",X"36",X"00",X"75",X"DD",X"36",
		X"08",X"85",X"DD",X"36",X"01",X"6A",X"DD",X"36",X"09",X"06",X"DD",X"36",X"03",X"F0",X"DD",X"36",
		X"0B",X"F0",X"21",X"88",X"63",X"C9",X"3A",X"27",X"62",X"FE",X"03",X"FD",X"36",X"01",X"3B",X"C0",
		X"FD",X"36",X"01",X"13",X"FD",X"36",X"02",X"0F",X"C9",X"3A",X"27",X"62",X"FE",X"03",X"3E",X"DD",
		X"28",X"02",X"3E",X"AD",X"DD",X"BE",X"03",X"D2",X"6C",X"2E",X"C3",X"5F",X"2E",X"00",X"00",X"00",
		X"00",X"00",X"00",X"CD",X"86",X"57",X"3D",X"CA",X"B2",X"1B",X"3A",X"1E",X"62",X"A7",X"C2",X"55",
		X"1B",X"3A",X"17",X"62",X"3D",X"CA",X"E6",X"1A",X"3A",X"15",X"62",X"3D",X"CA",X"B6",X"58",X"C3",
		X"31",X"58",X"17",X"DA",X"6E",X"1B",X"CD",X"1F",X"24",X"3A",X"10",X"60",X"1D",X"CA",X"F5",X"1A",
		X"CB",X"47",X"C2",X"8F",X"1C",X"15",X"CA",X"FE",X"1A",X"CB",X"4F",X"C2",X"AB",X"1C",X"3A",X"17",
		X"62",X"3D",X"C8",X"C9",X"05",X"62",X"C6",X"08",X"57",X"3A",X"03",X"62",X"F6",X"03",X"CB",X"97",
		X"01",X"15",X"00",X"CD",X"6E",X"23",X"F5",X"21",X"07",X"62",X"7E",X"E6",X"80",X"F6",X"06",X"77",
		X"21",X"1A",X"62",X"3E",X"04",X"B9",X"36",X"01",X"D2",X"2C",X"1B",X"35",X"F1",X"A7",X"CA",X"4E",
		X"1B",X"7E",X"A7",X"C0",X"2C",X"72",X"2C",X"70",X"3A",X"10",X"60",X"CB",X"5F",X"C2",X"86",X"40",
		X"3A",X"15",X"62",X"A7",X"C8",X"3A",X"10",X"60",X"CB",X"57",X"C3",X"F4",X"40",X"C9",X"2C",X"70",
		X"2C",X"72",X"C3",X"45",X"1B",X"21",X"1E",X"62",X"35",X"C0",X"3A",X"18",X"62",X"32",X"17",X"62",
		X"C3",X"A6",X"59",X"7E",X"E6",X"80",X"77",X"AF",X"32",X"02",X"62",X"C3",X"A6",X"1D",X"3E",X"01",
		X"CD",X"59",X"3A",X"21",X"10",X"62",X"3A",X"10",X"60",X"01",X"80",X"00",X"1F",X"DA",X"8A",X"1B",
		X"01",X"80",X"FF",X"1F",X"DA",X"8A",X"1B",X"01",X"00",X"00",X"AF",X"70",X"2C",X"71",X"2C",X"36",
		X"01",X"2C",X"36",X"48",X"2C",X"77",X"32",X"04",X"62",X"32",X"06",X"62",X"3A",X"07",X"62",X"E6",
		X"80",X"F6",X"0E",X"32",X"07",X"62",X"3A",X"05",X"62",X"32",X"0E",X"62",X"21",X"81",X"60",X"36",
		X"03",X"C9",X"DD",X"21",X"00",X"62",X"3A",X"03",X"62",X"DD",X"77",X"0B",X"3A",X"05",X"62",X"DD",
		X"77",X"0C",X"C3",X"92",X"47",X"CD",X"1F",X"24",X"15",X"C2",X"F2",X"1B",X"DD",X"36",X"10",X"00",
		X"DD",X"36",X"11",X"80",X"DD",X"CB",X"07",X"FE",X"3A",X"20",X"62",X"3D",X"CA",X"EC",X"1B",X"CD",
		X"07",X"24",X"DD",X"74",X"12",X"DD",X"75",X"13",X"DD",X"36",X"14",X"00",X"CD",X"9C",X"23",X"C3",
		X"05",X"1C",X"1D",X"C2",X"05",X"1C",X"DD",X"36",X"10",X"FF",X"DD",X"36",X"11",X"80",X"DD",X"CB",
		X"07",X"BE",X"C3",X"D8",X"1B",X"C3",X"5D",X"55",X"3D",X"CA",X"3A",X"1C",X"3A",X"1F",X"62",X"3D",
		X"CA",X"76",X"1C",X"3A",X"14",X"62",X"D6",X"14",X"C2",X"33",X"1C",X"3E",X"01",X"32",X"1F",X"62",
		X"CD",X"53",X"28",X"A7",X"CA",X"A6",X"1D",X"32",X"42",X"63",X"3E",X"01",X"32",X"40",X"63",X"CD",
		X"C2",X"0F",X"00",X"3C",X"CC",X"54",X"29",X"C3",X"78",X"44",X"05",X"CA",X"4F",X"1C",X"3C",X"32",
		X"1F",X"62",X"AF",X"21",X"10",X"62",X"06",X"05",X"77",X"2C",X"10",X"FC",X"C3",X"99",X"4A",X"CD",
		X"74",X"58",X"CD",X"84",X"58",X"EE",X"01",X"32",X"00",X"62",X"CD",X"C8",X"54",X"CD",X"FE",X"0B",
		X"F6",X"0F",X"77",X"00",X"00",X"C3",X"A2",X"58",X"AF",X"32",X"1F",X"62",X"3A",X"25",X"62",X"3D",
		X"CC",X"95",X"1D",X"C3",X"A1",X"4A",X"3A",X"05",X"62",X"21",X"0E",X"62",X"D6",X"18",X"BE",X"DA",
		X"78",X"44",X"3E",X"01",X"32",X"20",X"62",X"21",X"8C",X"60",X"36",X"03",X"C3",X"A6",X"1D",X"06",
		X"01",X"3A",X"0F",X"62",X"A7",X"C2",X"D2",X"1C",X"3A",X"02",X"62",X"47",X"3E",X"05",X"CD",X"09",
		X"30",X"32",X"02",X"62",X"E6",X"03",X"F6",X"80",X"C3",X"C2",X"1C",X"06",X"FF",X"3A",X"0F",X"62",
		X"A7",X"C2",X"D2",X"1C",X"3A",X"02",X"62",X"47",X"3E",X"01",X"CD",X"09",X"30",X"32",X"02",X"62",
		X"E6",X"03",X"21",X"07",X"62",X"77",X"1F",X"DC",X"8F",X"1D",X"3E",X"03",X"32",X"0F",X"62",X"C3",
		X"FA",X"11",X"21",X"03",X"62",X"7E",X"80",X"77",X"3A",X"27",X"62",X"3D",X"C2",X"EB",X"1C",X"CD",
		X"A9",X"49",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"0F",X"62",X"35",X"C3",
		X"A6",X"1D",X"3A",X"0F",X"62",X"A7",X"C2",X"8A",X"1D",X"CD",X"95",X"42",X"00",X"00",X"00",X"00",
		X"C3",X"11",X"1D",X"CD",X"96",X"56",X"A7",X"C2",X"76",X"1D",X"CD",X"A9",X"42",X"00",X"00",X"00",
		X"00",X"21",X"05",X"62",X"86",X"77",X"47",X"3A",X"22",X"62",X"EE",X"01",X"32",X"22",X"62",X"C2",
		X"51",X"1D",X"78",X"C6",X"08",X"21",X"1C",X"62",X"BE",X"CA",X"67",X"1D",X"2D",X"96",X"C3",X"C1",
		X"42",X"06",X"05",X"D6",X"08",X"CA",X"3F",X"1D",X"05",X"D6",X"04",X"CA",X"3F",X"1D",X"05",X"3E",
		X"80",X"21",X"07",X"62",X"A6",X"EE",X"80",X"B0",X"77",X"3E",X"01",X"32",X"15",X"62",X"C3",X"AC",
		X"1D",X"C3",X"6B",X"44",X"F6",X"03",X"CB",X"97",X"00",X"3A",X"24",X"62",X"EE",X"01",X"32",X"24",
		X"62",X"CC",X"8F",X"1D",X"C3",X"49",X"1D",X"3E",X"06",X"32",X"07",X"62",X"AF",X"32",X"19",X"62",
		X"32",X"15",X"62",X"C3",X"A6",X"1D",X"3A",X"1A",X"62",X"A7",X"CA",X"8A",X"1D",X"32",X"19",X"62",
		X"3A",X"1C",X"62",X"D6",X"13",X"21",X"05",X"62",X"BE",X"D0",X"21",X"0F",X"62",X"35",X"C9",X"3E",
		X"03",X"CD",X"84",X"2E",X"C9",X"32",X"25",X"62",X"3A",X"27",X"62",X"3D",X"C8",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C9",X"C3",X"AA",X"40",X"C3",X"AA",X"40",X"3A",X"10",X"60",X"E6",
		X"0C",X"CA",X"AA",X"40",X"C3",X"D0",X"42",X"3A",X"05",X"62",X"2C",X"77",X"C9",X"CD",X"0F",X"1E",
		X"EF",X"49",X"1E",X"C9",X"1D",X"4A",X"1E",X"00",X"00",X"C3",X"16",X"5D",X"3A",X"1A",X"60",X"E6",
		X"1F",X"20",X"08",X"3A",X"A8",X"63",X"EE",X"40",X"32",X"A8",X"63",X"3A",X"34",X"6A",X"F5",X"FE",
		X"44",X"CC",X"00",X"1E",X"FE",X"38",X"CC",X"0B",X"1E",X"F1",X"FE",X"28",X"20",X"0E",X"21",X"3C",
		X"6A",X"36",X"5B",X"23",X"36",X"4C",X"23",X"36",X"0B",X"23",X"36",X"14",X"21",X"08",X"69",X"C9",
		X"3E",X"06",X"32",X"4D",X"69",X"C6",X"64",X"32",X"55",X"69",X"C9",X"3E",X"05",X"18",X"F3",X"3A",
		X"1A",X"60",X"E6",X"0F",X"20",X"08",X"3A",X"3A",X"6A",X"EE",X"02",X"32",X"3A",X"6A",X"3A",X"40",
		X"63",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"CD",X"9F",X"30",X"3A",X"05",X"62",X"C6",X"14",
		X"4F",X"3A",X"03",X"62",X"00",X"00",X"21",X"30",X"6A",X"77",X"2C",X"70",X"2C",X"36",X"01",X"2C",
		X"71",X"3E",X"05",X"F7",X"00",X"00",X"00",X"00",X"00",X"C9",X"21",X"41",X"63",X"35",X"C0",X"AF",
		X"32",X"30",X"6A",X"C3",X"DD",X"18",X"C9",X"3A",X"27",X"62",X"FE",X"03",X"CA",X"80",X"1E",X"C3",
		X"0C",X"47",X"FD",X"21",X"58",X"69",X"3A",X"27",X"62",X"FE",X"01",X"06",X"05",X"C8",X"3A",X"29",
		X"62",X"C6",X"04",X"FE",X"0A",X"38",X"02",X"3E",X"0A",X"47",X"C9",X"00",X"00",X"00",X"00",X"00",
		X"3A",X"90",X"62",X"A7",X"C0",X"3E",X"16",X"32",X"0A",X"60",X"E1",X"C9",X"3A",X"50",X"63",X"A7",
		X"C8",X"CD",X"96",X"1E",X"E1",X"C9",X"3A",X"45",X"63",X"EF",X"A0",X"1E",X"09",X"1F",X"23",X"1F",
		X"3A",X"52",X"63",X"FE",X"65",X"21",X"58",X"69",X"CA",X"B4",X"1E",X"21",X"D0",X"69",X"DA",X"B4",
		X"1E",X"21",X"80",X"69",X"DD",X"2A",X"51",X"63",X"16",X"00",X"3A",X"53",X"63",X"5F",X"01",X"04",
		X"00",X"3A",X"54",X"63",X"A7",X"CA",X"CF",X"1E",X"09",X"DD",X"19",X"3D",X"C2",X"C8",X"1E",X"CD",
		X"C5",X"56",X"00",X"DD",X"7E",X"15",X"A7",X"3E",X"02",X"CA",X"DE",X"1E",X"3E",X"04",X"00",X"00",
		X"00",X"01",X"2C",X"6A",X"7E",X"36",X"00",X"02",X"0C",X"2C",X"3E",X"60",X"02",X"0C",X"2C",X"3E",
		X"0E",X"02",X"0C",X"2C",X"7E",X"02",X"21",X"45",X"63",X"34",X"2C",X"36",X"06",X"2C",X"36",X"05",
		X"3E",X"03",X"32",X"84",X"60",X"00",X"00",X"00",X"C9",X"21",X"46",X"63",X"35",X"C0",X"36",X"06",
		X"2C",X"35",X"CA",X"1D",X"1F",X"21",X"2D",X"6A",X"7E",X"EE",X"01",X"77",X"C9",X"36",X"04",X"2D",
		X"2D",X"34",X"C9",X"21",X"46",X"63",X"35",X"C0",X"36",X"0C",X"2C",X"35",X"CA",X"34",X"1F",X"21",
		X"2D",X"6A",X"34",X"C9",X"2D",X"2D",X"AF",X"77",X"32",X"50",X"63",X"3C",X"32",X"40",X"63",X"21",
		X"2C",X"6A",X"22",X"43",X"63",X"C9",X"3A",X"21",X"62",X"A7",X"C8",X"AF",X"32",X"04",X"62",X"32",
		X"06",X"62",X"32",X"21",X"62",X"32",X"10",X"62",X"32",X"11",X"62",X"32",X"12",X"62",X"32",X"13",
		X"62",X"32",X"14",X"62",X"3C",X"32",X"16",X"62",X"32",X"1F",X"62",X"3A",X"05",X"62",X"32",X"0E",
		X"62",X"C9",X"CD",X"7D",X"40",X"00",X"C0",X"DD",X"21",X"00",X"67",X"21",X"80",X"69",X"CD",X"33",
		X"11",X"00",X"00",X"DD",X"7E",X"00",X"3D",X"CA",X"93",X"1F",X"2C",X"2C",X"2C",X"2C",X"DD",X"19",
		X"10",X"F1",X"C9",X"DD",X"7E",X"01",X"3D",X"CA",X"EC",X"20",X"C3",X"A6",X"50",X"1F",X"DA",X"AC",
		X"1F",X"1F",X"DA",X"E5",X"1F",X"1F",X"DA",X"EF",X"1F",X"C3",X"8B",X"55",X"D9",X"C3",X"08",X"51",
		X"3A",X"27",X"62",X"06",X"09",X"FE",X"02",X"28",X"0B",X"04",X"FE",X"01",X"28",X"06",X"04",X"FE",
		X"04",X"28",X"01",X"04",X"70",X"23",X"C9",X"3E",X"03",X"32",X"82",X"6A",X"C9",X"76",X"DD",X"7E",
		X"0F",X"3D",X"C2",X"DF",X"1F",X"C3",X"59",X"51",X"EE",X"03",X"CD",X"30",X"0D",X"00",X"00",X"DD",
		X"77",X"0F",X"C3",X"BA",X"21",X"D9",X"01",X"00",X"01",X"DD",X"34",X"03",X"C3",X"F6",X"1F",X"D9",
		X"01",X"04",X"FF",X"DD",X"35",X"03",X"C3",X"16",X"29",X"DD",X"6E",X"05",X"7C",X"E6",X"07",X"FE",
		X"03",X"CA",X"5F",X"21",X"2D",X"2D",X"2D",X"CD",X"33",X"23",X"2C",X"2C",X"2C",X"7D",X"DD",X"77",
		X"05",X"CD",X"A5",X"4A",X"CD",X"B4",X"24",X"DD",X"7E",X"03",X"FE",X"0A",X"DA",X"57",X"16",X"FE",
		X"F8",X"DA",X"53",X"54",X"AF",X"DD",X"77",X"10",X"DD",X"36",X"11",X"60",X"C3",X"38",X"20",X"AF",
		X"DD",X"36",X"10",X"FF",X"DD",X"36",X"11",X"A0",X"DD",X"36",X"12",X"FF",X"DD",X"36",X"13",X"F0",
		X"DD",X"77",X"14",X"DD",X"77",X"0E",X"DD",X"77",X"04",X"DD",X"77",X"06",X"DD",X"36",X"02",X"08",
		X"C3",X"BA",X"21",X"D9",X"CD",X"9C",X"23",X"CD",X"76",X"51",X"A7",X"C2",X"83",X"20",X"DD",X"7E",
		X"03",X"C6",X"08",X"FE",X"10",X"DA",X"79",X"20",X"CD",X"B4",X"24",X"DD",X"7E",X"10",X"E6",X"01",
		X"07",X"07",X"4F",X"CD",X"DE",X"23",X"C3",X"BA",X"21",X"AF",X"DD",X"77",X"00",X"DD",X"77",X"03",
		X"C3",X"8C",X"51",X"DD",X"34",X"0E",X"DD",X"7E",X"0E",X"3D",X"CA",X"A2",X"20",X"3D",X"CA",X"C3",
		X"20",X"DD",X"7E",X"10",X"3D",X"3E",X"04",X"C2",X"9C",X"20",X"3E",X"02",X"DD",X"77",X"02",X"C3",
		X"BA",X"21",X"DD",X"7E",X"15",X"A7",X"C2",X"B5",X"20",X"21",X"05",X"62",X"DD",X"7E",X"05",X"D6",
		X"16",X"BE",X"D2",X"C3",X"20",X"DD",X"35",X"C9",X"00",X"C2",X"E1",X"20",X"DD",X"77",X"11",X"DD",
		X"36",X"10",X"FF",X"CD",X"07",X"24",X"CB",X"3C",X"CB",X"1D",X"CB",X"3C",X"CB",X"1D",X"DD",X"74",
		X"12",X"DD",X"75",X"13",X"AF",X"DD",X"77",X"14",X"DD",X"77",X"04",X"DD",X"77",X"06",X"C3",X"BA",
		X"21",X"DD",X"36",X"10",X"01",X"DD",X"36",X"11",X"00",X"C3",X"C3",X"20",X"D9",X"CD",X"9C",X"23",
		X"7C",X"D6",X"1A",X"DD",X"46",X"19",X"B8",X"DA",X"04",X"21",X"CD",X"80",X"55",X"A7",X"C2",X"18",
		X"21",X"CD",X"B4",X"24",X"DD",X"7E",X"03",X"C6",X"08",X"FE",X"10",X"D2",X"CE",X"1F",X"AF",X"DD",
		X"77",X"00",X"DD",X"77",X"03",X"C3",X"BA",X"21",X"C3",X"93",X"51",X"3A",X"08",X"69",X"D6",X"05",
		X"32",X"08",X"69",X"3A",X"0C",X"69",X"C6",X"05",X"32",X"0C",X"69",X"F1",X"FE",X"60",X"D8",X"3A",
		X"09",X"60",X"E6",X"1F",X"CB",X"47",X"0E",X"00",X"28",X"08",X"FE",X"10",X"0E",X"FF",X"30",X"02",
		X"0E",X"01",X"3A",X"80",X"6A",X"A7",X"C5",X"CC",X"EF",X"5B",X"C1",X"06",X"03",X"11",X"08",X"00",
		X"DD",X"21",X"4C",X"69",X"DD",X"34",X"00",X"DD",X"7E",X"00",X"E6",X"03",X"C3",X"FF",X"3E",X"CD",
		X"A6",X"51",X"57",X"7C",X"01",X"15",X"00",X"C3",X"87",X"5C",X"C3",X"BA",X"21",X"CD",X"6E",X"23",
		X"3D",X"C0",X"C3",X"B3",X"51",X"DD",X"77",X"17",X"3A",X"48",X"63",X"A7",X"CA",X"B2",X"21",X"3A",
		X"05",X"62",X"D6",X"10",X"BA",X"D8",X"3A",X"80",X"63",X"1F",X"3C",X"47",X"3A",X"18",X"60",X"4F",
		X"E6",X"03",X"B8",X"D0",X"21",X"10",X"60",X"3A",X"03",X"62",X"BB",X"CA",X"B2",X"21",X"D2",X"A9",
		X"21",X"CB",X"46",X"CA",X"AE",X"21",X"C3",X"B2",X"21",X"CB",X"4E",X"C2",X"B2",X"21",X"79",X"E6",
		X"18",X"C0",X"CD",X"D2",X"47",X"DD",X"36",X"02",X"01",X"C9",X"D9",X"DD",X"7E",X"03",X"77",X"2C",
		X"DD",X"7E",X"07",X"77",X"2C",X"DD",X"7E",X"08",X"77",X"2C",X"DD",X"7E",X"05",X"77",X"C3",X"8D",
		X"1F",X"80",X"50",X"04",X"05",X"01",X"AF",X"04",X"60",X"01",X"20",X"81",X"55",X"08",X"20",X"01",
		X"30",X"81",X"16",X"01",X"20",X"81",X"20",X"82",X"40",X"04",X"18",X"01",X"30",X"04",X"11",X"D1",
		X"21",X"21",X"CC",X"63",X"7E",X"07",X"83",X"5F",X"1A",X"32",X"10",X"60",X"2C",X"7E",X"35",X"A7",
		X"C0",X"1C",X"1A",X"77",X"2D",X"34",X"C9",X"3E",X"02",X"F7",X"3A",X"1A",X"60",X"1F",X"21",X"80",
		X"62",X"7E",X"DA",X"19",X"22",X"21",X"88",X"62",X"7E",X"E5",X"EF",X"27",X"22",X"59",X"22",X"99",
		X"22",X"A2",X"22",X"00",X"00",X"00",X"00",X"E1",X"2C",X"35",X"C2",X"3A",X"22",X"2D",X"34",X"2C",
		X"2C",X"CD",X"43",X"22",X"3E",X"01",X"32",X"1A",X"62",X"C9",X"2C",X"CD",X"43",X"22",X"AF",X"32",
		X"1A",X"62",X"C9",X"3A",X"05",X"62",X"FE",X"7A",X"D2",X"57",X"22",X"3A",X"16",X"62",X"A7",X"C2",
		X"57",X"22",X"3A",X"03",X"62",X"BE",X"C8",X"E1",X"C9",X"E1",X"2C",X"2C",X"2C",X"2C",X"35",X"C0",
		X"3E",X"04",X"77",X"2D",X"34",X"CD",X"BD",X"22",X"3E",X"78",X"BE",X"C2",X"75",X"22",X"2D",X"2D",
		X"2D",X"34",X"2C",X"2C",X"2C",X"2D",X"CD",X"43",X"22",X"3A",X"05",X"62",X"FE",X"68",X"D2",X"8A",
		X"22",X"21",X"05",X"62",X"34",X"21",X"4F",X"69",X"34",X"C9",X"1F",X"DA",X"81",X"22",X"1F",X"3E",
		X"01",X"DA",X"95",X"22",X"AF",X"32",X"22",X"62",X"C9",X"E1",X"3A",X"18",X"60",X"E6",X"3C",X"C0",
		X"34",X"C9",X"E1",X"2C",X"2C",X"2C",X"2C",X"35",X"C0",X"36",X"02",X"2D",X"35",X"CD",X"BD",X"22",
		X"3E",X"68",X"BE",X"C0",X"AF",X"06",X"80",X"2D",X"2D",X"70",X"2D",X"77",X"C9",X"7E",X"CB",X"5D",
		X"11",X"4B",X"69",X"C2",X"C9",X"22",X"11",X"47",X"69",X"12",X"C9",X"3A",X"48",X"63",X"A7",X"CA",
		X"E1",X"22",X"3A",X"80",X"63",X"3D",X"EF",X"F6",X"22",X"F6",X"22",X"03",X"23",X"03",X"23",X"1A",
		X"23",X"3A",X"29",X"62",X"47",X"05",X"3E",X"01",X"CA",X"F9",X"22",X"05",X"3E",X"B1",X"CA",X"F9",
		X"22",X"3E",X"E9",X"C3",X"F9",X"22",X"3A",X"18",X"60",X"DD",X"77",X"11",X"E6",X"01",X"3D",X"DD",
		X"77",X"10",X"C9",X"3A",X"18",X"60",X"DD",X"77",X"11",X"3A",X"03",X"62",X"DD",X"BE",X"03",X"3E",
		X"01",X"D2",X"16",X"23",X"3D",X"3D",X"DD",X"77",X"10",X"C9",X"3A",X"03",X"62",X"DD",X"96",X"03",
		X"0E",X"FF",X"DA",X"26",X"23",X"0C",X"07",X"CB",X"11",X"07",X"CB",X"11",X"DD",X"71",X"10",X"DD",
		X"77",X"11",X"C9",X"3E",X"0F",X"A4",X"05",X"CA",X"42",X"23",X"C3",X"23",X"58",X"06",X"FF",X"C3",
		X"47",X"23",X"FE",X"01",X"D0",X"06",X"01",X"3E",X"F0",X"BD",X"CA",X"60",X"23",X"3E",X"38",X"BD",
		X"DA",X"66",X"23",X"7D",X"CB",X"6F",X"CA",X"5C",X"23",X"00",X"6F",X"C9",X"00",X"C3",X"5A",X"23",
		X"CB",X"7C",X"C2",X"59",X"23",X"C9",X"C3",X"74",X"54",X"D8",X"7D",X"C3",X"C1",X"51",X"21",X"00",
		X"63",X"ED",X"B1",X"C2",X"9A",X"23",X"E5",X"C5",X"01",X"14",X"00",X"09",X"0C",X"5F",X"7A",X"BE",
		X"CA",X"8F",X"23",X"09",X"BE",X"CA",X"95",X"23",X"57",X"7B",X"C1",X"E1",X"C3",X"71",X"23",X"09",
		X"3E",X"01",X"C3",X"98",X"23",X"AF",X"ED",X"42",X"C1",X"46",X"E1",X"C9",X"DD",X"7E",X"04",X"DD",
		X"86",X"11",X"DD",X"77",X"04",X"DD",X"7E",X"03",X"DD",X"8E",X"10",X"DD",X"77",X"03",X"DD",X"7E",
		X"06",X"DD",X"96",X"13",X"6F",X"DD",X"7E",X"05",X"DD",X"9E",X"12",X"67",X"DD",X"7E",X"14",X"A7",
		X"17",X"3C",X"06",X"00",X"CB",X"10",X"CB",X"27",X"CB",X"10",X"CB",X"27",X"CB",X"10",X"CB",X"27",
		X"CB",X"10",X"4F",X"09",X"CD",X"DC",X"58",X"DD",X"75",X"06",X"DD",X"34",X"14",X"C9",X"DD",X"7E",
		X"0F",X"3D",X"C3",X"E2",X"51",X"AF",X"DD",X"CB",X"07",X"26",X"17",X"DD",X"CB",X"08",X"26",X"17",
		X"47",X"3E",X"03",X"B1",X"CD",X"09",X"30",X"1F",X"DD",X"CB",X"08",X"1E",X"1F",X"DD",X"CB",X"07",
		X"1E",X"3E",X"04",X"DD",X"77",X"0F",X"C9",X"DD",X"7E",X"14",X"07",X"07",X"07",X"07",X"4F",X"E6",
		X"0F",X"67",X"79",X"E6",X"F0",X"6F",X"DD",X"4E",X"13",X"DD",X"46",X"12",X"ED",X"42",X"C9",X"11",
		X"00",X"01",X"3A",X"03",X"62",X"FE",X"13",X"D8",X"15",X"1C",X"FE",X"EC",X"D0",X"1D",X"CD",X"49",
		X"40",X"00",X"C8",X"3A",X"05",X"62",X"FE",X"58",X"D0",X"3A",X"03",X"62",X"FE",X"50",X"D0",X"14",
		X"C9",X"21",X"FB",X"37",X"3E",X"88",X"06",X"07",X"86",X"23",X"10",X"FC",X"DD",X"21",X"00",X"63",
		X"A7",X"CA",X"58",X"24",X"DD",X"21",X"00",X"64",X"3A",X"27",X"62",X"3D",X"21",X"86",X"3B",X"CA",
		X"75",X"24",X"3D",X"21",X"C6",X"3A",X"CA",X"75",X"24",X"3D",X"21",X"BE",X"3F",X"CA",X"75",X"24",
		X"21",X"40",X"3C",X"00",X"00",X"11",X"05",X"00",X"7E",X"FE",X"04",X"38",X"0B",X"FE",X"AA",X"C8",
		X"FE",X"0E",X"28",X"04",X"19",X"18",X"F1",X"24",X"23",X"7E",X"DD",X"77",X"00",X"23",X"7E",X"DD",
		X"77",X"15",X"23",X"23",X"7E",X"DD",X"77",X"2A",X"DD",X"23",X"23",X"C3",X"78",X"24",X"23",X"7E",
		X"FD",X"77",X"00",X"23",X"7E",X"FD",X"77",X"15",X"23",X"23",X"7E",X"FD",X"77",X"2A",X"FD",X"23",
		X"23",X"C3",X"78",X"24",X"DD",X"7E",X"05",X"FE",X"FA",X"D8",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"DD",X"7E",X"15",X"A7",X"CA",X"D0",X"24",X"3E",X"03",X"32",X"B9",X"62",X"AF",
		X"DD",X"77",X"00",X"DD",X"77",X"03",X"00",X"00",X"00",X"00",X"00",X"E1",X"3A",X"48",X"63",X"A7",
		X"C2",X"BA",X"21",X"3C",X"32",X"48",X"63",X"C3",X"BA",X"21",X"3E",X"01",X"F7",X"CD",X"23",X"25",
		X"CD",X"91",X"25",X"DD",X"21",X"A0",X"65",X"06",X"05",X"21",X"30",X"69",X"DD",X"7E",X"00",X"A7",
		X"CA",X"1C",X"25",X"DD",X"7E",X"03",X"77",X"2C",X"DD",X"7E",X"07",X"77",X"2C",X"DD",X"7E",X"08",
		X"77",X"2C",X"DD",X"7E",X"05",X"77",X"2C",X"DD",X"19",X"10",X"E1",X"C3",X"56",X"53",X"04",X"6F",
		X"C3",X"17",X"25",X"21",X"9B",X"63",X"7E",X"A7",X"C2",X"8F",X"25",X"3A",X"9A",X"63",X"A7",X"C8",
		X"06",X"05",X"11",X"10",X"00",X"DD",X"21",X"B0",X"65",X"DD",X"CB",X"00",X"46",X"CA",X"45",X"25",
		X"DD",X"19",X"10",X"F5",X"C9",X"CD",X"57",X"00",X"3E",X"D0",X"32",X"B5",X"65",X"3E",X"F4",X"32",
		X"C5",X"65",X"3E",X"A3",X"32",X"E5",X"65",X"C3",X"76",X"25",X"05",X"CC",X"3A",X"A6",X"62",X"07",
		X"DD",X"36",X"03",X"07",X"D2",X"76",X"25",X"DD",X"36",X"03",X"F8",X"C3",X"76",X"25",X"CD",X"57",
		X"00",X"FE",X"68",X"C3",X"60",X"25",X"DD",X"36",X"00",X"01",X"DD",X"36",X"07",X"4B",X"DD",X"36",
		X"09",X"08",X"DD",X"36",X"0A",X"03",X"3E",X"7C",X"32",X"9B",X"63",X"AF",X"32",X"9A",X"63",X"35",
		X"C9",X"DD",X"21",X"B0",X"65",X"11",X"10",X"00",X"06",X"03",X"DD",X"CB",X"00",X"46",X"CA",X"BB",
		X"25",X"DD",X"7E",X"03",X"67",X"DD",X"7E",X"05",X"C3",X"53",X"49",X"25",X"DD",X"7E",X"05",X"FE",
		X"7C",X"CA",X"C0",X"25",X"3A",X"A6",X"63",X"84",X"CD",X"5F",X"4A",X"DD",X"19",X"10",X"DB",X"C9",
		X"7C",X"FE",X"80",X"CA",X"D6",X"25",X"3A",X"A5",X"63",X"D2",X"CF",X"25",X"3A",X"A4",X"63",X"84",
		X"DD",X"77",X"03",X"C3",X"BB",X"25",X"21",X"B8",X"69",X"3E",X"06",X"90",X"CA",X"E7",X"25",X"2C",
		X"2C",X"2C",X"2C",X"3D",X"C3",X"DC",X"25",X"AF",X"DD",X"77",X"00",X"DD",X"77",X"03",X"77",X"C3",
		X"BB",X"25",X"3E",X"01",X"F7",X"CD",X"25",X"59",X"CD",X"3B",X"59",X"CD",X"51",X"59",X"CD",X"D3",
		X"2A",X"C9",X"CD",X"84",X"49",X"0F",X"DA",X"16",X"26",X"21",X"A0",X"62",X"35",X"C2",X"16",X"26",
		X"36",X"53",X"2C",X"CD",X"DE",X"26",X"21",X"A1",X"62",X"CD",X"E9",X"26",X"32",X"A3",X"63",X"3A",
		X"1A",X"60",X"E6",X"1F",X"FE",X"01",X"C0",X"11",X"E4",X"69",X"EB",X"00",X"00",X"00",X"C9",X"3A",
		X"AA",X"63",X"3D",X"30",X"02",X"3E",X"02",X"32",X"AA",X"63",X"21",X"09",X"60",X"3A",X"1A",X"60",
		X"E6",X"01",X"20",X"10",X"3A",X"0D",X"6A",X"EE",X"0E",X"32",X"0D",X"6A",X"3C",X"32",X"11",X"6A",
		X"3C",X"32",X"15",X"6A",X"35",X"7E",X"E6",X"0F",X"20",X"13",X"2A",X"A8",X"63",X"7E",X"FE",X"7F",
		X"20",X"03",X"21",X"B0",X"27",X"7E",X"32",X"A7",X"63",X"23",X"22",X"A8",X"63",X"06",X"0C",X"21",
		X"A0",X"6A",X"CD",X"CF",X"5B",X"38",X"02",X"10",X"F9",X"06",X"0C",X"DD",X"21",X"A0",X"6A",X"11",
		X"3F",X"5C",X"1A",X"6F",X"13",X"1A",X"67",X"13",X"DD",X"7E",X"00",X"77",X"DD",X"23",X"23",X"23",
		X"23",X"3A",X"09",X"60",X"E6",X"01",X"3E",X"00",X"28",X"03",X"3A",X"A7",X"63",X"86",X"77",X"10",
		X"E1",X"3A",X"18",X"69",X"32",X"20",X"69",X"32",X"28",X"69",X"3A",X"1C",X"69",X"32",X"24",X"69",
		X"32",X"2C",X"69",X"3A",X"10",X"69",X"32",X"00",X"69",X"32",X"04",X"69",X"F5",X"3A",X"1B",X"69",
		X"D6",X"02",X"32",X"23",X"69",X"32",X"27",X"69",X"32",X"03",X"69",X"3A",X"1F",X"69",X"C6",X"10",
		X"32",X"2B",X"69",X"32",X"2F",X"69",X"32",X"07",X"69",X"C3",X"1B",X"21",X"00",X"00",X"CB",X"7E",
		X"CA",X"E6",X"26",X"36",X"02",X"C9",X"36",X"FE",X"C9",X"C3",X"8B",X"49",X"00",X"00",X"00",X"CB",
		X"7E",X"3E",X"FF",X"C3",X"3E",X"54",X"3E",X"01",X"77",X"C9",X"C3",X"B3",X"5A",X"CD",X"1C",X"01",
		X"DF",X"CD",X"74",X"08",X"3E",X"00",X"32",X"86",X"7D",X"3E",X"00",X"32",X"87",X"7D",X"11",X"9E",
		X"27",X"CD",X"A7",X"0D",X"06",X"04",X"21",X"A4",X"27",X"CD",X"42",X"0B",X"06",X"06",X"3E",X"54",
		X"0E",X"0E",X"21",X"0D",X"6A",X"77",X"23",X"36",X"0A",X"23",X"71",X"F5",X"78",X"FE",X"04",X"20",
		X"02",X"0E",X"1E",X"F1",X"23",X"23",X"3C",X"10",X"EC",X"21",X"F7",X"39",X"CD",X"4E",X"00",X"11",
		X"04",X"00",X"21",X"0B",X"69",X"01",X"10",X"0C",X"CD",X"3D",X"00",X"11",X"A0",X"6A",X"21",X"00",
		X"69",X"06",X"0C",X"AF",X"77",X"12",X"23",X"23",X"23",X"23",X"13",X"10",X"F6",X"3E",X"06",X"32",
		X"89",X"60",X"21",X"B0",X"27",X"22",X"A8",X"63",X"22",X"BB",X"63",X"7E",X"32",X"A7",X"63",X"3E",
		X"2D",X"32",X"01",X"69",X"32",X"05",X"69",X"3E",X"08",X"32",X"02",X"69",X"3E",X"88",X"32",X"06",
		X"69",X"3A",X"23",X"69",X"32",X"03",X"69",X"3A",X"2B",X"69",X"32",X"07",X"69",X"3E",X"02",X"32",
		X"AA",X"63",X"AF",X"32",X"80",X"6A",X"21",X"09",X"60",X"36",X"A0",X"23",X"34",X"C9",X"0A",X"EF",
		X"F8",X"10",X"F8",X"AA",X"F8",X"88",X"07",X"A8",X"08",X"EC",X"07",X"A8",X"00",X"4F",X"0F",X"9C",
		X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",
		X"6B",X"43",X"02",X"BE",X"93",X"43",X"02",X"BE",X"6B",X"43",X"02",X"50",X"93",X"43",X"02",X"50",
		X"A2",X"17",X"00",X"40",X"5C",X"97",X"00",X"40",X"67",X"4A",X"80",X"18",X"97",X"4A",X"80",X"18",
		X"00",X"00",X"00",X"00",X"DD",X"36",X"00",X"01",X"DD",X"36",X"03",X"37",X"DD",X"36",X"05",X"F8",
		X"DD",X"36",X"0D",X"08",X"36",X"34",X"35",X"C9",X"FD",X"21",X"00",X"62",X"3A",X"05",X"62",X"4F",
		X"21",X"08",X"0D",X"CD",X"6F",X"28",X"A7",X"C8",X"3D",X"32",X"00",X"62",X"C9",X"AF",X"32",X"99",
		X"6A",X"C3",X"FB",X"54",X"80",X"66",X"FD",X"CB",X"01",X"46",X"C2",X"32",X"28",X"FD",X"19",X"10",
		X"F5",X"C9",X"FD",X"4E",X"05",X"FD",X"66",X"09",X"FD",X"6E",X"0A",X"CD",X"6F",X"28",X"A7",X"C8",
		X"CD",X"16",X"55",X"3A",X"B9",X"63",X"90",X"32",X"54",X"63",X"7B",X"32",X"53",X"63",X"C3",X"1D",
		X"55",X"63",X"C9",X"CD",X"C4",X"17",X"00",X"3A",X"05",X"62",X"C6",X"0C",X"4F",X"3A",X"10",X"60",
		X"E6",X"03",X"21",X"0A",X"05",X"CA",X"6B",X"28",X"21",X"0A",X"13",X"CD",X"88",X"3E",X"C9",X"3A",
		X"27",X"62",X"E5",X"EF",X"00",X"00",X"E0",X"28",X"80",X"28",X"E0",X"28",X"80",X"28",X"00",X"00",
		X"E1",X"06",X"0A",X"78",X"32",X"B9",X"63",X"11",X"20",X"00",X"DD",X"21",X"00",X"67",X"CD",X"13",
		X"29",X"06",X"05",X"78",X"32",X"B9",X"63",X"1E",X"20",X"DD",X"21",X"00",X"64",X"CD",X"13",X"29",
		X"06",X"01",X"78",X"32",X"B9",X"63",X"1E",X"00",X"DD",X"21",X"A0",X"66",X"CD",X"13",X"29",X"C9",
		X"E1",X"06",X"05",X"78",X"32",X"B9",X"63",X"11",X"20",X"00",X"DD",X"21",X"00",X"64",X"CD",X"13",
		X"29",X"06",X"06",X"78",X"32",X"B9",X"63",X"1E",X"10",X"DD",X"21",X"A0",X"65",X"00",X"00",X"00",
		X"06",X"01",X"78",X"32",X"B9",X"63",X"1E",X"00",X"DD",X"21",X"A0",X"66",X"CD",X"13",X"29",X"C9",
		X"E1",X"06",X"05",X"78",X"32",X"B9",X"63",X"11",X"20",X"00",X"DD",X"21",X"00",X"64",X"CD",X"13",
		X"29",X"06",X"0A",X"78",X"32",X"B9",X"63",X"1E",X"10",X"DD",X"21",X"00",X"65",X"C3",X"11",X"53",
		X"C9",X"E1",X"06",X"05",X"78",X"32",X"B9",X"63",X"11",X"20",X"00",X"DD",X"21",X"00",X"64",X"CD",
		X"13",X"29",X"C9",X"C3",X"CD",X"4A",X"DD",X"7E",X"0C",X"A7",X"20",X"29",X"DD",X"7E",X"05",X"FE",
		X"47",X"20",X"03",X"DD",X"35",X"03",X"FE",X"58",X"20",X"03",X"DD",X"34",X"03",X"3A",X"29",X"62",
		X"FE",X"04",X"38",X"11",X"DD",X"7E",X"05",X"FE",X"7F",X"20",X"03",X"DD",X"34",X"03",X"FE",X"90",
		X"20",X"03",X"DD",X"35",X"03",X"CD",X"9A",X"55",X"C3",X"F9",X"1F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"3E",X"0B",X"F7",X"CD",X"74",X"29",X"32",X"18",X"62",X"0F",X"0F",X"32",
		X"85",X"60",X"78",X"A7",X"C8",X"FE",X"01",X"CA",X"6F",X"29",X"DD",X"36",X"01",X"01",X"C9",X"DD",
		X"36",X"11",X"01",X"C9",X"FD",X"21",X"00",X"62",X"3A",X"05",X"62",X"4F",X"21",X"08",X"04",X"06",
		X"02",X"11",X"10",X"00",X"DD",X"21",X"80",X"66",X"CD",X"13",X"29",X"C9",X"2A",X"C8",X"63",X"7D",
		X"C6",X"0E",X"6F",X"56",X"2C",X"7E",X"C6",X"0C",X"5F",X"EB",X"CD",X"F0",X"2F",X"7E",X"FE",X"B1",
		X"28",X"08",X"FE",X"D0",X"DA",X"AC",X"29",X"00",X"00",X"00",X"AF",X"C9",X"3E",X"01",X"C9",X"3E",
		X"05",X"F7",X"FD",X"21",X"00",X"62",X"3A",X"05",X"62",X"4F",X"21",X"08",X"02",X"CD",X"22",X"2A",
		X"A7",X"CA",X"20",X"2A",X"3E",X"04",X"90",X"CA",X"D0",X"29",X"DD",X"19",X"3D",X"C3",X"C7",X"29",
		X"DD",X"7E",X"05",X"D6",X"04",X"57",X"3A",X"0C",X"62",X"C6",X"05",X"BA",X"D2",X"EE",X"29",X"7A",
		X"D6",X"08",X"C3",X"8D",X"58",X"3E",X"01",X"47",X"CD",X"68",X"4A",X"33",X"33",X"C9",X"3A",X"0C",
		X"62",X"D6",X"0E",X"BA",X"D2",X"1B",X"2A",X"3A",X"10",X"62",X"A7",X"3A",X"03",X"62",X"CA",X"08",
		X"2A",X"F6",X"07",X"D6",X"04",X"C3",X"0E",X"2A",X"D6",X"08",X"F6",X"07",X"C6",X"04",X"32",X"03",
		X"62",X"32",X"4C",X"69",X"3E",X"01",X"06",X"00",X"33",X"33",X"C9",X"AF",X"32",X"00",X"62",X"C9",
		X"47",X"C9",X"06",X"04",X"C3",X"77",X"4A",X"CD",X"DC",X"17",X"00",X"CD",X"13",X"29",X"C9",X"DD",
		X"7E",X"03",X"67",X"DD",X"7E",X"05",X"C6",X"04",X"6F",X"E5",X"CD",X"F0",X"2F",X"D1",X"7E",X"FE",
		X"B0",X"DA",X"7B",X"2A",X"E6",X"0F",X"FE",X"08",X"D2",X"7B",X"2A",X"7E",X"FE",X"C0",X"CA",X"7B",
		X"2A",X"DA",X"69",X"2A",X"FE",X"D0",X"DA",X"6E",X"2A",X"FE",X"E0",X"DA",X"63",X"2A",X"FE",X"F0",
		X"DA",X"6E",X"2A",X"E6",X"0F",X"3D",X"C3",X"72",X"2A",X"3E",X"FF",X"C3",X"72",X"2A",X"E6",X"0F",
		X"D6",X"09",X"4F",X"7B",X"E6",X"F8",X"81",X"BB",X"DA",X"7D",X"2A",X"AF",X"C9",X"D6",X"04",X"DD",
		X"77",X"05",X"3E",X"01",X"C9",X"C3",X"64",X"58",X"A7",X"C0",X"3A",X"16",X"62",X"A7",X"C0",X"C3",
		X"95",X"49",X"FE",X"01",X"C8",X"3A",X"03",X"62",X"D6",X"03",X"67",X"3A",X"05",X"62",X"C6",X"08",
		X"6F",X"E5",X"CD",X"F0",X"2F",X"D1",X"7E",X"FE",X"D0",X"C3",X"68",X"16",X"3E",X"00",X"32",X"21",
		X"62",X"C3",X"8B",X"4A",X"7A",X"E6",X"07",X"CA",X"CD",X"2A",X"01",X"20",X"00",X"ED",X"42",X"7E",
		X"FE",X"D0",X"DA",X"CD",X"2A",X"3E",X"00",X"32",X"21",X"62",X"C9",X"00",X"00",X"3E",X"01",X"32",
		X"21",X"62",X"C9",X"C3",X"0F",X"4A",X"47",X"3A",X"05",X"62",X"FE",X"90",X"CA",X"EA",X"2A",X"FE",
		X"C0",X"CA",X"F6",X"2A",X"FE",X"D4",X"CA",X"F0",X"2A",X"C9",X"3A",X"A3",X"63",X"C3",X"02",X"2B",
		X"3A",X"A6",X"63",X"C3",X"02",X"2B",X"78",X"FE",X"80",X"3A",X"A5",X"63",X"D2",X"02",X"2B",X"3A",
		X"A4",X"63",X"80",X"32",X"03",X"62",X"CD",X"9C",X"40",X"CD",X"1F",X"24",X"21",X"03",X"62",X"1D",
		X"CA",X"18",X"2B",X"15",X"CA",X"1A",X"2B",X"C9",X"35",X"C9",X"34",X"C9",X"C3",X"2E",X"4E",X"62",
		X"CD",X"29",X"2B",X"CD",X"AF",X"29",X"AF",X"47",X"C9",X"3A",X"27",X"62",X"A7",X"C2",X"53",X"2B",
		X"3A",X"03",X"62",X"67",X"3A",X"05",X"62",X"C6",X"07",X"6F",X"CD",X"9B",X"2B",X"A7",X"CA",X"51",
		X"2B",X"7B",X"91",X"FE",X"04",X"D2",X"74",X"2B",X"79",X"D6",X"07",X"32",X"05",X"62",X"3E",X"01",
		X"47",X"E1",X"C9",X"3A",X"03",X"62",X"D6",X"03",X"67",X"3A",X"05",X"62",X"C6",X"07",X"6F",X"CD",
		X"9B",X"2B",X"FE",X"02",X"CA",X"7A",X"2B",X"7A",X"C6",X"07",X"67",X"6B",X"CD",X"9B",X"2B",X"A7",
		X"C8",X"C3",X"7A",X"2B",X"3E",X"00",X"06",X"00",X"E1",X"C9",X"3A",X"10",X"62",X"A7",X"3A",X"03",
		X"62",X"CA",X"8B",X"2B",X"F6",X"07",X"D6",X"04",X"C3",X"91",X"2B",X"D6",X"08",X"F6",X"07",X"C6",
		X"04",X"32",X"03",X"62",X"32",X"4C",X"69",X"3E",X"01",X"E1",X"C9",X"E5",X"CD",X"F0",X"2F",X"D1",
		X"7E",X"FE",X"D0",X"DA",X"D9",X"2B",X"E6",X"0F",X"FE",X"08",X"C3",X"32",X"52",X"7E",X"FE",X"C0",
		X"CA",X"D9",X"2B",X"DA",X"DC",X"2B",X"FE",X"D0",X"DA",X"CB",X"2B",X"FE",X"E0",X"DA",X"C5",X"2B",
		X"FE",X"F0",X"DA",X"CB",X"2B",X"E6",X"0F",X"3D",X"C3",X"CF",X"2B",X"E6",X"0F",X"D6",X"09",X"4F",
		X"7B",X"E6",X"F8",X"81",X"4F",X"BB",X"DA",X"E1",X"2B",X"AF",X"47",X"C9",X"7B",X"E6",X"F8",X"3D",
		X"4F",X"3A",X"0C",X"62",X"DD",X"96",X"05",X"83",X"B9",X"CA",X"EF",X"2B",X"D2",X"F8",X"2B",X"79",
		X"D6",X"07",X"32",X"05",X"62",X"C3",X"FD",X"2B",X"3E",X"02",X"06",X"00",X"C9",X"3E",X"01",X"47",
		X"C3",X"93",X"4A",X"3E",X"0A",X"F7",X"D7",X"3A",X"93",X"63",X"0F",X"D8",X"3A",X"B1",X"62",X"A7",
		X"C8",X"4F",X"3A",X"B0",X"62",X"D6",X"02",X"B9",X"DA",X"7B",X"2C",X"3A",X"82",X"63",X"CB",X"4F",
		X"C2",X"86",X"2C",X"3A",X"80",X"63",X"47",X"3A",X"1A",X"60",X"E6",X"1F",X"B8",X"CA",X"33",X"2C",
		X"10",X"FA",X"C9",X"3A",X"B0",X"62",X"CB",X"3F",X"B9",X"DA",X"41",X"2C",X"3A",X"19",X"60",X"0F",
		X"D0",X"CD",X"57",X"00",X"E6",X"0F",X"C2",X"86",X"2C",X"3E",X"01",X"32",X"82",X"63",X"3C",X"32",
		X"8F",X"63",X"3E",X"01",X"32",X"92",X"63",X"3A",X"B2",X"62",X"B9",X"C0",X"D6",X"08",X"32",X"B2",
		X"62",X"11",X"20",X"00",X"21",X"00",X"64",X"06",X"05",X"7E",X"A7",X"CA",X"72",X"2C",X"19",X"10",
		X"F8",X"C9",X"3A",X"82",X"63",X"F6",X"80",X"32",X"82",X"63",X"C9",X"C6",X"02",X"B9",X"CA",X"49",
		X"2C",X"3E",X"02",X"C3",X"4B",X"2C",X"AF",X"32",X"82",X"63",X"3E",X"03",X"C3",X"4F",X"2C",X"3E",
		X"0A",X"F7",X"D7",X"3A",X"93",X"63",X"0F",X"DA",X"15",X"2D",X"3A",X"92",X"63",X"0F",X"D0",X"DD",
		X"21",X"00",X"67",X"CD",X"33",X"11",X"00",X"00",X"DD",X"7E",X"00",X"0F",X"DA",X"B3",X"2C",X"0F",
		X"D2",X"B8",X"2C",X"DD",X"19",X"10",X"F1",X"C9",X"DD",X"22",X"AA",X"62",X"CD",X"E1",X"47",X"00",
		X"CD",X"41",X"11",X"00",X"90",X"87",X"87",X"5F",X"21",X"80",X"69",X"19",X"22",X"AC",X"62",X"3E",
		X"01",X"32",X"93",X"63",X"11",X"01",X"05",X"CD",X"9F",X"30",X"21",X"B1",X"62",X"35",X"C2",X"E6",
		X"2C",X"3E",X"01",X"32",X"86",X"63",X"7E",X"FE",X"04",X"D2",X"F6",X"2C",X"21",X"A8",X"69",X"87",
		X"87",X"5F",X"16",X"00",X"19",X"72",X"C3",X"08",X"52",X"00",X"DD",X"36",X"08",X"0D",X"DD",X"36",
		X"15",X"00",X"3A",X"82",X"63",X"07",X"D2",X"15",X"2D",X"CD",X"29",X"52",X"00",X"DD",X"36",X"08",
		X"0D",X"DD",X"36",X"15",X"01",X"21",X"AF",X"62",X"35",X"C0",X"36",X"18",X"3A",X"8F",X"63",X"A7",
		X"CA",X"51",X"2D",X"4F",X"21",X"32",X"39",X"3A",X"82",X"63",X"0F",X"DA",X"2F",X"2D",X"0D",X"79",
		X"87",X"87",X"87",X"4F",X"87",X"87",X"81",X"5F",X"16",X"00",X"19",X"CD",X"4E",X"00",X"21",X"8F",
		X"63",X"35",X"C2",X"51",X"2D",X"3E",X"01",X"32",X"AF",X"62",X"3A",X"82",X"63",X"0F",X"DA",X"83",
		X"2D",X"2A",X"A8",X"62",X"7E",X"DD",X"2A",X"AA",X"62",X"ED",X"5B",X"AC",X"62",X"FE",X"7F",X"C3",
		X"F6",X"56",X"79",X"CD",X"F1",X"18",X"C3",X"F8",X"51",X"CB",X"79",X"CA",X"70",X"2D",X"EE",X"03",
		X"13",X"12",X"DD",X"77",X"07",X"DD",X"7E",X"08",X"13",X"12",X"23",X"C3",X"D1",X"51",X"23",X"22",
		X"A8",X"62",X"C9",X"21",X"C3",X"39",X"22",X"A8",X"62",X"C3",X"54",X"2D",X"21",X"C3",X"39",X"22",
		X"A8",X"62",X"DD",X"36",X"01",X"01",X"3A",X"82",X"63",X"0F",X"00",X"00",X"00",X"DD",X"36",X"01",
		X"00",X"DD",X"36",X"02",X"02",X"CD",X"03",X"40",X"00",X"DD",X"36",X"0F",X"01",X"AF",X"DD",X"77",
		X"10",X"DD",X"77",X"11",X"DD",X"77",X"12",X"DD",X"77",X"13",X"DD",X"77",X"14",X"32",X"93",X"63",
		X"32",X"92",X"63",X"1A",X"DD",X"77",X"03",X"13",X"13",X"13",X"1A",X"DD",X"77",X"05",X"21",X"5C",
		X"38",X"CD",X"4E",X"00",X"21",X"0B",X"69",X"0E",X"00",X"FF",X"C9",X"3E",X"07",X"F7",X"D7",X"3A",
		X"80",X"63",X"3C",X"A7",X"1F",X"47",X"3A",X"27",X"62",X"FE",X"02",X"20",X"01",X"04",X"3E",X"FE",
		X"37",X"1F",X"A7",X"10",X"FC",X"47",X"3A",X"1A",X"60",X"A0",X"C0",X"3E",X"01",X"32",X"9A",X"63",
		X"C3",X"4A",X"49",X"C9",X"C3",X"41",X"4D",X"D7",X"DD",X"21",X"00",X"65",X"CD",X"62",X"1E",X"00",
		X"00",X"00",X"DD",X"7E",X"00",X"0F",X"D2",X"54",X"2E",X"3A",X"1A",X"60",X"E6",X"0F",X"C2",X"29",
		X"2E",X"C3",X"09",X"4D",X"EE",X"07",X"FD",X"77",X"01",X"DD",X"7E",X"0D",X"C3",X"B0",X"4B",X"00",
		X"00",X"00",X"00",X"00",X"DD",X"34",X"03",X"DD",X"6E",X"0E",X"DD",X"66",X"0F",X"7E",X"4F",X"FE",
		X"7F",X"CA",X"A1",X"2E",X"23",X"DD",X"86",X"05",X"DD",X"77",X"05",X"DD",X"75",X"0E",X"DD",X"74",
		X"0F",X"C3",X"A9",X"1A",X"DD",X"36",X"01",X"00",X"FD",X"36",X"14",X"00",X"C3",X"A7",X"2E",X"CD",
		X"27",X"4D",X"00",X"00",X"00",X"00",X"00",X"CD",X"24",X"11",X"00",X"00",X"DD",X"7E",X"03",X"FD",
		X"77",X"00",X"DD",X"7E",X"05",X"CD",X"CC",X"52",X"11",X"10",X"00",X"DD",X"19",X"1E",X"04",X"FD",
		X"19",X"10",X"8F",X"C9",X"F5",X"AF",X"32",X"8C",X"60",X"F1",X"C3",X"DA",X"0B",X"32",X"00",X"7C",
		X"32",X"81",X"7C",X"C9",X"00",X"00",X"3E",X"01",X"DD",X"86",X"05",X"DD",X"77",X"05",X"C3",X"6C",
		X"2E",X"21",X"AA",X"39",X"C3",X"4B",X"2E",X"3A",X"96",X"63",X"0F",X"D2",X"78",X"2E",X"AF",X"32",
		X"96",X"63",X"DD",X"36",X"05",X"43",X"DD",X"36",X"0D",X"01",X"3E",X"4C",X"DD",X"77",X"03",X"CD",
		X"96",X"1A",X"00",X"00",X"CD",X"09",X"59",X"00",X"21",X"AA",X"39",X"DD",X"75",X"0E",X"DD",X"74",
		X"0F",X"C3",X"78",X"2E",X"3E",X"0F",X"F7",X"00",X"3A",X"94",X"6A",X"A7",X"C8",X"2A",X"97",X"6A",
		X"E5",X"DD",X"E1",X"CD",X"00",X"2F",X"2A",X"95",X"6A",X"77",X"7E",X"FE",X"F0",X"D8",X"2D",X"2D",
		X"2D",X"AF",X"77",X"32",X"94",X"6A",X"DD",X"77",X"03",X"32",X"9C",X"6A",X"32",X"2C",X"6A",X"C9",
		X"DD",X"34",X"05",X"DD",X"34",X"05",X"DD",X"7E",X"05",X"C9",X"00",X"00",X"00",X"00",X"1E",X"3A",
		X"07",X"62",X"CB",X"27",X"D2",X"1B",X"2F",X"F6",X"80",X"CB",X"F8",X"F6",X"08",X"4F",X"3A",X"94",
		X"63",X"CB",X"5F",X"CA",X"43",X"2F",X"CB",X"C0",X"CB",X"C1",X"DD",X"36",X"09",X"05",X"DD",X"36",
		X"0A",X"06",X"DD",X"36",X"0F",X"00",X"DD",X"36",X"0E",X"F0",X"CB",X"79",X"CA",X"43",X"2F",X"DD",
		X"36",X"0E",X"10",X"79",X"32",X"4D",X"69",X"0E",X"07",X"21",X"94",X"63",X"34",X"C2",X"B7",X"2F",
		X"21",X"95",X"63",X"34",X"7E",X"FE",X"02",X"C2",X"BE",X"2F",X"AF",X"32",X"95",X"63",X"32",X"17",
		X"62",X"DD",X"77",X"01",X"3A",X"03",X"62",X"ED",X"44",X"DD",X"77",X"0E",X"3A",X"07",X"62",X"32",
		X"4D",X"69",X"DD",X"36",X"00",X"00",X"3A",X"89",X"63",X"32",X"89",X"60",X"EB",X"3A",X"03",X"62",
		X"DD",X"86",X"0E",X"77",X"DD",X"77",X"03",X"23",X"70",X"23",X"71",X"23",X"3A",X"05",X"62",X"DD",
		X"86",X"0F",X"77",X"DD",X"77",X"05",X"C9",X"3A",X"18",X"62",X"0F",X"D0",X"DD",X"36",X"09",X"06",
		X"DD",X"36",X"0A",X"03",X"3A",X"07",X"62",X"07",X"3E",X"3C",X"1F",X"47",X"0E",X"07",X"3A",X"89",
		X"60",X"32",X"89",X"63",X"C3",X"7C",X"2F",X"3A",X"95",X"63",X"A7",X"CA",X"7C",X"2F",X"3A",X"1A",
		X"60",X"CB",X"5F",X"CA",X"7C",X"2F",X"0E",X"01",X"C3",X"7C",X"2F",X"3E",X"05",X"F7",X"C3",X"9E",
		X"57",X"00",X"00",X"3E",X"03",X"32",X"B9",X"62",X"32",X"96",X"63",X"11",X"01",X"05",X"CD",X"9F",
		X"30",X"3A",X"B3",X"62",X"77",X"21",X"B1",X"62",X"35",X"C0",X"3E",X"01",X"32",X"86",X"63",X"C9",
		X"7D",X"0F",X"0F",X"0F",X"E6",X"1F",X"6F",X"7C",X"2F",X"E6",X"F8",X"5F",X"AF",X"67",X"CB",X"13",
		X"17",X"CB",X"13",X"17",X"C6",X"74",X"57",X"19",X"C9",X"57",X"0F",X"DA",X"22",X"30",X"0E",X"93",
		X"0F",X"0F",X"D2",X"17",X"30",X"0E",X"6C",X"07",X"DA",X"31",X"30",X"79",X"E6",X"F0",X"4F",X"C3",
		X"31",X"30",X"0E",X"B4",X"0F",X"0F",X"D2",X"2B",X"30",X"0E",X"1E",X"CB",X"50",X"CA",X"31",X"30",
		X"05",X"79",X"0F",X"0F",X"4F",X"E6",X"03",X"B8",X"C2",X"31",X"30",X"79",X"0F",X"0F",X"E6",X"03",
		X"FE",X"03",X"C0",X"CB",X"92",X"15",X"C0",X"3E",X"04",X"C9",X"11",X"C0",X"FF",X"3A",X"8E",X"63",
		X"4F",X"06",X"00",X"21",X"58",X"76",X"CD",X"64",X"30",X"21",X"B8",X"75",X"CD",X"64",X"30",X"21",
		X"8E",X"63",X"35",X"C9",X"09",X"7E",X"19",X"77",X"C9",X"DF",X"2A",X"C0",X"63",X"34",X"C9",X"21",
		X"AF",X"62",X"34",X"7E",X"E6",X"07",X"00",X"21",X"0B",X"69",X"0E",X"FC",X"FF",X"0E",X"81",X"21",
		X"09",X"69",X"CD",X"96",X"30",X"21",X"1D",X"69",X"CD",X"96",X"30",X"CD",X"57",X"00",X"E6",X"80",
		X"21",X"2D",X"69",X"AE",X"77",X"C9",X"06",X"02",X"79",X"AE",X"77",X"19",X"10",X"FA",X"C9",X"E5",
		X"21",X"C0",X"60",X"3A",X"B0",X"60",X"6F",X"CB",X"7E",X"CA",X"BB",X"30",X"72",X"2C",X"73",X"2C",
		X"7D",X"FE",X"C0",X"D2",X"B8",X"30",X"3E",X"C0",X"32",X"B0",X"60",X"E1",X"C9",X"21",X"50",X"69",
		X"06",X"01",X"CD",X"E4",X"30",X"2E",X"80",X"06",X"0A",X"CD",X"E4",X"30",X"2E",X"B8",X"06",X"0B",
		X"CD",X"E4",X"30",X"21",X"0C",X"6A",X"06",X"05",X"C3",X"E4",X"30",X"21",X"4C",X"69",X"36",X"00",
		X"2E",X"58",X"06",X"06",X"7D",X"36",X"00",X"C6",X"04",X"6F",X"10",X"F9",X"C9",X"CD",X"FA",X"30",
		X"CD",X"3C",X"31",X"CD",X"B1",X"31",X"CD",X"F3",X"34",X"C9",X"3A",X"80",X"63",X"FE",X"06",X"38",
		X"02",X"3E",X"05",X"EF",X"10",X"31",X"10",X"31",X"1B",X"31",X"26",X"31",X"26",X"31",X"31",X"31",
		X"3A",X"1A",X"60",X"E6",X"01",X"FE",X"01",X"C8",X"33",X"33",X"C9",X"3A",X"1A",X"60",X"E6",X"07",
		X"FE",X"05",X"F8",X"33",X"33",X"C9",X"3A",X"1A",X"60",X"E6",X"03",X"FE",X"03",X"F8",X"33",X"33",
		X"C9",X"3A",X"1A",X"60",X"E6",X"07",X"FE",X"07",X"F8",X"33",X"33",X"C9",X"DD",X"21",X"00",X"64",
		X"AF",X"32",X"A1",X"63",X"06",X"05",X"11",X"20",X"00",X"DD",X"7E",X"00",X"FE",X"00",X"CA",X"7C",
		X"31",X"3A",X"A1",X"63",X"3C",X"32",X"A1",X"63",X"3E",X"81",X"00",X"00",X"00",X"3A",X"17",X"62",
		X"FE",X"01",X"C2",X"6A",X"31",X"3E",X"00",X"DD",X"77",X"08",X"DD",X"19",X"10",X"DB",X"21",X"A0",
		X"63",X"36",X"00",X"3A",X"A1",X"63",X"FE",X"00",X"C0",X"33",X"33",X"C9",X"C3",X"AF",X"5B",X"00",
		X"00",X"CA",X"6A",X"31",X"3A",X"27",X"62",X"FE",X"02",X"C2",X"95",X"31",X"3A",X"A1",X"63",X"4F",
		X"3A",X"80",X"63",X"B9",X"C8",X"3A",X"A0",X"63",X"FE",X"01",X"C2",X"6A",X"31",X"C3",X"CE",X"56",
		X"DD",X"77",X"18",X"AF",X"32",X"A0",X"63",X"3A",X"A1",X"63",X"3C",X"32",X"A1",X"63",X"C3",X"6A",
		X"31",X"CD",X"DD",X"31",X"AF",X"32",X"A2",X"63",X"21",X"E0",X"63",X"22",X"C8",X"63",X"2A",X"C8",
		X"63",X"01",X"20",X"00",X"09",X"22",X"C8",X"63",X"7E",X"A7",X"CA",X"D0",X"31",X"CD",X"02",X"32",
		X"3A",X"A2",X"63",X"3C",X"32",X"A2",X"63",X"FE",X"05",X"C2",X"BE",X"31",X"C9",X"3A",X"80",X"63",
		X"FE",X"03",X"F8",X"CD",X"F6",X"31",X"FE",X"01",X"C0",X"21",X"39",X"64",X"3E",X"02",X"77",X"21",
		X"79",X"64",X"3E",X"02",X"77",X"C9",X"3A",X"18",X"60",X"E6",X"03",X"FE",X"01",X"C0",X"3A",X"1A",
		X"60",X"C9",X"DD",X"2A",X"C8",X"63",X"DD",X"7E",X"18",X"FE",X"01",X"CA",X"7A",X"32",X"DD",X"7E",
		X"0D",X"FE",X"04",X"F2",X"30",X"32",X"DD",X"7E",X"19",X"FE",X"02",X"CA",X"7E",X"32",X"CD",X"0F",
		X"33",X"3A",X"18",X"60",X"E6",X"02",X"C2",X"33",X"32",X"DD",X"7E",X"0D",X"A7",X"CA",X"57",X"32",
		X"CD",X"3D",X"33",X"DD",X"7E",X"0D",X"FE",X"04",X"F2",X"91",X"32",X"CD",X"AD",X"33",X"CD",X"8C",
		X"29",X"FE",X"01",X"CA",X"97",X"32",X"DD",X"2A",X"C8",X"63",X"DD",X"7E",X"0E",X"FE",X"10",X"DA",
		X"8C",X"32",X"FE",X"F0",X"D2",X"84",X"32",X"DD",X"7E",X"13",X"FE",X"00",X"C2",X"B9",X"32",X"3E",
		X"11",X"DD",X"77",X"13",X"16",X"00",X"5F",X"21",X"7A",X"3A",X"19",X"7E",X"DD",X"46",X"0E",X"DD",
		X"70",X"03",X"DD",X"4E",X"0F",X"81",X"DD",X"77",X"05",X"C9",X"CD",X"BD",X"32",X"C9",X"CD",X"D6",
		X"32",X"C3",X"29",X"32",X"3E",X"02",X"DD",X"77",X"0D",X"C3",X"57",X"32",X"3E",X"01",X"C3",X"86",
		X"32",X"CD",X"E7",X"33",X"C3",X"57",X"32",X"DD",X"2A",X"C8",X"63",X"DD",X"7E",X"0D",X"FE",X"01",
		X"C2",X"B1",X"32",X"3E",X"02",X"DD",X"35",X"0E",X"DD",X"77",X"0D",X"CD",X"C3",X"33",X"C3",X"57",
		X"32",X"3E",X"01",X"DD",X"34",X"0E",X"C3",X"A8",X"32",X"3D",X"C3",X"61",X"32",X"3A",X"27",X"62",
		X"FE",X"03",X"CA",X"CE",X"32",X"FE",X"02",X"CA",X"D2",X"32",X"CD",X"B9",X"34",X"C9",X"CD",X"2C",
		X"34",X"C9",X"CD",X"78",X"34",X"C9",X"DD",X"7E",X"1C",X"FE",X"00",X"C2",X"FD",X"32",X"DD",X"7E",
		X"1D",X"FE",X"01",X"C2",X"0B",X"33",X"DD",X"36",X"1D",X"00",X"3A",X"05",X"62",X"DD",X"46",X"0F",
		X"90",X"DA",X"03",X"33",X"DD",X"36",X"1C",X"FF",X"CD",X"30",X"47",X"00",X"C9",X"DD",X"35",X"1C",
		X"00",X"00",X"00",X"DD",X"36",X"19",X"00",X"DD",X"36",X"1C",X"00",X"CD",X"0F",X"33",X"C9",X"DD",
		X"7E",X"16",X"FE",X"00",X"C2",X"32",X"33",X"DD",X"36",X"16",X"4B",X"CD",X"30",X"47",X"00",X"3A",
		X"18",X"60",X"0F",X"D2",X"32",X"33",X"DD",X"7E",X"0D",X"FE",X"01",X"CA",X"36",X"33",X"CD",X"28",
		X"47",X"00",X"DD",X"35",X"16",X"C9",X"DD",X"36",X"0D",X"02",X"C3",X"32",X"33",X"DD",X"7E",X"0D",
		X"FE",X"08",X"CA",X"71",X"33",X"FE",X"04",X"CA",X"8A",X"33",X"CD",X"A1",X"33",X"DD",X"7E",X"0F",
		X"C6",X"08",X"57",X"DD",X"7E",X"0E",X"01",X"15",X"00",X"C3",X"AF",X"5D",X"A7",X"CA",X"99",X"33",
		X"DD",X"70",X"1F",X"3A",X"05",X"62",X"47",X"DD",X"7E",X"0F",X"90",X"00",X"C3",X"76",X"47",X"04",
		X"C9",X"DD",X"7E",X"0F",X"C6",X"08",X"DD",X"46",X"1F",X"B8",X"C0",X"CD",X"30",X"47",X"00",X"DD",
		X"7E",X"19",X"FE",X"02",X"C0",X"C3",X"28",X"47",X"00",X"C9",X"DD",X"7E",X"0F",X"C6",X"08",X"DD",
		X"46",X"1F",X"B8",X"C0",X"CD",X"30",X"47",X"00",X"C9",X"DD",X"70",X"1F",X"C3",X"66",X"47",X"00",
		X"C9",X"3E",X"07",X"F7",X"DD",X"7E",X"0F",X"FE",X"10",X"D0",X"33",X"33",X"C9",X"DD",X"7E",X"0D",
		X"FE",X"01",X"CA",X"D9",X"33",X"DD",X"7E",X"07",X"E6",X"7F",X"DD",X"77",X"07",X"DD",X"35",X"0E",
		X"CD",X"09",X"34",X"3A",X"27",X"62",X"FE",X"01",X"C0",X"DD",X"66",X"0E",X"DD",X"6E",X"0F",X"DD",
		X"46",X"0D",X"CD",X"33",X"23",X"DD",X"75",X"0F",X"C9",X"DD",X"7E",X"07",X"F6",X"80",X"DD",X"77",
		X"07",X"DD",X"34",X"0E",X"C3",X"C0",X"33",X"CD",X"09",X"34",X"DD",X"7E",X"0D",X"FE",X"08",X"C2",
		X"05",X"34",X"DD",X"7E",X"14",X"A7",X"C2",X"01",X"34",X"DD",X"36",X"14",X"02",X"DD",X"35",X"0F",
		X"C9",X"DD",X"35",X"14",X"C9",X"DD",X"34",X"0F",X"C9",X"DD",X"7E",X"15",X"A7",X"C2",X"28",X"34",
		X"DD",X"36",X"15",X"02",X"DD",X"34",X"07",X"DD",X"7E",X"07",X"E6",X"0F",X"FE",X"0F",X"C0",X"DD",
		X"7E",X"07",X"EE",X"02",X"DD",X"77",X"07",X"C9",X"DD",X"35",X"15",X"C9",X"DD",X"6E",X"1A",X"DD",
		X"66",X"1B",X"AF",X"01",X"00",X"00",X"ED",X"4A",X"C2",X"42",X"34",X"21",X"8C",X"3A",X"DD",X"36",
		X"03",X"40",X"DD",X"34",X"03",X"CD",X"8E",X"40",X"CA",X"56",X"34",X"DD",X"77",X"05",X"23",X"DD",
		X"75",X"1A",X"DD",X"74",X"1B",X"C9",X"AF",X"DD",X"77",X"13",X"DD",X"77",X"18",X"DD",X"77",X"0D",
		X"DD",X"77",X"1C",X"DD",X"7E",X"03",X"DD",X"77",X"0E",X"DD",X"7E",X"05",X"DD",X"77",X"0F",X"DD",
		X"36",X"1A",X"00",X"DD",X"36",X"1B",X"00",X"C9",X"DD",X"6E",X"1A",X"DD",X"66",X"1B",X"AF",X"01",
		X"00",X"00",X"ED",X"4A",X"C2",X"9A",X"34",X"21",X"AC",X"3A",X"3A",X"03",X"62",X"CB",X"7F",X"CA",
		X"A8",X"34",X"DD",X"36",X"0D",X"01",X"DD",X"36",X"03",X"4C",X"DD",X"7E",X"0D",X"FE",X"01",X"C2",
		X"B3",X"34",X"DD",X"34",X"03",X"C3",X"45",X"34",X"DD",X"36",X"0D",X"02",X"DD",X"36",X"03",X"48",
		X"C3",X"9A",X"34",X"DD",X"35",X"03",X"C3",X"45",X"34",X"3A",X"27",X"62",X"FE",X"04",X"C8",X"3A",
		X"03",X"62",X"CB",X"7F",X"C2",X"ED",X"34",X"21",X"C4",X"3A",X"06",X"00",X"3A",X"19",X"60",X"E6",
		X"06",X"4F",X"09",X"7E",X"DD",X"77",X"03",X"DD",X"77",X"0E",X"23",X"7E",X"DD",X"77",X"05",X"DD",
		X"77",X"0F",X"AF",X"DD",X"77",X"0D",X"DD",X"77",X"18",X"DD",X"77",X"1C",X"C9",X"21",X"D4",X"3A",
		X"C3",X"CA",X"34",X"21",X"00",X"64",X"11",X"D0",X"69",X"06",X"05",X"7E",X"A7",X"CA",X"1E",X"35",
		X"2C",X"2C",X"2C",X"7E",X"12",X"3E",X"04",X"85",X"6F",X"1C",X"7E",X"12",X"2C",X"1C",X"7E",X"12",
		X"2D",X"2D",X"2D",X"1C",X"7E",X"12",X"13",X"3E",X"1B",X"85",X"6F",X"10",X"DE",X"C9",X"3E",X"05",
		X"85",X"6F",X"3E",X"04",X"83",X"5F",X"C3",X"17",X"35",X"00",X"00",X"00",X"00",X"01",X"00",X"00",
		X"02",X"00",X"00",X"03",X"00",X"00",X"04",X"00",X"00",X"05",X"00",X"00",X"06",X"00",X"00",X"07",
		X"00",X"00",X"08",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"20",X"00",
		X"00",X"30",X"00",X"00",X"40",X"00",X"00",X"50",X"00",X"00",X"60",X"00",X"00",X"70",X"00",X"00",
		X"80",X"00",X"00",X"90",X"00",X"94",X"77",X"01",X"23",X"24",X"10",X"10",X"00",X"01",X"01",X"08",
		X"00",X"00",X"10",X"10",X"18",X"19",X"22",X"1F",X"23",X"18",X"19",X"10",X"23",X"2B",X"10",X"10",
		X"3F",X"00",X"00",X"18",X"01",X"F4",X"76",X"96",X"77",X"02",X"1E",X"14",X"10",X"10",X"00",X"00",
		X"09",X"05",X"00",X"00",X"10",X"10",X"1D",X"2B",X"10",X"29",X"1F",X"23",X"18",X"19",X"14",X"11",
		X"10",X"10",X"3F",X"00",X"00",X"95",X"00",X"F6",X"76",X"98",X"77",X"03",X"22",X"14",X"10",X"10",
		X"00",X"00",X"08",X"03",X"00",X"00",X"10",X"10",X"18",X"2B",X"10",X"29",X"11",X"1D",X"11",X"23",
		X"18",X"19",X"24",X"11",X"3F",X"00",X"00",X"83",X"00",X"F8",X"76",X"9A",X"77",X"04",X"24",X"18",
		X"10",X"10",X"00",X"00",X"06",X"02",X"00",X"00",X"10",X"10",X"18",X"19",X"23",X"11",X"1D",X"19",
		X"10",X"23",X"2B",X"10",X"10",X"10",X"3F",X"00",X"00",X"62",X"00",X"FA",X"76",X"9C",X"77",X"05",
		X"24",X"18",X"10",X"10",X"00",X"00",X"05",X"07",X"00",X"00",X"10",X"10",X"29",X"25",X"1B",X"1F",
		X"10",X"23",X"2B",X"10",X"10",X"10",X"10",X"10",X"3F",X"00",X"00",X"57",X"00",X"FC",X"76",X"3B",
		X"5C",X"4B",X"5C",X"5B",X"5C",X"6B",X"5C",X"7B",X"5C",X"8B",X"5C",X"9B",X"5C",X"AB",X"5C",X"BB",
		X"5C",X"CB",X"5C",X"3B",X"6C",X"4B",X"6C",X"5B",X"6C",X"6B",X"6C",X"7B",X"6C",X"8B",X"6C",X"9B",
		X"6C",X"AB",X"6C",X"BB",X"6C",X"CB",X"6C",X"3B",X"7C",X"4B",X"7C",X"5B",X"7C",X"6B",X"7C",X"7B",
		X"7C",X"8B",X"7C",X"9B",X"7C",X"AB",X"7C",X"BB",X"7C",X"CB",X"7C",X"8B",X"36",X"01",X"00",X"98",
		X"36",X"A5",X"36",X"B2",X"36",X"BF",X"36",X"06",X"00",X"CC",X"36",X"08",X"00",X"E6",X"36",X"FD",
		X"36",X"0B",X"00",X"15",X"37",X"1C",X"37",X"30",X"37",X"38",X"37",X"47",X"37",X"5D",X"37",X"73",
		X"37",X"8B",X"37",X"00",X"61",X"22",X"61",X"44",X"61",X"66",X"61",X"88",X"61",X"9E",X"37",X"B6",
		X"37",X"D2",X"37",X"E1",X"37",X"1D",X"00",X"F4",X"37",X"06",X"38",X"96",X"76",X"17",X"11",X"1D",
		X"15",X"10",X"10",X"1F",X"26",X"15",X"22",X"3F",X"94",X"76",X"20",X"1C",X"11",X"29",X"15",X"22",
		X"10",X"30",X"32",X"31",X"3F",X"94",X"76",X"20",X"1C",X"11",X"29",X"15",X"22",X"10",X"30",X"33",
		X"31",X"3F",X"80",X"76",X"18",X"19",X"17",X"18",X"10",X"23",X"13",X"1F",X"22",X"15",X"3F",X"9F",
		X"75",X"13",X"22",X"15",X"14",X"19",X"24",X"10",X"10",X"10",X"10",X"3F",X"5E",X"77",X"18",X"1F",
		X"27",X"10",X"18",X"19",X"17",X"18",X"10",X"13",X"11",X"1E",X"10",X"29",X"1F",X"25",X"10",X"17",
		X"15",X"24",X"10",X"FB",X"10",X"3F",X"29",X"77",X"1F",X"1E",X"1C",X"29",X"10",X"01",X"10",X"20",
		X"1C",X"11",X"29",X"15",X"22",X"10",X"12",X"25",X"24",X"24",X"1F",X"1E",X"3F",X"29",X"77",X"01",
		X"10",X"1F",X"22",X"10",X"02",X"10",X"20",X"1C",X"11",X"29",X"15",X"22",X"23",X"10",X"12",X"25",
		X"24",X"24",X"1F",X"1E",X"3F",X"27",X"76",X"20",X"25",X"23",X"18",X"3F",X"06",X"77",X"1E",X"11",
		X"1D",X"15",X"10",X"22",X"15",X"17",X"19",X"23",X"24",X"22",X"11",X"24",X"19",X"1F",X"1E",X"3F",
		X"88",X"76",X"1E",X"11",X"1D",X"15",X"2E",X"3F",X"E9",X"75",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",
		X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"3F",X"0B",X"77",X"11",X"10",X"12",X"10",X"13",X"10",X"14",
		X"10",X"15",X"10",X"16",X"10",X"17",X"10",X"18",X"10",X"19",X"10",X"1A",X"3F",X"0D",X"77",X"1B",
		X"10",X"1C",X"10",X"1D",X"10",X"1E",X"10",X"1F",X"10",X"20",X"10",X"21",X"10",X"22",X"10",X"23",
		X"10",X"24",X"3F",X"0F",X"77",X"25",X"10",X"26",X"10",X"27",X"10",X"28",X"10",X"29",X"10",X"2A",
		X"10",X"2B",X"10",X"2C",X"44",X"45",X"46",X"47",X"48",X"10",X"3F",X"F2",X"76",X"22",X"15",X"17",
		X"19",X"10",X"24",X"19",X"1D",X"15",X"10",X"10",X"30",X"06",X"00",X"31",X"10",X"3F",X"92",X"77",
		X"22",X"11",X"1E",X"1B",X"10",X"10",X"23",X"13",X"1F",X"22",X"15",X"10",X"10",X"10",X"10",X"10",
		X"10",X"1E",X"11",X"1D",X"15",X"3F",X"72",X"77",X"29",X"1F",X"25",X"22",X"10",X"1E",X"11",X"1D",
		X"15",X"10",X"27",X"11",X"23",X"10",X"22",X"15",X"17",X"19",X"23",X"24",X"15",X"22",X"15",X"14",
		X"42",X"3F",X"A7",X"76",X"19",X"1E",X"23",X"15",X"22",X"24",X"10",X"13",X"1F",X"19",X"1E",X"10",
		X"3F",X"0A",X"77",X"10",X"10",X"20",X"1C",X"11",X"29",X"15",X"22",X"10",X"10",X"10",X"10",X"13",
		X"1F",X"19",X"1E",X"3F",X"BC",X"76",X"C0",X"C1",X"C2",X"C3",X"C4",X"C5",X"C6",X"C7",X"C8",X"C9",
		X"CA",X"CB",X"3F",X"CD",X"CE",X"CF",X"D0",X"D1",X"D2",X"D3",X"D4",X"D5",X"3F",X"00",X"00",X"00",
		X"6B",X"C8",X"01",X"93",X"18",X"93",X"C0",X"01",X"63",X"18",X"63",X"48",X"01",X"9B",X"18",X"9B",
		X"48",X"01",X"6B",X"18",X"6B",X"C0",X"0A",X"EF",X"F8",X"10",X"F8",X"08",X"CF",X"48",X"10",X"48",
		X"AA",X"21",X"8D",X"60",X"11",X"81",X"7C",X"7E",X"A7",X"28",X"03",X"35",X"3E",X"01",X"12",X"21",
		X"8B",X"60",X"C9",X"00",X"90",X"91",X"92",X"7C",X"01",X"93",X"8D",X"7D",X"8C",X"7C",X"00",X"6F",
		X"7C",X"00",X"6E",X"7C",X"00",X"6D",X"7C",X"00",X"6C",X"8F",X"7F",X"8E",X"36",X"24",X"09",X"3F",
		X"20",X"23",X"09",X"3F",X"2B",X"22",X"09",X"3F",X"2B",X"20",X"07",X"2F",X"3B",X"27",X"09",X"30",
		X"1B",X"28",X"09",X"30",X"3B",X"2E",X"08",X"2E",X"1B",X"2C",X"08",X"2E",X"3B",X"30",X"08",X"40",
		X"1B",X"2F",X"08",X"40",X"2B",X"2D",X"08",X"2E",X"2B",X"2D",X"88",X"40",X"36",X"24",X"09",X"3F",
		X"20",X"23",X"09",X"3F",X"2B",X"22",X"09",X"3F",X"2B",X"20",X"08",X"2F",X"3B",X"27",X"09",X"30",
		X"1B",X"28",X"09",X"30",X"3B",X"2E",X"01",X"2E",X"1B",X"2C",X"01",X"2E",X"3B",X"30",X"01",X"40",
		X"1B",X"2F",X"01",X"40",X"FD",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"01",X"01",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"FF",X"00",X"00",X"01",X"00",X"01",X"01",X"01",X"01",X"01",X"7F",X"04",X"7F",X"F0",X"10",
		X"F0",X"02",X"DF",X"F2",X"70",X"F8",X"02",X"6F",X"F8",X"10",X"F8",X"AA",X"04",X"DF",X"D0",X"90",
		X"D0",X"02",X"DF",X"DC",X"20",X"D1",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"04",X"DF",X"A8",X"20",
		X"A8",X"04",X"5F",X"B0",X"20",X"B0",X"02",X"DF",X"B0",X"20",X"BB",X"AA",X"04",X"DF",X"88",X"30",
		X"88",X"04",X"DF",X"90",X"B0",X"90",X"02",X"DF",X"9A",X"20",X"8F",X"AA",X"04",X"BF",X"68",X"20",
		X"68",X"04",X"3F",X"70",X"20",X"70",X"02",X"DF",X"6E",X"20",X"79",X"AA",X"02",X"DF",X"58",X"A0",
		X"55",X"AA",X"36",X"A3",X"09",X"3F",X"20",X"A4",X"09",X"3F",X"2B",X"22",X"09",X"3F",X"2B",X"21",
		X"07",X"2F",X"3B",X"27",X"09",X"30",X"1B",X"28",X"09",X"30",X"3B",X"2E",X"08",X"2E",X"1B",X"2C",
		X"08",X"2E",X"3B",X"AF",X"08",X"40",X"1B",X"B0",X"08",X"40",X"36",X"A3",X"09",X"3F",X"20",X"A4",
		X"09",X"3F",X"2B",X"22",X"09",X"3F",X"2B",X"A0",X"07",X"2F",X"3B",X"A8",X"09",X"30",X"1B",X"A7",
		X"09",X"30",X"3B",X"AC",X"08",X"2E",X"1B",X"AE",X"08",X"2E",X"3B",X"AF",X"08",X"40",X"1B",X"B0",
		X"08",X"40",X"36",X"24",X"09",X"3F",X"20",X"23",X"09",X"3F",X"2B",X"22",X"09",X"3F",X"2B",X"21",
		X"07",X"2F",X"3B",X"27",X"09",X"30",X"1B",X"28",X"09",X"30",X"3B",X"2E",X"08",X"2E",X"1B",X"2C",
		X"08",X"2E",X"3B",X"30",X"08",X"40",X"1B",X"2F",X"08",X"40",X"FF",X"FF",X"00",X"00",X"01",X"01",
		X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"58",X"40",X"58",X"40",X"58",X"40",X"58",X"40",X"7F",X"58",X"40",X"7F",X"8A",
		X"24",X"09",X"2F",X"74",X"23",X"09",X"2F",X"7F",X"22",X"09",X"2F",X"7F",X"A0",X"07",X"1F",X"8F",
		X"A8",X"09",X"20",X"6F",X"A7",X"09",X"20",X"8F",X"AC",X"08",X"1E",X"6F",X"AE",X"08",X"1E",X"8F",
		X"30",X"08",X"30",X"6F",X"2F",X"08",X"30",X"8A",X"A3",X"09",X"2F",X"74",X"A4",X"09",X"2F",X"7F",
		X"22",X"09",X"2F",X"7F",X"21",X"07",X"1F",X"8F",X"27",X"09",X"20",X"6F",X"28",X"09",X"20",X"8F",
		X"2E",X"08",X"1E",X"6F",X"2C",X"08",X"1E",X"8F",X"AF",X"08",X"30",X"6F",X"B0",X"08",X"30",X"8A",
		X"24",X"89",X"20",X"74",X"23",X"89",X"20",X"7F",X"22",X"89",X"20",X"7F",X"A0",X"87",X"30",X"8F",
		X"A8",X"89",X"2F",X"6F",X"A7",X"89",X"2F",X"00",X"70",X"88",X"68",X"00",X"A9",X"88",X"6C",X"00",
		X"70",X"88",X"68",X"00",X"70",X"8A",X"68",X"00",X"3A",X"27",X"62",X"FE",X"03",X"21",X"A2",X"11",
		X"C0",X"21",X"55",X"3A",X"C9",X"3B",X"0F",X"04",X"04",X"32",X"16",X"62",X"32",X"8C",X"6A",X"3D",
		X"32",X"98",X"63",X"C9",X"00",X"02",X"01",X"04",X"03",X"02",X"01",X"04",X"03",X"02",X"01",X"04",
		X"03",X"02",X"01",X"04",X"03",X"02",X"01",X"04",X"03",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"78",X"77",X"77",X"76",
		X"76",X"75",X"75",X"74",X"74",X"73",X"72",X"72",X"71",X"71",X"72",X"72",X"73",X"74",X"74",X"75",
		X"76",X"78",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"80",X"7B",X"78",X"76",
		X"74",X"73",X"72",X"71",X"70",X"70",X"6F",X"6F",X"6F",X"70",X"70",X"71",X"72",X"73",X"74",X"75",
		X"76",X"77",X"78",X"AA",X"EE",X"F0",X"0D",X"6B",X"E0",X"6B",X"FF",X"0D",X"74",X"E0",X"74",X"FF",
		X"0D",X"94",X"E8",X"94",X"FF",X"0D",X"B4",X"E0",X"B4",X"FF",X"0D",X"BB",X"E0",X"BB",X"FF",X"0D",
		X"DB",X"D8",X"DB",X"FF",X"0D",X"E4",X"D8",X"E4",X"FF",X"00",X"6B",X"18",X"6B",X"30",X"00",X"9B",
		X"18",X"9B",X"30",X"00",X"13",X"48",X"13",X"E0",X"00",X"2B",X"48",X"2B",X"D8",X"00",X"43",X"78",
		X"43",X"A8",X"00",X"43",X"A8",X"43",X"E0",X"00",X"6B",X"48",X"6B",X"C8",X"00",X"8B",X"48",X"8B",
		X"98",X"00",X"A3",X"50",X"A3",X"C8",X"00",X"BB",X"50",X"BB",X"B8",X"00",X"D3",X"30",X"D3",X"90",
		X"00",X"D3",X"90",X"D3",X"C8",X"00",X"EB",X"30",X"3B",X"90",X"00",X"EB",X"90",X"EB",X"C8",X"08",
		X"5F",X"28",X"48",X"28",X"08",X"97",X"48",X"10",X"48",X"08",X"CF",X"50",X"90",X"50",X"08",X"4F",
		X"78",X"30",X"78",X"08",X"5F",X"A8",X"30",X"A8",X"08",X"EF",X"90",X"C0",X"90",X"05",X"47",X"F0",
		X"00",X"F0",X"05",X"7F",X"E0",X"60",X"E0",X"05",X"9F",X"E8",X"88",X"E8",X"05",X"C7",X"E0",X"A8",
		X"E0",X"05",X"EF",X"D8",X"D0",X"D8",X"0A",X"EF",X"F8",X"10",X"F8",X"AA",X"48",X"74",X"AC",X"74",
		X"0C",X"75",X"12",X"75",X"6F",X"75",X"73",X"75",X"CD",X"75",X"D1",X"75",X"51",X"76",X"F7",X"76",
		X"51",X"77",X"AD",X"77",X"B4",X"77",X"0D",X"14",X"C0",X"14",X"FF",X"0D",X"1B",X"70",X"1B",X"FF",
		X"0D",X"24",X"C0",X"24",X"FF",X"0D",X"64",X"E8",X"64",X"FF",X"0D",X"6B",X"E8",X"6B",X"FF",X"0D",
		X"CB",X"E8",X"CB",X"FF",X"0D",X"D4",X"E8",X"D4",X"FF",X"0D",X"DB",X"A8",X"DB",X"FF",X"0D",X"E4",
		X"A8",X"E4",X"FF",X"0D",X"74",X"E8",X"74",X"FF",X"02",X"6B",X"18",X"6B",X"30",X"0D",X"EB",X"E8",
		X"EB",X"FF",X"02",X"9B",X"18",X"9B",X"30",X"02",X"13",X"48",X"13",X"68",X"02",X"2B",X"48",X"2B",
		X"B0",X"02",X"43",X"48",X"43",X"98",X"02",X"5B",X"48",X"5B",X"78",X"02",X"73",X"48",X"73",X"80",
		X"02",X"8B",X"48",X"8B",X"78",X"02",X"A3",X"48",X"A3",X"98",X"02",X"BB",X"48",X"BB",X"78",X"02",
		X"D3",X"38",X"D3",X"78",X"02",X"EB",X"38",X"EB",X"78",X"01",X"D3",X"B0",X"D3",X"D8",X"01",X"EB",
		X"B0",X"EB",X"D8",X"02",X"13",X"70",X"13",X"B0",X"08",X"5F",X"28",X"48",X"28",X"08",X"A7",X"48",
		X"10",X"48",X"08",X"CF",X"48",X"B8",X"48",X"05",X"CF",X"C0",X"B0",X"C0",X"05",X"27",X"70",X"10",
		X"70",X"05",X"37",X"C0",X"00",X"C0",X"05",X"2F",X"E8",X"00",X"E8",X"05",X"7F",X"E8",X"58",X"E8",
		X"0B",X"D8",X"98",X"38",X"98",X"05",X"FF",X"E8",X"C0",X"E8",X"05",X"EF",X"A8",X"D0",X"A8",X"AA",
		X"04",X"40",X"E4",X"40",X"FF",X"04",X"90",X"5C",X"90",X"87",X"04",X"60",X"5C",X"60",X"87",X"04",
		X"40",X"5C",X"40",X"87",X"04",X"B8",X"BC",X"B8",X"E7",X"04",X"B0",X"5C",X"B0",X"87",X"04",X"40",
		X"94",X"40",X"AF",X"03",X"6B",X"18",X"6B",X"30",X"03",X"D3",X"30",X"D3",X"87",X"03",X"EB",X"30",
		X"EB",X"87",X"03",X"13",X"58",X"13",X"AF",X"03",X"2B",X"58",X"2B",X"AF",X"03",X"D3",X"90",X"D3",
		X"D8",X"03",X"EB",X"90",X"EB",X"D8",X"03",X"13",X"B8",X"13",X"E8",X"03",X"2B",X"B8",X"2B",X"E8",
		X"06",X"5F",X"28",X"40",X"28",X"06",X"2F",X"48",X"10",X"48",X"07",X"2F",X"50",X"10",X"50",X"06",
		X"C7",X"48",X"38",X"48",X"07",X"C7",X"50",X"38",X"50",X"06",X"C7",X"80",X"38",X"80",X"07",X"C7",
		X"88",X"38",X"88",X"06",X"C7",X"A8",X"38",X"A8",X"07",X"C7",X"B0",X"38",X"B0",X"06",X"EF",X"80",
		X"D0",X"80",X"07",X"EF",X"88",X"D0",X"88",X"06",X"2F",X"A8",X"10",X"A8",X"07",X"2F",X"B0",X"10",
		X"B0",X"06",X"C7",X"D0",X"38",X"D0",X"07",X"C7",X"D8",X"38",X"D8",X"06",X"47",X"F8",X"10",X"F8",
		X"0C",X"67",X"44",X"48",X"44",X"0F",X"BF",X"88",X"40",X"88",X"0F",X"BF",X"B0",X"40",X"B0",X"0F",
		X"BF",X"D8",X"40",X"D8",X"AA",X"16",X"75",X"F1",X"76",X"AA",X"75",X"6A",X"76",X"EA",X"76",X"FB",
		X"76",X"2A",X"75",X"11",X"75",X"1B",X"75",X"F6",X"76",X"00",X"10",X"10",X"10",X"10",X"30",X"31",
		X"32",X"33",X"34",X"35",X"36",X"37",X"38",X"39",X"3A",X"3B",X"3C",X"3D",X"3E",X"3F",X"40",X"41",
		X"42",X"43",X"38",X"44",X"45",X"46",X"47",X"48",X"49",X"4A",X"4B",X"4B",X"4B",X"4C",X"38",X"46",
		X"47",X"47",X"4D",X"4E",X"38",X"4F",X"4B",X"4B",X"50",X"51",X"38",X"52",X"10",X"53",X"54",X"55",
		X"56",X"57",X"10",X"58",X"59",X"5A",X"79",X"8A",X"10",X"A7",X"A9",X"AB",X"78",X"7F",X"90",X"A6",
		X"A8",X"AA",X"77",X"7E",X"8F",X"97",X"9E",X"A5",X"76",X"7D",X"8E",X"96",X"9D",X"A4",X"75",X"7C",
		X"8D",X"95",X"9C",X"A3",X"74",X"7B",X"8C",X"94",X"9B",X"A2",X"73",X"7A",X"8B",X"93",X"9A",X"A1",
		X"62",X"6A",X"72",X"92",X"99",X"A0",X"61",X"69",X"71",X"91",X"98",X"9F",X"60",X"68",X"70",X"5B",
		X"63",X"6B",X"5F",X"67",X"6F",X"5E",X"66",X"6E",X"5D",X"65",X"6D",X"5C",X"64",X"6C",X"5B",X"63",
		X"6B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"74",X"00",X"00",X"00",X"23",X"68",
		X"01",X"11",X"00",X"00",X"00",X"10",X"DB",X"68",X"01",X"40",X"00",X"00",X"06",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"01",X"20",X"01",
		X"FF",X"10",X"FF",X"34",X"C3",X"39",X"00",X"67",X"80",X"69",X"1A",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"1E",X"18",X"0B",X"4B",
		X"14",X"18",X"0B",X"4B",X"1E",X"18",X"0B",X"3B",X"14",X"18",X"0B",X"3B",X"3D",X"0E",X"01",X"01",
		X"4D",X"0E",X"04",X"01",X"27",X"70",X"01",X"E0",X"00",X"00",X"00",X"40",X"01",X"78",X"02",X"00",
		X"27",X"49",X"0C",X"F0",X"00",X"49",X"0C",X"88",X"1E",X"07",X"03",X"09",X"24",X"64",X"BB",X"C0",
		X"00",X"00",X"00",X"00",X"1B",X"8C",X"7C",X"64",X"44",X"02",X"08",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"30",X"70",X"00",X"98",X"D0",X"70",X"00",X"98",X"10",X"70",X"00",X"CC",
		X"98",X"70",X"00",X"CC",X"68",X"70",X"00",X"EC",X"D0",X"70",X"00",X"EC",X"2B",X"1A",X"0B",X"63",
		X"6B",X"1C",X"0C",X"63",X"8B",X"1B",X"0B",X"A3",X"A3",X"1A",X"0B",X"6B",X"9B",X"1C",X"0C",X"18",
		X"5B",X"1C",X"0C",X"60",X"A3",X"1A",X"0B",X"83",X"2B",X"1A",X"0B",X"60",X"6B",X"1C",X"0C",X"6B",
		X"8B",X"1C",X"0C",X"93",X"73",X"1C",X"0C",X"BB",X"6B",X"6B",X"8B",X"93",X"73",X"BB",X"00",X"00",
		X"11",X"01",X"00",X"06",X"79",X"1F",X"D2",X"28",X"1E",X"1E",X"03",X"06",X"7B",X"1F",X"D2",X"28",
		X"1E",X"1E",X"04",X"06",X"7C",X"C3",X"28",X"1E",X"3A",X"27",X"62",X"E5",X"EF",X"00",X"00",X"E0",
		X"28",X"99",X"3E",X"E0",X"28",X"99",X"3E",X"00",X"00",X"E1",X"AF",X"32",X"60",X"60",X"06",X"0A",
		X"11",X"20",X"00",X"DD",X"21",X"00",X"67",X"CD",X"C3",X"3E",X"06",X"05",X"DD",X"21",X"00",X"64",
		X"CD",X"C3",X"3E",X"3A",X"60",X"60",X"A7",X"C8",X"FE",X"01",X"C8",X"FE",X"03",X"3E",X"03",X"D8",
		X"3E",X"07",X"C9",X"DD",X"CB",X"00",X"46",X"CA",X"FA",X"3E",X"79",X"DD",X"96",X"05",X"D2",X"D3",
		X"3E",X"ED",X"44",X"3C",X"95",X"DA",X"DE",X"3E",X"DD",X"96",X"0A",X"D2",X"FA",X"3E",X"FD",X"7E",
		X"03",X"DD",X"96",X"03",X"D2",X"E9",X"3E",X"ED",X"44",X"94",X"DA",X"F3",X"3E",X"DD",X"96",X"09",
		X"D2",X"FA",X"3E",X"3A",X"60",X"60",X"3C",X"32",X"60",X"60",X"DD",X"19",X"10",X"C5",X"C9",X"20",
		X"0E",X"DD",X"CB",X"01",X"4E",X"20",X"08",X"3E",X"01",X"DD",X"AE",X"01",X"DD",X"77",X"01",X"79",
		X"DD",X"86",X"03",X"DD",X"77",X"03",X"DD",X"19",X"11",X"04",X"00",X"05",X"C2",X"54",X"21",X"3A",
		X"54",X"69",X"FE",X"07",X"C0",X"21",X"09",X"60",X"36",X"80",X"23",X"34",X"AF",X"32",X"89",X"60",
		X"21",X"B7",X"76",X"11",X"7A",X"5C",X"C3",X"65",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"21",X"BE",X"6A",X"34",X"7E",X"FE",X"05",X"C2",X"64",X"4C",X"36",X"00",X"C3",X"36",X"4C",X"21",
		X"BE",X"6A",X"34",X"7E",X"FE",X"03",X"C2",X"64",X"4C",X"36",X"00",X"C3",X"36",X"4C",X"00",X"73",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CD",X"A6",X"3F",X"C3",X"5F",X"0D",X"3E",X"00",X"F7",X"06",X"02",X"21",X"6C",X"77",X"36",X"10",
		X"23",X"23",X"36",X"C0",X"21",X"8C",X"74",X"10",X"F5",X"C9",X"00",X"00",X"00",X"00",X"02",X"2B",
		X"48",X"2B",X"E8",X"02",X"43",X"48",X"43",X"E8",X"02",X"5B",X"48",X"5B",X"E8",X"02",X"73",X"48",
		X"73",X"E8",X"02",X"8B",X"48",X"8B",X"E8",X"02",X"A3",X"48",X"A3",X"E8",X"02",X"BB",X"48",X"BB",
		X"E8",X"02",X"D3",X"48",X"D3",X"E8",X"09",X"E7",X"48",X"18",X"48",X"10",X"E7",X"50",X"18",X"50",
		X"09",X"EF",X"F8",X"10",X"F8",X"0E",X"18",X"58",X"18",X"F0",X"0E",X"E3",X"58",X"E3",X"F0",X"AA",
		X"08",X"03",X"88",X"DD",X"36",X"00",X"01",X"DD",X"36",X"0C",X"01",X"DD",X"36",X"09",X"04",X"3E",
		X"02",X"F7",X"3A",X"29",X"62",X"FE",X"01",X"28",X"20",X"3A",X"05",X"62",X"FE",X"58",X"21",X"BD",
		X"02",X"38",X"0F",X"CD",X"57",X"00",X"E6",X"0F",X"FE",X"04",X"21",X"BD",X"02",X"30",X"03",X"21",
		X"3D",X"04",X"DD",X"74",X"02",X"DD",X"75",X"07",X"C9",X"3A",X"05",X"62",X"FE",X"58",X"30",X"E3",
		X"CD",X"57",X"00",X"E6",X"0F",X"FE",X"0E",X"18",X"E1",X"3A",X"27",X"62",X"FE",X"02",X"20",X"27",
		X"3A",X"05",X"62",X"FE",X"41",X"38",X"20",X"FE",X"48",X"30",X"1C",X"3A",X"03",X"62",X"FE",X"9C",
		X"30",X"15",X"FE",X"98",X"38",X"11",X"E1",X"3A",X"07",X"62",X"E6",X"80",X"F6",X"01",X"32",X"07",
		X"62",X"32",X"A0",X"6A",X"C3",X"3A",X"1C",X"3A",X"27",X"62",X"EE",X"03",X"C9",X"3A",X"27",X"62",
		X"FE",X"02",X"C8",X"FE",X"04",X"C9",X"3A",X"15",X"62",X"A7",X"C8",X"C3",X"F2",X"1C",X"7E",X"FE",
		X"AA",X"C8",X"C6",X"C8",X"C9",X"CD",X"AA",X"40",X"21",X"0A",X"60",X"C9",X"32",X"4C",X"69",X"CD",
		X"AA",X"40",X"C9",X"32",X"4F",X"69",X"CD",X"AA",X"40",X"C9",X"21",X"4C",X"69",X"3A",X"03",X"62",
		X"C6",X"08",X"77",X"2C",X"3A",X"07",X"62",X"77",X"2C",X"3E",X"07",X"77",X"2C",X"3A",X"05",X"62",
		X"77",X"21",X"54",X"69",X"3A",X"03",X"62",X"D6",X"08",X"77",X"2C",X"3A",X"07",X"62",X"47",X"E6",
		X"80",X"4F",X"78",X"E6",X"7F",X"C6",X"64",X"B1",X"77",X"2C",X"07",X"30",X"0E",X"3A",X"4C",X"69",
		X"F5",X"3A",X"54",X"69",X"32",X"4C",X"69",X"F1",X"32",X"54",X"69",X"3E",X"07",X"77",X"2C",X"3A",
		X"05",X"62",X"77",X"C9",X"C2",X"03",X"1D",X"CB",X"47",X"20",X"03",X"CB",X"4F",X"C8",X"3A",X"0F",
		X"62",X"A7",X"C2",X"8A",X"1D",X"CD",X"10",X"41",X"3E",X"0C",X"32",X"0F",X"62",X"C3",X"49",X"1D",
		X"3A",X"07",X"62",X"47",X"E6",X"03",X"78",X"28",X"02",X"E6",X"7F",X"21",X"00",X"40",X"01",X"03",
		X"00",X"ED",X"B1",X"2B",X"3A",X"10",X"60",X"0F",X"38",X"6E",X"0F",X"30",X"68",X"CD",X"CA",X"41",
		X"CD",X"8F",X"41",X"7D",X"E6",X"FC",X"47",X"2D",X"7D",X"E6",X"03",X"FE",X"03",X"20",X"01",X"3D",
		X"4F",X"B0",X"6F",X"79",X"FE",X"02",X"7E",X"CD",X"59",X"41",X"F5",X"CD",X"66",X"41",X"F1",X"D0",
		X"3A",X"03",X"62",X"D6",X"0C",X"32",X"03",X"62",X"C9",X"F5",X"32",X"07",X"62",X"E6",X"7F",X"FE",
		X"08",X"CC",X"8F",X"1D",X"F1",X"C9",X"32",X"92",X"6A",X"4F",X"E6",X"80",X"EE",X"80",X"47",X"79",
		X"E6",X"7F",X"FE",X"03",X"28",X"05",X"AF",X"32",X"80",X"6A",X"C9",X"3E",X"04",X"B0",X"32",X"07",
		X"62",X"3E",X"01",X"32",X"91",X"6A",X"C9",X"3A",X"03",X"62",X"FE",X"EB",X"D8",X"18",X"06",X"3A",
		X"03",X"62",X"FE",X"14",X"D0",X"33",X"33",X"C9",X"CD",X"CA",X"41",X"CD",X"87",X"41",X"7D",X"E6",
		X"FC",X"47",X"2C",X"7D",X"E6",X"03",X"FE",X"03",X"20",X"01",X"AF",X"4F",X"B0",X"6F",X"79",X"FE",
		X"01",X"F5",X"7E",X"FE",X"03",X"20",X"02",X"F6",X"80",X"CD",X"59",X"41",X"CD",X"66",X"41",X"F1",
		X"D8",X"3A",X"03",X"62",X"C6",X"0C",X"32",X"03",X"62",X"C9",X"3A",X"07",X"62",X"47",X"E6",X"7F",
		X"FE",X"03",X"20",X"06",X"E5",X"CD",X"2E",X"42",X"E1",X"C9",X"E5",X"CD",X"E0",X"41",X"E1",X"C9",
		X"3A",X"07",X"62",X"CB",X"7F",X"20",X"3A",X"3A",X"10",X"60",X"CB",X"47",X"0E",X"F0",X"28",X"1E",
		X"0E",X"05",X"3A",X"03",X"62",X"81",X"67",X"57",X"3A",X"05",X"62",X"47",X"C6",X"F8",X"6F",X"78",
		X"C6",X"05",X"5F",X"01",X"01",X"00",X"CD",X"D3",X"46",X"A7",X"C8",X"C3",X"6E",X"42",X"3A",X"03",
		X"62",X"81",X"67",X"57",X"3A",X"05",X"62",X"47",X"C6",X"F8",X"6F",X"78",X"C6",X"05",X"5F",X"18",
		X"E2",X"3A",X"10",X"60",X"CB",X"47",X"0E",X"FB",X"28",X"C8",X"0E",X"10",X"18",X"E0",X"CD",X"42",
		X"46",X"3A",X"10",X"60",X"CB",X"47",X"3A",X"81",X"6A",X"28",X"03",X"3A",X"82",X"6A",X"A7",X"C0",
		X"AF",X"32",X"15",X"62",X"21",X"03",X"62",X"3A",X"03",X"62",X"67",X"3A",X"05",X"62",X"C6",X"0E",
		X"6F",X"CD",X"F0",X"2F",X"7E",X"FE",X"D0",X"3A",X"10",X"60",X"38",X"05",X"0F",X"3E",X"81",X"18",
		X"03",X"0F",X"3E",X"8E",X"32",X"07",X"62",X"38",X"05",X"E6",X"7F",X"32",X"07",X"62",X"33",X"33",
		X"33",X"33",X"33",X"33",X"33",X"33",X"3A",X"8D",X"6A",X"A7",X"3E",X"00",X"20",X"05",X"3C",X"32",
		X"A2",X"6A",X"3D",X"32",X"8D",X"6A",X"32",X"98",X"63",X"32",X"80",X"6A",X"3A",X"05",X"62",X"E6",
		X"FC",X"32",X"05",X"62",X"C9",X"3A",X"80",X"6A",X"A7",X"3E",X"03",X"20",X"02",X"3E",X"01",X"32",
		X"0F",X"62",X"3E",X"03",X"20",X"02",X"3E",X"03",X"C9",X"AF",X"32",X"9D",X"6A",X"3A",X"80",X"6A",
		X"A7",X"3E",X"04",X"20",X"02",X"3E",X"06",X"32",X"0F",X"62",X"3E",X"FD",X"20",X"02",X"3E",X"FE",
		X"C9",X"CA",X"67",X"1D",X"47",X"3A",X"80",X"6A",X"A7",X"78",X"C2",X"31",X"1D",X"C3",X"49",X"1D",
		X"3A",X"10",X"60",X"CB",X"57",X"C2",X"E6",X"43",X"AF",X"32",X"9D",X"6A",X"3A",X"8D",X"6A",X"A7",
		X"20",X"17",X"CD",X"42",X"46",X"4F",X"3A",X"80",X"6A",X"A7",X"20",X"37",X"79",X"A7",X"28",X"1B",
		X"CD",X"6E",X"43",X"A7",X"CA",X"A9",X"1D",X"18",X"40",X"CD",X"AD",X"43",X"4F",X"3A",X"07",X"62",
		X"E6",X"7F",X"FE",X"03",X"28",X"33",X"79",X"A7",X"C2",X"A9",X"1D",X"3A",X"8D",X"6A",X"A7",X"3E",
		X"00",X"20",X"03",X"32",X"8C",X"6A",X"32",X"15",X"62",X"32",X"80",X"6A",X"32",X"8D",X"6A",X"32",
		X"98",X"63",X"C9",X"3A",X"81",X"6A",X"4F",X"3A",X"82",X"6A",X"47",X"B1",X"28",X"DD",X"78",X"A1",
		X"28",X"1B",X"CD",X"6E",X"43",X"A7",X"CA",X"A9",X"1D",X"3A",X"4F",X"69",X"32",X"05",X"62",X"3A",
		X"4D",X"69",X"32",X"07",X"62",X"3E",X"00",X"32",X"24",X"62",X"C3",X"A9",X"1D",X"78",X"A7",X"3A",
		X"03",X"62",X"20",X"11",X"D6",X"0C",X"32",X"03",X"62",X"3E",X"08",X"32",X"07",X"62",X"AF",X"32",
		X"80",X"6A",X"C3",X"A9",X"1D",X"C6",X"0C",X"32",X"03",X"62",X"3E",X"88",X"18",X"ED",X"3A",X"80",
		X"6A",X"A7",X"28",X"26",X"01",X"20",X"00",X"C5",X"06",X"00",X"0E",X"07",X"3A",X"03",X"62",X"80",
		X"67",X"3A",X"05",X"62",X"81",X"6F",X"C1",X"CD",X"F0",X"2F",X"7E",X"FE",X"D0",X"3E",X"00",X"D8",
		X"7E",X"E6",X"0F",X"FE",X"08",X"3E",X"00",X"D0",X"3C",X"C9",X"01",X"01",X"00",X"C5",X"0E",X"07",
		X"3A",X"07",X"62",X"CB",X"7F",X"06",X"07",X"28",X"D3",X"06",X"F8",X"18",X"CF",X"DD",X"21",X"00",
		X"66",X"11",X"10",X"00",X"06",X"02",X"3A",X"03",X"62",X"4F",X"C6",X"FC",X"DD",X"BE",X"03",X"30",
		X"09",X"C6",X"08",X"DD",X"BE",X"03",X"38",X"02",X"18",X"06",X"DD",X"19",X"79",X"10",X"EB",X"C9",
		X"3A",X"05",X"62",X"47",X"DD",X"7E",X"05",X"C6",X"F8",X"B8",X"30",X"08",X"C6",X"15",X"B8",X"38",
		X"03",X"3E",X"01",X"C9",X"AF",X"C9",X"3A",X"8D",X"6A",X"A7",X"20",X"58",X"CD",X"42",X"46",X"4F",
		X"3A",X"80",X"6A",X"A7",X"79",X"20",X"63",X"A7",X"CA",X"39",X"43",X"3A",X"80",X"6A",X"A7",X"06",
		X"00",X"28",X"23",X"3A",X"03",X"62",X"47",X"C6",X"0C",X"67",X"78",X"C6",X"F4",X"57",X"3A",X"05",
		X"62",X"D6",X"08",X"6F",X"5F",X"C1",X"CD",X"D3",X"46",X"A7",X"CA",X"A9",X"1D",X"3A",X"4F",X"69",
		X"32",X"05",X"62",X"C3",X"A9",X"1D",X"01",X"01",X"00",X"C5",X"3A",X"07",X"62",X"CB",X"7F",X"06",
		X"08",X"28",X"02",X"06",X"F8",X"3A",X"03",X"62",X"80",X"67",X"57",X"3A",X"05",X"62",X"D6",X"08",
		X"6F",X"5F",X"18",X"D1",X"CD",X"AD",X"43",X"4F",X"3A",X"07",X"62",X"E6",X"7F",X"FE",X"03",X"CA",
		X"39",X"43",X"79",X"A7",X"C2",X"A9",X"1D",X"C3",X"39",X"43",X"01",X"20",X"00",X"C5",X"3A",X"81",
		X"6A",X"4F",X"3A",X"82",X"6A",X"A1",X"CA",X"39",X"43",X"18",X"90",X"2D",X"2D",X"3A",X"80",X"6A",
		X"B7",X"7E",X"CA",X"54",X"1D",X"C3",X"58",X"1D",X"E5",X"D5",X"C5",X"F5",X"08",X"3E",X"02",X"08",
		X"3A",X"16",X"62",X"A7",X"3A",X"03",X"62",X"CA",X"C2",X"45",X"C6",X"F7",X"57",X"3A",X"05",X"62",
		X"C6",X"FB",X"5F",X"3A",X"07",X"62",X"07",X"30",X"04",X"7A",X"C6",X"12",X"57",X"7A",X"F6",X"03",
		X"CB",X"97",X"57",X"21",X"00",X"63",X"3A",X"27",X"62",X"FE",X"03",X"01",X"15",X"00",X"20",X"02",
		X"0E",X"08",X"7A",X"ED",X"B1",X"C2",X"D9",X"45",X"E5",X"D5",X"C5",X"2B",X"7B",X"11",X"15",X"00",
		X"19",X"46",X"19",X"4E",X"CD",X"3A",X"46",X"C1",X"D1",X"E1",X"30",X"06",X"79",X"A7",X"20",X"E2",
		X"18",X"71",X"3A",X"16",X"62",X"A7",X"3A",X"07",X"62",X"CA",X"AF",X"45",X"E6",X"80",X"06",X"08",
		X"B0",X"4F",X"7A",X"FE",X"13",X"79",X"CB",X"BF",X"28",X"09",X"7A",X"FE",X"EB",X"79",X"CB",X"FF",
		X"28",X"01",X"79",X"32",X"07",X"62",X"7A",X"32",X"03",X"62",X"3E",X"0A",X"32",X"0F",X"62",X"3A",
		X"03",X"62",X"67",X"3A",X"05",X"62",X"C6",X"04",X"6F",X"CD",X"F0",X"2F",X"7E",X"FE",X"D0",X"38",
		X"0E",X"3E",X"01",X"32",X"21",X"62",X"32",X"8D",X"6A",X"3A",X"4D",X"69",X"32",X"07",X"62",X"AF",
		X"32",X"20",X"62",X"32",X"98",X"63",X"CD",X"4A",X"45",X"3C",X"32",X"15",X"62",X"CD",X"8F",X"1D",
		X"3A",X"05",X"62",X"FE",X"40",X"30",X"0C",X"3A",X"03",X"62",X"FE",X"70",X"30",X"05",X"3E",X"01",
		X"32",X"9E",X"6A",X"F1",X"C1",X"D1",X"E1",X"C3",X"A6",X"1D",X"AF",X"32",X"16",X"62",X"32",X"89",
		X"6A",X"32",X"8A",X"6A",X"32",X"8B",X"6A",X"C9",X"3A",X"27",X"62",X"FE",X"01",X"20",X"E4",X"3A",
		X"A2",X"6A",X"A7",X"20",X"DE",X"3A",X"8C",X"6A",X"A7",X"28",X"D8",X"3A",X"A2",X"6A",X"A7",X"20",
		X"D2",X"FD",X"21",X"00",X"62",X"FD",X"7E",X"05",X"C6",X"F8",X"4F",X"21",X"02",X"00",X"06",X"05",
		X"11",X"10",X"00",X"DD",X"21",X"D0",X"65",X"CD",X"FA",X"45",X"A7",X"28",X"B6",X"DD",X"7E",X"03",
		X"FD",X"77",X"03",X"FD",X"7E",X"07",X"E6",X"80",X"06",X"08",X"B0",X"FD",X"77",X"07",X"FD",X"36",
		X"0F",X"10",X"AF",X"CD",X"4A",X"45",X"3C",X"32",X"8D",X"6A",X"CD",X"F7",X"0B",X"18",X"94",X"E6",
		X"80",X"F6",X"08",X"32",X"07",X"62",X"7A",X"32",X"03",X"62",X"3E",X"10",X"32",X"0F",X"62",X"C3",
		X"FF",X"44",X"C6",X"F9",X"57",X"3A",X"05",X"62",X"C6",X"FB",X"5F",X"3A",X"07",X"62",X"07",X"D2",
		X"9D",X"44",X"7A",X"C6",X"10",X"57",X"C3",X"9D",X"44",X"08",X"3D",X"F5",X"08",X"F1",X"CA",X"58",
		X"45",X"3A",X"07",X"62",X"CB",X"7F",X"16",X"01",X"20",X"02",X"16",X"FF",X"3A",X"03",X"62",X"82",
		X"57",X"3A",X"05",X"62",X"C6",X"FB",X"5F",X"C3",X"9D",X"44",X"DD",X"CB",X"00",X"46",X"28",X"34",
		X"79",X"DD",X"96",X"05",X"30",X"02",X"ED",X"44",X"3C",X"95",X"38",X"05",X"DD",X"96",X"0A",X"30",
		X"23",X"C5",X"FD",X"7E",X"07",X"E6",X"80",X"0E",X"08",X"20",X"02",X"0E",X"F8",X"FD",X"7E",X"03",
		X"81",X"DD",X"96",X"03",X"C1",X"30",X"02",X"ED",X"44",X"94",X"38",X"05",X"DD",X"96",X"09",X"30",
		X"03",X"3E",X"01",X"C9",X"DD",X"19",X"10",X"C2",X"AF",X"C9",X"B8",X"D8",X"C5",X"47",X"79",X"B8",
		X"C1",X"C9",X"E5",X"D5",X"C5",X"3A",X"80",X"6A",X"B7",X"28",X"33",X"11",X"FB",X"F5",X"21",X"FB",
		X"0D",X"3A",X"07",X"62",X"07",X"30",X"06",X"11",X"FB",X"F3",X"21",X"FB",X"0B",X"3A",X"03",X"62",
		X"47",X"82",X"57",X"78",X"84",X"67",X"3A",X"05",X"62",X"47",X"83",X"5F",X"78",X"85",X"6F",X"CD",
		X"8F",X"46",X"32",X"81",X"6A",X"EB",X"CD",X"8F",X"46",X"32",X"82",X"6A",X"18",X"0D",X"3A",X"03",
		X"62",X"57",X"3A",X"05",X"62",X"C6",X"FB",X"5F",X"CD",X"8F",X"46",X"C1",X"D1",X"E1",X"C9",X"E5",
		X"C5",X"7A",X"F6",X"03",X"CB",X"97",X"57",X"21",X"00",X"63",X"01",X"15",X"00",X"7A",X"ED",X"B1",
		X"20",X"2D",X"E5",X"C5",X"D5",X"2B",X"11",X"15",X"00",X"19",X"46",X"19",X"4E",X"D1",X"7B",X"CD",
		X"3A",X"46",X"79",X"32",X"93",X"6A",X"C1",X"E1",X"38",X"E3",X"3A",X"8D",X"6A",X"A7",X"3E",X"01",
		X"28",X"0E",X"7A",X"C6",X"0C",X"32",X"03",X"62",X"AF",X"32",X"8D",X"6A",X"3C",X"18",X"01",X"AF",
		X"C1",X"E1",X"C9",X"DD",X"E5",X"D5",X"CD",X"F0",X"2F",X"D1",X"EB",X"D5",X"CD",X"F0",X"2F",X"D1",
		X"EB",X"DD",X"21",X"83",X"6A",X"7E",X"DD",X"77",X"00",X"09",X"DD",X"23",X"EB",X"E5",X"ED",X"52",
		X"E1",X"EB",X"30",X"F1",X"DD",X"36",X"00",X"00",X"21",X"83",X"6A",X"0E",X"00",X"7E",X"23",X"FE",
		X"00",X"28",X"05",X"FE",X"D0",X"38",X"F6",X"0C",X"79",X"DD",X"E1",X"C9",X"3A",X"05",X"62",X"FE",
		X"21",X"D0",X"3A",X"03",X"62",X"FE",X"50",X"D0",X"3E",X"05",X"32",X"07",X"62",X"3E",X"20",X"32",
		X"05",X"62",X"CD",X"A6",X"1D",X"C3",X"85",X"1E",X"DD",X"36",X"1D",X"01",X"CD",X"52",X"47",X"C9",
		X"3A",X"27",X"62",X"FE",X"02",X"20",X"0E",X"3A",X"03",X"62",X"DD",X"BE",X"03",X"38",X"0F",X"DD",
		X"36",X"0D",X"01",X"18",X"0D",X"E5",X"CD",X"57",X"00",X"E1",X"E6",X"03",X"20",X"F1",X"DD",X"36",
		X"0D",X"00",X"DD",X"7E",X"08",X"E6",X"7F",X"DD",X"77",X"08",X"0E",X"3E",X"DD",X"7E",X"07",X"E6",
		X"80",X"B1",X"DD",X"77",X"07",X"C9",X"DD",X"36",X"0D",X"08",X"DD",X"7E",X"08",X"F6",X"80",X"DD",
		X"77",X"08",X"0E",X"4E",X"18",X"E6",X"DD",X"36",X"0D",X"04",X"18",X"F6",X"CB",X"16",X"36",X"6F",
		X"38",X"02",X"36",X"6E",X"3E",X"01",X"AE",X"23",X"36",X"07",X"21",X"55",X"69",X"77",X"23",X"36",
		X"07",X"C9",X"CD",X"9C",X"23",X"3A",X"27",X"62",X"FE",X"02",X"20",X"21",X"3A",X"05",X"62",X"FE",
		X"F8",X"DA",X"C5",X"1B",X"3A",X"05",X"60",X"FE",X"01",X"3E",X"04",X"28",X"02",X"3E",X"0D",X"32",
		X"0A",X"60",X"3E",X"F8",X"32",X"05",X"62",X"3E",X"01",X"32",X"09",X"60",X"C9",X"FE",X"03",X"3A",
		X"05",X"62",X"20",X"07",X"FE",X"F9",X"DA",X"C5",X"1B",X"18",X"D9",X"FE",X"F8",X"DA",X"C5",X"1B",
		X"18",X"D2",X"3A",X"27",X"62",X"FE",X"04",X"DD",X"36",X"07",X"4E",X"C0",X"DD",X"36",X"07",X"3F",
		X"C9",X"3A",X"8F",X"6A",X"3D",X"20",X"0A",X"DD",X"36",X"00",X"02",X"3E",X"30",X"32",X"8F",X"6A",
		X"C9",X"32",X"8F",X"6A",X"33",X"33",X"C9",X"DD",X"7E",X"0C",X"A7",X"20",X"04",X"E1",X"C3",X"BA",
		X"21",X"DD",X"7E",X"03",X"C6",X"00",X"F6",X"03",X"CB",X"97",X"DD",X"77",X"03",X"DD",X"36",X"02",
		X"01",X"2C",X"2C",X"2C",X"67",X"7D",X"C6",X"08",X"57",X"7C",X"01",X"15",X"00",X"CD",X"2A",X"48",
		X"DD",X"70",X"17",X"CD",X"B2",X"21",X"E1",X"C3",X"BA",X"21",X"21",X"00",X"63",X"ED",X"B1",X"C2",
		X"53",X"48",X"E5",X"C5",X"01",X"14",X"00",X"09",X"0C",X"5F",X"7A",X"BE",X"30",X"0B",X"09",X"BE",
		X"CA",X"4E",X"48",X"57",X"7B",X"C1",X"E1",X"18",X"E4",X"09",X"3E",X"01",X"18",X"03",X"AF",X"ED",
		X"42",X"C1",X"46",X"E1",X"C9",X"DD",X"21",X"A0",X"65",X"21",X"30",X"69",X"11",X"10",X"00",X"06",
		X"06",X"CD",X"D3",X"11",X"DD",X"21",X"44",X"69",X"11",X"04",X"00",X"21",X"3C",X"69",X"06",X"02",
		X"7E",X"DD",X"77",X"00",X"23",X"23",X"DD",X"36",X"01",X"46",X"7E",X"DD",X"77",X"02",X"23",X"7E",
		X"DD",X"77",X"03",X"23",X"DD",X"19",X"10",X"E8",X"C9",X"21",X"18",X"3E",X"11",X"A7",X"65",X"01",
		X"0C",X"06",X"CD",X"2A",X"12",X"DD",X"E5",X"DD",X"21",X"00",X"66",X"21",X"DB",X"48",X"11",X"10",
		X"00",X"06",X"02",X"7E",X"DD",X"77",X"00",X"23",X"7E",X"DD",X"77",X"03",X"23",X"7E",X"DD",X"77",
		X"05",X"23",X"7E",X"DD",X"77",X"07",X"23",X"7E",X"DD",X"77",X"08",X"23",X"7E",X"DD",X"77",X"09",
		X"23",X"7E",X"DD",X"77",X"0A",X"23",X"DD",X"19",X"10",X"D9",X"21",X"B4",X"69",X"36",X"E0",X"23",
		X"36",X"4A",X"23",X"36",X"00",X"23",X"36",X"A0",X"DD",X"E1",X"C9",X"01",X"40",X"AB",X"46",X"02",
		X"08",X"04",X"01",X"60",X"B3",X"46",X"02",X"08",X"04",X"DD",X"21",X"A0",X"65",X"06",X"05",X"11",
		X"10",X"00",X"DD",X"E5",X"DD",X"36",X"00",X"01",X"DD",X"19",X"10",X"F8",X"DD",X"E1",X"DD",X"36",
		X"13",X"68",X"DD",X"36",X"15",X"D0",X"DD",X"36",X"23",X"95",X"DD",X"36",X"05",X"F4",X"DD",X"36",
		X"25",X"F4",X"DD",X"7E",X"23",X"C6",X"10",X"DD",X"77",X"03",X"3E",X"A3",X"DD",X"77",X"35",X"DD",
		X"77",X"45",X"3E",X"36",X"DD",X"77",X"33",X"C6",X"30",X"DD",X"77",X"43",X"DD",X"36",X"37",X"45",
		X"DD",X"36",X"47",X"45",X"3E",X"01",X"DD",X"77",X"1C",X"DD",X"77",X"2C",X"DD",X"77",X"3C",X"3E",
		X"60",X"32",X"A0",X"62",X"3E",X"B8",X"32",X"A3",X"62",X"C9",X"3E",X"0E",X"F7",X"3E",X"01",X"32",
		X"A0",X"63",X"C9",X"FE",X"A3",X"28",X"0B",X"FE",X"D0",X"C2",X"B4",X"25",X"3A",X"A4",X"63",X"C3",
		X"CF",X"25",X"3A",X"A3",X"63",X"84",X"DD",X"77",X"03",X"C6",X"30",X"DD",X"77",X"13",X"F5",X"E5",
		X"E6",X"07",X"20",X"0B",X"21",X"B5",X"69",X"CB",X"7E",X"36",X"CA",X"28",X"02",X"36",X"4A",X"E1",
		X"F1",X"C3",X"BB",X"25",X"3A",X"1A",X"60",X"00",X"00",X"00",X"C9",X"3A",X"1A",X"60",X"E6",X"03",
		X"CA",X"EF",X"26",X"AF",X"C9",X"3A",X"98",X"63",X"A7",X"CA",X"95",X"2A",X"3A",X"27",X"62",X"FE",
		X"01",X"C8",X"AF",X"32",X"16",X"62",X"C3",X"95",X"2A",X"3A",X"98",X"63",X"A7",X"C8",X"DD",X"21",
		X"B0",X"65",X"11",X"10",X"00",X"48",X"06",X"03",X"3A",X"05",X"62",X"C6",X"0C",X"DD",X"BE",X"05",
		X"28",X"05",X"DD",X"19",X"10",X"F7",X"C9",X"21",X"A3",X"63",X"7D",X"80",X"6F",X"78",X"FE",X"03",
		X"20",X"0E",X"16",X"0C",X"1E",X"18",X"7E",X"F2",X"ED",X"49",X"16",X"09",X"1E",X"13",X"18",X"0D",
		X"7E",X"B7",X"16",X"1C",X"1E",X"2A",X"F2",X"ED",X"49",X"16",X"18",X"1E",X"20",X"DD",X"7E",X"03",
		X"82",X"47",X"3A",X"03",X"62",X"B8",X"30",X"0B",X"78",X"93",X"47",X"3A",X"03",X"62",X"B8",X"38",
		X"02",X"AF",X"C9",X"AF",X"32",X"98",X"63",X"3C",X"32",X"16",X"62",X"32",X"21",X"62",X"C9",X"3A",
		X"98",X"63",X"47",X"3A",X"8D",X"6A",X"A7",X"20",X"3A",X"3A",X"03",X"62",X"47",X"3A",X"05",X"62",
		X"FE",X"9C",X"28",X"0F",X"FE",X"C4",X"28",X"13",X"FE",X"E8",X"C0",X"21",X"34",X"3E",X"11",X"A6",
		X"63",X"18",X"0E",X"21",X"24",X"3E",X"11",X"A3",X"63",X"18",X"06",X"21",X"2C",X"3E",X"11",X"A4",
		X"63",X"78",X"BE",X"D8",X"23",X"23",X"23",X"23",X"BE",X"D0",X"3A",X"98",X"63",X"A7",X"C8",X"1A",
		X"C3",X"02",X"2B",X"21",X"24",X"3E",X"11",X"A3",X"63",X"3A",X"03",X"62",X"47",X"18",X"F0",X"DD",
		X"77",X"03",X"C6",X"10",X"DD",X"77",X"E3",X"C9",X"32",X"98",X"63",X"3D",X"32",X"8E",X"6A",X"32",
		X"8D",X"6A",X"CD",X"75",X"4E",X"3C",X"C9",X"11",X"10",X"00",X"3A",X"8C",X"6A",X"A7",X"CA",X"27",
		X"2A",X"3A",X"8E",X"6A",X"A7",X"CA",X"EB",X"29",X"C3",X"27",X"2A",X"32",X"8D",X"6A",X"3C",X"32",
		X"8E",X"6A",X"C9",X"32",X"8E",X"6A",X"E1",X"E1",X"C9",X"3E",X"00",X"32",X"8E",X"6A",X"C3",X"A6",
		X"1D",X"3E",X"01",X"18",X"F6",X"DD",X"7E",X"0F",X"3D",X"20",X"1E",X"3A",X"27",X"62",X"FE",X"04",
		X"DD",X"7E",X"07",X"20",X"0D",X"DD",X"7E",X"0C",X"A7",X"DD",X"7E",X"07",X"28",X"04",X"EE",X"7F",
		X"18",X"02",X"EE",X"03",X"DD",X"77",X"07",X"3E",X"04",X"DD",X"77",X"0F",X"C9",X"DD",X"E5",X"DD",
		X"CB",X"00",X"46",X"28",X"58",X"CD",X"35",X"4B",X"7C",X"DD",X"86",X"0A",X"4F",X"FD",X"7E",X"05",
		X"91",X"DD",X"BE",X"05",X"28",X"02",X"30",X"45",X"7D",X"DD",X"86",X"0A",X"FD",X"86",X"05",X"DD",
		X"BE",X"05",X"38",X"39",X"CD",X"6C",X"4B",X"7C",X"DD",X"86",X"09",X"4F",X"FD",X"7E",X"03",X"91",
		X"DD",X"BE",X"03",X"28",X"02",X"30",X"26",X"7D",X"DD",X"86",X"09",X"FD",X"86",X"03",X"DD",X"BE",
		X"03",X"38",X"1A",X"3A",X"27",X"62",X"FE",X"02",X"20",X"08",X"DD",X"36",X"07",X"3D",X"DD",X"36",
		X"08",X"0E",X"DD",X"22",X"9A",X"6A",X"3E",X"01",X"DD",X"E1",X"33",X"33",X"C9",X"DD",X"19",X"10",
		X"9E",X"AF",X"DD",X"E1",X"C9",X"3A",X"07",X"62",X"E6",X"0F",X"21",X"05",X"05",X"C8",X"FE",X"01",
		X"21",X"05",X"05",X"C8",X"FE",X"02",X"21",X"05",X"05",X"C8",X"FE",X"03",X"21",X"05",X"07",X"C8",
		X"FE",X"04",X"21",X"07",X"05",X"C8",X"FE",X"08",X"21",X"05",X"06",X"C8",X"FE",X"09",X"21",X"05",
		X"06",X"C8",X"FE",X"0E",X"21",X"05",X"04",X"C8",X"21",X"05",X"05",X"C9",X"CD",X"79",X"4B",X"3A",
		X"07",X"62",X"CB",X"7F",X"C8",X"7C",X"65",X"6F",X"C9",X"3A",X"07",X"62",X"E6",X"0F",X"21",X"05",
		X"05",X"C8",X"FE",X"01",X"21",X"05",X"05",X"C8",X"FE",X"02",X"21",X"05",X"05",X"C8",X"FE",X"03",
		X"21",X"0B",X"0C",X"C8",X"FE",X"04",X"21",X"06",X"08",X"C8",X"FE",X"08",X"21",X"0B",X"02",X"C8",
		X"FE",X"09",X"21",X"0B",X"02",X"C8",X"FE",X"0E",X"21",X"04",X"04",X"C8",X"21",X"05",X"05",X"C9",
		X"FE",X"00",X"20",X"41",X"DD",X"35",X"03",X"3A",X"27",X"62",X"FE",X"03",X"20",X"22",X"DD",X"7E",
		X"05",X"FE",X"A0",X"30",X"1B",X"DD",X"7E",X"03",X"FE",X"20",X"D2",X"6C",X"2E",X"DD",X"36",X"0D",
		X"08",X"FD",X"36",X"01",X"11",X"DD",X"7E",X"05",X"C6",X"33",X"DD",X"77",X"06",X"C3",X"6C",X"2E",
		X"DD",X"7E",X"03",X"FE",X"08",X"D2",X"6C",X"2E",X"AF",X"DD",X"77",X"00",X"DD",X"77",X"03",X"DD",
		X"77",X"05",X"C3",X"6C",X"2E",X"FE",X"04",X"20",X"79",X"DD",X"7E",X"05",X"FE",X"58",X"DA",X"96",
		X"2E",X"78",X"FE",X"02",X"C2",X"C6",X"4C",X"3A",X"05",X"62",X"C6",X"FE",X"DD",X"BE",X"05",X"D2",
		X"DF",X"4C",X"C6",X"04",X"DD",X"BE",X"05",X"DA",X"DF",X"4C",X"AF",X"DD",X"77",X"0D",X"3A",X"27",
		X"62",X"FE",X"03",X"28",X"46",X"3A",X"29",X"62",X"3D",X"20",X"07",X"C3",X"40",X"3F",X"00",X"00",
		X"00",X"00",X"C3",X"4F",X"3F",X"00",X"3A",X"BF",X"6A",X"A7",X"20",X"28",X"3A",X"05",X"62",X"FE",
		X"43",X"30",X"07",X"3E",X"01",X"32",X"BF",X"6A",X"18",X"1A",X"DD",X"36",X"01",X"01",X"DD",X"7E",
		X"03",X"C6",X"08",X"DD",X"77",X"0B",X"DD",X"7E",X"05",X"DD",X"77",X"0C",X"DD",X"36",X"02",X"75",
		X"DD",X"36",X"04",X"0C",X"FD",X"36",X"01",X"BB",X"C3",X"6C",X"2E",X"FD",X"36",X"01",X"93",X"C3",
		X"6C",X"2E",X"FE",X"02",X"20",X"29",X"DD",X"34",X"03",X"DD",X"7E",X"03",X"FE",X"E0",X"DA",X"6C",
		X"2E",X"DD",X"36",X"0D",X"10",X"FD",X"36",X"01",X"11",X"3A",X"29",X"62",X"FE",X"03",X"DD",X"7E",
		X"05",X"38",X"04",X"C6",X"42",X"18",X"02",X"C6",X"2D",X"DD",X"77",X"06",X"C3",X"6C",X"2E",X"E6",
		X"18",X"CA",X"31",X"2E",X"DD",X"34",X"05",X"DD",X"7E",X"05",X"DD",X"BE",X"06",X"C2",X"6C",X"2E",
		X"DD",X"7E",X"0D",X"FE",X"08",X"21",X"93",X"00",X"20",X"03",X"21",X"13",X"02",X"DD",X"74",X"0D",
		X"FD",X"75",X"01",X"C3",X"6C",X"2E",X"DD",X"7E",X"05",X"FE",X"58",X"28",X"2C",X"FE",X"60",X"0E",
		X"02",X"28",X"17",X"FE",X"68",X"0E",X"05",X"28",X"11",X"FE",X"70",X"0E",X"03",X"28",X"0B",X"DD",
		X"7E",X"05",X"FE",X"78",X"CA",X"1A",X"4C",X"C3",X"96",X"2E",X"79",X"B8",X"CA",X"1A",X"4C",X"78",
		X"D6",X"05",X"B9",X"CA",X"1A",X"4C",X"C3",X"96",X"2E",X"3A",X"27",X"62",X"FE",X"03",X"20",X"05",
		X"DD",X"7E",X"05",X"18",X"C8",X"3E",X"04",X"18",X"E1",X"DD",X"7E",X"0D",X"E6",X"1C",X"C2",X"29",
		X"2E",X"3A",X"27",X"62",X"FE",X"03",X"FD",X"7E",X"01",X"20",X"04",X"EE",X"01",X"18",X"02",X"EE",
		X"07",X"FD",X"77",X"01",X"C3",X"29",X"2E",X"DD",X"36",X"0D",X"04",X"3A",X"27",X"62",X"FE",X"03",
		X"3E",X"3A",X"20",X"02",X"3E",X"11",X"FD",X"77",X"01",X"C9",X"3E",X"0E",X"F7",X"CD",X"ED",X"30",
		X"C9",X"3E",X"05",X"F7",X"21",X"A4",X"6A",X"7E",X"FE",X"70",X"28",X"01",X"34",X"C3",X"08",X"2E",
		X"CD",X"86",X"11",X"CD",X"69",X"4D",X"3E",X"01",X"32",X"60",X"66",X"3E",X"44",X"32",X"63",X"66",
		X"3E",X"F8",X"32",X"65",X"66",X"21",X"EC",X"3D",X"C9",X"21",X"75",X"4D",X"11",X"67",X"66",X"06",
		X"01",X"CD",X"2A",X"12",X"C9",X"50",X"0F",X"08",X"04",X"3A",X"90",X"6A",X"A7",X"28",X"05",X"3D",
		X"32",X"90",X"6A",X"C9",X"3E",X"01",X"32",X"90",X"6A",X"3A",X"10",X"60",X"1E",X"01",X"CB",X"47",
		X"20",X"08",X"1E",X"FF",X"CB",X"4F",X"20",X"02",X"1E",X"00",X"3A",X"03",X"62",X"83",X"32",X"03",
		X"62",X"3E",X"01",X"32",X"0F",X"62",X"3A",X"89",X"6A",X"A7",X"3A",X"67",X"66",X"20",X"54",X"FE",
		X"53",X"28",X"0B",X"3C",X"32",X"67",X"66",X"47",X"0E",X"00",X"3E",X"00",X"18",X"09",X"3D",X"32",
		X"67",X"66",X"47",X"0E",X"04",X"3E",X"01",X"32",X"89",X"6A",X"78",X"E6",X"03",X"B1",X"5F",X"16",
		X"00",X"21",X"26",X"4E",X"19",X"46",X"3A",X"05",X"62",X"80",X"32",X"05",X"62",X"32",X"4F",X"69",
		X"32",X"57",X"69",X"3A",X"87",X"6A",X"A7",X"C0",X"3A",X"10",X"60",X"07",X"D0",X"3A",X"67",X"66",
		X"32",X"8A",X"6A",X"3E",X"01",X"32",X"87",X"6A",X"3A",X"89",X"6A",X"A7",X"C0",X"3E",X"53",X"32",
		X"8A",X"6A",X"C9",X"FE",X"50",X"20",X"B7",X"3A",X"8A",X"6A",X"A7",X"20",X"05",X"3E",X"54",X"32",
		X"8A",X"6A",X"AF",X"32",X"8B",X"6A",X"32",X"98",X"63",X"3A",X"9F",X"6A",X"32",X"10",X"60",X"AF",
		X"32",X"9F",X"6A",X"C3",X"6E",X"1B",X"00",X"02",X"03",X"03",X"FB",X"FB",X"FD",X"00",X"DD",X"21",
		X"00",X"62",X"CD",X"29",X"2B",X"AF",X"32",X"88",X"6A",X"CD",X"AF",X"29",X"3A",X"27",X"62",X"3D",
		X"28",X"03",X"AF",X"47",X"C9",X"CD",X"4B",X"4E",X"AF",X"47",X"C9",X"3E",X"01",X"32",X"88",X"6A",
		X"FD",X"21",X"00",X"62",X"FD",X"7E",X"05",X"4F",X"21",X"08",X"08",X"CD",X"68",X"4E",X"A7",X"CA",
		X"20",X"2A",X"3E",X"01",X"90",X"C3",X"C7",X"29",X"06",X"01",X"11",X"10",X"00",X"DD",X"21",X"60",
		X"66",X"CD",X"13",X"29",X"C9",X"3A",X"88",X"6A",X"A7",X"C8",X"3E",X"01",X"32",X"8B",X"6A",X"3A",
		X"07",X"62",X"E6",X"80",X"07",X"A7",X"20",X"02",X"3E",X"02",X"32",X"9F",X"6A",X"AF",X"32",X"88",
		X"6A",X"C9",X"3A",X"15",X"62",X"A7",X"28",X"2B",X"3A",X"8F",X"60",X"FE",X"29",X"28",X"07",X"3E",
		X"01",X"32",X"8C",X"60",X"18",X"07",X"3E",X"01",X"32",X"82",X"60",X"18",X"16",X"21",X"4F",X"69",
		X"3E",X"F6",X"BE",X"38",X"27",X"34",X"34",X"21",X"57",X"69",X"34",X"34",X"3E",X"01",X"32",X"09",
		X"60",X"E1",X"C9",X"AF",X"32",X"8C",X"60",X"32",X"8F",X"60",X"21",X"54",X"69",X"36",X"00",X"21",
		X"63",X"66",X"36",X"00",X"21",X"FC",X"69",X"36",X"00",X"C3",X"DB",X"30",X"3E",X"29",X"32",X"8F",
		X"60",X"3E",X"20",X"32",X"09",X"60",X"21",X"4C",X"69",X"36",X"00",X"21",X"54",X"69",X"36",X"00",
		X"E1",X"C9",X"3A",X"91",X"6A",X"A7",X"C0",X"3A",X"15",X"62",X"A7",X"C0",X"CD",X"78",X"44",X"C9",
		X"3A",X"27",X"62",X"FE",X"04",X"CA",X"1F",X"16",X"FE",X"03",X"CA",X"41",X"16",X"C3",X"1B",X"16",
		X"11",X"07",X"67",X"21",X"2D",X"4F",X"01",X"1C",X"04",X"CD",X"2A",X"12",X"11",X"87",X"67",X"21",
		X"29",X"4F",X"01",X"1C",X"04",X"CD",X"2A",X"12",X"C9",X"3F",X"0E",X"02",X"02",X"41",X"0E",X"02",
		X"02",X"3A",X"27",X"62",X"3D",X"01",X"18",X"E0",X"C8",X"3D",X"01",X"18",X"E8",X"C8",X"3D",X"01",
		X"30",X"F0",X"C8",X"01",X"18",X"F0",X"C9",X"DD",X"7E",X"05",X"FE",X"41",X"38",X"07",X"CD",X"B6",
		X"4F",X"DD",X"66",X"03",X"C9",X"CD",X"77",X"4F",X"DD",X"36",X"02",X"02",X"18",X"F3",X"D9",X"01",
		X"00",X"00",X"DD",X"35",X"05",X"18",X"07",X"D9",X"01",X"00",X"00",X"DD",X"34",X"05",X"CD",X"B6",
		X"4F",X"DD",X"66",X"03",X"C3",X"F9",X"1F",X"DD",X"66",X"03",X"DD",X"7E",X"05",X"C6",X"FA",X"6F",
		X"E5",X"D1",X"C5",X"06",X"01",X"CD",X"D3",X"46",X"C1",X"A7",X"3E",X"10",X"20",X"24",X"DD",X"66",
		X"03",X"DD",X"7E",X"05",X"C6",X"06",X"6F",X"E5",X"D1",X"C5",X"06",X"01",X"CD",X"D3",X"46",X"C1",
		X"A7",X"3E",X"20",X"20",X"0D",X"DD",X"7E",X"0B",X"FE",X"00",X"20",X"02",X"3E",X"20",X"DD",X"77",
		X"02",X"C9",X"DD",X"77",X"0B",X"C9",X"DD",X"7E",X"03",X"C6",X"06",X"67",X"DD",X"6E",X"05",X"E5",
		X"D1",X"C5",X"06",X"01",X"CD",X"D3",X"46",X"C1",X"A7",X"3E",X"02",X"20",X"E5",X"DD",X"7E",X"03",
		X"C6",X"FA",X"67",X"DD",X"6E",X"05",X"E5",X"D1",X"C5",X"06",X"01",X"CD",X"D3",X"46",X"C1",X"A7",
		X"3E",X"04",X"20",X"CE",X"18",X"BF",X"DD",X"E5",X"E5",X"C5",X"D5",X"DD",X"66",X"03",X"DD",X"7E",
		X"05",X"C6",X"01",X"6F",X"CD",X"F0",X"2F",X"7E",X"FE",X"D0",X"38",X"23",X"DD",X"7E",X"05",X"FE",
		X"80",X"38",X"0E",X"FE",X"B0",X"38",X"04",X"FE",X"D8",X"38",X"06",X"DD",X"36",X"02",X"02",X"18",
		X"04",X"DD",X"36",X"02",X"04",X"DD",X"7E",X"05",X"D6",X"01",X"DD",X"77",X"05",X"18",X"04",X"DD",
		X"36",X"02",X"01",X"D1",X"C1",X"E1",X"DD",X"E1",X"C3",X"CE",X"1F",X"E5",X"DD",X"7E",X"0C",X"FE",
		X"00",X"28",X"1B",X"DD",X"7E",X"03",X"FE",X"13",X"28",X"09",X"CD",X"57",X"00",X"E6",X"0F",X"FE",
		X"05",X"38",X"0B",X"DD",X"36",X"02",X"40",X"DD",X"36",X"0E",X"90",X"DD",X"70",X"17",X"E1",X"C9",
		X"E5",X"DD",X"E5",X"D5",X"C5",X"DD",X"66",X"05",X"DD",X"6E",X"03",X"48",X"DD",X"21",X"00",X"67",
		X"11",X"20",X"00",X"06",X"0A",X"DD",X"7E",X"00",X"A7",X"28",X"06",X"DD",X"19",X"10",X"F6",X"18",
		X"2F",X"DD",X"36",X"00",X"01",X"DD",X"36",X"02",X"40",X"DD",X"75",X"03",X"DD",X"74",X"05",X"DD",
		X"36",X"07",X"3F",X"DD",X"36",X"08",X"0D",X"DD",X"36",X"0C",X"01",X"DD",X"36",X"0F",X"02",X"DD",
		X"71",X"17",X"3A",X"29",X"62",X"FE",X"01",X"3E",X"A0",X"28",X"02",X"3E",X"75",X"DD",X"77",X"1E",
		X"C1",X"D1",X"DD",X"E1",X"E1",X"C9",X"3A",X"27",X"62",X"FE",X"04",X"20",X"00",X"DD",X"7E",X"02",
		X"FE",X"01",X"20",X"0F",X"3A",X"27",X"62",X"FE",X"02",X"CA",X"AC",X"1F",X"D9",X"DD",X"34",X"05",
		X"C3",X"E6",X"4F",X"DD",X"7E",X"02",X"FE",X"40",X"20",X"28",X"DD",X"7E",X"1E",X"A7",X"20",X"10",
		X"DD",X"36",X"02",X"01",X"DD",X"36",X"1D",X"00",X"DD",X"36",X"1E",X"00",X"D9",X"C3",X"CE",X"1F",
		X"FE",X"19",X"30",X"1E",X"DD",X"7E",X"03",X"DD",X"86",X"1D",X"DD",X"77",X"03",X"DD",X"35",X"1E",
		X"18",X"EA",X"DD",X"7E",X"02",X"CB",X"67",X"C2",X"5E",X"4F",X"CB",X"6F",X"C2",X"67",X"4F",X"C3",
		X"9D",X"1F",X"FE",X"47",X"20",X"E7",X"18",X"C8",X"3A",X"27",X"62",X"DD",X"34",X"05",X"FE",X"04",
		X"20",X"10",X"DD",X"7E",X"17",X"DD",X"BE",X"05",X"C2",X"CE",X"1F",X"DD",X"36",X"02",X"00",X"C3",
		X"BA",X"21",X"DD",X"7E",X"05",X"FE",X"F4",X"DA",X"CE",X"1F",X"3A",X"27",X"62",X"FE",X"02",X"C2",
		X"C3",X"24",X"DD",X"36",X"05",X"F6",X"DD",X"34",X"11",X"DD",X"7E",X"11",X"FE",X"0A",X"30",X"07",
		X"DD",X"36",X"07",X"5D",X"C3",X"CE",X"1F",X"FE",X"1A",X"30",X"07",X"DD",X"36",X"07",X"5E",X"C3",
		X"CE",X"1F",X"DD",X"36",X"11",X"00",X"C3",X"C3",X"24",X"3A",X"27",X"62",X"FE",X"04",X"DD",X"7E",
		X"07",X"20",X"05",X"EE",X"7F",X"C3",X"DA",X"1F",X"DD",X"7E",X"05",X"FE",X"F6",X"DD",X"7E",X"07",
		X"C2",X"D8",X"1F",X"C3",X"DD",X"1F",X"DD",X"7E",X"05",X"D6",X"06",X"DD",X"77",X"05",X"CD",X"2F",
		X"2A",X"F5",X"DD",X"7E",X"05",X"C6",X"06",X"DD",X"77",X"05",X"F1",X"C9",X"DD",X"36",X"0C",X"03",
		X"C3",X"BA",X"21",X"3A",X"27",X"62",X"FE",X"04",X"DD",X"7E",X"05",X"C2",X"1B",X"21",X"DD",X"7E",
		X"07",X"EE",X"7F",X"C3",X"27",X"21",X"3A",X"27",X"62",X"FE",X"04",X"3E",X"00",X"28",X"02",X"3E",
		X"08",X"85",X"C9",X"3A",X"27",X"62",X"FE",X"04",X"CA",X"2B",X"50",X"78",X"D6",X"05",X"C3",X"75",
		X"21",X"3A",X"27",X"62",X"FE",X"04",X"C2",X"F7",X"47",X"CD",X"77",X"4F",X"E1",X"C3",X"BA",X"21",
		X"C9",X"3A",X"27",X"62",X"FE",X"04",X"7E",X"13",X"12",X"C2",X"7E",X"2D",X"C6",X"07",X"12",X"C3",
		X"7E",X"2D",X"C2",X"03",X"24",X"3A",X"27",X"62",X"FE",X"04",X"C2",X"E5",X"23",X"DD",X"7E",X"07",
		X"EE",X"7F",X"DD",X"77",X"07",X"C3",X"01",X"24",X"3A",X"27",X"62",X"FE",X"04",X"DD",X"7E",X"07",
		X"C2",X"69",X"2D",X"EE",X"7F",X"C3",X"70",X"2D",X"3A",X"27",X"62",X"FE",X"04",X"20",X"13",X"DD",
		X"36",X"07",X"3F",X"DD",X"36",X"08",X"0D",X"DD",X"36",X"0C",X"01",X"DD",X"36",X"15",X"00",X"C3",
		X"15",X"2D",X"DD",X"36",X"07",X"BD",X"C3",X"FA",X"2C",X"DD",X"36",X"07",X"BD",X"DD",X"36",X"09",
		X"04",X"C9",X"3A",X"8D",X"6A",X"A7",X"C2",X"D9",X"2B",X"D5",X"62",X"7B",X"D6",X"03",X"6F",X"CD",
		X"F0",X"2F",X"D1",X"7E",X"FE",X"D0",X"DA",X"FD",X"2B",X"3E",X"00",X"32",X"21",X"62",X"00",X"00",
		X"00",X"C3",X"D9",X"2B",X"DD",X"21",X"00",X"67",X"11",X"20",X"00",X"21",X"B7",X"52",X"06",X"07",
		X"DD",X"36",X"00",X"01",X"DD",X"36",X"0F",X"04",X"78",X"FE",X"04",X"30",X"14",X"DD",X"36",X"0C",
		X"01",X"DD",X"36",X"08",X"0D",X"DD",X"36",X"07",X"3F",X"DD",X"36",X"09",X"02",X"DD",X"36",X"0A",
		X"02",X"7E",X"DD",X"77",X"02",X"23",X"7E",X"DD",X"77",X"03",X"23",X"7E",X"DD",X"77",X"05",X"23",
		X"DD",X"19",X"10",X"CC",X"3A",X"29",X"62",X"FE",X"03",X"D8",X"DD",X"21",X"E0",X"67",X"DD",X"36",
		X"00",X"01",X"DD",X"36",X"03",X"7F",X"DD",X"36",X"05",X"B8",X"DD",X"36",X"07",X"41",X"DD",X"36",
		X"02",X"02",X"DD",X"36",X"0F",X"04",X"C9",X"04",X"68",X"47",X"02",X"60",X"7F",X"04",X"40",X"E0",
		X"04",X"A0",X"A8",X"02",X"90",X"47",X"04",X"70",X"CE",X"02",X"80",X"A7",X"FD",X"77",X"03",X"DD",
		X"7E",X"01",X"A7",X"C8",X"DD",X"34",X"0C",X"DD",X"7E",X"0C",X"FE",X"C3",X"30",X"2A",X"DD",X"7E",
		X"02",X"FD",X"77",X"15",X"DD",X"7E",X"04",X"FD",X"77",X"16",X"DD",X"7E",X"0B",X"FD",X"77",X"14",
		X"DD",X"7E",X"0C",X"FD",X"77",X"17",X"C9",X"AF",X"DD",X"77",X"01",X"FD",X"77",X"14",X"FD",X"77",
		X"15",X"FD",X"77",X"16",X"FD",X"77",X"17",X"C9",X"FE",X"CA",X"30",X"EB",X"FD",X"36",X"15",X"6B",
		X"C9",X"CD",X"13",X"29",X"3E",X"05",X"47",X"32",X"B9",X"63",X"1E",X"00",X"DD",X"21",X"00",X"67",
		X"DD",X"E5",X"E5",X"C5",X"11",X"10",X"00",X"21",X"6C",X"69",X"7E",X"DD",X"77",X"03",X"23",X"23",
		X"23",X"7E",X"DD",X"77",X"05",X"23",X"DD",X"36",X"00",X"01",X"DD",X"36",X"09",X"04",X"DD",X"36",
		X"0A",X"04",X"DD",X"19",X"10",X"E4",X"C1",X"E1",X"DD",X"E1",X"CD",X"13",X"29",X"06",X"05",X"DD",
		X"36",X"00",X"00",X"10",X"FA",X"C9",X"DD",X"21",X"00",X"66",X"11",X"10",X"00",X"21",X"D3",X"65",
		X"06",X"02",X"3A",X"8D",X"6A",X"A7",X"20",X"51",X"DD",X"34",X"0B",X"78",X"FE",X"02",X"20",X"5F",
		X"DD",X"7E",X"0B",X"FE",X"40",X"28",X"07",X"E6",X"07",X"28",X"16",X"C3",X"CF",X"53",X"DD",X"36",
		X"0B",X"00",X"DD",X"34",X"0C",X"DD",X"7E",X"0C",X"FE",X"04",X"C2",X"91",X"53",X"AF",X"DD",X"77",
		X"0C",X"DD",X"7E",X"0C",X"A7",X"CA",X"CF",X"53",X"FE",X"02",X"CA",X"CF",X"53",X"FE",X"01",X"28",
		X"0C",X"DD",X"7E",X"05",X"FE",X"AA",X"28",X"27",X"DD",X"34",X"05",X"18",X"22",X"DD",X"7E",X"05",
		X"FE",X"A5",X"28",X"1B",X"DD",X"35",X"05",X"18",X"16",X"DD",X"7E",X"03",X"C6",X"10",X"4F",X"3A",
		X"03",X"62",X"B9",X"30",X"A3",X"79",X"D6",X"20",X"4F",X"3A",X"03",X"62",X"B9",X"38",X"99",X"7E",
		X"DD",X"77",X"03",X"DD",X"19",X"19",X"05",X"20",X"89",X"DD",X"21",X"00",X"66",X"21",X"44",X"69",
		X"06",X"02",X"DD",X"7E",X"03",X"77",X"23",X"DD",X"7E",X"07",X"77",X"23",X"DD",X"7E",X"08",X"77",
		X"23",X"DD",X"7E",X"05",X"77",X"23",X"DD",X"19",X"10",X"E8",X"C9",X"32",X"B9",X"62",X"3E",X"02",
		X"32",X"80",X"63",X"DD",X"21",X"00",X"64",X"21",X"35",X"54",X"11",X"20",X"00",X"06",X"03",X"7E",
		X"23",X"DD",X"77",X"00",X"7E",X"23",X"DD",X"77",X"0E",X"7E",X"23",X"DD",X"77",X"0F",X"DD",X"19",
		X"10",X"ED",X"3A",X"29",X"62",X"FE",X"03",X"D8",X"DD",X"36",X"00",X"01",X"DD",X"36",X"0E",X"BA",
		X"DD",X"36",X"0F",X"48",X"C9",X"01",X"40",X"70",X"01",X"A0",X"48",X"01",X"D5",X"88",X"C2",X"F8",
		X"26",X"3A",X"0A",X"60",X"FE",X"16",X"C2",X"F6",X"26",X"3E",X"19",X"32",X"35",X"6A",X"3E",X"FF",
		X"C3",X"F8",X"26",X"3A",X"27",X"62",X"FE",X"02",X"C2",X"BA",X"21",X"DD",X"7E",X"03",X"FE",X"98",
		X"DA",X"BA",X"21",X"DD",X"7E",X"05",X"FE",X"48",X"D2",X"BA",X"21",X"DD",X"35",X"03",X"DD",X"34",
		X"05",X"C3",X"BA",X"21",X"7C",X"FE",X"14",X"38",X"05",X"FE",X"CF",X"C3",X"69",X"23",X"3A",X"27",
		X"62",X"B9",X"C2",X"F7",X"47",X"7D",X"FE",X"60",X"DA",X"69",X"23",X"E1",X"C3",X"2F",X"20",X"2A",
		X"43",X"63",X"3A",X"99",X"6A",X"A7",X"20",X"2C",X"E5",X"2C",X"2C",X"2C",X"22",X"95",X"6A",X"D5",
		X"C5",X"FD",X"21",X"80",X"66",X"2D",X"2D",X"2D",X"11",X"10",X"00",X"7E",X"06",X"05",X"FD",X"BE",
		X"03",X"28",X"04",X"FD",X"19",X"10",X"F7",X"FD",X"36",X"01",X"01",X"FD",X"22",X"97",X"6A",X"C1",
		X"D1",X"E1",X"7E",X"C9",X"7E",X"36",X"00",X"C9",X"3A",X"98",X"63",X"A7",X"20",X"08",X"3A",X"05",
		X"62",X"E6",X"FC",X"32",X"05",X"62",X"21",X"07",X"62",X"C9",X"21",X"30",X"6A",X"F5",X"3A",X"94",
		X"6A",X"A7",X"28",X"15",X"3A",X"9C",X"6A",X"06",X"7D",X"1E",X"08",X"3D",X"28",X"0B",X"06",X"7E",
		X"1E",X"15",X"3D",X"28",X"04",X"06",X"7F",X"1E",X"16",X"F1",X"C9",X"06",X"05",X"11",X"10",X"00",
		X"FD",X"21",X"80",X"66",X"FD",X"7E",X"03",X"A7",X"28",X"07",X"FD",X"CB",X"01",X"46",X"C2",X"32",
		X"28",X"FD",X"19",X"10",X"EF",X"C9",X"32",X"99",X"6A",X"32",X"50",X"63",X"C9",X"3E",X"80",X"32",
		X"42",X"63",X"DD",X"22",X"51",X"63",X"16",X"00",X"06",X"0A",X"FD",X"7E",X"03",X"DD",X"BE",X"03",
		X"28",X"04",X"DD",X"19",X"10",X"F7",X"3A",X"9C",X"6A",X"3C",X"32",X"9C",X"6A",X"C9",X"CD",X"2A",
		X"12",X"21",X"53",X"55",X"CD",X"A6",X"11",X"21",X"4C",X"3E",X"11",X"0C",X"6A",X"01",X"10",X"00",
		X"ED",X"B0",X"C9",X"9B",X"18",X"5B",X"60",X"A3",X"83",X"2B",X"60",X"00",X"00",X"3A",X"A0",X"6A",
		X"A7",X"20",X"17",X"CD",X"1C",X"2B",X"08",X"3A",X"8B",X"6A",X"A7",X"20",X"04",X"08",X"C3",X"08",
		X"1C",X"3E",X"00",X"32",X"20",X"62",X"08",X"C3",X"4F",X"1C",X"3E",X"48",X"32",X"05",X"62",X"AF",
		X"32",X"A0",X"6A",X"3E",X"A0",X"32",X"03",X"62",X"C3",X"A6",X"1D",X"3A",X"27",X"62",X"FE",X"02",
		X"C2",X"53",X"20",X"DD",X"34",X"05",X"D9",X"C3",X"5E",X"20",X"3A",X"27",X"62",X"FE",X"02",X"28",
		X"0A",X"DD",X"7E",X"05",X"FE",X"41",X"38",X"07",X"CD",X"77",X"4F",X"DD",X"66",X"03",X"C9",X"CD",
		X"77",X"4F",X"3E",X"02",X"DD",X"77",X"02",X"18",X"F2",X"3A",X"80",X"6A",X"A7",X"16",X"00",X"0E",
		X"01",X"28",X"0B",X"16",X"0C",X"0E",X"02",X"CD",X"CE",X"55",X"0E",X"02",X"16",X"F4",X"3A",X"03",
		X"62",X"82",X"06",X"05",X"21",X"0C",X"6A",X"BE",X"28",X"19",X"5F",X"38",X"03",X"96",X"18",X"02",
		X"7E",X"93",X"FE",X"0C",X"38",X"0D",X"7B",X"2C",X"2C",X"2C",X"2C",X"10",X"EA",X"16",X"F4",X"0D",
		X"20",X"DC",X"C9",X"D5",X"3A",X"80",X"6A",X"A7",X"28",X"1A",X"7A",X"B7",X"3A",X"07",X"62",X"16",
		X"F9",X"FA",X"0C",X"56",X"E6",X"80",X"20",X"1F",X"16",X"FD",X"18",X"1B",X"E6",X"80",X"28",X"17",
		X"16",X"FD",X"18",X"13",X"16",X"FD",X"3A",X"05",X"62",X"82",X"2C",X"D1",X"CD",X"4B",X"56",X"28",
		X"17",X"2D",X"2D",X"2D",X"D5",X"16",X"05",X"3A",X"05",X"62",X"82",X"2C",X"D1",X"CD",X"4B",X"56",
		X"7B",X"28",X"05",X"05",X"C8",X"2C",X"18",X"9F",X"2D",X"2D",X"2D",X"22",X"43",X"63",X"3E",X"02",
		X"32",X"42",X"63",X"3D",X"32",X"40",X"63",X"32",X"94",X"6A",X"C9",X"C5",X"E6",X"F8",X"F6",X"03",
		X"47",X"2C",X"2C",X"7E",X"E6",X"F8",X"F6",X"03",X"B8",X"C1",X"C9",X"3A",X"29",X"62",X"3C",X"C9",
		X"21",X"00",X"63",X"ED",X"B1",X"C0",X"E5",X"C5",X"01",X"14",X"00",X"09",X"0C",X"5F",X"7A",X"BE",
		X"28",X"12",X"09",X"BE",X"20",X"09",X"E5",X"CD",X"57",X"00",X"E1",X"E6",X"01",X"28",X"0E",X"7B",
		X"C1",X"E1",X"18",X"DF",X"09",X"3E",X"01",X"C1",X"46",X"E1",X"C3",X"60",X"33",X"AF",X"ED",X"42",
		X"C1",X"46",X"E1",X"C3",X"99",X"33",X"CD",X"9D",X"56",X"3A",X"0F",X"62",X"C9",X"3A",X"0F",X"62",
		X"CB",X"57",X"C8",X"3A",X"4D",X"69",X"E6",X"7F",X"FE",X"08",X"20",X"0E",X"3A",X"4D",X"69",X"EE",
		X"01",X"32",X"4D",X"69",X"C6",X"64",X"32",X"55",X"69",X"C9",X"FE",X"09",X"C0",X"3A",X"4F",X"69",
		X"CB",X"47",X"C0",X"18",X"E7",X"DD",X"36",X"00",X"00",X"DD",X"36",X"02",X"01",X"C9",X"3A",X"05",
		X"60",X"FE",X"01",X"28",X"1D",X"3A",X"29",X"62",X"FE",X"05",X"30",X"06",X"DD",X"7E",X"02",X"A7",
		X"20",X"10",X"DD",X"36",X"00",X"01",X"DD",X"36",X"18",X"01",X"DD",X"36",X"07",X"3D",X"DD",X"36",
		X"08",X"0E",X"AF",X"C3",X"A4",X"31",X"4F",X"7D",X"FE",X"CB",X"28",X"07",X"FE",X"C7",X"28",X"03",
		X"C3",X"62",X"2D",X"F5",X"3A",X"27",X"62",X"FE",X"04",X"3A",X"35",X"6A",X"20",X"0F",X"EE",X"01",
		X"32",X"35",X"6A",X"3A",X"3D",X"6A",X"EE",X"0F",X"32",X"3D",X"6A",X"18",X"05",X"EE",X"03",X"32",
		X"35",X"6A",X"F1",X"FE",X"CB",X"CA",X"8C",X"2D",X"C3",X"62",X"2D",X"7E",X"A7",X"CA",X"40",X"00",
		X"79",X"86",X"77",X"C3",X"40",X"00",X"11",X"04",X"00",X"CD",X"3B",X"00",X"3A",X"0A",X"60",X"FE",
		X"16",X"C0",X"3A",X"27",X"62",X"FE",X"03",X"3A",X"10",X"69",X"20",X"14",X"AF",X"32",X"00",X"69",
		X"32",X"04",X"69",X"32",X"20",X"69",X"32",X"24",X"69",X"32",X"28",X"69",X"32",X"2C",X"69",X"C9",
		X"81",X"32",X"00",X"69",X"32",X"04",X"69",X"3A",X"34",X"6A",X"81",X"32",X"34",X"6A",X"21",X"35",
		X"6A",X"3E",X"0D",X"32",X"3A",X"6A",X"3A",X"A3",X"63",X"A7",X"C8",X"7E",X"EE",X"0E",X"77",X"2C",
		X"36",X"00",X"2C",X"36",X"40",X"C9",X"3A",X"9E",X"6A",X"A7",X"28",X"09",X"11",X"99",X"57",X"21",
		X"CC",X"63",X"CD",X"F4",X"21",X"3A",X"16",X"62",X"C9",X"04",X"60",X"04",X"A0",X"02",X"21",X"B4",
		X"62",X"35",X"7E",X"A7",X"28",X"06",X"FE",X"10",X"CC",X"B7",X"57",X"C9",X"3E",X"03",X"32",X"96",
		X"63",X"CD",X"B7",X"57",X"C3",X"D3",X"2F",X"3A",X"35",X"6A",X"EE",X"03",X"32",X"35",X"6A",X"C9",
		X"CD",X"4E",X"00",X"3E",X"40",X"32",X"37",X"6A",X"3E",X"38",X"32",X"34",X"6A",X"3A",X"27",X"62",
		X"FE",X"03",X"C8",X"FE",X"04",X"28",X"07",X"3E",X"4C",X"32",X"34",X"6A",X"18",X"1C",X"3E",X"50",
		X"32",X"34",X"6A",X"3E",X"38",X"32",X"37",X"6A",X"3E",X"99",X"32",X"35",X"6A",X"E5",X"21",X"0B",
		X"58",X"11",X"3C",X"6A",X"01",X"04",X"00",X"ED",X"B0",X"E1",X"E5",X"21",X"38",X"6A",X"36",X"6B",
		X"2C",X"36",X"5F",X"2C",X"36",X"0D",X"2C",X"36",X"18",X"E1",X"C9",X"5C",X"48",X"00",X"38",X"32",
		X"A0",X"62",X"3A",X"3B",X"6A",X"FE",X"20",X"C8",X"3E",X"20",X"32",X"3B",X"6A",X"3E",X"40",X"32",
		X"38",X"6A",X"C9",X"FE",X"0F",X"D2",X"3D",X"23",X"3A",X"27",X"62",X"FE",X"02",X"CA",X"3D",X"23",
		X"C9",X"3A",X"8B",X"6A",X"A7",X"C2",X"79",X"4D",X"3A",X"10",X"60",X"CB",X"7F",X"CA",X"E2",X"1A",
		X"F5",X"AF",X"32",X"A2",X"6A",X"F1",X"C3",X"E2",X"1A",X"3A",X"27",X"62",X"3D",X"3A",X"00",X"62",
		X"C0",X"06",X"01",X"DD",X"21",X"60",X"66",X"21",X"FC",X"69",X"11",X"10",X"00",X"CD",X"D3",X"11",
		X"3A",X"00",X"62",X"C9",X"3A",X"8B",X"6A",X"A7",X"C0",X"3A",X"98",X"63",X"A7",X"C0",X"3A",X"15",
		X"62",X"C3",X"88",X"2A",X"32",X"16",X"62",X"32",X"89",X"6A",X"32",X"8A",X"6A",X"32",X"88",X"6A",
		X"32",X"87",X"6A",X"C9",X"3E",X"54",X"32",X"8A",X"6A",X"3A",X"20",X"62",X"C9",X"32",X"05",X"62",
		X"3A",X"88",X"6A",X"A7",X"CA",X"E5",X"29",X"3A",X"05",X"62",X"D6",X"04",X"32",X"05",X"62",X"C3",
		X"E5",X"29",X"3A",X"8B",X"6A",X"A7",X"3E",X"04",X"32",X"1E",X"62",X"CA",X"68",X"1C",X"3E",X"01",
		X"32",X"1E",X"62",X"C3",X"68",X"1C",X"3A",X"91",X"6A",X"A7",X"CA",X"38",X"1B",X"3A",X"0F",X"62",
		X"FE",X"08",X"28",X"07",X"3D",X"32",X"0F",X"62",X"C3",X"A6",X"1D",X"3A",X"92",X"6A",X"32",X"07",
		X"62",X"AF",X"32",X"91",X"6A",X"3C",X"32",X"80",X"6A",X"C3",X"A6",X"1D",X"DD",X"7E",X"10",X"A7",
		X"20",X"23",X"3A",X"8A",X"6A",X"FE",X"50",X"01",X"10",X"FF",X"28",X"18",X"FE",X"51",X"01",X"10",
		X"FF",X"28",X"11",X"FE",X"52",X"01",X"10",X"FF",X"28",X"0A",X"FE",X"53",X"01",X"10",X"FF",X"28",
		X"03",X"01",X"00",X"00",X"09",X"DD",X"74",X"05",X"C9",X"C5",X"3A",X"29",X"62",X"47",X"3E",X"40",
		X"D6",X"05",X"FE",X"2A",X"38",X"02",X"10",X"F8",X"C1",X"21",X"A4",X"6A",X"BE",X"D0",X"36",X"00",
		X"DD",X"36",X"00",X"01",X"C9",X"DD",X"21",X"D0",X"65",X"21",X"A3",X"63",X"11",X"6A",X"3A",X"3A",
		X"29",X"62",X"FE",X"03",X"38",X"27",X"11",X"63",X"40",X"18",X"22",X"DD",X"21",X"B0",X"65",X"21",
		X"A4",X"63",X"11",X"80",X"60",X"3A",X"29",X"62",X"FE",X"03",X"38",X"11",X"11",X"7A",X"6F",X"18",
		X"0C",X"DD",X"21",X"C0",X"65",X"21",X"A6",X"63",X"11",X"A5",X"89",X"18",X"00",X"CD",X"6C",X"59",
		X"3E",X"00",X"20",X"06",X"CD",X"7A",X"59",X"DD",X"7E",X"0C",X"77",X"C9",X"DD",X"34",X"0D",X"DD",
		X"7E",X"0D",X"FE",X"04",X"C0",X"DD",X"36",X"0D",X"00",X"C9",X"7A",X"DD",X"BE",X"03",X"3E",X"01",
		X"28",X"08",X"7B",X"DD",X"BE",X"03",X"3E",X"FF",X"20",X"03",X"DD",X"77",X"0C",X"C9",X"CD",X"1C",
		X"01",X"21",X"30",X"69",X"01",X"02",X"00",X"AF",X"77",X"23",X"10",X"FC",X"0D",X"20",X"F9",X"C9",
		X"00",X"12",X"00",X"00",X"16",X"00",X"00",X"00",X"CD",X"E0",X"5F",X"A7",X"CA",X"63",X"1B",X"C3",
		X"A6",X"1D",X"21",X"0A",X"60",X"3A",X"9E",X"6A",X"A7",X"C8",X"E1",X"C9",X"FE",X"03",X"C0",X"11",
		X"74",X"5A",X"1A",X"B7",X"C8",X"32",X"B3",X"63",X"13",X"1A",X"6F",X"13",X"1A",X"67",X"0E",X"B2",
		X"CD",X"87",X"5A",X"D5",X"3A",X"B3",X"63",X"FE",X"05",X"30",X"11",X"E6",X"01",X"0E",X"B3",X"11",
		X"E0",X"FF",X"28",X"05",X"0E",X"BB",X"11",X"20",X"00",X"CD",X"94",X"5A",X"D1",X"13",X"18",X"D2",
		X"CD",X"13",X"29",X"C9",X"F5",X"D9",X"DD",X"E5",X"CD",X"00",X"5A",X"DD",X"E1",X"D9",X"F1",X"C9",
		X"DD",X"77",X"05",X"21",X"B8",X"69",X"DD",X"21",X"A0",X"65",X"06",X"06",X"11",X"10",X"00",X"F5",
		X"DD",X"E5",X"CD",X"D3",X"11",X"DD",X"E1",X"F1",X"C9",X"F5",X"D9",X"3D",X"4F",X"06",X"00",X"21",
		X"B0",X"6A",X"09",X"36",X"01",X"87",X"4F",X"21",X"34",X"5A",X"09",X"5E",X"23",X"56",X"EB",X"36",
		X"00",X"D9",X"F1",X"C9",X"20",X"69",X"24",X"69",X"28",X"69",X"2C",X"69",X"00",X"69",X"04",X"69",
		X"3A",X"B3",X"63",X"4F",X"11",X"74",X"5A",X"1A",X"B7",X"C8",X"B9",X"28",X"05",X"13",X"13",X"13",
		X"18",X"F5",X"32",X"B3",X"63",X"13",X"1A",X"6F",X"13",X"1A",X"67",X"0E",X"EC",X"CD",X"87",X"5A",
		X"3A",X"B3",X"63",X"FE",X"05",X"D0",X"E6",X"01",X"11",X"E0",X"FF",X"28",X"03",X"11",X"20",X"00",
		X"CD",X"94",X"5A",X"C9",X"05",X"C8",X"75",X"06",X"28",X"76",X"03",X"68",X"75",X"04",X"88",X"76",
		X"01",X"A8",X"74",X"02",X"48",X"77",X"00",X"D5",X"E5",X"79",X"06",X"03",X"77",X"23",X"3D",X"10",
		X"FB",X"E1",X"D1",X"C9",X"19",X"79",X"77",X"EE",X"07",X"4F",X"3A",X"B3",X"63",X"FE",X"03",X"D0",
		X"E6",X"01",X"1B",X"06",X"03",X"19",X"79",X"77",X"EE",X"07",X"19",X"23",X"77",X"EE",X"07",X"4F",
		X"10",X"F3",X"C9",X"3E",X"04",X"F7",X"FD",X"21",X"00",X"62",X"DD",X"21",X"A0",X"65",X"06",X"06",
		X"78",X"32",X"B9",X"63",X"11",X"10",X"00",X"C5",X"CD",X"F0",X"59",X"A7",X"20",X"0D",X"C1",X"AF",
		X"32",X"9D",X"6A",X"DD",X"77",X"01",X"DD",X"19",X"10",X"F9",X"C9",X"3A",X"B9",X"63",X"4F",X"78",
		X"91",X"28",X"05",X"DD",X"19",X"04",X"18",X"F3",X"C1",X"DD",X"36",X"01",X"01",X"3A",X"10",X"60",
		X"1F",X"D8",X"1F",X"D8",X"1F",X"38",X"35",X"1F",X"30",X"20",X"DD",X"7E",X"0F",X"A7",X"20",X"1A",
		X"DD",X"36",X"02",X"00",X"3A",X"05",X"62",X"C6",X"10",X"FE",X"E2",X"38",X"02",X"3E",X"E2",X"CD",
		X"F4",X"59",X"FE",X"E2",X"38",X"10",X"DD",X"36",X"0F",X"01",X"AF",X"32",X"0F",X"62",X"DD",X"36",
		X"01",X"00",X"3C",X"32",X"9D",X"6A",X"DD",X"19",X"05",X"20",X"95",X"C9",X"AF",X"32",X"9D",X"6A",
		X"DD",X"77",X"0F",X"3C",X"DD",X"77",X"02",X"3A",X"05",X"62",X"D6",X"10",X"CD",X"F4",X"59",X"FE",
		X"5B",X"30",X"E3",X"3A",X"90",X"62",X"3D",X"32",X"90",X"62",X"E5",X"DD",X"E5",X"E1",X"7D",X"D6",
		X"A0",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"3C",X"32",X"B3",X"63",X"CD",X"19",X"5A",X"D9",X"3E",
		X"03",X"32",X"03",X"7D",X"32",X"83",X"60",X"CD",X"40",X"5A",X"D9",X"C5",X"3A",X"B3",X"63",X"3D",
		X"87",X"87",X"4F",X"06",X"00",X"21",X"B8",X"69",X"09",X"22",X"43",X"63",X"3E",X"04",X"32",X"42",
		X"63",X"3E",X"01",X"32",X"40",X"63",X"32",X"A1",X"6A",X"C1",X"E1",X"DD",X"36",X"08",X"07",X"DD",
		X"36",X"05",X"52",X"DD",X"E5",X"D9",X"CD",X"03",X"5A",X"D9",X"DD",X"E1",X"C9",X"21",X"35",X"6A",
		X"7E",X"1F",X"3E",X"02",X"1F",X"47",X"AE",X"77",X"2C",X"78",X"E6",X"80",X"AE",X"77",X"C9",X"3A",
		X"29",X"62",X"FE",X"01",X"3E",X"03",X"28",X"0B",X"3A",X"29",X"62",X"FE",X"02",X"3E",X"04",X"28",
		X"02",X"3E",X"05",X"E5",X"21",X"A1",X"63",X"BE",X"E1",X"CA",X"6A",X"31",X"C3",X"84",X"31",X"3A",
		X"AA",X"63",X"A7",X"20",X"05",X"23",X"7E",X"23",X"18",X"05",X"34",X"23",X"34",X"7E",X"23",X"FE",
		X"FE",X"30",X"03",X"FE",X"09",X"C9",X"2B",X"36",X"FE",X"2B",X"36",X"FE",X"23",X"23",X"C9",X"11",
		X"FE",X"5B",X"21",X"8F",X"76",X"CD",X"65",X"0B",X"3E",X"01",X"32",X"80",X"6A",X"C9",X"1B",X"15",
		X"15",X"20",X"10",X"17",X"1F",X"19",X"1E",X"17",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",X"24",X"1F",
		X"10",X"1D",X"11",X"22",X"19",X"1F",X"3A",X"23",X"10",X"18",X"19",X"14",X"15",X"1F",X"25",X"24",
		X"AA",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"01",X"02",X"01",X"00",X"00",X"FE",
		X"FE",X"FE",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"01",X"01",X"01",X"02",X"02",X"02",X"AA",X"18",
		X"69",X"08",X"69",X"0C",X"6A",X"18",X"6A",X"14",X"69",X"10",X"69",X"10",X"6A",X"1C",X"6A",X"1C",
		X"69",X"0C",X"69",X"14",X"6A",X"20",X"6A",X"1B",X"15",X"15",X"20",X"10",X"17",X"1F",X"19",X"1E",
		X"17",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",X"24",X"1F",X"10",X"1D",X"11",X"22",X"19",X"1F",X"3A",
		X"23",X"10",X"18",X"19",X"14",X"15",X"1F",X"25",X"24",X"AA",X"12",X"15",X"10",X"13",X"11",X"22",
		X"15",X"16",X"25",X"1C",X"10",X"39",X"AA",X"F5",X"3A",X"27",X"62",X"FE",X"04",X"28",X"07",X"F1",
		X"CD",X"6D",X"21",X"C3",X"BA",X"21",X"F1",X"DD",X"7E",X"0C",X"A7",X"CA",X"BA",X"21",X"DD",X"7E",
		X"02",X"E6",X"06",X"CA",X"BA",X"21",X"DD",X"66",X"03",X"DD",X"7E",X"05",X"D6",X"04",X"6F",X"CD",
		X"F0",X"2F",X"7E",X"FE",X"F7",X"20",X"25",X"DD",X"7E",X"05",X"FE",X"60",X"30",X"18",X"DD",X"7E",
		X"03",X"FE",X"4A",X"38",X"11",X"CD",X"57",X"00",X"E6",X"01",X"20",X"02",X"18",X"3B",X"CD",X"57",
		X"00",X"E6",X"01",X"C2",X"BA",X"21",X"DD",X"36",X"02",X"01",X"18",X"00",X"3A",X"29",X"62",X"C3",
		X"E7",X"5F",X"3A",X"05",X"62",X"FE",X"A0",X"D2",X"BA",X"21",X"3A",X"29",X"62",X"FE",X"05",X"0E",
		X"40",X"38",X"02",X"0E",X"20",X"3A",X"05",X"62",X"81",X"DD",X"BE",X"05",X"D2",X"BA",X"21",X"AF",
		X"DD",X"77",X"00",X"DD",X"77",X"03",X"C3",X"BA",X"21",X"3A",X"05",X"62",X"FE",X"90",X"30",X"BE",
		X"CD",X"50",X"50",X"C3",X"BA",X"21",X"3E",X"40",X"32",X"41",X"63",X"3E",X"02",X"32",X"40",X"63",
		X"3A",X"31",X"6A",X"FE",X"7A",X"20",X"0B",X"21",X"30",X"6A",X"11",X"28",X"6A",X"01",X"04",X"00",
		X"ED",X"B0",X"3A",X"42",X"63",X"1F",X"DA",X"70",X"3E",X"1F",X"DA",X"58",X"5D",X"1F",X"DA",X"4A",
		X"5D",X"16",X"00",X"A7",X"C8",X"CD",X"DA",X"54",X"18",X"05",X"06",X"7A",X"11",X"02",X"00",X"CD",
		X"9F",X"30",X"2A",X"43",X"63",X"7E",X"18",X"10",X"21",X"85",X"60",X"36",X"03",X"06",X"7C",X"11",
		X"04",X"00",X"CD",X"9F",X"30",X"CD",X"8F",X"54",X"2C",X"2C",X"2C",X"4E",X"F5",X"3A",X"A1",X"6A",
		X"F5",X"AF",X"32",X"A1",X"6A",X"F1",X"A7",X"28",X"04",X"3E",X"10",X"81",X"4F",X"F1",X"C3",X"36",
		X"1E",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",X"01",
		X"00",X"01",X"00",X"01",X"00",X"01",X"01",X"01",X"00",X"00",X"77",X"7A",X"77",X"77",X"AA",X"DB",
		X"33",X"09",X"D8",X"EB",X"32",X"09",X"D8",X"DB",X"35",X"09",X"E8",X"EB",X"34",X"09",X"E8",X"DD",
		X"36",X"11",X"00",X"DD",X"36",X"12",X"00",X"21",X"00",X"63",X"ED",X"B1",X"28",X"3E",X"DD",X"7E",
		X"11",X"A7",X"20",X"0C",X"DD",X"7E",X"12",X"A7",X"C8",X"DD",X"7E",X"12",X"47",X"C3",X"99",X"33",
		X"DD",X"7E",X"12",X"A7",X"20",X"07",X"DD",X"7E",X"11",X"47",X"C3",X"60",X"33",X"3A",X"05",X"62",
		X"C6",X"08",X"47",X"DD",X"7E",X"0F",X"90",X"30",X"E0",X"78",X"D6",X"10",X"47",X"DD",X"7E",X"0F",
		X"90",X"38",X"E3",X"DD",X"36",X"11",X"00",X"DD",X"36",X"12",X"00",X"C9",X"E5",X"C5",X"01",X"14",
		X"00",X"09",X"0C",X"5F",X"7A",X"BE",X"20",X"07",X"E5",X"09",X"7E",X"DD",X"77",X"11",X"E1",X"7A",
		X"09",X"BE",X"20",X"09",X"E5",X"AF",X"ED",X"42",X"7E",X"DD",X"77",X"12",X"E1",X"7B",X"C1",X"E1",
		X"C3",X"BA",X"5D",X"43",X"1C",X"0C",X"A3",X"BB",X"1C",X"0C",X"A3",X"43",X"A3",X"BB",X"A3",X"00",
		X"00",X"00",X"00",X"00",X"00",X"D3",X"D8",X"2B",X"D8",X"A3",X"D8",X"5B",X"D8",X"8B",X"D8",X"73",
		X"D8",X"5F",X"8D",X"02",X"02",X"3A",X"85",X"63",X"EF",X"4F",X"5E",X"E9",X"5E",X"EF",X"5E",X"21",
		X"F0",X"6A",X"34",X"7E",X"FE",X"01",X"20",X"08",X"21",X"81",X"5D",X"22",X"F1",X"6A",X"18",X"40",
		X"FE",X"40",X"38",X"3C",X"DD",X"21",X"34",X"6A",X"DD",X"34",X"00",X"DD",X"7E",X"00",X"FE",X"F0",
		X"20",X"23",X"3E",X"30",X"32",X"09",X"60",X"AF",X"32",X"80",X"6A",X"32",X"81",X"6A",X"32",X"83",
		X"6A",X"3E",X"1E",X"32",X"35",X"6A",X"21",X"85",X"63",X"34",X"3E",X"E0",X"32",X"37",X"6A",X"3E",
		X"F8",X"32",X"34",X"6A",X"C9",X"CB",X"57",X"3E",X"96",X"20",X"02",X"3E",X"95",X"DD",X"77",X"01",
		X"21",X"F4",X"6A",X"34",X"7E",X"FE",X"01",X"C0",X"36",X"00",X"2A",X"F1",X"6A",X"7E",X"FE",X"AA",
		X"28",X"A6",X"FE",X"77",X"28",X"09",X"FE",X"7A",X"20",X"0A",X"3E",X"03",X"32",X"82",X"60",X"23",
		X"22",X"F1",X"6A",X"C9",X"23",X"22",X"F1",X"6A",X"4F",X"21",X"4F",X"69",X"86",X"77",X"32",X"57",
		X"69",X"21",X"4C",X"69",X"7E",X"FE",X"F7",X"30",X"05",X"34",X"21",X"54",X"69",X"34",X"21",X"0B",
		X"69",X"FF",X"21",X"08",X"69",X"0E",X"01",X"FF",X"C9",X"DF",X"21",X"85",X"63",X"34",X"C9",X"21",
		X"34",X"6A",X"7E",X"FE",X"EE",X"30",X"1B",X"3A",X"A3",X"6A",X"A7",X"20",X"15",X"3E",X"01",X"32",
		X"A3",X"6A",X"CD",X"B7",X"5F",X"E5",X"21",X"9F",X"5D",X"11",X"08",X"69",X"01",X"10",X"00",X"ED",
		X"B0",X"E1",X"3A",X"83",X"6A",X"A7",X"CA",X"6F",X"5F",X"FE",X"02",X"28",X"2E",X"35",X"CB",X"46",
		X"C8",X"2A",X"84",X"6A",X"4E",X"23",X"22",X"84",X"6A",X"3E",X"AA",X"B9",X"28",X"0D",X"3A",X"37",
		X"6A",X"81",X"32",X"37",X"6A",X"FE",X"EE",X"D8",X"C3",X"B7",X"5F",X"3E",X"17",X"32",X"35",X"6A",
		X"3E",X"02",X"32",X"83",X"6A",X"3E",X"00",X"32",X"36",X"6A",X"C9",X"35",X"7E",X"28",X"0C",X"E6",
		X"03",X"C0",X"3A",X"35",X"6A",X"EE",X"0E",X"32",X"35",X"6A",X"C9",X"AF",X"32",X"85",X"63",X"2A",
		X"2A",X"62",X"7E",X"32",X"27",X"62",X"21",X"09",X"60",X"36",X"40",X"23",X"36",X"0A",X"C9",X"35",
		X"7E",X"FE",X"C0",X"06",X"03",X"28",X"0C",X"FE",X"B0",X"06",X"06",X"28",X"06",X"FE",X"A0",X"06",
		X"09",X"20",X"09",X"78",X"32",X"81",X"6A",X"3E",X"03",X"32",X"82",X"6A",X"21",X"82",X"6A",X"35",
		X"4E",X"20",X"02",X"36",X"03",X"06",X"00",X"3A",X"81",X"6A",X"81",X"4F",X"CD",X"BD",X"5F",X"21",
		X"21",X"5C",X"09",X"7E",X"21",X"37",X"6A",X"86",X"77",X"FE",X"EE",X"D8",X"21",X"2F",X"5C",X"22",
		X"84",X"6A",X"3E",X"01",X"32",X"83",X"6A",X"3E",X"03",X"32",X"82",X"60",X"C9",X"F5",X"C5",X"3A",
		X"34",X"6A",X"E6",X"03",X"CC",X"9D",X"5B",X"C1",X"F1",X"C9",X"06",X"09",X"C8",X"06",X"0A",X"C9",
		X"3E",X"09",X"C8",X"3E",X"0A",X"C9",X"3D",X"32",X"29",X"62",X"3C",X"C9",X"00",X"00",X"00",X"00",
		X"21",X"07",X"62",X"3A",X"15",X"62",X"C9",X"3D",X"CA",X"BA",X"21",X"C3",X"E2",X"5C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
