library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity VICTORY_1K is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of VICTORY_1K is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"7C",X"82",X"82",X"82",X"82",X"7C",X"00",X"00",X"02",X"02",X"FE",X"42",X"02",X"00",X"00",
		X"00",X"62",X"92",X"8A",X"86",X"86",X"42",X"00",X"00",X"8C",X"D2",X"B2",X"92",X"82",X"84",X"00",
		X"00",X"08",X"FE",X"48",X"28",X"18",X"08",X"00",X"00",X"1C",X"A2",X"A2",X"A2",X"A6",X"E4",X"00",
		X"00",X"8C",X"92",X"92",X"92",X"52",X"3C",X"00",X"00",X"C0",X"A0",X"90",X"8E",X"80",X"80",X"00",
		X"00",X"6C",X"92",X"92",X"92",X"92",X"6C",X"00",X"00",X"7C",X"92",X"92",X"92",X"92",X"60",X"00",
		X"3F",X"7F",X"FF",X"3F",X"3F",X"0E",X"0E",X"0C",X"08",X"0C",X"3E",X"3E",X"0F",X"0F",X"3F",X"3F",
		X"FF",X"FF",X"FF",X"E7",X"E7",X"FF",X"FF",X"FF",X"E7",X"BD",X"DB",X"7E",X"7E",X"DB",X"BD",X"E7",
		X"40",X"20",X"10",X"08",X"04",X"02",X"00",X"00",X"00",X"00",X"00",X"30",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",
		X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",X"44",X"C6",X"82",X"82",X"C6",X"7C",X"38",X"00",
		X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",X"82",X"92",X"92",X"92",X"FE",X"FE",X"00",X"00",
		X"80",X"90",X"90",X"90",X"90",X"FE",X"FE",X"00",X"9E",X"9E",X"92",X"82",X"C6",X"7C",X"38",X"00",
		X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",X"82",X"82",X"FE",X"FE",X"82",X"82",X"00",X"00",
		X"FC",X"FE",X"02",X"02",X"02",X"06",X"04",X"00",X"82",X"C6",X"6E",X"3C",X"18",X"FE",X"FE",X"00",
		X"02",X"02",X"02",X"02",X"FE",X"FE",X"00",X"00",X"FE",X"FE",X"70",X"38",X"70",X"FE",X"FE",X"00",
		X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",X"00",
		X"70",X"F8",X"88",X"88",X"88",X"FE",X"FE",X"00",X"7A",X"FC",X"8E",X"8A",X"82",X"FE",X"7C",X"00",
		X"72",X"F6",X"9E",X"8C",X"88",X"FE",X"FE",X"00",X"0C",X"5E",X"D2",X"92",X"92",X"F6",X"64",X"00",
		X"80",X"80",X"FE",X"FE",X"80",X"80",X"00",X"00",X"FC",X"FE",X"02",X"02",X"02",X"FE",X"FC",X"00",
		X"F0",X"F8",X"1C",X"0E",X"1C",X"F8",X"F0",X"00",X"F8",X"FE",X"1C",X"38",X"1C",X"FE",X"F8",X"00",
		X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",X"C0",X"F0",X"1E",X"1E",X"F0",X"C0",X"00",X"00",
		X"C2",X"E2",X"F2",X"BA",X"9E",X"8E",X"86",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"00",
		X"18",X"42",X"24",X"81",X"81",X"24",X"42",X"18",X"0D",X"53",X"31",X"19",X"08",X"04",X"F2",X"00",
		X"3C",X"42",X"A5",X"A5",X"A5",X"99",X"42",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"42",X"00",X"02",X"80",X"00",X"00",X"02",X"00",X"58",X"94",X"84",
		X"10",X"07",X"00",X"3C",X"50",X"97",X"50",X"3C",X"84",X"78",X"82",X"40",X"90",X"02",X"40",X"00",
		X"FF",X"FF",X"FF",X"C0",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"CF",X"C7",X"E3",X"F1",X"F8",X"FD",
		X"FF",X"F3",X"F3",X"F3",X"F9",X"F9",X"F9",X"FF",X"FF",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"FF",
		X"FF",X"FF",X"FF",X"C0",X"C0",X"FF",X"FF",X"FF",X"FD",X"F8",X"F1",X"E3",X"C7",X"CF",X"FF",X"FF",
		X"FF",X"F9",X"F9",X"F9",X"F3",X"F3",X"F3",X"FF",X"FF",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"FF",
		X"FF",X"FF",X"F9",X"F0",X"F0",X"F9",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",
		X"BE",X"E3",X"A1",X"CD",X"C2",X"F1",X"E7",X"FF",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"03",X"00",X"00",X"00",X"00",X"40",X"40",X"00",X"C0",X"00",X"00",X"00",X"00",X"02",X"02",
		X"40",X"40",X"00",X"00",X"00",X"00",X"03",X"00",X"02",X"02",X"00",X"00",X"00",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",
		X"03",X"03",X"01",X"0E",X"1C",X"08",X"00",X"00",X"E0",X"D0",X"30",X"70",X"F0",X"F0",X"70",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"40",X"40",
		X"00",X"01",X"03",X"07",X"07",X"00",X"00",X"00",X"40",X"40",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",
		X"01",X"03",X"01",X"01",X"01",X"01",X"00",X"00",X"FC",X"FC",X"F8",X"F0",X"F0",X"F8",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"1E",X"1E",X"0F",X"07",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"08",X"0A",X"09",X"08",X"0B",X"03",X"07",X"00",X"80",X"C0",X"80",X"80",X"C0",X"80",X"C0",X"00",
		X"00",X"0F",X"0F",X"0F",X"07",X"03",X"03",X"03",X"00",X"E0",X"E0",X"E0",X"C0",X"80",X"80",X"80",
		X"03",X"03",X"0F",X"07",X"03",X"03",X"01",X"00",X"80",X"80",X"E0",X"C0",X"80",X"80",X"00",X"00",
		X"06",X"07",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"40",X"00",
		X"00",X"00",X"01",X"01",X"02",X"07",X"06",X"07",X"00",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"06",X"07",X"06",X"03",X"01",X"01",X"00",X"00",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FC",X"F8",X"F0",X"F0",X"F0",X"FC",X"FE",X"F0",X"F0",X"E0",X"E0",X"F0",X"F8",X"FC",X"FE",
		X"80",X"C0",X"C0",X"F0",X"F0",X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FC",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"F0",X"F8",X"F0",X"E0",X"E0",X"F0",
		X"80",X"C0",X"E0",X"F0",X"E0",X"E0",X"F0",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FC",X"FC",X"F0",X"F0",X"E0",X"C0",X"00",X"E0",X"E0",X"C0",X"80",X"C0",X"80",X"00",X"00",
		X"00",X"80",X"80",X"C0",X"80",X"C0",X"80",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"1F",X"0F",X"07",X"03",X"01",
		X"01",X"03",X"07",X"0F",X"1F",X"3F",X"7F",X"FF",X"80",X"C0",X"E0",X"F0",X"F8",X"FC",X"FE",X"FF",
		X"FF",X"FE",X"FC",X"F8",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F9",X"F6",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",
		X"EF",X"F6",X"F9",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FC",X"FB",X"F7",X"F7",X"FF",X"FF",X"FF",X"FF",X"3F",X"DF",X"EF",X"EF",
		X"F7",X"F7",X"FB",X"FC",X"FF",X"FF",X"FF",X"FF",X"EF",X"EF",X"DF",X"3F",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FC",X"FB",X"F7",X"EF",X"EF",X"EF",X"FF",X"FF",X"0F",X"F7",X"FB",X"FD",X"DD",X"BD",
		X"EF",X"EF",X"EF",X"F7",X"FB",X"FC",X"FF",X"FF",X"7D",X"FD",X"BD",X"FB",X"F7",X"0F",X"FF",X"FF",
		X"F0",X"EF",X"DF",X"BF",X"3F",X"7F",X"7D",X"7D",X"0F",X"F7",X"FB",X"FD",X"FE",X"FE",X"FE",X"7E",
		X"7F",X"7E",X"7D",X"3F",X"BF",X"DF",X"EF",X"F0",X"FE",X"7E",X"FE",X"FD",X"FB",X"F7",X"EF",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"02",X"0A",X"07",X"00",X"00",X"00",X"00",X"00",X"40",X"80",X"00",
		X"1F",X"07",X"0A",X"02",X"00",X"00",X"00",X"00",X"E0",X"00",X"80",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"09",X"05",X"07",X"27",X"00",X"00",X"00",X"20",X"40",X"00",X"80",X"C0",
		X"17",X"03",X"05",X"09",X"00",X"00",X"00",X"00",X"D0",X"90",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"08",X"00",X"21",X"18",X"1A",X"00",X"10",X"20",X"40",X"00",X"00",X"C8",X"42",
		X"04",X"00",X"02",X"00",X"08",X"11",X"21",X"00",X"5C",X"40",X"48",X"60",X"08",X"04",X"00",X"00",
		X"08",X"08",X"08",X"04",X"14",X"23",X"11",X"12",X"00",X"80",X"84",X"98",X"A0",X"A0",X"00",X"44",
		X"04",X"06",X"06",X"01",X"04",X"10",X"20",X"00",X"62",X"4C",X"70",X"88",X"40",X"44",X"40",X"40");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
