library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity rom4t33 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of rom4t33 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"41",X"9F",X"41",X"BE",X"41",X"DD",X"41",X"FC",X"1A",X"A5",X"1A",X"B8",X"1A",X"D3",X"41",X"80",
		X"3A",X"1A",X"20",X"DB",X"A7",X"CD",X"D2",X"06",X"DC",X"3A",X"CD",X"20",X"06",X"9D",X"29",X"D2",
		X"3A",X"19",X"20",X"FB",X"E6",X"C3",X"00",X"1D",X"1A",X"29",X"1F",X"E6",X"03",X"FE",X"F0",X"DA",
		X"01",X"07",X"F0",X"FF",X"01",X"F0",X"FF",X"01",X"F0",X"00",X"05",X"B0",X"FF",X"07",X"F0",X"F0",
		X"00",X"40",X"FF",X"FF",X"FF",X"FF",X"F8",X"D8",X"E0",X"B0",X"00",X"01",X"E0",X"FF",X"FF",X"40",
		X"F8",X"F8",X"F8",X"FF",X"FF",X"50",X"20",X"70",X"03",X"02",X"F8",X"FF",X"03",X"F8",X"FF",X"00",
		X"FF",X"00",X"7C",X"FF",X"01",X"FC",X"FF",X"01",X"20",X"FF",X"FF",X"00",X"7F",X"FF",X"00",X"00",
		X"38",X"6C",X"38",X"FF",X"FF",X"10",X"00",X"10",X"7C",X"FC",X"00",X"01",X"7C",X"FF",X"FF",X"7C",
		X"FE",X"BE",X"FE",X"FF",X"FF",X"36",X"3E",X"36",X"FF",X"FF",X"00",X"3F",X"00",X"00",X"FF",X"FF",
		X"FF",X"00",X"00",X"FF",X"F8",X"FE",X"1F",X"00",X"3E",X"FF",X"FF",X"1C",X"08",X"1C",X"08",X"FF",
		X"BD",X"EF",X"BF",X"FF",X"FF",X"EA",X"6C",X"AE",X"00",X"00",X"FF",X"00",X"EF",X"FF",X"FF",X"EF",
		X"D2",X"DE",X"01",X"01",X"DE",X"FF",X"01",X"7E",X"6C",X"FF",X"FF",X"28",X"00",X"28",X"FF",X"FF",
		X"01",X"D8",X"FF",X"00",X"50",X"D8",X"50",X"FF",X"FF",X"01",X"DC",X"7E",X"01",X"01",X"DC",X"FF",
		X"FC",X"A4",X"02",X"02",X"FC",X"FF",X"02",X"B8",X"FF",X"00",X"BC",X"FF",X"03",X"BC",X"FF",X"03",
		X"01",X"A0",X"FF",X"00",X"00",X"A0",X"FF",X"FF",X"FF",X"03",X"B0",X"B8",X"01",X"03",X"B0",X"FF",
		X"28",X"CD",X"C3",X"0A",X"17",X"E7",X"FF",X"FF",X"A3",X"3A",X"FE",X"20",X"D2",X"01",X"1E",X"5F",
		X"32",X"F1",X"20",X"DF",X"88",X"CD",X"C3",X"17",X"FF",X"FF",X"FF",X"FF",X"CD",X"FF",X"18",X"8D",
		X"FE",X"1B",X"CA",X"80",X"1B",X"C0",X"8E",X"C3",X"16",X"E6",X"D1",X"3A",X"A7",X"20",X"C0",X"CA",
		X"A7",X"E1",X"10",X"CA",X"FE",X"19",X"CA",X"01",X"E5",X"1B",X"7E",X"24",X"B6",X"23",X"B6",X"23",
		X"67",X"00",X"49",X"C3",X"EB",X"18",X"C3",X"2B",X"19",X"10",X"D6",X"7D",X"6F",X"20",X"DE",X"7C",
		X"18",X"49",X"15",X"FE",X"5C",X"D2",X"FE",X"1B",X"1B",X"DD",X"E6",X"7D",X"FE",X"1F",X"D2",X"19",
		X"C3",X"1B",X"18",X"49",X"25",X"E5",X"23",X"7E",X"D2",X"10",X"18",X"49",X"09",X"FE",X"21",X"DA",
		X"D6",X"7D",X"6F",X"20",X"DE",X"7C",X"67",X"00",X"23",X"B6",X"E1",X"B6",X"C2",X"A7",X"18",X"81",
		X"20",X"D8",X"2D",X"C3",X"3A",X"16",X"20",X"D7",X"49",X"C3",X"32",X"18",X"20",X"D9",X"32",X"97",
		X"CF",X"32",X"C3",X"20",X"05",X"5E",X"0F",X"3E",X"CA",X"A7",X"16",X"2D",X"7D",X"C3",X"3D",X"16",
		X"C3",X"20",X"1B",X"7D",X"06",X"C5",X"11",X"00",X"CF",X"32",X"C3",X"20",X"16",X"5F",X"D5",X"32",
		X"1F",X"1A",X"79",X"12",X"47",X"B0",X"FE",X"7B",X"20",X"B0",X"1A",X"B7",X"12",X"1F",X"13",X"4F",
		X"C1",X"78",X"C0",X"A7",X"C3",X"2B",X"17",X"CC",X"CA",X"BF",X"1B",X"B8",X"C3",X"13",X"1B",X"A2",
		X"EB",X"77",X"23",X"23",X"23",X"23",X"3C",X"7E",X"08",X"3E",X"90",X"C3",X"00",X"1B",X"03",X"3E",
		X"77",X"23",X"D6",X"7D",X"6F",X"0A",X"00",X"00",X"70",X"23",X"71",X"23",X"72",X"23",X"73",X"23",
		X"32",X"05",X"22",X"00",X"81",X"C9",X"0F",X"E6",X"C2",X"A7",X"19",X"26",X"00",X"3A",X"C6",X"22",
		X"32",X"0F",X"20",X"ED",X"21",X"C3",X"00",X"1B",X"12",X"4F",X"ED",X"3A",X"3C",X"20",X"E6",X"3C",
		X"12",X"D8",X"10",X"D8",X"0F",X"D8",X"11",X"D8",X"1A",X"88",X"1A",X"6B",X"1A",X"4E",X"1A",X"31",
		X"42",X"C2",X"3A",X"1B",X"20",X"F4",X"00",X"85",X"E6",X"81",X"4F",X"0F",X"1B",X"D1",X"A7",X"12",
		X"3D",X"20",X"ED",X"C3",X"D1",X"1B",X"24",X"24",X"3A",X"6F",X"20",X"F3",X"67",X"8C",X"F4",X"3A",
		X"DF",X"3A",X"F5",X"20",X"32",X"97",X"20",X"DF",X"D2",X"C3",X"CD",X"1F",X"17",X"88",X"20",X"26",
		X"1B",X"00",X"12",X"7C",X"7D",X"1B",X"3A",X"12",X"00",X"3A",X"6F",X"22",X"05",X"C3",X"00",X"1B",
		X"1D",X"A5",X"EE",X"3A",X"A7",X"20",X"C5",X"C2",X"20",X"DF",X"01",X"FE",X"EE",X"C3",X"CD",X"13",
		X"22",X"05",X"ED",X"3A",X"5F",X"20",X"19",X"16",X"3E",X"06",X"32",X"0C",X"20",X"EE",X"32",X"97",
		X"FE",X"22",X"D2",X"02",X"19",X"1B",X"54",X"C3",X"32",X"1A",X"22",X"02",X"1A",X"13",X"01",X"32",
		X"00",X"18",X"26",X"6F",X"7E",X"22",X"FE",X"2B",X"FE",X"19",X"CA",X"01",X"1B",X"68",X"49",X"C3",
		X"F9",X"CA",X"57",X"1F",X"77",X"97",X"4E",X"2B",X"CA",X"0C",X"1F",X"7A",X"2B",X"5E",X"A7",X"7E",
		X"A7",X"00",X"F8",X"C2",X"09",X"18",X"FE",X"7C",X"46",X"2B",X"95",X"C3",X"3A",X"06",X"20",X"DF",
		X"26",X"18",X"7E",X"27",X"C2",X"A7",X"02",X"06",X"DA",X"25",X"18",X"C3",X"3E",X"FE",X"BB",X"DA",
		X"01",X"3E",X"DF",X"32",X"3A",X"20",X"20",X"EF",X"98",X"C3",X"26",X"04",X"C3",X"3E",X"18",X"BB",
		X"01",X"3E",X"F4",X"32",X"3E",X"20",X"32",X"02",X"32",X"3C",X"20",X"EF",X"32",X"97",X"20",X"F3",
		X"18",X"ED",X"8A",X"CD",X"97",X"18",X"F6",X"32",X"20",X"F0",X"00",X"3A",X"FE",X"22",X"CA",X"05",
		X"2B",X"EB",X"C3",X"7D",X"1B",X"E0",X"00",X"00",X"32",X"20",X"20",X"DF",X"C2",X"C3",X"C9",X"04",
		X"00",X"01",X"FF",X"01",X"FF",X"00",X"FE",X"FF",X"FF",X"FF",X"FF",X"00",X"01",X"00",X"01",X"01",
		X"49",X"C3",X"79",X"18",X"04",X"32",X"78",X"22",X"C6",X"7D",X"6F",X"20",X"CE",X"7C",X"67",X"00",
		X"18",X"94",X"EB",X"22",X"C3",X"20",X"1B",X"C6",X"03",X"32",X"C3",X"22",X"19",X"5C",X"C3",X"2B",
		X"06",X"9D",X"10",X"D2",X"3A",X"1A",X"20",X"EB",X"32",X"97",X"20",X"DF",X"EC",X"3A",X"CD",X"20",
		X"03",X"FE",X"F0",X"DA",X"00",X"19",X"10",X"C3",X"A7",X"CD",X"D2",X"06",X"1A",X"10",X"1F",X"E6",
		X"32",X"7C",X"22",X"03",X"00",X"3A",X"CD",X"22",X"C3",X"1A",X"1D",X"E6",X"32",X"7D",X"22",X"04",
		X"23",X"23",X"F9",X"3A",X"BD",X"20",X"41",X"C3",X"18",X"8A",X"CA",X"C9",X"19",X"D0",X"23",X"23",
		X"7E",X"23",X"13",X"12",X"7E",X"23",X"13",X"12",X"00",X"02",X"16",X"5F",X"7E",X"21",X"13",X"12",
		X"19",X"9D",X"F9",X"3A",X"CD",X"20",X"19",X"72",X"C9",X"23",X"BC",X"CD",X"FE",X"00",X"DA",X"0D",
		X"20",X"F9",X"D9",X"C3",X"23",X"1E",X"77",X"97",X"77",X"78",X"12",X"3D",X"23",X"13",X"32",X"7B",
		X"CA",X"DA",X"3A",X"19",X"20",X"F8",X"72",X"CD",X"D6",X"C3",X"CD",X"1E",X"00",X"BC",X"07",X"FE",
		X"43",X"60",X"FF",X"FF",X"FF",X"FF",X"3C",X"77",X"78",X"19",X"0B",X"FE",X"BE",X"C2",X"C3",X"19",
		X"1F",X"17",X"97",X"23",X"C3",X"77",X"1F",X"14",X"13",X"12",X"7B",X"23",X"F8",X"32",X"C3",X"20",
		X"F7",X"3A",X"CD",X"20",X"19",X"72",X"77",X"78",X"BC",X"CD",X"FE",X"00",X"DA",X"0C",X"13",X"38",
		X"6A",X"C3",X"3E",X"19",X"C3",X"30",X"04",X"8F",X"12",X"3C",X"23",X"13",X"32",X"7B",X"20",X"F7",
		X"DB",X"32",X"32",X"20",X"20",X"DC",X"00",X"C9",X"57",X"97",X"EB",X"32",X"32",X"20",X"20",X"EC",
		X"20",X"FE",X"67",X"8C",X"25",X"FE",X"25",X"DA",X"1C",X"0A",X"FF",X"3A",X"85",X"20",X"3A",X"6F",
		X"26",X"1E",X"1B",X"25",X"12",X"7C",X"7D",X"1B",X"FE",X"1E",X"DA",X"3E",X"1E",X"1B",X"1B",X"CA",
		X"1E",X"1B",X"5F",X"1A",X"B3",X"0A",X"BC",X"C3",X"CD",X"12",X"1D",X"A5",X"26",X"C9",X"C3",X"3E",
		X"0F",X"07",X"00",X"FF",X"00",X"00",X"FF",X"07",X"80",X"1D",X"09",X"80",X"FF",X"0B",X"80",X"00",
		X"01",X"07",X"C0",X"FF",X"01",X"C0",X"FF",X"01",X"FE",X"FF",X"3F",X"F0",X"FF",X"07",X"C0",X"F0",
		X"80",X"80",X"80",X"FF",X"FF",X"00",X"21",X"FF",X"80",X"C0",X"00",X"01",X"80",X"FF",X"FF",X"80",
		X"C2",X"19",X"18",X"49",X"23",X"23",X"FE",X"7E",X"40",X"7F",X"11",X"3E",X"6F",X"85",X"FE",X"7E",
		X"FF",X"FF",X"00",X"00",X"02",X"05",X"80",X"FF",X"C2",X"08",X"06",X"A7",X"F8",X"C3",X"FF",X"1A",
		X"FF",X"FF",X"C0",X"00",X"07",X"01",X"00",X"FF",X"08",X"00",X"FF",X"05",X"80",X"00",X"08",X"00",
		X"FF",X"FF",X"80",X"40",X"00",X"01",X"20",X"FF",X"01",X"00",X"FF",X"01",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"EB",X"97",X"00",X"E9",X"02",X"3E",X"02",X"40",X"FF",X"01",X"20",X"00",X"02",X"00",
		X"21",X"20",X"E0",X"FF",X"FE",X"22",X"CD",X"20",X"FB",X"32",X"21",X"20",X"01",X"00",X"FC",X"22",
		X"00",X"1E",X"E5",X"2B",X"75",X"CD",X"E1",X"02",X"02",X"7F",X"23",X"00",X"A7",X"7E",X"D6",X"CA",
		X"3A",X"23",X"20",X"F7",X"C2",X"BD",X"1E",X"C2",X"A7",X"7A",X"82",X"CA",X"23",X"19",X"23",X"23",
		X"20",X"FE",X"87",X"CD",X"23",X"02",X"A7",X"7E",X"CD",X"00",X"1F",X"92",X"00",X"21",X"22",X"20",
		X"7A",X"E1",X"C3",X"A7",X"1F",X"10",X"00",X"00",X"14",X"CA",X"2B",X"1F",X"CD",X"E5",X"02",X"6B",
		X"FF",X"01",X"00",X"00",X"00",X"01",X"FF",X"FF",X"80",X"80",X"03",X"07",X"80",X"FF",X"03",X"00",
		X"20",X"FA",X"C3",X"BD",X"02",X"48",X"02",X"3E",X"A3",X"CA",X"23",X"19",X"23",X"23",X"3A",X"23",
		X"CD",X"20",X"05",X"A2",X"7E",X"23",X"CA",X"A7",X"FB",X"32",X"21",X"20",X"FF",X"FF",X"FC",X"22",
		X"A7",X"7A",X"3E",X"CA",X"23",X"13",X"23",X"23",X"1F",X"3E",X"E5",X"2B",X"61",X"CD",X"E1",X"02",
		X"92",X"CD",X"21",X"1F",X"E0",X"FF",X"FE",X"22",X"3A",X"23",X"20",X"F8",X"C2",X"BD",X"1F",X"2C",
		X"19",X"67",X"E5",X"2B",X"57",X"CD",X"E1",X"02",X"CD",X"20",X"05",X"AA",X"7E",X"23",X"CA",X"A7",
		X"1F",X"74",X"03",X"FE",X"E9",X"CA",X"3E",X"13",X"A7",X"7A",X"63",X"C3",X"00",X"19",X"CA",X"A7",
		X"1D",X"70",X"2B",X"5E",X"97",X"56",X"CA",X"BA",X"32",X"01",X"20",X"DF",X"13",X"03",X"C3",X"23",
		X"03",X"AA",X"2B",X"1C",X"2B",X"2B",X"C3",X"7D",X"1F",X"8B",X"77",X"12",X"8B",X"C3",X"1E",X"1F",
		X"3A",X"04",X"20",X"F6",X"06",X"C3",X"3A",X"04",X"1F",X"EA",X"F5",X"3A",X"A7",X"20",X"10",X"C2",
		X"CA",X"02",X"1F",X"B8",X"C8",X"21",X"C3",X"20",X"20",X"EF",X"01",X"FE",X"B2",X"CA",X"FE",X"1F",
		X"C4",X"21",X"5E",X"20",X"56",X"23",X"4E",X"23",X"1F",X"BB",X"C0",X"21",X"C3",X"20",X"1F",X"BB",
		X"E1",X"1D",X"C1",X"D1",X"E6",X"7D",X"CA",X"1F",X"46",X"23",X"C5",X"EB",X"E5",X"D5",X"53",X"CD",
		X"5F",X"8B",X"F3",X"3A",X"8A",X"20",X"1A",X"57",X"04",X"2A",X"54",X"D5",X"3A",X"5D",X"20",X"F4",
		X"18",X"10",X"00",X"32",X"C3",X"22",X"1B",X"DE",X"C2",X"A7",X"18",X"2D",X"F0",X"3A",X"C3",X"20",
		X"2B",X"1D",X"2B",X"2B",X"C3",X"7D",X"1B",X"DE",X"FE",X"79",X"DA",X"20",X"1D",X"A1",X"97",X"C3",
		X"C9",X"09",X"00",X"D3",X"02",X"D3",X"A6",X"C3",X"00",X"CD",X"CD",X"40",X"05",X"B2",X"CB",X"CD",
		X"FF",X"0F",X"0F",X"F0",X"FF",X"FF",X"FF",X"FF",X"F0",X"08",X"FF",X"0F",X"0F",X"F0",X"F0",X"FF",
		X"60",X"FF",X"FF",X"18",X"18",X"60",X"60",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"18",X"60",
		X"FF",X"FF",X"30",X"FF",X"FF",X"C0",X"C0",X"30",X"FF",X"18",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"30",X"FF",X"FF",X"C0",X"C0",X"30",X"FF",X"FF",
		X"FF",X"07",X"80",X"78",X"07",X"00",X"78",X"FF",X"80",X"78",X"07",X"00",X"78",X"FF",X"00",X"80",
		X"FF",X"0F",X"00",X"F0",X"0F",X"00",X"F0",X"FF",X"00",X"80",X"FF",X"07",X"F0",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"E0",X"1E",X"01",X"E0",X"FF",X"00",X"00",X"FF",X"0F",X"00",X"F0",X"0F",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"01",X"00",X"FF",X"1E",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3C",X"C0",X"FF",X"03",X"C0",X"00",X"03",X"3C",
		X"00",X"FF",X"78",X"80",X"FF",X"07",X"80",X"00",X"FF",X"FF",X"FF",X"FF",X"80",X"00",X"07",X"78",
		X"11",X"FF",X"FF",X"1F",X"1F",X"0E",X"00",X"FF",X"07",X"78",X"00",X"FF",X"78",X"80",X"FF",X"07",
		X"32",X"FF",X"FF",X"3A",X"3E",X"1C",X"00",X"FF",X"FF",X"0E",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"74",X"FF",X"FF",X"74",X"74",X"38",X"00",X"FF",X"FF",X"1C",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"02",X"FF",X"D1",X"B6",X"66",X"C3",X"00",X"1F",X"FF",X"38",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7C",X"23",X"40",X"FE",X"F6",X"C2",X"C9",X"1C",X"00",X"00",X"21",X"00",X"24",X"00",X"00",X"36",
		X"FF",X"00",X"00",X"80",X"FF",X"FF",X"FF",X"FF",X"C0",X"C0",X"01",X"03",X"C0",X"FF",X"01",X"80",
		X"FF",X"70",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"00",X"FF",X"E8",X"C8",X"70",X"00",X"FF",
		X"01",X"00",X"00",X"FF",X"FF",X"E0",X"FF",X"FF",X"F0",X"FF",X"01",X"F0",X"FF",X"01",X"10",X"E0",
		X"02",X"01",X"00",X"FF",X"00",X"C0",X"FF",X"01",X"E0",X"FF",X"03",X"E0",X"FF",X"02",X"60",X"C0",
		X"05",X"03",X"00",X"FF",X"00",X"80",X"FF",X"03",X"C0",X"FF",X"05",X"C0",X"FF",X"05",X"C0",X"80",
		X"D6",X"7D",X"4F",X"20",X"DE",X"7C",X"47",X"00",X"00",X"FF",X"0A",X"00",X"03",X"5F",X"57",X"0A",
		X"2F",X"1A",X"0A",X"5F",X"C3",X"A3",X"1C",X"E9",X"C5",X"E5",X"2F",X"1A",X"77",X"A6",X"D5",X"13",
		X"81",X"CD",X"FE",X"1D",X"C2",X"FF",X"1D",X"60",X"FE",X"1A",X"C2",X"FF",X"1D",X"63",X"E1",X"C1",
		X"67",X"00",X"D6",X"79",X"4F",X"20",X"DE",X"78",X"13",X"C9",X"C6",X"7D",X"6F",X"20",X"CE",X"7C",
		X"40",X"FE",X"9F",X"DA",X"26",X"1D",X"1A",X"25",X"47",X"00",X"25",X"FE",X"F0",X"DA",X"7C",X"1F",
		X"57",X"0A",X"D6",X"7D",X"4F",X"20",X"DE",X"7C",X"06",X"C9",X"1A",X"3E",X"0A",X"C9",X"03",X"5F",
		X"C3",X"D5",X"1E",X"2A",X"D1",X"02",X"13",X"03",X"47",X"00",X"C5",X"E5",X"B6",X"1A",X"13",X"77",
		X"CD",X"E1",X"1D",X"81",X"FF",X"FE",X"B2",X"C2",X"1A",X"23",X"FF",X"FE",X"B5",X"C2",X"C1",X"1D",
		X"EB",X"46",X"D5",X"C5",X"CD",X"E5",X"1D",X"53",X"C9",X"1D",X"23",X"5E",X"23",X"56",X"23",X"4E",
		X"1B",X"0F",X"4F",X"12",X"02",X"C2",X"3A",X"1E",X"D1",X"E1",X"C3",X"C1",X"19",X"30",X"E6",X"81",
		X"C3",X"67",X"1E",X"02",X"3A",X"C6",X"C3",X"6F",X"20",X"FD",X"6F",X"85",X"FC",X"3A",X"8C",X"20");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
