library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity cclimber_big_sprite_tile_bit1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of cclimber_big_sprite_tile_bit1 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"7F",
		X"00",X"01",X"03",X"06",X"0C",X"18",X"31",X"33",X"FF",X"FF",X"BF",X"3F",X"7F",X"FF",X"FF",X"FF",
		X"33",X"39",X"3D",X"3F",X"1F",X"1F",X"0F",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"1F",X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"F8",
		X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"1F",X"00",X"00",X"80",X"00",X"80",X"00",X"00",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"7C",X"76",X"7E",X"60",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"FE",X"F6",X"FE",X"C0",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"BF",X"7F",X"FF",X"FF",X"FF",X"FE",X"FC",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"1F",X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"F8",
		X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"1F",X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"E0",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"F8",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"C0",
		X"FE",X"F8",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"01",X"03",X"02",X"06",X"FC",X"F8",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"01",X"03",X"02",X"06",X"FC",X"F8",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7C",X"76",X"7E",X"60",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"7C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"76",X"7E",X"60",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"01",X"03",X"02",X"06",X"FC",X"F8",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"01",X"03",X"02",X"06",X"FC",X"F8",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"01",X"00",X"01",X"01",X"C0",X"C0",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"01",X"03",X"02",X"06",X"FC",X"F8",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"F0",X"18",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"F0",X"18",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"07",X"0F",X"1F",X"1F",X"07",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"3F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"3F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"1F",X"1F",X"0F",X"07",X"03",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"02",X"01",X"01",X"01",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"7F",X"FF",X"F9",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F9",X"FF",X"7F",X"3F",X"00",
		X"00",X"1F",X"3F",X"7C",X"78",X"78",X"78",X"78",X"00",X"E3",X"F3",X"FB",X"7B",X"7B",X"7B",X"7B",
		X"78",X"78",X"78",X"78",X"78",X"7C",X"3F",X"1F",X"03",X"7B",X"7B",X"7B",X"7B",X"FB",X"F3",X"E3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3C",X"3C",X"EA",X"D5",X"6B",X"75",X"7B",X"7D",X"F3",X"F3",X"AA",X"55",X"BA",X"F7",X"AF",X"F7",
		X"EF",X"F7",X"EB",X"F5",X"2A",X"15",X"F3",X"F3",X"BE",X"F7",X"BF",X"F7",X"AA",X"55",X"CF",X"CF",
		X"CF",X"CF",X"FF",X"F5",X"2A",X"35",X"EA",X"F5",X"3C",X"3C",X"FF",X"55",X"AA",X"55",X"AB",X"57",
		X"EA",X"F5",X"2A",X"35",X"EA",X"F5",X"EA",X"F5",X"AB",X"55",X"AA",X"55",X"AA",X"5F",X"BF",X"7D",
		X"2A",X"35",X"EA",X"F5",X"EA",X"FF",X"3C",X"3C",X"BA",X"7D",X"BF",X"5F",X"AA",X"FF",X"F3",X"F3",
		X"E0",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"C0",X"E0",X"F0",X"F8",X"F8",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"E0",X"E0",X"C0",X"C0",X"80",X"80",X"00",
		X"FE",X"FC",X"FC",X"F8",X"F8",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C7",X"E7",X"F7",X"F7",X"F7",X"F7",X"F7",X"07",X"FC",X"FE",X"9F",X"8F",X"8F",X"8F",X"9F",X"FE",
		X"F7",X"F7",X"F7",X"F7",X"F7",X"E7",X"C7",X"00",X"FC",X"BC",X"BE",X"9E",X"9F",X"8F",X"8F",X"00",
		X"00",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"00",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"FE",X"FE",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CF",X"CF",X"AA",X"55",X"AE",X"DD",X"EE",X"7D",X"3C",X"3C",X"AA",X"55",X"BB",X"5F",X"AB",X"DF",
		X"AF",X"7D",X"EE",X"DD",X"AA",X"55",X"3C",X"3C",X"FB",X"DF",X"FB",X"DF",X"AA",X"55",X"F3",X"F3",
		X"F3",X"F3",X"FF",X"55",X"FB",X"DF",X"AB",X"D7",X"CF",X"CF",X"FF",X"55",X"EA",X"75",X"BB",X"77",
		X"AB",X"DF",X"FB",X"55",X"AA",X"75",X"BB",X"F5",X"EB",X"77",X"BB",X"55",X"AA",X"F5",X"BB",X"FF",
		X"BB",X"F5",X"BB",X"7D",X"AA",X"FF",X"CF",X"CF",X"BF",X"F5",X"BB",X"F5",X"AA",X"FF",X"3C",X"3C",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"F7",X"F7",X"F7",X"F1",X"FF",X"FF",X"FF",X"FF",X"B4",X"5D",X"36",X"94",
		X"FF",X"FF",X"FF",X"FF",X"A9",X"AB",X"AD",X"89",X"FF",X"FF",X"FF",X"FF",X"BD",X"5B",X"1B",X"5D",
		X"FF",X"FF",X"FF",X"FF",X"57",X"55",X"53",X"15",X"FF",X"FF",X"FF",X"FF",X"DA",X"DA",X"DA",X"4A",
		X"07",X"07",X"07",X"8E",X"8E",X"8E",X"DC",X"DC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DC",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"07",X"07",X"0F",X"0F",X"0F",X"1F",X"1E",X"F0",X"F0",X"F0",X"F8",X"78",X"78",X"7C",X"3C",
		X"1E",X"3E",X"3F",X"3F",X"7C",X"78",X"F8",X"00",X"3C",X"3E",X"FE",X"FE",X"1F",X"0F",X"0F",X"00",
		X"00",X"E0",X"E0",X"E0",X"F1",X"F1",X"F1",X"FB",X"00",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",
		X"FB",X"FB",X"BF",X"BF",X"BF",X"9F",X"9F",X"9F",X"FD",X"FD",X"BD",X"BD",X"BD",X"3D",X"3D",X"3D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3C",X"3C",X"AA",X"55",X"AA",X"55",X"AE",X"77",X"F3",X"F3",X"AA",X"55",X"AA",X"57",X"EF",X"7F",
		X"FE",X"57",X"FF",X"77",X"AA",X"55",X"CF",X"CF",X"EE",X"77",X"EF",X"F7",X"AA",X"55",X"3C",X"3C",
		X"F3",X"F3",X"FF",X"55",X"EB",X"F5",X"BA",X"5D",X"CF",X"CF",X"FF",X"55",X"FE",X"77",X"EA",X"D7",
		X"FB",X"5F",X"BB",X"55",X"AA",X"FF",X"BB",X"F7",X"AB",X"55",X"FB",X"55",X"AA",X"7D",X"EB",X"75",
		X"BE",X"F7",X"BB",X"FF",X"AA",X"FF",X"3C",X"3C",X"FF",X"75",X"EB",X"7D",X"AA",X"FF",X"F3",X"F3",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FA",X"A9",X"AB",X"8B",X"FF",X"FF",X"FF",X"FF",X"DF",X"AF",X"9F",X"CF",
		X"FF",X"FF",X"FF",X"FF",X"BD",X"5D",X"5D",X"B4",X"FF",X"FF",X"FF",X"FF",X"13",X"B5",X"B5",X"B3",
		X"FF",X"FF",X"FF",X"FF",X"A8",X"2D",X"2D",X"AD",X"FF",X"FF",X"FF",X"FF",X"89",X"9A",X"9A",X"89",
		X"00",X"EF",X"EF",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"F8",X"FC",X"3E",X"1E",X"1E",X"1E",X"3E",
		X"EF",X"0F",X"0F",X"0F",X"0F",X"0F",X"EF",X"EF",X"FC",X"F8",X"78",X"7C",X"3C",X"3E",X"1E",X"1E",
		X"7F",X"7F",X"7F",X"07",X"07",X"0F",X"0F",X"1F",X"FF",X"EF",X"EF",X"EF",X"C7",X"C7",X"87",X"83",
		X"1F",X"3F",X"3E",X"7E",X"7F",X"7F",X"FF",X"00",X"03",X"03",X"01",X"00",X"E0",X"E0",X"E0",X"00",
		X"00",X"FF",X"FF",X"E7",X"E3",X"E3",X"E3",X"E7",X"00",X"1F",X"9F",X"DE",X"DE",X"DE",X"DE",X"9E",
		X"FF",X"E7",X"E3",X"E3",X"E3",X"E7",X"FF",X"FF",X"1F",X"9E",X"DE",X"DE",X"DE",X"DE",X"9F",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CF",X"CF",X"AA",X"55",X"AA",X"5F",X"BB",X"F5",X"3C",X"3C",X"AB",X"57",X"A8",X"54",X"EE",X"76",
		X"BE",X"D7",X"BB",X"5F",X"AA",X"55",X"F3",X"F3",X"EF",X"77",X"FF",X"7F",X"A8",X"54",X"CF",X"CF",
		X"3C",X"3C",X"FF",X"55",X"EA",X"75",X"EA",X"D5",X"F3",X"F3",X"FF",X"57",X"AC",X"54",X"AF",X"57",
		X"AA",X"D5",X"AA",X"55",X"AA",X"F5",X"BA",X"DD",X"AF",X"57",X"AC",X"54",X"AF",X"57",X"AF",X"57",
		X"BA",X"F5",X"BA",X"DD",X"AA",X"FF",X"CF",X"CF",X"AC",X"54",X"AF",X"57",X"AF",X"FF",X"3C",X"3C");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
