library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity tropical_chr_bit1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of tropical_chr_bit1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FD",X"F9",X"FB",X"FB",X"FB",X"FB",X"F3",X"F7",
		X"00",X"00",X"00",X"C0",X"80",X"C0",X"C0",X"60",X"7F",X"3F",X"3F",X"3C",X"74",X"20",X"60",X"20",
		X"FF",X"FF",X"FF",X"BF",X"1F",X"1F",X"3F",X"BF",X"FF",X"FE",X"FC",X"FE",X"FC",X"FB",X"FF",X"FE",
		X"40",X"00",X"1C",X"7D",X"E0",X"80",X"0A",X"BF",X"20",X"00",X"3D",X"3D",X"1E",X"3E",X"7C",X"E0",
		X"21",X"53",X"DF",X"FF",X"FF",X"7F",X"3F",X"1F",X"FF",X"FF",X"FF",X"FF",X"FC",X"FE",X"FC",X"FC",
		X"F8",X"FC",X"99",X"30",X"38",X"73",X"77",X"E7",X"1F",X"3F",X"1F",X"5F",X"DF",X"DF",X"9F",X"BF",
		X"FC",X"F9",X"F3",X"FB",X"F7",X"F7",X"EF",X"FF",X"00",X"01",X"03",X"04",X"14",X"30",X"20",X"20",
		X"FE",X"FF",X"FF",X"FB",X"FC",X"FE",X"FC",X"F8",X"9B",X"11",X"81",X"C3",X"C3",X"01",X"01",X"01",
		X"FF",X"FF",X"EF",X"CF",X"DF",X"BF",X"3F",X"3F",X"FF",X"FC",X"FF",X"FF",X"8F",X"43",X"F4",X"A8",
		X"38",X"E0",X"C0",X"80",X"80",X"90",X"D0",X"C8",X"00",X"00",X"00",X"01",X"01",X"07",X"07",X"0F",
		X"50",X"60",X"60",X"E0",X"E0",X"E0",X"F0",X"F8",X"0F",X"0F",X"17",X"17",X"1B",X"1B",X"01",X"03",
		X"F8",X"F8",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"0F",X"0F",X"1F",X"0F",X"1C",X"00",X"00",X"00",
		X"E0",X"D8",X"BC",X"7C",X"7C",X"FC",X"FC",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"FC",X"7C",X"1E",X"0E",X"0E",X"06",X"06",X"46",X"D1",X"F1",X"B0",X"10",X"00",X"02",X"03",X"03",
		X"C7",X"E2",X"82",X"82",X"80",X"84",X"86",X"06",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"00",X"00",X"10",X"00",
		X"28",X"28",X"28",X"00",X"00",X"00",X"00",X"00",X"28",X"28",X"7C",X"28",X"7C",X"28",X"28",X"00",
		X"10",X"3C",X"50",X"38",X"14",X"78",X"10",X"00",X"60",X"64",X"08",X"10",X"20",X"4C",X"0C",X"00",
		X"30",X"48",X"50",X"20",X"54",X"48",X"34",X"00",X"30",X"10",X"20",X"00",X"00",X"00",X"00",X"00",
		X"08",X"10",X"20",X"20",X"20",X"10",X"08",X"00",X"20",X"10",X"08",X"08",X"08",X"10",X"20",X"00",
		X"00",X"10",X"54",X"38",X"54",X"10",X"00",X"00",X"00",X"10",X"10",X"7C",X"10",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"30",X"10",X"20",X"00",X"00",X"00",X"00",X"7C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"30",X"30",X"00",X"00",X"04",X"08",X"10",X"20",X"40",X"00",X"00",
		X"38",X"4C",X"C6",X"C6",X"C6",X"64",X"38",X"00",X"30",X"70",X"30",X"30",X"30",X"30",X"FC",X"00",
		X"7C",X"C6",X"0E",X"3C",X"78",X"E0",X"FE",X"00",X"7E",X"0C",X"18",X"3C",X"06",X"C6",X"7C",X"00",
		X"1C",X"3C",X"6C",X"CC",X"FE",X"0C",X"0C",X"00",X"F8",X"C0",X"F8",X"0C",X"0C",X"CC",X"78",X"00",
		X"3C",X"60",X"C0",X"FC",X"C6",X"C6",X"7C",X"00",X"FE",X"C6",X"0C",X"18",X"30",X"30",X"30",X"00",
		X"78",X"C4",X"E4",X"78",X"9E",X"86",X"7C",X"00",X"7C",X"C6",X"C6",X"7E",X"06",X"0C",X"78",X"00",
		X"00",X"30",X"30",X"00",X"30",X"30",X"00",X"00",X"00",X"30",X"30",X"00",X"30",X"10",X"20",X"00",
		X"04",X"08",X"10",X"20",X"10",X"08",X"04",X"00",X"00",X"00",X"7E",X"00",X"7E",X"00",X"00",X"00",
		X"20",X"10",X"08",X"04",X"08",X"10",X"20",X"00",X"38",X"44",X"04",X"08",X"10",X"00",X"10",X"00",
		X"3C",X"42",X"99",X"A1",X"A1",X"99",X"42",X"3C",X"38",X"6C",X"C6",X"C6",X"FE",X"C6",X"C6",X"00",
		X"FC",X"C6",X"C6",X"FC",X"C6",X"C6",X"FC",X"00",X"3C",X"66",X"C0",X"C0",X"C0",X"66",X"3C",X"00",
		X"F8",X"CC",X"C6",X"C6",X"C6",X"CC",X"F8",X"00",X"FC",X"C0",X"C0",X"F8",X"C0",X"C0",X"FE",X"00",
		X"FE",X"C0",X"C0",X"FC",X"C0",X"C0",X"C0",X"00",X"3E",X"60",X"C0",X"CE",X"C6",X"66",X"3E",X"00",
		X"C6",X"C6",X"C6",X"FE",X"C6",X"C6",X"C6",X"00",X"FC",X"30",X"30",X"30",X"30",X"30",X"FC",X"00",
		X"06",X"06",X"06",X"06",X"06",X"C6",X"78",X"00",X"C6",X"CC",X"D8",X"F0",X"F8",X"DC",X"CE",X"00",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"FE",X"00",X"C6",X"EE",X"FE",X"FE",X"D6",X"C6",X"C6",X"00",
		X"C6",X"E6",X"F6",X"FE",X"DE",X"CE",X"C6",X"00",X"7C",X"C6",X"C6",X"C6",X"C6",X"C6",X"7C",X"00",
		X"FC",X"C6",X"C6",X"C6",X"FC",X"C0",X"C0",X"00",X"7C",X"C6",X"C6",X"C6",X"DE",X"CC",X"7A",X"00",
		X"FC",X"C6",X"C6",X"CE",X"F8",X"DC",X"CE",X"00",X"78",X"CC",X"C0",X"7C",X"06",X"C6",X"7C",X"00",
		X"FC",X"30",X"30",X"30",X"30",X"30",X"30",X"00",X"C6",X"C6",X"C6",X"C6",X"C6",X"C6",X"7C",X"00",
		X"C6",X"C6",X"C6",X"EE",X"7C",X"38",X"10",X"00",X"C6",X"C6",X"D6",X"FE",X"FE",X"EE",X"C6",X"00",
		X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",X"CC",X"CC",X"CC",X"78",X"30",X"30",X"30",X"00",
		X"FC",X"FC",X"18",X"30",X"60",X"FC",X"FC",X"00",X"38",X"20",X"20",X"20",X"20",X"20",X"38",X"00",
		X"80",X"40",X"20",X"10",X"08",X"04",X"02",X"00",X"38",X"08",X"08",X"08",X"08",X"08",X"38",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"FF",X"FF",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"0E",X"0C",X"0C",X"0C",X"0C",X"08",X"18",X"18",X"FF",X"FF",X"7F",X"1D",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"F8",X"C0",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"7F",X"01",X"00",X"00",X"0C",X"18",X"31",X"FC",X"FE",
		X"10",X"B0",X"B0",X"90",X"90",X"C8",X"44",X"F8",X"F9",X"FF",X"FF",X"F8",X"EC",X"C0",X"00",X"00",
		X"E6",X"FF",X"FC",X"CF",X"E3",X"C0",X"00",X"58",X"70",X"F8",X"E0",X"80",X"E0",X"00",X"04",X"B2",
		X"F9",X"FF",X"FF",X"F8",X"EC",X"C0",X"00",X"00",X"3F",X"00",X"00",X"00",X"00",X"40",X"EE",X"FF",
		X"FF",X"00",X"00",X"00",X"68",X"3D",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"40",X"F6",X"AF",X"FF",
		X"FF",X"03",X"00",X"01",X"0B",X"BF",X"EF",X"FF",X"FE",X"FF",X"FF",X"5E",X"EB",X"44",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"81",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"81",
		X"81",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"81",
		X"00",X"00",X"00",X"00",X"03",X"01",X"03",X"07",X"03",X"01",X"08",X"19",X"3D",X"78",X"3B",X"3F",
		X"00",X"06",X"8F",X"9F",X"BF",X"7F",X"FF",X"FE",X"EE",X"E5",X"F8",X"71",X"FB",X"FD",X"EE",X"CE",
		X"00",X"00",X"00",X"0A",X"9E",X"9D",X"3F",X"5F",X"BF",X"FD",X"FB",X"F4",X"E6",X"DF",X"FF",X"7E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"B0",X"B0",X"A0",X"40",X"00",X"0C",X"18",X"00",X"00",
		X"00",X"02",X"06",X"0F",X"0F",X"1F",X"0E",X"2F",X"77",X"7E",X"7D",X"75",X"2A",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"40",X"80",X"00",X"20",X"60",X"48",X"00",X"A0",X"40",X"80",X"00",
		X"1E",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"BC",X"8C",X"51",X"B3",X"62",X"60",X"F0",X"00",
		X"BC",X"78",X"ED",X"92",X"03",X"00",X"00",X"00",X"16",X"2D",X"5D",X"1A",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"98",X"30",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"02",X"04",X"00",X"04",X"08",X"18",X"00",X"00",
		X"02",X"0F",X"1F",X"3F",X"2D",X"5E",X"79",X"30",X"07",X"23",X"72",X"D1",X"EA",X"EA",X"D4",X"76",
		X"00",X"00",X"D0",X"B8",X"F8",X"F0",X"E0",X"80",X"BF",X"FD",X"FB",X"F4",X"E6",X"DF",X"FF",X"7F",
		X"21",X"73",X"FB",X"E9",X"F3",X"FB",X"77",X"3F",X"7E",X"FF",X"77",X"6B",X"31",X"00",X"00",X"00",
		X"FF",X"FE",X"BF",X"D7",X"CF",X"BF",X"BF",X"5F",X"4F",X"EF",X"F2",X"61",X"83",X"04",X"01",X"00",
		X"00",X"00",X"00",X"01",X"03",X"01",X"23",X"67",X"77",X"3F",X"7F",X"FF",X"7F",X"BF",X"BF",X"7E",
		X"00",X"00",X"20",X"70",X"E0",X"C0",X"80",X"C0",X"E0",X"F0",X"F0",X"F8",X"E0",X"40",X"81",X"83",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"8E",X"1C",X"18",X"38",X"28",X"50",X"00",X"02",X"1C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"B0",X"A0",X"40",X"08",X"1E",X"3D",X"DE",X"EF",X"DF",X"8E",X"57",X"FE",X"F8",X"FE",X"FF",X"FF",
		X"1E",X"00",X"01",X"00",X"00",X"00",X"C3",X"F1",X"E8",X"94",X"00",X"80",X"14",X"FE",X"DF",X"00",
		X"BC",X"78",X"ED",X"92",X"07",X"C3",X"B1",X"E2",X"44",X"1E",X"0D",X"00",X"44",X"EE",X"93",X"04",
		X"BC",X"8C",X"5D",X"F9",X"F3",X"E2",X"07",X"88",X"00",X"00",X"02",X"80",X"44",X"EE",X"FF",X"0F",
		X"16",X"2D",X"5D",X"9A",X"D0",X"80",X"00",X"04",X"1D",X"23",X"76",X"FC",X"26",X"FF",X"FF",X"F0",
		X"00",X"00",X"00",X"08",X"1E",X"3D",X"DE",X"EF",X"1D",X"23",X"76",X"FC",X"26",X"FF",X"FF",X"F0",
		X"00",X"00",X"00",X"40",X"E8",X"FD",X"9E",X"00",X"BC",X"78",X"ED",X"92",X"8F",X"FF",X"E3",X"00",
		X"00",X"00",X"00",X"00",X"E0",X"F0",X"78",X"00",X"BF",X"8E",X"5F",X"FD",X"FF",X"FF",X"FB",X"07",
		X"00",X"00",X"00",X"00",X"04",X"09",X"1C",X"00",X"00",X"00",X"00",X"00",X"82",X"1D",X"73",X"00",
		X"00",X"00",X"00",X"00",X"82",X"1D",X"63",X"08",X"00",X"00",X"00",X"00",X"41",X"B8",X"CE",X"00",
		X"00",X"00",X"00",X"00",X"20",X"90",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C3",X"F1",
		X"1E",X"00",X"01",X"00",X"07",X"0F",X"1F",X"00",X"00",X"00",X"00",X"00",X"01",X"C3",X"B1",X"E2",
		X"00",X"00",X"1C",X"79",X"F3",X"E2",X"07",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"C3",X"F1",
		X"00",X"00",X"00",X"80",X"C0",X"80",X"00",X"04",X"00",X"00",X"00",X"00",X"01",X"C3",X"B1",X"E2",
		X"A0",X"CC",X"1A",X"BD",X"7A",X"BE",X"6D",X"DF",X"00",X"8C",X"5C",X"BC",X"EE",X"77",X"AC",X"F9",
		X"3C",X"38",X"25",X"C4",X"ED",X"EF",X"DB",X"EE",X"00",X"00",X"20",X"74",X"99",X"5B",X"FD",X"EF",
		X"00",X"00",X"00",X"80",X"00",X"80",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"A0",X"B0",X"E8",X"78",X"E8",X"DF",X"60",X"00",X"05",X"0D",X"17",X"1E",X"17",X"FB",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"5C",X"EC",X"7F",X"FA",X"67",X"F7",X"9D",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"87",X"CC",X"BE",X"F7",X"FF",X"7A",X"30",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"11",X"7A",X"F3",X"EF",X"FF",X"FF",X"6E",X"38",X"30",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"83",X"87",X"C7",X"6F",X"CD",X"EB",X"FF",X"13",X"00",
		X"00",X"00",X"00",X"01",X"00",X"00",X"01",X"80",X"D4",X"EA",X"F0",X"D8",X"B2",X"FD",X"03",X"00",
		X"00",X"00",X"40",X"30",X"80",X"C0",X"80",X"80",X"00",X"00",X"40",X"2E",X"F3",X"7C",X"E9",X"00",
		X"C0",X"80",X"0A",X"04",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"90",X"62",X"0D",X"03",X"00",
		X"01",X"03",X"01",X"11",X"0C",X"08",X"00",X"00",X"01",X"09",X"9B",X"4F",X"7F",X"BB",X"F7",X"E7",
		X"FD",X"FE",X"BF",X"D7",X"0F",X"00",X"00",X"00",X"82",X"C5",X"1F",X"AF",X"F7",X"E7",X"BD",X"7E",
		X"07",X"23",X"72",X"D1",X"EA",X"6A",X"04",X"16",X"38",X"74",X"BE",X"FD",X"F6",X"D9",X"BD",X"0F",
		X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"01",X"03",X"07",X"E3",X"F7",X"CE",X"7C",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"08",X"00",
		X"3C",X"38",X"C5",X"61",X"F8",X"F4",X"FA",X"E0",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",
		X"00",X"8C",X"9C",X"80",X"00",X"00",X"20",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"87",X"CF",X"FD",X"6E",X"BF",X"77",X"21",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F7",X"F7",X"E7",X"EF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"D9",X"64",X"C0",X"40",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"DE",X"F6",X"BD",X"F6",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"ED",X"BF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"6F",X"18",X"00",X"00",X"00",X"00",X"00",X"FE",X"EE",X"BB",X"E6",X"38",X"10",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"51",X"A4",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"53",X"FF",
		X"FF",X"F7",X"BF",X"ED",X"52",X"14",X"00",X"00",X"FF",X"FB",X"AE",X"5B",X"17",X"06",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"BC",X"EF",X"FB",X"6C",X"DF",X"CA",X"90",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"7B",X"2E",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"FD",X"B3",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"B4",X"FF",X"E7",X"EF",X"DE",X"DE",X"DE",X"9D",X"BF",X"BF",
		X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"BF",X"BF",X"BF",X"3F",X"7F",X"7F",X"7F",
		X"FF",X"FE",X"FE",X"FE",X"FE",X"FC",X"FD",X"FD",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"70",X"7C",X"7E",X"7C",X"70",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"0C",X"1E",X"37",X"FC",X"7F",X"1F",X"09",X"04",X"00",X"18",X"63",X"04",X"00",
		X"1E",X"7B",X"FC",X"AE",X"10",X"00",X"00",X"41",X"8C",X"18",X"A0",X"78",X"F1",X"EE",X"FC",X"68",
		X"CC",X"86",X"D1",X"08",X"5C",X"3F",X"37",X"4F",X"FC",X"36",X"0D",X"1C",X"36",X"71",X"F8",X"44",
		X"01",X"08",X"1F",X"2C",X"01",X"03",X"C5",X"9F",X"8F",X"DD",X"1B",X"3F",X"66",X"0C",X"0F",X"1C",
		X"EE",X"7D",X"38",X"08",X"E4",X"D0",X"00",X"88",X"F0",X"C0",X"00",X"80",X"43",X"00",X"00",X"80",
		X"60",X"48",X"07",X"01",X"03",X"01",X"03",X"04",X"18",X"30",X"60",X"E0",X"04",X"03",X"00",X"00",
		X"00",X"09",X"03",X"80",X"C1",X"87",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"04",X"03",X"07",
		X"E0",X"C0",X"E0",X"C0",X"8F",X"03",X"01",X"03",X"07",X"03",X"1E",X"F8",X"44",X"80",X"E0",X"00",
		X"01",X"03",X"05",X"8F",X"1E",X"FF",X"F9",X"BF",X"F3",X"00",X"A0",X"18",X"7C",X"3F",X"3F",X"7B",
		X"C6",X"80",X"00",X"08",X"F0",X"CA",X"EC",X"C8",X"01",X"F6",X"7C",X"08",X"FC",X"F8",X"9C",X"2E",
		X"0C",X"0B",X"1E",X"34",X"40",X"04",X"28",X"79",X"37",X"16",X"3F",X"69",X"3E",X"1C",X"0F",X"07",
		X"17",X"01",X"67",X"09",X"93",X"78",X"25",X"83",X"E6",X"37",X"8C",X"9B",X"41",X"03",X"E1",X"80",
		X"80",X"C4",X"B9",X"F0",X"A0",X"08",X"32",X"FC",X"9A",X"E0",X"F1",X"CC",X"9B",X"FE",X"E4",X"6F",
		X"E1",X"B1",X"8A",X"46",X"1E",X"3F",X"99",X"7F",X"36",X"FD",X"7F",X"33",X"47",X"0E",X"FC",X"FF",
		X"E0",X"91",X"C4",X"20",X"00",X"80",X"C0",X"20",X"00",X"00",X"C0",X"80",X"40",X"00",X"00",X"10",
		X"60",X"B9",X"1E",X"20",X"01",X"00",X"00",X"00",X"18",X"34",X"78",X"D0",X"00",X"00",X"00",X"00",
		X"04",X"03",X"02",X"0F",X"9C",X"78",X"32",X"1C",X"0F",X"08",X"50",X"3E",X"0D",X"1F",X"23",X"06",
		X"E0",X"93",X"47",X"03",X"47",X"3F",X"18",X"10",X"20",X"80",X"09",X"07",X"03",X"8F",X"FD",X"70",
		X"3F",X"02",X"DE",X"F7",X"67",X"FF",X"FC",X"38",X"0E",X"40",X"80",X"00",X"C8",X"F0",X"BB",X"FF",
		X"00",X"00",X"00",X"00",X"20",X"C8",X"F0",X"00",X"80",X"60",X"30",X"A0",X"70",X"C0",X"C0",X"80",
		X"C2",X"88",X"7E",X"F3",X"F9",X"E4",X"F0",X"3E",X"FE",X"ED",X"B0",X"45",X"13",X"04",X"23",X"61",
		X"F1",X"7E",X"FA",X"9C",X"FA",X"35",X"7F",X"3F",X"CF",X"73",X"A7",X"88",X"F5",X"E3",X"BB",X"C6",
		X"1F",X"1B",X"3F",X"3E",X"1D",X"07",X"BF",X"FE",X"3F",X"DE",X"84",X"F2",X"E8",X"C4",X"F8",X"C0",
		X"00",X"80",X"40",X"00",X"01",X"80",X"00",X"00",X"60",X"08",X"07",X"03",X"01",X"06",X"08",X"30",
		X"01",X"00",X"20",X"C2",X"E1",X"00",X"00",X"01",X"03",X"26",X"0F",X"86",X"18",X"00",X"00",X"00",
		X"E2",X"C4",X"70",X"C0",X"E0",X"7F",X"FF",X"A6",X"00",X"00",X"88",X"F1",X"3F",X"1F",X"7B",X"3E",
		X"3F",X"0F",X"19",X"30",X"E0",X"FC",X"BF",X"1F",X"38",X"60",X"E2",X"FC",X"F2",X"3B",X"F0",X"60",
		X"E4",X"F8",X"E0",X"38",X"58",X"30",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"1F",X"3E",X"17",X"79",X"F3",X"A9",X"67",
		X"64",X"FF",X"5F",X"F9",X"3C",X"0F",X"3F",X"FE",X"ED",X"13",X"01",X"93",X"E1",X"FB",X"FC",X"68",
		X"FC",X"7A",X"FE",X"D8",X"F6",X"3F",X"FF",X"EF",X"C7",X"F1",X"E3",X"B7",X"CF",X"F3",X"7E",X"2C",
		X"D8",X"7C",X"3C",X"76",X"3C",X"FE",X"7C",X"B8",X"24",X"F0",X"F0",X"C9",X"E3",X"BD",X"C0",X"00",
		X"00",X"00",X"03",X"06",X"00",X"00",X"80",X"38",X"1C",X"39",X"60",X"C0",X"80",X"D0",X"EC",X"03",
		X"3C",X"1E",X"0C",X"1F",X"1F",X"3E",X"78",X"FC",X"7E",X"8F",X"07",X"4F",X"3E",X"78",X"F1",X"C3",
		X"7F",X"9F",X"0E",X"1C",X"FF",X"EF",X"1E",X"3C",X"7F",X"FC",X"FE",X"DC",X"07",X"61",X"FF",X"E9",
		X"F0",X"F8",X"70",X"18",X"B8",X"E0",X"00",X"80",X"00",X"C0",X"00",X"40",X"80",X"80",X"C0",X"E0",
		X"03",X"0F",X"3F",X"67",X"CB",X"FF",X"FF",X"73",X"3B",X"1D",X"7F",X"F7",X"CE",X"87",X"DB",X"FF",
		X"FF",X"DE",X"FF",X"7C",X"FF",X"EE",X"77",X"C3",X"F1",X"FF",X"FF",X"99",X"CF",X"1F",X"EF",X"FE",
		X"FC",X"E8",X"7C",X"F9",X"F0",X"C0",X"E0",X"C0",X"F0",X"E0",X"C3",X"01",X"87",X"3F",X"ED",X"07",
		X"19",X"3C",X"F0",X"79",X"03",X"03",X"21",X"C3",X"07",X"03",X"8F",X"C7",X"80",X"81",X"27",X"DF",
		X"F1",X"7F",X"FC",X"E7",X"DF",X"9F",X"C7",X"EF",X"FF",X"F1",X"C3",X"EF",X"FF",X"FF",X"C3",X"1C",
		X"FE",X"F8",X"F8",X"3C",X"FC",X"FC",X"98",X"0C",X"FC",X"F0",X"C0",X"80",X"C0",X"80",X"C0",X"E0",
		X"06",X"03",X"3F",X"FF",X"66",X"FF",X"AF",X"F9",X"FF",X"FD",X"FC",X"CC",X"F8",X"7C",X"10",X"F8",
		X"B8",X"FC",X"E8",X"E0",X"C0",X"E0",X"00",X"80",X"C0",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"02",X"01",X"00",X"05",X"03",X"07",X"0E",X"DD",X"8F",X"1F",X"3B",X"17",X"32",X"7F",X"7C",
		X"FF",X"D7",X"BD",X"BD",X"FB",X"FF",X"FF",X"DF",X"FD",X"7F",X"FF",X"FF",X"E7",X"F3",X"FF",X"FF",
		X"00",X"01",X"0F",X"1F",X"0F",X"3E",X"FC",X"F8",X"D0",X"E1",X"A0",X"81",X"03",X"82",X"01",X"03",
		X"3F",X"FE",X"F0",X"C0",X"00",X"00",X"07",X"1F",X"77",X"FF",X"FD",X"BF",X"FF",X"EF",X"FF",X"7F",
		X"00",X"02",X"0C",X"1B",X"1E",X"BC",X"64",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",
		X"01",X"03",X"03",X"01",X"03",X"01",X"00",X"00",X"00",X"03",X"0F",X"3C",X"6E",X"F8",X"FC",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"01",X"07",X"07",X"03",X"00",
		X"00",X"00",X"00",X"00",X"03",X"07",X"03",X"00",X"03",X"1F",X"79",X"B7",X"FF",X"FA",X"9F",X"DF",
		X"00",X"00",X"00",X"03",X"0F",X"1F",X"3A",X"71",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"07",X"1D",X"3F",X"1F",X"FF",X"94",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"01",X"07",X"03",X"00",X"10",X"60",
		X"01",X"00",X"00",X"00",X"00",X"00",X"03",X"0F",X"65",X"F0",X"B8",X"E0",X"FA",X"FC",X"48",X"24",
		X"F9",X"F0",X"DF",X"7E",X"3C",X"F6",X"DC",X"E6",X"70",X"81",X"00",X"00",X"05",X"33",X"61",X"80",
		X"06",X"0F",X"87",X"07",X"01",X"30",X"18",X"44",X"20",X"70",X"FC",X"FF",X"3E",X"F2",X"BB",X"74",
		X"6D",X"F8",X"F3",X"9F",X"BF",X"07",X"21",X"7C",X"B0",X"07",X"0F",X"14",X"7E",X"37",X"6F",X"7C",
		X"1D",X"1C",X"B8",X"F0",X"FC",X"B9",X"F5",X"E0",X"20",X"90",X"40",X"00",X"20",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"80",X"20",X"1C",X"02",X"07",X"03",X"06",X"08",X"30",X"60",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"01",X"13",X"07",X"01",X"83",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"1A",X"1F",X"3F",X"47",X"0C",X"C0",X"80",X"C0",X"81",X"1E",X"07",X"03",X"07",X"0F",X"06",X"3D",
		X"07",X"1F",X"FE",X"FB",X"E1",X"03",X"07",X"0B",X"1F",X"3E",X"FF",X"F9",X"7F",X"E6",X"01",X"00",
		X"C0",X"90",X"E1",X"F7",X"FF",X"8C",X"00",X"00",X"00",X"F0",X"8A",X"CC",X"88",X"02",X"EC",X"F8",
		X"70",X"E0",X"C0",X"C0",X"80",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"07",X"3F",X"7F",
		X"01",X"07",X"03",X"10",X"60",X"58",X"F1",X"A0",X"02",X"21",X"40",X"CC",X"BF",X"B8",X"FE",X"A6",
		X"B8",X"E0",X"F0",X"FD",X"5E",X"07",X"9E",X"27",X"4E",X"E0",X"94",X"0F",X"1A",X"9F",X"33",X"6F",
		X"4F",X"13",X"8E",X"87",X"03",X"12",X"E6",X"C1",X"80",X"20",X"CA",X"F1",X"68",X"83",X"C5",X"30",
		X"D7",X"8F",X"EF",X"1B",X"87",X"C7",X"29",X"1C",X"7C",X"FF",X"73",X"FE",X"D8",X"F4",X"FF",X"CE",
		X"A0",X"10",X"E0",X"80",X"C0",X"23",X"88",X"40",X"00",X"00",X"80",X"40",X"00",X"00",X"00",X"00",
		X"02",X"0C",X"10",X"60",X"C0",X"72",X"2C",X"40",X"03",X"00",X"00",X"00",X"30",X"68",X"D0",X"A0",
		X"30",X"00",X"00",X"00",X"09",X"07",X"04",X"1E",X"38",X"F0",X"64",X"38",X"1E",X"11",X"A0",X"7C",
		X"7F",X"3E",X"F7",X"7C",X"C0",X"26",X"8F",X"07",X"8E",X"7F",X"31",X"20",X"40",X"00",X"11",X"0F",
		X"F2",X"7B",X"F0",X"E0",X"7F",X"06",X"BE",X"FF",X"F7",X"E7",X"FC",X"78",X"0E",X"40",X"80",X"00",
		X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"20",X"C8",X"F0",X"00",X"80",X"60",X"30",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"00",X"01",X"03",X"01",X"00",X"00",X"01",
		X"03",X"06",X"01",X"07",X"0E",X"0D",X"07",X"0F",X"07",X"03",X"01",X"00",X"03",X"0F",X"3E",X"F1",
		X"CF",X"A7",X"9D",X"0B",X"20",X"FD",X"E7",X"F3",X"C8",X"80",X"E0",X"F8",X"FB",X"B5",X"C2",X"16",
		X"F7",X"F8",X"D0",X"E2",X"FC",X"F4",X"38",X"F4",X"6A",X"FF",X"FF",X"7F",X"3C",X"CF",X"9E",X"23",
		X"E7",X"FD",X"5C",X"3E",X"37",X"7E",X"7C",X"3A",X"0F",X"7E",X"FC",X"F8",X"FC",X"78",X"10",X"C8",
		X"3B",X"81",X"00",X"00",X"00",X"80",X"01",X"02",X"00",X"00",X"00",X"00",X"C0",X"10",X"0E",X"07",
		X"80",X"D9",X"07",X"03",X"01",X"C0",X"85",X"C3",X"00",X"00",X"01",X"03",X"06",X"4C",X"1F",X"0D",
		X"F0",X"E3",X"87",X"E4",X"C8",X"E0",X"80",X"C1",X"FF",X"FF",X"FF",X"4C",X"00",X"00",X"11",X"E3",
		X"C1",X"FF",X"E9",X"3F",X"0F",X"19",X"30",X"E0",X"FC",X"FF",X"7F",X"3F",X"78",X"E0",X"E2",X"FC",
		X"80",X"C0",X"E0",X"E4",X"F8",X"E0",X"38",X"78",X"30",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"01",X"01",X"03",X"01",X"03",X"00",X"00",X"00",X"00",X"07",X"1F",X"7E",X"FC",X"5F",X"E7",
		X"F5",X"E3",X"C9",X"FE",X"7F",X"F3",X"F9",X"79",X"3C",X"FF",X"FB",X"B7",X"4F",X"07",X"27",X"C3",
		X"B7",X"FF",X"F9",X"F4",X"FC",X"F0",X"6C",X"FE",X"FF",X"FE",X"DF",X"8E",X"E3",X"C7",X"6F",X"9F",
		X"DF",X"FC",X"B0",X"F8",X"78",X"EC",X"78",X"FC",X"F8",X"F9",X"70",X"48",X"E0",X"E0",X"93",X"C7",
		X"DE",X"0F",X"00",X"00",X"06",X"0C",X"00",X"00",X"00",X"00",X"71",X"38",X"73",X"C0",X"80",X"00",
		X"0F",X"BE",X"7C",X"1E",X"0C",X"3F",X"1F",X"3F",X"7D",X"F8",X"FC",X"FE",X"1F",X"0F",X"9F",X"7F",
		X"C3",X"1C",X"7F",X"9F",X"0E",X"1C",X"FF",X"FF",X"EF",X"1E",X"3C",X"7F",X"FC",X"FE",X"DC",X"07",
		X"C0",X"E0",X"F0",X"F8",X"70",X"38",X"18",X"B8",X"E0",X"00",X"80",X"00",X"C0",X"00",X"40",X"80",
		X"01",X"07",X"1F",X"7F",X"FE",X"CE",X"97",X"FF",X"FE",X"E7",X"77",X"3B",X"FF",X"EF",X"9D",X"0E",
		X"DF",X"FF",X"BD",X"7E",X"7C",X"F9",X"FF",X"DD",X"EF",X"87",X"E3",X"FF",X"FF",X"32",X"9F",X"3E",
		X"F8",X"F8",X"D0",X"F0",X"F3",X"E4",X"E0",X"80",X"C0",X"80",X"C0",X"C0",X"87",X"03",X"0F",X"7C",
		X"00",X"31",X"18",X"70",X"C1",X"FB",X"03",X"03",X"41",X"C7",X"0F",X"07",X"1F",X"8F",X"00",X"01",
		X"7C",X"F1",X"F7",X"FF",X"FC",X"E7",X"DF",X"1F",X"87",X"CF",X"FF",X"F1",X"C3",X"EF",X"FF",X"FF",
		X"FE",X"FE",X"F8",X"F0",X"FC",X"3C",X"FC",X"FC",X"98",X"0C",X"FC",X"F0",X"C0",X"80",X"C0",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"03",X"0F",X"0F",X"07",
		X"00",X"00",X"00",X"00",X"01",X"06",X"0F",X"07",X"01",X"03",X"3F",X"F3",X"2F",X"FF",X"F4",X"9F",
		X"1F",X"1D",X"0F",X"7F",X"FF",X"CD",X"FF",X"5E",X"F3",X"FF",X"FD",X"FC",X"CC",X"F8",X"7C",X"10",
		X"FC",X"70",X"F8",X"D0",X"C0",X"80",X"C0",X"00",X"80",X"01",X"07",X"0C",X"00",X"00",X"00",X"00",
		X"06",X"0F",X"05",X"03",X"01",X"0B",X"07",X"0F",X"1D",X"3B",X"1F",X"3F",X"77",X"2F",X"65",X"FF",
		X"FF",X"FF",X"FF",X"AD",X"7D",X"7B",X"FF",X"FF",X"FF",X"F3",X"79",X"FF",X"FF",X"E7",X"F3",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0F",X"F0",X"A0",X"C3",X"41",X"03",X"07",X"05",X"03",
		X"07",X"03",X"1F",X"75",X"FF",X"7E",X"FF",X"28",X"3F",X"EF",X"FF",X"FB",X"7F",X"FF",X"DF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0D",X"1F",X"05",X"72",X"00",X"00",X"00",X"00",X"00",
		X"06",X"03",X"1F",X"6F",X"FF",X"7A",X"FC",X"54",X"F0",X"A0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"E0",X"41",X"87",X"83",X"06",X"0F",X"0B",X"07",X"0E",X"04",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"7D",X"DF",X"FF",X"F7",X"FF",X"ED",X"FA",X"55",X"FC",X"B0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"09",X"F1",X"A0",X"C0",X"42",X"01",X"00",X"01",X"00",
		X"07",X"33",X"5F",X"35",X"FF",X"7E",X"EC",X"40",X"3D",X"EF",X"7F",X"FB",X"7E",X"F5",X"D8",X"B0",
		X"0A",X"17",X"0F",X"1D",X"0B",X"01",X"00",X"00",X"37",X"5F",X"3A",X"55",X"08",X"00",X"00",X"00",
		X"50",X"E0",X"A0",X"80",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"EB",X"F6",X"C4",X"80",X"80",X"FF",X"FF",X"FF",X"3F",X"9F",X"47",X"63",X"F1",
		X"02",X"02",X"01",X"0F",X"07",X"00",X"00",X"18",X"78",X"71",X"E1",X"E3",X"F3",X"E7",X"E7",X"2F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"BE",X"5E",X"08",X"BC",X"B1",X"7F",X"7F",X"77",X"73",X"61",X"61",
		X"61",X"E0",X"F0",X"F8",X"B8",X"B0",X"C0",X"E1",X"FF",X"6F",X"1F",X"1E",X"3E",X"7C",X"FC",X"F8",
		X"EC",X"FF",X"2A",X"70",X"18",X"18",X"0C",X"0C",X"00",X"00",X"01",X"07",X"0F",X"0F",X"07",X"02",
		X"60",X"68",X"C8",X"98",X"9C",X"1C",X"3C",X"3E",X"21",X"6C",X"5E",X"76",X"FF",X"FF",X"DF",X"E7",
		X"F0",X"60",X"03",X"07",X"0F",X"3C",X"BD",X"FF",X"06",X"03",X"10",X"E1",X"C4",X"8F",X"80",X"80",
		X"00",X"00",X"F0",X"78",X"38",X"80",X"00",X"00",X"00",X"00",X"00",X"08",X"79",X"43",X"32",X"04",
		X"7E",X"7E",X"FF",X"DF",X"9F",X"0F",X"07",X"01",X"ED",X"7B",X"7F",X"3F",X"8F",X"C0",X"F0",X"FF",
		X"FC",X"FF",X"FF",X"FF",X"FF",X"FE",X"01",X"FE",X"C0",X"C0",X"E0",X"E0",X"C0",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"03",X"06",X"08",X"00",X"05",X"0F",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"0D",
		X"0E",X"0D",X"05",X"07",X"0D",X"0F",X"07",X"06",X"03",X"01",X"07",X"1E",X"7F",X"2B",X"84",X"C0",
		X"60",X"F8",X"C4",X"F1",X"31",X"C8",X"80",X"FC",X"F0",X"E0",X"B0",X"E0",X"31",X"80",X"05",X"03",
		X"69",X"7E",X"FF",X"CF",X"BC",X"19",X"3F",X"1F",X"1E",X"06",X"C0",X"60",X"11",X"82",X"C0",X"F0",
		X"A3",X"03",X"0F",X"17",X"C3",X"B4",X"E0",X"CE",X"7F",X"FF",X"1E",X"87",X"F3",X"C0",X"1E",X"3D",
		X"F9",X"60",X"D0",X"FC",X"38",X"74",X"70",X"E0",X"C0",X"F1",X"E6",X"D4",X"80",X"80",X"40",X"00",
		X"00",X"01",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"30",X"08",X"1E",X"0C",
		X"60",X"50",X"C0",X"A1",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"27",X"0F",X"03",X"06",X"1C",
		X"3C",X"22",X"00",X"40",X"F8",X"34",X"3E",X"7F",X"8F",X"19",X"80",X"00",X"80",X"02",X"3C",X"0F",
		X"40",X"00",X"00",X"23",X"1E",X"0F",X"3F",X"FD",X"F7",X"C3",X"07",X"0E",X"16",X"3E",X"7D",X"FF",
		X"0E",X"00",X"80",X"00",X"01",X"80",X"31",X"C3",X"EF",X"FF",X"18",X"00",X"00",X"00",X"F0",X"88",
		X"80",X"60",X"30",X"20",X"70",X"E0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"06",X"1F",X"0F",X"43",X"81",X"60",X"C6",X"80",X"09",X"87",X"02",X"00",
		X"0F",X"3E",X"FB",X"C4",X"E1",X"80",X"C2",X"F6",X"78",X"1C",X"7B",X"9F",X"3A",X"80",X"53",X"3F",
		X"EC",X"D7",X"0A",X"58",X"3F",X"4E",X"3B",X"1C",X"0E",X"4B",X"98",X"04",X"01",X"83",X"29",X"C7",
		X"F3",X"3D",X"78",X"8F",X"5E",X"3C",X"BF",X"6E",X"1F",X"1C",X"AC",X"76",X"F1",X"F0",X"FC",X"CE",
		X"BB",X"F0",X"40",X"20",X"80",X"40",X"80",X"00",X"01",X"86",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"20",X"18",X"0C",X"06",X"1C",X"20",X"C0",X"80",X"60",X"48",X"80",X"06",X"01",X"00",X"00",
		X"0C",X"98",X"3E",X"1B",X"60",X"00",X"01",X"00",X"13",X"0E",X"09",X"3C",X"70",X"E0",X"C8",X"70",
		X"00",X"00",X"23",X"C7",X"FF",X"7E",X"EF",X"F8",X"80",X"06",X"0F",X"07",X"8E",X"7F",X"31",X"20",
		X"78",X"E0",X"E2",X"FC",X"F2",X"7B",X"F0",X"E0",X"7F",X"06",X"BE",X"FF",X"EF",X"CF",X"FC",X"78",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"20",X"C8",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"02",X"03",X"01",X"00",X"00",X"01",X"0F",
		X"03",X"01",X"07",X"0F",X"1A",X"06",X"1C",X"38",X"37",X"3F",X"1F",X"3F",X"1F",X"0E",X"07",X"03",
		X"F0",X"7C",X"9F",X"3F",X"9F",X"7B",X"17",X"41",X"FB",X"9F",X"8C",X"CF",X"01",X"03",X"83",X"E1",
		X"1F",X"9D",X"0E",X"DF",X"E3",X"41",X"88",X"F0",X"F1",X"D1",X"E1",X"D0",X"A8",X"FD",X"FF",X"FF",
		X"1F",X"BF",X"7F",X"9E",X"FB",X"78",X"FC",X"EE",X"FD",X"B8",X"F8",X"F4",X"3E",X"FC",X"F8",X"F0",
		X"C1",X"27",X"8E",X"37",X"03",X"00",X"00",X"00",X"01",X"03",X"07",X"05",X"00",X"00",X"00",X"00",
		X"80",X"01",X"00",X"01",X"B3",X"0F",X"07",X"01",X"80",X"01",X"8B",X"07",X"01",X"01",X"03",X"07",
		X"07",X"0F",X"FE",X"F0",X"E3",X"87",X"E4",X"C8",X"80",X"C0",X"00",X"83",X"FF",X"FF",X"FF",X"4C",
		X"FE",X"DC",X"07",X"C1",X"FF",X"EF",X"39",X"1F",X"0F",X"1B",X"30",X"E0",X"FC",X"DF",X"7F",X"3F",
		X"00",X"40",X"80",X"80",X"C0",X"E0",X"E4",X"F8",X"E0",X"F0",X"38",X"78",X"30",X"E0",X"E0",X"C0",
		X"00",X"00",X"01",X"03",X"03",X"07",X"06",X"03",X"07",X"03",X"01",X"00",X"03",X"1F",X"7E",X"F9",
		X"7F",X"FE",X"EB",X"C7",X"93",X"3D",X"FF",X"FF",X"CF",X"E5",X"E7",X"73",X"FF",X"EF",X"DE",X"3F",
		X"3B",X"1C",X"6F",X"FF",X"F3",X"EB",X"F9",X"F8",X"E1",X"D8",X"FD",X"FF",X"FD",X"7E",X"3C",X"8F",
		X"3E",X"7C",X"BF",X"F8",X"60",X"F0",X"F0",X"F0",X"D8",X"F0",X"F8",X"F0",X"F2",X"E0",X"80",X"C0",
		X"1E",X"F8",X"BC",X"1F",X"00",X"00",X"04",X"08",X"1C",X"00",X"00",X"00",X"01",X"E3",X"71",X"E6",
		X"01",X"03",X"0F",X"BF",X"7E",X"38",X"0C",X"18",X"7F",X"3F",X"7F",X"FD",X"F0",X"F8",X"FC",X"1F",
		X"FF",X"FF",X"C3",X"1C",X"7F",X"9F",X"06",X"0C",X"1E",X"FF",X"FF",X"EF",X"1E",X"3C",X"7F",X"FC",
		X"C0",X"80",X"C0",X"E0",X"F0",X"F8",X"70",X"30",X"38",X"18",X"F0",X"E0",X"00",X"80",X"00",X"C0",
		X"1F",X"0F",X"03",X"0F",X"3F",X"FE",X"FC",X"9D",X"2F",X"FF",X"FD",X"CF",X"EE",X"67",X"FF",X"DE",
		X"38",X"BE",X"FF",X"FF",X"7B",X"FD",X"79",X"F3",X"FF",X"BB",X"DF",X"0F",X"C7",X"FF",X"FF",X"64",
		X"F0",X"30",X"F8",X"F0",X"A0",X"E0",X"E7",X"DC",X"C0",X"00",X"80",X"01",X"80",X"80",X"0E",X"07",
		X"00",X"00",X"01",X"63",X"31",X"61",X"E3",X"F7",X"07",X"07",X"83",X"87",X"0F",X"07",X"1F",X"0F",
		X"FF",X"FF",X"FF",X"F1",X"F7",X"FF",X"FC",X"E7",X"DF",X"1F",X"87",X"CF",X"FF",X"F1",X"C3",X"EF",
		X"FF",X"FF",X"FE",X"F8",X"F8",X"F0",X"F0",X"38",X"FC",X"FC",X"98",X"0C",X"FC",X"F0",X"C0",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"01",X"06",X"0F",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"03",X"0D",X"1F",X"0E",X"03",X"0F",X"7F",X"F3",X"6F",X"FF",X"EF",
		X"1E",X"3F",X"3A",X"1F",X"FF",X"FF",X"9B",X"FF",X"A6",X"F3",X"FF",X"FD",X"FC",X"CC",X"F8",X"FC",
		X"50",X"F8",X"E0",X"F0",X"A0",X"80",X"00",X"80",X"00",X"00",X"06",X"1C",X"38",X"00",X"00",X"00",
		X"07",X"0D",X"1D",X"0B",X"07",X"03",X"17",X"0E",X"1F",X"3B",X"77",X"3E",X"FF",X"6F",X"DF",X"CB",
		X"DF",X"FF",X"FF",X"FF",X"FD",X"DD",X"7B",X"7B",X"7F",X"FF",X"F3",X"F9",X"FF",X"FF",X"FF",X"E7",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"07",X"F0",X"E0",X"41",X"87",X"83",X"06",X"0F",X"0B",
		X"07",X"0F",X"07",X"3F",X"EA",X"FE",X"FC",X"FE",X"FF",X"7F",X"DF",X"FF",X"F7",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"06",X"05",X"07",X"03",X"01",X"00",
		X"40",X"00",X"04",X"28",X"78",X"73",X"6F",X"2E",X"3F",X"69",X"7E",X"3C",X"37",X"1F",X"0F",X"3F",
		X"24",X"1E",X"09",X"00",X"01",X"03",X"C3",X"27",X"8E",X"8D",X"40",X"01",X"E0",X"C0",X"80",X"C0",
		X"E8",X"00",X"02",X"4C",X"FF",X"26",X"F8",X"FC",X"7C",X"F3",X"E6",X"FF",X"FF",X"F3",X"37",X"00",
		X"81",X"07",X"0F",X"A7",X"1F",X"8F",X"0D",X"3F",X"5F",X"0C",X"D1",X"03",X"3B",X"FF",X"FF",X"7B",
		X"C4",X"C0",X"C0",X"F0",X"38",X"E4",X"80",X"00",X"F0",X"E0",X"D0",X"80",X"80",X"00",X"C4",X"98",
		X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"03",X"06",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"03",X"01",X"00",X"C0",X"20",X"80",X"43",X"01",X"00",X"00",X"00",X"01",X"00",X"07",
		X"E0",X"E1",X"C0",X"90",X"E0",X"78",X"44",X"00",X"80",X"F0",X"68",X"7C",X"FF",X"1F",X"33",X"00",
		X"0C",X"1F",X"FF",X"63",X"40",X"80",X"00",X"01",X"46",X"3C",X"1F",X"7E",X"FB",X"EF",X"83",X"07",
		X"FF",X"EF",X"C7",X"FC",X"F8",X"0E",X"00",X"00",X"00",X"02",X"01",X"61",X"83",X"EF",X"FF",X"18",
		X"00",X"00",X"C8",X"F0",X"00",X"80",X"60",X"30",X"20",X"E0",X"C0",X"C0",X"80",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"0F",X"1B",X"7E",X"3F",X"0F",X"05",X"80",X"19",X"02",
		X"FC",X"78",X"3E",X"1F",X"3E",X"FB",X"AC",X"10",X"84",X"01",X"08",X"98",X"60",X"71",X"EE",X"7C",
		X"06",X"0F",X"0F",X"87",X"32",X"5C",X"28",X"62",X"FC",X"38",X"EE",X"71",X"38",X"2C",X"62",X"11",
		X"A0",X"F6",X"FF",X"FF",X"CE",X"37",X"E1",X"0E",X"7A",X"F1",X"FE",X"B8",X"7C",X"72",X"B0",X"98",
		X"78",X"F0",X"E0",X"C0",X"E6",X"C0",X"00",X"80",X"00",X"00",X"00",X"01",X"07",X"18",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"41",X"30",X"18",X"1C",X"38",X"40",X"80",X"00",X"00",X"00",X"00",
		X"03",X"03",X"07",X"0E",X"18",X"30",X"78",X"33",X"E1",X"00",X"03",X"01",X"27",X"1C",X"12",X"78",
		X"E3",X"FF",X"FE",X"98",X"00",X"01",X"47",X"8F",X"FF",X"FE",X"DF",X"F0",X"00",X"0C",X"1F",X"0F",
		X"F8",X"BD",X"FF",X"7F",X"FF",X"E0",X"E2",X"FC",X"F2",X"7B",X"F0",X"E0",X"7F",X"06",X"7E",X"FD",
		X"70",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"0C",X"0F",X"1F",X"36",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"01",
		X"00",X"01",X"07",X"0F",X"01",X"1E",X"3C",X"6A",X"11",X"73",X"E0",X"C2",X"B7",X"FA",X"FC",X"D7",
		X"7F",X"FB",X"64",X"C0",X"F2",X"7C",X"FF",X"7F",X"FD",X"EE",X"5F",X"07",X"ED",X"7F",X"3F",X"37",
		X"9E",X"78",X"FF",X"1E",X"7B",X"3C",X"7F",X"8E",X"04",X"01",X"23",X"C3",X"C7",X"46",X"87",X"43",
		X"FD",X"79",X"3F",X"3F",X"7E",X"FF",X"3C",X"F6",X"E0",X"E0",X"F0",X"B8",X"F4",X"E0",X"E0",X"D0",
		X"C0",X"00",X"81",X"83",X"4E",X"1C",X"6E",X"07",X"00",X"00",X"00",X"00",X"03",X"06",X"0F",X"1F",
		X"C7",X"E3",X"CC",X"00",X"02",X"01",X"03",X"67",X"1F",X"0E",X"07",X"03",X"01",X"82",X"16",X"0F",
		X"B8",X"1C",X"1F",X"3F",X"1F",X"FC",X"E0",X"C3",X"17",X"0F",X"C8",X"90",X"00",X"80",X"00",X"01",
		X"3C",X"7F",X"FC",X"FE",X"DC",X"07",X"C1",X"FF",X"FF",X"DF",X"79",X"1F",X"0F",X"A3",X"60",X"C0",
		X"00",X"00",X"C0",X"00",X"40",X"80",X"80",X"C0",X"E0",X"C0",X"E4",X"F8",X"C0",X"B0",X"18",X"38",
		X"00",X"00",X"00",X"01",X"00",X"07",X"0F",X"0E",X"1C",X"1F",X"0F",X"1F",X"0F",X"07",X"00",X"0F",
		X"03",X"1F",X"FC",X"F8",X"CE",X"AF",X"3E",X"07",X"4F",X"F7",X"FF",X"9F",X"CB",X"8F",X"E7",X"F9",
		X"FF",X"BC",X"76",X"38",X"DF",X"FF",X"CF",X"07",X"D7",X"E3",X"E1",X"83",X"60",X"FB",X"FF",X"FB",
		X"FE",X"C8",X"7C",X"F8",X"7F",X"F4",X"F0",X"C0",X"60",X"E0",X"F0",X"E0",X"C0",X"F0",X"E0",X"E5",
		X"1C",X"0E",X"3C",X"F0",X"BA",X"1D",X"00",X"00",X"00",X"08",X"10",X"38",X"00",X"00",X"01",X"03",
		X"1F",X"0F",X"01",X"03",X"0F",X"BF",X"7E",X"3C",X"31",X"18",X"30",X"FC",X"7F",X"FF",X"F5",X"E0",
		X"0F",X"9F",X"FF",X"FF",X"C1",X"18",X"7F",X"F6",X"3F",X"0C",X"18",X"3E",X"FF",X"FF",X"8F",X"1E",
		X"C0",X"80",X"C0",X"80",X"C0",X"E0",X"F0",X"F0",X"F8",X"F0",X"30",X"28",X"18",X"F0",X"E0",X"00",
		X"1F",X"1E",X"0F",X"03",X"0F",X"3E",X"F9",X"F0",X"7B",X"3F",X"4F",X"FF",X"FB",X"9E",X"DD",X"CF",
		X"EF",X"78",X"7E",X"FF",X"FF",X"FE",X"E7",X"FB",X"73",X"E7",X"FF",X"76",X"BF",X"1E",X"8F",X"FF",
		X"FC",X"F0",X"38",X"F0",X"F0",X"40",X"E0",X"C3",X"DF",X"F3",X"80",X"00",X"01",X"01",X"00",X"00",
		X"00",X"20",X"00",X"01",X"63",X"31",X"E0",X"C1",X"6B",X"F7",X"07",X"07",X"82",X"87",X"0F",X"07",
		X"FF",X"7F",X"FF",X"FC",X"E1",X"F7",X"FF",X"FF",X"F0",X"E7",X"DF",X"1F",X"07",X"8E",X"FF",X"C7",
		X"FC",X"FE",X"FE",X"FC",X"F8",X"E0",X"F0",X"E0",X"F0",X"38",X"FC",X"FC",X"38",X"0C",X"FC",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"0C",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"03",X"0F",X"3B",X"7F",X"3C",X"0F",X"7F",X"FF",X"E7",X"DF",X"FF",
		X"0F",X"3C",X"FF",X"F5",X"7F",X"FF",X"FF",X"39",X"FF",X"A6",X"F3",X"FE",X"FE",X"FC",X"CC",X"F8",
		X"FC",X"A0",X"F0",X"C0",X"60",X"C0",X"80",X"00",X"80",X"00",X"00",X"0E",X"78",X"3C",X"00",X"00",
		X"07",X"02",X"01",X"00",X"05",X"03",X"07",X"0E",X"DD",X"8F",X"1F",X"3B",X"17",X"32",X"7F",X"7C",
		X"FF",X"D7",X"BD",X"BD",X"FB",X"FF",X"FF",X"6F",X"F9",X"7D",X"FF",X"FF",X"E7",X"F3",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"01",X"D0",X"E1",X"A0",X"81",X"03",X"82",X"01",X"03",
		X"07",X"1F",X"3F",X"1E",X"FF",X"D5",X"FC",X"F8",X"77",X"FF",X"FD",X"BF",X"FF",X"EF",X"FF",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"64",X"76",X"3E",X"0C",X"04",X"00",X"00",X"0C",X"1C",X"D8",X"78",X"70",X"10",X"00",X"00",
		X"01",X"01",X"03",X"03",X"07",X"06",X"06",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"82",X"1B",
		X"1F",X"3F",X"32",X"70",X"60",X"E0",X"C0",X"C0",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"06",X"07",X"06",X"0C",X"0C",X"1C",X"18",X"38",X"31",X"F1",X"E3",X"6B",X"07",X"06",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"30",X"73",X"63",X"E3",X"C6",X"C6",X"8E",X"8C",X"1C",X"38",
		X"38",X"30",X"20",X"60",X"60",X"E0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"07",X"06",X"06",X"0C",X"0C",X"1C",X"18",X"38",X"11",
		X"01",X"83",X"47",X"7F",X"3E",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"31",X"73",X"63",
		X"E3",X"C6",X"C6",X"8E",X"8C",X"9C",X"18",X"18",X"30",X"30",X"70",X"60",X"E0",X"C0",X"C0",X"80",
		X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"07",X"07",X"0C",X"0C",X"1C",X"18",X"38",
		X"30",X"70",X"60",X"E0",X"C0",X"40",X"00",X"00",X"38",X"F0",X"F0",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"0C",X"1C",X"18",X"18",X"30",X"30",X"70",X"60",X"E0",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"02",X"00",X"00",X"01",X"03",X"03",X"03",X"01",X"01",X"03",X"03",
		X"10",X"60",X"5C",X"F8",X"90",X"41",X"00",X"20",X"40",X"C0",X"98",X"7E",X"71",X"FC",X"4C",X"F2",
		X"15",X"01",X"01",X"67",X"09",X"23",X"F0",X"48",X"02",X"0F",X"18",X"1F",X"3E",X"73",X"6F",X"07",
		X"80",X"E0",X"C4",X"B9",X"F0",X"A2",X"00",X"10",X"62",X"FC",X"3A",X"80",X"C0",X"E1",X"98",X"36",
		X"C1",X"E1",X"B1",X"8A",X"46",X"07",X"1F",X"3F",X"9F",X"7C",X"3F",X"36",X"FD",X"7F",X"33",X"47",
		X"E0",X"F0",X"C8",X"C1",X"60",X"10",X"00",X"00",X"C0",X"E0",X"90",X"00",X"00",X"C0",X"80",X"40",
		X"0E",X"1C",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"17",X"0C",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"19",X"07",X"03",X"01",X"80",X"40",X"00",X"85",X"03",X"00",
		X"9F",X"78",X"24",X"40",X"F0",X"C0",X"C2",X"81",X"00",X"C0",X"F1",X"88",X"00",X"00",X"E0",X"D0",
		X"00",X"0C",X"3E",X"1F",X"0F",X"1C",X"3F",X"FF",X"C7",X"81",X"00",X"00",X"02",X"8C",X"78",X"3F",
		X"77",X"3E",X"06",X"7C",X"FE",X"FF",X"EF",X"C7",X"FC",X"F8",X"1E",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C8",X"F0",X"00",X"80",X"60",X"30",X"20",X"70",X"E0",
		X"06",X"03",X"03",X"07",X"03",X"01",X"00",X"00",X"00",X"03",X"0A",X"3C",X"6E",X"F8",X"FC",X"3E",
		X"DF",X"F9",X"F0",X"5C",X"F0",X"C0",X"F8",X"7E",X"F8",X"ED",X"B0",X"41",X"13",X"04",X"23",X"61",
		X"BB",X"ED",X"FE",X"D9",X"1A",X"3F",X"3F",X"1F",X"CB",X"70",X"A1",X"88",X"F0",X"E3",X"BB",X"C6",
		X"9F",X"2D",X"17",X"0F",X"81",X"D3",X"FF",X"FF",X"9D",X"6F",X"C2",X"19",X"F4",X"E2",X"FC",X"B0",
		X"E8",X"C0",X"C0",X"A0",X"F0",X"E0",X"C0",X"80",X"CC",X"89",X"00",X"00",X"00",X"00",X"00",X"03",
		X"06",X"0D",X"1E",X"34",X"00",X"00",X"00",X"00",X"00",X"02",X"C0",X"60",X"31",X"60",X"80",X"00",
		X"02",X"01",X"28",X"1E",X"07",X"07",X"0F",X"05",X"30",X"60",X"F0",X"67",X"C3",X"01",X"07",X"03",
		X"00",X"00",X"00",X"01",X"C7",X"FF",X"FE",X"38",X"01",X"07",X"8F",X"1F",X"FF",X"FC",X"FF",X"F0",
		X"07",X"A0",X"60",X"C0",X"F8",X"BD",X"FF",X"7F",X"F3",X"E0",X"C2",X"FC",X"F2",X"FB",X"F0",X"C0",
		X"80",X"30",X"18",X"38",X"70",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"03",X"07",
		X"00",X"00",X"00",X"00",X"07",X"1D",X"3F",X"07",X"40",X"59",X"F3",X"A1",X"07",X"4F",X"82",X"08",
		X"1E",X"03",X"1F",X"FF",X"EE",X"99",X"00",X"C9",X"F0",X"F0",X"EC",X"FE",X"D4",X"F0",X"64",X"1F",
		X"1F",X"8F",X"D3",X"1D",X"A0",X"FE",X"7C",X"F8",X"6C",X"F0",X"7D",X"29",X"13",X"07",X"8B",X"4F",
		X"77",X"FF",X"F7",X"FB",X"F0",X"3E",X"7F",X"FC",X"FC",X"7E",X"B8",X"AC",X"C0",X"C0",X"E0",X"30",
		X"E0",X"C0",X"DA",X"81",X"00",X"00",X"01",X"82",X"0C",X"18",X"6C",X"06",X"00",X"00",X"00",X"00",
		X"01",X"03",X"07",X"CF",X"E6",X"58",X"80",X"04",X"03",X"03",X"07",X"CF",X"3E",X"1C",X"0F",X"07",
		X"FF",X"E9",X"C0",X"78",X"1C",X"3F",X"7F",X"3D",X"FF",X"F8",X"41",X"87",X"2F",X"1F",X"90",X"20",
		X"FF",X"8F",X"1C",X"38",X"7F",X"FC",X"BE",X"FC",X"BF",X"0F",X"83",X"EF",X"FF",X"DF",X"79",X"1F",
		X"F0",X"E0",X"00",X"00",X"00",X"C0",X"00",X"40",X"80",X"00",X"00",X"80",X"80",X"E4",X"F8",X"40",
		X"00",X"00",X"00",X"00",X"01",X"07",X"07",X"03",X"1E",X"0C",X"38",X"71",X"6F",X"3F",X"7E",X"3F",
		X"03",X"01",X"0F",X"7F",X"F8",X"F0",X"9D",X"3F",X"9F",X"FD",X"1E",X"3F",X"DF",X"F3",X"7F",X"2E",
		X"BB",X"9F",X"FF",X"79",X"EC",X"71",X"3A",X"7F",X"FC",X"9F",X"0F",X"A6",X"C7",X"C3",X"07",X"C1",
		X"1E",X"FE",X"FC",X"90",X"F8",X"F0",X"FC",X"F7",X"E0",X"E0",X"80",X"C0",X"C0",X"E0",X"C0",X"80",
		X"00",X"00",X"1C",X"0E",X"1C",X"70",X"E0",X"74",X"3B",X"00",X"00",X"00",X"10",X"20",X"71",X"00",
		X"1F",X"3F",X"7E",X"3F",X"03",X"17",X"0F",X"1F",X"7C",X"F8",X"71",X"62",X"30",X"60",X"F8",X"FF",
		X"FF",X"8F",X"1F",X"3F",X"FF",X"FF",X"EF",X"03",X"30",X"FF",X"ED",X"3F",X"0E",X"1C",X"38",X"FF",
		X"BC",X"F0",X"C0",X"80",X"C0",X"80",X"C0",X"C0",X"E0",X"F0",X"F4",X"F8",X"F0",X"10",X"28",X"18",
		X"19",X"3F",X"3F",X"3C",X"1E",X"07",X"3F",X"FD",X"F3",X"E1",X"36",X"7F",X"9F",X"FC",X"F7",X"3C",
		X"BF",X"FF",X"DF",X"F0",X"FC",X"FF",X"FF",X"FC",X"CF",X"F7",X"A7",X"CF",X"FF",X"F4",X"7E",X"3C",
		X"98",X"F0",X"B8",X"E0",X"70",X"E0",X"E1",X"80",X"C3",X"9F",X"F6",X"03",X"00",X"00",X"01",X"03",
		X"01",X"01",X"00",X"61",X"03",X"01",X"C7",X"E3",X"C0",X"C1",X"93",X"EF",X"0E",X"0F",X"86",X"0F",
		X"EF",X"DF",X"C7",X"EF",X"FF",X"F8",X"E1",X"F7",X"7F",X"FF",X"F0",X"C7",X"1F",X"3F",X"07",X"8E",
		X"FE",X"FE",X"DC",X"8E",X"FE",X"FC",X"F8",X"E0",X"F0",X"E0",X"F0",X"38",X"FC",X"FC",X"38",X"0C",
		X"03",X"03",X"06",X"06",X"0C",X"0B",X"0F",X"07",X"00",X"00",X"01",X"00",X"00",X"00",X"03",X"0F",
		X"00",X"00",X"00",X"01",X"01",X"00",X"03",X"0F",X"36",X"FF",X"FF",X"F3",X"3F",X"FF",X"FF",X"CF",
		X"03",X"1F",X"79",X"FF",X"EB",X"FE",X"FF",X"FF",X"73",X"FF",X"4E",X"E3",X"FE",X"FE",X"FC",X"F8",
		X"F0",X"F8",X"40",X"E0",X"C0",X"60",X"C0",X"80",X"00",X"80",X"00",X"0C",X"1E",X"78",X"BC",X"00",
		X"06",X"0F",X"05",X"03",X"01",X"0B",X"07",X"0F",X"1D",X"3B",X"1F",X"3F",X"77",X"2F",X"65",X"FF",
		X"FF",X"FF",X"FF",X"AD",X"7D",X"7B",X"FF",X"FF",X"FF",X"F3",X"79",X"FF",X"FF",X"E7",X"F3",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"F0",X"A0",X"C3",X"41",X"03",X"07",X"05",X"03",
		X"01",X"0F",X"3F",X"7F",X"3D",X"FE",X"AA",X"F8",X"3F",X"EF",X"FF",X"FB",X"7F",X"FF",X"DF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"17",X"0C",X"02",X"00",X"01",X"0A",X"1E",X"1C",
		X"01",X"07",X"03",X"00",X"40",X"80",X"60",X"C1",X"86",X"80",X"09",X"07",X"02",X"00",X"00",X"C0",
		X"B8",X"E0",X"F4",X"F8",X"51",X"0A",X"07",X"87",X"1E",X"0E",X"80",X"40",X"13",X"7F",X"C1",X"C1",
		X"07",X"0F",X"13",X"CE",X"87",X"03",X"83",X"12",X"E6",X"80",X"00",X"00",X"12",X"E1",X"D0",X"C0",
		X"C3",X"C7",X"8F",X"EF",X"1A",X"07",X"87",X"C7",X"2D",X"1C",X"1C",X"7C",X"FF",X"73",X"FE",X"D8",
		X"D0",X"88",X"F0",X"C0",X"80",X"C0",X"20",X"01",X"80",X"40",X"00",X"00",X"00",X"80",X"40",X"00",
		X"00",X"01",X"02",X"0C",X"18",X"38",X"70",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"80",X"00",X"00",X"00",X"01",X"00",X"00",X"04",X"03",X"07",X"67",X"1E",X"0F",X"07",X"03",
		X"07",X"03",X"01",X"07",X"03",X"1E",X"F8",X"44",X"80",X"E0",X"00",X"04",X"03",X"81",X"C1",X"F2",
		X"FF",X"FF",X"B9",X"FF",X"81",X"00",X"18",X"78",X"3C",X"3F",X"79",X"7F",X"FF",X"01",X"01",X"00",
		X"78",X"E4",X"F6",X"E4",X"01",X"F6",X"7C",X"0C",X"FC",X"FE",X"CF",X"9F",X"0F",X"FC",X"F8",X"1E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C8",X"F0",X"00",X"00",
		X"00",X"15",X"1E",X"1C",X"1B",X"0F",X"0F",X"1D",X"0F",X"07",X"03",X"01",X"03",X"0F",X"2A",X"F1",
		X"24",X"1E",X"09",X"20",X"7E",X"E5",X"C3",X"73",X"A0",X"00",X"E0",X"F8",X"E3",X"B5",X"C0",X"02",
		X"50",X"C0",X"12",X"7D",X"EE",X"B4",X"F8",X"64",X"6A",X"FF",X"FF",X"7F",X"2E",X"C1",X"87",X"20",
		X"4F",X"1F",X"2F",X"3C",X"7F",X"B7",X"1F",X"3E",X"07",X"4F",X"FF",X"FE",X"77",X"BE",X"08",X"60",
		X"00",X"00",X"80",X"C0",X"A0",X"00",X"00",X"80",X"C0",X"80",X"00",X"00",X"34",X"23",X"00",X"01",
		X"01",X"00",X"00",X"00",X"0C",X"1A",X"3C",X"68",X"00",X"00",X"00",X"00",X"00",X"84",X"C0",X"E0",
		X"9C",X"78",X"32",X"1C",X"0F",X"08",X"50",X"3E",X"0D",X"1F",X"23",X"06",X"00",X"00",X"00",X"0F",
		X"47",X"3F",X"18",X"10",X"20",X"80",X"04",X"03",X"07",X"8F",X"FD",X"70",X"03",X"05",X"8F",X"0F",
		X"BF",X"F3",X"7E",X"1C",X"07",X"40",X"80",X"80",X"E4",X"78",X"FD",X"FF",X"E3",X"C0",X"80",X"84",
		X"80",X"E4",X"78",X"00",X"40",X"30",X"18",X"10",X"38",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"06",
		X"00",X"01",X"00",X"00",X"00",X"00",X"07",X"1F",X"37",X"7E",X"3C",X"9F",X"03",X"67",X"C7",X"83",
		X"FF",X"F9",X"FC",X"7C",X"0E",X"FE",X"FC",X"B8",X"61",X"07",X"01",X"A7",X"C3",X"E1",X"DC",X"F8",
		X"CF",X"FC",X"BB",X"7D",X"3F",X"CF",X"67",X"B3",X"83",X"F8",X"F1",X"E3",X"B6",X"C1",X"F6",X"A6",
		X"0F",X"1F",X"07",X"DF",X"FF",X"9F",X"EE",X"C0",X"F8",X"F0",X"FC",X"F2",X"F0",X"F8",X"E4",X"B0",
		X"C0",X"80",X"00",X"C0",X"80",X"34",X"03",X"01",X"00",X"03",X"04",X"18",X"30",X"DC",X"0E",X"00",
		X"62",X"F1",X"00",X"03",X"07",X"0F",X"9E",X"CC",X"B0",X"00",X"00",X"00",X"04",X"03",X"02",X"0F",
		X"E0",X"F0",X"FF",X"FF",X"D3",X"80",X"C4",X"78",X"3F",X"1F",X"7B",X"3E",X"E0",X"93",X"47",X"03",
		X"30",X"E0",X"FC",X"FF",X"1F",X"3E",X"78",X"FF",X"FC",X"3E",X"FC",X"78",X"1F",X"03",X"DF",X"FF",
		X"38",X"58",X"30",X"E0",X"C0",X"80",X"80",X"00",X"80",X"C0",X"00",X"40",X"80",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"1F",X"1E",X"0C",X"7A",X"33",X"E0",X"C4",X"BF",
		X"3F",X"1C",X"0E",X"03",X"1F",X"7E",X"F1",X"E0",X"C1",X"74",X"FD",X"7F",X"F6",X"78",X"FE",X"7F",
		X"EE",X"F8",X"76",X"BF",X"FF",X"F3",X"DB",X"E1",X"E3",X"F5",X"CF",X"F3",X"7F",X"3F",X"9D",X"1F",
		X"FE",X"7C",X"3E",X"FC",X"F8",X"20",X"E0",X"F0",X"E0",X"F9",X"EE",X"C0",X"C0",X"00",X"80",X"80",
		X"03",X"06",X"00",X"40",X"1C",X"0E",X"1C",X"30",X"E0",X"C0",X"E8",X"74",X"03",X"01",X"00",X"10",
		X"0C",X"1F",X"3F",X"7E",X"F8",X"7E",X"0F",X"07",X"4F",X"3F",X"7C",X"F9",X"E3",X"F2",X"E0",X"78",
		X"0E",X"1C",X"FF",X"FF",X"1F",X"3F",X"FF",X"FF",X"DE",X"07",X"61",X"FF",X"F6",X"3F",X"0F",X"19",
		X"70",X"18",X"B8",X"E0",X"80",X"10",X"C0",X"00",X"40",X"80",X"80",X"C0",X"E0",X"E4",X"F8",X"E0",
		X"0F",X"19",X"33",X"7F",X"7F",X"79",X"3D",X"0F",X"7F",X"FB",X"E7",X"C3",X"6D",X"FF",X"3F",X"FC",
		X"CF",X"DF",X"FF",X"F7",X"BB",X"E1",X"F8",X"FF",X"FF",X"F9",X"9F",X"E7",X"4F",X"97",X"FF",X"EC",
		X"DC",X"38",X"F8",X"60",X"F0",X"E0",X"F0",X"F0",X"E3",X"C1",X"C7",X"BF",X"ED",X"07",X"00",X"00",
		X"BC",X"01",X"03",X"03",X"01",X"63",X"07",X"03",X"8F",X"C7",X"80",X"81",X"27",X"DF",X"3C",X"1E",
		X"FC",X"EF",X"DF",X"9F",X"C7",X"EF",X"FF",X"F8",X"E1",X"F7",X"FF",X"FF",X"C3",X"1C",X"7F",X"9F",
		X"FC",X"7E",X"FE",X"FE",X"CC",X"86",X"FE",X"FC",X"F0",X"C0",X"E0",X"C0",X"E0",X"F0",X"F8",X"F8",
		X"00",X"01",X"07",X"0F",X"1C",X"1C",X"39",X"17",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"03",
		X"00",X"00",X"00",X"01",X"03",X"03",X"01",X"07",X"1F",X"6C",X"FF",X"FE",X"E7",X"37",X"FF",X"FF",
		X"1F",X"07",X"7F",X"B3",X"FF",X"D7",X"FE",X"FF",X"FF",X"F2",X"FF",X"9E",X"C7",X"FE",X"FE",X"B4",
		X"F0",X"E0",X"F0",X"40",X"E0",X"C0",X"70",X"C0",X"00",X"00",X"80",X"00",X"00",X"0C",X"1E",X"78",
		X"07",X"0D",X"1D",X"0B",X"07",X"03",X"17",X"0E",X"1F",X"3B",X"77",X"3E",X"FF",X"6F",X"DF",X"CB",
		X"DF",X"FF",X"FF",X"FF",X"FD",X"DD",X"7B",X"7B",X"7F",X"FF",X"F3",X"F9",X"FF",X"FF",X"FF",X"E7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0F",X"F0",X"E0",X"41",X"87",X"83",X"06",X"0F",X"0B",
		X"07",X"01",X"1F",X"7F",X"FF",X"7A",X"FC",X"54",X"FF",X"7F",X"DF",X"FF",X"F7",X"FF",X"FF",X"FF",
		X"06",X"06",X"0C",X"0C",X"1C",X"18",X"38",X"11",X"E3",X"C6",X"F6",X"9E",X"9C",X"84",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"06",X"06",X"0C",X"0C",X"1C",X"98",X"78",X"71",X"35",X"03",X"03",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"03",X"13",X"26",X"26",X"46",X"4C",X"CC",X"8C",X"98",X"18",X"18",
		X"30",X"30",X"30",X"60",X"60",X"60",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"03",X"03",X"03",X"06",X"06",X"0E",X"0C",X"04",X"00",X"00",X"00",X"08",X"0C",X"1C",X"18",X"38",
		X"30",X"70",X"60",X"60",X"C0",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"04",X"04",X"08",X"08",X"18",X"18",X"30",X"31",X"31",
		X"00",X"00",X"00",X"20",X"30",X"30",X"22",X"63",X"47",X"46",X"4E",X"8C",X"8C",X"98",X"18",X"38",
		X"30",X"70",X"60",X"60",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"01",X"01",X"02",X"02",X"04",
		X"01",X"83",X"43",X"77",X"3E",X"1E",X"04",X"00",X"E3",X"C6",X"F6",X"9E",X"9C",X"84",X"00",X"00",
		X"20",X"30",X"70",X"60",X"E0",X"C0",X"C0",X"80",X"F3",X"E3",X"7B",X"0E",X"0E",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"12",X"1B",X"3F",X"36",X"72",X"60",X"60",X"C0",X"00",X"00",X"20",
		X"B0",X"F0",X"60",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
