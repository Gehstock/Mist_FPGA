library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity monitor is
    generic(
        AddrWidth   : integer := 14
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(AddrWidth-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end monitor;

architecture rtl of monitor is
    type rom16384x8 is array (0 to 2**AddrWidth-1) of std_logic_vector(7 downto 0); 
    constant romData : rom16384x8 := (
         x"31",  x"c0",  x"eb",  x"21",  x"78",  x"00",  x"11",  x"00", -- 0000
         x"f0",  x"cd",  x"2c",  x"00",  x"21",  x"ba",  x"0e",  x"11", -- 0008
         x"00",  x"c0",  x"cd",  x"2c",  x"00",  x"21",  x"5b",  x"31", -- 0010
         x"11",  x"00",  x"80",  x"cd",  x"2c",  x"00",  x"01",  x"07", -- 0018
         x"00",  x"11",  x"00",  x"ec",  x"21",  x"71",  x"00",  x"ed", -- 0020
         x"b0",  x"c3",  x"00",  x"ec",  x"3e",  x"80",  x"ed",  x"a0", -- 0028
         x"cd",  x"6b",  x"00",  x"30",  x"f9",  x"d5",  x"01",  x"00", -- 0030
         x"00",  x"50",  x"14",  x"cd",  x"6b",  x"00",  x"30",  x"fa", -- 0038
         x"d4",  x"6b",  x"00",  x"cb",  x"11",  x"cb",  x"10",  x"38", -- 0040
         x"1f",  x"15",  x"20",  x"f4",  x"03",  x"5e",  x"23",  x"cb", -- 0048
         x"33",  x"30",  x"0c",  x"16",  x"10",  x"cd",  x"6b",  x"00", -- 0050
         x"cb",  x"12",  x"30",  x"f9",  x"14",  x"cb",  x"3a",  x"cb", -- 0058
         x"1b",  x"e3",  x"e5",  x"ed",  x"52",  x"d1",  x"ed",  x"b0", -- 0060
         x"e1",  x"30",  x"c5",  x"87",  x"c0",  x"7e",  x"23",  x"17", -- 0068
         x"c9",  x"3e",  x"05",  x"d3",  x"02",  x"c3",  x"00",  x"f0", -- 0070
         x"c3",  x"0c",  x"64",  x"f6",  x"c3",  x"ae",  x"02",  x"56", -- 0078
         x"f7",  x"36",  x"c3",  x"7f",  x"02",  x"83",  x"02",  x"9e", -- 0080
         x"db",  x"02",  x"ae",  x"02",  x"a8",  x"02",  x"60",  x"c4", -- 0088
         x"02",  x"de",  x"f5",  x"c3",  x"0b",  x"f8",  x"36",  x"c3", -- 0090
         x"fc",  x"08",  x"df",  x"02",  x"34",  x"1b",  x"f4",  x"c3", -- 0098
         x"6f",  x"02",  x"a4",  x"08",  x"69",  x"33",  x"02",  x"37", -- 00A0
         x"1b",  x"1a",  x"d2",  x"05",  x"d9",  x"02",  x"66",  x"e5", -- 00A8
         x"02",  x"f4",  x"f7",  x"43",  x"09",  x"00",  x"f0",  x"0c", -- 00B0
         x"f0",  x"15",  x"f0",  x"12",  x"f0",  x"0f",  x"00",  x"f0", -- 00B8
         x"18",  x"f0",  x"39",  x"f0",  x"3c",  x"f0",  x"e2",  x"00", -- 00C0
         x"f3",  x"65",  x"f3",  x"06",  x"f0",  x"f3",  x"f3",  x"f8", -- 00C8
         x"00",  x"f3",  x"2d",  x"f4",  x"45",  x"f4",  x"6a",  x"f4", -- 00D0
         x"3c",  x"18",  x"f7",  x"3b",  x"f7",  x"33",  x"27",  x"f0", -- 00D8
         x"2a",  x"00",  x"f0",  x"1e",  x"f0",  x"21",  x"f0",  x"a8", -- 00E0
         x"f4",  x"e3",  x"00",  x"fa",  x"24",  x"f0",  x"3f",  x"f0", -- 00E8
         x"42",  x"f0",  x"3e",  x"06",  x"f7",  x"3d",  x"f7",  x"b9", -- 00F0
         x"f5",  x"19",  x"d8",  x"00",  x"f4",  x"21",  x"89",  x"f0", -- 00F8
         x"e5",  x"21",  x"80",  x"00",  x"00",  x"22",  x"1b",  x"00", -- 0100
         x"3e",  x"3e",  x"cd",  x"05",  x"f3",  x"03",  x"cd",  x"5c", -- 0108
         x"f3",  x"38",  x"23",  x"cd",  x"1a",  x"00",  x"d8",  x"21", -- 0110
         x"ea",  x"f5",  x"e5",  x"cd",  x"ea",  x"f1",  x"00",  x"ca", -- 0118
         x"e6",  x"f5",  x"c5",  x"cd",  x"8e",  x"f2",  x"c1",  x"0c", -- 0120
         x"28",  x"07",  x"cd",  x"26",  x"14",  x"2a",  x"71",  x"00", -- 0128
         x"00",  x"e9",  x"08",  x"30",  x"2a",  x"cd",  x"fe",  x"f2", -- 0130
         x"60",  x"da",  x"bc",  x"06",  x"00",  x"04",  x"21",  x"e9", -- 0138
         x"ef",  x"11",  x"d5",  x"fb",  x"cd",  x"ca",  x"74",  x"3e", -- 0140
         x"3a",  x"3a",  x"07",  x"d5",  x"5e",  x"23",  x"56",  x"23", -- 0148
         x"33",  x"8e",  x"0d",  x"e1",  x"d1",  x"13",  x"00",  x"85", -- 0150
         x"23",  x"10",  x"e5",  x"c9",  x"05",  x"41",  x"28",  x"2c", -- 0158
         x"08",  x"da",  x"1d",  x"44",  x"01",  x"09",  x"2e",  x"00", -- 0160
         x"2b",  x"b8",  x"f2",  x"58",  x"c1",  x"20",  x"50",  x"3e", -- 0168
         x"06",  x"04",  x"93",  x"87",  x"32",  x"33",  x"74",  x"40", -- 0170
         x"00",  x"00",  x"79",  x"fe",  x"3a",  x"20",  x"05",  x"cd", -- 0178
         x"c4",  x"02",  x"f1",  x"fe",  x"3d",  x"c2",  x"e2",  x"f5", -- 0180
         x"da",  x"2d",  x"5b",  x"6e",  x"b2",  x"80",  x"6e",  x"17", -- 0188
         x"cd",  x"ab",  x"f0",  x"d8",  x"00",  x"00",  x"e5",  x"d5", -- 0190
         x"7c",  x"84",  x"85",  x"87",  x"16",  x"00",  x"00",  x"5f", -- 0198
         x"21",  x"c9",  x"ef",  x"19",  x"71",  x"23",  x"70",  x"06", -- 01A0
         x"d1",  x"e1",  x"3a",  x"04",  x"00",  x"80",  x"06",  x"37", -- 01A8
         x"3a",  x"3b",  x"47",  x"00",  x"4d",  x"bc",  x"28",  x"0a", -- 01B0
         x"95",  x"3c",  x"fe",  x"06",  x"00",  x"28",  x"04",  x"3d", -- 01B8
         x"b8",  x"20",  x"25",  x"d5",  x"58",  x"60",  x"21",  x"19", -- 01C0
         x"06",  x"09",  x"3c",  x"cb",  x"1e",  x"07",  x"3d",  x"20", -- 01C8
         x"07",  x"cb",  x"39",  x"06",  x"80",  x"03",  x"05",  x"10", -- 01D0
         x"f2",  x"43",  x"cd",  x"ce",  x"f2",  x"07",  x"d1",  x"30", -- 01D8
         x"0b",  x"08",  x"32",  x"1b",  x"8c",  x"72",  x"37",  x"c9", -- 01E0
         x"c3",  x"87",  x"18",  x"2a",  x"72",  x"73",  x"23",  x"72", -- 01E8
         x"00",  x"c3",  x"bd",  x"f0",  x"08",  x"38",  x"34",  x"06", -- 01F0
         x"03",  x"07",  x"3e",  x"17",  x"32",  x"2f",  x"00",  x"70", -- 01F8
         x"e0",  x"76",  x"93",  x"e3",  x"18",  x"d8",  x"5f",  x"3a", -- 0200
         x"0b",  x"bb",  x"3e",  x"03",  x"0c",  x"d8",  x"4d",  x"6c", -- 0208
         x"63",  x"1c",  x"10",  x"3e",  x"0c",  x"3b",  x"10",  x"e3", -- 0210
         x"c3",  x"92",  x"0c",  x"22",  x"1e",  x"a2",  x"01",  x"32", -- 0218
         x"1d",  x"00",  x"b7",  x"c9",  x"b0",  x"07",  x"08",  x"cf", -- 0220
         x"c4",  x"e4",  x"11",  x"01",  x"31",  x"01",  x"cd",  x"c6", -- 0228
         x"a0",  x"e4",  x"60",  x"c3",  x"df",  x"21",  x"00",  x"81", -- 0230
         x"00",  x"23",  x"7e",  x"fe",  x"20",  x"28",  x"fa",  x"00", -- 0238
         x"cd",  x"d7",  x"f1",  x"4f",  x"c0",  x"fe",  x"01",  x"d8", -- 0240
         x"00",  x"bf",  x"c9",  x"7e",  x"b7",  x"c8",  x"e5",  x"c5", -- 0248
         x"21",  x"00",  x"ab",  x"fc",  x"01",  x"05",  x"00",  x"ed", -- 0250
         x"b1",  x"c1",  x"00",  x"e1",  x"36",  x"20",  x"23",  x"c9", -- 0258
         x"11",  x"52",  x"01",  x"00",  x"af",  x"06",  x"51",  x"12", -- 0260
         x"1b",  x"10",  x"fc",  x"e5",  x"a0",  x"e7",  x"01",  x"38", -- 0268
         x"0d",  x"28",  x"0b",  x"12",  x"04",  x"13",  x"40",  x"31", -- 0270
         x"20",  x"f8",  x"cd",  x"d0",  x"f1",  x"00",  x"78",  x"32", -- 0278
         x"00",  x"01",  x"79",  x"e1",  x"08",  x"3a",  x"c3",  x"55", -- 0280
         x"fe",  x"30",  x"38",  x"16",  x"8b",  x"13",  x"30",  x"12", -- 0288
         x"3e",  x"63",  x"11",  x"12",  x"cd",  x"15",  x"f8",  x"3c", -- 0290
         x"35",  x"38",  x"02",  x"4f",  x"bf",  x"00",  x"82",  x"fe", -- 0298
         x"40",  x"38",  x"61",  x"f8",  x"bb",  x"86",  x"17",  x"cd", -- 02A0
         x"4d",  x"f2",  x"f5",  x"d5",  x"04",  x"18",  x"06",  x"a1", -- 02A8
         x"09",  x"cd",  x"69",  x"f2",  x"f1",  x"83",  x"23",  x"f5", -- 02B0
         x"b7",  x"ed",  x"52",  x"f1",  x"62",  x"18",  x"00",  x"04", -- 02B8
         x"af",  x"07",  x"3c",  x"30",  x"fb",  x"03",  x"21",  x"c1", -- 02C0
         x"ef",  x"d6",  x"08",  x"23",  x"07",  x"06",  x"c6",  x"08", -- 02C8
         x"2b",  x"28",  x"fb",  x"8d",  x"20",  x"cb",  x"16",  x"3d", -- 02D0
         x"c8",  x"10",  x"62",  x"fa",  x"3a",  x"d5",  x"eb",  x"1a", -- 02D8
         x"81",  x"a6",  x"04",  x"e0",  x"48",  x"52",  x"e6",  x"df", -- 02E0
         x"be",  x"13",  x"23",  x"00",  x"20",  x"0c",  x"10",  x"ee", -- 02E8
         x"d1",  x"d1",  x"6b",  x"62",  x"03",  x"2b",  x"7e",  x"2b", -- 02F0
         x"6e",  x"67",  x"c9",  x"d4",  x"11",  x"c9",  x"21",  x"00", -- 02F8
         x"80",  x"9c",  x"3e",  x"c3",  x"ed",  x"06",  x"a1",  x"20", -- 0300
         x"12",  x"23",  x"23",  x"a9",  x"4d",  x"0b",  x"7f",  x"b8", -- 0308
         x"44",  x"82",  x"0c",  x"00",  x"af",  x"2b",  x"2b",  x"be", -- 0310
         x"20",  x"e8",  x"e1",  x"25",  x"c4",  x"9b",  x"24",  x"c9", -- 0318
         x"00",  x"c1",  x"c9",  x"01",  x"06",  x"02",  x"21",  x"26", -- 0320
         x"fc",  x"a0",  x"ff",  x"19",  x"c5",  x"41",  x"05",  x"b1", -- 0328
         x"31",  x"6c",  x"20",  x"c8",  x"79",  x"23",  x"88",  x"eb", -- 0330
         x"fc",  x"10",  x"f0",  x"0c",  x"f6",  x"01",  x"c9",  x"f5", -- 0338
         x"a2",  x"85",  x"58",  x"78",  x"b7",  x"16",  x"9b",  x"64", -- 0340
         x"cb",  x"60",  x"3f",  x"e8",  x"cb",  x"0b",  x"23",  x"e6", -- 0348
         x"03",  x"83",  x"b3",  x"20",  x"f1",  x"19",  x"19",  x"e5", -- 0350
         x"a3",  x"95",  x"00",  x"21",  x"ff",  x"ff",  x"eb",  x"cd", -- 0358
         x"bc",  x"fc",  x"d1",  x"50",  x"3f",  x"8a",  x"00",  x"c5", -- 0360
         x"ed",  x"b0",  x"18",  x"0e",  x"3e",  x"0d",  x"a3",  x"af", -- 0368
         x"28",  x"3e",  x"0a",  x"0d",  x"4f",  x"cd",  x"d1",  x"fc", -- 0370
         x"c1",  x"40",  x"81",  x"3e",  x"00",  x"20",  x"18",  x"f1", -- 0378
         x"ed",  x"73",  x"0b",  x"00",  x"31",  x"0c",  x"c0",  x"01", -- 0380
         x"37",  x"3f",  x"17",  x"f5",  x"ed",  x"00",  x"43",  x"0d", -- 0388
         x"00",  x"32",  x"0f",  x"00",  x"21",  x"45",  x"60",  x"f3", -- 0390
         x"98",  x"21",  x"34",  x"b9",  x"da",  x"a9",  x"50",  x"06", -- 0398
         x"0b",  x"f0",  x"09",  x"09",  x"01",  x"7e",  x"23",  x"66", -- 03A0
         x"6f",  x"4b",  x"42",  x"3a",  x"81",  x"19",  x"e5",  x"2e", -- 03A8
         x"03",  x"c9",  x"30",  x"06",  x"90",  x"ba",  x"f5",  x"f1", -- 03B0
         x"37",  x"fa",  x"02",  x"40",  x"11",  x"33",  x"ed",  x"4b", -- 03B8
         x"32",  x"ed",  x"7b",  x"42",  x"c7",  x"8e",  x"ce",  x"41", -- 03C0
         x"3e",  x"50",  x"12",  x"58",  x"11",  x"e1",  x"03",  x"23", -- 03C8
         x"4d",  x"44",  x"03",  x"36",  x"48",  x"79",  x"35",  x"2e", -- 03D0
         x"6a",  x"cd",  x"7f",  x"6d",  x"69",  x"d8",  x"ed",  x"00", -- 03D8
         x"17",  x"00",  x"34",  x"35",  x"e1",  x"20",  x"03",  x"2b", -- 03E0
         x"fe",  x"03",  x"20",  x"03",  x"af",  x"d8",  x"10",  x"fe", -- 03E8
         x"1f",  x"28",  x"1b",  x"33",  x"fe",  x"02",  x"b4",  x"00", -- 03F0
         x"cd",  x"c6",  x"f3",  x"20",  x"fb",  x"18",  x"d7",  x"fe", -- 03F8
         x"c8",  x"a0",  x"20",  x"fe",  x"00",  x"0b",  x"28",  x"cf", -- 0400
         x"fe",  x"0a",  x"28",  x"cb",  x"fe",  x"52",  x"08",  x"9b", -- 0408
         x"60",  x"16",  x"18",  x"c2",  x"fe",  x"10",  x"28",  x"0a", -- 0410
         x"03",  x"34",  x"02",  x"03",  x"b4",  x"03",  x"d8",  x"1a", -- 0418
         x"92",  x"11",  x"b3",  x"3a",  x"35",  x"61",  x"9b",  x"47", -- 0420
         x"81",  x"83",  x"47",  x"c8",  x"0b",  x"0a",  x"fe",  x"09", -- 0428
         x"aa",  x"1c",  x"de",  x"42",  x"38",  x"f4",  x"3e",  x"08", -- 0430
         x"d4",  x"bf",  x"10",  x"f3",  x"90",  x"07",  x"35",  x"c9", -- 0438
         x"07",  x"1a",  x"b7",  x"20",  x"06",  x"3a",  x"6a",  x"9a", -- 0440
         x"90",  x"af",  x"c0",  x"36",  x"13",  x"18",  x"ef",  x"21", -- 0448
         x"03",  x"01",  x"03",  x"18",  x"38",  x"cd",  x"93",  x"f5", -- 0450
         x"3c",  x"82",  x"00",  x"af",  x"32",  x"6c",  x"00",  x"6c", -- 0458
         x"cd",  x"da",  x"e1",  x"a5",  x"f5",  x"d9",  x"0c",  x"11", -- 0460
         x"be",  x"0c",  x"19",  x"11",  x"6d",  x"f4",  x"98",  x"08", -- 0468
         x"bd",  x"06",  x"b0",  x"d1",  x"21",  x"5c",  x"c5",  x"8a", -- 0470
         x"0b",  x"dd",  x"1c",  x"a1",  x"42",  x"37",  x"c0",  x"3a", -- 0478
         x"73",  x"86",  x"3d",  x"32",  x"c0",  x"ef",  x"9e",  x"5b", -- 0480
         x"1d",  x"22",  x"db",  x"0d",  x"cc",  x"76",  x"ad",  x"53", -- 0488
         x"d8",  x"31",  x"21",  x"3b",  x"2b",  x"34",  x"f5",  x"67", -- 0490
         x"f7",  x"29",  x"6a",  x"4c",  x"32",  x"db",  x"bd",  x"92", -- 0498
         x"0c",  x"2e",  x"01",  x"70",  x"6d",  x"17",  x"5a",  x"6b", -- 04A0
         x"0b",  x"02",  x"69",  x"5f",  x"72",  x"31",  x"5f",  x"d9", -- 04A8
         x"7b",  x"ff",  x"11",  x"18",  x"a0",  x"5c",  x"6d",  x"5b", -- 04B0
         x"0c",  x"3a",  x"4c",  x"b7",  x"91",  x"a2",  x"3e",  x"09", -- 04B8
         x"83",  x"f5",  x"2a",  x"95",  x"11",  x"d5",  x"11",  x"7f", -- 04C0
         x"94",  x"14",  x"52",  x"d1",  x"98",  x"59",  x"89",  x"19", -- 04C8
         x"38",  x"ed",  x"a0",  x"0d",  x"3b",  x"f2",  x"30",  x"a1", -- 04D0
         x"0b",  x"d6",  x"fe",  x"61",  x"d8",  x"30",  x"7e",  x"e0", -- 04D8
         x"6d",  x"65",  x"c3",  x"ae",  x"cd",  x"d5",  x"01",  x"fc", -- 04E0
         x"06",  x"16",  x"03",  x"21",  x"f5",  x"40",  x"e5",  x"2b", -- 04E8
         x"36",  x"3a",  x"23",  x"30",  x"0a",  x"c5",  x"3e",  x"07", -- 04F0
         x"47",  x"af",  x"c6",  x"00",  x"01",  x"27",  x"10",  x"fb", -- 04F8
         x"77",  x"3e",  x"33",  x"ed",  x"0c",  x"67",  x"23",  x"77", -- 0500
         x"23",  x"48",  x"c1",  x"03",  x"1b",  x"15",  x"20",  x"e2", -- 0508
         x"f4",  x"02",  x"0e",  x"08",  x"c3",  x"f7",  x"f2",  x"a4", -- 0510
         x"57",  x"56",  x"b9",  x"6d",  x"17",  x"59",  x"d8",  x"58", -- 0518
         x"99",  x"71",  x"30",  x"1d",  x"a5",  x"07",  x"cd",  x"59", -- 0520
         x"ff",  x"cd",  x"51",  x"bd",  x"d6",  x"03",  x"c0",  x"3a", -- 0528
         x"61",  x"30",  x"be",  x"e1",  x"74",  x"28",  x"09",  x"fe", -- 0530
         x"ff",  x"06",  x"28",  x"05",  x"f1",  x"3e",  x"0b",  x"90", -- 0538
         x"19",  x"04",  x"0c",  x"d8",  x"4c",  x"15",  x"3c",  x"c7", -- 0540
         x"05",  x"20",  x"01",  x"3c",  x"5b",  x"7c",  x"ba",  x"8d", -- 0548
         x"c8",  x"21",  x"e6",  x"2d",  x"3a",  x"86",  x"bc",  x"e1", -- 0550
         x"26",  x"d0",  x"11",  x"e4",  x"14",  x"d7",  x"26",  x"88", -- 0558
         x"f5",  x"fc",  x"d8",  x"66",  x"21",  x"43",  x"4f",  x"30", -- 0560
         x"22",  x"64",  x"0e",  x"4d",  x"32",  x"66",  x"00",  x"37", -- 0568
         x"18",  x"16",  x"c0",  x"37",  x"2e",  x"e1",  x"ba",  x"ef", -- 0570
         x"26",  x"2e",  x"bc",  x"61",  x"b8",  x"d8",  x"11",  x"d6", -- 0578
         x"19",  x"26",  x"d2",  x"aa",  x"d2",  x"ce",  x"7e",  x"85", -- 0580
         x"40",  x"30",  x"09",  x"b7",  x"37",  x"c8",  x"cd",  x"70", -- 0588
         x"a3",  x"b9",  x"18",  x"c1",  x"99",  x"6d",  x"63",  x"a6", -- 0590
         x"42",  x"f5",  x"30",  x"5b",  x"05",  x"10",  x"af",  x"c9", -- 0598
         x"09",  x"1b",  x"c3",  x"d9",  x"03",  x"47",  x"7e",  x"f5", -- 05A0
         x"45",  x"13",  x"28",  x"a6",  x"11",  x"48",  x"fc",  x"da", -- 05A8
         x"d7",  x"e5",  x"80",  x"2a",  x"b1",  x"26",  x"d0",  x"b5", -- 05B0
         x"a0",  x"80",  x"dd",  x"41",  x"99",  x"28",  x"1f",  x"c7", -- 05B8
         x"7f",  x"a1",  x"93",  x"c0",  x"0e",  x"a9",  x"95",  x"31", -- 05C0
         x"f2",  x"b9",  x"87",  x"13",  x"1a",  x"b3",  x"38",  x"1e", -- 05C8
         x"d8",  x"60",  x"e5",  x"32",  x"47",  x"0e",  x"00",  x"eb", -- 05D0
         x"3e",  x"30",  x"1f",  x"be",  x"4e",  x"ed",  x"a0",  x"03", -- 05D8
         x"03",  x"18",  x"2b",  x"23",  x"10",  x"74",  x"71",  x"eb", -- 05E0
         x"79",  x"60",  x"b7",  x"ff",  x"c0",  x"c0",  x"cc",  x"3e", -- 05E8
         x"07",  x"a5",  x"03",  x"02",  x"36",  x"03",  x"01",  x"03", -- 05F0
         x"d0",  x"e2",  x"18",  x"82",  x"50",  x"d0",  x"50",  x"88", -- 05F8
         x"32",  x"f5",  x"9c",  x"61",  x"15",  x"81",  x"80",  x"74", -- 0600
         x"f1",  x"11",  x"5b",  x"fc",  x"d6",  x"05",  x"30",  x"78", -- 0608
         x"0c",  x"5f",  x"6f",  x"f1",  x"c6",  x"35",  x"a3",  x"9f", -- 0610
         x"00",  x"18",  x"4d",  x"d6",  x"02",  x"d8",  x"f5",  x"11", -- 0618
         x"56",  x"4f",  x"fc",  x"cc",  x"36",  x"df",  x"40",  x"20", -- 0620
         x"04",  x"06",  x"08",  x"18",  x"6a",  x"03",  x"e3",  x"0f", -- 0628
         x"00",  x"21",  x"cc",  x"fb",  x"11",  x"09",  x"00",  x"cb", -- 0630
         x"38",  x"00",  x"04",  x"19",  x"10",  x"fd",  x"eb",  x"18", -- 0638
         x"1f",  x"11",  x"0c",  x"62",  x"fc",  x"3d",  x"28",  x"b2", -- 0640
         x"d4",  x"73",  x"05",  x"13",  x"28",  x"11",  x"81",  x"05", -- 0648
         x"0d",  x"11",  x"50",  x"92",  x"05",  x"07",  x"11",  x"9d", -- 0650
         x"a2",  x"05",  x"01",  x"1b",  x"aa",  x"42",  x"63",  x"90", -- 0658
         x"d9",  x"f3",  x"31",  x"30",  x"00",  x"02",  x"a3",  x"a2", -- 0660
         x"91",  x"06",  x"5d",  x"54",  x"13",  x"06",  x"01",  x"dc", -- 0668
         x"78",  x"91",  x"00",  x"ed",  x"47",  x"3c",  x"d3",  x"8a", -- 0670
         x"3e",  x"cf",  x"d9",  x"03",  x"af",  x"02",  x"d3",  x"88", -- 0678
         x"4c",  x"f5",  x"06",  x"03",  x"40",  x"7e",  x"2f",  x"77", -- 0680
         x"56",  x"ba",  x"03",  x"c0",  x"dd",  x"28",  x"06",  x"1a", -- 0688
         x"0d",  x"2b",  x"22",  x"2b",  x"23",  x"80",  x"e5",  x"10", -- 0690
         x"ea",  x"0d",  x"21",  x"14",  x"f3",  x"22",  x"f1",  x"41", -- 0698
         x"cd",  x"e0",  x"f6",  x"11",  x"30",  x"61",  x"92",  x"7b", -- 06A0
         x"49",  x"9f",  x"f1",  x"ab",  x"9f",  x"e3",  x"d7",  x"0e", -- 06A8
         x"21",  x"f9",  x"85",  x"22",  x"01",  x"00",  x"31",  x"eb", -- 06B0
         x"e6",  x"fc",  x"b0",  x"f9",  x"cd",  x"12",  x"f7",  x"2e", -- 06B8
         x"11",  x"f7",  x"81",  x"cc",  x"21",  x"23",  x"dd",  x"5e", -- 06C0
         x"82",  x"30",  x"84",  x"55",  x"ac",  x"6e",  x"c2",  x"d2", -- 06C8
         x"d4",  x"e9",  x"fc",  x"c0",  x"11",  x"ca",  x"ef",  x"01", -- 06D0
         x"1f",  x"1b",  x"00",  x"36",  x"ff",  x"78",  x"11",  x"3d", -- 06D8
         x"06",  x"21",  x"b0",  x"fc",  x"0e",  x"0c",  x"09",  x"21", -- 06E0
         x"01",  x"24",  x"fc",  x"22",  x"eb",  x"ef",  x"22",  x"ed", -- 06E8
         x"b5",  x"02",  x"ef",  x"8f",  x"06",  x"b4",  x"f7",  x"22", -- 06F0
         x"cd",  x"ef",  x"92",  x"2f",  x"27",  x"55",  x"96",  x"4c", -- 06F8
         x"a9",  x"6a",  x"a3",  x"b7",  x"df",  x"d8",  x"1d",  x"e9", -- 0700
         x"17",  x"f1",  x"f8",  x"22",  x"60",  x"cb",  x"20",  x"e3", -- 0708
         x"ef",  x"ed",  x"5e",  x"11",  x"dc",  x"b8",  x"1b",  x"7b", -- 0710
         x"6d",  x"b2",  x"96",  x"42",  x"b6",  x"3d",  x"00",  x"e9", -- 0718
         x"2e",  x"07",  x"18",  x"07",  x"2e",  x"05",  x"59",  x"30", -- 0720
         x"50",  x"2c",  x"00",  x"7d",  x"cd",  x"58",  x"f7",  x"6c", -- 0728
         x"d8",  x"bf",  x"c8",  x"db",  x"dd",  x"ff",  x"a5",  x"d0", -- 0730
         x"28",  x"9a",  x"fe",  x"04",  x"c8",  x"1c",  x"ed",  x"53", -- 0738
         x"bc",  x"87",  x"67",  x"bc",  x"81",  x"b4",  x"c5",  x"d5", -- 0740
         x"25",  x"f4",  x"19",  x"04",  x"c1",  x"af",  x"ee",  x"ee", -- 0748
         x"21",  x"15",  x"6f",  x"f7",  x"e3",  x"e2",  x"40",  x"e9", -- 0750
         x"c1",  x"4f",  x"38",  x"f0",  x"aa",  x"de",  x"d8",  x"e7", -- 0758
         x"d0",  x"79",  x"b2",  x"8a",  x"f6",  x"28",  x"8a",  x"66", -- 0760
         x"d5",  x"b9",  x"10",  x"73",  x"20",  x"f9",  x"bf",  x"59", -- 0768
         x"ee",  x"7a",  x"04",  x"9b",  x"15",  x"c5",  x"0a",  x"53", -- 0770
         x"e1",  x"4d",  x"d8",  x"10",  x"d7",  x"f4",  x"0d",  x"0c", -- 0778
         x"06",  x"06",  x"18",  x"b6",  x"4d",  x"18",  x"f8",  x"f8", -- 0780
         x"28",  x"f6",  x"28",  x"18",  x"ac",  x"0f",  x"04",  x"18", -- 0788
         x"74",  x"a6",  x"e1",  x"28",  x"64",  x"f0",  x"cc",  x"20", -- 0790
         x"1e",  x"e4",  x"cd",  x"aa",  x"7c",  x"9f",  x"60",  x"18", -- 0798
         x"dc",  x"cd",  x"8f",  x"fe",  x"dc",  x"f3",  x"13",  x"00", -- 07A0
         x"b8",  x"aa",  x"14",  x"c3",  x"e9",  x"fa",  x"91",  x"34", -- 07A8
         x"5a",  x"4f",  x"ff",  x"5f",  x"07",  x"5f",  x"13",  x"51", -- 07B0
         x"1b",  x"05",  x"69",  x"60",  x"68",  x"fb",  x"01",  x"12", -- 07B8
         x"38",  x"01",  x"3d",  x"69",  x"74",  x"0e",  x"4f",  x"0c", -- 07C0
         x"c2",  x"3a",  x"1d",  x"b7",  x"29",  x"2a",  x"d1",  x"64", -- 07C8
         x"4c",  x"45",  x"91",  x"e6",  x"95",  x"0e",  x"68",  x"61", -- 07D0
         x"e7",  x"7a",  x"18",  x"1a",  x"8f",  x"a3",  x"6a",  x"00", -- 07D8
         x"cd",  x"36",  x"f8",  x"d8",  x"01",  x"02",  x"00",  x"1a", -- 07E0
         x"18",  x"13",  x"d6",  x"30",  x"e3",  x"00",  x"0a",  x"3f", -- 07E8
         x"d8",  x"80",  x"0d",  x"c8",  x"87",  x"01",  x"47",  x"87", -- 07F0
         x"87",  x"80",  x"47",  x"18",  x"ec",  x"98",  x"f7",  x"13", -- 07F8
         x"be",  x"c8",  x"c0",  x"e2",  x"4e",  x"38",  x"0a",  x"13", -- 0800
         x"77",  x"91",  x"09",  x"d5",  x"2e",  x"cc",  x"40",  x"b8", -- 0808
         x"c1",  x"eb",  x"36",  x"30",  x"eb",  x"a3",  x"a4",  x"75", -- 0810
         x"f0",  x"84",  x"d7",  x"bb",  x"e6",  x"43",  x"30",  x"20", -- 0818
         x"0a",  x"db",  x"9d",  x"86",  x"80",  x"1b",  x"79",  x"12", -- 0820
         x"f1",  x"18",  x"d1",  x"e4",  x"9a",  x"c9",  x"d6",  x"19", -- 0828
         x"14",  x"38",  x"15",  x"d9",  x"00",  x"06",  x"f8",  x"7b", -- 0830
         x"a0",  x"b1",  x"c9",  x"7b",  x"09",  x"06",  x"8f",  x"cb", -- 0838
         x"21",  x"7c",  x"01",  x"c8",  x"01",  x"db",  x"88",  x"06", -- 0840
         x"c7",  x"cd",  x"79",  x"f8",  x"9e",  x"85",  x"27",  x"0e", -- 0848
         x"64",  x"3a",  x"82",  x"5f",  x"f3",  x"b9",  x"8c",  x"61", -- 0850
         x"cd",  x"68",  x"f8",  x"44",  x"8d",  x"af",  x"1a",  x"77", -- 0858
         x"c9",  x"79",  x"9d",  x"18",  x"28",  x"39",  x"53",  x"05", -- 0860
         x"7b",  x"ee",  x"1b",  x"80",  x"18",  x"ed",  x"07",  x"1d", -- 0868
         x"d0",  x"37",  x"c4",  x"ad",  x"81",  x"0d",  x"ff",  x"01", -- 0870
         x"30",  x"93",  x"e1",  x"31",  x"cf",  x"21",  x"a1",  x"ea", -- 0878
         x"b8",  x"88",  x"97",  x"03",  x"d3",  x"80",  x"ff",  x"42", -- 0880
         x"1e",  x"3f",  x"62",  x"71",  x"0a",  x"e8",  x"de",  x"c9", -- 0888
         x"c5",  x"39",  x"36",  x"d6",  x"03",  x"ce",  x"a6",  x"2d", -- 0890
         x"02",  x"34",  x"79",  x"77",  x"86",  x"02",  x"0a",  x"cd", -- 0898
         x"7d",  x"f9",  x"3a",  x"16",  x"84",  x"ca",  x"18",  x"c3", -- 08A0
         x"6e",  x"7b",  x"d4",  x"fa",  x"2a",  x"18",  x"a7",  x"f5", -- 08A8
         x"5e",  x"3c",  x"8d",  x"e7",  x"a7",  x"c0",  x"eb",  x"22", -- 08B0
         x"3b",  x"00",  x"0f",  x"26",  x"29",  x"22",  x"3d",  x"04", -- 08B8
         x"b1",  x"3a",  x"b4",  x"36",  x"25",  x"02",  x"13",  x"fc", -- 08C0
         x"02",  x"29",  x"4c",  x"e6",  x"38",  x"e9",  x"4c",  x"f1", -- 08C8
         x"f3",  x"40",  x"04",  x"3a",  x"14",  x"6f",  x"c9",  x"06", -- 08D0
         x"21",  x"06",  x"3f",  x"f6",  x"dc",  x"97",  x"b4",  x"07", -- 08D8
         x"67",  x"32",  x"23",  x"32",  x"14",  x"94",  x"1b",  x"0e", -- 08E0
         x"0a",  x"a9",  x"f0",  x"39",  x"30",  x"e6",  x"d6",  x"36", -- 08E8
         x"31",  x"38",  x"de",  x"63",  x"f1",  x"23",  x"ca",  x"8d", -- 08F0
         x"f8",  x"e0",  x"4d",  x"05",  x"33",  x"8d",  x"34",  x"ca", -- 08F8
         x"f3",  x"f9",  x"31",  x"08",  x"5b",  x"74",  x"f8",  x"bd", -- 0900
         x"2b",  x"3c",  x"7f",  x"18",  x"4a",  x"a1",  x"3d",  x"67", -- 0908
         x"c0",  x"6d",  x"ec",  x"eb",  x"8b",  x"1b",  x"93",  x"92", -- 0910
         x"28",  x"00",  x"68",  x"9e",  x"19",  x"2c",  x"67",  x"db", -- 0918
         x"0e",  x"53",  x"1f",  x"21",  x"2c",  x"df",  x"af",  x"34", -- 0920
         x"c0",  x"e5",  x"08",  x"d8",  x"36",  x"28",  x"4e",  x"28", -- 0928
         x"30",  x"02",  x"3b",  x"d4",  x"02",  x"53",  x"c7",  x"b8", -- 0930
         x"02",  x"1e",  x"fe",  x"13",  x"28",  x"d8",  x"71",  x"8f", -- 0938
         x"43",  x"12",  x"18",  x"1a",  x"3a",  x"a7",  x"0e",  x"88", -- 0940
         x"1f",  x"2c",  x"e8",  x"83",  x"3a",  x"3c",  x"00",  x"90", -- 0948
         x"47",  x"9d",  x"30",  x"4f",  x"fa",  x"c1",  x"10",  x"c3", -- 0950
         x"d2",  x"b6",  x"05",  x"32",  x"6c",  x"3f",  x"02",  x"11", -- 0958
         x"9c",  x"dd",  x"34",  x"8a",  x"81",  x"c0",  x"1b",  x"1a", -- 0960
         x"3c",  x"77",  x"21",  x"a8",  x"23",  x"34",  x"23",  x"3d", -- 0968
         x"be",  x"0b",  x"d0",  x"77",  x"18",  x"77",  x"1a",  x"d5", -- 0970
         x"23",  x"35",  x"1a",  x"ba",  x"a8",  x"3d",  x"d4",  x"1a", -- 0978
         x"35",  x"46",  x"be",  x"63",  x"d8",  x"25",  x"18",  x"5d", -- 0980
         x"3a",  x"1a",  x"29",  x"4f",  x"3a",  x"4f",  x"21",  x"cd", -- 0988
         x"92",  x"05",  x"90",  x"33",  x"ca",  x"41",  x"b4",  x"7c", -- 0990
         x"04",  x"22",  x"2d",  x"d4",  x"cb",  x"c8",  x"ef",  x"31", -- 0998
         x"cb",  x"6f",  x"c3",  x"e5",  x"f2",  x"3f",  x"4b",  x"ad", -- 09A0
         x"5c",  x"cb",  x"e5",  x"c3",  x"ac",  x"0b",  x"78",  x"34", -- 09A8
         x"16",  x"85",  x"62",  x"df",  x"47",  x"06",  x"ae",  x"e6", -- 09B0
         x"f0",  x"78",  x"cc",  x"c0",  x"2f",  x"77",  x"a2",  x"53", -- 09B8
         x"2a",  x"e3",  x"29",  x"9f",  x"ae",  x"28",  x"77",  x"27", -- 09C0
         x"b9",  x"fc",  x"3a",  x"95",  x"27",  x"77",  x"eb",  x"be", -- 09C8
         x"a4",  x"af",  x"f5",  x"b6",  x"56",  x"b4",  x"0b",  x"4f", -- 09D0
         x"8d",  x"02",  x"47",  x"f1",  x"a8",  x"ab",  x"01",  x"41", -- 09D8
         x"a0",  x"66",  x"c1",  x"f5",  x"78",  x"91",  x"3f",  x"28", -- 09E0
         x"37",  x"0f",  x"2e",  x"9d",  x"21",  x"19",  x"18",  x"02", -- 09E8
         x"55",  x"f2",  x"cb",  x"ad",  x"c5",  x"c8",  x"0c",  x"27", -- 09F0
         x"47",  x"2b",  x"54",  x"1b",  x"f8",  x"3c",  x"fc",  x"2e", -- 09F8
         x"cb",  x"0a",  x"91",  x"4f",  x"b4",  x"3f",  x"f9",  x"bc", -- 0A00
         x"53",  x"9f",  x"54",  x"42",  x"02",  x"c1",  x"db",  x"a9", -- 0A08
         x"db",  x"fa",  x"4d",  x"16",  x"10",  x"ca",  x"f1",  x"28", -- 0A10
         x"4f",  x"50",  x"47",  x"a8",  x"66",  x"ee",  x"2b",  x"90", -- 0A18
         x"28",  x"0d",  x"36",  x"0e",  x"20",  x"c5",  x"f5",  x"c4", -- 0A20
         x"2d",  x"82",  x"80",  x"b0",  x"7e",  x"a3",  x"0f",  x"cb", -- 0A28
         x"bf",  x"77",  x"f1",  x"8b",  x"e9",  x"8c",  x"33",  x"33", -- 0A30
         x"c9",  x"0e",  x"0d",  x"0c",  x"27",  x"cb",  x"19",  x"07", -- 0A38
         x"00",  x"e6",  x"7f",  x"cc",  x"ee",  x"f3",  x"f5",  x"cc", -- 0A40
         x"53",  x"fa",  x"f1",  x"04",  x"15",  x"fb",  x"0d",  x"3e", -- 0A48
         x"83",  x"d3",  x"93",  x"f1",  x"c2",  x"90",  x"f1",  x"fb", -- 0A50
         x"c9",  x"cc",  x"b6",  x"d3",  x"82",  x"b7",  x"ff",  x"01", -- 0A58
         x"80",  x"3e",  x"c7",  x"d3",  x"83",  x"3e",  x"40",  x"4c", -- 0A60
         x"03",  x"27",  x"10",  x"3e",  x"96",  x"af",  x"03",  x"cf", -- 0A68
         x"aa",  x"99",  x"1b",  x"92",  x"19",  x"92",  x"b8",  x"6e", -- 0A70
         x"2e",  x"b5",  x"0a",  x"03",  x"ff",  x"2c",  x"03",  x"17", -- 0A78
         x"3a",  x"93",  x"3d",  x"c0",  x"3d",  x"c9",  x"18",  x"1e", -- 0A80
         x"1f",  x"5d",  x"00",  x"03",  x"08",  x"09",  x"0a",  x"0b", -- 0A88
         x"02",  x"0d",  x"b9",  x"e6",  x"19",  x"de",  x"29",  x"5e", -- 0A90
         x"14",  x"0c",  x"1b",  x"0c",  x"00",  x"a3",  x"9a",  x"00", -- 0A98
         x"1c",  x"1d",  x"7d",  x"ab",  x"8d",  x"82",  x"85",  x"86", -- 0AA0
         x"00",  x"84",  x"cf",  x"c3",  x"96",  x"90",  x"9b",  x"9c", -- 0AA8
         x"af",  x"00",  x"c4",  x"95",  x"92",  x"ae",  x"87",  x"ac", -- 0AB0
         x"8c",  x"91",  x"03",  x"83",  x"ad",  x"80",  x"81",  x"c2", -- 0AB8
         x"00",  x"00",  x"60",  x"93",  x"02",  x"ec",  x"ed",  x"ee", -- 0AC0
         x"ef",  x"f0",  x"0f",  x"ca",  x"cc",  x"d0",  x"d1",  x"ce", -- 0AC8
         x"c0",  x"fc",  x"df",  x"fd",  x"db",  x"b3",  x"a0",  x"00", -- 0AD0
         x"a1",  x"9e",  x"9f",  x"c0",  x"c7",  x"b4",  x"b0",  x"b1", -- 0AD8
         x"d8",  x"c7",  x"dc",  x"ff",  x"00",  x"dd",  x"be",  x"b2", -- 0AE0
         x"a3",  x"f9",  x"aa",  x"a5",  x"a9",  x"00",  x"88",  x"c8", -- 0AE8
         x"c6",  x"bc",  x"b6",  x"bb",  x"ba",  x"fb",  x"00",  x"fa", -- 0AF0
         x"bd",  x"b8",  x"a8",  x"c1",  x"a6",  x"89",  x"b5",  x"00", -- 0AF8
         x"f8",  x"a4",  x"a2",  x"a7",  x"c5",  x"98",  x"00",  x"d7", -- 0B00
         x"00",  x"b9",  x"d2",  x"d3",  x"f2",  x"e0",  x"e2",  x"f4", -- 0B08
         x"e8",  x"01",  x"f5",  x"f6",  x"8a",  x"d4",  x"8b",  x"d8", -- 0B10
         x"d9",  x"b8",  x"e3",  x"d5",  x"d6",  x"ea",  x"00",  x"e7", -- 0B18
         x"f3",  x"e6",  x"c9",  x"e1",  x"e9",  x"e3",  x"e4",  x"03", -- 0B20
         x"cb",  x"94",  x"9d",  x"97",  x"9a",  x"99",  x"b9",  x"8f", -- 0B28
         x"97",  x"06",  x"4e",  x"53",  x"54",  x"8d",  x"1c",  x"e0", -- 0B30
         x"01",  x"52",  x"45",  x"41",  x"44",  x"45",  x"52",  x"98", -- 0B38
         x"f4",  x"ef",  x"50",  x"55",  x"1f",  x"4e",  x"43",  x"48", -- 0B40
         x"11",  x"ec",  x"05",  x"4c",  x"49",  x"7b",  x"19",  x"08", -- 0B48
         x"9c",  x"1b",  x"4f",  x"53",  x"03",  x"00",  x"d6",  x"80", -- 0B50
         x"c3",  x"ba",  x"f0",  x"41",  x"1d",  x"53",  x"47",  x"4e", -- 0B58
         x"12",  x"00",  x"14",  x"c3",  x"81",  x"f1",  x"54",  x"49", -- 0B60
         x"4d",  x"45",  x"94",  x"0b",  x"22",  x"f5",  x"1d",  x"43", -- 0B68
         x"4c",  x"4f",  x"3d",  x"e4",  x"0b",  x"8e",  x"43",  x"39", -- 0B70
         x"52",  x"54",  x"ba",  x"18",  x"00",  x"42",  x"41",  x"05", -- 0B78
         x"14",  x"01",  x"0c",  x"06",  x"72",  x"6f",  x"62",  x"6f", -- 0B80
         x"74",  x"04",  x"6e",  x"cd",  x"19",  x"5a",  x"20",  x"83", -- 0B88
         x"4d",  x"30",  x"31",  x"47",  x"14",  x"80",  x"1b",  x"0a", -- 0B90
         x"73",  x"74",  x"61",  x"72",  x"74",  x"20",  x"ca",  x"04", -- 0B98
         x"70",  x"65",  x"57",  x"31",  x"07",  x"42",  x"5e",  x"2d", -- 0BA0
         x"65",  x"72",  x"81",  x"24",  x"72",  x"07",  x"00",  x"6d", -- 0BA8
         x"65",  x"6d",  x"8c",  x"06",  x"79",  x"20",  x"70",  x"0c", -- 0BB0
         x"74",  x"65",  x"7e",  x"63",  x"02",  x"96",  x"80",  x"65", -- 0BB8
         x"6e",  x"64",  x"20",  x"6f",  x"66",  x"20",  x"94",  x"17", -- 0BC0
         x"00",  x"72",  x"fd",  x"14",  x"06",  x"10",  x"6e",  x"86", -- 0BC8
         x"1d",  x"20",  x"66",  x"6f",  x"75",  x"1a",  x"00",  x"39", -- 0BD0
         x"62",  x"61",  x"0d",  x"41",  x"14",  x"00",  x"66",  x"69", -- 0BD8
         x"6c",  x"65",  x"14",  x"19",  x"20",  x"06",  x"2c",  x"2e", -- 0BE0
         x"3a",  x"43",  x"ff",  x"bf",  x"20",  x"fb",  x"fc",  x"c2", -- 0BE8
         x"fc",  x"e4",  x"16",  x"fc",  x"bd",  x"ff",  x"f7",  x"79", -- 0BF0
         x"f2",  x"b3",  x"fb",  x"c4",  x"cf",  x"f3",  x"a4",  x"0e", -- 0BF8
         x"9e",  x"40",  x"3e",  x"3c",  x"2b",  x"34",  x"be",  x"20", -- 0C00
         x"cf",  x"96",  x"ad",  x"31",  x"f7",  x"3e",  x"18",  x"6f", -- 0C08
         x"0a",  x"02",  x"0a",  x"91",  x"30",  x"e1",  x"ed",  x"4d", -- 0C10
         x"f5",  x"f9",  x"fd",  x"32",  x"b0",  x"e1",  x"3e",  x"7f", -- 0C18
         x"32",  x"69",  x"24",  x"04",  x"a5",  x"4b",  x"e4",  x"82", -- 0C20
         x"3d",  x"16",  x"fb",  x"5f",  x"81",  x"bc",  x"16",  x"35", -- 0C28
         x"bb",  x"f4",  x"a5",  x"a6",  x"20",  x"dc",  x"82",  x"cd", -- 0C30
         x"30",  x"0d",  x"fd",  x"28",  x"1c",  x"be",  x"ad",  x"bf", -- 0C38
         x"df",  x"d8",  x"b4",  x"07",  x"36",  x"6d",  x"06",  x"97", -- 0C40
         x"bf",  x"0e",  x"0d",  x"d6",  x"a6",  x"fb",  x"e8",  x"df", -- 0C48
         x"28",  x"04",  x"d7",  x"87",  x"07",  x"5e",  x"e1",  x"34", -- 0C50
         x"fa",  x"c0",  x"c8",  x"e5",  x"d5",  x"c5",  x"21",  x"15", -- 0C58
         x"68",  x"fe",  x"e5",  x"f5",  x"2d",  x"7a",  x"0c",  x"7b", -- 0C60
         x"94",  x"02",  x"3a",  x"26",  x"9e",  x"e0",  x"06",  x"cb", -- 0C68
         x"c3",  x"cb",  x"fa",  x"37",  x"cb",  x"bd",  x"1b",  x"5a", -- 0C70
         x"97",  x"e0",  x"cd",  x"81",  x"fe",  x"67",  x"cd",  x"01", -- 0C78
         x"89",  x"fe",  x"6f",  x"d1",  x"c1",  x"c0",  x"c5",  x"e0", -- 0C80
         x"cf",  x"af",  x"cd",  x"83",  x"01",  x"fe",  x"f5",  x"84", -- 0C88
         x"67",  x"f1",  x"85",  x"bf",  x"7e",  x"13",  x"12",  x"e0", -- 0C90
         x"e0",  x"5f",  x"7d",  x"fe",  x"48",  x"28",  x"19",  x"6e", -- 0C98
         x"fe",  x"41",  x"34",  x"fe",  x"46",  x"80",  x"af",  x"3e", -- 0CA0
         x"a9",  x"d6",  x"00",  x"2c",  x"6f",  x"7c",  x"fe",  x"38", -- 0CA8
         x"c0",  x"7d",  x"c3",  x"00",  x"38",  x"fe",  x"fe",  x"40", -- 0CB0
         x"28",  x"6b",  x"d0",  x"d6",  x"00",  x"39",  x"d8",  x"84", -- 0CB8
         x"cb",  x"78",  x"28",  x"2d",  x"01",  x"71",  x"90",  x"9b", -- 0CC0
         x"f3",  x"d4",  x"61",  x"ae",  x"c0",  x"60",  x"0d",  x"ed", -- 0CC8
         x"41",  x"00",  x"cb",  x"7c",  x"c8",  x"3c",  x"fe",  x"0c", -- 0CD0
         x"38",  x"64",  x"00",  x"28",  x"60",  x"fe",  x"0e",  x"38", -- 0CD8
         x"5e",  x"28",  x"5a",  x"00",  x"fe",  x"0f",  x"28",  x"58", -- 0CE0
         x"d6",  x"2b",  x"38",  x"4e",  x"00",  x"fe",  x"0d",  x"d0", -- 0CE8
         x"21",  x"33",  x"fb",  x"18",  x"55",  x"70",  x"3d",  x"fe", -- 0CF0
         x"d8",  x"01",  x"d6",  x"06",  x"c8",  x"30",  x"0d",  x"fe", -- 0CF8
         x"fa",  x"80",  x"f8",  x"d6",  x"1f",  x"cb",  x"1c",  x"73", -- 0D00
         x"c8",  x"d6",  x"b3",  x"e0",  x"50",  x"1b",  x"38",  x"34", -- 0D08
         x"fe",  x"1e",  x"1e",  x"c0",  x"18",  x"2f",  x"60",  x"3b", -- 0D10
         x"26",  x"28",  x"28",  x"26",  x"3b",  x"20",  x"28",  x"50", -- 0D18
         x"20",  x"37",  x"18",  x"21",  x"40",  x"c1",  x"34",  x"20", -- 0D20
         x"78",  x"a9",  x"ba",  x"c0",  x"a0",  x"ef",  x"a4",  x"7c", -- 0D28
         x"20",  x"00",  x"c2",  x"b7",  x"20",  x"a2",  x"3e",  x"5f", -- 0D30
         x"18",  x"08",  x"03",  x"c6",  x"20",  x"c6",  x"2b",  x"c6", -- 0D38
         x"10",  x"05",  x"c1",  x"3e",  x"28",  x"1d",  x"21",  x"53", -- 0D40
         x"fb",  x"d0",  x"e2",  x"4f",  x"09",  x"7e",  x"7d",  x"fe", -- 0D48
         x"6d",  x"ee",  x"83",  x"5d",  x"28",  x"ec",  x"b7",  x"e1", -- 0D50
         x"d3",  x"a9",  x"44",  x"c4",  x"0a",  x"18",  x"0c",  x"43", -- 0D58
         x"e1",  x"fe",  x"7e",  x"ba",  x"3a",  x"96",  x"d4",  x"b7", -- 0D60
         x"88",  x"af",  x"bc",  x"11",  x"b2",  x"47",  x"31",  x"fe", -- 0D68
         x"7d",  x"1e",  x"8d",  x"8a",  x"e6",  x"c5",  x"04",  x"18", -- 0D70
         x"1f",  x"ea",  x"c1",  x"d1",  x"21",  x"33",  x"80",  x"e0", -- 0D78
         x"60",  x"20",  x"03",  x"1d",  x"d6",  x"21",  x"3c",  x"d2", -- 0D80
         x"cc",  x"fa",  x"a4",  x"3e",  x"25",  x"a3",  x"ff",  x"74", -- 0D88
         x"34",  x"93",  x"40",  x"af",  x"18",  x"d7",  x"3e",  x"f7", -- 0D90
         x"fc",  x"dc",  x"81",  x"cb",  x"01",  x"3b",  x"d8",  x"10", -- 0D98
         x"fa",  x"c0",  x"81",  x"bf",  x"b0",  x"ab",  x"db",  x"91", -- 0DA0
         x"2f",  x"53",  x"57",  x"9c",  x"6a",  x"ef",  x"fb",  x"f1", -- 0DA8
         x"2c",  x"0b",  x"67",  x"3e",  x"fe",  x"6b",  x"06",  x"6f", -- 0DB0
         x"90",  x"6a",  x"85",  x"6f",  x"03",  x"07",  x"b6",  x"85", -- 0DB8
         x"00",  x"d3",  x"91",  x"db",  x"90",  x"2f",  x"5f",  x"3e", -- 0DC0
         x"80",  x"92",  x"07",  x"ab",  x"92",  x"be",  x"69",  x"75", -- 0DC8
         x"09",  x"fe",  x"a6",  x"e4",  x"af",  x"65",  x"46",  x"5f", -- 0DD0
         x"6d",  x"69",  x"0b",  x"0a",  x"43",  x"93",  x"57",  x"ad", -- 0DD8
         x"2d",  x"aa",  x"80",  x"e3",  x"fe",  x"cd",  x"29",  x"ff", -- 0DE0
         x"3a",  x"6b",  x"c7",  x"15",  x"18",  x"ff",  x"2a",  x"93", -- 0DE8
         x"a3",  x"06",  x"80",  x"7e",  x"08",  x"f5",  x"0e",  x"24", -- 0DF0
         x"86",  x"6e",  x"28",  x"d4",  x"f2",  x"a6",  x"0c",  x"7a", -- 0DF8
         x"b3",  x"66",  x"3e",  x"85",  x"8e",  x"fe",  x"4b",  x"03", -- 0E00
         x"fb",  x"0c",  x"57",  x"c9",  x"c5",  x"4f",  x"96",  x"03", -- 0E08
         x"cb",  x"09",  x"f5",  x"dc",  x"3b",  x"00",  x"f1",  x"d4", -- 0E10
         x"2d",  x"ff",  x"10",  x"f4",  x"c1",  x"1e",  x"c4",  x"cd", -- 0E18
         x"06",  x"1e",  x"70",  x"20",  x"b6",  x"1e",  x"0c",  x"40", -- 0E20
         x"7a",  x"cd",  x"38",  x"2c",  x"32",  x"6a",  x"e3",  x"e2", -- 0E28
         x"02",  x"c4",  x"b5",  x"fa",  x"53",  x"f2",  x"ef",  x"de", -- 0E30
         x"cc",  x"eb",  x"3a",  x"10",  x"04",  x"fb",  x"79",  x"05", -- 0E38
         x"a8",  x"34",  x"f3",  x"9b",  x"7e",  x"e1",  x"94",  x"3e", -- 0E40
         x"05",  x"1c",  x"b0",  x"a5",  x"03",  x"0f",  x"29",  x"0b", -- 0E48
         x"0a",  x"03",  x"e7",  x"e2",  x"03",  x"d7",  x"16",  x"00", -- 0E50
         x"cd",  x"d1",  x"ff",  x"38",  x"f9",  x"fe",  x"90",  x"38", -- 0E58
         x"1a",  x"f5",  x"10",  x"f5",  x"b9",  x"58",  x"ad",  x"28", -- 0E60
         x"4f",  x"37",  x"cd",  x"e0",  x"00",  x"ff",  x"fe",  x"52", -- 0E68
         x"30",  x"f1",  x"10",  x"ef",  x"cd",  x"05",  x"e8",  x"ff", -- 0E70
         x"d8",  x"32",  x"6b",  x"05",  x"a5",  x"05",  x"aa",  x"a2", -- 0E78
         x"0b",  x"77",  x"01",  x"a9",  x"f1",  x"6a",  x"0e",  x"47", -- 0E80
         x"0e",  x"19",  x"b8",  x"c8",  x"37",  x"79",  x"db",  x"80", -- 0E88
         x"a5",  x"7c",  x"07",  x"5f",  x"4c",  x"f1",  x"77",  x"af", -- 0E90
         x"98",  x"99",  x"3c",  x"b0",  x"44",  x"4f",  x"81",  x"0a", -- 0E98
         x"81",  x"c9",  x"16",  x"08",  x"af",  x"5f",  x"43",  x"73", -- 0EA0
         x"3f",  x"30",  x"04",  x"74",  x"03",  x"d8",  x"37",  x"cb", -- 0EA8
         x"1b",  x"15",  x"20",  x"49",  x"c8",  x"0e",  x"7b",  x"c9", -- 0EB0
         x"00",  x"04",  x"18",  x"00",  x"0b",  x"c3",  x"8c",  x"c0", -- 0EB8
         x"7f",  x"7f",  x"42",  x"41",  x"00",  x"53",  x"49",  x"43", -- 0EC0
         x"00",  x"21",  x"bd",  x"c0",  x"11",  x"00",  x"00",  x"03", -- 0EC8
         x"01",  x"67",  x"00",  x"ed",  x"b0",  x"eb",  x"00",  x"f9", -- 0ED0
         x"cd",  x"69",  x"c6",  x"32",  x"ab",  x"03",  x"32",  x"00", -- 0ED8
         x"00",  x"04",  x"21",  x"92",  x"c0",  x"cd",  x"c9",  x"d1", -- 0EE0
         x"2c",  x"21",  x"ae",  x"05",  x"cd",  x"ae",  x"00",  x"c5", -- 0EE8
         x"21",  x"62",  x"03",  x"cd",  x"86",  x"c9",  x"7a",  x"18", -- 0EF0
         x"d6",  x"06",  x"21",  x"2a",  x"2b",  x"30",  x"03",  x"00", -- 0EF8
         x"11",  x"ff",  x"bf",  x"23",  x"cd",  x"89",  x"c6",  x"28", -- 0F00
         x"00",  x"09",  x"7e",  x"47",  x"2f",  x"77",  x"be",  x"70", -- 0F08
         x"28",  x"30",  x"f2",  x"2b",  x"42",  x"ff",  x"22",  x"b0", -- 0F10
         x"03",  x"18",  x"19",  x"22",  x"56",  x"27",  x"41",  x"c6", -- 0F18
         x"2a",  x"c0",  x"05",  x"11",  x"ef",  x"fb",  x"19",  x"cd", -- 0F20
         x"29",  x"16",  x"d8",  x"21",  x"a0",  x"40",  x"2a",  x"00", -- 0F28
         x"04",  x"e0",  x"7e",  x"fe",  x"78",  x"20",  x"01",  x"3e", -- 0F30
         x"00",  x"af",  x"32",  x"fc",  x"03",  x"31",  x"67",  x"03", -- 0F38
         x"18",  x"64",  x"0a",  x"7c",  x"52",  x"45",  x"b4",  x"7e", -- 0F40
         x"71",  x"c3",  x"00",  x"88",  x"c3",  x"0c",  x"0a",  x"0d", -- 0F48
         x"48",  x"43",  x"2d",  x"93",  x"11",  x"09",  x"00",  x"00", -- 0F50
         x"20",  x"42",  x"59",  x"54",  x"45",  x"53",  x"20",  x"6a", -- 0F58
         x"46",  x"23",  x"45",  x"0d",  x"00",  x"4d",  x"45",  x"4d", -- 0F60
         x"4f",  x"52",  x"59",  x"20",  x"45",  x"00",  x"4e",  x"44", -- 0F68
         x"20",  x"3f",  x"20",  x"3a",  x"00",  x"c3",  x"02",  x"89", -- 0F70
         x"c0",  x"c3",  x"67",  x"c9",  x"00",  x"c0",  x"00",  x"d6", -- 0F78
         x"00",  x"6f",  x"7c",  x"de",  x"00",  x"31",  x"67",  x"78", -- 0F80
         x"03",  x"47",  x"3e",  x"00",  x"60",  x"12",  x"35",  x"4a", -- 0F88
         x"ca",  x"99",  x"39",  x"00",  x"1c",  x"76",  x"98",  x"22", -- 0F90
         x"95",  x"b3",  x"98",  x"0a",  x"00",  x"dd",  x"47",  x"98", -- 0F98
         x"53",  x"d1",  x"99",  x"99",  x"0a",  x"00",  x"1a",  x"9f", -- 0FA0
         x"98",  x"65",  x"bc",  x"cd",  x"98",  x"d6",  x"00",  x"77", -- 0FA8
         x"3e",  x"98",  x"52",  x"c7",  x"4f",  x"80",  x"0b",  x"0f", -- 0FB0
         x"ff",  x"1b",  x"00",  x"0a",  x"01",  x"2c",  x"f0",  x"49", -- 0FB8
         x"d7",  x"4e",  x"00",  x"00",  x"65",  x"0b",  x"04",  x"fe", -- 0FC0
         x"ff",  x"00",  x"43",  x"29",  x"01",  x"04",  x"0d",  x"c5", -- 0FC8
         x"b0",  x"6b",  x"c6",  x"73",  x"ce",  x"45",  x"58",  x"54", -- 0FD0
         x"00",  x"c4",  x"41",  x"54",  x"41",  x"c9",  x"4e",  x"50", -- 0FD8
         x"55",  x"c0",  x"08",  x"49",  x"4d",  x"d2",  x"45",  x"41", -- 0FE0
         x"44",  x"18",  x"cc",  x"45",  x"54",  x"43",  x"54",  x"4f", -- 0FE8
         x"d2",  x"0d",  x"55",  x"4e",  x"c9",  x"46",  x"0f",  x"53", -- 0FF0
         x"e1",  x"09",  x"a3",  x"8c",  x"0f",  x"53",  x"55",  x"42", -- 0FF8
         x"0b",  x"54",  x"55",  x"33",  x"52",  x"4e",  x"05",  x"4d", -- 1000
         x"d3",  x"12",  x"30",  x"50",  x"cf",  x"2e",  x"cf",  x"4e", -- 1008
         x"ce",  x"55",  x"06",  x"4c",  x"4c",  x"d7",  x"41",  x"49", -- 1010
         x"38",  x"45",  x"02",  x"46",  x"d0",  x"4f",  x"4b",  x"45", -- 1018
         x"c4",  x"98",  x"03",  x"c1",  x"17",  x"4f",  x"cc",  x"49", -- 1020
         x"60",  x"4e",  x"36",  x"c3",  x"4c",  x"53",  x"d7",  x"49", -- 1028
         x"00",  x"44",  x"54",  x"48",  x"c2",  x"59",  x"45",  x"a1", -- 1030
         x"c3",  x"66",  x"41",  x"27",  x"d0",  x"52",  x"15",  x"54", -- 1038
         x"3f",  x"c3",  x"4f",  x"03",  x"1d",  x"52",  x"f6",  x"1c", -- 1040
         x"67",  x"52",  x"04",  x"4f",  x"c1",  x"6c",  x"c3",  x"53", -- 1048
         x"41",  x"56",  x"45",  x"80",  x"85",  x"57",  x"d4",  x"41", -- 1050
         x"00",  x"42",  x"28",  x"d4",  x"4f",  x"c6",  x"4e",  x"d3", -- 1058
         x"50",  x"67",  x"43",  x"07",  x"48",  x"45",  x"5a",  x"86", -- 1060
         x"81",  x"66",  x"45",  x"01",  x"50",  x"ab",  x"ad",  x"aa", -- 1068
         x"af",  x"de",  x"c1",  x"80",  x"aa",  x"cf",  x"52",  x"be", -- 1070
         x"0c",  x"bd",  x"bc",  x"d3",  x"47",  x"91",  x"30",  x"3f", -- 1078
         x"c1",  x"42",  x"53",  x"d5",  x"18",  x"53",  x"52",  x"c6", -- 1080
         x"94",  x"50",  x"b3",  x"60",  x"75",  x"53",  x"d3",  x"51", -- 1088
         x"52",  x"d2",  x"c1",  x"1f",  x"cc",  x"4e",  x"c5",  x"58", -- 1090
         x"50",  x"fe",  x"5d",  x"0d",  x"64",  x"49",  x"4e",  x"0c", -- 1098
         x"c1",  x"54",  x"4e",  x"d0",  x"d7",  x"4a",  x"4b",  x"c4", -- 10A0
         x"03",  x"1e",  x"d0",  x"49",  x"cc",  x"4c",  x"49",  x"52", -- 10A8
         x"30",  x"24",  x"d6",  x"83",  x"07",  x"c1",  x"53",  x"43", -- 10B0
         x"c3",  x"48",  x"09",  x"80",  x"10",  x"46",  x"54",  x"24", -- 10B8
         x"d2",  x"49",  x"47",  x"48",  x"d8",  x"05",  x"cd",  x"a1", -- 10C0
         x"74",  x"0e",  x"85",  x"06",  x"d4",  x"52",  x"98",  x"14", -- 10C8
         x"03",  x"46",  x"18",  x"46",  x"c5",  x"44",  x"cd",  x"30", -- 10D0
         x"c5",  x"b9",  x"00",  x"45",  x"80",  x"1a",  x"c9",  x"de", -- 10D8
         x"c7",  x"dc",  x"cc",  x"00",  x"48",  x"ca",  x"ec",  x"cb", -- 10E0
         x"01",  x"cf",  x"1f",  x"cc",  x"00",  x"5d",  x"ca",  x"07", -- 10E8
         x"ca",  x"eb",  x"c9",  x"cf",  x"ca",  x"03",  x"df",  x"c8", -- 10F0
         x"f6",  x"c9",  x"25",  x"ca",  x"81",  x"20",  x"18",  x"c9", -- 10F8
         x"ec",  x"d3",  x"00",  x"b3",  x"ca",  x"c0",  x"cb",  x"f7", -- 1100
         x"d3",  x"c4",  x"d0",  x"30",  x"37",  x"d4",  x"3a",  x"fa", -- 1108
         x"c5",  x"ea",  x"c6",  x"03",  x"d0",  x"dd",  x"b9",  x"cb", -- 1110
         x"f4",  x"df",  x"1b",  x"00",  x"38",  x"db",  x"fa",  x"ca", -- 1118
         x"48",  x"c9",  x"f2",  x"c6",  x"00",  x"aa",  x"c9",  x"43", -- 1120
         x"dc",  x"41",  x"dd",  x"40",  x"c6",  x"00",  x"2d",  x"c6", -- 1128
         x"b7",  x"c7",  x"b8",  x"c7",  x"e7",  x"c3",  x"c0",  x"19", -- 1130
         x"a6",  x"d6",  x"70",  x"d7",  x"bc",  x"d6",  x"00",  x"03", -- 1138
         x"03",  x"90",  x"d0",  x"e3",  x"d3",  x"bd",  x"d0",  x"00", -- 1140
         x"1f",  x"d9",  x"fd",  x"d9",  x"59",  x"d5",  x"6d",  x"d9", -- 1148
         x"00",  x"70",  x"da",  x"76",  x"da",  x"d7",  x"da",  x"ec", -- 1150
         x"da",  x"30",  x"31",  x"d4",  x"86",  x"00",  x"d5",  x"d6", -- 1158
         x"2c",  x"d3",  x"56",  x"d1",  x"bf",  x"d3",  x"00",  x"3b", -- 1160
         x"d3",  x"4b",  x"d3",  x"5b",  x"d3",  x"89",  x"d3",  x"00", -- 1168
         x"92",  x"d3",  x"79",  x"11",  x"d8",  x"79",  x"6a",  x"d4", -- 1170
         x"00",  x"7c",  x"98",  x"d5",  x"7c",  x"f3",  x"d5",  x"7f", -- 1178
         x"28",  x"00",  x"d9",  x"50",  x"5e",  x"ce",  x"46",  x"5d", -- 1180
         x"ce",  x"4e",  x"00",  x"46",  x"53",  x"4e",  x"52",  x"47", -- 1188
         x"4f",  x"44",  x"46",  x"06",  x"43",  x"4f",  x"56",  x"4f", -- 1190
         x"4d",  x"84",  x"58",  x"91",  x"85",  x"44",  x"44",  x"2f", -- 1198
         x"30",  x"0e",  x"ed",  x"c5",  x"6c",  x"53",  x"bc",  x"31", -- 11A0
         x"de",  x"0c",  x"43",  x"4e",  x"55",  x"46",  x"0a",  x"49", -- 11A8
         x"4f",  x"cd",  x"d0",  x"52",  x"81",  x"d4",  x"52",  x"07", -- 11B0
         x"9e",  x"ec",  x"95",  x"21",  x"20",  x"00",  x"46",  x"49", -- 11B8
         x"8e",  x"f4",  x"ef",  x"6c",  x"4f",  x"d5",  x"8c",  x"44", -- 11C0
         x"0d",  x"a7",  x"b3",  x"f2",  x"62",  x"42",  x"c0",  x"41", -- 11C8
         x"00",  x"4b",  x"00",  x"e5",  x"2a",  x"db",  x"03",  x"06", -- 11D0
         x"00",  x"00",  x"09",  x"09",  x"3e",  x"e5",  x"3e",  x"d0", -- 11D8
         x"95",  x"6f",  x"00",  x"3e",  x"ff",  x"9c",  x"38",  x"04", -- 11E0
         x"67",  x"39",  x"e1",  x"00",  x"d8",  x"1e",  x"0c",  x"18", -- 11E8
         x"14",  x"2a",  x"ca",  x"03",  x"00",  x"22",  x"58",  x"03", -- 11F0
         x"1e",  x"02",  x"01",  x"1e",  x"14",  x"db",  x"02",  x"00", -- 11F8
         x"02",  x"12",  x"02",  x"5a",  x"22",  x"bb",  x"b4",  x"43", -- 1200
         x"fe",  x"00",  x"55",  x"cb",  x"21",  x"dd",  x"c2",  x"57", -- 1208
         x"19",  x"44",  x"06",  x"4d",  x"0b",  x"3e",  x"3f",  x"1e", -- 1210
         x"0e",  x"d6",  x"d4",  x"c4",  x"05",  x"c3",  x"b5",  x"83", -- 1218
         x"d9",  x"2e",  x"11",  x"e2",  x"d2",  x"b4",  x"80",  x"ca", -- 1220
         x"0d",  x"c0",  x"7c",  x"a5",  x"3c",  x"c4",  x"04",  x"21", -- 1228
         x"d8",  x"3e",  x"c1",  x"af",  x"cb",  x"2f",  x"1d",  x"20", -- 1230
         x"00",  x"37",  x"dc",  x"fd",  x"dd",  x"cd",  x"df",  x"c6", -- 1238
         x"2b",  x"a0",  x"57",  x"21",  x"ea",  x"03",  x"3a",  x"00", -- 1240
         x"4d",  x"03",  x"b7",  x"28",  x"6b",  x"ed",  x"5b",  x"4e", -- 1248
         x"00",  x"03",  x"f2",  x"f0",  x"c3",  x"d5",  x"cd",  x"2a", -- 1250
         x"d8",  x"60",  x"d1",  x"04",  x"bb",  x"c4",  x"3e",  x"2a", -- 1258
         x"38",  x"1b",  x"02",  x"3e",  x"20",  x"8f",  x"29",  x"c6", -- 1260
         x"92",  x"87",  x"d1",  x"30",  x"06",  x"3f",  x"86",  x"25", -- 1268
         x"18",  x"ba",  x"2a",  x"50",  x"f7",  x"a0",  x"38",  x"f4", -- 1270
         x"d5",  x"11",  x"f9",  x"bc",  x"5d",  x"15",  x"ea",  x"22", -- 1278
         x"e9",  x"33",  x"ae",  x"80",  x"f5",  x"18",  x"47",  x"c8", -- 1280
         x"cd",  x"97",  x"f6",  x"28",  x"b5",  x"28",  x"c0",  x"c1", -- 1288
         x"39",  x"30",  x"58",  x"03",  x"d5",  x"7e",  x"23",  x"b6", -- 1290
         x"23",  x"28",  x"3e",  x"56",  x"7f",  x"34",  x"0a",  x"66", -- 1298
         x"56",  x"6f",  x"26",  x"94",  x"a0",  x"de",  x"d1",  x"c2", -- 12A0
         x"96",  x"c3",  x"01",  x"38",  x"b7",  x"3f",  x"18",  x"cd", -- 12A8
         x"3e",  x"3e",  x"2b",  x"56",  x"da",  x"0f",  x"30",  x"21", -- 12B0
         x"61",  x"19",  x"bd",  x"c8",  x"3c",  x"3d",  x"6a",  x"ca", -- 12B8
         x"0a",  x"f5",  x"3f",  x"c0",  x"78",  x"da",  x"c4",  x"47", -- 12C0
         x"d1",  x"f1",  x"d2",  x"0d",  x"8a",  x"c8",  x"d5",  x"c5", -- 12C8
         x"71",  x"cd",  x"6f",  x"1b",  x"b7",  x"17",  x"52",  x"00", -- 12D0
         x"38",  x"08",  x"f1",  x"f5",  x"b7",  x"20",  x"03",  x"c3", -- 12D8
         x"00",  x"20",  x"ca",  x"c5",  x"30",  x"11",  x"eb",  x"2a", -- 12E0
         x"d7",  x"05",  x"03",  x"1a",  x"02",  x"03",  x"13",  x"00", -- 12E8
         x"82",  x"20",  x"f7",  x"ed",  x"79",  x"43",  x"0c",  x"30", -- 12F0
         x"28",  x"22",  x"40",  x"13",  x"e3",  x"c1",  x"09",  x"e5", -- 12F8
         x"cd",  x"0c",  x"ab",  x"c4",  x"e1",  x"22",  x"0a",  x"eb", -- 1300
         x"36",  x"00",  x"ff",  x"d1",  x"23",  x"23",  x"73",  x"23", -- 1308
         x"72",  x"23",  x"31",  x"11",  x"62",  x"2b",  x"77",  x"23", -- 1310
         x"13",  x"ef",  x"3c",  x"ef",  x"a0",  x"d5",  x"23",  x"eb", -- 1318
         x"21",  x"c5",  x"67",  x"e5",  x"62",  x"6b",  x"01",  x"9e", -- 1320
         x"c8",  x"23",  x"98",  x"04",  x"a6",  x"3c",  x"05",  x"af", -- 1328
         x"be",  x"23",  x"14",  x"20",  x"fc",  x"eb",  x"29",  x"18", -- 1330
         x"07",  x"e8",  x"cd",  x"30",  x"c3",  x"c5",  x"43",  x"40", -- 1338
         x"55",  x"7e",  x"02",  x"c8",  x"0b",  x"2b",  x"06",  x"18", -- 1340
         x"f6",  x"2a",  x"5f",  x"03",  x"d9",  x"34",  x"2a",  x"2b", -- 1348
         x"d6",  x"25",  x"23",  x"c5",  x"14",  x"19",  x"60",  x"58", -- 1350
         x"69",  x"08",  x"3f",  x"c8",  x"3f",  x"18",  x"d0",  x"18", -- 1358
         x"e4",  x"9f",  x"05",  x"af",  x"03",  x"0e",  x"05",  x"6c", -- 1360
         x"5f",  x"08",  x"fb",  x"e5",  x"18",  x"fe",  x"9a",  x"00", -- 1368
         x"71",  x"c5",  x"47",  x"fe",  x"22",  x"ca",  x"91",  x"03", -- 1370
         x"c5",  x"b7",  x"ca",  x"97",  x"c5",  x"3a",  x"1b",  x"00", -- 1378
         x"b7",  x"7e",  x"20",  x"73",  x"fe",  x"3f",  x"3e",  x"9e", -- 1380
         x"36",  x"28",  x"6d",  x"1c",  x"30",  x"ce",  x"41",  x"fe", -- 1388
         x"3c",  x"38",  x"64",  x"88",  x"b8",  x"20",  x"c1",  x"c5", -- 1390
         x"03",  x"01",  x"6d",  x"c5",  x"c5",  x"06",  x"7f",  x"13", -- 1398
         x"07",  x"61",  x"38",  x"07",  x"fe",  x"7b",  x"df",  x"00", -- 13A0
         x"e6",  x"5f",  x"77",  x"4e",  x"eb",  x"c0",  x"64",  x"f2", -- 13A8
         x"26",  x"c5",  x"04",  x"7e",  x"e6",  x"0e",  x"7f",  x"20", -- 13B0
         x"15",  x"3a",  x"b6",  x"06",  x"a7",  x"c8",  x"3a",  x"51", -- 13B8
         x"a7",  x"28",  x"c0",  x"3c",  x"57",  x"2a",  x"0c",  x"50", -- 13C0
         x"e0",  x"15",  x"c8",  x"b9",  x"20",  x"00",  x"dd",  x"eb", -- 13C8
         x"e5",  x"13",  x"1a",  x"b7",  x"fa",  x"69",  x"01",  x"c5", -- 13D0
         x"4f",  x"78",  x"fe",  x"88",  x"20",  x"04",  x"42",  x"98", -- 13D8
         x"2b",  x"5b",  x"23",  x"43",  x"02",  x"3f",  x"00",  x"b9", -- 13E0
         x"28",  x"e5",  x"e1",  x"18",  x"bb",  x"48",  x"f1",  x"d4", -- 13E8
         x"98",  x"eb",  x"79",  x"60",  x"c1",  x"f6",  x"12",  x"06", -- 13F0
         x"13",  x"0c",  x"d6",  x"3a",  x"28",  x"6f",  x"49",  x"c6", -- 13F8
         x"af",  x"80",  x"a1",  x"d6",  x"54",  x"03",  x"28",  x"05", -- 1400
         x"d6",  x"0e",  x"c2",  x"e3",  x"d6",  x"16",  x"7e",  x"e4", -- 1408
         x"41",  x"09",  x"b8",  x"28",  x"e0",  x"85",  x"1f",  x"0c", -- 1410
         x"13",  x"18",  x"f3",  x"0f",  x"f7",  x"27",  x"45",  x"01", -- 1418
         x"c9",  x"4c",  x"39",  x"85",  x"00",  x"52",  x"a1",  x"8c", -- 1420
         x"00",  x"43",  x"4f",  x"92",  x"a5",  x"86",  x"10",  x"cd", -- 1428
         x"e3",  x"cd",  x"e4",  x"00",  x"dd",  x"e3",  x"fe",  x"1c", -- 1430
         x"11",  x"9f",  x"c5",  x"28",  x"07",  x"0e",  x"fe",  x"1d", -- 1438
         x"11",  x"a4",  x"06",  x"80",  x"a7",  x"1e",  x"11",  x"a8", -- 1440
         x"15",  x"c5",  x"20",  x"14",  x"34",  x"8e",  x"c9",  x"cd", -- 1448
         x"2c",  x"a7",  x"cb",  x"6e",  x"a3",  x"80",  x"f1",  x"c5", -- 1450
         x"e1",  x"c3",  x"5e",  x"cb",  x"00",  x"cd",  x"0f",  x"df", -- 1458
         x"20",  x"02",  x"e1",  x"c9",  x"cd",  x"18",  x"27",  x"df", -- 1460
         x"38",  x"e1",  x"87",  x"32",  x"df",  x"18",  x"c1",  x"66", -- 1468
         x"98",  x"8b",  x"d5",  x"dd",  x"23",  x"1c",  x"18",  x"f7", -- 1470
         x"11",  x"f7",  x"0a",  x"d5",  x"28",  x"17",  x"d4",  x"21", -- 1478
         x"eb",  x"e3",  x"28",  x"96",  x"b3",  x"9c",  x"8c",  x"c8", -- 1480
         x"e1",  x"f3",  x"bd",  x"28",  x"28",  x"06",  x"10",  x"c2", -- 1488
         x"48",  x"07",  x"c3",  x"eb",  x"7d",  x"b4",  x"ca",  x"d9", -- 1490
         x"2c",  x"22",  x"10",  x"cb",  x"ff",  x"a3",  x"a3",  x"51", -- 1498
         x"e1",  x"a0",  x"99",  x"c1",  x"c3",  x"9a",  x"03",  x"cd", -- 14A0
         x"5f",  x"de",  x"3a",  x"09",  x"91",  x"1c",  x"25",  x"f3", -- 14A8
         x"3e",  x"cc",  x"89",  x"b2",  x"dc",  x"05",  x"f1",  x"af", -- 14B0
         x"18",  x"ea",  x"c0",  x"16",  x"85",  x"e0",  x"26",  x"5e", -- 14B8
         x"03",  x"c3",  x"5d",  x"01",  x"15",  x"d8",  x"68",  x"0d", -- 14C0
         x"b5",  x"cf",  x"fa",  x"06",  x"ff",  x"3d",  x"22",  x"c4", -- 14C8
         x"17",  x"c3",  x"19",  x"c8",  x"f7",  x"6d",  x"09",  x"d9", -- 14D0
         x"02",  x"db",  x"d5",  x"3f",  x"89",  x"e0",  x"97",  x"b4", -- 14D8
         x"d8",  x"0a",  x"b2",  x"9a",  x"00",  x"1d",  x"de",  x"af", -- 14E0
         x"6f",  x"67",  x"22",  x"d5",  x"c1",  x"ff",  x"cc",  x"83", -- 14E8
         x"0e",  x"df",  x"03",  x"e5",  x"c5",  x"2a",  x"31",  x"3b", -- 14F0
         x"c9",  x"7c",  x"e5",  x"18",  x"7d",  x"93",  x"c9",  x"b2", -- 14F8
         x"80",  x"41",  x"d8",  x"fe",  x"5b",  x"3f",  x"c9",  x"3a", -- 1500
         x"f1",  x"51",  x"e5",  x"bb",  x"8f",  x"79",  x"6e",  x"74", -- 1508
         x"d6",  x"0a",  x"3e",  x"08",  x"18",  x"eb",  x"4d",  x"fb", -- 1510
         x"0c",  x"dd",  x"f5",  x"de",  x"72",  x"c8",  x"00",  x"38", -- 1518
         x"13",  x"3a",  x"41",  x"03",  x"47",  x"3a",  x"ac",  x"31", -- 1520
         x"03",  x"04",  x"ba",  x"06",  x"05",  x"b8",  x"cc",  x"61", -- 1528
         x"cb",  x"88",  x"5a",  x"0b",  x"79",  x"80",  x"d4",  x"c1", -- 1530
         x"f1",  x"6b",  x"c9",  x"e7",  x"a6",  x"b7",  x"2e",  x"09", -- 1538
         x"af",  x"04",  x"7b",  x"3c",  x"69",  x"4a",  x"fd",  x"b1", -- 1540
         x"d3",  x"22",  x"61",  x"8c",  x"64",  x"63",  x"03",  x"65", -- 1548
         x"82",  x"41",  x"6c",  x"c9",  x"ed",  x"53",  x"46",  x"da", -- 1550
         x"68",  x"89",  x"80",  x"25",  x"de",  x"cd",  x"c8",  x"dd", -- 1558
         x"28",  x"12",  x"90",  x"c5",  x"1d",  x"2a",  x"13",  x"ab", -- 1560
         x"a6",  x"ff",  x"b4",  x"cd",  x"08",  x"e1",  x"3a",  x"a3", -- 1568
         x"80",  x"c5",  x"cd",  x"91",  x"c7",  x"e1",  x"4e",  x"23", -- 1570
         x"00",  x"46",  x"23",  x"78",  x"b1",  x"28",  x"59",  x"cd", -- 1578
         x"67",  x"00",  x"c7",  x"cd",  x"f9",  x"c8",  x"c5",  x"5e", -- 1580
         x"23",  x"56",  x"29",  x"23",  x"e5",  x"8f",  x"9d",  x"cd", -- 1588
         x"71",  x"36",  x"84",  x"8f",  x"1f",  x"2c",  x"65",  x"9e", -- 1590
         x"ee",  x"d2",  x"66",  x"28",  x"14",  x"b9",  x"43",  x"d3", -- 1598
         x"f2",  x"3c",  x"23",  x"7b",  x"9a",  x"02",  x"11",  x"1a", -- 15A0
         x"cb",  x"40",  x"f2",  x"4e",  x"c7",  x"18",  x"49",  x"e6", -- 15A8
         x"1c",  x"a8",  x"18",  x"ba",  x"1f",  x"d7",  x"18",  x"6e", -- 15B0
         x"f2",  x"bf",  x"44",  x"63",  x"03",  x"d2",  x"8e",  x"9a", -- 15B8
         x"05",  x"e1",  x"55",  x"c0",  x"5a",  x"10",  x"c2",  x"fe", -- 15C0
         x"03",  x"20",  x"58",  x"ea",  x"84",  x"2f",  x"0c",  x"4e", -- 15C8
         x"ee",  x"66",  x"2a",  x"82",  x"15",  x"7f",  x"5d",  x"8b", -- 15D0
         x"f6",  x"29",  x"06",  x"26",  x"c9",  x"0d",  x"d6",  x"7f", -- 15D8
         x"fe",  x"56",  x"d7",  x"4c",  x"d6",  x"55",  x"96",  x"b3", -- 15E0
         x"e3",  x"6e",  x"18",  x"b0",  x"21",  x"2c",  x"c1",  x"47", -- 15E8
         x"5a",  x"ac",  x"c7",  x"33",  x"10",  x"f8",  x"f0",  x"56", -- 15F0
         x"c9",  x"be",  x"b0",  x"0a",  x"ca",  x"78",  x"21",  x"a0", -- 15F8
         x"39",  x"a0",  x"81",  x"2c",  x"81",  x"c0",  x"a9",  x"00", -- 1600
         x"e5",  x"69",  x"60",  x"7a",  x"b3",  x"eb",  x"cd",  x"d8", -- 1608
         x"eb",  x"42",  x"b0",  x"01",  x"e0",  x"b7",  x"e1",  x"c8", -- 1610
         x"05",  x"09",  x"18",  x"e3",  x"3e",  x"64",  x"0b",  x"e2", -- 1618
         x"cd",  x"95",  x"a6",  x"c1",  x"f8",  x"bd",  x"a2",  x"18", -- 1620
         x"22",  x"c8",  x"e5",  x"30",  x"02",  x"30",  x"cd",  x"c1", -- 1628
         x"c7",  x"d1",  x"cc",  x"ab",  x"09",  x"d5",  x"18",  x"2b", -- 1630
         x"56",  x"2b",  x"d1",  x"6e",  x"35",  x"2a",  x"15",  x"80", -- 1638
         x"30",  x"e1",  x"20",  x"e8",  x"d1",  x"f9",  x"eb",  x"33", -- 1640
         x"0e",  x"08",  x"a7",  x"5b",  x"c3",  x"11",  x"e3",  x"04", -- 1648
         x"7f",  x"58",  x"04",  x"b4",  x"00",  x"cd",  x"cd",  x"cc", -- 1650
         x"c8",  x"a6",  x"cd",  x"26",  x"60",  x"cd",  x"3e",  x"eb", -- 1658
         x"d6",  x"e1",  x"c5",  x"d5",  x"06",  x"01",  x"00",  x"81", -- 1660
         x"51",  x"5a",  x"a2",  x"40",  x"ab",  x"3e",  x"01",  x"20", -- 1668
         x"0e",  x"a4",  x"e1",  x"9b",  x"18",  x"d0",  x"1b",  x"1b", -- 1670
         x"36",  x"f5",  x"33",  x"33",  x"cf",  x"33",  x"06",  x"02", -- 1678
         x"81",  x"c5",  x"33",  x"cd",  x"16",  x"de",  x"86",  x"af", -- 1680
         x"8f",  x"86",  x"2a",  x"d0",  x"e8",  x"28",  x"b7",  x"a3", -- 1688
         x"ce",  x"a6",  x"9f",  x"65",  x"b6",  x"7f",  x"c9",  x"23", -- 1690
         x"0e",  x"c2",  x"83",  x"59",  x"59",  x"3a",  x"0a",  x"50", -- 1698
         x"d1",  x"0f",  x"e5",  x"ca",  x"3c",  x"65",  x"a7",  x"43", -- 16A0
         x"ca",  x"6e",  x"ef",  x"e1",  x"a3",  x"50",  x"11",  x"54", -- 16A8
         x"d7",  x"70",  x"c8",  x"d6",  x"80",  x"da",  x"c0",  x"b0", -- 16B0
         x"fe",  x"25",  x"00",  x"38",  x"14",  x"d6",  x"50",  x"38", -- 16B8
         x"34",  x"fe",  x"05",  x"16",  x"38",  x"0a",  x"47",  x"f2", -- 16C0
         x"a0",  x"28",  x"29",  x"c3",  x"03",  x"e0",  x"0e",  x"c6", -- 16C8
         x"25",  x"07",  x"4f",  x"85",  x"b7",  x"a4",  x"14",  x"40", -- 16D0
         x"c2",  x"09",  x"f1",  x"0d",  x"c5",  x"96",  x"a9",  x"60", -- 16D8
         x"d0",  x"99",  x"90",  x"28",  x"f7",  x"b3",  x"c0",  x"3f", -- 16E0
         x"a3",  x"8c",  x"bc",  x"db",  x"e3",  x"ac",  x"e8",  x"cb", -- 16E8
         x"ea",  x"63",  x"c3",  x"6f",  x"3e",  x"2c",  x"be",  x"9f", -- 16F0
         x"71",  x"3e",  x"29",  x"18",  x"85",  x"d2",  x"26",  x"90", -- 16F8
         x"a6",  x"aa",  x"eb",  x"d6",  x"25",  x"e5",  x"16",  x"d5", -- 1700
         x"9e",  x"e6",  x"d1",  x"d2",  x"87",  x"f9",  x"85",  x"38", -- 1708
         x"dd",  x"80",  x"cc",  x"86",  x"f3",  x"dd",  x"06",  x"c0", -- 1710
         x"fe",  x"13",  x"28",  x"08",  x"87",  x"4a",  x"c0",  x"8d", -- 1718
         x"22",  x"18",  x"0f",  x"c8",  x"92",  x"1e",  x"c8",  x"3c", -- 1720
         x"fe",  x"0a",  x"02",  x"30",  x"02",  x"18",  x"0a",  x"f1", -- 1728
         x"c0",  x"f6",  x"c0",  x"c0",  x"00",  x"21",  x"f6",  x"ff", -- 1730
         x"c1",  x"a1",  x"89",  x"0d",  x"f5",  x"7d",  x"a4",  x"3c", -- 1738
         x"9c",  x"8d",  x"22",  x"d3",  x"d7",  x"3a",  x"12",  x"b6", -- 1740
         x"49",  x"2b",  x"ab",  x"c3",  x"4a",  x"ae",  x"a0",  x"f1", -- 1748
         x"21",  x"21",  x"c3",  x"01",  x"c2",  x"71",  x"c3",  x"c3", -- 1750
         x"88",  x"c3",  x"2a",  x"8c",  x"16",  x"7c",  x"b5",  x"1e", -- 1758
         x"5c",  x"56",  x"c3",  x"d7",  x"72",  x"d3",  x"90",  x"7c", -- 1760
         x"61",  x"a3",  x"a1",  x"42",  x"9d",  x"f2",  x"07",  x"6f", -- 1768
         x"c9",  x"1e",  x"08",  x"c3",  x"19",  x"40",  x"0d",  x"3a", -- 1770
         x"e8",  x"03",  x"fe",  x"90",  x"01",  x"da",  x"45",  x"d7", -- 1778
         x"01",  x"80",  x"90",  x"11",  x"fe",  x"db",  x"93",  x"00", -- 1780
         x"18",  x"d7",  x"e1",  x"51",  x"c8",  x"15",  x"18",  x"e1", -- 1788
         x"2b",  x"0c",  x"40",  x"2e",  x"d0",  x"e5",  x"f5",  x"21", -- 1790
         x"98",  x"51",  x"19",  x"8e",  x"30",  x"da",  x"c2",  x"e4", -- 1798
         x"85",  x"19",  x"29",  x"c0",  x"01",  x"f1",  x"d6",  x"30", -- 17A0
         x"5f",  x"16",  x"00",  x"37",  x"19",  x"eb",  x"c0",  x"31", -- 17A8
         x"e0",  x"28",  x"ad",  x"62",  x"5e",  x"53",  x"be",  x"c8", -- 17B0
         x"e5",  x"94",  x"dc",  x"28",  x"10",  x"53",  x"e1",  x"b0", -- 17B8
         x"68",  x"bd",  x"6c",  x"ba",  x"10",  x"df",  x"16",  x"e3", -- 17C0
         x"af",  x"c0",  x"93",  x"5f",  x"7c",  x"9a",  x"57",  x"28", -- 17C8
         x"da",  x"3e",  x"be",  x"b5",  x"f1",  x"3c",  x"01",  x"28", -- 17D0
         x"aa",  x"a6",  x"45",  x"d2",  x"0d",  x"eb",  x"29",  x"22", -- 17D8
         x"56",  x"bd",  x"bd",  x"30",  x"8a",  x"dd",  x"53",  x"ed", -- 17E0
         x"f2",  x"e0",  x"cd",  x"cc",  x"05",  x"01",  x"54",  x"6f", -- 17E8
         x"10",  x"0e",  x"51",  x"03",  x"e8",  x"67",  x"94",  x"21", -- 17F0
         x"e5",  x"19",  x"3e",  x"8c",  x"ba",  x"68",  x"ee",  x"86", -- 17F8
         x"fd",  x"49",  x"f8",  x"bb",  x"0f",  x"8c",  x"30",  x"23", -- 1800
         x"dc",  x"be",  x"c4",  x"58",  x"d4",  x"ae",  x"bc",  x"2b", -- 1808
         x"e1",  x"50",  x"0e",  x"b8",  x"1d",  x"c0",  x"16",  x"cf", -- 1810
         x"80",  x"bd",  x"c7",  x"f9",  x"fe",  x"8c",  x"1e",  x"04", -- 1818
         x"3d",  x"20",  x"f0",  x"4e",  x"24",  x"23",  x"80",  x"eb", -- 1820
         x"20",  x"07",  x"3a",  x"eb",  x"ff",  x"db",  x"27",  x"87", -- 1828
         x"a2",  x"7e",  x"50",  x"43",  x"e1",  x"0c",  x"01",  x"3a", -- 1830
         x"0e",  x"00",  x"9a",  x"8a",  x"79",  x"48",  x"c6",  x"81", -- 1838
         x"c8",  x"b8",  x"c8",  x"6a",  x"95",  x"f3",  x"05",  x"18", -- 1840
         x"f4",  x"cd",  x"06",  x"cf",  x"18",  x"c0",  x"b4",  x"d5", -- 1848
         x"3a",  x"62",  x"ae",  x"c2",  x"cd",  x"ca",  x"2e",  x"f1", -- 1850
         x"e3",  x"d2",  x"10",  x"1f",  x"cd",  x"2b",  x"cd",  x"36", -- 1858
         x"28",  x"35",  x"69",  x"e5",  x"f7",  x"cb",  x"23",  x"8f", -- 1860
         x"3c",  x"a0",  x"ac",  x"72",  x"30",  x"12",  x"a7",  x"9e", -- 1868
         x"93",  x"b3",  x"34",  x"e8",  x"49",  x"c0",  x"10",  x"e8", -- 1870
         x"ea",  x"d1",  x"cd",  x"1b",  x"64",  x"d3",  x"b9",  x"66", -- 1878
         x"bc",  x"06",  x"ed",  x"19",  x"fa",  x"e3",  x"d1",  x"c2", -- 1880
         x"3d",  x"f7",  x"c2",  x"a8",  x"cb",  x"1d",  x"21",  x"d4", -- 1888
         x"7e",  x"c9",  x"36",  x"8c",  x"fc",  x"a3",  x"5b",  x"88", -- 1890
         x"2b",  x"a2",  x"e1",  x"78",  x"ca",  x"92",  x"88",  x"e8", -- 1898
         x"87",  x"c9",  x"fe",  x"39",  x"2c",  x"c0",  x"b7",  x"ac", -- 18A0
         x"65",  x"93",  x"d2",  x"88",  x"35",  x"1a",  x"a9",  x"67", -- 18A8
         x"29",  x"88",  x"fd",  x"20",  x"08",  x"23",  x"a0",  x"93", -- 18B0
         x"0a",  x"fe",  x"d4",  x"20",  x"f8",  x"e1",  x"10",  x"da", -- 18B8
         x"07",  x"ca",  x"c3",  x"78",  x"91",  x"2d",  x"b4",  x"99", -- 18C0
         x"18",  x"07",  x"c5",  x"3d",  x"fd",  x"68",  x"88",  x"cc", -- 18C8
         x"28",  x"5e",  x"1b",  x"d5",  x"38",  x"48",  x"09",  x"e3", -- 18D0
         x"78",  x"0f",  x"06",  x"e0",  x"fe",  x"60",  x"a5",  x"4e", -- 18D8
         x"cb",  x"fe",  x"a8",  x"28",  x"78",  x"60",  x"e5",  x"50", -- 18E0
         x"28",  x"5d",  x"fe",  x"3b",  x"ca",  x"14",  x"b2",  x"cb", -- 18E8
         x"c1",  x"55",  x"e5",  x"a0",  x"c3",  x"f3",  x"a4",  x"ef", -- 18F0
         x"d0",  x"34",  x"d8",  x"cd",  x"8a",  x"14",  x"d1",  x"36", -- 18F8
         x"20",  x"be",  x"0a",  x"34",  x"03",  x"b8",  x"88",  x"e0", -- 1900
         x"85",  x"0a",  x"04",  x"a8",  x"8c",  x"0d",  x"86",  x"3d", -- 1908
         x"b8",  x"d4",  x"c9",  x"bc",  x"77",  x"a0",  x"0f",  x"18", -- 1910
         x"a0",  x"0e",  x"2b",  x"c5",  x"61",  x"05",  x"36",  x"00", -- 1918
         x"51",  x"91",  x"3e",  x"0d",  x"70",  x"91",  x"0a",  x"af", -- 1920
         x"04",  x"70",  x"16",  x"01",  x"3a",  x"40",  x"03",  x"3d", -- 1928
         x"c8",  x"f5",  x"af",  x"4d",  x"0d",  x"f1",  x"a0",  x"09", -- 1930
         x"3a",  x"42",  x"22",  x"c6",  x"c3",  x"37",  x"30",  x"29", -- 1938
         x"d6",  x"0d",  x"ab",  x"b0",  x"20",  x"fa",  x"2f",  x"18", -- 1940
         x"62",  x"15",  x"a9",  x"1e",  x"1d",  x"d4",  x"cd",  x"db", -- 1948
         x"be",  x"e4",  x"fa",  x"a8",  x"61",  x"e5",  x"91",  x"41", -- 1950
         x"1f",  x"2f",  x"83",  x"30",  x"0b",  x"99",  x"fe",  x"08", -- 1958
         x"47",  x"27",  x"ed",  x"16",  x"10",  x"fb",  x"a8",  x"ba", -- 1960
         x"8b",  x"f8",  x"69",  x"85",  x"bb",  x"32",  x"7d",  x"8c", -- 1968
         x"1a",  x"88",  x"cc",  x"55",  x"c9",  x"3f",  x"00",  x"52", -- 1970
         x"45",  x"44",  x"4f",  x"20",  x"46",  x"52",  x"4f",  x"3b", -- 1978
         x"4d",  x"20",  x"b1",  x"1b",  x"41",  x"52",  x"54",  x"81", -- 1980
         x"94",  x"3a",  x"ce",  x"9f",  x"4c",  x"42",  x"e6",  x"8f", -- 1988
         x"21",  x"c9",  x"2c",  x"d3",  x"f3",  x"c3",  x"85",  x"fd", -- 1990
         x"22",  x"37",  x"d1",  x"aa",  x"c1",  x"d3",  x"bd",  x"a3", -- 1998
         x"10",  x"22",  x"20",  x"10",  x"cd",  x"78",  x"8b",  x"0e", -- 19A0
         x"a6",  x"9e",  x"3b",  x"e5",  x"04",  x"07",  x"d4",  x"18", -- 19A8
         x"c6",  x"18",  x"04",  x"08",  x"cf",  x"c6",  x"c1",  x"2a", -- 19B0
         x"38",  x"36",  x"bb",  x"f1",  x"af",  x"76",  x"2b",  x"d5", -- 19B8
         x"37",  x"30",  x"36",  x"2c",  x"c2",  x"cb",  x"a7",  x"ab", -- 19C0
         x"57",  x"f6",  x"31",  x"b8",  x"49",  x"e3",  x"82",  x"a3", -- 19C8
         x"f1",  x"a2",  x"d0",  x"7f",  x"e3",  x"bc",  x"42",  x"98", -- 19D0
         x"1e",  x"b2",  x"5c",  x"20",  x"7d",  x"49",  x"ee",  x"a0", -- 19D8
         x"36",  x"d1",  x"c1",  x"da",  x"1f",  x"4c",  x"c9",  x"38", -- 19E0
         x"ca",  x"2c",  x"47",  x"ca",  x"f0",  x"b6",  x"e0",  x"50", -- 19E8
         x"21",  x"a8",  x"2b",  x"57",  x"f2",  x"78",  x"e2",  x"b6", -- 19F0
         x"2c",  x"57",  x"d5",  x"a1",  x"16",  x"3a",  x"06",  x"2c", -- 19F8
         x"91",  x"94",  x"8e",  x"d1",  x"b1",  x"c0",  x"88",  x"cc", -- 1A00
         x"8b",  x"46",  x"c3",  x"77",  x"ca",  x"a1",  x"51",  x"a1", -- 1A08
         x"d7",  x"e3",  x"44",  x"d6",  x"e1",  x"a2",  x"92",  x"cb", -- 1A10
         x"b5",  x"58",  x"1e",  x"c2",  x"db",  x"cb",  x"0e",  x"0a", -- 1A18
         x"20",  x"2c",  x"93",  x"d1",  x"33",  x"eb",  x"c2",  x"68", -- 1A20
         x"f4",  x"e4",  x"b6",  x"05",  x"21",  x"ab",  x"cc",  x"c4", -- 1A28
         x"c9",  x"10",  x"f7",  x"3f",  x"45",  x"58",  x"00",  x"54", -- 1A30
         x"52",  x"41",  x"20",  x"49",  x"47",  x"4e",  x"4f",  x"a0", -- 1A38
         x"eb",  x"c2",  x"df",  x"a3",  x"d2",  x"82",  x"05",  x"11", -- 1A40
         x"b9",  x"da",  x"1e",  x"06",  x"4b",  x"f7",  x"2b",  x"dc", -- 1A48
         x"94",  x"ca",  x"03",  x"54",  x"fe",  x"1a",  x"83",  x"20", -- 1A50
         x"e2",  x"b6",  x"29",  x"cc",  x"d4",  x"58",  x"c4",  x"b0", -- 1A58
         x"51",  x"f3",  x"d2",  x"bc",  x"03",  x"c2",  x"4e",  x"c3", -- 1A60
         x"f9",  x"d5",  x"2a",  x"6a",  x"f5",  x"b3",  x"dd",  x"71", -- 1A68
         x"d6",  x"dd",  x"cb",  x"f3",  x"d4",  x"71",  x"b2",  x"75", -- 1A70
         x"ee",  x"d6",  x"46",  x"83",  x"2b",  x"c1",  x"90",  x"09", -- 1A78
         x"e1",  x"6b",  x"9b",  x"8e",  x"c5",  x"41",  x"c3",  x"50", -- 1A80
         x"c8",  x"f9",  x"2a",  x"71",  x"bc",  x"86",  x"8d",  x"da", -- 1A88
         x"96",  x"a2",  x"05",  x"df",  x"cc",  x"19",  x"80",  x"f6", -- 1A90
         x"37",  x"40",  x"d4",  x"8f",  x"0b",  x"b7",  x"e8",  x"1e", -- 1A98
         x"18",  x"c9",  x"6c",  x"b7",  x"4d",  x"28",  x"2b",  x"97", -- 1AA0
         x"86",  x"d5",  x"0e",  x"01",  x"c7",  x"b8",  x"0c",  x"ad", -- 1AA8
         x"cd",  x"22",  x"6f",  x"d1",  x"9a",  x"be",  x"02",  x"c1", -- 1AB0
         x"fa",  x"33",  x"78",  x"d4",  x"f3",  x"61",  x"7e",  x"18", -- 1AB8
         x"d6",  x"b3",  x"38",  x"15",  x"be",  x"c7",  x"cb",  x"80", -- 1AC0
         x"fe",  x"01",  x"17",  x"aa",  x"ba",  x"53",  x"57",  x"cd", -- 1AC8
         x"16",  x"22",  x"c6",  x"97",  x"03",  x"18",  x"e7",  x"7a", -- 1AD0
         x"91",  x"21",  x"84",  x"ce",  x"7e",  x"47",  x"0d",  x"d6", -- 1AD8
         x"ac",  x"e7",  x"82",  x"07",  x"d0",  x"5f",  x"80",  x"53", -- 1AE0
         x"3d",  x"b3",  x"7b",  x"ca",  x"b3",  x"d2",  x"0d",  x"07", -- 1AE8
         x"83",  x"5f",  x"21",  x"c9",  x"80",  x"19",  x"78",  x"56", -- 1AF0
         x"ba",  x"d0",  x"23",  x"a4",  x"b7",  x"19",  x"c5",  x"01", -- 1AF8
         x"49",  x"03",  x"43",  x"4a",  x"d8",  x"a0",  x"d6",  x"58", -- 1B00
         x"51",  x"ba",  x"dc",  x"f7",  x"a2",  x"32",  x"32",  x"18", -- 1B08
         x"90",  x"88",  x"59",  x"ae",  x"46",  x"1e",  x"24",  x"40", -- 1B10
         x"ee",  x"da",  x"c4",  x"b8",  x"cd",  x"8f",  x"d4",  x"a6", -- 1B18
         x"37",  x"fe",  x"03",  x"ac",  x"28",  x"e8",  x"fe",  x"2e", -- 1B20
         x"ca",  x"0d",  x"0c",  x"fe",  x"ad",  x"28",  x"19",  x"ec", -- 1B28
         x"59",  x"ca",  x"d4",  x"00",  x"fe",  x"aa",  x"ca",  x"e3", -- 1B30
         x"ce",  x"fe",  x"a7",  x"00",  x"ca",  x"f0",  x"d0",  x"d6", -- 1B38
         x"b6",  x"30",  x"28",  x"cd",  x"19",  x"36",  x"cd",  x"c3", -- 1B40
         x"cd",  x"82",  x"16",  x"7d",  x"cd",  x"3d",  x"cd",  x"83", -- 1B48
         x"a2",  x"ed",  x"02",  x"c0",  x"d6",  x"a9",  x"5e",  x"c4", -- 1B50
         x"71",  x"98",  x"6f",  x"e5",  x"9c",  x"a5",  x"c1",  x"93", -- 1B58
         x"a9",  x"cc",  x"92",  x"1f",  x"10",  x"bc",  x"6e",  x"db", -- 1B60
         x"54",  x"c5",  x"5c",  x"79",  x"0b",  x"fe",  x"33",  x"38", -- 1B68
         x"07",  x"8d",  x"5e",  x"e3",  x"5e",  x"e0",  x"4e",  x"e8", -- 1B70
         x"41",  x"fe",  x"2d",  x"38",  x"17",  x"56",  x"43",  x"fc", -- 1B78
         x"4e",  x"2a",  x"ec",  x"a9",  x"f3",  x"1d",  x"e3",  x"37", -- 1B80
         x"1f",  x"f4",  x"b4",  x"e6",  x"18",  x"08",  x"46",  x"cd", -- 1B88
         x"35",  x"e3",  x"11",  x"f2",  x"ed",  x"96",  x"94",  x"74", -- 1B90
         x"8f",  x"66",  x"30",  x"69",  x"e9",  x"f3",  x"30",  x"ad", -- 1B98
         x"c8",  x"2f",  x"c8",  x"14",  x"fe",  x"2b",  x"da",  x"06", -- 1BA0
         x"ac",  x"c1",  x"33",  x"c9",  x"b9",  x"5b",  x"f5",  x"83", -- 1BA8
         x"70",  x"fe",  x"f1",  x"18",  x"eb",  x"c1",  x"e3",  x"35", -- 1BB0
         x"e0",  x"d6",  x"f5",  x"b0",  x"0b",  x"c1",  x"79",  x"21", -- 1BB8
         x"b0",  x"00",  x"d0",  x"20",  x"05",  x"a3",  x"4f",  x"78", -- 1BC0
         x"a2",  x"e9",  x"60",  x"b3",  x"04",  x"b2",  x"e9",  x"21", -- 1BC8
         x"96",  x"ce",  x"a0",  x"86",  x"1c",  x"1f",  x"7a",  x"17", -- 1BD0
         x"ea",  x"18",  x"64",  x"78",  x"ff",  x"00",  x"c3",  x"97", -- 1BD8
         x"cd",  x"98",  x"ce",  x"79",  x"b7",  x"1b",  x"1f",  x"c1", -- 1BE0
         x"d1",  x"2e",  x"2b",  x"6a",  x"0c",  x"d9",  x"ce",  x"e5", -- 1BE8
         x"ca",  x"a2",  x"ac",  x"fa",  x"32",  x"bb",  x"32",  x"fe", -- 1BF0
         x"d2",  x"c2",  x"50",  x"23",  x"8f",  x"99",  x"d1",  x"c5", -- 1BF8
         x"1a",  x"02",  x"d3",  x"44",  x"b3",  x"f1",  x"00",  x"57", -- 1C00
         x"e1",  x"7b",  x"b2",  x"c8",  x"7a",  x"d6",  x"01",  x"00", -- 1C08
         x"d8",  x"af",  x"bb",  x"3c",  x"d0",  x"15",  x"1d",  x"0a", -- 1C10
         x"ef",  x"81",  x"9c",  x"90",  x"ed",  x"3f",  x"c3",  x"a2", -- 1C18
         x"00",  x"d6",  x"3c",  x"8f",  x"c1",  x"a0",  x"c6",  x"ff", -- 1C20
         x"9f",  x"05",  x"c3",  x"a9",  x"d6",  x"16",  x"5a",  x"04", -- 1C28
         x"fb",  x"a0",  x"87",  x"7b",  x"06",  x"2f",  x"4f",  x"7a", -- 1C30
         x"2f",  x"cd",  x"7d",  x"c1",  x"63",  x"c3",  x"de",  x"46", -- 1C38
         x"e6",  x"c8",  x"a0",  x"d5",  x"0a",  x"01",  x"fa",  x"ce", -- 1C40
         x"c5",  x"e1",  x"41",  x"ad",  x"03",  x"46",  x"8d",  x"ce", -- 1C48
         x"c9",  x"f7",  x"af",  x"4f",  x"28",  x"e4",  x"94",  x"38", -- 1C50
         x"05",  x"0f",  x"38",  x"2d",  x"0b",  x"4f",  x"0a",  x"fb", -- 1C58
         x"62",  x"e9",  x"f6",  x"05",  x"d6",  x"24",  x"20",  x"0a", -- 1C60
         x"3c",  x"16",  x"1c",  x"0f",  x"81",  x"14",  x"3a",  x"f4", -- 1C68
         x"d8",  x"3d",  x"ca",  x"03",  x"dd",  x"cf",  x"f2",  x"48", -- 1C70
         x"cf",  x"7e",  x"b9",  x"33",  x"28",  x"6f",  x"41",  x"c1", -- 1C78
         x"0f",  x"e5",  x"50",  x"59",  x"2a",  x"df",  x"70",  x"bc", -- 1C80
         x"11",  x"01",  x"e1",  x"03",  x"ca",  x"e0",  x"d5",  x"2a", -- 1C88
         x"d9",  x"df",  x"84",  x"8c",  x"57",  x"0f",  x"d0",  x"ae", -- 1C90
         x"79",  x"96",  x"23",  x"18",  x"20",  x"02",  x"78",  x"04", -- 1C98
         x"28",  x"38",  x"23",  x"a7",  x"00",  x"18",  x"cf",  x"5a", -- 1CA0
         x"ff",  x"3b",  x"11",  x"55",  x"f0",  x"8f",  x"d8",  x"31", -- 1CA8
         x"d0",  x"cb",  x"ed",  x"fd",  x"13",  x"2a",  x"db",  x"3f", -- 1CB0
         x"57",  x"09",  x"a7",  x"1c",  x"ab",  x"c4",  x"e0",  x"fc", -- 1CB8
         x"0a",  x"fa",  x"b6",  x"22",  x"3d",  x"2b",  x"c0",  x"f5", -- 1CC0
         x"21",  x"c0",  x"b7",  x"d1",  x"73",  x"23",  x"33",  x"72", -- 1CC8
         x"23",  x"32",  x"c9",  x"32",  x"bc",  x"b1",  x"21",  x"20", -- 1CD0
         x"c3",  x"45",  x"b4",  x"ed",  x"0a",  x"97",  x"80",  x"b0", -- 1CD8
         x"e3",  x"57",  x"d5",  x"c8",  x"b0",  x"5b",  x"c9",  x"63", -- 1CE0
         x"c1",  x"dc",  x"44",  x"92",  x"3c",  x"5b",  x"57",  x"96", -- 1CE8
         x"29",  x"ee",  x"b8",  x"e9",  x"8b",  x"3c",  x"41",  x"1d", -- 1CF0
         x"1e",  x"00",  x"fb",  x"61",  x"ce",  x"a0",  x"83",  x"3f", -- 1CF8
         x"3e",  x"19",  x"c1",  x"ec",  x"50",  x"85",  x"35",  x"aa", -- 1D00
         x"50",  x"b9",  x"85",  x"16",  x"7e",  x"b8",  x"a9",  x"b9", -- 1D08
         x"08",  x"e8",  x"3a",  x"e8",  x"24",  x"8d",  x"51",  x"00", -- 1D10
         x"c3",  x"f1",  x"44",  x"4d",  x"ca",  x"aa",  x"cf",  x"96", -- 1D18
         x"0a",  x"28",  x"5f",  x"1e",  x"10",  x"d9",  x"47",  x"11", -- 1D20
         x"d2",  x"e0",  x"f1",  x"ca",  x"67",  x"c9",  x"71",  x"0a", -- 1D28
         x"23",  x"70",  x"23",  x"4f",  x"db",  x"4c",  x"ab",  x"29", -- 1D30
         x"ab",  x"3a",  x"0c",  x"2a",  x"00",  x"17",  x"79",  x"01", -- 1D38
         x"0b",  x"00",  x"30",  x"02",  x"c1",  x"59",  x"03",  x"1a", -- 1D40
         x"f5",  x"e5",  x"b0",  x"4f",  x"d7",  x"91",  x"00",  x"f1", -- 1D48
         x"3d",  x"20",  x"ea",  x"f5",  x"42",  x"4b",  x"eb",  x"55", -- 1D50
         x"19",  x"f7",  x"98",  x"cd",  x"30",  x"99",  x"73",  x"66", -- 1D58
         x"81",  x"b2",  x"03",  x"57",  x"48",  x"b0",  x"5e",  x"02", -- 1D60
         x"eb",  x"29",  x"09",  x"eb",  x"2b",  x"2b",  x"c0",  x"bd", -- 1D68
         x"f1",  x"38",  x"19",  x"22",  x"47",  x"4f",  x"bb",  x"16", -- 1D70
         x"16",  x"e1",  x"7a",  x"e3",  x"5d",  x"f5",  x"e0",  x"2c", -- 1D78
         x"90",  x"43",  x"d1",  x"19",  x"fc",  x"43",  x"7f",  x"8b", -- 1D80
         x"07",  x"29",  x"29",  x"c1",  x"2a",  x"48",  x"9f",  x"c9", -- 1D88
         x"b0",  x"ab",  x"6c",  x"21",  x"b7",  x"39",  x"91",  x"c1", -- 1D90
         x"d4",  x"0d",  x"f0",  x"43",  x"cd",  x"09",  x"d2",  x"13", -- 1D98
         x"ec",  x"9b",  x"2a",  x"c4",  x"78",  x"03",  x"e2",  x"4f", -- 1DA0
         x"f0",  x"e2",  x"41",  x"50",  x"c1",  x"d8",  x"21",  x"81", -- 1DA8
         x"1b",  x"73",  x"06",  x"90",  x"c3",  x"ae",  x"d6",  x"52", -- 1DB0
         x"9c",  x"47",  x"02",  x"af",  x"18",  x"ed",  x"cd",  x"45", -- 1DB8
         x"d1",  x"a1",  x"da",  x"01",  x"b9",  x"8e",  x"c5",  x"d5", -- 1DC0
         x"6d",  x"98",  x"69",  x"da",  x"85",  x"76",  x"56",  x"2b", -- 1DC8
         x"5e",  x"e1",  x"96",  x"f4",  x"90",  x"37",  x"82",  x"9a", -- 1DD0
         x"63",  x"e3",  x"80",  x"b7",  x"c3",  x"84",  x"ff",  x"28", -- 1DD8
         x"2b",  x"24",  x"18",  x"a5",  x"19",  x"e3",  x"80",  x"8a", -- 1DE0
         x"7a",  x"b3",  x"ca",  x"30",  x"54",  x"c3",  x"97",  x"14", -- 1DE8
         x"66",  x"6f",  x"e5",  x"b9",  x"5e",  x"9e",  x"63",  x"03", -- 1DF0
         x"2a",  x"e3",  x"03",  x"0a",  x"6f",  x"e1",  x"03",  x"21", -- 1DF8
         x"03",  x"27",  x"b7",  x"a1",  x"fa",  x"b3",  x"5d",  x"e2", -- 1E00
         x"c7",  x"d3",  x"11",  x"ff",  x"03",  x"1d",  x"03",  x"24", -- 1E08
         x"b1",  x"ff",  x"93",  x"84",  x"42",  x"e1",  x"c0",  x"1e", -- 1E10
         x"16",  x"57",  x"8e",  x"14",  x"a7",  x"3e",  x"80",  x"81", -- 1E18
         x"60",  x"b6",  x"47",  x"cd",  x"0b",  x"cf",  x"2e",  x"c3", -- 1E20
         x"29",  x"5e",  x"5b",  x"a9",  x"a0",  x"c0",  x"0a",  x"01", -- 1E28
         x"57",  x"d3",  x"c5",  x"b5",  x"47",  x"e5",  x"75",  x"c5", -- 1E30
         x"c3",  x"26",  x"ba",  x"9e",  x"e0",  x"d1",  x"e5",  x"6f", -- 1E38
         x"cd",  x"f2",  x"15",  x"d2",  x"d1",  x"c9",  x"10",  x"e6", -- 1E40
         x"eb",  x"69",  x"77",  x"e8",  x"1b",  x"a1",  x"70",  x"52", -- 1E48
         x"2b",  x"06",  x"22",  x"50",  x"19",  x"e5",  x"0e",  x"ff", -- 1E50
         x"a4",  x"30",  x"0c",  x"f8",  x"3a",  x"06",  x"ba",  x"f9", -- 1E58
         x"1a",  x"b8",  x"20",  x"f4",  x"ff",  x"b3",  x"cc",  x"e8", -- 1E60
         x"64",  x"e3",  x"fa",  x"79",  x"a6",  x"34",  x"11",  x"2a", -- 1E68
         x"2a",  x"28",  x"b2",  x"03",  x"fc",  x"8b",  x"3e",  x"01", -- 1E70
         x"a0",  x"4f",  x"8f",  x"68",  x"c3",  x"59",  x"22",  x"10", -- 1E78
         x"e1",  x"7e",  x"82",  x"82",  x"1e",  x"81",  x"82",  x"23", -- 1E80
         x"2d",  x"6c",  x"28",  x"92",  x"1c",  x"1d",  x"c8",  x"bb", -- 1E88
         x"ed",  x"06",  x"fe",  x"0d",  x"cc",  x"66",  x"cb",  x"b3", -- 1E90
         x"e0",  x"f2",  x"b7",  x"0e",  x"f1",  x"f5",  x"98",  x"c0", -- 1E98
         x"74",  x"fc",  x"1f",  x"06",  x"ff",  x"09",  x"28",  x"37", -- 1EA0
         x"b3",  x"e0",  x"22",  x"0d",  x"db",  x"56",  x"f1",  x"8b", -- 1EA8
         x"00",  x"1e",  x"1a",  x"28",  x"c2",  x"bf",  x"f5",  x"01", -- 1EB0
         x"6b",  x"e3",  x"d0",  x"5f",  x"d5",  x"d8",  x"14",  x"fa", -- 1EB8
         x"e1",  x"da",  x"e0",  x"2c",  x"fe",  x"b4",  x"7d",  x"03", -- 1EC0
         x"34",  x"5d",  x"02",  x"2b",  x"01",  x"1a",  x"d2",  x"20", -- 1EC8
         x"3f",  x"93",  x"c6",  x"0e",  x"5f",  x"d9",  x"0e",  x"ec", -- 1ED0
         x"94",  x"cb",  x"00",  x"b7",  x"cd",  x"68",  x"d2",  x"18", -- 1ED8
         x"27",  x"ee",  x"c1",  x"d7",  x"35",  x"49",  x"34",  x"75", -- 1EE0
         x"7b",  x"bc",  x"0a",  x"b7",  x"f2",  x"3b",  x"d2",  x"ad", -- 1EE8
         x"3c",  x"e4",  x"34",  x"cc",  x"7f",  x"09",  x"66",  x"1c", -- 1EF0
         x"0a",  x"61",  x"1c",  x"da",  x"01",  x"59",  x"d2",  x"aa", -- 1EF8
         x"e0",  x"80",  x"ac",  x"35",  x"ef",  x"5e",  x"f0",  x"97", -- 1F00
         x"e5",  x"8a",  x"85",  x"8a",  x"e8",  x"19",  x"e2",  x"d8", -- 1F08
         x"d6",  x"85",  x"b4",  x"07",  x"bc",  x"f6",  x"09",  x"90", -- 1F10
         x"1a",  x"f1",  x"f1",  x"e5",  x"cd",  x"55",  x"e5",  x"1b", -- 1F18
         x"7d",  x"b4",  x"b7",  x"86",  x"46",  x"2b",  x"4e",  x"e5", -- 1F20
         x"b6",  x"67",  x"6e",  x"26",  x"46",  x"aa",  x"d0",  x"2b", -- 1F28
         x"56",  x"2e",  x"ae",  x"95",  x"b4",  x"bf",  x"5d",  x"9b", -- 1F30
         x"0e",  x"2b",  x"c3",  x"0c",  x"4d",  x"ff",  x"bc",  x"39", -- 1F38
         x"e7",  x"f5",  x"03",  x"e1",  x"91",  x"7e",  x"27",  x"c9", -- 1F40
         x"85",  x"86",  x"1e",  x"1c",  x"da",  x"10",  x"86",  x"7b", -- 1F48
         x"d1",  x"d1",  x"a7",  x"96",  x"cd",  x"16",  x"01",  x"d3", -- 1F50
         x"15",  x"c2",  x"a8",  x"fc",  x"cd",  x"e9",  x"d2",  x"a6", -- 1F58
         x"02",  x"21",  x"f2",  x"39",  x"62",  x"18",  x"6f",  x"ca", -- 1F60
         x"6b",  x"ba",  x"e7",  x"6f",  x"2c",  x"a0",  x"00",  x"0a", -- 1F68
         x"12",  x"03",  x"13",  x"18",  x"57",  x"f8",  x"3d",  x"3b", -- 1F70
         x"df",  x"25",  x"e5",  x"99",  x"c0",  x"d5",  x"69",  x"1b", -- 1F78
         x"4e",  x"28",  x"97",  x"70",  x"99",  x"47",  x"50",  x"09", -- 1F80
         x"89",  x"e5",  x"90",  x"43",  x"ee",  x"61",  x"8a",  x"85", -- 1F88
         x"89",  x"28",  x"14",  x"c0",  x"ea",  x"43",  x"c9",  x"01", -- 1F90
         x"c0",  x"d0",  x"f0",  x"50",  x"fb",  x"d2",  x"af",  x"57", -- 1F98
         x"a2",  x"80",  x"f2",  x"e9",  x"50",  x"0e",  x"30",  x"d3", -- 1FA0
         x"28",  x"55",  x"90",  x"da",  x"0c",  x"1a",  x"c9",  x"98", -- 1FA8
         x"b0",  x"80",  x"ca",  x"7f",  x"24",  x"d4",  x"7a",  x"6e", -- 1FB0
         x"73",  x"e0",  x"a9",  x"c0",  x"0a",  x"da",  x"d3",  x"af", -- 1FB8
         x"e3",  x"4f",  x"e5",  x"d7",  x"ef",  x"d8",  x"e0",  x"78", -- 1FC0
         x"11",  x"0e",  x"00",  x"f2",  x"2b",  x"ef",  x"1f",  x"c1", -- 1FC8
         x"e1",  x"e5",  x"2c",  x"cd",  x"45",  x"66",  x"68",  x"0e", -- 1FD0
         x"a2",  x"d8",  x"14",  x"d5",  x"56",  x"89",  x"76",  x"b3", -- 1FD8
         x"05",  x"18",  x"cf",  x"68",  x"2d",  x"99",  x"1a",  x"39", -- 1FE0
         x"90",  x"18",  x"e3",  x"02",  x"7e",  x"cd",  x"de",  x"d3", -- 1FE8
         x"04",  x"05",  x"98",  x"84",  x"c5",  x"1e",  x"19",  x"ff", -- 1FF0
         x"fe",  x"29",  x"8b",  x"dc",  x"fa",  x"af",  x"21",  x"92", -- 1FF8
         x"c3",  x"f1",  x"e3",  x"01",  x"61",  x"cb",  x"33",  x"3d", -- 2000
         x"be",  x"3c",  x"6a",  x"d0",  x"cb",  x"91",  x"05",  x"bb", -- 2008
         x"47",  x"d8",  x"43",  x"c9",  x"07",  x"7f",  x"ca",  x"cf", -- 2010
         x"d4",  x"5f",  x"54",  x"22",  x"c3",  x"06",  x"19",  x"46", -- 2018
         x"72",  x"e3",  x"eb",  x"75",  x"d2",  x"b8",  x"67",  x"70", -- 2020
         x"c9",  x"eb",  x"ae",  x"31",  x"c2",  x"55",  x"c5",  x"23", -- 2028
         x"80",  x"92",  x"4f",  x"ed",  x"78",  x"60",  x"c3",  x"ad", -- 2030
         x"cd",  x"3e",  x"14",  x"d4",  x"81",  x"07",  x"03",  x"4f", -- 2038
         x"7b",  x"ed",  x"79",  x"13",  x"b5",  x"0a",  x"f5",  x"c8", -- 2040
         x"bd",  x"f4",  x"99",  x"5e",  x"c1",  x"78",  x"19",  x"25", -- 2048
         x"ab",  x"a0",  x"28",  x"5f",  x"fa",  x"d3",  x"ba",  x"32", -- 2050
         x"0d",  x"17",  x"5e",  x"2b",  x"fd",  x"52",  x"80",  x"95", -- 2058
         x"61",  x"c9",  x"b7",  x"98",  x"8f",  x"53",  x"2e",  x"7b", -- 2060
         x"04",  x"e4",  x"c5",  x"1a",  x"18",  x"04",  x"b2",  x"cd", -- 2068
         x"6c",  x"c9",  x"d5",  x"a5",  x"38",  x"d1",  x"12",  x"b0", -- 2070
         x"12",  x"eb",  x"d4",  x"09",  x"7e",  x"c3",  x"b1",  x"d0", -- 2078
         x"f4",  x"16",  x"06",  x"e3",  x"88",  x"d3",  x"21",  x"28", -- 2080
         x"04",  x"d9",  x"9b",  x"ca",  x"18",  x"09",  x"04",  x"61", -- 2088
         x"21",  x"8b",  x"56",  x"fb",  x"78",  x"c9",  x"ff",  x"3a", -- 2090
         x"c3",  x"c5",  x"b7",  x"9d",  x"90",  x"d6",  x"90",  x"30", -- 2098
         x"0c",  x"15",  x"2f",  x"3c",  x"eb",  x"e0",  x"97",  x"97", -- 20A0
         x"78",  x"1b",  x"fe",  x"19",  x"d0",  x"dc",  x"95",  x"03", -- 20A8
         x"d7",  x"32",  x"67",  x"f1",  x"93",  x"19",  x"d5",  x"b4", -- 20B0
         x"21",  x"96",  x"18",  x"f2",  x"ab",  x"f1",  x"00",  x"0a", -- 20B8
         x"d5",  x"30",  x"4b",  x"23",  x"34",  x"28",  x"31",  x"63", -- 20C0
         x"2e",  x"d8",  x"00",  x"3e",  x"d5",  x"18",  x"40",  x"af", -- 20C8
         x"90",  x"47",  x"7e",  x"33",  x"9b",  x"5f",  x"67",  x"9a", -- 20D0
         x"57",  x"03",  x"00",  x"99",  x"4f",  x"dc",  x"16",  x"d5", -- 20D8
         x"68",  x"63",  x"af",  x"76",  x"47",  x"a7",  x"20",  x"00", -- 20E0
         x"16",  x"4a",  x"54",  x"65",  x"6f",  x"78",  x"d6",  x"08", -- 20E8
         x"0e",  x"fe",  x"e0",  x"20",  x"f0",  x"86",  x"b0",  x"5d", -- 20F0
         x"c9",  x"05",  x"29",  x"cb",  x"00",  x"12",  x"cb",  x"11", -- 20F8
         x"f2",  x"d4",  x"d4",  x"78",  x"5c",  x"6a",  x"45",  x"cb", -- 2100
         x"08",  x"60",  x"21",  x"12",  x"86",  x"77",  x"30",  x"e5", -- 2108
         x"c8",  x"78",  x"78",  x"08",  x"79",  x"fc",  x"fd",  x"d4", -- 2110
         x"a0",  x"aa",  x"06",  x"e6",  x"80",  x"a9",  x"4f",  x"c3", -- 2118
         x"76",  x"1c",  x"00",  x"c0",  x"14",  x"c0",  x"0c",  x"c0", -- 2120
         x"0e",  x"80",  x"34",  x"02",  x"c0",  x"c3",  x"53",  x"d6", -- 2128
         x"7e",  x"83",  x"94",  x"5b",  x"8a",  x"5b",  x"89",  x"60", -- 2130
         x"4f",  x"b7",  x"e9",  x"c8",  x"e0",  x"2f",  x"77",  x"36", -- 2138
         x"af",  x"6f",  x"71",  x"7d",  x"71",  x"7d",  x"dd",  x"70", -- 2140
         x"7d",  x"6f",  x"6f",  x"a0",  x"62",  x"a8",  x"b8",  x"43", -- 2148
         x"5a",  x"51",  x"c8",  x"ca",  x"18",  x"f5",  x"3a",  x"c6", -- 2150
         x"09",  x"f1",  x"cc",  x"c7",  x"79",  x"1f",  x"01",  x"4f", -- 2158
         x"cb",  x"1a",  x"cb",  x"1b",  x"cb",  x"18",  x"ab",  x"e6", -- 2160
         x"00",  x"00",  x"00",  x"81",  x"03",  x"aa",  x"56",  x"19", -- 2168
         x"80",  x"f1",  x"22",  x"00",  x"76",  x"80",  x"45",  x"aa", -- 2170
         x"38",  x"82",  x"cd",  x"97",  x"18",  x"d6",  x"b7",  x"ea", -- 2178
         x"b3",  x"f8",  x"73",  x"49",  x"01",  x"35",  x"80",  x"f4", -- 2180
         x"a6",  x"04",  x"90",  x"2a",  x"f5",  x"70",  x"af",  x"98", -- 2188
         x"6f",  x"e9",  x"80",  x"d1",  x"04",  x"cd",  x"f5",  x"d5", -- 2190
         x"21",  x"48",  x"c4",  x"a8",  x"66",  x"d4",  x"30",  x"21", -- 2198
         x"4c",  x"05",  x"ce",  x"d9",  x"01",  x"80",  x"fa",  x"1f", -- 21A0
         x"3e",  x"1a",  x"c0",  x"fc",  x"0b",  x"d8",  x"32",  x"01", -- 21A8
         x"31",  x"0c",  x"18",  x"72",  x"c7",  x"ad",  x"40",  x"30", -- 21B0
         x"c8",  x"2e",  x"15",  x"58",  x"d6",  x"79",  x"32",  x"68", -- 21B8
         x"f7",  x"a5",  x"22",  x"e5",  x"d2",  x"01",  x"81",  x"23", -- 21C0
         x"50",  x"58",  x"21",  x"bc",  x"d4",  x"e5",  x"9b",  x"03", -- 21C8
         x"d5",  x"e5",  x"04",  x"e5",  x"58",  x"d9",  x"88",  x"28", -- 21D0
         x"80",  x"06",  x"2e",  x"08",  x"1f",  x"67",  x"79",  x"30", -- 21D8
         x"0b",  x"d3",  x"f1",  x"21",  x"74",  x"19",  x"92",  x"3a", -- 21E0
         x"d3",  x"2b",  x"89",  x"80",  x"95",  x"2d",  x"7c",  x"20", -- 21E8
         x"65",  x"e4",  x"83",  x"41",  x"b1",  x"85",  x"bc",  x"08", -- 21F0
         x"e7",  x"01",  x"20",  x"84",  x"bb",  x"65",  x"ec",  x"1a", -- 21F8
         x"5a",  x"05",  x"ca",  x"4b",  x"c3",  x"2e",  x"ff",  x"00", -- 2200
         x"5c",  x"34",  x"34",  x"2b",  x"7e",  x"32",  x"14",  x"03", -- 2208
         x"a5",  x"04",  x"10",  x"87",  x"04",  x"0c",  x"03",  x"41", -- 2210
         x"eb",  x"81",  x"a1",  x"57",  x"5f",  x"32",  x"17",  x"ab", -- 2218
         x"d4",  x"c5",  x"b3",  x"f0",  x"0b",  x"03",  x"de",  x"00", -- 2220
         x"15",  x"3f",  x"30",  x"07",  x"0d",  x"b1",  x"9f",  x"37", -- 2228
         x"d2",  x"98",  x"d5",  x"79",  x"3c",  x"3d",  x"01",  x"1f", -- 2230
         x"fa",  x"ec",  x"d4",  x"17",  x"cb",  x"13",  x"63",  x"e1", -- 2238
         x"89",  x"e6",  x"10",  x"3a",  x"a8",  x"19",  x"17",  x"1d", -- 2240
         x"79",  x"b2",  x"39",  x"b3",  x"20",  x"f4",  x"a0",  x"eb", -- 2248
         x"02",  x"35",  x"e1",  x"20",  x"c7",  x"1e",  x"0a",  x"a3", -- 2250
         x"8f",  x"e8",  x"20",  x"ca",  x"7c",  x"d6",  x"7d",  x"a0", -- 2258
         x"11",  x"ae",  x"80",  x"47",  x"1f",  x"00",  x"a8",  x"78", -- 2260
         x"f2",  x"7b",  x"d6",  x"c6",  x"80",  x"77",  x"ad",  x"94", -- 2268
         x"a2",  x"e3",  x"7f",  x"77",  x"98",  x"40",  x"80",  x"2f", -- 2270
         x"0d",  x"e1",  x"b7",  x"e1",  x"f2",  x"ba",  x"18",  x"18", -- 2278
         x"8c",  x"2c",  x"eb",  x"95",  x"c1",  x"c6",  x"02",  x"38", -- 2280
         x"c7",  x"47",  x"43",  x"82",  x"59",  x"31",  x"8d",  x"16", -- 2288
         x"18",  x"bc",  x"a4",  x"79",  x"a9",  x"80",  x"e7",  x"03", -- 2290
         x"fe",  x"2f",  x"17",  x"9f",  x"c0",  x"59",  x"3c",  x"2f", -- 2298
         x"06",  x"88",  x"41",  x"bd",  x"46",  x"1d",  x"4f",  x"70", -- 22A0
         x"88",  x"40",  x"23",  x"36",  x"80",  x"17",  x"c3",  x"28", -- 22A8
         x"b9",  x"d4",  x"15",  x"f0",  x"21",  x"cf",  x"23",  x"7e", -- 22B0
         x"ee",  x"59",  x"80",  x"4b",  x"93",  x"7c",  x"83",  x"7a", -- 22B8
         x"0d",  x"8b",  x"dd",  x"99",  x"80",  x"49",  x"82",  x"11", -- 22C0
         x"db",  x"0f",  x"18",  x"51",  x"03",  x"f6",  x"99",  x"ed", -- 22C8
         x"53",  x"17",  x"ed",  x"43",  x"ed",  x"16",  x"df",  x"97", -- 22D0
         x"8a",  x"09",  x"71",  x"82",  x"4e",  x"83",  x"23",  x"30", -- 22D8
         x"c9",  x"11",  x"0b",  x"06",  x"04",  x"1a",  x"77",  x"1a", -- 22E0
         x"13",  x"23",  x"10",  x"ee",  x"58",  x"42",  x"07",  x"37", -- 22E8
         x"1f",  x"1a",  x"77",  x"3f",  x"1f",  x"c6",  x"94",  x"77", -- 22F0
         x"79",  x"09",  x"4f",  x"14",  x"1f",  x"ae",  x"c9",  x"bf", -- 22F8
         x"18",  x"5d",  x"21",  x"a0",  x"d6",  x"51",  x"e5",  x"64", -- 2300
         x"79",  x"c8",  x"46",  x"22",  x"ae",  x"79",  x"b0",  x"e0", -- 2308
         x"32",  x"d7",  x"1f",  x"a9",  x"c9",  x"02",  x"23",  x"78", -- 2310
         x"be",  x"c0",  x"2b",  x"79",  x"94",  x"03",  x"7a",  x"03", -- 2318
         x"7b",  x"18",  x"96",  x"c0",  x"e1",  x"e2",  x"a8",  x"47", -- 2320
         x"b1",  x"70",  x"ae",  x"f0",  x"2a",  x"c9",  x"a0",  x"de", -- 2328
         x"00",  x"ae",  x"67",  x"fc",  x"69",  x"d7",  x"3e",  x"98", -- 2330
         x"90",  x"a4",  x"c8",  x"19",  x"7c",  x"17",  x"dc",  x"ee", -- 2338
         x"e1",  x"ae",  x"49",  x"aa",  x"81",  x"23",  x"1b",  x"7a", -- 2340
         x"a3",  x"3c",  x"c0",  x"0b",  x"21",  x"8f",  x"8d",  x"fe", -- 2348
         x"98",  x"3a",  x"7e",  x"d0",  x"b0",  x"a7",  x"45",  x"d7", -- 2350
         x"36",  x"03",  x"98",  x"7b",  x"f5",  x"79",  x"17",  x"cd", -- 2358
         x"ca",  x"0e",  x"8a",  x"aa",  x"f9",  x"40",  x"78",  x"b1", -- 2360
         x"c8",  x"3e",  x"10",  x"29",  x"3d",  x"38",  x"06",  x"b6", -- 2368
         x"01",  x"eb",  x"30",  x"04",  x"09",  x"da",  x"0b",  x"d0", -- 2370
         x"ee",  x"de",  x"17",  x"fe",  x"00",  x"2d",  x"f5",  x"28", -- 2378
         x"05",  x"fe",  x"2b",  x"28",  x"01",  x"db",  x"8c",  x"ad", -- 2380
         x"16",  x"47",  x"67",  x"2f",  x"bf",  x"fc",  x"00",  x"38", -- 2388
         x"3d",  x"fe",  x"2e",  x"28",  x"16",  x"fe",  x"45",  x"2d", -- 2390
         x"20",  x"15",  x"a1",  x"8b",  x"4d",  x"ce",  x"12",  x"00", -- 2398
         x"4b",  x"14",  x"20",  x"07",  x"af",  x"93",  x"5f",  x"0c", -- 23A0
         x"00",  x"0c",  x"28",  x"de",  x"e5",  x"7b",  x"90",  x"f4", -- 23A8
         x"ed",  x"0d",  x"d7",  x"f2",  x"e4",  x"d7",  x"d2",  x"40", -- 23B0
         x"e7",  x"d5",  x"f1",  x"3c",  x"20",  x"f2",  x"1a",  x"d1", -- 23B8
         x"f1",  x"cc",  x"fb",  x"e2",  x"97",  x"c8",  x"cf",  x"0f", -- 23C0
         x"82",  x"d6",  x"f0",  x"76",  x"a3",  x"0e",  x"57",  x"78", -- 23C8
         x"89",  x"47",  x"c6",  x"56",  x"d5",  x"0d",  x"d6",  x"51", -- 23D0
         x"30",  x"f4",  x"b3",  x"e1",  x"93",  x"28",  x"18",  x"a8", -- 23D8
         x"a3",  x"ca",  x"cd",  x"a9",  x"9d",  x"36",  x"c3",  x"85", -- 23E0
         x"40",  x"7b",  x"07",  x"07",  x"83",  x"07",  x"63",  x"86", -- 23E8
         x"1a",  x"5f",  x"18",  x"a5",  x"d5",  x"27",  x"0d",  x"d8", -- 23F0
         x"35",  x"98",  x"59",  x"96",  x"9d",  x"06",  x"98",  x"86", -- 23F8
         x"62",  x"92",  x"c8",  x"65",  x"d1",  x"11",  x"ea",  x"03", -- 2400
         x"8b",  x"96",  x"36",  x"57",  x"0c",  x"42",  x"d8",  x"36", -- 2408
         x"2d",  x"8c",  x"80",  x"30",  x"ca",  x"ef",  x"d8",  x"e5", -- 2410
         x"fc",  x"db",  x"60",  x"af",  x"5e",  x"f5",  x"bf",  x"40", -- 2418
         x"43",  x"91",  x"11",  x"f8",  x"c0",  x"a3",  x"18",  x"d7", -- 2420
         x"0d",  x"b7",  x"e2",  x"6e",  x"d8",  x"d0",  x"18",  x"ee", -- 2428
         x"83",  x"12",  x"18",  x"ec",  x"05",  x"85",  x"85",  x"1c", -- 2430
         x"cd",  x"5e",  x"d4",  x"3c",  x"05",  x"f6",  x"23",  x"84", -- 2438
         x"01",  x"e0",  x"70",  x"f1",  x"81",  x"3c",  x"fa",  x"0c", -- 2440
         x"89",  x"d8",  x"fe",  x"08",  x"eb",  x"00",  x"3c",  x"47", -- 2448
         x"3e",  x"02",  x"3d",  x"3d",  x"00",  x"e1",  x"f5",  x"11", -- 2450
         x"08",  x"d9",  x"05",  x"20",  x"06",  x"28",  x"36",  x"2e", -- 2458
         x"52",  x"23",  x"05",  x"c5",  x"06",  x"cc",  x"f5",  x"d6", -- 2460
         x"86",  x"a4",  x"d5",  x"21",  x"e1",  x"06",  x"2f",  x"04", -- 2468
         x"8e",  x"e9",  x"9e",  x"c6",  x"7a",  x"9e",  x"9e",  x"c3", -- 2470
         x"79",  x"9e",  x"4f",  x"91",  x"a2",  x"30",  x"f0",  x"9d", -- 2478
         x"9c",  x"23",  x"5a",  x"46",  x"f0",  x"00",  x"70",  x"23", -- 2480
         x"c1",  x"0d",  x"20",  x"d2",  x"05",  x"34",  x"28",  x"0b", -- 2488
         x"bd",  x"38",  x"fe",  x"30",  x"bc",  x"c5",  x"97",  x"c4", -- 2490
         x"83",  x"35",  x"f1",  x"28",  x"1a",  x"36",  x"45",  x"44", -- 2498
         x"63",  x"2b",  x"81",  x"41",  x"9f",  x"bd",  x"e5",  x"00", -- 24A0
         x"3d",  x"d6",  x"0a",  x"30",  x"fb",  x"c6",  x"3a",  x"23", -- 24A8
         x"fd",  x"2c",  x"ed",  x"64",  x"71",  x"8b",  x"01",  x"05", -- 24B0
         x"74",  x"94",  x"11",  x"f7",  x"23",  x"80",  x"a3",  x"e1", -- 24B8
         x"e2",  x"65",  x"29",  x"d8",  x"e9",  x"bb",  x"80",  x"80", -- 24C0
         x"a0",  x"86",  x"01",  x"10",  x"27",  x"64",  x"00",  x"9c", -- 24C8
         x"00",  x"6e",  x"64",  x"0c",  x"0a",  x"02",  x"97",  x"eb", -- 24D0
         x"9b",  x"e1",  x"d6",  x"e3",  x"e9",  x"43",  x"93",  x"70", -- 24D8
         x"c3",  x"dd",  x"95",  x"b4",  x"40",  x"78",  x"ca",  x"6d", -- 24E0
         x"d9",  x"f2",  x"38",  x"29",  x"d9",  x"b7",  x"bc",  x"73", -- 24E8
         x"03",  x"d0",  x"d4",  x"ce",  x"61",  x"79",  x"f6",  x"7f", -- 24F0
         x"40",  x"9e",  x"f2",  x"29",  x"55",  x"d9",  x"d9",  x"8d", -- 24F8
         x"70",  x"d7",  x"23",  x"f5",  x"43",  x"53",  x"e1",  x"7c", -- 2500
         x"1f",  x"a3",  x"fc",  x"af",  x"fc",  x"03",  x"e3",  x"85", -- 2508
         x"dc",  x"1a",  x"d9",  x"0d",  x"f7",  x"14",  x"1b",  x"59", -- 2510
         x"d5",  x"3f",  x"9a",  x"5b",  x"d5",  x"85",  x"02",  x"38", -- 2518
         x"81",  x"11",  x"3b",  x"aa",  x"a9",  x"0b",  x"e1",  x"01", -- 2520
         x"fe",  x"88",  x"d2",  x"76",  x"d6",  x"5a",  x"37",  x"99", -- 2528
         x"e8",  x"fd",  x"da",  x"d6",  x"09",  x"f5",  x"93",  x"ed", -- 2530
         x"61",  x"d5",  x"18",  x"91",  x"ac",  x"db",  x"49",  x"6c", -- 2538
         x"09",  x"ca",  x"3b",  x"21",  x"ad",  x"7c",  x"52",  x"d9", -- 2540
         x"f9",  x"0c",  x"c1",  x"4a",  x"c3",  x"33",  x"08",  x"40", -- 2548
         x"00",  x"2e",  x"94",  x"74",  x"70",  x"4f",  x"2e",  x"77", -- 2550
         x"6e",  x"00",  x"02",  x"88",  x"7a",  x"e6",  x"a0",  x"2a", -- 2558
         x"7c",  x"50",  x"01",  x"aa",  x"aa",  x"7e",  x"ff",  x"ff", -- 2560
         x"7f",  x"7f",  x"40",  x"c0",  x"81",  x"b8",  x"81",  x"a0", -- 2568
         x"60",  x"11",  x"98",  x"d5",  x"d5",  x"91",  x"89",  x"35", -- 2570
         x"2e",  x"e1",  x"6f",  x"0e",  x"a3",  x"eb",  x"3f",  x"bb", -- 2578
         x"46",  x"50",  x"3d",  x"c8",  x"87",  x"0e",  x"f5",  x"18", -- 2580
         x"f5",  x"15",  x"95",  x"f2",  x"07",  x"e3",  x"30",  x"e1", -- 2588
         x"18",  x"dd",  x"a4",  x"e2",  x"00",  x"1b",  x"03",  x"fa", -- 2590
         x"5d",  x"da",  x"21",  x"3c",  x"03",  x"ec",  x"26",  x"0b", -- 2598
         x"c8",  x"86",  x"34",  x"e6",  x"07",  x"b0",  x"c4",  x"a4", -- 25A0
         x"87",  x"87",  x"5d",  x"4f",  x"b4",  x"58",  x"a7",  x"03", -- 25A8
         x"1a",  x"03",  x"3c",  x"e6",  x"03",  x"13",  x"0c",  x"fe", -- 25B0
         x"01",  x"88",  x"32",  x"0a",  x"21",  x"60",  x"5d",  x"da", -- 25B8
         x"1a",  x"86",  x"a6",  x"62",  x"7b",  x"0d",  x"59",  x"ee", -- 25C0
         x"4f",  x"4f",  x"8a",  x"bd",  x"a4",  x"cd",  x"03",  x"21", -- 25C8
         x"19",  x"b6",  x"80",  x"7e",  x"d6",  x"ab",  x"20",  x"04", -- 25D0
         x"77",  x"0e",  x"0c",  x"15",  x"1c",  x"cd",  x"a3",  x"28", -- 25D8
         x"50",  x"c3",  x"f7",  x"6d",  x"d6",  x"e9",  x"4e",  x"01", -- 25E0
         x"18",  x"a7",  x"80",  x"b1",  x"46",  x"68",  x"99",  x"e9", -- 25E8
         x"92",  x"00",  x"69",  x"10",  x"d1",  x"75",  x"68",  x"21", -- 25F0
         x"ba",  x"da",  x"ba",  x"3c",  x"88",  x"12",  x"49",  x"83", -- 25F8
         x"9a",  x"a3",  x"58",  x"8e",  x"58",  x"f5",  x"99",  x"c8", -- 2600
         x"c0",  x"38",  x"f5",  x"6d",  x"3a",  x"be",  x"21",  x"66", -- 2608
         x"6c",  x"db",  x"37",  x"35",  x"f2",  x"a6",  x"09",  x"5e", -- 2610
         x"8c",  x"09",  x"b7",  x"f5",  x"f4",  x"8a",  x"6f",  x"17", -- 2618
         x"39",  x"28",  x"f1",  x"d4",  x"09",  x"c2",  x"da",  x"73", -- 2620
         x"c3",  x"b5",  x"ac",  x"3c",  x"49",  x"f3",  x"00",  x"7f", -- 2628
         x"05",  x"ba",  x"d7",  x"1e",  x"86",  x"03",  x"64",  x"26", -- 2630
         x"99",  x"87",  x"58",  x"34",  x"b6",  x"00",  x"e0",  x"5d", -- 2638
         x"a5",  x"86",  x"6b",  x"da",  x"18",  x"83",  x"4f",  x"38", -- 2640
         x"76",  x"da",  x"b0",  x"9a",  x"df",  x"fd",  x"5b",  x"31", -- 2648
         x"f3",  x"ec",  x"64",  x"49",  x"fc",  x"91",  x"a9",  x"a8", -- 2650
         x"2c",  x"fb",  x"43",  x"81",  x"da",  x"09",  x"db",  x"e5", -- 2658
         x"21",  x"81",  x"51",  x"59",  x"75",  x"8c",  x"e8",  x"6f", -- 2660
         x"d4",  x"13",  x"55",  x"db",  x"8a",  x"50",  x"9e",  x"00", -- 2668
         x"c9",  x"09",  x"4a",  x"d7",  x"3b",  x"78",  x"02",  x"00", -- 2670
         x"6e",  x"84",  x"7b",  x"fe",  x"c1",  x"2f",  x"7c",  x"74", -- 2678
         x"00",  x"31",  x"9a",  x"7d",  x"84",  x"3d",  x"5a",  x"7d", -- 2680
         x"c8",  x"00",  x"7f",  x"91",  x"7e",  x"e4",  x"bb",  x"4c", -- 2688
         x"7e",  x"6c",  x"c5",  x"f1",  x"7f",  x"20",  x"e9",  x"85", -- 2690
         x"49",  x"db",  x"28",  x"03",  x"66",  x"e7",  x"37",  x"47", -- 2698
         x"6e",  x"db",  x"f1",  x"e9",  x"cc",  x"d3",  x"fe",  x"ae", -- 26A0
         x"5c",  x"c0",  x"de",  x"ed",  x"88",  x"b0",  x"89",  x"0b", -- 26A8
         x"fe",  x"94",  x"a6",  x"9c",  x"03",  x"47",  x"d2",  x"48", -- 26B0
         x"c3",  x"d6",  x"07",  x"c3",  x"57",  x"da",  x"06",  x"b5", -- 26B8
         x"d0",  x"00",  x"00",  x"b5",  x"6f",  x"eb",  x"18",  x"e0", -- 26C0
         x"7b",  x"87",  x"a0",  x"00",  x"f6",  x"0d",  x"57",  x"1e", -- 26C8
         x"33",  x"ef",  x"18",  x"be",  x"38",  x"e5",  x"36",  x"c9", -- 26D0
         x"bf",  x"f0",  x"70",  x"f8",  x"b3",  x"cd",  x"03",  x"fe", -- 26D8
         x"d2",  x"cd",  x"09",  x"d2",  x"2a",  x"f6",  x"f0",  x"ed", -- 26E0
         x"5b",  x"56",  x"03",  x"07",  x"af",  x"ed",  x"52",  x"d1", -- 26E8
         x"e3",  x"03",  x"9a",  x"14",  x"28",  x"dd",  x"c8",  x"85", -- 26F0
         x"e4",  x"dd",  x"47",  x"e1",  x"00",  x"04",  x"12",  x"13", -- 26F8
         x"2b",  x"7d",  x"b4",  x"20",  x"f6",  x"b5",  x"0a",  x"5f", -- 2700
         x"28",  x"03",  x"57",  x"23",  x"38",  x"44",  x"7f",  x"2a", -- 2708
         x"2b",  x"40",  x"0c",  x"90",  x"ae",  x"1b",  x"7b",  x"b2", -- 2710
         x"fc",  x"1b",  x"33",  x"e8",  x"cc",  x"f8",  x"dc",  x"38", -- 2718
         x"42",  x"20",  x"60",  x"2d",  x"26",  x"77",  x"dd",  x"e3", -- 2720
         x"2b",  x"d5",  x"e9",  x"4c",  x"50",  x"b8",  x"ce",  x"82", -- 2728
         x"05",  x"e1",  x"00",  x"42",  x"4b",  x"03",  x"d1",  x"2b", -- 2730
         x"70",  x"2b",  x"71",  x"06",  x"2b",  x"35",  x"03",  x"20", -- 2738
         x"fc",  x"ab",  x"b6",  x"76",  x"f0",  x"ca",  x"25",  x"fd", -- 2740
         x"dd",  x"d9",  x"69",  x"c0",  x"85",  x"18",  x"29",  x"00", -- 2748
         x"cd",  x"87",  x"dc",  x"e5",  x"e2",  x"7b",  x"db",  x"eb", -- 2750
         x"85",  x"ad",  x"7b",  x"5e",  x"e1",  x"80",  x"5e",  x"e1", -- 2758
         x"28",  x"c7",  x"cd",  x"1d",  x"de",  x"21",  x"00",  x"3f", -- 2760
         x"dc",  x"c3",  x"71",  x"c3",  x"42",  x"41",  x"44",  x"cc", -- 2768
         x"99",  x"ae",  x"28",  x"0c",  x"c6",  x"cd",  x"b0",  x"dc", -- 2770
         x"6c",  x"d7",  x"03",  x"2a",  x"1b",  x"1b",  x"c6",  x"03", -- 2778
         x"39",  x"01",  x"d1",  x"ff",  x"41",  x"14",  x"09",  x"44", -- 2780
         x"4d",  x"43",  x"6f",  x"a2",  x"3e",  x"67",  x"e5",  x"84", -- 2788
         x"33",  x"d2",  x"3e",  x"c3",  x"4e",  x"49",  x"91",  x"19", -- 2790
         x"2a",  x"21",  x"12",  x"6e",  x"d6",  x"c3",  x"0e",  x"8a", -- 2798
         x"c4",  x"1e",  x"26",  x"ae",  x"f6",  x"0a",  x"ac",  x"59", -- 27A0
         x"cd",  x"01",  x"cc",  x"c8",  x"3b",  x"3e",  x"01",  x"32", -- 27A8
         x"cc",  x"89",  x"d6",  x"06",  x"cf",  x"58",  x"05",  x"94", -- 27B0
         x"8f",  x"60",  x"69",  x"eb",  x"d1",  x"19",  x"4e",  x"fa", -- 27B8
         x"83",  x"09",  x"09",  x"23",  x"3a",  x"ae",  x"8f",  x"b0", -- 27C0
         x"c9",  x"3e",  x"d4",  x"23",  x"00",  x"01",  x"3e",  x"d3", -- 27C8
         x"f5",  x"3a",  x"5d",  x"03",  x"a7",  x"18",  x"3e",  x"00", -- 27D0
         x"32",  x"05",  x"28",  x"04",  x"f1",  x"35",  x"c6",  x"04", -- 27D8
         x"a8",  x"72",  x"be",  x"81",  x"3a",  x"3c",  x"cd",  x"f1", -- 27E0
         x"2e",  x"09",  x"3f",  x"d3",  x"78",  x"21",  x"fe",  x"06", -- 27E8
         x"38",  x"0d",  x"2b",  x"99",  x"00",  x"10",  x"fb",  x"d5", -- 27F0
         x"11",  x"82",  x"dc",  x"73",  x"23",  x"0c",  x"72",  x"d1", -- 27F8
         x"23",  x"f1",  x"9e",  x"6d",  x"01",  x"eb",  x"80",  x"47", -- 2800
         x"79",  x"fe",  x"09",  x"38",  x"04",  x"0d",  x"23",  x"0c", -- 2808
         x"18",  x"f7",  x"ed",  x"b0",  x"b7",  x"bf",  x"ba",  x"74", -- 2810
         x"86",  x"ac",  x"dd",  x"32",  x"20",  x"fa",  x"b9",  x"0b", -- 2818
         x"4f",  x"30",  x"01",  x"04",  x"81",  x"13",  x"79",  x"c9", -- 2820
         x"5a",  x"1e",  x"07",  x"03",  x"cb",  x"bc",  x"f8",  x"7d", -- 2828
         x"06",  x"3e",  x"13",  x"20",  x"02",  x"02",  x"c6",  x"08", -- 2830
         x"32",  x"08",  x"03",  x"a0",  x"ec",  x"f1",  x"c3",  x"2c", -- 2838
         x"d5",  x"dd",  x"19",  x"47",  x"cb",  x"5a",  x"c7",  x"19", -- 2840
         x"12",  x"45",  x"19",  x"09",  x"b0",  x"19",  x"c3",  x"d2", -- 2848
         x"a0",  x"fd",  x"67",  x"24",  x"d8",  x"62",  x"80",  x"2a", -- 2850
         x"c0",  x"d4",  x"11",  x"ff",  x"30",  x"fb",  x"19",  x"f7", -- 2858
         x"61",  x"11",  x"4f",  x"cd",  x"b5",  x"dd",  x"e1",  x"9d", -- 2860
         x"9a",  x"0c",  x"33",  x"8e",  x"11",  x"43",  x"cf",  x"0e", -- 2868
         x"f6",  x"df",  x"65",  x"84",  x"db",  x"e2",  x"89",  x"50", -- 2870
         x"dd",  x"c1",  x"d0",  x"dd",  x"e6",  x"87",  x"e5",  x"a7", -- 2878
         x"e0",  x"d8",  x"9a",  x"77",  x"34",  x"77",  x"81",  x"f2", -- 2880
         x"60",  x"85",  x"f4",  x"ac",  x"1f",  x"b1",  x"92",  x"c5", -- 2888
         x"d0",  x"1d",  x"3b",  x"c1",  x"79",  x"cd",  x"ca",  x"72", -- 2890
         x"78",  x"eb",  x"04",  x"e3",  x"eb",  x"95",  x"b0",  x"28", -- 2898
         x"b4",  x"56",  x"2b",  x"64",  x"5e",  x"b8",  x"28",  x"28", -- 28A0
         x"f3",  x"1a",  x"10",  x"13",  x"0b",  x"fc",  x"fd",  x"23", -- 28A8
         x"e5",  x"da",  x"1f",  x"0d",  x"1f",  x"e1",  x"f1",  x"1f", -- 28B0
         x"cf",  x"60",  x"1a",  x"aa",  x"f6",  x"30",  x"c9",  x"3a", -- 28B8
         x"a9",  x"db",  x"b9",  x"d4",  x"5f",  x"46",  x"99",  x"23", -- 28C0
         x"3e",  x"0c",  x"d1",  x"45",  x"57",  x"14",  x"0f",  x"5f", -- 28C8
         x"7a",  x"78",  x"7b",  x"e9",  x"d8",  x"3c",  x"b3",  x"c3", -- 28D0
         x"09",  x"0c",  x"ba",  x"0b",  x"b4",  x"00",  x"7a",  x"18", -- 28D8
         x"06",  x"d5",  x"29",  x"1e",  x"80",  x"0c",  x"cb",  x"e1", -- 28E0
         x"19",  x"ef",  x"c8",  x"dd",  x"c5",  x"11",  x"42",  x"c4", -- 28E8
         x"b1",  x"06",  x"7a",  x"b0",  x"aa",  x"31",  x"3e",  x"dc", -- 28F0
         x"15",  x"1c",  x"10",  x"f8",  x"b0",  x"84",  x"e1",  x"3e", -- 28F8
         x"f5",  x"a1",  x"df",  x"eb",  x"2b",  x"06",  x"8e",  x"2f", -- 2900
         x"47",  x"83",  x"ce",  x"d9",  x"45",  x"23",  x"20",  x"31", -- 2908
         x"21",  x"da",  x"30",  x"38",  x"ee",  x"79",  x"8b",  x"28", -- 2910
         x"50",  x"12",  x"2d",  x"87",  x"fe",  x"04",  x"c0",  x"07", -- 2918
         x"30",  x"16",  x"cb",  x"4e",  x"cb",  x"ce",  x"b1",  x"8e", -- 2920
         x"51",  x"3c",  x"27",  x"e1",  x"c3",  x"90",  x"89",  x"cb", -- 2928
         x"5e",  x"cb",  x"00",  x"de",  x"18",  x"ee",  x"cb",  x"6e", -- 2930
         x"cb",  x"ee",  x"18",  x"63",  x"e8",  x"e2",  x"da",  x"03", -- 2938
         x"39",  x"30",  x"a9",  x"39",  x"8b",  x"63",  x"00",  x"3a", -- 2940
         x"10",  x"38",  x"14",  x"cb",  x"66",  x"cb",  x"4c",  x"e6", -- 2948
         x"c9",  x"3c",  x"8a",  x"00",  x"c4",  x"cb",  x"56",  x"cb", -- 2950
         x"d6",  x"18",  x"f0",  x"03",  x"cb",  x"46",  x"cb",  x"c6", -- 2958
         x"18",  x"ea",  x"38",  x"f1",  x"03",  x"8b",  x"78",  x"2a", -- 2960
         x"95",  x"23",  x"a0",  x"00",  x"01",  x"61",  x"03",  x"c5", -- 2968
         x"ae",  x"c9",  x"31",  x"d7",  x"de",  x"ae",  x"35",  x"fe", -- 2970
         x"22",  x"d6",  x"03",  x"b7",  x"28",  x"1f",  x"f2",  x"a7", -- 2978
         x"de",  x"1d",  x"15",  x"9a",  x"c7",  x"c1",  x"13",  x"80", -- 2980
         x"fa",  x"b7",  x"f2",  x"bb",  x"d3",  x"70",  x"e4",  x"98", -- 2988
         x"1e",  x"d8",  x"b7",  x"ca",  x"80",  x"3e",  x"20",  x"03", -- 2990
         x"18",  x"0c",  x"03",  x"02",  x"c4",  x"fd",  x"56",  x"fc", -- 2998
         x"18",  x"09",  x"e1",  x"d0",  x"cb",  x"28",  x"2a",  x"a5", -- 29A0
         x"43",  x"af",  x"02",  x"e1",  x"77",  x"7f",  x"cd",  x"a4", -- 29A8
         x"c5",  x"9e",  x"8e",  x"ed",  x"94",  x"9e",  x"74",  x"8a", -- 29B0
         x"80",  x"fe",  x"0a",  x"20",  x"05",  x"cd",  x"2b",  x"12", -- 29B8
         x"df",  x"db",  x"cc",  x"0f",  x"df",  x"c0",  x"cf",  x"27", -- 29C0
         x"df",  x"9b",  x"00",  x"32",  x"df",  x"18",  x"e7",  x"fe", -- 29C8
         x"0d",  x"14",  x"c0",  x"3e",  x"09",  x"30",  x"23",  x"6a", -- 29D0
         x"7e",  x"49",  x"f6",  x"d1",  x"b6",  x"20",  x"a1",  x"1b", -- 29D8
         x"30",  x"c3",  x"d4",  x"06",  x"fe",  x"ba",  x"07",  x"02", -- 29E0
         x"a7",  x"2a",  x"b6",  x"2f",  x"37",  x"e8",  x"19",  x"08", -- 29E8
         x"28",  x"44",  x"c8",  x"80",  x"28",  x"2a",  x"fe",  x"1f", -- 29F0
         x"28",  x"47",  x"fe",  x"00",  x"19",  x"ca",  x"c5",  x"df", -- 29F8
         x"fe",  x"18",  x"ca",  x"cf",  x"c6",  x"04",  x"02",  x"ca", -- 2A00
         x"db",  x"04",  x"1a",  x"07",  x"28",  x"48",  x"fe",  x"0b", -- 2A08
         x"c8",  x"5a",  x"bc",  x"02",  x"01",  x"02",  x"f8",  x"0a", -- 2A10
         x"05",  x"3f",  x"4a",  x"25",  x"c9",  x"77",  x"4f",  x"dc", -- 2A18
         x"9e",  x"ab",  x"03",  x"a3",  x"e5",  x"3a",  x"28",  x"07", -- 2A20
         x"7e",  x"84",  x"0a",  x"d2",  x"03",  x"a2",  x"c6",  x"60", -- 2A28
         x"f0",  x"15",  x"6e",  x"18",  x"df",  x"e5",  x"23",  x"a0", -- 2A30
         x"9a",  x"f4",  x"fb",  x"c6",  x"d1",  x"73",  x"af",  x"cb", -- 2A38
         x"e3",  x"2d",  x"17",  x"78",  x"20",  x"f7",  x"6b",  x"ec", -- 2A40
         x"0e",  x"b0",  x"25",  x"34",  x"2a",  x"20",  x"0c",  x"15", -- 2A48
         x"af",  x"11",  x"33",  x"3b",  x"67",  x"d1",  x"e2",  x"f9", -- 2A50
         x"c4",  x"02",  x"0b",  x"7e",  x"0c",  x"28",  x"4b",  x"20", -- 2A58
         x"4b",  x"c9",  x"4a",  x"4c",  x"c1",  x"b2",  x"89",  x"bc", -- 2A60
         x"00",  x"18",  x"90",  x"cd",  x"c5",  x"ff",  x"58",  x"09", -- 2A68
         x"bc",  x"eb",  x"6f",  x"f2",  x"45",  x"e1",  x"f6",  x"61", -- 2A70
         x"10",  x"fe",  x"00",  x"c9",  x"1e",  x"ff",  x"c3",  x"0e", -- 2A78
         x"27",  x"e0",  x"ff",  x"00",  x"ce",  x"0c",  x"d2",  x"e0", -- 2A80
         x"9c",  x"71",  x"02",  x"57",  x"e1",  x"11",  x"80",  x"04", -- 2A88
         x"00",  x"e6",  x"c9",  x"4e",  x"4b",  x"45",  x"59",  x"00", -- 2A90
         x"24",  x"ca",  x"4f",  x"59",  x"53",  x"54",  x"d3",  x"54", -- 2A98
         x"07",  x"52",  x"49",  x"4e",  x"47",  x"24",  x"11",  x"80", -- 2AA0
         x"0a",  x"52",  x"d2",  x"45",  x"4e",  x"55",  x"4d",  x"c4", -- 2AA8
         x"00",  x"45",  x"4c",  x"45",  x"54",  x"45",  x"d0",  x"41", -- 2AB0
         x"55",  x"01",  x"53",  x"45",  x"c2",  x"45",  x"45",  x"50", -- 2AB8
         x"d7",  x"80",  x"1d",  x"44",  x"4f",  x"57",  x"c2",  x"4f", -- 2AC0
         x"52",  x"44",  x"2b",  x"45",  x"52",  x"36",  x"17",  x"63", -- 2AC8
         x"50",  x"07",  x"c1",  x"54",  x"d0",  x"1c",  x"30",  x"54", -- 2AD0
         x"cc",  x"19",  x"45",  x"c3",  x"49",  x"52",  x"6f",  x"43", -- 2AD8
         x"2e",  x"a1",  x"15",  x"0b",  x"cc",  x"0f",  x"41",  x"42", -- 2AE0
         x"3a",  x"d3",  x"49",  x"18",  x"5a",  x"45",  x"da",  x"21", -- 2AE8
         x"4f",  x"c8",  x"4f",  x"6c",  x"4d",  x"16",  x"c7",  x"1b", -- 2AF0
         x"53",  x"d3",  x"3d",  x"43",  x"41",  x"20",  x"04",  x"52", -- 2AF8
         x"8a",  x"4a",  x"4e",  x"d0",  x"4f",  x"25",  x"02",  x"d8", -- 2B00
         x"50",  x"4f",  x"53",  x"a1",  x"d9",  x"80",  x"04",  x"80", -- 2B08
         x"19",  x"e4",  x"f5",  x"e4",  x"3c",  x"0c",  x"e4",  x"c1", -- 2B10
         x"e4",  x"f8",  x"b6",  x"00",  x"e5",  x"a7",  x"e3",  x"34", -- 2B18
         x"e4",  x"b5",  x"00",  x"e1",  x"79",  x"e1",  x"7d",  x"e1", -- 2B20
         x"7e",  x"e1",  x"17",  x"00",  x"e5",  x"d6",  x"a7",  x"d9", -- 2B28
         x"a7",  x"dc",  x"a7",  x"4a",  x"06",  x"ca",  x"df",  x"a7", -- 2B30
         x"e2",  x"a7",  x"1a",  x"e8",  x"28",  x"a7",  x"eb",  x"0b", -- 2B38
         x"ee",  x"a7",  x"01",  x"f1",  x"a7",  x"f4",  x"a7",  x"f7", -- 2B40
         x"a7",  x"fa",  x"41",  x"0b",  x"fd",  x"a7",  x"78",  x"d6", -- 2B48
         x"b2",  x"e5",  x"6d",  x"99",  x"e9",  x"07",  x"80",  x"f1", -- 2B50
         x"e5",  x"fe",  x"16",  x"0d",  x"30",  x"62",  x"07",  x"4f", -- 2B58
         x"f9",  x"80",  x"eb",  x"21",  x"9e",  x"e0",  x"09",  x"4e", -- 2B60
         x"06",  x"23",  x"46",  x"c5",  x"eb",  x"c3",  x"8b",  x"99", -- 2B68
         x"d5",  x"64",  x"ec",  x"fe",  x"06",  x"e2",  x"d0",  x"fe", -- 2B70
         x"e1",  x"ca",  x"4e",  x"3a",  x"6e",  x"fd",  x"cb",  x"20", -- 2B78
         x"69",  x"3f",  x"bd",  x"be",  x"06",  x"3a",  x"fd",  x"51", -- 2B80
         x"f5",  x"19",  x"28",  x"0d",  x"48",  x"ad",  x"cd",  x"f0", -- 2B88
         x"69",  x"0a",  x"3b",  x"28",  x"35",  x"18",  x"5f",  x"25", -- 2B90
         x"0c",  x"78",  x"63",  x"0c",  x"28",  x"cd",  x"d6",  x"d2", -- 2B98
         x"21",  x"e0",  x"20",  x"13",  x"2d",  x"1e",  x"c6",  x"ab", -- 2BA0
         x"b8",  x"c3",  x"cb",  x"f1",  x"32",  x"35",  x"70",  x"c1", -- 2BA8
         x"97",  x"e2",  x"1a",  x"d3",  x"b8",  x"c3",  x"e0",  x"48", -- 2BB0
         x"06",  x"67",  x"56",  x"c9",  x"20",  x"90",  x"80",  x"79", -- 2BB8
         x"d6",  x"3e",  x"38",  x"e8",  x"3b",  x"fe",  x"07",  x"8a", -- 2BC0
         x"b0",  x"84",  x"18",  x"32",  x"38",  x"dd",  x"40",  x"30", -- 2BC8
         x"d9",  x"eb",  x"05",  x"01",  x"96",  x"e0",  x"e1",  x"6f", -- 2BD0
         x"01",  x"86",  x"66",  x"69",  x"de",  x"b1",  x"34",  x"01", -- 2BD8
         x"0e",  x"18",  x"02",  x"f6",  x"af",  x"b3",  x"0c",  x"21", -- 2BE0
         x"d4",  x"ab",  x"cc",  x"38",  x"6e",  x"af",  x"01",  x"30", -- 2BE8
         x"6a",  x"3d",  x"4f",  x"f1",  x"90",  x"ad",  x"0b",  x"cb", -- 2BF0
         x"21",  x"b1",  x"01",  x"3d",  x"28",  x"17",  x"94",  x"04", -- 2BF8
         x"41",  x"b7",  x"94",  x"06",  x"28",  x"0a",  x"d7",  x"ca", -- 2C00
         x"b0",  x"66",  x"00",  x"32",  x"28",  x"00",  x"c9",  x"e6", -- 2C08
         x"70",  x"18",  x"f4",  x"00",  x"79",  x"d3",  x"88",  x"c9", -- 2C10
         x"0e",  x"1d",  x"cd",  x"05",  x"54",  x"00",  x"f7",  x"03", -- 2C18
         x"28",  x"2d",  x"cd",  x"f7",  x"e7",  x"42",  x"9f",  x"03", -- 2C20
         x"4a",  x"00",  x"3c",  x"3c",  x"57",  x"fe",  x"2a",  x"30", -- 2C28
         x"20",  x"f1",  x"3d",  x"5f",  x"f1",  x"09",  x"9c",  x"1b", -- 2C30
         x"1a",  x"9f",  x"00",  x"f1",  x"4f",  x"3c",  x"b8",  x"30", -- 2C38
         x"10",  x"7b",  x"1b",  x"3c",  x"ba",  x"30",  x"b6",  x"b7", -- 2C40
         x"06",  x"f3",  x"78",  x"19",  x"a2",  x"29",  x"00",  x"c3", -- 2C48
         x"e6",  x"e7",  x"c3",  x"4b",  x"e1",  x"01",  x"0a",  x"00", -- 2C50
         x"00",  x"c5",  x"50",  x"58",  x"28",  x"27",  x"fe",  x"2c", -- 2C58
         x"3d",  x"28",  x"09",  x"98",  x"3b",  x"86",  x"c9",  x"9f", -- 2C60
         x"14",  x"d1",  x"28",  x"1a",  x"e2",  x"15",  x"0a",  x"b2", -- 2C68
         x"a4",  x"f1",  x"ac",  x"08",  x"14",  x"c2",  x"44",  x"00", -- 2C70
         x"e1",  x"7a",  x"b3",  x"28",  x"d1",  x"eb",  x"e3",  x"eb", -- 2C78
         x"dc",  x"a7",  x"cd",  x"bb",  x"24",  x"c4",  x"d1",  x"05", -- 2C80
         x"e9",  x"95",  x"d1",  x"48",  x"91",  x"eb",  x"1f",  x"38", -- 2C88
         x"ba",  x"d1",  x"d5",  x"86",  x"d5",  x"f5",  x"18",  x"0e", -- 2C90
         x"e9",  x"26",  x"f4",  x"eb",  x"ec",  x"a5",  x"f9",  x"ff", -- 2C98
         x"00",  x"14",  x"e1",  x"38",  x"e9",  x"d5",  x"5e",  x"23", -- 2CA0
         x"56",  x"db",  x"33",  x"eb",  x"4c",  x"07",  x"90",  x"60", -- 2CA8
         x"b6",  x"2b",  x"eb",  x"20",  x"ed",  x"b4",  x"0e",  x"b8", -- 2CB0
         x"ed",  x"27",  x"c3",  x"af",  x"d8",  x"b0",  x"e2",  x"af", -- 2CB8
         x"56",  x"3c",  x"04",  x"dd",  x"f2",  x"e9",  x"43",  x"07", -- 2CC0
         x"f1",  x"71",  x"2a",  x"f0",  x"a5",  x"5e",  x"23",  x"50", -- 2CC8
         x"a9",  x"eb",  x"09",  x"eb",  x"dc",  x"87",  x"eb",  x"3d", -- 2CD0
         x"a7",  x"23",  x"01",  x"94",  x"60",  x"c5",  x"3e",  x"02", -- 2CD8
         x"32",  x"4e",  x"00",  x"03",  x"2a",  x"5f",  x"03",  x"2b", -- 2CE0
         x"c5",  x"c5",  x"23",  x"34",  x"c1",  x"c1",  x"f0",  x"90", -- 2CE8
         x"2b",  x"c8",  x"c5",  x"54",  x"d5",  x"af",  x"e3",  x"df", -- 2CF0
         x"88",  x"a6",  x"eb",  x"4f",  x"3a",  x"c3",  x"1e",  x"b7", -- 2CF8
         x"79",  x"28",  x"5f",  x"b0",  x"61",  x"20",  x"ee",  x"e5", -- 2D00
         x"ad",  x"bf",  x"56",  x"1e",  x"10",  x"b5",  x"2d",  x"7e", -- 2D08
         x"02",  x"0e",  x"fa",  x"4d",  x"8f",  x"ed",  x"78",  x"a0", -- 2D10
         x"01",  x"84",  x"78",  x"f1",  x"18",  x"c0",  x"b3",  x"eb", -- 2D18
         x"13",  x"aa",  x"98",  x"e7",  x"d5",  x"42",  x"6e",  x"e1", -- 2D20
         x"67",  x"c5",  x"f9",  x"be",  x"78",  x"98",  x"80",  x"c5", -- 2D28
         x"af",  x"06",  x"98",  x"cd",  x"ae",  x"fc",  x"95",  x"34", -- 2D30
         x"d8",  x"f5",  x"0d",  x"ac",  x"33",  x"eb",  x"2b",  x"4f", -- 2D38
         x"aa",  x"23",  x"1b",  x"c8",  x"94",  x"09",  x"54",  x"2f", -- 2D40
         x"5d",  x"13",  x"9b",  x"0f",  x"1b",  x"2b",  x"b5",  x"58", -- 2D48
         x"e1",  x"40",  x"c1",  x"18",  x"e3",  x"00",  x"fe",  x"88", -- 2D50
         x"28",  x"19",  x"fe",  x"8c",  x"28",  x"15",  x"03",  x"fe", -- 2D58
         x"8b",  x"28",  x"11",  x"fe",  x"d4",  x"ab",  x"03",  x"fe", -- 2D60
         x"da",  x"ae",  x"13",  x"fe",  x"d3",  x"d3",  x"50",  x"fe", -- 2D68
         x"a9",  x"c2",  x"b2",  x"75",  x"e2",  x"d2",  x"dd",  x"c6", -- 2D70
         x"06",  x"cc",  x"f5",  x"05",  x"14",  x"7e",  x"0b",  x"c6", -- 2D78
         x"f1",  x"6c",  x"58",  x"eb",  x"0d",  x"23",  x"71",  x"23", -- 2D80
         x"79",  x"70",  x"d7",  x"f2",  x"1d",  x"78",  x"6e",  x"77", -- 2D88
         x"f6",  x"c1",  x"0a",  x"62",  x"6b",  x"1b",  x"1a",  x"20", -- 2D90
         x"07",  x"10",  x"fe",  x"3a",  x"30",  x"0c",  x"a7",  x"83", -- 2D98
         x"2b",  x"e3",  x"f5",  x"c6",  x"0c",  x"87",  x"3a",  x"97", -- 2DA0
         x"49",  x"e7",  x"6f",  x"cb",  x"00",  x"72",  x"95",  x"71", -- 2DA8
         x"3e",  x"0d",  x"a6",  x"8b",  x"d1",  x"b3",  x"c5",  x"e3", -- 2DB0
         x"56",  x"14",  x"07",  x"29",  x"d5",  x"d4",  x"5f",  x"93", -- 2DB8
         x"51",  x"18",  x"51",  x"9f",  x"ec",  x"07",  x"20",  x"11", -- 2DC0
         x"cd",  x"f3",  x"a9",  x"6a",  x"fb",  x"89",  x"80",  x"07", -- 2DC8
         x"fe",  x"1e",  x"20",  x"54",  x"f3",  x"c2",  x"66",  x"ea", -- 2DD0
         x"5e",  x"50",  x"c9",  x"94",  x"e3",  x"fc",  x"90",  x"d8", -- 2DD8
         x"dd",  x"21",  x"0b",  x"00",  x"e4",  x"3e",  x"05",  x"0e", -- 2DE0
         x"8d",  x"06",  x"0a",  x"dd",  x"3c",  x"86",  x"00",  x"fc", -- 2DE8
         x"c4",  x"94",  x"f6",  x"3d",  x"cf",  x"85",  x"9c",  x"5c", -- 2DF0
         x"7e",  x"eb",  x"28",  x"55",  x"1b",  x"6e",  x"ba",  x"39", -- 2DF8
         x"08",  x"35",  x"bb",  x"0c",  x"3d",  x"08",  x"d1",  x"0a", -- 2E00
         x"c1",  x"f1",  x"18",  x"cf",  x"3e",  x"ae",  x"07",  x"f6", -- 2E08
         x"dc",  x"c3",  x"f0",  x"7c",  x"c3",  x"53",  x"1f",  x"49", -- 2E10
         x"43",  x"20",  x"00",  x"e7",  x"02",  x"8c",  x"c0",  x"57", -- 2E18
         x"6f",  x"0c",  x"9d",  x"16",  x"e5",  x"33",  x"0f",  x"d1", -- 2E20
         x"a5",  x"cd",  x"dd",  x"a7",  x"01",  x"2b",  x"2a",  x"c2", -- 2E28
         x"03",  x"77",  x"c3",  x"a9",  x"c5",  x"9f",  x"6e",  x"0d", -- 2E30
         x"cb",  x"0e",  x"14",  x"02",  x"1e",  x"07",  x"80",  x"9e", -- 2E38
         x"7e",  x"84",  x"a9",  x"28",  x"0c",  x"f8",  x"8e",  x"e4", -- 2E40
         x"cc",  x"03",  x"db",  x"c8",  x"da",  x"1f",  x"44",  x"83", -- 2E48
         x"00",  x"d5",  x"4f",  x"af",  x"b9",  x"28",  x"0c",  x"b8", -- 2E50
         x"cc",  x"69",  x"79",  x"05",  x"a5",  x"46",  x"81",  x"38", -- 2E58
         x"29",  x"8b",  x"06",  x"47",  x"0e",  x"aa",  x"8f",  x"e1", -- 2E60
         x"6b",  x"f6",  x"26",  x"7e",  x"f9",  x"26",  x"e3",  x"7c", -- 2E68
         x"02",  x"6f",  x"32",  x"24",  x"25",  x"80",  x"63",  x"28", -- 2E70
         x"40",  x"f2",  x"d2",  x"c1",  x"ef",  x"27",  x"f4",  x"03", -- 2E78
         x"94",  x"5e",  x"02",  x"d3",  x"5a",  x"1e",  x"5f",  x"1c", -- 2E80
         x"86",  x"fd",  x"c8",  x"8b",  x"77",  x"30",  x"d3",  x"23", -- 2E88
         x"cf",  x"2c",  x"9b",  x"31",  x"ba",  x"06",  x"2b",  x"0d", -- 2E90
         x"c5",  x"0c",  x"13",  x"48",  x"11",  x"31",  x"23",  x"0d", -- 2E98
         x"50",  x"1a",  x"be",  x"28",  x"63",  x"2d",  x"18",  x"2c", -- 2EA0
         x"e1",  x"36",  x"79",  x"31",  x"4a",  x"dc",  x"30",  x"a7", -- 2EA8
         x"dd",  x"12",  x"7d",  x"18",  x"2a",  x"06",  x"84",  x"80", -- 2EB0
         x"1a",  x"89",  x"5a",  x"bc",  x"4c",  x"88",  x"1a",  x"c9", -- 2EB8
         x"33",  x"4f",  x"03",  x"6d",  x"47",  x"ef",  x"2f",  x"df", -- 2EC0
         x"29",  x"35",  x"b8",  x"8d",  x"3d",  x"20",  x"f9",  x"af", -- 2EC8
         x"35",  x"11",  x"89",  x"b3",  x"d5",  x"18",  x"88",  x"e0", -- 2ED0
         x"e3",  x"18",  x"f6",  x"c3",  x"8f",  x"66",  x"b0",  x"0d", -- 2ED8
         x"cd",  x"24",  x"d4",  x"a7",  x"31",  x"28",  x"45",  x"93", -- 2EE0
         x"0a",  x"30",  x"41",  x"0e",  x"06",  x"d0",  x"03",  x"38", -- 2EE8
         x"3a",  x"8a",  x"60",  x"28",  x"01",  x"48",  x"79",  x"1b", -- 2EF0
         x"c3",  x"c0",  x"d0",  x"97",  x"cb",  x"88",  x"fa",  x"06", -- 2EF8
         x"20",  x"de",  x"83",  x"e6",  x"64",  x"e2",  x"5b",  x"60", -- 2F00
         x"b6",  x"fd",  x"63",  x"f1",  x"62",  x"e5",  x"47",  x"78", -- 2F08
         x"fb",  x"ae",  x"e4",  x"bf",  x"d6",  x"14",  x"28",  x"38", -- 2F10
         x"03",  x"d2",  x"a1",  x"2e",  x"00",  x"65",  x"55",  x"8b", -- 2F18
         x"e2",  x"04",  x"ae",  x"00",  x"03",  x"19",  x"10",  x"fd", -- 2F20
         x"52",  x"59",  x"ea",  x"99",  x"ec",  x"19",  x"df",  x"65", -- 2F28
         x"9a",  x"e6",  x"85",  x"c6",  x"40",  x"fe",  x"d5",  x"38", -- 2F30
         x"09",  x"3a",  x"6f",  x"fc",  x"ea",  x"8b",  x"1a",  x"cd", -- 2F38
         x"06",  x"e0",  x"e4",  x"03",  x"3a",  x"ae",  x"bd",  x"4a", -- 2F40
         x"d4",  x"ad",  x"80",  x"07",  x"cd",  x"8a",  x"d1",  x"9f", -- 2F48
         x"40",  x"2a",  x"e5",  x"03",  x"34",  x"cd",  x"03",  x"fe", -- 2F50
         x"d2",  x"cd",  x"ee",  x"d6",  x"e1",  x"b6",  x"f2",  x"fd", -- 2F58
         x"e1",  x"98",  x"f5",  x"57",  x"1c",  x"00",  x"1d",  x"28", -- 2F60
         x"13",  x"0a",  x"cd",  x"bf",  x"e5",  x"30",  x"f8",  x"e7", -- 2F68
         x"77",  x"00",  x"32",  x"fd",  x"72",  x"e0",  x"1e",  x"23", -- 2F70
         x"fd",  x"23",  x"d7",  x"2c",  x"ea",  x"87",  x"db",  x"02", -- 2F78
         x"f1",  x"d0",  x"eb",  x"01",  x"fd",  x"e5",  x"dd",  x"e5", -- 2F80
         x"18",  x"a7",  x"40",  x"04",  x"e1",  x"d5",  x"11",  x"c0", -- 2F88
         x"ef",  x"a1",  x"8b",  x"c5",  x"92",  x"c9",  x"6c",  x"bd", -- 2F90
         x"ca",  x"26",  x"42",  x"c4",  x"bd",  x"61",  x"e1",  x"c0", -- 2F98
         x"eb",  x"68",  x"9e",  x"d2",  x"e9",  x"b6",  x"d1",  x"9e", -- 2FA0
         x"82",  x"38",  x"c4",  x"00",  x"30",  x"f5",  x"c1",  x"c3", -- 2FA8
         x"50",  x"c4",  x"47",  x"e5",  x"0f",  x"2a",  x"b0",  x"e0", -- 2FB0
         x"3e",  x"aa",  x"bf",  x"bd",  x"36",  x"c8",  x"c3",  x"de", -- 2FB8
         x"0c",  x"ff",  x"cb",  x"6b",  x"c2",  x"eb",  x"9e",  x"22", -- 2FC0
         x"62",  x"92",  x"40",  x"21",  x"1e",  x"e6",  x"e5",  x"7b", -- 2FC8
         x"dd",  x"eb",  x"17",  x"52",  x"ae",  x"21",  x"1b",  x"42", -- 2FD0
         x"e6",  x"09",  x"be",  x"06",  x"66",  x"6f",  x"e9",  x"c1", -- 2FD8
         x"53",  x"0a",  x"00",  x"0d",  x"56",  x"65",  x"72",  x"69", -- 2FE0
         x"66",  x"79",  x"20",  x"e4",  x"81",  x"59",  x"29",  x"00", -- 2FE8
         x"2f",  x"4e",  x"29",  x"3f",  x"3a",  x"00",  x"0a",  x"52", -- 2FF0
         x"00",  x"65",  x"77",  x"69",  x"6e",  x"64",  x"20",  x"3c", -- 2FF8
         x"3d",  x"60",  x"3d",  x"1d",  x"00",  x"52",  x"e6",  x"72", -- 3000
         x"e6",  x"01",  x"34",  x"e7",  x"85",  x"e6",  x"82",  x"dc", -- 3008
         x"6e",  x"5f",  x"03",  x"01",  x"d8",  x"f9",  x"af",  x"14", -- 3010
         x"0e",  x"0b",  x"ce",  x"3a",  x"d5",  x"83",  x"0e",  x"cb", -- 3018
         x"bb",  x"18",  x"0a",  x"a0",  x"7a",  x"0b",  x"29",  x"0e", -- 3020
         x"01",  x"04",  x"57",  x"c3",  x"b8",  x"05",  x"f4",  x"8c", -- 3028
         x"bd",  x"ca",  x"d5",  x"5a",  x"0c",  x"60",  x"d1",  x"1b", -- 3030
         x"c9",  x"16",  x"0a",  x"18",  x"f1",  x"00",  x"16",  x"0d", -- 3038
         x"18",  x"ed",  x"d5",  x"cb",  x"5b",  x"28",  x"0a",  x"22", -- 3040
         x"d5",  x"0e",  x"0f",  x"16",  x"7d",  x"16",  x"9b",  x"86", -- 3048
         x"4e",  x"01",  x"0b",  x"00",  x"2a",  x"92",  x"19",  x"85", -- 3050
         x"80",  x"7e",  x"32",  x"75",  x"00",  x"11",  x"80",  x"00", -- 3058
         x"a5",  x"ac",  x"03",  x"21",  x"6e",  x"00",  x"36",  x"0b", -- 3060
         x"21",  x"0a",  x"74",  x"3a",  x"07",  x"9f",  x"07",  x"09", -- 3068
         x"72",  x"b1",  x"59",  x"08",  x"cb",  x"73",  x"a5",  x"d3", -- 3070
         x"01",  x"0f",  x"fe",  x"80",  x"c2",  x"7d",  x"e7",  x"3a", -- 3078
         x"e2",  x"28",  x"e3",  x"20",  x"4a",  x"1a",  x"21",  x"47", -- 3080
         x"50",  x"56",  x"43",  x"23",  x"10",  x"f9",  x"61",  x"21", -- 3088
         x"d9",  x"f8",  x"2b",  x"79",  x"9b",  x"bd",  x"42",  x"a6", -- 3090
         x"a3",  x"19",  x"22",  x"1b",  x"0c",  x"53",  x"15",  x"62", -- 3098
         x"af",  x"3b",  x"97",  x"66",  x"40",  x"36",  x"28",  x"74", -- 30A0
         x"0c",  x"5a",  x"62",  x"21",  x"1f",  x"e6",  x"cd",  x"62", -- 30A8
         x"02",  x"10",  x"d6",  x"ea",  x"02",  x"81",  x"01",  x"e6", -- 30B0
         x"fe",  x"4e",  x"28",  x"66",  x"11",  x"34",  x"72",  x"12", -- 30B8
         x"9e",  x"0f",  x"3a",  x"6b",  x"51",  x"26",  x"6c",  x"e4", -- 30C0
         x"af",  x"cd",  x"83",  x"31",  x"e7",  x"c1",  x"55",  x"18", -- 30C8
         x"49",  x"d5",  x"4a",  x"79",  x"44",  x"b2",  x"05",  x"1b", -- 30D0
         x"6b",  x"1f",  x"a0",  x"54",  x"19",  x"18",  x"cd",  x"30", -- 30D8
         x"9d",  x"e7",  x"a4",  x"0b",  x"8b",  x"00",  x"56",  x"d5", -- 30E0
         x"a9",  x"01",  x"0c",  x"18",  x"1c",  x"12",  x"ab",  x"0e", -- 30E8
         x"d1",  x"13",  x"c3",  x"ad",  x"a6",  x"02",  x"20",  x"10", -- 30F0
         x"ae",  x"27",  x"7c",  x"41",  x"9d",  x"a6",  x"89",  x"50", -- 30F8
         x"1d",  x"83",  x"89",  x"cb",  x"9b",  x"c9",  x"81",  x"9a", -- 3100
         x"14",  x"43",  x"14",  x"d0",  x"cd",  x"67",  x"7e",  x"d1", -- 3108
         x"eb",  x"ed",  x"8c",  x"1c",  x"20",  x"f5",  x"c3",  x"ca", -- 3110
         x"68",  x"19",  x"06",  x"0b",  x"98",  x"cc",  x"31",  x"90", -- 3118
         x"cc",  x"22",  x"0c",  x"09",  x"0e",  x"11",  x"8a",  x"68", -- 3120
         x"00",  x"d3",  x"1b",  x"00",  x"20",  x"04",  x"2b",  x"10", -- 3128
         x"f8",  x"c9",  x"d6",  x"04",  x"01",  x"be",  x"20",  x"d8", -- 3130
         x"3e",  x"ff",  x"32",  x"5e",  x"99",  x"99",  x"f0",  x"ff", -- 3138
         x"0d",  x"ee",  x"00",  x"e1",  x"3d",  x"c4",  x"c5",  x"43", -- 3140
         x"3b",  x"02",  x"00",  x"51",  x"14",  x"1c",  x"0e",  x"12", -- 3148
         x"46",  x"ba",  x"b4",  x"c8",  x"cc",  x"a6",  x"f1",  x"c9", -- 3150
         x"80",  x"00",  x"40",  x"c3",  x"02",  x"0c",  x"80",  x"4d", -- 3158
         x"4f",  x"4e",  x"20",  x"c0",  x"00",  x"00",  x"31",  x"c0", -- 3160
         x"eb",  x"cd",  x"cb",  x"00",  x"86",  x"cd",  x"d7",  x"80", -- 3168
         x"c3",  x"03",  x"f0",  x"00",  x"98",  x"00",  x"3e",  x"02", -- 3170
         x"00",  x"cf",  x"c9",  x"3e",  x"00",  x"cf",  x"76",  x"18", -- 3178
         x"fd",  x"00",  x"c1",  x"e1",  x"31",  x"00",  x"02",  x"e9", -- 3180
         x"c9",  x"2a",  x"c0",  x"00",  x"20",  x"4d",  x"6f",  x"6e", -- 3188
         x"69",  x"74",  x"00",  x"6f",  x"72",  x"20",  x"56",  x"30", -- 3190
         x"2e",  x"30",  x"30",  x"28",  x"31",  x"20",  x"12",  x"0a", -- 3198
         x"00",  x"18",  x"fd",  x"21",  x"02",  x"03",  x"39",  x"fd", -- 31A0
         x"66",  x"00",  x"00",  x"7c",  x"57",  x"d6",  x"30",  x"38", -- 31A8
         x"0a",  x"3e",  x"00",  x"39",  x"94",  x"38",  x"05",  x"7a", -- 31B0
         x"c6",  x"d0",  x"6f",  x"0a",  x"c9",  x"7c",  x"d6",  x"41", -- 31B8
         x"0e",  x"48",  x"46",  x"0e",  x"c9",  x"b5",  x"0e",  x"61", -- 31C0
         x"24",  x"0e",  x"66",  x"0e",  x"66",  x"a9",  x"0e",  x"2e", -- 31C8
         x"ff",  x"5e",  x"3e",  x"03",  x"f5",  x"33",  x"cd",  x"c2", -- 31D0
         x"83",  x"33",  x"60",  x"06",  x"e5",  x"c5",  x"2e",  x"00", -- 31D8
         x"e5",  x"0b",  x"0f",  x"27",  x"84",  x"33",  x"4d",  x"98", -- 31E0
         x"0e",  x"3e",  x"0a",  x"94",  x"22",  x"c9",  x"dd",  x"18", -- 31E8
         x"e5",  x"dd",  x"21",  x"94",  x"00",  x"dd",  x"39",  x"dd", -- 31F0
         x"6e",  x"04",  x"dd",  x"66",  x"00",  x"05",  x"e5",  x"56", -- 31F8
         x"23",  x"5e",  x"e1",  x"7a",  x"e6",  x"00",  x"03",  x"28", -- 3200
         x"04",  x"d6",  x"03",  x"20",  x"02",  x"cb",  x"00",  x"fb", -- 3208
         x"cb",  x"3b",  x"cb",  x"1a",  x"72",  x"23",  x"73",  x"22", -- 3210
         x"dd",  x"e1",  x"00",  x"27",  x"21",  x"ee",  x"ff",  x"39", -- 3218
         x"f9",  x"dd",  x"1b",  x"36",  x"f6",  x"d2",  x"03",  x"f7", -- 3220
         x"31",  x"29",  x"36",  x"f4",  x"07",  x"f5",  x"4c",  x"07", -- 3228
         x"f2",  x"1a",  x"36",  x"f3",  x"a3",  x"03",  x"f1",  x"01", -- 3230
         x"03",  x"52",  x"f0",  x"07",  x"ef",  x"94",  x"03",  x"ee", -- 3238
         x"03",  x"f8",  x"c0",  x"ef",  x"03",  x"d3",  x"00",  x"02", -- 3240
         x"21",  x"31",  x"80",  x"e5",  x"cd",  x"d8",  x"83",  x"00", -- 3248
         x"f1",  x"cd",  x"cf",  x"83",  x"dd",  x"75",  x"ff",  x"7d", -- 3250
         x"18",  x"b7",  x"28",  x"f6",  x"6b",  x"ff",  x"7c",  x"fe", -- 3258
         x"02",  x"0a",  x"ca",  x"ca",  x"81",  x"fe",  x"0d",  x"c6", -- 3260
         x"04",  x"3a",  x"ca",  x"e2",  x"04",  x"67",  x"00",  x"28", -- 3268
         x"72",  x"fe",  x"6b",  x"ca",  x"bc",  x"81",  x"d6",  x"0c", -- 3270
         x"6d",  x"ca",  x"e9",  x"81",  x"1d",  x"70",  x"28",  x"00", -- 3278
         x"55",  x"d6",  x"72",  x"28",  x"3f",  x"dd",  x"7e",  x"f2", -- 3280
         x"66",  x"c6",  x"54",  x"77",  x"fd",  x"07",  x"f3",  x"66", -- 3288
         x"ce",  x"50",  x"77",  x"fe",  x"18",  x"73",  x"01",  x"28", -- 3290
         x"0f",  x"d6",  x"74",  x"c2",  x"9b",  x"82",  x"4b",  x"65", -- 3298
         x"01",  x"71",  x"30",  x"18",  x"a8",  x"bc",  x"67",  x"f2", -- 32A0
         x"50",  x"f3",  x"66",  x"22",  x"b3",  x"25",  x"77",  x"09", -- 32A8
         x"7e",  x"fe",  x"05",  x"4a",  x"f3",  x"e6",  x"01",  x"18", -- 32B0
         x"8d",  x"3e",  x"05",  x"cb",  x"7e",  x"1e",  x"80",  x"81", -- 32B8
         x"2a",  x"80",  x"f1",  x"13",  x"c3",  x"1c",  x"81",  x"a4", -- 32C0
         x"0d",  x"83",  x"0d",  x"ba",  x"1f",  x"86",  x"21",  x"c3", -- 32C8
         x"89",  x"f0",  x"14",  x"1a",  x"18",  x"5c",  x"86",  x"1a", -- 32D0
         x"a0",  x"c1",  x"ef",  x"90",  x"c5",  x"34",  x"54",  x"ff", -- 32D8
         x"a3",  x"b0",  x"2f",  x"17",  x"2f",  x"b5",  x"06",  x"f3", -- 32E0
         x"07",  x"fb",  x"0c",  x"1b",  x"fc",  x"00",  x"11",  x"97", -- 32E8
         x"40",  x"7a",  x"d6",  x"80",  x"30",  x"12",  x"21",  x"0d", -- 32F0
         x"08",  x"00",  x"39",  x"d5",  x"3c",  x"af",  x"b0",  x"57", -- 32F8
         x"d1",  x"2e",  x"f6",  x"12",  x"13",  x"18",  x"44",  x"e9", -- 3300
         x"0e",  x"97",  x"bb",  x"14",  x"20",  x"59",  x"39",  x"21", -- 3308
         x"06",  x"20",  x"25",  x"1f",  x"67",  x"00",  x"56",  x"dd", -- 3310
         x"5e",  x"f4",  x"7a",  x"93",  x"28",  x"38",  x"89",  x"90", -- 3318
         x"01",  x"26",  x"20",  x"e3",  x"24",  x"64",  x"c1",  x"cf", -- 3320
         x"31",  x"aa",  x"25",  x"20",  x"79",  x"d1",  x"11",  x"f4", -- 3328
         x"a4",  x"bb",  x"dd",  x"0c",  x"34",  x"f2",  x"20",  x"a5", -- 3330
         x"04",  x"f3",  x"18",  x"69",  x"a0",  x"1a",  x"fc",  x"cb", -- 3338
         x"e7",  x"0a",  x"4c",  x"fb",  x"08",  x"34",  x"18",  x"fb", -- 3340
         x"20",  x"03",  x"04",  x"fc",  x"21",  x"bd",  x"48",  x"83", -- 3348
         x"fb",  x"22",  x"c3",  x"f2",  x"81",  x"50",  x"c4",  x"01", -- 3350
         x"49",  x"80",  x"33",  x"7d",  x"3c",  x"ca",  x"1c",  x"45", -- 3358
         x"0d",  x"f0",  x"07",  x"06",  x"00",  x"e6",  x"f0",  x"4f", -- 3360
         x"09",  x"94",  x"4c",  x"f0",  x"0d",  x"f1",  x"d6",  x"0c", -- 3368
         x"02",  x"20",  x"04",  x"3e",  x"cd",  x"4c",  x"01",  x"af", -- 3370
         x"be",  x"58",  x"fb",  x"0e",  x"ef",  x"3d",  x"20",  x"6c", -- 3378
         x"5f",  x"05",  x"fb",  x"ab",  x"95",  x"21",  x"28",  x"d1", -- 3380
         x"11",  x"f3",  x"28",  x"fa",  x"c7",  x"33",  x"06",  x"77", -- 3388
         x"fa",  x"09",  x"76",  x"f9",  x"09",  x"d9",  x"0f",  x"7e", -- 3390
         x"0a",  x"e8",  x"11",  x"c3",  x"b7",  x"83",  x"65",  x"3b", -- 3398
         x"04",  x"c2",  x"65",  x"07",  x"8c",  x"58",  x"14",  x"ba", -- 33A0
         x"29",  x"86",  x"2f",  x"f2",  x"31",  x"af",  x"27",  x"f3", -- 33A8
         x"8c",  x"4b",  x"c9",  x"1d",  x"13",  x"ee",  x"9c",  x"d7", -- 33B0
         x"84",  x"28",  x"ee",  x"04",  x"9a",  x"37",  x"5e",  x"ca", -- 33B8
         x"7c",  x"36",  x"19",  x"02",  x"28",  x"58",  x"17",  x"06", -- 33C0
         x"04",  x"28",  x"28",  x"b1",  x"06",  x"05",  x"28",  x"3b", -- 33C8
         x"60",  x"06",  x"06",  x"28",  x"2a",  x"18",  x"45",  x"26", -- 33D0
         x"3e",  x"2a",  x"43",  x"b0",  x"89",  x"4a",  x"f8",  x"f7", -- 33D8
         x"41",  x"ee",  x"03",  x"18",  x"4b",  x"4a",  x"05",  x"05", -- 33E0
         x"13",  x"c1",  x"a3",  x"41",  x"40",  x"09",  x"06",  x"18", -- 33E8
         x"3b",  x"3e",  x"3a",  x"94",  x"27",  x"18",  x"31",  x"c6", -- 33F0
         x"15",  x"f8",  x"b7",  x"20",  x"95",  x"a9",  x"2d",  x"b0", -- 33F8
         x"0f",  x"c3",  x"25",  x"35",  x"f8",  x"d4",  x"1a",  x"2e", -- 3400
         x"45",  x"77",  x"99",  x"a7",  x"3e",  x"2e",  x"38",  x"cc", -- 3408
         x"d9",  x"f2",  x"0d",  x"20",  x"4f",  x"6b",  x"f8",  x"4d", -- 3410
         x"db",  x"00",  x"3a",  x"fb",  x"4a",  x"ae",  x"39",  x"03", -- 3418
         x"7e",  x"d3",  x"00",  x"c9",  x"db",  x"01",  x"5d",  x"1a", -- 3420
         x"02",  x"d3",  x"01",  x"d7",  x"da",  x"cc",  x"82",  x"7e", -- 3428
         x"b7",  x"c8",  x"23",  x"e5",  x"50",  x"2f",  x"e1",  x"18", -- 3430
         x"f2",  x"c9",  x"99",  x"d3",  x"58",  x"56",  x"04",  x"7e", -- 3438
         x"00",  x"d6",  x"1a",  x"0a",  x"30",  x"0a",  x"ff",  x"a6", -- 3440
         x"30",  x"d5",  x"5d",  x"09",  x"37",  x"34",  x"09",  x"92", -- 3448
         x"47",  x"0a",  x"e7",  x"0f",  x"9c",  x"11",  x"eb",  x"11", -- 3450
         x"93",  x"10",  x"ce",  x"0c",  x"42",  x"66",  x"42",  x"01", -- 3458
         x"cd",  x"a7",  x"86",  x"3f",  x"25",  x"00",  x"56",  x"7a", -- 3460
         x"82",  x"0a",  x"05",  x"07",  x"19",  x"36",  x"00",  x"6a", -- 3468
         x"0e",  x"00",  x"b0",  x"e0",  x"06",  x"04",  x"ec",  x"36", -- 3470
         x"20",  x"5d",  x"54",  x"03",  x"13",  x"01",  x"bf",  x"03", -- 3478
         x"ed",  x"b0",  x"0c",  x"44",  x"e8",  x"ca",  x"0c",  x"6e", -- 3480
         x"32",  x"e2",  x"24",  x"18",  x"af",  x"ed",  x"4b",  x"f3", -- 3488
         x"0c",  x"f6",  x"06",  x"69",  x"60",  x"29",  x"29",  x"09", -- 3490
         x"02",  x"29",  x"6c",  x"11",  x"2c",  x"19",  x"f5",  x"c1", -- 3498
         x"04",  x"16",  x"00",  x"d5",  x"01",  x"b3",  x"28",  x"c5", -- 34A0
         x"97",  x"69",  x"9f",  x"e8",  x"db",  x"00",  x"dd",  x"43", -- 34A8
         x"e8",  x"2d",  x"20",  x"4c",  x"2d",  x"f5",  x"f5",  x"8f", -- 34B0
         x"2f",  x"0c",  x"ec",  x"19",  x"33",  x"33",  x"1c",  x"7e", -- 34B8
         x"04",  x"a6",  x"a7",  x"db",  x"05",  x"05",  x"05",  x"ff", -- 34C0
         x"f4",  x"1f",  x"08",  x"ea",  x"6c",  x"b7",  x"76",  x"cb", -- 34C8
         x"c5",  x"e0",  x"fe",  x"68",  x"8f",  x"ff",  x"03",  x"5f", -- 34D0
         x"d6",  x"09",  x"28",  x"20",  x"7b",  x"ae",  x"12",  x"20", -- 34D8
         x"36",  x"a8",  x"2e",  x"ce",  x"11",  x"34",  x"b6",  x"43", -- 34E0
         x"40",  x"18",  x"42",  x"c9",  x"21",  x"57",  x"01",  x"0f", -- 34E8
         x"00",  x"09",  x"6c",  x"1a",  x"ae",  x"86",  x"94",  x"73", -- 34F0
         x"d5",  x"86",  x"20",  x"a6",  x"04",  x"fd",  x"05",  x"18", -- 34F8
         x"a1",  x"3e",  x"17",  x"fd",  x"02",  x"42",  x"fd",  x"96", -- 3500
         x"00",  x"30",  x"05",  x"41",  x"99",  x"22",  x"dd",  x"f9", -- 3508
         x"81",  x"9e",  x"3b",  x"09",  x"3c",  x"45",  x"12",  x"45", -- 3510
         x"aa",  x"de",  x"ff",  x"1c",  x"a2",  x"19",  x"82",  x"31", -- 3518
         x"4f",  x"b5",  x"14",  x"1b",  x"79",  x"47",  x"b8",  x"46", -- 3520
         x"07",  x"78",  x"b8",  x"41",  x"77",  x"eb",  x"18",  x"05", -- 3528
         x"b6",  x"06",  x"37",  x"06",  x"06",  x"bc",  x"03",  x"cb", -- 3530
         x"05",  x"3e",  x"03",  x"0a",  x"04",  x"1e",  x"10",  x"f6", -- 3538
         x"ae",  x"0a",  x"b3",  x"5d",  x"91",  x"05",  x"38",  x"cf", -- 3540
         x"33",  x"42",  x"57",  x"3a",  x"4e",  x"9c",  x"62",  x"fa", -- 3548
         x"23",  x"02",  x"10",  x"fb",  x"c9",  x"01",  x"07",  x"00", -- 3550
         x"c0",  x"cc",  x"02",  x"86",  x"c9",  x"81",  x"c3",  x"db", -- 3558
         x"07",  x"d2",  x"e0",  x"06",  x"f0",  x"c9",  x"cd",  x"4f", -- 3560
         x"84",  x"89",  x"dd",  x"75",  x"c9",  x"81",  x"0a",  x"c1", -- 3568
         x"d1",  x"ed",  x"53",  x"d7",  x"03",  x"b3",  x"91",  x"c0", -- 3570
         x"2d",  x"0c",  x"03",  x"01",  x"67",  x"00",  x"2d",  x"eb", -- 3578
         x"f9",  x"0c",  x"af",  x"32",  x"ab",  x"03",  x"af",  x"85", -- 3580
         x"04",  x"2a",  x"36",  x"00",  x"41",  x"ff",  x"22",  x"b0", -- 3588
         x"03",  x"19",  x"22",  x"56",  x"33",  x"03",  x"3e",  x"14", -- 3590
         x"fc",  x"03",  x"3d",  x"3b",  x"c6",  x"23",  x"bd",  x"00", -- 3598
         x"93",  x"c4",  x"cd",  x"69",  x"c6",  x"c3",  x"54",  x"c8", -- 35A0
         x"42",  x"c9",  x"42",  x"3a",  x"21",  x"c0",  x"01",  x"aa", -- 35A8
         x"2c",  x"1f",  x"12",  x"42",  x"d7",  x"41",  x"5e",  x"41", -- 35B0
         x"21",  x"49",  x"31",  x"67",  x"7d",  x"24",  x"0d",  x"c7", -- 35B8
         x"47",  x"50",  x"ef",  x"dd",  x"4e",  x"08",  x"00",  x"dd", -- 35C0
         x"46",  x"09",  x"51",  x"58",  x"0b",  x"7b",  x"b2",  x"30", -- 35C8
         x"28",  x"07",  x"ea",  x"1a",  x"06",  x"77",  x"23",  x"d6", -- 35D0
         x"4d",  x"19",  x"80",  x"ef",  x"00",  x"01",  x"01",  x"07", -- 35D8
         x"00",  x"78",  x"b1",  x"28",  x"08",  x"55",  x"9a",  x"e4", -- 35E0
         x"ca",  x"81",  x"da",  x"c9",  x"00",  x"00",  x"80",  x"00", -- 35E8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 35F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 35F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3600
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3608
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3610
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3618
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3620
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3628
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3630
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3638
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3640
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3648
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3650
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3658
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3660
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3668
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3670
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3678
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3680
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3688
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3690
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3698
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 36A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 36A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 36B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 36B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 36C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 36C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 36D0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 36D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 36E0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 36E8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 36F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 36F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3700
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3708
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3710
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3718
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3720
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3728
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3730
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3738
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3740
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3748
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3750
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3758
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3760
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3768
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3770
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3778
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3780
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3788
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3790
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3798
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 37A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 37A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 37B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 37B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 37C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 37C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 37D0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 37D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 37E0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 37E8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 37F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 37F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3800
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3808
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3810
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3818
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3820
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3828
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3830
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3838
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3840
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3848
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3850
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3858
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3860
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3868
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3870
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3878
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3880
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3888
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3890
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3898
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 38A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 38A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 38B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 38B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 38C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 38C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 38D0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 38D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 38E0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 38E8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 38F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 38F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3900
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3908
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3910
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3918
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3920
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3928
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3930
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3938
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3940
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3948
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3950
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3958
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3960
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3968
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3970
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3978
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3980
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3988
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3990
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3998
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 39A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 39A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 39B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 39B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 39C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 39C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 39D0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 39D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 39E0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 39E8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 39F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 39F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A10
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A28
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A30
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A38
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A40
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A48
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A50
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A58
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A60
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A68
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A70
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A78
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A80
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A88
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A90
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3AA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3AA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3AB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3AB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3AC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3AC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3AD0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3AD8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3AE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3AE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3AF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3AF8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B10
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B28
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B30
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B38
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B40
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B48
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B50
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B58
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B60
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B68
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B70
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B78
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B80
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B88
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B90
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3BA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3BA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3BB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3BB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3BC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3BC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3BD0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3BD8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3BE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3BE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3BF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3BF8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C10
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C28
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C30
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C38
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C40
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C48
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C50
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C58
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C60
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C68
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C70
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C78
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C80
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C88
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C90
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3CA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3CA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3CB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3CB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3CC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3CC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3CD0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3CD8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3CE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3CE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3CF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3CF8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D10
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D28
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D30
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D38
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D40
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D48
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D50
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D58
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D60
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D68
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D70
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D78
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D80
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D88
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D90
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3DA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3DA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3DB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3DB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3DC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3DC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3DD0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3DD8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3DE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3DE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3DF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3DF8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E10
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E28
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E30
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E38
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E40
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E48
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E50
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E58
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E60
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E68
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E70
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E78
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E80
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E88
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E90
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3EA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3EA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3EB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3EB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3EC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3EC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3ED0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3ED8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3EE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3EE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3EF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3EF8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F10
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F28
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F30
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F38
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F40
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F48
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F50
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F58
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F60
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F68
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F70
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F78
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F80
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F88
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F90
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3FA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3FA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3FB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3FB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3FC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3FC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3FD0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3FD8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3FE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3FE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3FF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00"  -- 3FF8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
