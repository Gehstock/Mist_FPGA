library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity domino_sp_bits is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of domino_sp_bits is
	type rom is array(0 to  32767) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"29",X"99",
		X"00",X"99",X"29",X"11",X"00",X"92",X"24",X"49",X"00",X"72",X"24",X"59",X"00",X"72",X"44",X"69",
		X"00",X"92",X"44",X"11",X"00",X"99",X"24",X"11",X"00",X"00",X"29",X"99",X"00",X"00",X"29",X"90",
		X"00",X"00",X"90",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"C9",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"A9",X"00",X"00",X"CC",X"29",X"00",X"00",X"C9",X"99",X"00",X"00",X"CC",X"9C",X"00",
		X"00",X"9C",X"94",X"00",X"00",X"9C",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"9C",X"00",
		X"00",X"99",X"CC",X"00",X"00",X"44",X"C9",X"00",X"00",X"44",X"99",X"90",X"00",X"49",X"44",X"90",
		X"00",X"99",X"44",X"90",X"00",X"94",X"94",X"90",X"00",X"94",X"44",X"90",X"00",X"94",X"44",X"90",
		X"00",X"99",X"44",X"90",X"00",X"92",X"99",X"90",X"00",X"92",X"22",X"90",X"00",X"99",X"22",X"00",
		X"00",X"91",X"22",X"00",X"00",X"11",X"22",X"00",X"00",X"11",X"22",X"00",X"00",X"11",X"99",X"00",
		X"00",X"99",X"91",X"00",X"00",X"11",X"91",X"00",X"00",X"91",X"99",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"09",X"C9",X"00",X"00",X"09",X"CC",X"00",X"00",X"09",X"99",X"00",
		X"00",X"99",X"AA",X"00",X"00",X"9C",X"2A",X"00",X"00",X"9C",X"99",X"00",X"00",X"9C",X"C9",X"00",
		X"00",X"99",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"99",X"9C",X"00",X"00",X"44",X"CC",X"00",X"00",X"44",X"99",X"00",X"00",X"99",X"44",X"90",
		X"00",X"99",X"44",X"90",X"00",X"94",X"94",X"90",X"00",X"94",X"44",X"90",X"00",X"94",X"44",X"90",
		X"00",X"94",X"44",X"90",X"00",X"99",X"99",X"90",X"00",X"99",X"22",X"90",X"00",X"92",X"99",X"90",
		X"00",X"92",X"91",X"00",X"00",X"92",X"11",X"00",X"00",X"92",X"11",X"00",X"00",X"99",X"11",X"00",
		X"00",X"91",X"99",X"00",X"00",X"91",X"11",X"00",X"00",X"99",X"91",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"C9",X"00",X"00",X"09",X"CC",X"00",
		X"00",X"09",X"44",X"00",X"00",X"00",X"94",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"9C",X"00",X"00",X"00",X"C9",X"00",X"00",X"99",X"99",X"99",X"00",X"99",X"D9",X"99",
		X"00",X"F9",X"D4",X"99",X"00",X"99",X"44",X"99",X"00",X"99",X"94",X"99",X"00",X"99",X"94",X"99",
		X"00",X"99",X"49",X"99",X"00",X"99",X"D9",X"99",X"00",X"99",X"D9",X"99",X"00",X"99",X"D9",X"99",
		X"00",X"99",X"D9",X"99",X"00",X"99",X"D9",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"09",X"11",
		X"00",X"19",X"00",X"11",X"00",X"99",X"00",X"19",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"C9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"9C",X"99",X"00",X"00",X"9C",X"CC",X"00",
		X"00",X"99",X"44",X"00",X"00",X"09",X"94",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9C",X"00",
		X"00",X"00",X"CC",X"90",X"00",X"00",X"CC",X"90",X"00",X"00",X"99",X"90",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"F9",X"99",X"99",X"00",X"99",X"94",X"99",X"00",X"99",X"49",X"99",
		X"00",X"99",X"44",X"99",X"00",X"99",X"C9",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"09",X"99",X"00",X"00",X"09",X"11",X"00",X"00",X"09",X"11",X"00",X"00",X"09",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"99",X"00",
		X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",
		X"00",X"09",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"99",X"99",X"00",X"09",X"44",X"44",X"00",X"99",X"44",X"44",X"00",X"94",X"44",X"94",
		X"00",X"44",X"44",X"99",X"00",X"49",X"44",X"94",X"00",X"49",X"44",X"99",X"00",X"44",X"44",X"9C",
		X"00",X"44",X"99",X"9C",X"00",X"99",X"22",X"99",X"00",X"44",X"22",X"00",X"00",X"99",X"29",X"00",
		X"00",X"9C",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"90",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"9C",X"00",
		X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",
		X"00",X"00",X"CC",X"90",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"09",X"99",X"90",X"00",X"99",X"44",X"99",X"00",X"94",X"44",X"49",X"00",X"44",X"44",X"44",
		X"00",X"49",X"44",X"44",X"00",X"49",X"44",X"99",X"00",X"44",X"44",X"09",X"00",X"44",X"99",X"09",
		X"00",X"99",X"99",X"09",X"00",X"44",X"22",X"09",X"00",X"99",X"22",X"09",X"00",X"9C",X"99",X"09",
		X"00",X"9C",X"29",X"99",X"00",X"09",X"99",X"90",X"00",X"00",X"90",X"90",X"00",X"00",X"90",X"90",
		X"00",X"00",X"90",X"90",X"00",X"00",X"90",X"90",X"00",X"00",X"90",X"90",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"A9",
		X"00",X"00",X"CC",X"99",X"00",X"00",X"C9",X"99",X"00",X"00",X"CC",X"9C",X"00",X"00",X"99",X"CC",
		X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"99",X"00",X"00",X"C9",X"99",X"00",X"00",X"CC",X"99",
		X"00",X"00",X"CC",X"99",X"00",X"00",X"9C",X"44",X"00",X"00",X"99",X"99",X"00",X"00",X"44",X"94",
		X"99",X"09",X"44",X"94",X"91",X"09",X"99",X"99",X"91",X"99",X"99",X"90",X"91",X"99",X"44",X"99",
		X"91",X"99",X"44",X"29",X"91",X"92",X"99",X"22",X"91",X"92",X"99",X"92",X"91",X"22",X"00",X"22",
		X"99",X"29",X"00",X"22",X"00",X"99",X"00",X"22",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"91",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",
		X"00",X"00",X"99",X"C9",X"00",X"00",X"CC",X"99",X"00",X"00",X"C9",X"C9",X"00",X"00",X"CC",X"CC",
		X"00",X"00",X"99",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"99",X"00",X"00",X"C9",X"99",
		X"00",X"00",X"CC",X"99",X"00",X"00",X"CC",X"C9",X"00",X"00",X"9C",X"99",X"00",X"00",X"99",X"99",
		X"00",X"09",X"44",X"94",X"00",X"99",X"44",X"94",X"00",X"29",X"99",X"99",X"00",X"29",X"99",X"00",
		X"00",X"29",X"44",X"00",X"00",X"29",X"99",X"00",X"00",X"22",X"29",X"00",X"00",X"99",X"29",X"00",
		X"00",X"99",X"99",X"00",X"00",X"22",X"90",X"00",X"00",X"22",X"00",X"00",X"00",X"29",X"00",X"00",
		X"00",X"29",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"C9",X"00",X"00",X"99",X"C9",X"00",
		X"00",X"99",X"99",X"00",X"00",X"C9",X"A9",X"00",X"00",X"CC",X"9C",X"00",X"00",X"CC",X"9C",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"CC",X"99",X"00",X"00",X"CC",X"99",X"00",X"00",X"C9",X"99",X"00",X"00",X"CC",X"49",X"00",
		X"00",X"CC",X"49",X"00",X"00",X"99",X"44",X"00",X"00",X"99",X"99",X"00",X"00",X"94",X"49",X"00",
		X"00",X"99",X"44",X"00",X"00",X"92",X"99",X"00",X"00",X"99",X"22",X"00",X"00",X"91",X"22",X"00",
		X"00",X"11",X"22",X"00",X"00",X"11",X"92",X"00",X"00",X"11",X"99",X"00",X"00",X"99",X"91",X"00",
		X"00",X"11",X"99",X"00",X"00",X"91",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"09",X"CC",X"99",X"00",X"09",X"CC",X"99",X"00",X"00",X"99",X"90",
		X"00",X"00",X"29",X"90",X"00",X"00",X"A9",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"CC",X"90",
		X"00",X"09",X"9C",X"99",X"00",X"00",X"99",X"90",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"90",
		X"00",X"09",X"CC",X"90",X"00",X"99",X"9C",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"44",X"94",
		X"00",X"99",X"94",X"94",X"00",X"94",X"99",X"94",X"00",X"99",X"94",X"44",X"00",X"00",X"44",X"99",
		X"00",X"00",X"44",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"90",
		X"00",X"00",X"90",X"90",X"00",X"00",X"90",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"CC",X"90",X"00",X"00",X"CC",X"00",X"00",X"00",X"99",X"00",
		X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",
		X"00",X"99",X"CC",X"00",X"00",X"CC",X"CC",X"90",X"00",X"CC",X"99",X"90",X"00",X"C9",X"44",X"90",
		X"00",X"99",X"44",X"90",X"00",X"94",X"44",X"90",X"00",X"94",X"44",X"90",X"00",X"99",X"94",X"90",
		X"00",X"09",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"22",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"99",X"C9",X"00",X"00",X"99",X"CC",X"00",X"00",X"09",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"9C",X"99",X"00",X"00",X"9C",X"99",X"00",X"00",X"9C",X"99",X"00",
		X"00",X"99",X"CC",X"90",X"00",X"99",X"CC",X"90",X"00",X"C9",X"99",X"90",X"00",X"CC",X"44",X"90",
		X"00",X"C9",X"44",X"90",X"00",X"99",X"44",X"90",X"00",X"44",X"44",X"00",X"00",X"94",X"44",X"00",
		X"00",X"94",X"44",X"00",X"00",X"94",X"99",X"00",X"00",X"94",X"44",X"00",X"00",X"94",X"99",X"00",
		X"00",X"99",X"22",X"00",X"00",X"92",X"22",X"00",X"00",X"92",X"99",X"00",X"00",X"92",X"91",X"00",
		X"00",X"99",X"11",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"11",X"00",X"00",X"91",X"11",X"00",
		X"00",X"99",X"11",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"CC",X"90",X"00",X"00",X"99",X"90",X"09",X"99",X"9A",X"90",
		X"9D",X"DD",X"92",X"90",X"99",X"99",X"99",X"90",X"99",X"99",X"CC",X"90",X"99",X"F9",X"CC",X"90",
		X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"9C",X"00",
		X"CC",X"99",X"C9",X"00",X"CC",X"99",X"CC",X"00",X"CC",X"F9",X"99",X"90",X"99",X"99",X"99",X"90",
		X"99",X"99",X"44",X"90",X"9D",X"D9",X"44",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"49",X"00",
		X"99",X"99",X"44",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"22",X"00",X"99",X"99",X"29",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"29",X"00",X"99",X"99",X"99",X"00",X"99",X"F9",X"29",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"19",X"99",X"00",X"00",X"19",X"19",X"00",X"00",X"99",X"99",
		X"00",X"00",X"99",X"00",X"00",X"00",X"CC",X"90",X"00",X"00",X"2A",X"90",X"00",X"00",X"99",X"90",
		X"00",X"00",X"DD",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"49",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"C9",
		X"00",X"00",X"99",X"C9",X"00",X"00",X"DD",X"C9",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"19",X"19",X"00",X"00",X"99",X"99",
		X"00",X"00",X"99",X"90",X"00",X"00",X"CC",X"90",X"00",X"09",X"CC",X"90",X"00",X"09",X"99",X"90",
		X"00",X"09",X"99",X"90",X"00",X"09",X"99",X"90",X"00",X"09",X"99",X"90",X"00",X"09",X"99",X"90",
		X"00",X"09",X"CC",X"90",X"00",X"00",X"CC",X"90",X"00",X"99",X"CC",X"99",X"00",X"94",X"CC",X"94",
		X"00",X"94",X"99",X"44",X"00",X"94",X"99",X"44",X"00",X"99",X"44",X"49",X"00",X"09",X"44",X"99",
		X"00",X"00",X"44",X"90",X"00",X"00",X"49",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"44",X"90",
		X"00",X"00",X"99",X"90",X"00",X"00",X"22",X"90",X"00",X"00",X"22",X"90",X"00",X"00",X"22",X"90",
		X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"22",X"00",
		X"00",X"00",X"22",X"90",X"00",X"00",X"99",X"19",X"00",X"00",X"19",X"19",X"00",X"00",X"99",X"99",
		X"00",X"00",X"99",X"40",X"00",X"09",X"99",X"40",X"00",X"09",X"9A",X"40",X"00",X"09",X"9A",X"04",
		X"00",X"09",X"AA",X"04",X"00",X"09",X"AA",X"40",X"00",X"9C",X"99",X"40",X"00",X"9C",X"CC",X"40",
		X"00",X"9C",X"CC",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"44",X"CC",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"94",X"00",
		X"00",X"49",X"44",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"94",X"00",X"00",X"94",X"44",X"00",
		X"00",X"99",X"44",X"00",X"00",X"09",X"44",X"00",X"00",X"09",X"99",X"09",X"00",X"09",X"99",X"09",
		X"00",X"00",X"99",X"09",X"00",X"00",X"29",X"99",X"00",X"00",X"22",X"91",X"00",X"00",X"22",X"91",
		X"00",X"00",X"22",X"11",X"00",X"00",X"92",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"99",X"00",X"00",X"09",X"CC",X"00",X"00",X"09",X"CC",X"00",X"00",X"09",X"CC",X"00",
		X"00",X"09",X"C9",X"00",X"00",X"09",X"99",X"00",X"00",X"9C",X"9C",X"00",X"00",X"9C",X"CC",X"00",
		X"00",X"9C",X"CC",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"49",X"00",
		X"00",X"99",X"99",X"09",X"00",X"44",X"CC",X"99",X"00",X"44",X"99",X"49",X"00",X"44",X"94",X"49",
		X"00",X"49",X"44",X"99",X"00",X"49",X"99",X"00",X"00",X"49",X"94",X"00",X"00",X"49",X"44",X"09",
		X"00",X"49",X"94",X"09",X"00",X"49",X"94",X"09",X"00",X"49",X"99",X"99",X"00",X"49",X"99",X"29",
		X"00",X"49",X"99",X"29",X"00",X"49",X"99",X"99",X"00",X"99",X"90",X"00",X"00",X"09",X"90",X"00",
		X"00",X"09",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"90",X"AA",X"00",X"99",X"C9",X"00",X"00",X"99",X"CC",X"00",X"00",X"99",X"CC",X"AA",
		X"00",X"99",X"99",X"00",X"00",X"99",X"9C",X"AA",X"00",X"C9",X"CC",X"0A",X"00",X"C9",X"CC",X"00",
		X"00",X"CC",X"99",X"00",X"00",X"9C",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"9C",X"00",X"00",X"49",X"CC",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"44",X"00",
		X"00",X"49",X"44",X"00",X"00",X"49",X"99",X"00",X"00",X"49",X"94",X"00",X"00",X"49",X"44",X"09",
		X"00",X"49",X"94",X"09",X"00",X"49",X"94",X"09",X"00",X"49",X"99",X"99",X"00",X"99",X"99",X"29",
		X"00",X"49",X"99",X"29",X"00",X"49",X"99",X"99",X"00",X"99",X"90",X"00",X"00",X"09",X"90",X"00",
		X"00",X"09",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"DD",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"9F",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"9D",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"D9",X"00",X"00",X"09",X"9D",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",
		X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"D9",X"90",X"00",X"99",X"D9",X"99",
		X"00",X"99",X"D9",X"99",X"00",X"DD",X"DD",X"DD",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",
		X"00",X"00",X"9D",X"00",X"00",X"00",X"9D",X"00",X"00",X"00",X"9D",X"00",X"00",X"00",X"9D",X"00",
		X"00",X"00",X"9D",X"00",X"00",X"00",X"9D",X"00",X"00",X"00",X"9D",X"00",X"00",X"00",X"9D",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9D",X"00",
		X"00",X"00",X"9D",X"00",X"00",X"00",X"9D",X"00",X"00",X"00",X"9D",X"00",X"00",X"00",X"9D",X"00",
		X"00",X"00",X"9D",X"00",X"00",X"00",X"9D",X"00",X"00",X"00",X"9D",X"00",X"00",X"00",X"9D",X"00",
		X"00",X"00",X"9D",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"D9",X"90",X"00",X"00",X"9D",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"D9",X"00",X"00",X"00",X"9D",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",
		X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"99",
		X"00",X"00",X"9D",X"99",X"00",X"00",X"9D",X"99",X"00",X"00",X"99",X"9D",X"00",X"00",X"99",X"DD",
		X"00",X"00",X"99",X"D9",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",
		X"00",X"00",X"D9",X"99",X"00",X"00",X"DD",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"DD",X"DD",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"FF",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"DD",X"D9",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"00",X"00",
		X"00",X"F9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"DD",X"00",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"09",X"9F",X"99",X"00",X"09",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"9D",X"DD",X"DD",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"F9",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"F9",X"90",X"00",
		X"00",X"99",X"99",X"00",X"00",X"DD",X"D9",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"FF",X"00",X"00",X"99",X"99",X"00",
		X"00",X"DD",X"DD",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"CC",X"00",X"00",X"9C",X"99",X"00",X"00",X"9C",X"9E",X"99",
		X"00",X"CC",X"EC",X"C9",X"00",X"9C",X"EC",X"C9",X"00",X"CC",X"C9",X"C9",X"00",X"9C",X"99",X"99",
		X"00",X"9C",X"CC",X"99",X"00",X"9C",X"99",X"99",X"00",X"9C",X"9F",X"99",X"00",X"9C",X"99",X"99",
		X"09",X"99",X"9F",X"99",X"09",X"99",X"99",X"99",X"09",X"99",X"44",X"99",X"09",X"D9",X"CC",X"99",
		X"09",X"D9",X"99",X"99",X"09",X"D9",X"99",X"99",X"09",X"D9",X"99",X"99",X"09",X"99",X"99",X"99",
		X"09",X"99",X"44",X"CC",X"09",X"99",X"44",X"CC",X"09",X"99",X"44",X"CC",X"09",X"99",X"49",X"CC",
		X"09",X"99",X"99",X"9C",X"99",X"99",X"99",X"99",X"9C",X"99",X"99",X"CC",X"99",X"99",X"C9",X"CC",
		X"09",X"99",X"C9",X"CE",X"09",X"99",X"CC",X"CE",X"09",X"99",X"CC",X"EC",X"09",X"99",X"CC",X"99",
		X"09",X"99",X"CC",X"99",X"09",X"C9",X"99",X"BB",X"09",X"CC",X"BB",X"BB",X"09",X"99",X"BB",X"BB",
		X"09",X"BB",X"BB",X"BB",X"09",X"BB",X"9B",X"BB",X"09",X"BB",X"9B",X"BB",X"00",X"BB",X"9B",X"BB",
		X"00",X"BB",X"9B",X"BB",X"00",X"BB",X"9B",X"BB",X"00",X"BB",X"9B",X"BB",X"00",X"BB",X"99",X"BB",
		X"00",X"99",X"9B",X"BB",X"00",X"EE",X"9B",X"B9",X"00",X"77",X"9B",X"B9",X"00",X"77",X"99",X"B9",
		X"00",X"77",X"99",X"B9",X"00",X"77",X"9B",X"B9",X"00",X"99",X"9B",X"B9",X"00",X"77",X"9B",X"B9",
		X"00",X"77",X"B9",X"99",X"00",X"99",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"99",X"99",
		X"00",X"00",X"97",X"79",X"00",X"00",X"99",X"99",X"00",X"00",X"97",X"90",X"00",X"00",X"99",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"95",X"55",X"00",X"00",X"22",X"59",X"00",X"00",X"99",X"59",X"00",
		X"09",X"22",X"99",X"00",X"09",X"55",X"90",X"00",X"99",X"55",X"00",X"90",X"9F",X"59",X"99",X"99",
		X"99",X"59",X"95",X"99",X"99",X"99",X"55",X"99",X"95",X"99",X"55",X"99",X"99",X"55",X"55",X"59",
		X"09",X"99",X"99",X"59",X"00",X"00",X"99",X"55",X"00",X"00",X"99",X"55",X"00",X"00",X"55",X"55",
		X"00",X"00",X"55",X"55",X"00",X"00",X"55",X"55",X"00",X"00",X"99",X"55",X"00",X"00",X"59",X"59",
		X"00",X"00",X"55",X"99",X"00",X"00",X"55",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"77",
		X"00",X"00",X"95",X"99",X"00",X"00",X"95",X"59",X"00",X"00",X"55",X"99",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"95",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"92",X"00",X"00",X"09",X"99",X"00",X"00",
		X"09",X"55",X"99",X"00",X"99",X"55",X"59",X"00",X"9F",X"99",X"95",X"90",X"99",X"59",X"99",X"99",
		X"99",X"59",X"55",X"99",X"95",X"99",X"55",X"99",X"99",X"94",X"55",X"99",X"09",X"44",X"59",X"59",
		X"00",X"44",X"99",X"59",X"00",X"44",X"55",X"55",X"00",X"99",X"99",X"55",X"00",X"99",X"99",X"55",
		X"00",X"99",X"55",X"55",X"99",X"55",X"55",X"55",X"97",X"59",X"99",X"55",X"99",X"99",X"00",X"55",
		X"99",X"90",X"00",X"95",X"95",X"00",X"00",X"99",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"CC",X"00",X"00",X"09",X"9C",X"00",X"00",X"09",X"9C",X"00",
		X"00",X"09",X"9C",X"00",X"00",X"09",X"9C",X"00",X"00",X"09",X"CC",X"00",X"00",X"09",X"CC",X"00",
		X"00",X"09",X"CC",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"44",X"CC",X"00",X"00",X"44",X"99",X"00",X"00",X"94",X"94",X"99",
		X"00",X"99",X"44",X"99",X"00",X"99",X"44",X"99",X"00",X"97",X"94",X"99",X"00",X"97",X"99",X"99",
		X"00",X"99",X"9C",X"99",X"00",X"99",X"CC",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"22",X"99",
		X"00",X"9F",X"22",X"99",X"00",X"99",X"22",X"99",X"00",X"99",X"22",X"99",X"00",X"99",X"22",X"99",
		X"00",X"00",X"99",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"09",X"C9",X"00",X"00",X"99",X"CC",X"00",X"00",X"99",X"C9",X"00",
		X"00",X"99",X"C9",X"00",X"00",X"99",X"C9",X"00",X"00",X"9C",X"CC",X"00",X"00",X"9C",X"CC",X"00",
		X"00",X"9C",X"CC",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"44",X"CC",X"00",X"00",X"44",X"99",X"99",X"00",X"49",X"94",X"99",
		X"00",X"99",X"44",X"99",X"00",X"99",X"44",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"44",X"99",
		X"00",X"99",X"44",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"22",X"99",X"00",X"F9",X"22",X"99",
		X"00",X"99",X"99",X"91",X"00",X"99",X"99",X"91",X"00",X"92",X"99",X"11",X"00",X"92",X"00",X"19",
		X"00",X"19",X"00",X"19",X"00",X"11",X"00",X"99",X"00",X"11",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"99",X"C9",X"00",X"00",X"09",X"CC",X"00",X"09",X"99",X"C9",X"00",
		X"99",X"99",X"C9",X"00",X"9C",X"99",X"C9",X"00",X"9C",X"9C",X"C9",X"00",X"99",X"9C",X"CC",X"00",
		X"09",X"9C",X"CC",X"00",X"09",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"94",X"99",X"00",X"00",X"44",X"CC",X"00",X"00",X"44",X"99",X"00",X"00",X"99",X"94",X"00",
		X"00",X"99",X"44",X"00",X"00",X"09",X"44",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"44",X"00",
		X"00",X"09",X"44",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"22",X"09",X"00",X"00",X"22",X"99",
		X"00",X"09",X"99",X"91",X"00",X"99",X"09",X"91",X"00",X"92",X"00",X"11",X"00",X"92",X"00",X"19",
		X"00",X"19",X"00",X"19",X"00",X"11",X"00",X"99",X"00",X"11",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"60",X"99",X"06",X"00",X"00",X"99",X"06",X"05",X"09",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"9C",X"00",X"00",X"99",X"9F",X"00",X"00",X"99",X"FF",X"99",
		X"03",X"C9",X"FF",X"C9",X"00",X"99",X"9F",X"C9",X"00",X"CC",X"C9",X"C9",X"00",X"9C",X"C9",X"99",
		X"00",X"9C",X"9C",X"99",X"00",X"99",X"CC",X"99",X"00",X"9C",X"C9",X"99",X"00",X"9C",X"99",X"99",
		X"09",X"99",X"49",X"99",X"09",X"99",X"44",X"99",X"09",X"99",X"99",X"99",X"09",X"D9",X"C9",X"99",
		X"09",X"D9",X"99",X"99",X"09",X"D9",X"99",X"99",X"09",X"D9",X"99",X"9C",X"09",X"99",X"99",X"CC",
		X"09",X"99",X"94",X"CC",X"09",X"99",X"94",X"CC",X"09",X"99",X"44",X"CC",X"09",X"99",X"99",X"99",
		X"99",X"09",X"99",X"00",X"90",X"99",X"09",X"90",X"00",X"09",X"09",X"99",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"44",X"00",X"00",X"94",X"4A",X"00",X"00",X"94",X"4A",X"99",
		X"00",X"44",X"EA",X"49",X"00",X"94",X"E4",X"49",X"00",X"44",X"49",X"49",X"00",X"94",X"99",X"99",
		X"00",X"94",X"44",X"99",X"00",X"94",X"99",X"99",X"00",X"94",X"F9",X"99",X"00",X"94",X"99",X"99",
		X"09",X"99",X"F9",X"99",X"09",X"99",X"F9",X"99",X"09",X"99",X"99",X"99",X"09",X"D9",X"44",X"99",
		X"09",X"D9",X"99",X"99",X"09",X"D9",X"99",X"99",X"09",X"D9",X"99",X"99",X"09",X"99",X"99",X"99",
		X"09",X"99",X"44",X"CC",X"09",X"99",X"44",X"CC",X"09",X"99",X"44",X"CC",X"09",X"99",X"49",X"CC",
		X"09",X"99",X"99",X"9C",X"99",X"99",X"99",X"99",X"9C",X"99",X"99",X"CC",X"99",X"99",X"C9",X"CC",
		X"09",X"99",X"C9",X"CE",X"09",X"99",X"CC",X"CE",X"09",X"99",X"CC",X"EC",X"09",X"99",X"CC",X"99",
		X"09",X"99",X"CC",X"99",X"09",X"C9",X"99",X"FF",X"09",X"CC",X"FF",X"44",X"09",X"99",X"FF",X"44",
		X"09",X"44",X"FF",X"FF",X"09",X"FF",X"F9",X"FF",X"09",X"F4",X"F9",X"44",X"09",X"F4",X"99",X"44",
		X"09",X"99",X"09",X"99",X"00",X"EE",X"09",X"EE",X"00",X"EE",X"99",X"CC",X"00",X"CE",X"9E",X"99",
		X"00",X"CE",X"9C",X"90",X"00",X"CC",X"9E",X"90",X"00",X"CE",X"9C",X"99",X"00",X"CC",X"9E",X"CC",
		X"09",X"EC",X"99",X"EC",X"09",X"CE",X"09",X"CE",X"99",X"9C",X"00",X"E9",X"91",X"9C",X"00",X"99",
		X"9B",X"99",X"99",X"9B",X"9B",X"BB",X"9B",X"BB",X"99",X"9B",X"B9",X"BB",X"09",X"BB",X"99",X"BB",
		X"09",X"9B",X"99",X"9B",X"09",X"BB",X"BB",X"99",X"0B",X"B9",X"BB",X"BB",X"09",X"99",X"99",X"B9",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"12",
		X"00",X"99",X"00",X"22",X"90",X"CC",X"00",X"99",X"40",X"C9",X"00",X"9B",X"40",X"99",X"09",X"99",
		X"40",X"C9",X"99",X"E9",X"22",X"C9",X"99",X"99",X"A0",X"C9",X"97",X"45",X"A0",X"99",X"97",X"45",
		X"A0",X"96",X"97",X"45",X"F0",X"66",X"97",X"45",X"00",X"66",X"97",X"45",X"00",X"69",X"97",X"45",
		X"00",X"99",X"97",X"45",X"00",X"92",X"97",X"45",X"00",X"26",X"97",X"45",X"00",X"66",X"97",X"45",
		X"00",X"99",X"99",X"47",X"00",X"AA",X"09",X"47",X"00",X"AA",X"00",X"47",X"00",X"A9",X"00",X"99",
		X"00",X"99",X"00",X"95",X"00",X"9E",X"00",X"95",X"00",X"99",X"00",X"99",X"00",X"9E",X"09",X"99",
		X"00",X"99",X"99",X"59",X"00",X"99",X"9B",X"59",X"00",X"99",X"99",X"99",X"00",X"99",X"09",X"00",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"12",
		X"F0",X"99",X"00",X"22",X"A0",X"CC",X"00",X"99",X"A0",X"C9",X"00",X"9B",X"A0",X"99",X"09",X"99",
		X"22",X"C9",X"99",X"99",X"40",X"C9",X"97",X"45",X"40",X"C9",X"97",X"45",X"40",X"99",X"97",X"45",
		X"90",X"96",X"97",X"45",X"00",X"66",X"97",X"45",X"00",X"66",X"97",X"45",X"00",X"69",X"97",X"45",
		X"00",X"99",X"97",X"45",X"00",X"92",X"97",X"45",X"00",X"26",X"97",X"45",X"00",X"66",X"99",X"47",
		X"00",X"66",X"09",X"47",X"00",X"99",X"00",X"47",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"95",
		X"00",X"A9",X"90",X"95",X"00",X"AA",X"90",X"99",X"09",X"9A",X"90",X"90",X"99",X"9A",X"90",X"99",
		X"99",X"99",X"00",X"59",X"99",X"09",X"00",X"59",X"09",X"00",X"00",X"99",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"42",X"00",X"00",X"00",X"C2",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"99",X"CC",X"90",X"00",X"9A",X"C9",X"99",X"00",X"AA",X"CC",X"A9",X"00",X"AA",X"CC",X"AA",
		X"00",X"AA",X"99",X"A9",X"00",X"9A",X"A9",X"99",X"00",X"C9",X"A9",X"9C",X"00",X"99",X"29",X"99",
		X"00",X"92",X"A2",X"99",X"99",X"92",X"AA",X"90",X"90",X"9A",X"AA",X"90",X"99",X"9A",X"AA",X"99",
		X"94",X"9A",X"A2",X"09",X"94",X"9A",X"2A",X"99",X"94",X"99",X"AA",X"99",X"94",X"59",X"99",X"99",
		X"94",X"59",X"00",X"09",X"94",X"59",X"00",X"09",X"94",X"59",X"00",X"09",X"99",X"99",X"00",X"09",
		X"00",X"22",X"00",X"09",X"00",X"99",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"C4",X"00",X"00",X"00",X"CC",X"00",X"00",X"99",X"CC",X"90",
		X"00",X"9A",X"CC",X"99",X"00",X"AA",X"CC",X"A9",X"00",X"AA",X"CC",X"AA",X"00",X"AA",X"CC",X"A9",
		X"00",X"9A",X"99",X"99",X"00",X"C9",X"A9",X"9C",X"00",X"99",X"A9",X"99",X"00",X"92",X"29",X"99",
		X"99",X"92",X"A2",X"90",X"90",X"92",X"AA",X"90",X"99",X"9A",X"AA",X"99",X"94",X"99",X"AA",X"99",
		X"94",X"99",X"A2",X"99",X"94",X"99",X"2A",X"99",X"94",X"9A",X"AA",X"99",X"94",X"99",X"99",X"99",
		X"94",X"90",X"09",X"09",X"94",X"90",X"00",X"09",X"99",X"90",X"00",X"09",X"00",X"90",X"00",X"99",
		X"00",X"90",X"00",X"29",X"00",X"00",X"00",X"99",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"99",X"E4",X"00",X"00",X"9A",X"E4",X"90",
		X"00",X"AA",X"EE",X"99",X"00",X"AA",X"EE",X"A9",X"00",X"AA",X"4E",X"AA",X"00",X"AA",X"49",X"A9",
		X"00",X"9A",X"99",X"99",X"00",X"C9",X"9A",X"9C",X"00",X"99",X"AA",X"99",X"00",X"09",X"AA",X"99",
		X"00",X"99",X"99",X"90",X"00",X"92",X"AA",X"90",X"00",X"9A",X"A9",X"99",X"00",X"99",X"A9",X"A9",
		X"00",X"99",X"A9",X"A9",X"00",X"99",X"A9",X"99",X"00",X"9A",X"AA",X"A9",X"00",X"99",X"99",X"99",
		X"00",X"90",X"09",X"09",X"00",X"90",X"00",X"09",X"00",X"90",X"00",X"09",X"00",X"90",X"00",X"99",
		X"00",X"90",X"00",X"29",X"00",X"00",X"00",X"99",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"55",X"00",X"00",X"95",X"99",X"00",
		X"00",X"55",X"FF",X"00",X"00",X"55",X"FF",X"90",X"00",X"59",X"99",X"90",X"00",X"99",X"99",X"90",
		X"00",X"9F",X"99",X"90",X"00",X"99",X"49",X"90",X"00",X"99",X"49",X"90",X"00",X"9F",X"49",X"90",
		X"00",X"9F",X"99",X"90",X"00",X"99",X"FF",X"90",X"00",X"59",X"FF",X"90",X"00",X"55",X"FF",X"90",
		X"00",X"95",X"FF",X"00",X"00",X"95",X"FF",X"00",X"00",X"99",X"99",X"99",X"00",X"09",X"55",X"99",
		X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"92",X"99",X"99",X"00",X"22",X"22",X"44",X"00",X"99",X"29",X"44",
		X"00",X"C9",X"99",X"55",X"00",X"9C",X"49",X"99",X"00",X"CC",X"99",X"C9",X"0D",X"9C",X"00",X"99",
		X"0D",X"99",X"90",X"94",X"09",X"09",X"90",X"94",X"00",X"09",X"99",X"44",X"DD",X"99",X"93",X"99",
		X"D9",X"93",X"33",X"00",X"D9",X"93",X"39",X"00",X"09",X"93",X"99",X"00",X"09",X"93",X"99",X"00",
		X"09",X"99",X"9A",X"90",X"09",X"69",X"9A",X"99",X"00",X"69",X"99",X"66",X"09",X"69",X"96",X"66",
		X"09",X"66",X"66",X"66",X"09",X"22",X"22",X"22",X"09",X"22",X"22",X"22",X"99",X"99",X"22",X"99",
		X"9D",X"77",X"22",X"77",X"9D",X"75",X"66",X"57",X"9D",X"99",X"66",X"97",X"9D",X"D9",X"66",X"99",
		X"99",X"99",X"99",X"97",X"00",X"77",X"00",X"77",X"00",X"77",X"00",X"74",X"00",X"99",X"00",X"99",
		X"00",X"99",X"09",X"00",X"00",X"92",X"92",X"00",X"00",X"22",X"29",X"99",X"00",X"99",X"99",X"49",
		X"00",X"CE",X"99",X"49",X"00",X"9E",X"49",X"49",X"00",X"CC",X"99",X"49",X"0D",X"9C",X"55",X"99",
		X"0D",X"99",X"58",X"00",X"09",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"DD",X"99",X"93",X"00",
		X"D9",X"93",X"33",X"00",X"D9",X"93",X"33",X"00",X"09",X"93",X"99",X"00",X"09",X"93",X"99",X"00",
		X"09",X"93",X"99",X"00",X"09",X"99",X"9A",X"90",X"09",X"69",X"9A",X"99",X"00",X"69",X"99",X"66",
		X"09",X"69",X"96",X"66",X"09",X"66",X"66",X"66",X"09",X"99",X"22",X"99",X"09",X"77",X"22",X"79",
		X"99",X"77",X"22",X"77",X"9D",X"97",X"22",X"77",X"9D",X"D9",X"66",X"97",X"9D",X"99",X"66",X"97",
		X"9D",X"97",X"66",X"75",X"09",X"77",X"99",X"55",X"00",X"77",X"00",X"59",X"00",X"99",X"00",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"09",X"99",X"00",X"99",X"9E",X"E9",X"00",X"E9",X"9E",X"E9",
		X"00",X"E9",X"9E",X"99",X"00",X"E9",X"99",X"90",X"00",X"EE",X"E9",X"90",X"00",X"EE",X"EE",X"99",
		X"00",X"9E",X"EE",X"E9",X"00",X"9E",X"E9",X"E9",X"00",X"9E",X"E9",X"E9",X"00",X"9E",X"99",X"99",
		X"00",X"EE",X"99",X"00",X"00",X"99",X"E9",X"00",X"00",X"99",X"EE",X"00",X"00",X"90",X"9E",X"00",
		X"00",X"90",X"99",X"00",X"00",X"90",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"99",X"00",X"00",X"9E",X"E9",X"00",X"90",X"9E",X"E9",X"00",X"99",X"9E",X"99",
		X"00",X"E9",X"99",X"90",X"00",X"EE",X"E9",X"90",X"00",X"9E",X"EE",X"99",X"00",X"EE",X"EE",X"99",
		X"00",X"EE",X"E9",X"E9",X"00",X"9E",X"E9",X"E9",X"00",X"9E",X"E9",X"99",X"00",X"9E",X"EE",X"99",
		X"00",X"99",X"E9",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"09",X"9E",X"00",
		X"00",X"09",X"9E",X"00",X"00",X"09",X"E9",X"00",X"00",X"09",X"E9",X"00",X"00",X"00",X"E9",X"00",
		X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"EE",X"00",X"00",X"99",X"9E",X"00",
		X"00",X"9E",X"99",X"00",X"00",X"9E",X"90",X"00",X"00",X"EE",X"90",X"00",X"00",X"E9",X"99",X"00",
		X"00",X"E9",X"E9",X"00",X"00",X"E9",X"E9",X"00",X"00",X"EE",X"E9",X"00",X"00",X"EE",X"99",X"00",
		X"00",X"99",X"90",X"00",X"00",X"E9",X"90",X"00",X"00",X"EE",X"99",X"00",X"00",X"9E",X"EE",X"00",
		X"00",X"E9",X"EE",X"00",X"00",X"EE",X"99",X"00",X"00",X"EE",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"09",
		X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"AA",X"00",X"99",X"9D",X"99",X"00",X"AA",X"99",X"AA",
		X"00",X"99",X"99",X"AA",X"00",X"AA",X"99",X"99",X"00",X"99",X"55",X"09",X"00",X"90",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"99",X"00",X"FF",X"00",X"44",X"00",X"FF",X"00",X"99",X"00",X"FF",X"00",X"99",X"00",
		X"00",X"F0",X"9A",X"00",X"00",X"F0",X"C9",X"00",X"00",X"99",X"C9",X"00",X"00",X"C9",X"99",X"00",
		X"00",X"C9",X"44",X"00",X"00",X"99",X"C9",X"00",X"00",X"C9",X"99",X"00",X"00",X"99",X"55",X"00",
		X"00",X"95",X"99",X"00",X"00",X"95",X"99",X"00",X"00",X"95",X"55",X"00",X"00",X"99",X"55",X"00",
		X"00",X"09",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"44",X"92",X"00",X"00",X"94",X"99",X"00",X"00",X"99",X"29",X"00",
		X"00",X"EE",X"22",X"00",X"00",X"EE",X"22",X"00",X"00",X"99",X"92",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"C9",X"00",
		X"00",X"00",X"C9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"79",X"00",X"00",X"00",X"79",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"C9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"C9",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"00",
		X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"09",X"92",X"00",X"00",X"09",X"92",X"00",
		X"00",X"09",X"99",X"00",X"00",X"09",X"FF",X"00",X"00",X"09",X"FF",X"00",X"00",X"09",X"FF",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"49",X"00",X"00",X"99",X"44",X"00",X"09",X"99",X"94",X"00",
		X"09",X"94",X"A9",X"00",X"09",X"99",X"99",X"00",X"09",X"9C",X"CC",X"00",X"00",X"99",X"CC",X"00",
		X"00",X"99",X"44",X"00",X"00",X"99",X"44",X"00",X"09",X"99",X"C9",X"00",X"09",X"92",X"99",X"00",
		X"09",X"29",X"22",X"00",X"09",X"29",X"22",X"00",X"00",X"99",X"29",X"00",X"00",X"92",X"29",X"00",
		X"00",X"92",X"29",X"00",X"00",X"92",X"29",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"99",X"00",
		X"00",X"96",X"99",X"00",X"00",X"96",X"69",X"00",X"00",X"96",X"69",X"00",X"00",X"96",X"66",X"00",
		X"00",X"99",X"69",X"00",X"00",X"11",X"69",X"00",X"00",X"11",X"69",X"00",X"00",X"11",X"69",X"00",
		X"00",X"99",X"99",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"99",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"CC",X"00",X"99",X"99",X"CC",X"99",X"99",X"99",X"99",X"99",
		X"00",X"90",X"22",X"90",X"00",X"90",X"22",X"90",X"00",X"90",X"22",X"90",X"00",X"90",X"22",X"90",
		X"00",X"90",X"22",X"90",X"99",X"99",X"22",X"99",X"99",X"99",X"22",X"99",X"00",X"00",X"29",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",
		X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"90",
		X"00",X"00",X"99",X"99",X"00",X"00",X"66",X"69",X"00",X"00",X"66",X"66",X"00",X"09",X"99",X"96",
		X"00",X"09",X"66",X"96",X"00",X"09",X"66",X"99",X"00",X"09",X"99",X"00",X"00",X"09",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"99",X"00",X"00",X"77",X"9C",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"99",
		X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"09",X"00",X"00",X"94",X"09",X"00",X"00",X"99",X"09",
		X"00",X"00",X"44",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"CC",X"99",X"00",X"00",X"99",X"99",
		X"00",X"00",X"22",X"29",X"00",X"00",X"29",X"99",X"00",X"00",X"29",X"99",X"00",X"00",X"29",X"00",
		X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"69",X"00",
		X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"69",X"19",X"00",X"00",X"69",X"99",
		X"00",X"00",X"99",X"19",X"00",X"00",X"19",X"19",X"00",X"00",X"19",X"99",X"00",X"00",X"99",X"90",
		X"00",X"99",X"99",X"00",X"00",X"CC",X"44",X"00",X"99",X"C9",X"44",X"99",X"99",X"99",X"44",X"99",
		X"00",X"29",X"44",X"00",X"00",X"29",X"94",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"C9",X"00",
		X"00",X"00",X"CC",X"00",X"99",X"99",X"CC",X"99",X"99",X"99",X"99",X"99",X"00",X"00",X"99",X"00",
		X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"09",X"29",X"00",
		X"00",X"09",X"29",X"00",X"00",X"09",X"29",X"00",X"00",X"09",X"29",X"00",X"00",X"09",X"99",X"00",
		X"00",X"09",X"C9",X"00",X"00",X"09",X"C9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"09",X"69",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"19",X"00",
		X"00",X"11",X"19",X"00",X"00",X"91",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"09",X"99",X"00",X"49",X"09",X"69",X"09",X"44",X"09",X"99",X"99",X"44",X"96",X"99",
		X"99",X"99",X"96",X"90",X"09",X"EE",X"96",X"90",X"09",X"CC",X"99",X"99",X"09",X"CC",X"00",X"11",
		X"00",X"9C",X"00",X"91",X"00",X"99",X"00",X"91",X"00",X"CC",X"00",X"11",X"00",X"99",X"00",X"91",
		X"00",X"55",X"00",X"91",X"00",X"99",X"00",X"91",X"00",X"59",X"00",X"91",X"00",X"99",X"00",X"91",
		X"00",X"9C",X"90",X"91",X"00",X"99",X"90",X"91",X"00",X"55",X"99",X"99",X"00",X"55",X"99",X"44",
		X"00",X"99",X"90",X"44",X"00",X"11",X"00",X"44",X"00",X"19",X"99",X"44",X"00",X"11",X"99",X"44",
		X"09",X"11",X"99",X"44",X"09",X"99",X"99",X"44",X"99",X"99",X"90",X"99",X"99",X"09",X"90",X"95",
		X"99",X"00",X"00",X"59",X"99",X"00",X"00",X"7A",X"99",X"00",X"00",X"97",X"99",X"00",X"00",X"99",
		X"00",X"99",X"00",X"99",X"00",X"44",X"00",X"79",X"00",X"44",X"00",X"79",X"09",X"44",X"00",X"7A",
		X"09",X"99",X"00",X"7A",X"00",X"EE",X"00",X"96",X"00",X"EC",X"00",X"96",X"00",X"CC",X"00",X"96",
		X"00",X"99",X"00",X"99",X"00",X"C9",X"00",X"91",X"00",X"CC",X"00",X"91",X"00",X"99",X"00",X"91",
		X"00",X"99",X"00",X"11",X"00",X"59",X"00",X"91",X"00",X"99",X"00",X"91",X"00",X"9C",X"90",X"91",
		X"00",X"99",X"90",X"91",X"00",X"55",X"99",X"99",X"00",X"55",X"99",X"44",X"00",X"99",X"90",X"44",
		X"00",X"11",X"00",X"44",X"00",X"11",X"00",X"44",X"00",X"11",X"00",X"44",X"00",X"19",X"00",X"44",
		X"00",X"19",X"00",X"44",X"00",X"19",X"00",X"99",X"00",X"19",X"00",X"57",X"00",X"19",X"00",X"55",
		X"00",X"19",X"00",X"9A",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"55",X"00",X"99",X"00",X"99",
		X"00",X"00",X"99",X"00",X"00",X"00",X"CC",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"9A",X"90",
		X"00",X"00",X"9A",X"90",X"00",X"90",X"99",X"90",X"00",X"90",X"CC",X"90",X"00",X"90",X"CC",X"90",
		X"00",X"99",X"99",X"90",X"00",X"99",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"9C",X"00",
		X"00",X"94",X"C9",X"00",X"00",X"99",X"CC",X"90",X"00",X"09",X"99",X"99",X"00",X"00",X"44",X"49",
		X"00",X"00",X"49",X"44",X"00",X"00",X"99",X"44",X"00",X"00",X"9C",X"49",X"00",X"00",X"9C",X"99",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"22",X"00",X"00",X"19",X"29",X"00",
		X"00",X"11",X"99",X"00",X"00",X"11",X"99",X"00",X"00",X"91",X"09",X"00",X"00",X"91",X"09",X"00",
		X"00",X"99",X"09",X"00",X"00",X"09",X"09",X"99",X"00",X"00",X"09",X"19",X"00",X"00",X"09",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F9",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"F9",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"49",X"00",X"00",X"09",X"44",X"00",
		X"00",X"94",X"44",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"A9",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"9C",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"C4",X"00",X"00",X"00",X"94",X"00",
		X"00",X"00",X"99",X"00",X"00",X"09",X"97",X"00",X"00",X"99",X"77",X"00",X"00",X"97",X"97",X"00",
		X"00",X"99",X"77",X"00",X"00",X"C9",X"99",X"00",X"00",X"C9",X"97",X"00",X"00",X"99",X"77",X"00",
		X"00",X"09",X"99",X"00",X"00",X"99",X"DD",X"90",X"00",X"94",X"D9",X"90",X"00",X"94",X"99",X"90",
		X"00",X"94",X"D9",X"90",X"00",X"99",X"99",X"99",X"00",X"94",X"09",X"99",X"00",X"99",X"09",X"99",
		X"00",X"09",X"00",X"99",X"00",X"09",X"00",X"99",X"00",X"09",X"00",X"90",X"00",X"0A",X"09",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",
		X"00",X"90",X"99",X"11",X"09",X"99",X"11",X"44",X"09",X"41",X"11",X"55",X"09",X"41",X"77",X"66",
		X"09",X"99",X"77",X"11",X"00",X"90",X"11",X"11",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"91",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"91",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"9C",X"00",X"00",X"C9",X"C9",X"00",X"00",X"CC",X"CC",X"00",
		X"00",X"44",X"4C",X"00",X"00",X"49",X"4C",X"00",X"00",X"C9",X"C9",X"00",X"00",X"CC",X"C9",X"00",
		X"00",X"9C",X"99",X"00",X"00",X"99",X"94",X"00",X"00",X"49",X"99",X"00",X"00",X"44",X"99",X"00",
		X"09",X"44",X"99",X"00",X"09",X"44",X"99",X"00",X"09",X"44",X"99",X"00",X"09",X"44",X"99",X"00",
		X"09",X"99",X"99",X"00",X"09",X"29",X"99",X"00",X"09",X"22",X"99",X"00",X"09",X"99",X"99",X"00",
		X"09",X"19",X"99",X"00",X"00",X"11",X"99",X"00",X"00",X"11",X"99",X"00",X"00",X"11",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"11",X"99",X"00",X"00",X"19",X"99",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"C9",X"99",X"00",X"00",X"9C",X"9C",X"00",X"00",X"CC",X"CC",X"00",
		X"00",X"44",X"44",X"00",X"00",X"C9",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"9C",X"CC",X"00",
		X"00",X"99",X"C9",X"00",X"00",X"99",X"99",X"00",X"00",X"49",X"94",X"00",X"00",X"44",X"99",X"00",
		X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",
		X"00",X"44",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"99",X"00",
		X"00",X"22",X"19",X"00",X"00",X"99",X"11",X"00",X"00",X"29",X"11",X"00",X"00",X"99",X"11",X"00",
		X"00",X"19",X"99",X"00",X"00",X"19",X"11",X"00",X"00",X"99",X"19",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",
		X"00",X"09",X"9C",X"00",X"00",X"99",X"99",X"00",X"00",X"CC",X"9C",X"00",X"00",X"CC",X"C9",X"00",
		X"00",X"9C",X"CC",X"00",X"00",X"99",X"44",X"00",X"00",X"09",X"9C",X"00",X"00",X"09",X"CC",X"00",
		X"00",X"00",X"C9",X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"94",X"99",X"00",X"99",X"44",X"99",
		X"00",X"99",X"44",X"9F",X"00",X"99",X"44",X"99",X"00",X"99",X"49",X"99",X"00",X"99",X"99",X"99",
		X"00",X"F9",X"99",X"99",X"09",X"99",X"99",X"99",X"09",X"99",X"99",X"99",X"09",X"99",X"99",X"99",
		X"09",X"99",X"99",X"9F",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"29",X"99",X"00",
		X"00",X"99",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"90",X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"9A",X"CC",X"00",X"00",X"9A",X"9C",X"00",X"00",X"C9",X"CC",X"00",X"00",X"CC",X"99",X"00",
		X"00",X"CC",X"CC",X"00",X"00",X"99",X"44",X"00",X"00",X"99",X"9C",X"00",X"00",X"99",X"CC",X"00",
		X"00",X"09",X"CC",X"00",X"00",X"00",X"C9",X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"99",X"99",
		X"09",X"99",X"94",X"99",X"09",X"99",X"44",X"F9",X"09",X"99",X"44",X"99",X"09",X"99",X"49",X"99",
		X"09",X"99",X"99",X"99",X"09",X"F9",X"99",X"99",X"09",X"99",X"99",X"99",X"09",X"99",X"99",X"99",
		X"09",X"99",X"99",X"99",X"09",X"99",X"F9",X"F9",X"09",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"91",X"00",X"00",X"11",X"91",X"00",X"00",X"11",X"91",X"00",X"00",X"99",X"99",X"00",
		X"00",X"00",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"C9",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"CC",X"99",X"00",X"00",X"CC",X"99",X"00",X"00",X"CC",X"9C",X"00",
		X"00",X"9C",X"CC",X"00",X"00",X"9C",X"CC",X"00",X"00",X"99",X"CC",X"00",X"00",X"09",X"C9",X"00",
		X"00",X"99",X"99",X"90",X"00",X"94",X"44",X"99",X"00",X"44",X"44",X"49",X"00",X"99",X"44",X"49",
		X"00",X"99",X"44",X"99",X"00",X"99",X"44",X"49",X"00",X"99",X"44",X"99",X"00",X"99",X"44",X"C9",
		X"00",X"99",X"99",X"C9",X"00",X"99",X"22",X"99",X"00",X"99",X"92",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"92",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"09",X"C9",X"00",X"00",X"09",X"CC",X"00",X"00",X"09",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"9C",X"99",X"00",X"00",X"9C",X"99",X"00",X"00",X"9C",X"99",X"00",
		X"00",X"99",X"CC",X"00",X"00",X"09",X"CC",X"00",X"00",X"09",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"99",X"99",X"00",X"00",X"44",X"44",X"00",X"00",X"99",X"44",X"90",X"00",X"99",X"44",X"99",
		X"00",X"99",X"44",X"49",X"00",X"99",X"44",X"44",X"00",X"99",X"44",X"44",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"44",X"00",X"99",X"22",X"99",X"00",X"99",X"92",X"CC",X"00",X"99",X"99",X"CC",
		X"00",X"99",X"29",X"99",X"00",X"99",X"99",X"00",X"00",X"99",X"09",X"00",X"00",X"99",X"09",X"00",
		X"00",X"99",X"09",X"00",X"00",X"99",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"C9",X"00",X"00",X"CC",X"C9",
		X"00",X"00",X"CC",X"99",X"00",X"00",X"CC",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"99",
		X"00",X"09",X"C9",X"9C",X"00",X"09",X"CC",X"9C",X"09",X"09",X"99",X"9C",X"99",X"99",X"49",X"9C",
		X"91",X"99",X"44",X"9C",X"11",X"49",X"99",X"99",X"19",X"44",X"94",X"00",X"99",X"44",X"44",X"00",
		X"92",X"99",X"49",X"90",X"99",X"29",X"99",X"90",X"99",X"22",X"99",X"99",X"90",X"29",X"00",X"29",
		X"90",X"99",X"00",X"29",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"09",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"C9",
		X"00",X"00",X"CC",X"C9",X"00",X"00",X"CC",X"99",X"00",X"00",X"CC",X"90",X"00",X"00",X"99",X"99",
		X"00",X"00",X"99",X"9C",X"00",X"09",X"C9",X"C9",X"00",X"09",X"CC",X"99",X"00",X"99",X"99",X"9C",
		X"00",X"99",X"49",X"9C",X"00",X"49",X"44",X"99",X"00",X"49",X"99",X"99",X"00",X"44",X"94",X"00",
		X"00",X"99",X"49",X"00",X"00",X"99",X"99",X"00",X"00",X"22",X"90",X"00",X"00",X"22",X"00",X"00",
		X"00",X"22",X"00",X"00",X"00",X"29",X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"92",X"00",X"00",
		X"91",X"22",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"91",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"C9",X"C9",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"C9",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"C9",X"00",X"00",X"9C",X"CC",X"00",X"00",X"CC",X"CC",X"00",
		X"00",X"CC",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"44",X"00",X"00",X"44",X"99",X"00",
		X"00",X"99",X"44",X"00",X"00",X"29",X"99",X"00",X"00",X"99",X"22",X"00",X"00",X"19",X"22",X"00",
		X"00",X"11",X"99",X"00",X"00",X"11",X"29",X"00",X"00",X"11",X"99",X"00",X"00",X"99",X"19",X"00",
		X"00",X"11",X"99",X"00",X"00",X"19",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"99",X"C9",X"00",X"00",X"99",X"CC",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"A9",X"00",X"00",X"9C",X"29",X"00",X"00",X"9C",X"99",X"00",X"00",X"94",X"C9",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"CC",X"99",X"00",
		X"00",X"CC",X"CC",X"00",X"00",X"C9",X"99",X"00",X"00",X"CC",X"99",X"90",X"00",X"CC",X"49",X"90",
		X"00",X"99",X"49",X"90",X"00",X"99",X"99",X"90",X"00",X"94",X"44",X"90",X"00",X"94",X"44",X"00",
		X"00",X"94",X"44",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"22",X"00",X"00",X"09",X"99",X"00",
		X"00",X"09",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"C9",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"CC",X"99",X"00",X"00",X"CC",X"99",X"00",X"00",X"CC",X"9C",X"00",
		X"00",X"9C",X"CC",X"00",X"00",X"9C",X"CC",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"49",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"94",X"44",X"00",X"00",X"94",X"44",X"00",
		X"00",X"94",X"99",X"00",X"00",X"94",X"99",X"00",X"00",X"94",X"44",X"00",X"00",X"94",X"99",X"00",
		X"00",X"99",X"22",X"00",X"00",X"92",X"92",X"00",X"00",X"92",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"09",X"09",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"C9",X"99",X"00",X"00",X"CC",X"9C",X"00",X"00",X"CC",X"CC",X"00",
		X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"9C",X"9C",X"00",X"00",X"99",X"99",X"00",
		X"00",X"94",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"49",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"99",X"94",X"00",
		X"00",X"92",X"99",X"00",X"00",X"22",X"22",X"00",X"00",X"29",X"99",X"00",X"00",X"22",X"19",X"00",
		X"00",X"99",X"11",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"11",X"00",X"00",X"19",X"11",X"00",
		X"00",X"99",X"11",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"9C",X"00",X"99",X"00",X"A9",X"00",
		X"DD",X"90",X"A9",X"00",X"99",X"90",X"9C",X"00",X"99",X"90",X"C9",X"00",X"F9",X"90",X"99",X"00",
		X"99",X"90",X"99",X"00",X"99",X"90",X"99",X"00",X"99",X"90",X"9C",X"00",X"99",X"90",X"C9",X"00",
		X"99",X"99",X"99",X"00",X"99",X"94",X"CC",X"00",X"F9",X"99",X"99",X"00",X"99",X"9C",X"99",X"00",
		X"99",X"CC",X"44",X"00",X"DD",X"CC",X"44",X"00",X"99",X"99",X"99",X"00",X"99",X"90",X"99",X"00",
		X"F9",X"90",X"44",X"00",X"99",X"90",X"99",X"00",X"99",X"90",X"22",X"00",X"99",X"90",X"92",X"00",
		X"99",X"90",X"22",X"00",X"99",X"90",X"99",X"00",X"99",X"90",X"99",X"00",X"99",X"90",X"22",X"00",
		X"99",X"90",X"99",X"00",X"99",X"99",X"11",X"00",X"00",X"91",X"11",X"00",X"00",X"99",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"CC",X"00",X"00",X"09",X"C2",X"00",X"00",X"09",X"99",X"00",
		X"00",X"09",X"DD",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"09",X"99",X"00",X"00",X"94",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"9C",X"99",X"00",
		X"00",X"9C",X"99",X"00",X"00",X"9C",X"DD",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"F9",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"91",X"11",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"C9",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"CC",X"99",X"00",X"00",X"CC",X"99",X"00",X"00",X"CC",X"9C",X"00",
		X"00",X"9C",X"CC",X"00",X"00",X"9C",X"CC",X"00",X"00",X"99",X"CC",X"90",X"00",X"99",X"C9",X"90",
		X"00",X"49",X"99",X"90",X"00",X"44",X"99",X"90",X"00",X"44",X"44",X"90",X"00",X"99",X"44",X"00",
		X"00",X"99",X"44",X"00",X"00",X"99",X"44",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"44",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"99",X"00",
		X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"00",
		X"00",X"99",X"92",X"00",X"00",X"91",X"99",X"00",X"00",X"91",X"09",X"00",X"00",X"09",X"09",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"AA",X"00",X"00",X"99",X"99",X"40",
		X"00",X"9C",X"99",X"70",X"00",X"9C",X"AA",X"00",X"00",X"9C",X"99",X"00",X"00",X"99",X"CC",X"00",
		X"00",X"CC",X"9C",X"00",X"00",X"CC",X"99",X"00",X"00",X"CC",X"99",X"00",X"00",X"CC",X"99",X"00",
		X"00",X"9C",X"99",X"00",X"00",X"99",X"94",X"00",X"00",X"49",X"94",X"00",X"00",X"99",X"99",X"00",
		X"00",X"94",X"49",X"00",X"09",X"94",X"99",X"00",X"99",X"44",X"44",X"00",X"9C",X"44",X"44",X"00",
		X"9C",X"44",X"99",X"00",X"9C",X"99",X"44",X"00",X"99",X"22",X"99",X"99",X"00",X"92",X"92",X"19",
		X"00",X"99",X"22",X"19",X"00",X"09",X"92",X"19",X"00",X"00",X"99",X"19",X"00",X"00",X"29",X"19",
		X"00",X"00",X"29",X"19",X"00",X"00",X"99",X"99",X"00",X"00",X"91",X"00",X"00",X"00",X"99",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"C9",X"00",X"00",X"99",X"9C",X"00",
		X"00",X"9C",X"99",X"00",X"00",X"9C",X"CC",X"00",X"00",X"9C",X"CC",X"00",X"00",X"99",X"CC",X"00",
		X"00",X"CC",X"9C",X"00",X"00",X"CC",X"99",X"00",X"00",X"CC",X"99",X"00",X"00",X"C9",X"99",X"00",
		X"00",X"9C",X"99",X"99",X"00",X"99",X"99",X"CC",X"00",X"49",X"99",X"C9",X"00",X"49",X"99",X"CC",
		X"00",X"44",X"49",X"99",X"00",X"94",X"99",X"00",X"00",X"94",X"44",X"99",X"00",X"99",X"44",X"91",
		X"00",X"99",X"99",X"11",X"00",X"11",X"44",X"11",X"00",X"11",X"99",X"11",X"09",X"11",X"92",X"11",
		X"99",X"11",X"22",X"11",X"9C",X"11",X"99",X"99",X"99",X"99",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"91",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"C9",X"00",
		X"00",X"CC",X"99",X"00",X"00",X"C9",X"C9",X"00",X"00",X"CC",X"CC",X"A0",X"00",X"99",X"C9",X"00",
		X"00",X"CC",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"CC",X"99",X"00",X"00",X"9C",X"94",X"00",X"00",X"99",X"94",X"00",X"00",X"49",X"99",X"00",
		X"00",X"44",X"49",X"00",X"00",X"94",X"99",X"00",X"00",X"94",X"44",X"99",X"00",X"99",X"44",X"91",
		X"00",X"99",X"99",X"11",X"00",X"11",X"44",X"11",X"00",X"11",X"99",X"11",X"09",X"11",X"92",X"11",
		X"99",X"11",X"22",X"11",X"9C",X"11",X"99",X"99",X"99",X"99",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"91",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"90",X"00",X"00",
		X"09",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"9D",X"99",X"00",X"00",X"9D",X"D9",X"00",X"00",
		X"09",X"9D",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"D9",X"00",
		X"00",X"09",X"9D",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F9",X"F9",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"90",X"09",X"DD",X"DD",X"D9",X"09",X"99",X"99",X"99",X"09",X"99",X"99",X"99",
		X"09",X"99",X"99",X"99",X"09",X"99",X"99",X"99",X"09",X"99",X"99",X"99",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"99",X"00",X"00",X"9D",X"99",X"00",X"00",X"99",X"9D",X"00",X"00",X"9F",X"D9",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"9F",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"9D",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"9F",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"9D",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"9D",X"90",X"00",
		X"00",X"99",X"99",X"00",X"00",X"F9",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"09",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"9D",X"90",
		X"00",X"00",X"F9",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",
		X"00",X"00",X"99",X"99",X"00",X"00",X"DD",X"DD",X"00",X"09",X"9D",X"D9",X"00",X"99",X"99",X"99",
		X"00",X"9D",X"9F",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"9D",X"90",X"00",X"99",X"9D",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"D9",X"00",
		X"00",X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"9D",X"DD",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"9D",X"DD",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"09",X"99",X"90",X"00",X"09",X"99",X"90",X"00",X"99",X"99",X"99",X"00",X"9D",X"DD",X"D9",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"09",X"99",X"90",X"00",X"09",X"9F",X"90",X"00",
		X"09",X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"DD",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"9F",X"99",X"00",X"00",
		X"99",X"99",X"90",X"00",X"DD",X"DD",X"90",X"00",X"99",X"99",X"90",X"00",X"99",X"99",X"90",X"00",
		X"99",X"99",X"90",X"00",X"99",X"99",X"90",X"00",X"99",X"99",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"99",X"90",X"00",
		X"09",X"9F",X"90",X"00",X"09",X"99",X"90",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"9D",X"DD",X"D9",X"00",X"99",X"99",X"99",X"00",X"09",X"99",X"90",X"00",X"09",X"99",X"90",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"9C",X"9C",X"00",
		X"00",X"9C",X"CC",X"00",X"00",X"C9",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"EE",X"42",X"00",
		X"00",X"EE",X"42",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"9C",X"99",X"00",X"CC",X"CC",X"99",
		X"00",X"CC",X"CC",X"99",X"09",X"CC",X"99",X"99",X"09",X"C9",X"9F",X"99",X"99",X"C9",X"99",X"99",
		X"99",X"C9",X"9C",X"99",X"99",X"9C",X"9C",X"99",X"99",X"9C",X"CC",X"99",X"99",X"99",X"CC",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"EE",X"99",X"99",X"9C",X"EC",X"99",X"99",X"CC",
		X"CE",X"99",X"99",X"CE",X"EC",X"99",X"99",X"CC",X"EE",X"99",X"99",X"CE",X"EC",X"99",X"99",X"EC",
		X"CE",X"99",X"99",X"CE",X"CC",X"99",X"99",X"CC",X"CC",X"99",X"99",X"CC",X"CC",X"99",X"99",X"CC",
		X"EC",X"C9",X"99",X"CC",X"CE",X"C9",X"CC",X"E9",X"EC",X"CC",X"CC",X"C9",X"CC",X"CC",X"CE",X"99",
		X"CC",X"99",X"99",X"90",X"CC",X"99",X"9B",X"90",X"C9",X"9B",X"BB",X"90",X"C9",X"9B",X"BB",X"90",
		X"C9",X"BB",X"BB",X"90",X"C9",X"BB",X"BB",X"90",X"99",X"BB",X"BB",X"90",X"00",X"BB",X"BB",X"90",
		X"00",X"BB",X"BB",X"90",X"00",X"BB",X"BB",X"90",X"00",X"BB",X"BB",X"90",X"00",X"BB",X"BB",X"90",
		X"00",X"99",X"BB",X"90",X"00",X"E9",X"BB",X"90",X"00",X"7E",X"BB",X"00",X"00",X"77",X"BB",X"00",
		X"00",X"77",X"9B",X"00",X"00",X"77",X"BB",X"00",X"00",X"99",X"BB",X"00",X"00",X"77",X"BB",X"00",
		X"00",X"79",X"9B",X"90",X"00",X"99",X"BB",X"90",X"00",X"00",X"BB",X"90",X"00",X"00",X"99",X"90",
		X"00",X"00",X"7E",X"90",X"00",X"00",X"9E",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"95",X"00",X"99",X"00",X"95",X"00",X"99",X"00",
		X"95",X"99",X"99",X"00",X"99",X"55",X"95",X"00",X"09",X"52",X"55",X"00",X"00",X"59",X"55",X"00",
		X"99",X"52",X"99",X"00",X"55",X"55",X"00",X"00",X"99",X"55",X"99",X"00",X"99",X"99",X"95",X"00",
		X"99",X"44",X"55",X"99",X"95",X"44",X"55",X"55",X"55",X"44",X"55",X"95",X"55",X"44",X"55",X"99",
		X"95",X"95",X"55",X"90",X"99",X"95",X"95",X"90",X"00",X"95",X"55",X"90",X"00",X"99",X"55",X"90",
		X"00",X"09",X"55",X"90",X"00",X"09",X"55",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"97",X"90",
		X"00",X"00",X"99",X"00",X"00",X"00",X"59",X"00",X"00",X"09",X"99",X"90",X"00",X"99",X"55",X"90",
		X"00",X"95",X"55",X"90",X"00",X"99",X"59",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"55",X"00",X"00",X"09",X"52",X"00",X"00",X"09",X"59",X"00",X"00",X"99",X"52",X"00",X"00",
		X"55",X"55",X"00",X"00",X"99",X"55",X"90",X"00",X"99",X"95",X"99",X"00",X"99",X"95",X"99",X"09",
		X"95",X"95",X"95",X"99",X"55",X"95",X"95",X"95",X"55",X"95",X"95",X"99",X"95",X"99",X"95",X"90",
		X"99",X"99",X"55",X"90",X"00",X"95",X"55",X"90",X"00",X"55",X"95",X"99",X"00",X"59",X"55",X"97",
		X"09",X"55",X"55",X"99",X"99",X"59",X"55",X"95",X"99",X"99",X"99",X"55",X"95",X"00",X"00",X"55",
		X"95",X"00",X"00",X"59",X"55",X"00",X"00",X"99",X"95",X"00",X"00",X"99",X"95",X"00",X"00",X"09",
		X"99",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"CC",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"9A",X"00",X"00",X"99",X"92",X"00",X"00",X"99",X"C9",X"00",X"00",X"99",X"CC",X"00",
		X"00",X"CC",X"C9",X"00",X"00",X"9C",X"99",X"00",X"00",X"9C",X"99",X"00",X"00",X"9C",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"C9",X"00",X"00",X"49",X"99",X"00",X"09",X"44",X"99",X"99",
		X"09",X"44",X"99",X"9D",X"09",X"94",X"49",X"9D",X"09",X"99",X"44",X"9D",X"09",X"79",X"94",X"9D",
		X"09",X"77",X"94",X"9D",X"09",X"99",X"99",X"9D",X"09",X"92",X"92",X"9D",X"09",X"99",X"22",X"9D",
		X"09",X"99",X"22",X"9D",X"09",X"92",X"22",X"9D",X"09",X"92",X"22",X"9D",X"09",X"99",X"29",X"99",
		X"00",X"09",X"99",X"00",X"00",X"09",X"11",X"00",X"00",X"09",X"11",X"00",X"00",X"09",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"C9",X"00",X"00",X"99",X"99",X"00",
		X"00",X"9C",X"AA",X"00",X"00",X"9C",X"A2",X"00",X"00",X"9C",X"99",X"00",X"00",X"99",X"CC",X"00",
		X"00",X"CC",X"9C",X"00",X"00",X"CC",X"99",X"00",X"00",X"CC",X"99",X"00",X"00",X"CC",X"99",X"00",
		X"00",X"9C",X"99",X"00",X"00",X"99",X"90",X"00",X"99",X"49",X"99",X"90",X"99",X"94",X"99",X"D9",
		X"99",X"94",X"99",X"D9",X"99",X"44",X"49",X"D9",X"99",X"44",X"94",X"D9",X"99",X"44",X"44",X"D9",
		X"99",X"99",X"44",X"D9",X"99",X"99",X"99",X"99",X"99",X"99",X"22",X"91",X"99",X"92",X"22",X"11",
		X"99",X"92",X"22",X"19",X"99",X"22",X"99",X"19",X"99",X"22",X"99",X"99",X"00",X"22",X"09",X"90",
		X"00",X"99",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"CC",X"9C",X"A9",X"00",X"C9",X"9C",X"A2",X"00",X"C9",X"9C",X"99",X"00",X"C9",X"99",X"CC",X"00",
		X"99",X"CC",X"9C",X"00",X"94",X"CC",X"99",X"00",X"99",X"CC",X"99",X"00",X"09",X"9C",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"49",X"90",X"00",X"00",X"44",X"90",X"00",X"00",X"44",X"90",X"00",
		X"00",X"99",X"99",X"00",X"00",X"94",X"49",X"00",X"00",X"44",X"94",X"00",X"00",X"44",X"44",X"00",
		X"00",X"99",X"44",X"00",X"00",X"99",X"99",X"99",X"00",X"99",X"22",X"91",X"00",X"92",X"22",X"11",
		X"00",X"92",X"22",X"19",X"00",X"22",X"99",X"19",X"00",X"22",X"09",X"99",X"00",X"22",X"09",X"90",
		X"00",X"99",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"09",X"99",X"00",X"00",X"99",X"99",X"00",X"50",X"99",X"99",X"05",X"55",X"9C",X"9C",X"05",
		X"00",X"9C",X"CC",X"00",X"00",X"F9",X"99",X"00",X"00",X"F9",X"FF",X"00",X"00",X"FF",X"FF",X"0A",
		X"30",X"FF",X"99",X"00",X"00",X"9F",X"99",X"00",X"00",X"99",X"FF",X"00",X"00",X"CC",X"99",X"00",
		X"00",X"9C",X"CC",X"90",X"09",X"99",X"CC",X"99",X"09",X"99",X"99",X"99",X"99",X"CC",X"99",X"99",
		X"99",X"CC",X"49",X"99",X"99",X"9C",X"94",X"99",X"99",X"9C",X"49",X"99",X"99",X"99",X"44",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"EE",X"99",X"99",X"CC",X"EC",X"99",X"99",X"CC",
		X"CE",X"99",X"49",X"CE",X"EC",X"99",X"49",X"CC",X"99",X"99",X"49",X"99",X"90",X"99",X"99",X"90",
		X"09",X"99",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"90",X"99",X"09",X"90",X"90",X"00",
		X"00",X"09",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"94",X"94",X"00",
		X"00",X"94",X"44",X"00",X"00",X"44",X"A9",X"00",X"00",X"49",X"AA",X"00",X"00",X"99",X"99",X"00",
		X"00",X"9A",X"AA",X"00",X"00",X"4A",X"44",X"00",X"00",X"44",X"94",X"99",X"00",X"94",X"44",X"99",
		X"00",X"99",X"49",X"99",X"09",X"9F",X"99",X"99",X"09",X"9F",X"FF",X"99",X"99",X"99",X"99",X"99",
		X"99",X"49",X"F9",X"99",X"99",X"99",X"F9",X"99",X"99",X"94",X"94",X"99",X"99",X"99",X"44",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"EE",X"99",X"99",X"9C",X"EC",X"99",X"99",X"CC",
		X"CE",X"99",X"99",X"CE",X"EC",X"99",X"99",X"CC",X"EE",X"99",X"99",X"CE",X"EC",X"99",X"99",X"EC",
		X"CE",X"99",X"99",X"CE",X"CC",X"99",X"99",X"CC",X"CC",X"99",X"99",X"CC",X"CC",X"99",X"99",X"CC",
		X"EC",X"C9",X"99",X"CC",X"CE",X"C9",X"CC",X"E9",X"CC",X"CC",X"CC",X"C9",X"CC",X"CC",X"CE",X"99",
		X"CC",X"99",X"99",X"90",X"CC",X"99",X"94",X"90",X"C9",X"9F",X"F4",X"90",X"C9",X"9F",X"FF",X"90",
		X"C9",X"F4",X"F4",X"90",X"C9",X"F4",X"94",X"99",X"99",X"4F",X"FF",X"F9",X"FF",X"4F",X"FF",X"F9",
		X"99",X"99",X"99",X"99",X"09",X"EE",X"CE",X"90",X"00",X"EC",X"CE",X"90",X"00",X"CC",X"CE",X"90",
		X"00",X"CE",X"EC",X"00",X"00",X"EC",X"CE",X"00",X"00",X"CE",X"CE",X"99",X"00",X"EC",X"EC",X"E9",
		X"99",X"EC",X"CE",X"E9",X"B9",X"CE",X"99",X"CC",X"1B",X"EC",X"09",X"99",X"BB",X"99",X"00",X"BB",
		X"BB",X"BB",X"99",X"B9",X"BB",X"BB",X"B9",X"99",X"99",X"B9",X"99",X"9B",X"99",X"99",X"9B",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"99",X"BB",X"BB",X"9B",X"BB",X"9B",X"99",X"BB",X"99",X"BB",X"9B",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"77",
		X"00",X"90",X"00",X"77",X"00",X"90",X"09",X"99",X"02",X"90",X"99",X"BB",X"22",X"00",X"9E",X"BB",
		X"22",X"99",X"EE",X"BB",X"22",X"CC",X"99",X"99",X"22",X"CC",X"47",X"45",X"02",X"C9",X"47",X"45",
		X"00",X"99",X"47",X"45",X"00",X"90",X"47",X"45",X"00",X"90",X"47",X"45",X"00",X"90",X"47",X"45",
		X"00",X"90",X"47",X"45",X"00",X"90",X"47",X"45",X"00",X"90",X"47",X"45",X"00",X"90",X"47",X"45",
		X"00",X"90",X"47",X"47",X"00",X"90",X"97",X"47",X"00",X"90",X"99",X"47",X"00",X"00",X"09",X"99",
		X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"09",
		X"00",X"00",X"BA",X"99",X"00",X"90",X"55",X"9A",X"00",X"99",X"BB",X"99",X"00",X"99",X"99",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"77",
		X"00",X"90",X"00",X"77",X"00",X"90",X"09",X"99",X"02",X"90",X"99",X"BB",X"22",X"00",X"9E",X"BB",
		X"22",X"99",X"99",X"99",X"22",X"CC",X"47",X"45",X"22",X"CC",X"47",X"45",X"02",X"C9",X"47",X"45",
		X"00",X"99",X"47",X"45",X"00",X"90",X"47",X"45",X"00",X"90",X"47",X"45",X"00",X"90",X"47",X"45",
		X"00",X"90",X"47",X"45",X"00",X"90",X"47",X"45",X"00",X"90",X"47",X"45",X"00",X"90",X"47",X"47",
		X"00",X"90",X"97",X"47",X"09",X"90",X"99",X"47",X"09",X"90",X"09",X"99",X"09",X"00",X"00",X"59",
		X"09",X"90",X"00",X"99",X"09",X"99",X"00",X"90",X"99",X"AA",X"09",X"99",X"22",X"AA",X"99",X"9B",
		X"92",X"AA",X"9B",X"B5",X"99",X"99",X"9A",X"B5",X"99",X"99",X"99",X"9A",X"99",X"09",X"09",X"99",
		X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"49",X"00",X"00",X"09",X"44",X"00",
		X"00",X"99",X"AA",X"00",X"00",X"94",X"22",X"00",X"00",X"94",X"CC",X"00",X"00",X"94",X"CC",X"00",
		X"00",X"94",X"44",X"00",X"00",X"94",X"99",X"00",X"00",X"94",X"44",X"90",X"00",X"99",X"CC",X"99",
		X"00",X"AA",X"99",X"C9",X"09",X"99",X"AA",X"CC",X"99",X"99",X"AA",X"CC",X"9C",X"99",X"99",X"CC",
		X"9C",X"29",X"99",X"9C",X"9C",X"AA",X"AA",X"9C",X"99",X"AA",X"AA",X"9C",X"90",X"AA",X"AA",X"99",
		X"99",X"AA",X"22",X"44",X"95",X"22",X"AA",X"99",X"95",X"AA",X"AA",X"55",X"95",X"99",X"99",X"55",
		X"95",X"CC",X"09",X"55",X"95",X"CC",X"09",X"54",X"95",X"CC",X"09",X"54",X"95",X"99",X"09",X"54",
		X"95",X"22",X"09",X"55",X"99",X"99",X"09",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"92",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"49",X"00",X"00",X"09",X"44",X"00",
		X"00",X"99",X"44",X"00",X"00",X"9C",X"44",X"00",X"00",X"9C",X"44",X"00",X"00",X"99",X"C4",X"00",
		X"00",X"A9",X"CC",X"00",X"00",X"A9",X"CC",X"90",X"00",X"A9",X"C9",X"99",X"00",X"A9",X"99",X"C9",
		X"09",X"AA",X"9A",X"CC",X"99",X"AA",X"AA",X"CC",X"9C",X"9A",X"AA",X"CC",X"9C",X"99",X"9A",X"9C",
		X"9C",X"99",X"99",X"9C",X"99",X"AA",X"AA",X"9C",X"90",X"AA",X"AA",X"99",X"99",X"AA",X"AA",X"04",
		X"95",X"9A",X"22",X"99",X"95",X"A2",X"AA",X"55",X"95",X"AA",X"AA",X"55",X"95",X"99",X"99",X"54",
		X"95",X"9C",X"CC",X"54",X"95",X"9C",X"99",X"54",X"95",X"9C",X"09",X"55",X"95",X"9C",X"09",X"55",
		X"99",X"9C",X"09",X"99",X"00",X"99",X"09",X"00",X"00",X"92",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"49",X"00",X"00",X"09",X"44",X"00",
		X"00",X"99",X"44",X"00",X"00",X"94",X"44",X"00",X"00",X"94",X"44",X"00",X"00",X"99",X"44",X"00",
		X"00",X"99",X"44",X"00",X"00",X"A9",X"49",X"90",X"00",X"AA",X"99",X"99",X"09",X"AA",X"9A",X"C9",
		X"99",X"9A",X"AA",X"CC",X"9C",X"9A",X"AA",X"CC",X"99",X"AA",X"AA",X"CC",X"9C",X"AA",X"AA",X"9C",
		X"99",X"AA",X"99",X"9C",X"99",X"A9",X"AA",X"9C",X"90",X"AA",X"AA",X"99",X"99",X"AA",X"AA",X"00",
		X"95",X"9A",X"AA",X"99",X"95",X"AA",X"9A",X"55",X"95",X"AA",X"AA",X"55",X"95",X"99",X"99",X"55",
		X"95",X"9C",X"CC",X"54",X"95",X"9C",X"99",X"54",X"95",X"9C",X"00",X"54",X"95",X"9C",X"09",X"55",
		X"99",X"9C",X"09",X"55",X"00",X"99",X"09",X"99",X"00",X"92",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"09",X"99",X"00",X"00",X"09",X"59",X"00",X"00",X"09",X"59",X"00",X"00",X"09",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"95",X"55",X"00",X"00",X"55",X"95",X"00",
		X"00",X"99",X"99",X"00",X"00",X"9F",X"99",X"00",X"00",X"9F",X"99",X"00",X"00",X"FF",X"9F",X"00",
		X"00",X"FF",X"FF",X"00",X"00",X"99",X"FF",X"00",X"00",X"99",X"FF",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"99",X"00",X"9F",X"FF",X"92",
		X"00",X"99",X"F9",X"92",X"00",X"59",X"99",X"92",X"00",X"55",X"95",X"92",X"00",X"95",X"55",X"92",
		X"00",X"99",X"99",X"92",X"00",X"09",X"99",X"99",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"22",X"99",X"90",X"00",X"22",X"22",X"99",X"00",X"99",X"99",X"49",
		X"00",X"E9",X"00",X"49",X"00",X"CD",X"00",X"49",X"DD",X"44",X"00",X"49",X"DD",X"49",X"00",X"49",
		X"D0",X"CC",X"00",X"49",X"90",X"C9",X"09",X"49",X"9D",X"99",X"99",X"49",X"99",X"39",X"39",X"99",
		X"09",X"33",X"99",X"00",X"0D",X"33",X"9A",X"00",X"99",X"39",X"AA",X"00",X"95",X"39",X"AA",X"00",
		X"55",X"33",X"A2",X"00",X"95",X"33",X"99",X"90",X"95",X"13",X"96",X"99",X"99",X"99",X"66",X"69",
		X"66",X"69",X"66",X"99",X"22",X"22",X"22",X"95",X"22",X"22",X"22",X"95",X"22",X"99",X"22",X"99",
		X"92",X"79",X"22",X"99",X"96",X"57",X"69",X"79",X"96",X"75",X"69",X"77",X"96",X"95",X"69",X"77",
		X"99",X"77",X"99",X"74",X"00",X"77",X"09",X"49",X"00",X"79",X"00",X"99",X"00",X"99",X"00",X"90",
		X"00",X"99",X"29",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"90",X"00",X"00",X"99",X"99",X"00",
		X"00",X"E9",X"44",X"00",X"00",X"CC",X"44",X"00",X"DD",X"99",X"49",X"00",X"DD",X"94",X"59",X"00",
		X"D0",X"C9",X"99",X"00",X"90",X"C9",X"99",X"00",X"90",X"CC",X"93",X"00",X"99",X"99",X"33",X"00",
		X"09",X"39",X"39",X"00",X"09",X"33",X"99",X"00",X"00",X"39",X"9A",X"00",X"99",X"39",X"AA",X"00",
		X"95",X"33",X"AA",X"00",X"55",X"33",X"AA",X"00",X"95",X"13",X"99",X"90",X"95",X"33",X"96",X"99",
		X"99",X"99",X"66",X"69",X"66",X"69",X"66",X"99",X"22",X"92",X"22",X"95",X"22",X"99",X"22",X"95",
		X"22",X"79",X"29",X"99",X"92",X"77",X"29",X"79",X"96",X"77",X"69",X"79",X"96",X"77",X"69",X"79",
		X"96",X"77",X"69",X"59",X"99",X"79",X"99",X"99",X"00",X"99",X"00",X"90",X"00",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"E9",X"00",
		X"00",X"09",X"E9",X"00",X"00",X"9E",X"EE",X"00",X"00",X"E9",X"EE",X"00",X"00",X"EE",X"EE",X"00",
		X"00",X"EE",X"E9",X"00",X"00",X"9E",X"EE",X"00",X"00",X"99",X"EE",X"00",X"00",X"E9",X"9E",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"E9",X"00",X"00",X"99",X"EE",X"00",
		X"00",X"99",X"E9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"E9",X"00",X"00",X"09",X"E9",X"00",
		X"00",X"99",X"EE",X"00",X"00",X"9E",X"EE",X"00",X"00",X"E9",X"EE",X"00",X"00",X"EE",X"E9",X"00",
		X"00",X"9E",X"EE",X"00",X"00",X"99",X"EE",X"00",X"00",X"99",X"9E",X"00",X"00",X"E9",X"99",X"00",
		X"00",X"E9",X"99",X"00",X"00",X"E9",X"99",X"00",X"00",X"EE",X"90",X"00",X"00",X"9E",X"00",X"00",
		X"00",X"9E",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"EE",X"90",X"00",
		X"00",X"EE",X"90",X"00",X"00",X"EE",X"90",X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",
		X"00",X"EE",X"90",X"00",X"00",X"EE",X"90",X"00",X"00",X"9E",X"90",X"00",X"00",X"9E",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"E9",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"9E",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"E9",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"EE",X"90",X"00",X"00",X"EE",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"44",X"09",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"90",X"99",
		X"00",X"00",X"99",X"AA",X"00",X"00",X"D9",X"AA",X"09",X"90",X"FD",X"9A",X"99",X"99",X"99",X"99",
		X"9A",X"92",X"99",X"AA",X"99",X"22",X"99",X"AA",X"9A",X"99",X"55",X"99",X"99",X"00",X"99",X"00",
		X"09",X"00",X"99",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"99",X"00",
		X"00",X"09",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"99",X"00",X"F0",X"09",X"49",X"00",X"F0",X"99",X"44",X"00",X"FF",X"94",X"99",X"00",
		X"00",X"9C",X"9C",X"00",X"00",X"99",X"9C",X"00",X"00",X"09",X"CC",X"00",X"00",X"99",X"4C",X"00",
		X"00",X"55",X"C9",X"00",X"00",X"55",X"99",X"00",X"00",X"95",X"55",X"00",X"00",X"99",X"55",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"59",X"00",X"00",X"59",X"55",X"00",
		X"00",X"99",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"22",X"00",X"00",X"09",X"22",X"00",
		X"00",X"99",X"29",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"00",X"00",
		X"00",X"90",X"99",X"00",X"00",X"90",X"29",X"00",X"00",X"90",X"29",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"0F",X"09",X"00",X"00",X"FF",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"49",X"00",X"00",X"09",X"44",X"00",
		X"00",X"09",X"94",X"00",X"00",X"09",X"49",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"99",X"00",
		X"00",X"99",X"77",X"00",X"00",X"97",X"77",X"00",X"00",X"95",X"79",X"00",X"00",X"95",X"99",X"00",
		X"00",X"95",X"95",X"00",X"00",X"97",X"97",X"00",X"00",X"99",X"77",X"00",X"00",X"09",X"77",X"00",
		X"00",X"09",X"79",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"22",X"00",X"00",X"09",X"22",X"00",
		X"00",X"09",X"22",X"00",X"00",X"09",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"29",X"00",X"00",X"E9",X"22",X"00",
		X"00",X"E9",X"99",X"00",X"00",X"E9",X"09",X"00",X"00",X"EE",X"09",X"00",X"00",X"99",X"09",X"00",
		X"09",X"99",X"00",X"00",X"09",X"94",X"90",X"00",X"09",X"44",X"90",X"00",X"99",X"49",X"99",X"00",
		X"99",X"9A",X"49",X"00",X"99",X"99",X"99",X"00",X"99",X"CC",X"C9",X"00",X"09",X"CC",X"99",X"00",
		X"09",X"44",X"90",X"00",X"99",X"44",X"90",X"00",X"99",X"99",X"99",X"00",X"99",X"29",X"22",X"00",
		X"99",X"92",X"22",X"00",X"99",X"92",X"22",X"00",X"00",X"22",X"92",X"00",X"00",X"29",X"92",X"00",
		X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"99",X"99",X"00",
		X"00",X"69",X"CC",X"00",X"00",X"66",X"CC",X"00",X"00",X"66",X"9C",X"00",X"00",X"66",X"99",X"00",
		X"00",X"96",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"19",X"00",X"00",
		X"00",X"99",X"99",X"00",X"00",X"19",X"19",X"00",X"00",X"99",X"11",X"00",X"00",X"90",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"94",X"00",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"00",X"09",X"9C",X"00",X"00",X"09",X"9C",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"9C",X"00",
		X"00",X"09",X"94",X"00",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"00",X"00",X"99",X"00",
		X"00",X"00",X"29",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"92",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"66",X"90",X"00",X"00",X"66",X"99",X"00",X"99",X"96",X"69",
		X"00",X"19",X"66",X"99",X"00",X"19",X"99",X"91",X"00",X"19",X"90",X"91",X"00",X"19",X"00",X"99",
		X"00",X"19",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"99",X"00",X"00",X"44",X"CC",X"00",X"00",X"44",X"CC",X"00",X"00",X"44",X"99",
		X"00",X"00",X"44",X"99",X"00",X"00",X"49",X"99",X"00",X"00",X"99",X"92",X"00",X"00",X"94",X"92",
		X"00",X"00",X"49",X"92",X"00",X"00",X"99",X"99",X"00",X"00",X"CC",X"99",X"00",X"09",X"99",X"99",
		X"00",X"99",X"22",X"99",X"00",X"92",X"22",X"99",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",
		X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"92",X"99",X"00",
		X"00",X"99",X"69",X"00",X"00",X"9C",X"66",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"99",X"99",X"49",X"99",X"99",X"99",X"44",X"99",
		X"09",X"CC",X"44",X"09",X"09",X"CC",X"44",X"09",X"09",X"99",X"44",X"09",X"09",X"29",X"94",X"09",
		X"09",X"09",X"94",X"09",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"00",X"09",X"90",X"00",
		X"00",X"09",X"90",X"00",X"00",X"09",X"20",X"00",X"00",X"99",X"20",X"00",X"00",X"99",X"20",X"00",
		X"00",X"29",X"20",X"00",X"00",X"22",X"20",X"00",X"00",X"92",X"20",X"00",X"00",X"99",X"90",X"00",
		X"00",X"69",X"60",X"00",X"00",X"96",X"60",X"00",X"00",X"99",X"90",X"00",X"00",X"09",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"77",X"00",X"09",X"90",X"77",X"00",X"99",X"99",X"99",X"00",X"44",X"44",X"66",X"00",
		X"99",X"99",X"66",X"00",X"9E",X"EC",X"66",X"00",X"CE",X"9C",X"99",X"99",X"9C",X"99",X"00",X"33",
		X"9C",X"C9",X"00",X"93",X"99",X"C9",X"09",X"93",X"09",X"99",X"93",X"99",X"99",X"90",X"31",X"90",
		X"95",X"90",X"93",X"90",X"99",X"90",X"99",X"90",X"99",X"99",X"00",X"90",X"99",X"CE",X"00",X"90",
		X"95",X"CE",X"00",X"99",X"95",X"9C",X"00",X"99",X"95",X"99",X"99",X"99",X"99",X"90",X"99",X"44",
		X"99",X"90",X"09",X"44",X"91",X"90",X"09",X"44",X"99",X"90",X"09",X"44",X"99",X"99",X"00",X"44",
		X"99",X"11",X"00",X"44",X"11",X"11",X"00",X"49",X"11",X"11",X"00",X"99",X"11",X"91",X"00",X"59",
		X"11",X"99",X"00",X"95",X"19",X"09",X"00",X"95",X"99",X"00",X"00",X"59",X"99",X"00",X"00",X"99",
		X"00",X"90",X"00",X"66",X"00",X"99",X"00",X"66",X"99",X"49",X"00",X"66",X"94",X"44",X"00",X"AA",
		X"99",X"99",X"00",X"AA",X"99",X"EC",X"00",X"66",X"9C",X"C9",X"00",X"66",X"99",X"C9",X"00",X"66",
		X"09",X"CC",X"00",X"99",X"09",X"99",X"09",X"90",X"99",X"CC",X"99",X"90",X"95",X"99",X"93",X"99",
		X"99",X"90",X"93",X"11",X"99",X"99",X"99",X"99",X"99",X"CE",X"00",X"90",X"95",X"CE",X"00",X"99",
		X"95",X"9C",X"00",X"99",X"95",X"99",X"99",X"99",X"99",X"90",X"99",X"44",X"99",X"90",X"09",X"44",
		X"91",X"90",X"09",X"44",X"91",X"90",X"09",X"44",X"91",X"90",X"00",X"44",X"99",X"90",X"00",X"44",
		X"09",X"00",X"00",X"49",X"09",X"00",X"00",X"99",X"09",X"00",X"00",X"99",X"09",X"00",X"00",X"79",
		X"09",X"00",X"00",X"79",X"09",X"99",X"00",X"59",X"09",X"99",X"00",X"99",X"09",X"99",X"00",X"90",
		X"00",X"00",X"99",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"9C",X"00",X"00",X"00",X"A9",X"00",
		X"00",X"00",X"29",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"C9",X"00",X"09",X"00",X"99",X"00",
		X"09",X"00",X"99",X"00",X"09",X"90",X"99",X"00",X"00",X"99",X"9C",X"00",X"00",X"94",X"C9",X"00",
		X"00",X"44",X"99",X"00",X"00",X"44",X"CC",X"00",X"00",X"94",X"99",X"00",X"00",X"99",X"44",X"90",
		X"00",X"00",X"99",X"90",X"00",X"00",X"C9",X"90",X"00",X"00",X"C9",X"90",X"00",X"00",X"C9",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"22",X"00",X"00",X"99",X"92",X"00",
		X"00",X"99",X"22",X"00",X"00",X"92",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"19",X"22",X"00",
		X"00",X"11",X"99",X"00",X"00",X"91",X"11",X"00",X"00",X"99",X"11",X"00",X"00",X"09",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"94",X"99",X"00",
		X"00",X"44",X"44",X"00",X"00",X"99",X"99",X"00",X"00",X"9A",X"C9",X"00",X"00",X"9A",X"C9",X"00",
		X"00",X"99",X"99",X"00",X"00",X"9C",X"90",X"00",X"00",X"94",X"99",X"00",X"00",X"99",X"97",X"00",
		X"00",X"99",X"97",X"00",X"00",X"97",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"79",X"79",X"00",
		X"00",X"79",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"77",X"00",X"00",X"99",X"79",X"00",
		X"00",X"90",X"9D",X"00",X"00",X"99",X"DD",X"00",X"00",X"49",X"9D",X"00",X"00",X"49",X"DD",X"00",
		X"00",X"49",X"DD",X"00",X"00",X"99",X"D9",X"00",X"00",X"49",X"DD",X"00",X"00",X"99",X"9D",X"00",
		X"00",X"90",X"99",X"00",X"00",X"90",X"09",X"00",X"00",X"90",X"99",X"00",X"00",X"90",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"91",X"00",X"00",X"99",X"91",
		X"99",X"00",X"91",X"11",X"92",X"99",X"11",X"91",X"52",X"11",X"11",X"91",X"52",X"11",X"11",X"91",
		X"99",X"99",X"11",X"19",X"00",X"00",X"11",X"91",X"00",X"00",X"99",X"19",X"00",X"00",X"00",X"91",
		X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"91",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"9C",X"90",X"00",X"00",X"CC",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"AA",X"99",X"00",X"00",X"A2",X"C9",X"00",X"00",X"99",X"C9",X"00",X"00",X"9C",X"C9",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"00",X"00",
		X"00",X"C9",X"99",X"00",X"00",X"CC",X"44",X"00",X"09",X"99",X"99",X"00",X"99",X"44",X"99",X"00",
		X"94",X"44",X"99",X"00",X"44",X"99",X"99",X"00",X"44",X"44",X"99",X"00",X"99",X"44",X"99",X"00",
		X"44",X"44",X"99",X"00",X"99",X"99",X"99",X"00",X"CC",X"22",X"99",X"00",X"CC",X"29",X"99",X"00",
		X"99",X"92",X"99",X"00",X"00",X"92",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"90",X"99",X"00",
		X"00",X"90",X"99",X"00",X"00",X"90",X"99",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"9C",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"9A",X"99",X"00",X"00",X"92",X"CC",X"00",X"00",X"99",X"9C",X"00",X"00",X"C9",X"CC",X"00",
		X"00",X"49",X"49",X"00",X"00",X"99",X"C9",X"00",X"00",X"99",X"99",X"00",X"00",X"C9",X"90",X"00",
		X"09",X"CC",X"99",X"00",X"99",X"9C",X"49",X"00",X"94",X"99",X"44",X"00",X"94",X"44",X"99",X"00",
		X"94",X"44",X"99",X"00",X"94",X"99",X"99",X"00",X"99",X"44",X"99",X"00",X"9C",X"44",X"99",X"00",
		X"9C",X"44",X"99",X"00",X"99",X"99",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"29",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"9C",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"AA",X"C9",X"00",X"00",X"2A",X"C9",X"00",X"00",X"99",X"C9",X"00",X"00",X"CC",X"99",X"00",
		X"00",X"C9",X"CC",X"00",X"00",X"99",X"CC",X"00",X"00",X"99",X"CC",X"00",X"00",X"99",X"CC",X"00",
		X"00",X"99",X"99",X"00",X"00",X"09",X"44",X"00",X"09",X"99",X"44",X"99",X"9D",X"99",X"44",X"99",
		X"9D",X"99",X"4F",X"99",X"9D",X"99",X"99",X"99",X"9D",X"CC",X"99",X"99",X"9D",X"CC",X"99",X"99",
		X"9D",X"CC",X"99",X"99",X"9D",X"99",X"99",X"99",X"9D",X"99",X"99",X"99",X"9D",X"99",X"99",X"99",
		X"9D",X"9F",X"F9",X"99",X"9D",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"09",X"90",X"22",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"99",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"CC",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"A9",X"99",X"00",X"00",X"29",X"99",X"00",X"00",X"9C",X"99",X"00",X"00",X"CC",X"99",X"00",
		X"00",X"9C",X"CC",X"00",X"00",X"99",X"C9",X"00",X"00",X"99",X"C9",X"00",X"00",X"99",X"C9",X"00",
		X"00",X"99",X"99",X"00",X"00",X"9C",X"99",X"00",X"00",X"99",X"94",X"00",X"99",X"99",X"44",X"90",
		X"D9",X"99",X"44",X"90",X"D9",X"99",X"49",X"90",X"D9",X"99",X"99",X"90",X"D9",X"99",X"99",X"90",
		X"D9",X"99",X"99",X"90",X"D9",X"99",X"99",X"90",X"D9",X"99",X"99",X"90",X"D9",X"99",X"99",X"90",
		X"D9",X"99",X"99",X"90",X"D9",X"F9",X"99",X"90",X"D9",X"99",X"99",X"90",X"99",X"99",X"99",X"90",
		X"00",X"99",X"90",X"00",X"00",X"11",X"90",X"00",X"00",X"11",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"9C",X"00",X"00",X"C9",X"CC",X"00",X"00",X"CC",X"CC",X"00",
		X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"C9",X"00",X"00",X"99",X"99",X"00",
		X"00",X"49",X"49",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"99",X"44",X"00",
		X"00",X"99",X"44",X"00",X"00",X"99",X"44",X"00",X"00",X"99",X"44",X"00",X"00",X"99",X"44",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"92",X"00",X"00",X"99",X"92",X"00",
		X"00",X"91",X"22",X"00",X"00",X"11",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"11",X"99",X"00",
		X"00",X"11",X"91",X"00",X"00",X"11",X"91",X"00",X"00",X"91",X"99",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"C9",X"99",X"00",X"00",X"CC",X"9C",X"00",
		X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"9C",X"CC",X"00",X"00",X"99",X"99",X"00",
		X"00",X"94",X"94",X"00",X"00",X"44",X"44",X"00",X"00",X"99",X"44",X"00",X"00",X"99",X"44",X"00",
		X"00",X"99",X"44",X"90",X"00",X"99",X"44",X"90",X"00",X"99",X"44",X"90",X"00",X"99",X"94",X"90",
		X"00",X"99",X"99",X"90",X"00",X"99",X"22",X"90",X"00",X"99",X"29",X"90",X"00",X"99",X"99",X"90",
		X"00",X"99",X"91",X"90",X"00",X"99",X"11",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"11",X"00",
		X"00",X"99",X"11",X"00",X"00",X"99",X"11",X"00",X"00",X"09",X"91",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"99",X"CC",X"00",X"00",X"99",X"9C",X"00",X"00",X"99",X"9C",X"00",
		X"00",X"09",X"9C",X"00",X"00",X"09",X"9C",X"00",X"00",X"09",X"CC",X"00",X"00",X"09",X"CC",X"00",
		X"00",X"09",X"CC",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",
		X"00",X"99",X"44",X"99",X"00",X"44",X"CC",X"C9",X"99",X"44",X"99",X"C9",X"19",X"44",X"94",X"C9",
		X"11",X"44",X"44",X"C9",X"99",X"99",X"99",X"99",X"92",X"99",X"44",X"00",X"22",X"44",X"94",X"00",
		X"22",X"44",X"99",X"99",X"22",X"99",X"99",X"91",X"92",X"29",X"99",X"91",X"99",X"99",X"00",X"11",
		X"09",X"00",X"00",X"11",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"CC",X"00",X"00",X"99",X"9C",X"00",
		X"00",X"99",X"9C",X"00",X"00",X"99",X"9C",X"00",X"00",X"09",X"9C",X"00",X"00",X"09",X"CC",X"00",
		X"00",X"09",X"CC",X"00",X"00",X"09",X"CC",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"99",X"99",
		X"00",X"00",X"99",X"9C",X"00",X"99",X"44",X"9C",X"00",X"44",X"CC",X"CC",X"00",X"44",X"99",X"C9",
		X"00",X"44",X"94",X"C9",X"00",X"44",X"44",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"00",
		X"00",X"44",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"29",X"00",X"00",
		X"00",X"99",X"00",X"00",X"09",X"92",X"00",X"00",X"99",X"22",X"00",X"00",X"19",X"29",X"00",X"00",
		X"11",X"99",X"00",X"00",X"11",X"99",X"00",X"00",X"99",X"11",X"00",X"00",X"99",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"9C",X"99",X"00",X"00",X"CC",X"99",X"00",X"00",X"CC",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"A9",X"C9",X"00",X"00",X"99",X"C9",X"00",X"00",X"9C",X"C9",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"9F",X"CC",X"00",
		X"00",X"99",X"CC",X"00",X"00",X"9C",X"9C",X"00",X"09",X"99",X"CC",X"00",X"09",X"94",X"CC",X"00",
		X"09",X"94",X"99",X"00",X"09",X"99",X"99",X"00",X"09",X"44",X"49",X"00",X"09",X"44",X"49",X"00",
		X"00",X"44",X"49",X"00",X"00",X"99",X"99",X"00",X"00",X"22",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"92",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"C9",X"00",
		X"00",X"99",X"C9",X"00",X"00",X"99",X"C9",X"00",X"00",X"CC",X"CC",X"00",X"00",X"4C",X"CC",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"9C",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"9C",X"99",X"00",X"00",X"CC",X"C9",X"00",X"00",X"CC",X"CC",X"00",
		X"00",X"99",X"CC",X"00",X"00",X"99",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"99",X"44",X"00",
		X"00",X"44",X"99",X"00",X"00",X"99",X"92",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"91",X"00",
		X"00",X"99",X"11",X"00",X"00",X"92",X"11",X"00",X"00",X"99",X"11",X"00",X"00",X"91",X"99",X"00",
		X"00",X"99",X"11",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"9C",X"00",X"00",X"C9",X"CC",X"00",X"00",X"CC",X"CC",X"00",
		X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"C9",X"C9",X"00",X"00",X"99",X"99",X"00",
		X"00",X"44",X"49",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"94",X"00",X"00",X"44",X"44",X"00",X"00",X"49",X"99",X"00",
		X"00",X"99",X"29",X"00",X"00",X"22",X"22",X"00",X"00",X"99",X"92",X"00",X"00",X"91",X"22",X"00",
		X"00",X"11",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"11",X"99",X"00",X"00",X"11",X"91",X"00",
		X"00",X"11",X"99",X"00",X"00",X"91",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"9C",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"CC",X"00",X"00",X"99",X"CC",X"00",X"00",X"C9",X"CC",X"00",
		X"00",X"CC",X"C9",X"00",X"00",X"CC",X"C9",X"00",X"00",X"99",X"99",X"00",X"00",X"94",X"99",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"49",X"00",X"00",X"44",X"49",X"00",
		X"00",X"99",X"49",X"00",X"00",X"99",X"49",X"00",X"00",X"44",X"49",X"00",X"00",X"99",X"49",X"00",
		X"00",X"22",X"99",X"00",X"00",X"29",X"29",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"99",X"00",
		X"00",X"90",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"DD",X"9C",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"CC",X"00",X"99",X"99",X"9C",X"00",
		X"99",X"99",X"94",X"00",X"99",X"99",X"44",X"00",X"9F",X"9C",X"9C",X"00",X"99",X"99",X"9C",X"00",
		X"99",X"99",X"C9",X"00",X"99",X"49",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"94",X"00",
		X"99",X"94",X"49",X"00",X"DD",X"94",X"44",X"00",X"99",X"99",X"99",X"00",X"99",X"94",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"92",X"00",X"99",X"09",X"22",X"00",X"99",X"09",X"22",X"00",
		X"9F",X"09",X"22",X"00",X"99",X"09",X"92",X"00",X"99",X"09",X"29",X"00",X"99",X"09",X"22",X"00",
		X"99",X"99",X"99",X"00",X"99",X"91",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"99",X"99",X"00",
		X"00",X"00",X"90",X"00",X"00",X"99",X"C9",X"00",X"00",X"99",X"AC",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"DD",X"00",X"00",X"99",X"99",X"00",X"00",X"C9",X"99",X"00",X"00",X"C9",X"F9",X"00",
		X"00",X"99",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"49",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"C9",X"F9",X"00",X"00",X"C9",X"99",X"00",
		X"00",X"CC",X"99",X"00",X"00",X"CC",X"DD",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"99",X"00",
		X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",
		X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"F9",X"00",X"00",X"09",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"11",X"11",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"9C",X"00",X"00",X"C9",X"CC",X"00",X"00",X"CC",X"CC",X"00",
		X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"C9",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"94",X"00",X"00",X"49",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"99",X"44",X"00",X"00",X"99",X"44",X"00",X"00",X"94",X"44",X"00",X"00",X"94",X"44",X"00",
		X"00",X"44",X"99",X"00",X"00",X"99",X"22",X"00",X"00",X"92",X"22",X"00",X"00",X"92",X"92",X"00",
		X"00",X"92",X"22",X"00",X"00",X"92",X"22",X"00",X"00",X"92",X"22",X"00",X"00",X"99",X"22",X"00",
		X"00",X"99",X"22",X"00",X"00",X"19",X"99",X"00",X"00",X"11",X"11",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"CC",X"00",X"00",X"99",X"9C",X"00",X"00",X"99",X"9C",X"00",
		X"00",X"CC",X"97",X"00",X"00",X"9C",X"99",X"00",X"00",X"CC",X"CC",X"00",X"00",X"9C",X"CC",X"00",
		X"00",X"CC",X"C9",X"00",X"00",X"CC",X"94",X"00",X"00",X"CC",X"94",X"00",X"00",X"CC",X"94",X"00",
		X"00",X"C9",X"49",X"00",X"00",X"CC",X"49",X"00",X"00",X"99",X"99",X"00",X"09",X"44",X"90",X"00",
		X"99",X"44",X"00",X"00",X"94",X"44",X"99",X"00",X"49",X"44",X"49",X"00",X"44",X"44",X"44",X"00",
		X"CC",X"44",X"44",X"00",X"C9",X"94",X"49",X"00",X"99",X"99",X"99",X"00",X"00",X"22",X"91",X"00",
		X"00",X"22",X"91",X"00",X"00",X"92",X"91",X"00",X"00",X"99",X"91",X"00",X"00",X"09",X"91",X"00",
		X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"99",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"CC",X"90",X"00",X"00",X"9C",X"99",X"00",X"00",X"CC",X"CC",X"00",X"00",X"9C",X"CC",X"00",
		X"00",X"CC",X"C9",X"00",X"00",X"CC",X"90",X"00",X"00",X"C9",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"C9",X"00",X"90",X"00",X"CC",X"99",X"99",X"00",X"99",X"44",X"CC",X"00",X"44",X"94",X"C9",
		X"00",X"44",X"99",X"99",X"00",X"44",X"99",X"00",X"00",X"44",X"49",X"90",X"00",X"99",X"44",X"90",
		X"00",X"11",X"44",X"90",X"00",X"11",X"49",X"90",X"00",X"11",X"99",X"90",X"99",X"11",X"22",X"90",
		X"CC",X"11",X"22",X"90",X"CC",X"11",X"99",X"90",X"99",X"99",X"00",X"00",X"09",X"11",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"CC",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"C9",X"00",X"00",X"CC",X"C9",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"94",X"00",X"00",X"99",X"99",X"00",X"00",X"94",X"99",X"00",
		X"00",X"94",X"94",X"00",X"00",X"99",X"44",X"00",X"00",X"CC",X"99",X"00",X"00",X"99",X"90",X"00",
		X"00",X"44",X"90",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"49",X"90",X"00",X"99",X"44",X"90",
		X"00",X"11",X"44",X"90",X"00",X"11",X"49",X"90",X"00",X"11",X"99",X"90",X"99",X"11",X"22",X"90",
		X"CC",X"11",X"22",X"90",X"CC",X"11",X"99",X"90",X"99",X"99",X"00",X"00",X"09",X"11",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9F",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9D",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"9F",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9D",X"00",X"00",X"00",
		X"D9",X"00",X"00",X"00",X"D9",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"9F",X"00",X"00",X"99",X"D9",X"00",X"00",X"09",X"9D",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"F9",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"D9",X"00",X"00",X"09",X"9D",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"09",X"99",X"99",X"00",
		X"99",X"9F",X"99",X"00",X"DD",X"DD",X"DD",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"90",X"00",X"00",X"DD",X"D0",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"DD",X"90",X"00",
		X"00",X"9D",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"09",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"D9",X"00",X"00",
		X"09",X"D9",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"D9",X"00",X"00",X"00",X"9D",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"9F",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"9D",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"D9",X"00",X"00",X"00",X"9D",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",
		X"00",X"00",X"99",X"D9",X"00",X"09",X"99",X"99",X"00",X"99",X"DD",X"99",X"00",X"99",X"9D",X"99",
		X"00",X"D9",X"99",X"99",X"00",X"DD",X"99",X"99",X"00",X"9D",X"9D",X"90",X"00",X"99",X"DD",X"00",
		X"00",X"99",X"D9",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"09",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"DD",X"DD",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"F9",X"F9",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"F9",X"F9",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"DD",X"DD",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"F9",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"F9",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"DD",X"DD",X"00",X"00",
		X"99",X"99",X"00",X"00",X"FF",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"9D",X"DD",X"00",X"00",X"99",X"99",X"00",X"00",
		X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"F9",X"00",X"00",X"99",X"99",X"00",X"00",X"DD",X"DD",X"00",X"00",
		X"9F",X"9F",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"DD",X"DD",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"9D",X"DD",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"DD",X"DD",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"C9",X"C9",X"00",
		X"00",X"CC",X"C9",X"00",X"00",X"99",X"9C",X"00",X"00",X"99",X"99",X"00",X"00",X"2A",X"AE",X"00",
		X"00",X"22",X"2E",X"00",X"00",X"CC",X"CC",X"00",X"00",X"C9",X"CC",X"00",X"00",X"CC",X"CC",X"90",
		X"09",X"CC",X"CC",X"90",X"99",X"99",X"CC",X"99",X"99",X"F9",X"9C",X"99",X"99",X"99",X"9C",X"99",
		X"99",X"9F",X"CC",X"99",X"99",X"99",X"C9",X"99",X"99",X"CC",X"C9",X"99",X"99",X"CC",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"C9",X"C9",X"99",X"99",X"CE",X"EC",X"99",X"99",X"EE",
		X"EE",X"94",X"99",X"CC",X"EC",X"94",X"99",X"EE",X"CE",X"94",X"99",X"CC",X"EC",X"99",X"99",X"EC",
		X"EE",X"99",X"99",X"CC",X"EC",X"99",X"99",X"C9",X"CE",X"99",X"99",X"C9",X"EC",X"9C",X"CC",X"99",
		X"EE",X"CC",X"CC",X"90",X"CC",X"99",X"CC",X"90",X"CE",X"CC",X"EC",X"00",X"CC",X"CC",X"CE",X"00",
		X"CC",X"CC",X"99",X"00",X"CC",X"99",X"BB",X"00",X"C9",X"BB",X"BB",X"00",X"C9",X"BB",X"BB",X"00",
		X"C9",X"BB",X"BB",X"00",X"C9",X"BB",X"BB",X"00",X"99",X"BB",X"BB",X"00",X"99",X"BB",X"BB",X"00",
		X"9B",X"BB",X"BB",X"00",X"9B",X"B9",X"BB",X"00",X"99",X"B9",X"BB",X"00",X"09",X"B9",X"BB",X"00",
		X"99",X"B9",X"BB",X"00",X"99",X"99",X"BB",X"00",X"99",X"99",X"BB",X"00",X"97",X"79",X"BB",X"00",
		X"97",X"79",X"BB",X"00",X"97",X"79",X"BB",X"00",X"99",X"99",X"BB",X"00",X"99",X"99",X"BB",X"00",
		X"09",X"90",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"E7",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"90",X"00",X"99",X"00",X"99",X"00",
		X"95",X"99",X"59",X"00",X"55",X"59",X"59",X"00",X"57",X"25",X"59",X"00",X"97",X"9E",X"99",X"00",
		X"99",X"2E",X"90",X"00",X"55",X"E5",X"00",X"00",X"55",X"55",X"99",X"00",X"55",X"55",X"55",X"00",
		X"55",X"95",X"99",X"99",X"55",X"45",X"99",X"59",X"55",X"44",X"99",X"55",X"55",X"44",X"59",X"95",
		X"59",X"45",X"55",X"95",X"99",X"55",X"55",X"95",X"00",X"55",X"55",X"95",X"00",X"55",X"55",X"95",
		X"00",X"55",X"55",X"99",X"00",X"99",X"55",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",
		X"00",X"99",X"95",X"00",X"00",X"97",X"55",X"00",X"00",X"99",X"55",X"00",X"00",X"59",X"59",X"00",
		X"00",X"55",X"99",X"00",X"00",X"55",X"99",X"00",X"00",X"95",X"09",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",
		X"99",X"59",X"00",X"00",X"95",X"25",X"00",X"00",X"57",X"25",X"00",X"99",X"99",X"25",X"00",X"95",
		X"55",X"55",X"00",X"95",X"55",X"59",X"00",X"95",X"55",X"59",X"99",X"95",X"55",X"59",X"55",X"95",
		X"55",X"59",X"55",X"55",X"55",X"59",X"99",X"59",X"55",X"59",X"99",X"99",X"59",X"55",X"99",X"00",
		X"99",X"95",X"59",X"00",X"00",X"55",X"55",X"00",X"00",X"55",X"55",X"99",X"99",X"55",X"55",X"79",
		X"97",X"95",X"55",X"97",X"77",X"99",X"55",X"99",X"99",X"09",X"99",X"59",X"99",X"00",X"00",X"55",
		X"95",X"00",X"00",X"55",X"55",X"00",X"00",X"55",X"59",X"00",X"00",X"55",X"59",X"00",X"00",X"55",
		X"99",X"00",X"00",X"59",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"CC",X"A9",X"00",X"00",X"C9",X"A9",X"00",X"00",X"CC",X"9C",X"00",X"00",X"99",X"CC",X"00",
		X"00",X"CC",X"CC",X"00",X"00",X"44",X"99",X"00",X"00",X"C9",X"99",X"00",X"00",X"CC",X"99",X"00",
		X"00",X"CC",X"90",X"00",X"00",X"9C",X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"99",X"99",X"00",
		X"99",X"49",X"99",X"90",X"9F",X"44",X"99",X"90",X"99",X"44",X"49",X"90",X"99",X"94",X"44",X"90",
		X"99",X"99",X"44",X"90",X"99",X"99",X"99",X"90",X"99",X"22",X"22",X"90",X"99",X"22",X"29",X"90",
		X"9F",X"92",X"29",X"90",X"99",X"99",X"99",X"90",X"99",X"29",X"99",X"90",X"99",X"99",X"99",X"00",
		X"00",X"19",X"99",X"00",X"00",X"19",X"11",X"00",X"00",X"19",X"11",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"C9",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"C9",X"CC",X"00",X"00",X"9C",X"CC",X"00",
		X"00",X"CC",X"C9",X"00",X"00",X"44",X"99",X"00",X"00",X"C9",X"90",X"00",X"00",X"CC",X"90",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"99",X"99",X"99",X"00",X"99",X"49",X"99",X"00",
		X"94",X"44",X"99",X"00",X"44",X"44",X"99",X"00",X"44",X"44",X"49",X"00",X"99",X"44",X"44",X"00",
		X"44",X"44",X"44",X"00",X"99",X"99",X"99",X"90",X"CC",X"99",X"29",X"90",X"CC",X"99",X"22",X"90",
		X"99",X"29",X"22",X"90",X"99",X"22",X"92",X"00",X"99",X"22",X"22",X"00",X"00",X"99",X"92",X"00",
		X"00",X"90",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"99",X"99",X"90",X"00",
		X"C9",X"C9",X"90",X"00",X"C9",X"99",X"99",X"00",X"99",X"C9",X"CC",X"00",X"99",X"9C",X"CC",X"00",
		X"44",X"CC",X"C9",X"00",X"44",X"44",X"99",X"00",X"44",X"C9",X"90",X"00",X"94",X"CC",X"90",X"00",
		X"99",X"CC",X"00",X"00",X"09",X"9C",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"49",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"44",X"90",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"49",X"00",
		X"00",X"44",X"49",X"00",X"00",X"99",X"99",X"90",X"00",X"99",X"29",X"90",X"00",X"99",X"22",X"90",
		X"00",X"29",X"22",X"90",X"00",X"22",X"92",X"00",X"00",X"22",X"22",X"00",X"00",X"99",X"92",X"00",
		X"00",X"90",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"99",X"00",X"00",
		X"05",X"99",X"90",X"00",X"05",X"99",X"99",X"55",X"55",X"99",X"99",X"50",X"50",X"C9",X"C9",X"00",
		X"00",X"CC",X"C9",X"00",X"00",X"9F",X"9C",X"00",X"A0",X"9F",X"F9",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"99",X"99",X"00",X"00",X"CC",X"9C",X"00",
		X"09",X"CC",X"C9",X"00",X"99",X"CC",X"C9",X"90",X"99",X"9C",X"99",X"90",X"99",X"99",X"99",X"99",
		X"99",X"99",X"9C",X"99",X"99",X"CC",X"99",X"99",X"99",X"CC",X"49",X"99",X"99",X"CC",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"CC",X"99",X"99",X"CE",X"EC",X"99",X"99",X"EE",
		X"CC",X"94",X"99",X"CC",X"EC",X"94",X"99",X"EE",X"99",X"94",X"99",X"99",X"09",X"99",X"99",X"09",
		X"00",X"00",X"99",X"90",X"90",X"00",X"00",X"00",X"99",X"09",X"00",X"00",X"00",X"09",X"09",X"90",
		X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"49",X"49",X"00",
		X"00",X"44",X"49",X"00",X"00",X"99",X"94",X"00",X"00",X"9A",X"99",X"00",X"00",X"A9",X"A9",X"00",
		X"00",X"AA",X"AA",X"00",X"00",X"A4",X"AA",X"00",X"00",X"49",X"44",X"00",X"00",X"44",X"49",X"90",
		X"09",X"94",X"99",X"90",X"99",X"99",X"F9",X"99",X"99",X"FF",X"99",X"99",X"99",X"99",X"94",X"99",
		X"99",X"FF",X"44",X"99",X"99",X"9F",X"49",X"99",X"99",X"49",X"49",X"99",X"99",X"44",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"C9",X"C9",X"99",X"99",X"CE",X"EC",X"99",X"99",X"EE",
		X"EE",X"94",X"99",X"CC",X"EC",X"94",X"99",X"EE",X"CE",X"94",X"99",X"CC",X"EC",X"99",X"99",X"EC",
		X"EE",X"99",X"99",X"CC",X"EC",X"99",X"99",X"C9",X"CE",X"99",X"99",X"C9",X"EC",X"9C",X"CC",X"99",
		X"EE",X"CC",X"CC",X"90",X"CC",X"99",X"CC",X"90",X"CC",X"CC",X"EC",X"00",X"CC",X"CC",X"CE",X"00",
		X"CC",X"CC",X"99",X"00",X"CC",X"99",X"4F",X"00",X"C9",X"F4",X"4F",X"00",X"C9",X"FF",X"FF",X"00",
		X"C9",X"4F",X"44",X"00",X"C9",X"49",X"44",X"00",X"99",X"FF",X"FF",X"00",X"F9",X"FF",X"FF",X"00",
		X"99",X"99",X"99",X"00",X"9E",X"EC",X"EE",X"00",X"9C",X"CC",X"CC",X"00",X"99",X"EE",X"CE",X"00",
		X"09",X"CE",X"EE",X"00",X"00",X"EC",X"CC",X"00",X"00",X"CE",X"CE",X"00",X"00",X"EC",X"EC",X"00",
		X"09",X"C9",X"CE",X"90",X"99",X"99",X"EC",X"90",X"B1",X"90",X"9C",X"99",X"BB",X"90",X"99",X"B9",
		X"BB",X"99",X"00",X"99",X"BB",X"B9",X"99",X"1B",X"9B",X"99",X"BB",X"BB",X"99",X"9B",X"BB",X"BB",
		X"99",X"BB",X"BB",X"B9",X"99",X"B9",X"99",X"B9",X"BB",X"99",X"99",X"99",X"99",X"BB",X"BB",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"09",X"77",
		X"00",X"00",X"99",X"77",X"99",X"00",X"9E",X"99",X"9C",X"00",X"EE",X"BB",X"9C",X"00",X"EE",X"BB",
		X"9C",X"99",X"EE",X"BB",X"9C",X"97",X"99",X"99",X"9C",X"99",X"45",X"45",X"9C",X"90",X"45",X"45",
		X"9C",X"00",X"45",X"45",X"99",X"00",X"45",X"45",X"09",X"00",X"45",X"45",X"09",X"00",X"45",X"45",
		X"09",X"00",X"45",X"45",X"09",X"00",X"45",X"45",X"99",X"00",X"45",X"45",X"96",X"00",X"47",X"45",
		X"99",X"00",X"47",X"47",X"9A",X"00",X"47",X"49",X"9A",X"00",X"47",X"99",X"99",X"00",X"99",X"90",
		X"09",X"00",X"95",X"90",X"99",X"00",X"99",X"00",X"9A",X"00",X"99",X"00",X"9A",X"00",X"90",X"99",
		X"9A",X"00",X"99",X"AB",X"99",X"00",X"A9",X"55",X"99",X"00",X"99",X"BB",X"99",X"00",X"90",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"09",X"77",
		X"00",X"00",X"99",X"77",X"99",X"00",X"9E",X"99",X"9C",X"00",X"EE",X"BB",X"9C",X"00",X"EE",X"BB",
		X"9C",X"99",X"99",X"99",X"9C",X"97",X"45",X"45",X"9C",X"99",X"45",X"45",X"9C",X"90",X"45",X"45",
		X"9C",X"00",X"45",X"45",X"99",X"00",X"45",X"45",X"09",X"00",X"45",X"45",X"09",X"00",X"45",X"45",
		X"09",X"00",X"45",X"45",X"09",X"00",X"45",X"45",X"09",X"00",X"47",X"45",X"99",X"00",X"47",X"47",
		X"96",X"00",X"47",X"49",X"99",X"00",X"47",X"99",X"AA",X"00",X"99",X"90",X"9A",X"00",X"95",X"00",
		X"99",X"00",X"99",X"00",X"99",X"99",X"09",X"00",X"29",X"A9",X"99",X"90",X"22",X"A9",X"B9",X"99",
		X"29",X"99",X"5B",X"B9",X"99",X"99",X"5B",X"A9",X"99",X"99",X"A9",X"99",X"99",X"90",X"99",X"90",
		X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"94",X"99",X"00",
		X"00",X"44",X"49",X"00",X"00",X"44",X"CC",X"00",X"00",X"44",X"CC",X"00",X"00",X"44",X"99",X"00",
		X"00",X"4C",X"C9",X"00",X"00",X"4C",X"C9",X"00",X"00",X"49",X"C9",X"00",X"09",X"99",X"99",X"00",
		X"99",X"AA",X"9A",X"90",X"9C",X"AA",X"AA",X"99",X"CC",X"AA",X"AA",X"C9",X"CC",X"99",X"99",X"CC",
		X"CC",X"99",X"99",X"CC",X"CC",X"AA",X"AA",X"CC",X"99",X"AA",X"AA",X"C9",X"00",X"AA",X"AA",X"99",
		X"99",X"AA",X"AA",X"44",X"55",X"22",X"22",X"99",X"55",X"AA",X"AA",X"55",X"55",X"99",X"99",X"55",
		X"45",X"CC",X"CC",X"55",X"45",X"99",X"CC",X"54",X"45",X"90",X"CC",X"54",X"55",X"99",X"CC",X"54",
		X"55",X"29",X"CC",X"55",X"99",X"99",X"99",X"99",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"94",X"99",X"00",
		X"00",X"4A",X"49",X"00",X"00",X"C2",X"44",X"00",X"00",X"CC",X"44",X"00",X"00",X"9C",X"44",X"00",
		X"00",X"C4",X"44",X"00",X"00",X"C9",X"44",X"00",X"09",X"C4",X"44",X"00",X"99",X"9C",X"99",X"90",
		X"9C",X"99",X"AA",X"99",X"CC",X"AA",X"AA",X"C9",X"CC",X"AA",X"AA",X"CC",X"CC",X"AA",X"AA",X"CC",
		X"CC",X"99",X"99",X"CC",X"99",X"AA",X"99",X"C9",X"00",X"AA",X"AA",X"99",X"99",X"AA",X"AA",X"44",
		X"55",X"AA",X"AA",X"99",X"55",X"22",X"22",X"55",X"55",X"AA",X"AA",X"55",X"45",X"99",X"99",X"54",
		X"45",X"C9",X"CC",X"54",X"45",X"C9",X"9C",X"54",X"55",X"C9",X"9C",X"55",X"55",X"C9",X"99",X"55",
		X"99",X"C9",X"22",X"99",X"00",X"99",X"99",X"00",X"00",X"29",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"94",X"99",X"00",
		X"00",X"44",X"49",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"49",X"00",
		X"00",X"94",X"99",X"00",X"09",X"99",X"9A",X"00",X"99",X"99",X"AA",X"00",X"9C",X"A9",X"AA",X"90",
		X"CC",X"AA",X"AA",X"99",X"CC",X"AA",X"AA",X"C9",X"9C",X"AA",X"AA",X"CC",X"CC",X"AA",X"AA",X"99",
		X"CC",X"A9",X"9A",X"CC",X"99",X"99",X"99",X"C9",X"00",X"AA",X"AA",X"99",X"99",X"AA",X"AA",X"00",
		X"55",X"AA",X"AA",X"99",X"55",X"AA",X"AA",X"55",X"55",X"AA",X"AA",X"55",X"45",X"99",X"99",X"55",
		X"45",X"C9",X"CC",X"54",X"45",X"C9",X"9C",X"54",X"55",X"C9",X"9C",X"54",X"55",X"C9",X"99",X"55",
		X"99",X"C9",X"22",X"55",X"00",X"99",X"99",X"99",X"00",X"29",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"55",X"99",X"00",X"00",X"99",X"55",X"00",
		X"00",X"9F",X"95",X"00",X"00",X"FF",X"95",X"00",X"00",X"FF",X"99",X"00",X"00",X"FF",X"F9",X"00",
		X"00",X"FF",X"FF",X"00",X"00",X"99",X"FF",X"00",X"00",X"99",X"FF",X"00",X"00",X"F9",X"FF",X"00",
		X"00",X"FF",X"FF",X"00",X"00",X"FF",X"F9",X"00",X"00",X"FF",X"F9",X"90",X"00",X"FF",X"95",X"90",
		X"00",X"FF",X"95",X"90",X"00",X"9F",X"55",X"90",X"00",X"99",X"59",X"90",X"00",X"55",X"99",X"90",
		X"00",X"99",X"99",X"90",X"00",X"99",X"99",X"90",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"AA",X"00",X"00",X"00",X"D9",X"09",X"00",X"00",X"CC",X"09",X"00",X"00",X"9C",X"09",X"00",
		X"9D",X"99",X"99",X"00",X"9D",X"C4",X"93",X"00",X"90",X"CC",X"33",X"00",X"90",X"9C",X"33",X"00",
		X"99",X"99",X"99",X"00",X"95",X"33",X"29",X"00",X"55",X"93",X"29",X"00",X"55",X"99",X"29",X"00",
		X"55",X"99",X"99",X"00",X"55",X"99",X"96",X"00",X"55",X"99",X"66",X"00",X"99",X"33",X"66",X"90",
		X"66",X"99",X"66",X"99",X"22",X"22",X"22",X"55",X"22",X"22",X"22",X"55",X"22",X"22",X"29",X"59",
		X"29",X"92",X"99",X"99",X"99",X"99",X"97",X"96",X"97",X"79",X"77",X"96",X"97",X"79",X"75",X"96",
		X"97",X"79",X"77",X"99",X"99",X"99",X"97",X"90",X"09",X"90",X"99",X"00",X"00",X"00",X"09",X"00",
		X"00",X"99",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"99",X"00",X"00",X"99",X"94",X"00",
		X"00",X"A9",X"44",X"00",X"00",X"CC",X"99",X"00",X"00",X"9C",X"9C",X"00",X"00",X"99",X"CC",X"00",
		X"9D",X"44",X"C9",X"00",X"9D",X"99",X"9C",X"00",X"90",X"CC",X"99",X"00",X"90",X"CC",X"90",X"00",
		X"90",X"99",X"90",X"00",X"99",X"33",X"99",X"00",X"95",X"93",X"29",X"00",X"55",X"99",X"29",X"00",
		X"55",X"99",X"A9",X"00",X"55",X"99",X"99",X"00",X"55",X"99",X"96",X"00",X"55",X"33",X"66",X"00",
		X"99",X"33",X"66",X"90",X"66",X"99",X"66",X"99",X"22",X"22",X"29",X"55",X"29",X"22",X"99",X"55",
		X"99",X"92",X"97",X"59",X"97",X"92",X"77",X"99",X"97",X"96",X"77",X"96",X"97",X"96",X"77",X"96",
		X"95",X"96",X"77",X"96",X"99",X"99",X"97",X"99",X"09",X"00",X"99",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"99",X"EE",X"00",X"00",X"EE",X"AE",X"00",X"00",X"99",X"EE",X"00",X"00",X"EE",X"EE",X"00",
		X"00",X"EE",X"9E",X"00",X"00",X"EE",X"9E",X"00",X"00",X"EE",X"99",X"00",X"00",X"E9",X"E9",X"00",
		X"09",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"9E",X"90",X"99",X"00",X"99",X"00",X"99",X"00",
		X"09",X"00",X"99",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"99",X"00",X"09",X"99",X"EE",X"00",
		X"09",X"EE",X"AE",X"00",X"00",X"99",X"AE",X"00",X"00",X"9E",X"EE",X"00",X"00",X"EE",X"9E",X"00",
		X"00",X"EE",X"9E",X"00",X"00",X"EE",X"99",X"00",X"00",X"EE",X"E9",X"00",X"00",X"9E",X"99",X"00",
		X"00",X"99",X"09",X"00",X"00",X"EE",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"EA",X"00",X"00",X"00",X"EA",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"E9",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"E9",X"00",X"00",
		X"00",X"E9",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"9E",X"00",X"00",
		X"99",X"99",X"00",X"00",X"9E",X"9E",X"00",X"00",X"9E",X"EE",X"00",X"00",X"99",X"EE",X"00",X"00",
		X"09",X"99",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"00",X"00",X"99",X"94",X"00",X"00",X"09",X"09",X"00",X"00",X"00",X"00",X"90",
		X"00",X"09",X"00",X"99",X"99",X"99",X"90",X"A9",X"9A",X"9D",X"99",X"A9",X"AA",X"99",X"99",X"9A",
		X"AA",X"99",X"92",X"AA",X"99",X"99",X"99",X"99",X"AA",X"95",X"90",X"90",X"AA",X"99",X"90",X"00",
		X"99",X"99",X"90",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"94",X"90",X"00",X"00",X"44",X"99",X"00",X"FF",X"99",X"49",X"00",
		X"00",X"C9",X"C9",X"00",X"00",X"C9",X"99",X"00",X"00",X"CC",X"90",X"00",X"00",X"94",X"90",X"00",
		X"00",X"9C",X"99",X"00",X"00",X"99",X"59",X"00",X"00",X"55",X"55",X"00",X"00",X"55",X"55",X"00",
		X"00",X"99",X"99",X"00",X"00",X"59",X"99",X"00",X"00",X"55",X"99",X"00",X"00",X"55",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"22",X"90",X"00",X"00",X"22",X"90",X"00",
		X"00",X"22",X"90",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"99",X"00",
		X"00",X"09",X"9E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"9E",X"00",
		X"00",X"00",X"9E",X"00",X"00",X"00",X"99",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"94",X"90",X"00",X"00",X"44",X"90",X"00",
		X"00",X"49",X"90",X"00",X"00",X"94",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"95",X"00",X"00",X"79",X"97",X"00",X"00",X"79",X"57",X"00",
		X"00",X"99",X"79",X"00",X"00",X"77",X"79",X"00",X"00",X"77",X"99",X"00",X"00",X"97",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"22",X"90",X"00",X"00",X"22",X"90",X"00",
		X"00",X"22",X"90",X"00",X"00",X"92",X"90",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"92",X"99",X"00",X"00",X"22",X"9E",X"00",
		X"00",X"99",X"9E",X"00",X"00",X"90",X"9E",X"00",X"00",X"90",X"EE",X"00",X"00",X"90",X"99",X"00",
		X"99",X"99",X"00",X"00",X"CC",X"44",X"00",X"00",X"CC",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"9C",X"00",X"00",X"99",X"9C",X"00",X"00",X"29",X"CC",X"00",X"00",X"29",X"99",X"00",X"00",
		X"29",X"CC",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"CC",X"90",X"00",X"99",X"99",X"90",X"00",
		X"99",X"22",X"90",X"00",X"99",X"22",X"90",X"00",X"00",X"22",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"22",X"90",X"00",X"00",X"22",X"90",X"00",X"00",X"22",X"90",X"00",X"00",X"22",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"66",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",
		X"00",X"09",X"90",X"00",X"00",X"99",X"99",X"00",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"90",X"94",X"9C",X"90",X"90",X"94",X"9C",X"90",X"90",X"94",X"99",X"90",X"90",X"99",X"90",X"90",
		X"90",X"99",X"90",X"90",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"00",X"09",X"90",X"00",
		X"00",X"09",X"90",X"00",X"00",X"09",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"92",X"92",X"00",X"00",X"92",X"22",X"00",X"00",X"92",X"29",X"00",X"00",X"92",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"96",X"99",X"09",X"00",X"99",X"99",X"99",X"00",X"99",X"90",X"11",
		X"00",X"66",X"90",X"11",X"00",X"66",X"90",X"19",X"00",X"99",X"00",X"19",X"00",X"99",X"00",X"90",
		X"00",X"19",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"90",X"00",X"09",X"49",X"90",X"00",X"09",X"44",X"90",X"00",X"99",X"44",X"99",
		X"00",X"94",X"44",X"99",X"00",X"94",X"94",X"99",X"00",X"94",X"44",X"99",X"00",X"99",X"99",X"90",
		X"00",X"09",X"9C",X"90",X"00",X"09",X"CC",X"99",X"00",X"99",X"99",X"99",X"00",X"29",X"92",X"99",
		X"00",X"29",X"29",X"99",X"00",X"99",X"22",X"99",X"00",X"92",X"22",X"00",X"00",X"22",X"22",X"00",
		X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"92",X"22",X"00",X"00",X"99",X"29",X"00",
		X"00",X"99",X"99",X"00",X"00",X"96",X"66",X"00",X"00",X"96",X"99",X"00",X"00",X"99",X"66",X"00",
		X"00",X"09",X"69",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"99",X"00",
		X"00",X"99",X"91",X"00",X"00",X"91",X"91",X"00",X"00",X"11",X"99",X"00",X"00",X"99",X"09",X"00",
		X"00",X"99",X"00",X"00",X"00",X"44",X"00",X"00",X"99",X"99",X"99",X"99",X"99",X"C9",X"99",X"99",
		X"00",X"C9",X"90",X"00",X"00",X"C9",X"90",X"00",X"00",X"9C",X"90",X"00",X"00",X"CC",X"90",X"00",
		X"00",X"49",X"90",X"00",X"99",X"9C",X"99",X"99",X"99",X"99",X"99",X"99",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",
		X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"00",X"79",X"00",X"94",X"00",X"79",X"00",X"44",X"90",X"AA",X"00",X"44",X"99",X"AA",X"00",
		X"99",X"99",X"97",X"00",X"EE",X"C9",X"97",X"00",X"EE",X"CC",X"97",X"90",X"C4",X"99",X"99",X"99",
		X"C4",X"00",X"00",X"39",X"CC",X"00",X"99",X"99",X"99",X"00",X"33",X"90",X"55",X"00",X"11",X"00",
		X"55",X"00",X"33",X"00",X"55",X"00",X"99",X"00",X"95",X"90",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"EE",X"00",X"00",X"55",X"CC",X"09",X"99",X"55",X"9C",X"99",X"99",X"55",X"9C",X"77",X"44",
		X"99",X"99",X"77",X"44",X"11",X"00",X"74",X"44",X"11",X"00",X"94",X"44",X"91",X"90",X"99",X"49",
		X"99",X"99",X"09",X"99",X"99",X"11",X"00",X"90",X"19",X"11",X"00",X"00",X"99",X"19",X"00",X"90",
		X"90",X"99",X"00",X"90",X"99",X"99",X"00",X"90",X"99",X"00",X"00",X"90",X"99",X"00",X"00",X"00",
		X"09",X"00",X"00",X"69",X"99",X"00",X"09",X"97",X"94",X"99",X"09",X"77",X"44",X"49",X"09",X"77",
		X"99",X"99",X"09",X"77",X"EE",X"CC",X"09",X"99",X"EE",X"CC",X"09",X"69",X"EC",X"99",X"00",X"69",
		X"CC",X"90",X"00",X"99",X"9C",X"90",X"99",X"09",X"99",X"90",X"33",X"99",X"55",X"00",X"11",X"93",
		X"55",X"00",X"31",X"31",X"95",X"90",X"99",X"99",X"99",X"99",X"00",X"00",X"99",X"EE",X"00",X"90",
		X"55",X"CC",X"99",X"99",X"55",X"9C",X"99",X"99",X"55",X"9C",X"77",X"44",X"99",X"99",X"77",X"44",
		X"11",X"00",X"44",X"44",X"11",X"00",X"94",X"44",X"11",X"00",X"99",X"49",X"99",X"00",X"09",X"99",
		X"19",X"00",X"00",X"90",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"19",X"00",X"00",X"00",
		X"19",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"9C",X"99",X"00",X"00",X"99",X"99",X"00",X"99",X"99",X"CC",X"00",X"9C",X"99",X"9C",X"00",
		X"CC",X"99",X"94",X"00",X"9C",X"99",X"44",X"00",X"99",X"9C",X"9C",X"00",X"00",X"99",X"9C",X"00",
		X"00",X"49",X"C9",X"00",X"00",X"44",X"99",X"00",X"00",X"99",X"94",X"00",X"00",X"99",X"44",X"00",
		X"00",X"99",X"49",X"00",X"00",X"94",X"99",X"00",X"00",X"94",X"44",X"00",X"00",X"94",X"44",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"92",X"00",X"00",X"92",X"22",X"00",X"00",X"92",X"22",X"00",
		X"00",X"22",X"22",X"00",X"00",X"22",X"92",X"00",X"00",X"22",X"29",X"00",X"00",X"92",X"22",X"00",
		X"00",X"99",X"99",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"99",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"94",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"A9",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"C9",X"00",X"00",X"00",X"CC",X"90",X"00",X"00",X"49",X"99",X"00",
		X"00",X"9C",X"79",X"00",X"00",X"99",X"79",X"00",X"00",X"97",X"99",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"99",X"00",X"99",X"CC",X"99",X"00",X"49",X"CC",X"79",X"00",X"00",X"99",X"99",X"00",
		X"00",X"09",X"D9",X"00",X"00",X"09",X"D9",X"00",X"00",X"09",X"D9",X"00",X"00",X"09",X"99",X"00",
		X"00",X"00",X"9D",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"DD",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"09",X"00",X"99",X"00",X"92",X"99",X"90",
		X"90",X"92",X"11",X"99",X"99",X"92",X"94",X"19",X"41",X"72",X"95",X"19",X"41",X"72",X"96",X"99",
		X"99",X"92",X"11",X"19",X"00",X"92",X"11",X"99",X"00",X"92",X"91",X"19",X"00",X"92",X"91",X"99",
		X"00",X"09",X"99",X"19",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"99",X"00",X"00",
		X"09",X"9A",X"00",X"00",X"09",X"9A",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"CC",X"00",X"00",
		X"09",X"C9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"09",X"99",X"90",X"00",X"99",X"CC",X"99",X"00",X"94",X"99",X"49",X"00",X"44",X"44",X"44",X"00",
		X"44",X"94",X"94",X"00",X"99",X"99",X"94",X"00",X"99",X"44",X"44",X"00",X"90",X"94",X"44",X"00",
		X"90",X"94",X"99",X"00",X"90",X"99",X"44",X"00",X"90",X"22",X"99",X"00",X"90",X"92",X"C9",X"00",
		X"99",X"99",X"C9",X"00",X"09",X"92",X"90",X"00",X"09",X"99",X"00",X"00",X"09",X"09",X"00",X"00",
		X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"A9",X"90",X"00",X"00",X"A9",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"CC",X"90",X"00",
		X"00",X"9C",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"44",X"CC",X"90",X"00",X"44",X"99",X"99",X"00",X"49",X"44",X"49",X"00",
		X"49",X"94",X"44",X"00",X"49",X"99",X"94",X"00",X"99",X"44",X"94",X"00",X"C9",X"94",X"44",X"00",
		X"C9",X"94",X"44",X"00",X"99",X"99",X"99",X"00",X"00",X"22",X"44",X"00",X"00",X"92",X"99",X"00",
		X"00",X"99",X"C9",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"90",X"00",X"00",X"09",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"9C",X"90",X"00",X"00",X"CC",X"99",X"00",X"00",X"9C",X"99",X"00",
		X"00",X"9C",X"99",X"00",X"00",X"9C",X"99",X"00",X"00",X"CC",X"C9",X"00",X"00",X"CC",X"C9",X"00",
		X"00",X"CC",X"C9",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"99",X"00",X"00",X"CC",X"49",X"00",X"99",X"99",X"49",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"94",X"99",X"00",X"99",X"94",X"99",X"00",
		X"99",X"94",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"91",X"00",X"29",X"00",
		X"91",X"00",X"91",X"00",X"99",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"99",X"00",
		X"00",X"99",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"C9",X"90",X"00",X"00",X"C9",X"90",X"00",
		X"00",X"C9",X"90",X"00",X"00",X"C9",X"90",X"00",X"00",X"CC",X"90",X"00",X"00",X"CC",X"90",X"00",
		X"00",X"CC",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"99",X"00",X"00",X"CC",X"44",X"00",X"00",X"99",X"44",X"00",X"99",X"99",X"49",X"00",
		X"99",X"9D",X"99",X"00",X"99",X"9D",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"C9",X"99",X"00",X"99",X"CC",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"9D",X"99",X"00",
		X"99",X"9D",X"99",X"00",X"99",X"9D",X"99",X"00",X"99",X"9D",X"99",X"00",X"99",X"99",X"99",X"00",
		X"00",X"99",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"9C",X"90",X"00",X"00",X"CC",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"C9",X"00",X"00",X"99",X"C9",X"00",X"00",X"99",X"C9",X"00",
		X"00",X"CC",X"99",X"00",X"00",X"CC",X"90",X"00",X"00",X"CC",X"90",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"99",X"99",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"09",X"44",X"99",X"00",
		X"09",X"44",X"99",X"00",X"09",X"44",X"49",X"00",X"09",X"44",X"49",X"00",X"09",X"44",X"49",X"00",
		X"09",X"49",X"49",X"00",X"09",X"99",X"99",X"00",X"09",X"22",X"99",X"00",X"09",X"99",X"29",X"00",
		X"00",X"19",X"29",X"00",X"00",X"11",X"29",X"00",X"00",X"99",X"99",X"00",X"00",X"11",X"99",X"00",
		X"00",X"11",X"19",X"00",X"00",X"11",X"19",X"00",X"00",X"19",X"99",X"00",X"00",X"99",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"9C",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"9C",X"00",X"00",X"99",X"CC",X"00",X"00",X"99",X"CC",X"00",
		X"00",X"CC",X"C9",X"00",X"00",X"CC",X"C9",X"00",X"00",X"CC",X"99",X"00",X"00",X"9C",X"90",X"00",
		X"00",X"99",X"99",X"00",X"00",X"44",X"44",X"00",X"09",X"44",X"44",X"00",X"09",X"44",X"44",X"00",
		X"09",X"44",X"99",X"00",X"09",X"44",X"99",X"00",X"09",X"44",X"49",X"00",X"09",X"49",X"49",X"00",
		X"09",X"99",X"99",X"00",X"09",X"22",X"29",X"00",X"09",X"92",X"29",X"00",X"00",X"99",X"99",X"00",
		X"00",X"22",X"19",X"00",X"00",X"99",X"11",X"00",X"00",X"22",X"99",X"00",X"00",X"99",X"11",X"00",
		X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"99",X"19",X"00",X"00",X"00",X"99",X"00",
		X"00",X"09",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"9A",X"00",X"00",X"99",X"9A",X"00",
		X"00",X"99",X"9A",X"00",X"00",X"99",X"9A",X"00",X"00",X"C9",X"99",X"00",X"00",X"C9",X"CC",X"00",
		X"00",X"CC",X"C9",X"00",X"00",X"9C",X"99",X"00",X"00",X"9C",X"99",X"00",X"00",X"9C",X"99",X"00",
		X"00",X"99",X"49",X"00",X"00",X"49",X"C9",X"00",X"00",X"99",X"99",X"00",X"90",X"44",X"44",X"00",
		X"90",X"44",X"44",X"00",X"90",X"99",X"99",X"00",X"99",X"99",X"49",X"00",X"29",X"44",X"99",X"00",
		X"29",X"44",X"92",X"90",X"99",X"99",X"29",X"99",X"29",X"99",X"99",X"19",X"22",X"00",X"99",X"19",
		X"92",X"00",X"99",X"99",X"99",X"00",X"09",X"90",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"CC",X"00",
		X"00",X"99",X"9A",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"9A",X"00",X"00",X"C9",X"CC",X"00",
		X"00",X"C9",X"CC",X"00",X"00",X"CC",X"C9",X"00",X"00",X"9C",X"99",X"00",X"00",X"9C",X"99",X"90",
		X"00",X"9C",X"99",X"90",X"00",X"99",X"44",X"90",X"00",X"99",X"CC",X"90",X"00",X"49",X"99",X"90",
		X"00",X"44",X"44",X"00",X"09",X"44",X"44",X"00",X"09",X"99",X"99",X"00",X"09",X"99",X"00",X"00",
		X"09",X"44",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",
		X"99",X"92",X"00",X"00",X"92",X"29",X"00",X"00",X"22",X"99",X"00",X"00",X"92",X"90",X"00",X"00",
		X"99",X"00",X"00",X"00",X"19",X"99",X"00",X"00",X"11",X"19",X"00",X"00",X"99",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"99",X"CC",X"90",X"00",X"09",X"CC",X"00",X"00",X"09",X"CC",X"00",X"00",
		X"09",X"C9",X"00",X"00",X"09",X"C9",X"00",X"00",X"09",X"C9",X"00",X"00",X"09",X"CC",X"00",X"00",
		X"99",X"C9",X"90",X"00",X"09",X"99",X"00",X"00",X"00",X"49",X"90",X"00",X"09",X"9F",X"90",X"00",
		X"09",X"99",X"90",X"00",X"99",X"CC",X"99",X"00",X"99",X"99",X"99",X"00",X"49",X"44",X"99",X"00",
		X"49",X"49",X"99",X"00",X"49",X"99",X"99",X"00",X"44",X"49",X"99",X"00",X"99",X"44",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"22",X"00",X"00",X"09",X"99",X"00",X"00",
		X"09",X"09",X"00",X"00",X"09",X"09",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"9C",X"99",X"00",X"00",X"C9",X"99",X"00",
		X"00",X"C9",X"99",X"00",X"00",X"C9",X"9C",X"00",X"00",X"C9",X"CC",X"00",X"00",X"C9",X"44",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"9C",X"CC",X"00",X"00",X"99",X"CC",X"00",X"00",X"99",X"9C",X"00",X"00",X"94",X"CC",X"00",
		X"00",X"94",X"CC",X"00",X"00",X"44",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"94",X"99",X"00",
		X"00",X"44",X"99",X"00",X"00",X"99",X"29",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"19",X"00",
		X"00",X"22",X"11",X"00",X"00",X"29",X"11",X"00",X"00",X"99",X"11",X"00",X"00",X"19",X"99",X"00",
		X"00",X"99",X"11",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"9C",X"99",X"00",X"00",X"CC",X"99",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"C9",X"00",X"00",X"99",X"C9",X"00",X"00",X"99",X"C9",X"00",
		X"09",X"CC",X"99",X"00",X"09",X"CC",X"99",X"00",X"09",X"99",X"9C",X"00",X"09",X"44",X"CC",X"00",
		X"09",X"44",X"9C",X"00",X"09",X"44",X"99",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"49",X"00",
		X"00",X"44",X"49",X"00",X"00",X"99",X"49",X"00",X"00",X"44",X"49",X"00",X"00",X"99",X"49",X"00",
		X"00",X"22",X"99",X"00",X"00",X"22",X"29",X"00",X"00",X"99",X"29",X"00",X"00",X"19",X"29",X"00",
		X"00",X"11",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"11",X"99",X"00",X"00",X"11",X"19",X"00",
		X"00",X"11",X"99",X"00",X"00",X"19",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"09",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"CC",X"99",X"00",X"09",X"CC",X"CC",X"00",X"09",X"99",X"CC",X"00",X"09",X"44",X"9C",X"00",
		X"09",X"44",X"99",X"00",X"09",X"44",X"49",X"00",X"09",X"44",X"49",X"00",X"09",X"49",X"99",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"22",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"99",X"9A",X"99",X"00",
		X"DD",X"92",X"99",X"00",X"99",X"99",X"CC",X"00",X"99",X"CC",X"9C",X"00",X"99",X"CC",X"CC",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"C9",X"00",X"99",X"99",X"99",X"00",X"99",X"CC",X"90",X"00",
		X"99",X"9C",X"99",X"00",X"99",X"99",X"49",X"00",X"99",X"49",X"49",X"00",X"99",X"99",X"44",X"00",
		X"99",X"94",X"49",X"00",X"DD",X"94",X"49",X"00",X"99",X"99",X"99",X"00",X"99",X"44",X"99",X"00",
		X"99",X"44",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"22",X"29",X"00",X"99",X"22",X"29",X"00",
		X"99",X"22",X"29",X"00",X"99",X"22",X"29",X"00",X"99",X"92",X"99",X"00",X"99",X"22",X"29",X"00",
		X"99",X"99",X"99",X"00",X"99",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"99",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"9C",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"DD",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"9C",X"00",X"00",X"9F",X"9C",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"94",X"00",X"00",X"99",X"94",X"00",X"00",X"9F",X"9C",X"00",X"00",X"99",X"9C",X"00",
		X"00",X"99",X"CC",X"00",X"00",X"DD",X"CC",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"9F",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"91",X"00",X"00",X"11",X"11",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"9C",X"99",X"00",X"00",X"CC",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"C9",X"00",X"00",X"99",X"C9",X"00",X"00",X"99",X"C9",X"00",
		X"00",X"CC",X"99",X"00",X"00",X"CC",X"99",X"00",X"00",X"CC",X"99",X"00",X"00",X"CC",X"99",X"00",
		X"00",X"99",X"49",X"00",X"00",X"99",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"49",X"00",
		X"00",X"44",X"99",X"00",X"00",X"94",X"99",X"00",X"00",X"44",X"49",X"00",X"00",X"44",X"49",X"00",
		X"00",X"99",X"49",X"00",X"00",X"92",X"99",X"00",X"00",X"22",X"29",X"00",X"00",X"22",X"29",X"00",
		X"00",X"22",X"29",X"00",X"00",X"22",X"29",X"00",X"00",X"22",X"29",X"00",X"00",X"22",X"29",X"00",
		X"00",X"22",X"29",X"00",X"00",X"99",X"99",X"00",X"00",X"11",X"11",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"90",X"00",X"00",X"9C",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"CC",X"90",X"00",
		X"00",X"CC",X"90",X"00",X"00",X"CC",X"90",X"00",X"00",X"C9",X"90",X"00",X"00",X"99",X"90",X"00",
		X"09",X"99",X"90",X"00",X"09",X"CC",X"00",X"00",X"99",X"99",X"00",X"00",X"94",X"99",X"00",X"00",
		X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"49",X"49",X"90",X"00",X"99",X"44",X"90",X"00",
		X"90",X"44",X"90",X"00",X"90",X"44",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"22",X"99",X"00",
		X"00",X"22",X"19",X"00",X"00",X"22",X"19",X"00",X"00",X"22",X"19",X"00",X"00",X"92",X"19",X"00",
		X"00",X"99",X"19",X"00",X"00",X"09",X"19",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"99",X"00",
		X"00",X"99",X"00",X"00",X"00",X"9C",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9C",X"00",X"00",
		X"00",X"9C",X"00",X"00",X"00",X"9C",X"90",X"00",X"00",X"9C",X"90",X"00",X"00",X"CC",X"90",X"00",
		X"00",X"CC",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"94",X"00",X"00",
		X"09",X"99",X"00",X"00",X"09",X"CC",X"99",X"99",X"09",X"99",X"49",X"C9",X"09",X"99",X"49",X"99",
		X"09",X"44",X"99",X"00",X"09",X"44",X"00",X"00",X"09",X"49",X"90",X"00",X"09",X"94",X"90",X"00",
		X"09",X"99",X"90",X"00",X"09",X"11",X"90",X"00",X"99",X"11",X"99",X"00",X"99",X"11",X"22",X"00",
		X"C9",X"11",X"22",X"00",X"CC",X"11",X"99",X"00",X"C9",X"99",X"00",X"00",X"99",X"11",X"00",X"00",
		X"00",X"19",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"0A",X"00",X"00",X"CC",X"0A",X"00",X"09",X"9C",X"00",X"00",X"09",X"CC",X"99",X"00",
		X"09",X"CC",X"C9",X"00",X"09",X"C9",X"C9",X"00",X"09",X"C9",X"99",X"00",X"09",X"CC",X"49",X"00",
		X"09",X"99",X"99",X"00",X"09",X"99",X"49",X"00",X"00",X"94",X"49",X"00",X"00",X"44",X"49",X"00",
		X"09",X"49",X"49",X"00",X"09",X"99",X"99",X"00",X"09",X"CC",X"90",X"00",X"09",X"99",X"00",X"00",
		X"09",X"44",X"00",X"00",X"09",X"44",X"00",X"00",X"09",X"49",X"90",X"00",X"09",X"94",X"90",X"00",
		X"09",X"99",X"90",X"00",X"09",X"11",X"90",X"00",X"99",X"11",X"99",X"00",X"99",X"11",X"22",X"00",
		X"C9",X"11",X"22",X"00",X"CC",X"11",X"99",X"00",X"C9",X"99",X"00",X"00",X"99",X"11",X"00",X"00",
		X"00",X"19",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"9D",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",X"00",
		X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",X"00",
		X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",X"00",
		X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",X"00",
		X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",X"00",
		X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",X"00",
		X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",
		X"9D",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"9D",X"00",X"00",X"99",X"9D",X"00",X"00",X"99",X"D9",X"00",X"00",
		X"09",X"9D",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"D9",X"00",
		X"00",X"09",X"9D",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"09",X"9F",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"9F",X"99",X"9F",X"00",X"DD",X"DD",X"DD",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"D9",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9F",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"90",X"00",X"00",
		X"99",X"99",X"00",X"00",X"DD",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"9F",X"99",X"00",X"00",
		X"09",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"9D",X"90",X"00",
		X"00",X"99",X"99",X"00",X"00",X"DD",X"99",X"00",X"00",X"D9",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"09",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"9D",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"F9",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"F9",X"D9",X"00",
		X"00",X"99",X"9D",X"00",X"00",X"99",X"DD",X"00",X"00",X"D9",X"D9",X"00",X"00",X"DD",X"99",X"00",
		X"00",X"9D",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"DD",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"DD",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"DD",X"DD",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"F9",X"9F",X"00",X"00",X"99",X"99",X"00",X"00",X"DD",X"DD",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"F9",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"F9",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"DD",X"D9",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"F9",X"00",X"00",
		X"99",X"99",X"00",X"00",X"DD",X"DD",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"F9",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"F9",X"00",X"00",
		X"99",X"99",X"00",X"00",X"DD",X"DD",X"00",X"00",X"99",X"99",X"00",X"00",X"F9",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"DD",X"DD",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"CC",X"99",X"00",X"00",X"99",X"C9",X"00",X"99",X"4E",X"C9",X"00",
		X"9C",X"4C",X"CC",X"00",X"9C",X"CC",X"C9",X"00",X"9C",X"9C",X"CC",X"00",X"99",X"99",X"C9",X"00",
		X"99",X"CC",X"C9",X"00",X"99",X"99",X"C9",X"00",X"99",X"F9",X"C9",X"90",X"99",X"99",X"C9",X"90",
		X"99",X"9F",X"99",X"90",X"99",X"99",X"99",X"90",X"99",X"44",X"99",X"90",X"99",X"CC",X"99",X"90",
		X"99",X"99",X"99",X"90",X"99",X"99",X"D9",X"90",X"99",X"99",X"D9",X"90",X"99",X"99",X"99",X"90",
		X"CC",X"49",X"9C",X"90",X"CC",X"49",X"9C",X"90",X"CC",X"44",X"9C",X"90",X"CC",X"44",X"99",X"90",
		X"CC",X"94",X"99",X"90",X"C9",X"99",X"9C",X"90",X"99",X"99",X"CC",X"00",X"C9",X"CC",X"CC",X"00",
		X"C9",X"CC",X"CC",X"00",X"C9",X"CC",X"EC",X"00",X"C9",X"CC",X"CE",X"00",X"CC",X"CC",X"CC",X"00",
		X"CC",X"CC",X"99",X"00",X"CC",X"99",X"BB",X"00",X"C9",X"BB",X"BB",X"00",X"C9",X"BB",X"BB",X"00",
		X"C9",X"BB",X"BB",X"00",X"C9",X"B9",X"BB",X"00",X"C9",X"99",X"BB",X"00",X"9B",X"B9",X"BB",X"00",
		X"BB",X"99",X"BB",X"00",X"BB",X"90",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",
		X"B9",X"00",X"BB",X"00",X"99",X"00",X"BB",X"00",X"EE",X"00",X"BB",X"00",X"77",X"00",X"BB",X"00",
		X"77",X"00",X"BB",X"00",X"77",X"00",X"BB",X"00",X"99",X"00",X"BB",X"00",X"77",X"09",X"BB",X"00",
		X"97",X"09",X"99",X"00",X"99",X"09",X"BB",X"00",X"00",X"09",X"BB",X"00",X"00",X"09",X"99",X"00",
		X"00",X"09",X"77",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"59",X"09",X"00",X"00",X"79",X"99",X"00",X"00",X"79",X"95",X"00",X"00",X"79",X"55",X"00",X"00",
		X"99",X"55",X"00",X"00",X"55",X"59",X"00",X"00",X"55",X"99",X"99",X"00",X"55",X"99",X"55",X"00",
		X"55",X"95",X"55",X"00",X"55",X"55",X"95",X"90",X"59",X"55",X"95",X"90",X"59",X"55",X"95",X"90",
		X"99",X"55",X"55",X"90",X"00",X"59",X"55",X"90",X"00",X"59",X"55",X"90",X"00",X"55",X"55",X"90",
		X"00",X"55",X"95",X"90",X"00",X"55",X"95",X"00",X"00",X"55",X"99",X"00",X"00",X"95",X"55",X"00",
		X"00",X"95",X"55",X"00",X"00",X"99",X"59",X"00",X"00",X"79",X"99",X"00",X"00",X"97",X"99",X"00",
		X"00",X"99",X"59",X"00",X"00",X"59",X"55",X"00",X"00",X"55",X"99",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"90",X"00",X"00",X"79",X"90",X"00",X"00",X"79",X"99",X"00",X"90",X"99",X"59",X"00",X"90",
		X"55",X"59",X"00",X"90",X"55",X"59",X"00",X"90",X"55",X"59",X"99",X"90",X"55",X"59",X"55",X"90",
		X"55",X"55",X"55",X"90",X"59",X"55",X"55",X"90",X"59",X"95",X"95",X"00",X"99",X"95",X"95",X"00",
		X"09",X"99",X"95",X"00",X"09",X"55",X"55",X"00",X"99",X"59",X"55",X"00",X"77",X"59",X"55",X"90",
		X"79",X"55",X"95",X"99",X"99",X"55",X"95",X"79",X"95",X"99",X"99",X"99",X"59",X"00",X"09",X"99",
		X"59",X"00",X"09",X"99",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"9C",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"C9",X"00",X"00",X"CC",X"C9",X"00",
		X"00",X"44",X"99",X"00",X"00",X"49",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"C9",X"00",X"00",
		X"09",X"CC",X"00",X"00",X"09",X"CC",X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"99",X"99",X"00",
		X"99",X"94",X"99",X"00",X"99",X"99",X"9F",X"00",X"99",X"49",X"99",X"00",X"99",X"94",X"99",X"00",
		X"99",X"44",X"99",X"00",X"99",X"9C",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"22",X"99",X"00",
		X"99",X"22",X"99",X"00",X"99",X"22",X"99",X"00",X"99",X"22",X"99",X"00",X"99",X"22",X"99",X"00",
		X"00",X"99",X"90",X"00",X"00",X"11",X"90",X"00",X"00",X"11",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"9C",X"90",X"00",X"00",X"CC",X"90",X"00",
		X"00",X"44",X"90",X"00",X"00",X"49",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"99",X"C9",X"00",X"00",X"94",X"CC",X"00",X"00",X"94",X"99",X"99",X"00",X"44",X"99",X"99",X"00",
		X"44",X"44",X"F9",X"00",X"49",X"44",X"99",X"00",X"99",X"44",X"99",X"00",X"99",X"44",X"99",X"00",
		X"99",X"44",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"22",X"99",X"00",X"99",X"92",X"99",X"00",
		X"99",X"99",X"29",X"00",X"99",X"99",X"29",X"00",X"99",X"99",X"29",X"00",X"11",X"90",X"99",X"00",
		X"11",X"00",X"91",X"00",X"91",X"00",X"99",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"90",X"99",X"00",X"00",X"99",X"99",X"90",X"00",X"44",X"9C",X"90",X"00",X"94",X"CC",X"90",X"00",
		X"99",X"44",X"90",X"00",X"49",X"49",X"00",X"00",X"44",X"99",X"00",X"00",X"49",X"99",X"00",X"00",
		X"44",X"C9",X"00",X"00",X"94",X"CC",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"99",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"22",X"90",X"00",X"00",X"92",X"99",X"00",
		X"00",X"99",X"29",X"00",X"00",X"90",X"29",X"00",X"99",X"90",X"29",X"00",X"11",X"90",X"99",X"00",
		X"11",X"00",X"91",X"00",X"91",X"00",X"99",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"CC",X"99",X"30",X"00",X"F9",X"99",X"00",X"99",X"F9",X"99",X"00",
		X"9C",X"F9",X"9C",X"00",X"9C",X"F9",X"99",X"00",X"9C",X"9C",X"CC",X"00",X"99",X"9C",X"C9",X"00",
		X"99",X"C9",X"C9",X"00",X"99",X"CC",X"99",X"00",X"99",X"CC",X"C9",X"00",X"99",X"99",X"C9",X"00",
		X"99",X"94",X"99",X"90",X"99",X"99",X"99",X"90",X"99",X"C9",X"99",X"90",X"99",X"CC",X"9D",X"90",
		X"99",X"99",X"9D",X"90",X"99",X"99",X"9D",X"90",X"C9",X"99",X"9D",X"90",X"CC",X"99",X"99",X"90",
		X"CC",X"49",X"99",X"90",X"CC",X"49",X"99",X"90",X"CC",X"44",X"99",X"90",X"99",X"99",X"99",X"90",
		X"00",X"99",X"90",X"99",X"09",X"90",X"99",X"09",X"99",X"90",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"A4",X"99",X"00",X"00",X"AA",X"49",X"00",X"99",X"9A",X"99",X"00",
		X"94",X"AA",X"94",X"00",X"94",X"44",X"49",X"00",X"94",X"94",X"44",X"00",X"99",X"99",X"49",X"00",
		X"99",X"44",X"49",X"00",X"99",X"99",X"49",X"00",X"99",X"9F",X"49",X"90",X"99",X"99",X"49",X"90",
		X"99",X"9F",X"99",X"90",X"99",X"9F",X"99",X"90",X"99",X"99",X"99",X"90",X"99",X"44",X"99",X"90",
		X"99",X"99",X"99",X"90",X"99",X"99",X"D9",X"90",X"99",X"99",X"D9",X"90",X"99",X"99",X"99",X"90",
		X"CC",X"49",X"9C",X"90",X"CC",X"49",X"9C",X"90",X"CC",X"44",X"9C",X"90",X"CC",X"44",X"99",X"90",
		X"CC",X"94",X"99",X"90",X"C9",X"99",X"9C",X"90",X"99",X"99",X"CC",X"00",X"C9",X"CC",X"CC",X"00",
		X"C9",X"CC",X"CC",X"00",X"C9",X"CC",X"EC",X"00",X"C9",X"CC",X"CE",X"00",X"CC",X"CC",X"CC",X"00",
		X"CC",X"CC",X"99",X"00",X"CC",X"99",X"FF",X"00",X"C9",X"44",X"F4",X"00",X"C9",X"FF",X"F4",X"00",
		X"C9",X"FF",X"FF",X"00",X"C9",X"9F",X"FF",X"00",X"C9",X"99",X"F4",X"00",X"99",X"99",X"F4",X"00",
		X"99",X"90",X"99",X"00",X"EE",X"90",X"EE",X"00",X"CC",X"99",X"EC",X"00",X"CC",X"C9",X"CE",X"00",
		X"9C",X"C9",X"C9",X"00",X"99",X"E9",X"E9",X"00",X"09",X"C9",X"CC",X"00",X"99",X"90",X"CE",X"00",
		X"9C",X"90",X"EC",X"00",X"99",X"00",X"CE",X"00",X"B9",X"00",X"EC",X"00",X"3B",X"00",X"9C",X"90",
		X"BB",X"90",X"99",X"90",X"BB",X"99",X"99",X"B0",X"99",X"BB",X"31",X"90",X"9B",X"BB",X"BB",X"90",
		X"99",X"B9",X"B9",X"90",X"99",X"99",X"99",X"00",X"BB",X"9B",X"9B",X"00",X"99",X"B9",X"BB",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",
		X"09",X"00",X"91",X"00",X"99",X"00",X"99",X"90",X"2C",X"00",X"E9",X"90",X"2A",X"00",X"EE",X"90",
		X"2C",X"99",X"EE",X"99",X"CC",X"55",X"99",X"99",X"CC",X"99",X"45",X"49",X"CC",X"00",X"45",X"49",
		X"99",X"00",X"45",X"49",X"99",X"00",X"45",X"49",X"99",X"00",X"45",X"49",X"69",X"00",X"45",X"49",
		X"66",X"00",X"45",X"49",X"99",X"00",X"45",X"49",X"99",X"00",X"45",X"49",X"66",X"00",X"45",X"09",
		X"99",X"00",X"47",X"99",X"AA",X"00",X"47",X"90",X"AA",X"00",X"47",X"00",X"AA",X"00",X"99",X"00",
		X"AA",X"00",X"59",X"00",X"AA",X"00",X"59",X"00",X"AA",X"00",X"99",X"00",X"AA",X"00",X"99",X"90",
		X"AA",X"00",X"95",X"99",X"99",X"00",X"95",X"B9",X"99",X"00",X"99",X"99",X"99",X"00",X"00",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",
		X"09",X"00",X"91",X"00",X"99",X"00",X"99",X"90",X"2C",X"00",X"E9",X"90",X"2A",X"00",X"EE",X"90",
		X"2C",X"99",X"99",X"99",X"CC",X"55",X"45",X"49",X"CC",X"99",X"45",X"49",X"CC",X"00",X"45",X"49",
		X"99",X"00",X"45",X"49",X"99",X"00",X"45",X"49",X"99",X"00",X"45",X"49",X"69",X"00",X"45",X"49",
		X"66",X"00",X"45",X"49",X"99",X"00",X"45",X"49",X"99",X"00",X"45",X"49",X"66",X"00",X"47",X"99",
		X"66",X"00",X"47",X"90",X"99",X"00",X"47",X"00",X"AA",X"00",X"99",X"00",X"AA",X"00",X"59",X"00",
		X"AA",X"99",X"59",X"00",X"9A",X"99",X"99",X"00",X"99",X"99",X"09",X"00",X"99",X"99",X"99",X"00",
		X"90",X"99",X"95",X"00",X"00",X"90",X"95",X"00",X"90",X"00",X"99",X"00",X"90",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"94",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"90",X"00",X"00",X"44",X"90",X"00",X"00",X"4C",X"90",X"00",X"00",X"CC",X"90",X"00",
		X"00",X"CC",X"09",X"00",X"09",X"CC",X"9A",X"00",X"99",X"CC",X"AA",X"00",X"9A",X"9C",X"AA",X"00",
		X"C9",X"99",X"AA",X"00",X"CC",X"AA",X"99",X"00",X"CC",X"A9",X"99",X"90",X"CC",X"99",X"99",X"90",
		X"C9",X"92",X"92",X"90",X"C9",X"AA",X"A2",X"90",X"99",X"AA",X"AA",X"99",X"00",X"AA",X"A9",X"09",
		X"99",X"AA",X"99",X"49",X"55",X"22",X"29",X"99",X"55",X"AA",X"AA",X"59",X"55",X"99",X"99",X"59",
		X"45",X"C9",X"90",X"59",X"45",X"90",X"90",X"59",X"45",X"00",X"90",X"59",X"59",X"00",X"90",X"59",
		X"59",X"00",X"90",X"59",X"99",X"00",X"90",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"29",X"00",
		X"00",X"99",X"00",X"00",X"00",X"94",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"A2",X"90",X"00",X"00",X"22",X"90",X"00",X"00",X"CC",X"90",X"00",X"00",X"CC",X"99",X"00",
		X"09",X"4C",X"9A",X"00",X"99",X"99",X"9A",X"00",X"9A",X"4C",X"9A",X"00",X"C9",X"CC",X"9A",X"00",
		X"CC",X"99",X"99",X"00",X"CC",X"AA",X"A9",X"90",X"CC",X"A9",X"99",X"90",X"C9",X"99",X"99",X"90",
		X"C9",X"92",X"92",X"90",X"99",X"AA",X"22",X"90",X"00",X"AA",X"A2",X"99",X"99",X"AA",X"AA",X"49",
		X"55",X"AA",X"AA",X"99",X"55",X"22",X"29",X"59",X"55",X"AA",X"AA",X"59",X"45",X"99",X"99",X"59",
		X"45",X"00",X"C9",X"59",X"45",X"00",X"C9",X"59",X"55",X"00",X"C9",X"59",X"55",X"00",X"99",X"59",
		X"99",X"00",X"22",X"99",X"00",X"00",X"99",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"94",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"90",X"00",X"00",X"44",X"90",X"00",X"00",X"44",X"90",X"00",X"09",X"44",X"99",X"00",
		X"99",X"44",X"AA",X"00",X"9A",X"44",X"AA",X"00",X"9A",X"94",X"AA",X"00",X"C9",X"99",X"AA",X"00",
		X"CC",X"99",X"99",X"00",X"CC",X"A9",X"A9",X"90",X"99",X"AA",X"A9",X"90",X"90",X"AA",X"AA",X"90",
		X"90",X"99",X"AA",X"90",X"90",X"AA",X"9A",X"90",X"00",X"AA",X"AA",X"99",X"99",X"AA",X"AA",X"09",
		X"55",X"AA",X"AA",X"99",X"55",X"AA",X"A9",X"59",X"55",X"AA",X"AA",X"59",X"45",X"99",X"99",X"59",
		X"45",X"00",X"C9",X"59",X"45",X"00",X"C9",X"59",X"55",X"00",X"C9",X"59",X"55",X"00",X"99",X"59",
		X"99",X"00",X"22",X"59",X"00",X"00",X"99",X"99",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"95",X"00",X"00",
		X"00",X"95",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"55",X"90",X"00",X"09",X"99",X"90",X"00",
		X"09",X"FF",X"99",X"00",X"99",X"FF",X"59",X"00",X"95",X"FF",X"55",X"00",X"95",X"FF",X"95",X"00",
		X"95",X"99",X"95",X"00",X"95",X"44",X"95",X"00",X"95",X"44",X"95",X"00",X"95",X"44",X"95",X"00",
		X"95",X"99",X"95",X"00",X"95",X"FF",X"95",X"00",X"95",X"FF",X"55",X"00",X"99",X"FF",X"59",X"00",
		X"09",X"FF",X"99",X"00",X"00",X"FF",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"55",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"90",X"99",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"90",X"00",X"00",X"09",X"90",X"00",X"00",X"09",X"90",X"00",X"00",X"09",X"90",X"00",X"00",
		X"00",X"99",X"00",X"00",X"09",X"29",X"09",X"00",X"09",X"92",X"99",X"00",X"09",X"99",X"94",X"00",
		X"09",X"A9",X"94",X"00",X"09",X"9C",X"99",X"00",X"09",X"C9",X"CC",X"00",X"09",X"C9",X"C9",X"00",
		X"D0",X"99",X"9C",X"00",X"D0",X"4C",X"99",X"00",X"00",X"CC",X"39",X"00",X"00",X"C9",X"99",X"00",
		X"90",X"99",X"90",X"00",X"99",X"39",X"00",X"00",X"55",X"39",X"00",X"00",X"55",X"39",X"90",X"00",
		X"99",X"33",X"99",X"00",X"96",X"39",X"66",X"00",X"96",X"99",X"66",X"00",X"96",X"39",X"66",X"00",
		X"66",X"99",X"66",X"90",X"22",X"22",X"22",X"99",X"22",X"22",X"22",X"99",X"99",X"22",X"99",X"99",
		X"97",X"22",X"77",X"29",X"77",X"66",X"75",X"D9",X"77",X"66",X"79",X"D9",X"79",X"66",X"9D",X"99",
		X"47",X"99",X"79",X"90",X"77",X"00",X"77",X"00",X"97",X"00",X"77",X"00",X"99",X"00",X"99",X"00",
		X"00",X"99",X"00",X"00",X"09",X"29",X"00",X"00",X"09",X"92",X"99",X"00",X"09",X"99",X"44",X"00",
		X"09",X"A9",X"54",X"00",X"09",X"CC",X"99",X"00",X"09",X"C9",X"C9",X"00",X"09",X"99",X"99",X"00",
		X"D0",X"45",X"90",X"00",X"D0",X"99",X"90",X"00",X"00",X"CC",X"90",X"00",X"00",X"C9",X"00",X"00",
		X"00",X"99",X"00",X"00",X"90",X"39",X"00",X"00",X"99",X"39",X"00",X"00",X"55",X"39",X"00",X"00",
		X"55",X"33",X"90",X"00",X"99",X"39",X"99",X"00",X"96",X"99",X"66",X"00",X"96",X"33",X"66",X"00",
		X"96",X"39",X"66",X"00",X"66",X"99",X"66",X"90",X"99",X"22",X"99",X"99",X"97",X"22",X"77",X"99",
		X"77",X"22",X"77",X"99",X"77",X"22",X"79",X"D9",X"79",X"66",X"9D",X"D9",X"79",X"66",X"99",X"69",
		X"57",X"66",X"79",X"99",X"55",X"99",X"77",X"90",X"95",X"00",X"77",X"00",X"99",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"09",X"00",X"99",X"00",
		X"09",X"99",X"EE",X"00",X"09",X"EE",X"AE",X"00",X"09",X"99",X"EE",X"00",X"09",X"EE",X"99",X"00",
		X"09",X"EE",X"EE",X"00",X"00",X"EE",X"E9",X"00",X"09",X"EE",X"99",X"00",X"99",X"EE",X"F9",X"00",
		X"9E",X"9E",X"F9",X"00",X"EE",X"9E",X"99",X"00",X"EE",X"99",X"90",X"00",X"EE",X"09",X"99",X"00",
		X"EE",X"00",X"99",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"00",X"09",X"00",X"99",X"00",X"99",X"00",X"EE",X"99",X"EE",X"00",
		X"9E",X"EE",X"AE",X"00",X"99",X"99",X"AE",X"00",X"09",X"EE",X"99",X"00",X"09",X"EE",X"E9",X"00",
		X"09",X"EE",X"E9",X"00",X"09",X"EE",X"99",X"00",X"00",X"9E",X"F9",X"00",X"00",X"9E",X"F9",X"00",
		X"00",X"9E",X"99",X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",
		X"00",X"9E",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EA",X"00",X"00",X"00",X"EA",X"00",X"00",
		X"00",X"E9",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"9F",X"00",X"00",X"09",X"9F",X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"9E",X"99",X"00",X"00",X"9E",X"9E",X"00",X"00",X"9E",X"9E",X"00",X"00",X"9E",X"99",X"00",X"00",
		X"9E",X"99",X"00",X"00",X"9E",X"E9",X"00",X"00",X"9E",X"E9",X"00",X"00",X"EE",X"99",X"00",X"00",
		X"9E",X"9E",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"40",X"00",X"00",X"90",X"90",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"99",X"00",X"99",X"D9",X"9A",X"00",X"A9",X"FD",X"99",X"90",X"AA",X"99",X"AA",X"90",
		X"99",X"99",X"2A",X"90",X"9A",X"99",X"99",X"90",X"AA",X"55",X"00",X"00",X"99",X"99",X"00",X"00",
		X"90",X"99",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"99",X"00",X"00",X"FF",X"99",X"00",X"00",
		X"0F",X"A9",X"00",X"00",X"00",X"9C",X"00",X"00",X"09",X"9C",X"00",X"00",X"09",X"99",X"00",X"00",
		X"09",X"44",X"00",X"00",X"09",X"9C",X"90",X"00",X"09",X"99",X"90",X"00",X"09",X"55",X"90",X"00",
		X"09",X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"99",X"00",X"00",
		X"09",X"29",X"00",X"00",X"09",X"22",X"00",X"00",X"09",X"22",X"00",X"00",X"09",X"22",X"90",X"00",
		X"09",X"92",X"E9",X"00",X"09",X"99",X"E9",X"00",X"09",X"09",X"E9",X"00",X"00",X"00",X"E9",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9C",X"00",X"00",
		X"00",X"9C",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"77",X"90",X"00",X"00",X"77",X"90",X"00",
		X"00",X"97",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"79",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"9C",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9C",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"2F",X"00",X"00",X"00",X"2F",X"00",X"00",X"00",X"2F",X"00",X"00",X"00",X"2F",X"00",X"00",
		X"00",X"2F",X"00",X"00",X"00",X"2F",X"00",X"00",X"00",X"2F",X"90",X"00",X"00",X"2F",X"90",X"00",
		X"00",X"9F",X"90",X"00",X"00",X"0F",X"90",X"00",X"00",X"0F",X"90",X"00",X"00",X"0F",X"90",X"00",
		X"99",X"99",X"00",X"00",X"C9",X"44",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"C9",X"00",X"00",X"90",X"C9",X"00",X"00",X"90",X"CC",X"00",X"00",X"90",X"99",X"00",X"00",
		X"99",X"CC",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"CC",X"00",X"00",X"99",X"99",X"00",X"00",
		X"92",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"29",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"96",X"00",X"00",
		X"09",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"91",X"96",X"00",X"00",X"91",X"96",X"00",X"00",
		X"91",X"99",X"00",X"00",X"91",X"91",X"00",X"00",X"99",X"91",X"00",X"00",X"09",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"9C",X"00",X"00",X"99",X"9C",X"99",X"99",X"99",X"99",X"99",X"99",
		X"00",X"92",X"90",X"00",X"00",X"92",X"90",X"00",X"00",X"92",X"90",X"00",X"00",X"92",X"00",X"00",
		X"00",X"92",X"00",X"00",X"99",X"92",X"99",X"99",X"99",X"92",X"99",X"99",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"92",X"00",X"00",
		X"00",X"22",X"90",X"00",X"00",X"22",X"90",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"69",X"00",
		X"00",X"99",X"66",X"99",X"00",X"66",X"66",X"99",X"00",X"99",X"99",X"19",X"00",X"99",X"99",X"19",
		X"00",X"66",X"09",X"99",X"00",X"66",X"00",X"90",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"00",X"00",X"97",X"99",X"00",X"00",X"77",X"99",X"00",X"00",X"74",X"99",X"90",
		X"00",X"44",X"49",X"90",X"00",X"99",X"49",X"90",X"00",X"49",X"99",X"90",X"00",X"44",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"C9",X"99",X"00",X"00",X"9C",X"99",X"90",X"00",X"99",X"29",X"90",
		X"00",X"22",X"92",X"90",X"00",X"22",X"92",X"90",X"00",X"22",X"99",X"00",X"00",X"22",X"29",X"00",
		X"00",X"22",X"29",X"00",X"00",X"22",X"29",X"00",X"00",X"22",X"99",X"00",X"00",X"29",X"99",X"00",
		X"00",X"99",X"69",X"00",X"00",X"66",X"69",X"00",X"00",X"69",X"69",X"00",X"00",X"66",X"69",X"00",
		X"00",X"96",X"99",X"00",X"00",X"96",X"11",X"00",X"00",X"96",X"11",X"00",X"00",X"96",X"99",X"00",
		X"00",X"99",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"99",X"99",X"00",
		X"99",X"99",X"00",X"00",X"9C",X"44",X"00",X"00",X"9C",X"44",X"99",X"99",X"99",X"94",X"99",X"99",
		X"09",X"A9",X"09",X"00",X"09",X"99",X"09",X"00",X"09",X"CC",X"09",X"00",X"09",X"C4",X"09",X"00",
		X"09",X"94",X"09",X"00",X"99",X"CC",X"99",X"99",X"99",X"99",X"99",X"99",X"00",X"92",X"00",X"00",
		X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"92",X"00",X"00",
		X"00",X"92",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"69",X"00",X"00",X"09",X"99",X"00",X"00",
		X"09",X"19",X"00",X"00",X"09",X"19",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"00",X"66",X"00",X"44",X"00",X"66",X"00",X"44",X"00",X"66",X"00",X"44",X"00",X"99",X"00",
		X"99",X"00",X"77",X"00",X"EE",X"90",X"77",X"00",X"EE",X"90",X"77",X"00",X"4C",X"90",X"99",X"00",
		X"49",X"00",X"09",X"00",X"CC",X"00",X"90",X"00",X"9C",X"00",X"99",X"00",X"99",X"00",X"11",X"00",
		X"99",X"00",X"99",X"00",X"59",X"00",X"90",X"00",X"55",X"00",X"00",X"00",X"95",X"90",X"00",X"00",
		X"99",X"99",X"09",X"00",X"59",X"9C",X"99",X"00",X"55",X"CC",X"99",X"99",X"55",X"CC",X"77",X"49",
		X"99",X"99",X"44",X"49",X"11",X"00",X"44",X"49",X"11",X"09",X"44",X"99",X"11",X"99",X"44",X"90",
		X"11",X"99",X"94",X"00",X"99",X"99",X"99",X"00",X"00",X"99",X"09",X"00",X"00",X"99",X"09",X"00",
		X"00",X"99",X"09",X"00",X"00",X"90",X"09",X"00",X"90",X"00",X"09",X"00",X"90",X"00",X"00",X"00",
		X"99",X"00",X"09",X"99",X"44",X"00",X"97",X"79",X"44",X"00",X"77",X"79",X"44",X"90",X"77",X"79",
		X"99",X"90",X"77",X"79",X"EE",X"99",X"77",X"99",X"EE",X"C9",X"99",X"00",X"44",X"99",X"00",X"00",
		X"44",X"00",X"00",X"00",X"CC",X"00",X"90",X"99",X"99",X"00",X"99",X"39",X"59",X"00",X"33",X"19",
		X"59",X"00",X"11",X"39",X"55",X"00",X"99",X"99",X"95",X"90",X"00",X"00",X"95",X"99",X"99",X"00",
		X"99",X"9C",X"99",X"90",X"55",X"CC",X"99",X"99",X"55",X"CC",X"77",X"49",X"99",X"99",X"44",X"49",
		X"11",X"00",X"44",X"49",X"11",X"00",X"44",X"99",X"11",X"00",X"44",X"90",X"11",X"00",X"94",X"00",
		X"11",X"00",X"99",X"00",X"91",X"00",X"09",X"00",X"91",X"00",X"99",X"00",X"11",X"00",X"95",X"00",
		X"11",X"00",X"95",X"00",X"99",X"00",X"95",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"09",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"9A",X"99",X"00",
		X"00",X"92",X"99",X"00",X"99",X"99",X"CC",X"00",X"9C",X"CC",X"9C",X"00",X"9C",X"CC",X"CC",X"00",
		X"CC",X"99",X"99",X"00",X"C9",X"99",X"C9",X"00",X"99",X"99",X"99",X"00",X"99",X"CC",X"90",X"00",
		X"09",X"9C",X"99",X"00",X"00",X"99",X"49",X"00",X"00",X"49",X"44",X"00",X"00",X"44",X"94",X"00",
		X"00",X"44",X"94",X"00",X"00",X"44",X"94",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"49",X"00",
		X"00",X"44",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"22",X"29",X"00",X"09",X"22",X"29",X"00",
		X"09",X"92",X"29",X"00",X"09",X"99",X"29",X"00",X"09",X"99",X"99",X"00",X"00",X"29",X"29",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"11",X"00",X"00",X"90",X"11",X"00",X"00",X"90",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9F",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"9F",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"A9",X"00",X"00",
		X"00",X"A9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"79",X"00",X"00",X"09",X"99",X"00",X"00",
		X"99",X"97",X"00",X"00",X"9C",X"99",X"00",X"00",X"9C",X"94",X"00",X"00",X"99",X"99",X"00",X"00",
		X"00",X"77",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"DD",X"99",X"00",X"00",X"9D",X"D9",X"00",
		X"00",X"99",X"D9",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",
		X"00",X"00",X"D9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
