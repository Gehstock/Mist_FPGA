library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_SND_2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_SND_2 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"21",X"50",X"80",X"C3",X"70",X"0D",X"DD",X"21",X"58",X"80",X"C3",X"70",X"0D",X"CD",X"5C",X"07",
		X"3E",X"01",X"32",X"A0",X"80",X"3E",X"20",X"32",X"A1",X"80",X"3E",X"10",X"32",X"A2",X"80",X"AF",
		X"32",X"A5",X"80",X"32",X"A6",X"80",X"21",X"00",X"01",X"22",X"A3",X"80",X"21",X"00",X"05",X"22",
		X"A7",X"80",X"CD",X"B3",X"04",X"CD",X"FA",X"04",X"06",X"0D",X"CD",X"D8",X"05",X"C9",X"2A",X"A3",
		X"80",X"2B",X"7C",X"B5",X"28",X"5C",X"22",X"A3",X"80",X"3A",X"A5",X"80",X"B7",X"28",X"06",X"FE",
		X"01",X"28",X"24",X"AF",X"C9",X"21",X"A0",X"80",X"35",X"20",X"F8",X"36",X"01",X"CD",X"5A",X"06",
		X"B7",X"11",X"04",X"00",X"ED",X"52",X"CD",X"B3",X"04",X"21",X"A1",X"80",X"35",X"20",X"E4",X"36",
		X"20",X"21",X"A5",X"80",X"34",X"18",X"DC",X"2A",X"A7",X"80",X"11",X"50",X"00",X"3A",X"A6",X"80",
		X"E6",X"01",X"20",X"1B",X"B7",X"ED",X"52",X"22",X"A7",X"80",X"CD",X"B3",X"04",X"21",X"A2",X"80",
		X"35",X"20",X"06",X"36",X"10",X"21",X"A6",X"80",X"34",X"21",X"A5",X"80",X"35",X"18",X"B4",X"19",
		X"18",X"E5",X"3E",X"FF",X"C9",X"CD",X"A1",X"06",X"3E",X"18",X"32",X"B0",X"80",X"21",X"00",X"01",
		X"22",X"B1",X"80",X"AF",X"32",X"B3",X"80",X"21",X"00",X"02",X"22",X"B4",X"80",X"16",X"06",X"1E",
		X"00",X"CD",X"34",X"05",X"CD",X"68",X"05",X"06",X"03",X"CD",X"D8",X"05",X"C9",X"2A",X"B4",X"80",
		X"2B",X"7C",X"B5",X"28",X"4B",X"22",X"B4",X"80",X"3A",X"B3",X"80",X"FE",X"00",X"28",X"1B",X"2A",
		X"B1",X"80",X"2B",X"7C",X"B5",X"20",X"34",X"21",X"00",X"01",X"22",X"B1",X"80",X"16",X"06",X"1E",
		X"00",X"CD",X"34",X"05",X"AF",X"32",X"B3",X"80",X"AF",X"C9",X"21",X"B0",X"80",X"35",X"20",X"F8",
		X"36",X"18",X"16",X"06",X"CD",X"0F",X"06",X"1C",X"7B",X"FE",X"08",X"28",X"05",X"CD",X"34",X"05",
		X"18",X"E6",X"CD",X"34",X"05",X"21",X"B3",X"80",X"34",X"18",X"DD",X"22",X"B1",X"80",X"18",X"D8",
		X"3E",X"FF",X"C9",X"CD",X"96",X"07",X"3E",X"01",X"32",X"C0",X"80",X"21",X"00",X"08",X"22",X"C3",
		X"80",X"AF",X"32",X"C5",X"80",X"21",X"00",X"02",X"22",X"C6",X"80",X"21",X"00",X"05",X"CD",X"B3",
		X"04",X"CD",X"FA",X"04",X"06",X"08",X"CD",X"D8",X"05",X"C9",X"2A",X"C6",X"80",X"2B",X"7C",X"B5",
		X"28",X"43",X"22",X"C6",X"80",X"21",X"C0",X"80",X"35",X"20",X"2C",X"36",X"01",X"CD",X"5A",X"06",
		X"11",X"08",X"00",X"19",X"ED",X"5B",X"C3",X"80",X"7C",X"BA",X"20",X"18",X"7D",X"BB",X"20",X"14",
		X"3A",X"C5",X"80",X"B7",X"20",X"13",X"21",X"00",X"0B",X"22",X"C3",X"80",X"3E",X"FF",X"32",X"C5",
		X"80",X"21",X"00",X"05",X"CD",X"B3",X"04",X"AF",X"C9",X"21",X"00",X"08",X"22",X"C3",X"80",X"AF",
		X"32",X"C5",X"80",X"18",X"EC",X"3E",X"FF",X"C9",X"CD",X"22",X"07",X"3E",X"08",X"32",X"D0",X"80",
		X"3E",X"05",X"32",X"D1",X"80",X"3E",X"0C",X"32",X"D2",X"80",X"AF",X"32",X"D3",X"80",X"21",X"50",
		X"00",X"CD",X"B3",X"04",X"CD",X"FA",X"04",X"06",X"00",X"CD",X"D8",X"05",X"C9",X"3A",X"D3",X"80",
		X"FE",X"00",X"28",X"18",X"FE",X"01",X"28",X"26",X"FE",X"02",X"28",X"27",X"FE",X"03",X"28",X"33",
		X"21",X"D2",X"80",X"35",X"28",X"32",X"AF",X"32",X"D3",X"80",X"AF",X"C9",X"CD",X"25",X"06",X"3C",
		X"FE",X"0A",X"20",X"04",X"21",X"D3",X"80",X"34",X"47",X"CD",X"D8",X"05",X"18",X"EC",X"CD",X"0B",
		X"12",X"18",X"E7",X"CD",X"25",X"06",X"3D",X"20",X"04",X"21",X"D3",X"80",X"34",X"47",X"CD",X"D8",
		X"05",X"18",X"D7",X"CD",X"18",X"12",X"18",X"D2",X"3E",X"FF",X"C9",X"21",X"D0",X"80",X"35",X"C0",
		X"3E",X"08",X"77",X"21",X"D3",X"80",X"34",X"C9",X"21",X"D1",X"80",X"35",X"C0",X"3E",X"05",X"77",
		X"21",X"D3",X"80",X"34",X"C9",X"00",X"01",X"04",X"00",X"80",X"00",X"04",X"00",X"00",X"02",X"08",
		X"08",X"00",X"20",X"21",X"2F",X"12",X"11",X"00",X"81",X"01",X"04",X"00",X"ED",X"B0",X"CD",X"96",
		X"07",X"CD",X"FA",X"04",X"2A",X"25",X"12",X"CD",X"B3",X"04",X"3E",X"0D",X"47",X"C3",X"D8",X"05",
		X"DD",X"E5",X"FD",X"E5",X"DD",X"21",X"00",X"81",X"FD",X"21",X"2F",X"12",X"CD",X"75",X"12",X"CD",
		X"5A",X"06",X"22",X"18",X"81",X"CD",X"CA",X"12",X"AF",X"FD",X"E1",X"DD",X"E1",X"21",X"02",X"81",
		X"CB",X"4E",X"C8",X"3D",X"C9",X"DD",X"CB",X"02",X"46",X"C2",X"A3",X"12",X"C3",X"7F",X"12",X"DD",
		X"35",X"00",X"C0",X"FD",X"7E",X"00",X"DD",X"77",X"00",X"CD",X"5A",X"06",X"ED",X"5B",X"27",X"12",
		X"B7",X"ED",X"52",X"CD",X"B3",X"04",X"EB",X"2A",X"29",X"12",X"B7",X"ED",X"52",X"D8",X"DD",X"CB",
		X"02",X"C6",X"C9",X"DD",X"35",X"01",X"C0",X"FD",X"7E",X"01",X"DD",X"77",X"01",X"CD",X"5A",X"06",
		X"ED",X"5B",X"2B",X"12",X"19",X"CD",X"B3",X"04",X"ED",X"5B",X"2D",X"12",X"B7",X"ED",X"52",X"D8",
		X"DD",X"CB",X"02",X"86",X"2A",X"25",X"12",X"C3",X"B3",X"04",X"DD",X"35",X"03",X"C0",X"FD",X"7E",
		X"03",X"DD",X"77",X"03",X"CD",X"25",X"06",X"3D",X"47",X"CD",X"D8",X"05",X"78",X"B7",X"C0",X"DD",
		X"CB",X"02",X"CE",X"C9",X"DD",X"35",X"03",X"C0",X"FD",X"7E",X"03",X"DD",X"77",X"03",X"CD",X"25",
		X"06",X"3C",X"47",X"CD",X"D8",X"05",X"FE",X"0C",X"C0",X"DD",X"CB",X"02",X"CE",X"06",X"00",X"C3",
		X"D8",X"05",X"21",X"1E",X"13",X"11",X"10",X"81",X"01",X"04",X"00",X"ED",X"B0",X"CD",X"96",X"07",
		X"CD",X"FA",X"04",X"2A",X"18",X"81",X"CD",X"B3",X"04",X"06",X"03",X"C3",X"D8",X"05",X"08",X"08",
		X"01",X"30",X"DD",X"E5",X"FD",X"E5",X"DD",X"21",X"10",X"81",X"FD",X"21",X"1E",X"13",X"CD",X"75",
		X"12",X"CD",X"E4",X"12",X"AF",X"FD",X"E1",X"DD",X"E1",X"21",X"12",X"81",X"CB",X"4E",X"C8",X"3D",
		X"C9",X"CD",X"A1",X"06",X"AF",X"32",X"24",X"81",X"3E",X"02",X"32",X"23",X"81",X"CD",X"FA",X"04",
		X"3E",X"08",X"32",X"20",X"81",X"21",X"20",X"00",X"22",X"21",X"81",X"21",X"80",X"00",X"CD",X"B3",
		X"04",X"06",X"08",X"CD",X"D8",X"05",X"C9",X"3A",X"24",X"81",X"B7",X"20",X"0B",X"2A",X"21",X"81",
		X"2B",X"7C",X"B5",X"28",X"37",X"22",X"21",X"81",X"21",X"20",X"81",X"35",X"28",X"1A",X"CD",X"5A",
		X"06",X"11",X"20",X"00",X"19",X"11",X"00",X"05",X"7C",X"BA",X"20",X"07",X"7D",X"BB",X"20",X"03",
		X"21",X"80",X"00",X"CD",X"B3",X"04",X"AF",X"C9",X"3E",X"08",X"32",X"20",X"81",X"CD",X"25",X"06",
		X"3D",X"28",X"06",X"47",X"CD",X"D8",X"05",X"18",X"D5",X"3E",X"FF",X"C9",X"21",X"20",X"00",X"22",
		X"21",X"81",X"21",X"23",X"81",X"35",X"20",X"05",X"3E",X"01",X"32",X"24",X"81",X"CD",X"50",X"13",
		X"18",X"A5",X"00",X"04",X"00",X"01",X"01",X"20",X"01",X"00",X"01",X"20",X"01",X"21",X"C2",X"13",
		X"11",X"85",X"80",X"01",X"0B",X"00",X"ED",X"B0",X"CD",X"96",X"07",X"2A",X"C2",X"13",X"CD",X"B3",
		X"04",X"CD",X"FA",X"04",X"06",X"0D",X"C3",X"D8",X"05",X"2A",X"87",X"80",X"2B",X"22",X"87",X"80",
		X"7D",X"B4",X"3E",X"FF",X"C8",X"DD",X"E5",X"DD",X"21",X"85",X"80",X"DD",X"CB",X"07",X"46",X"CD",
		X"05",X"14",X"DD",X"E1",X"C9",X"CA",X"0B",X"14",X"C3",X"33",X"14",X"AF",X"DD",X"35",X"04",X"C0",
		X"DD",X"7E",X"08",X"DD",X"77",X"04",X"CD",X"5A",X"06",X"B7",X"11",X"08",X"00",X"ED",X"52",X"CD",
		X"B3",X"04",X"AF",X"DD",X"35",X"05",X"C0",X"DD",X"7E",X"09",X"DD",X"77",X"05",X"DD",X"CB",X"07",
		X"C6",X"AF",X"C9",X"2A",X"85",X"80",X"11",X"30",X"00",X"DD",X"CB",X"07",X"4E",X"20",X"04",X"B7",
		X"ED",X"52",X"06",X"19",X"22",X"85",X"80",X"CD",X"B3",X"04",X"DD",X"35",X"06",X"20",X"0E",X"DD",
		X"7E",X"0A",X"DD",X"77",X"06",X"3E",X"02",X"DD",X"AE",X"07",X"DD",X"77",X"07",X"DD",X"CB",X"07",
		X"86",X"AF",X"DD",X"CB",X"07",X"56",X"C8",X"DD",X"CB",X"07",X"8E",X"C9",X"21",X"7A",X"14",X"11",
		X"85",X"80",X"01",X"0B",X"00",X"ED",X"B0",X"C3",X"D8",X"13",X"00",X"03",X"E0",X"00",X"01",X"10",
		X"01",X"04",X"01",X"10",X"01",X"80",X"01",X"20",X"00",X"00",X"10",X"10",X"00",X"00",X"02",X"00",
		X"02",X"08",X"08",X"10",X"10",X"00",X"04",X"0F",X"0F",X"21",X"8F",X"14",X"11",X"60",X"81",X"01",
		X"07",X"00",X"ED",X"B0",X"CD",X"5C",X"07",X"CD",X"FA",X"04",X"2A",X"85",X"14",X"CD",X"B3",X"04",
		X"3A",X"97",X"14",X"47",X"C3",X"D8",X"05",X"2A",X"60",X"81",X"2B",X"22",X"60",X"81",X"7D",X"B4",
		X"3E",X"FF",X"C8",X"DD",X"E5",X"FD",X"E5",X"DD",X"21",X"60",X"81",X"FD",X"21",X"8F",X"14",X"CD",
		X"DB",X"14",X"CD",X"E5",X"14",X"FD",X"E1",X"DD",X"E1",X"AF",X"C9",X"DD",X"CB",X"06",X"46",X"C2",
		X"13",X"15",X"C3",X"EF",X"14",X"DD",X"CB",X"06",X"4E",X"CA",X"3A",X"15",X"C3",X"55",X"15",X"DD",
		X"35",X"02",X"C0",X"FD",X"7E",X"02",X"DD",X"77",X"02",X"CD",X"5A",X"06",X"ED",X"5B",X"87",X"14",
		X"B7",X"ED",X"52",X"CD",X"B3",X"04",X"EB",X"B7",X"2A",X"89",X"14",X"ED",X"52",X"D8",X"DD",X"CB",
		X"06",X"C6",X"C9",X"DD",X"35",X"03",X"C0",X"FD",X"7E",X"03",X"DD",X"77",X"03",X"CD",X"5A",X"06",
		X"ED",X"5B",X"8B",X"14",X"19",X"CD",X"B3",X"04",X"ED",X"5B",X"8D",X"14",X"B7",X"ED",X"52",X"D8",
		X"DD",X"CB",X"06",X"86",X"2A",X"85",X"14",X"C3",X"B3",X"04",X"DD",X"35",X"04",X"C0",X"FD",X"7E",
		X"04",X"DD",X"77",X"04",X"CD",X"25",X"06",X"3D",X"47",X"CD",X"D8",X"05",X"FD",X"BE",X"07",X"C0",
		X"DD",X"CB",X"06",X"CE",X"C9",X"DD",X"35",X"05",X"C0",X"FD",X"7E",X"05",X"DD",X"77",X"05",X"CD",
		X"25",X"06",X"3C",X"47",X"CD",X"D8",X"05",X"FD",X"BE",X"09",X"C0",X"DD",X"CB",X"06",X"8E",X"FD",
		X"46",X"08",X"C3",X"D8",X"05",X"1F",X"0F",X"3F",X"0F",X"5F",X"0A",X"82",X"83",X"82",X"85",X"82",
		X"83",X"82",X"85",X"82",X"83",X"82",X"85",X"82",X"83",X"82",X"85",X"8E",X"8F",X"8E",X"91",X"8E",
		X"8F",X"8E",X"91",X"8E",X"8F",X"8E",X"91",X"8E",X"8F",X"8E",X"91",X"FF",X"1F",X"01",X"3F",X"0F",
		X"5F",X"0A",X"84",X"85",X"84",X"87",X"84",X"85",X"84",X"87",X"84",X"85",X"84",X"87",X"84",X"85",
		X"84",X"87",X"90",X"91",X"90",X"93",X"90",X"91",X"90",X"93",X"90",X"91",X"90",X"93",X"90",X"91",
		X"90",X"93",X"FF",X"FF",X"1F",X"0E",X"3F",X"0F",X"5F",X"09",X"A2",X"A6",X"A9",X"89",X"89",X"8B",
		X"8D",X"8E",X"90",X"B2",X"AE",X"B3",X"93",X"93",X"B2",X"95",X"93",X"B2",X"B0",X"AE",X"A0",X"FF",
		X"1F",X"0E",X"3F",X"0F",X"5F",X"09",X"A2",X"A6",X"A9",X"89",X"89",X"8B",X"8D",X"8E",X"90",X"B2",
		X"AE",X"AE",X"8E",X"8E",X"AE",X"8D",X"8E",X"AD",X"AB",X"A9",X"FF",X"1F",X"07",X"3F",X"0F",X"5F",
		X"09",X"A2",X"A6",X"A9",X"89",X"89",X"8B",X"8D",X"8E",X"90",X"B2",X"AE",X"AB",X"8B",X"8B",X"A9",
		X"89",X"8B",X"A9",X"A7",X"A6",X"A0",X"FF",X"1F",X"0E",X"3F",X"0F",X"5F",X"0B",X"94",X"8D",X"96",
		X"8D",X"94",X"8D",X"96",X"8D",X"94",X"99",X"98",X"96",X"B4",X"B2",X"94",X"8D",X"96",X"8D",X"94",
		X"8D",X"96",X"8D",X"94",X"99",X"98",X"96",X"B4",X"B2",X"94",X"8D",X"96",X"8D",X"94",X"8D",X"96",
		X"8D",X"94",X"99",X"98",X"96",X"B4",X"B2",X"D1",X"CF",X"CD",X"FF",X"1F",X"08",X"3F",X"0F",X"5F",
		X"0A",X"A8",X"AA",X"A8",X"AA",X"E8",X"A8",X"AA",X"A8",X"AA",X"E8",X"A8",X"AA",X"A8",X"AA",X"E8",
		X"C8",X"C6",X"C5",X"FF",X"1F",X"08",X"3F",X"0F",X"5F",X"0A",X"A5",X"A6",X"A5",X"A6",X"E5",X"A5",
		X"A6",X"A5",X"A6",X"E5",X"A5",X"A6",X"A5",X"A6",X"E5",X"C5",X"C3",X"C1",X"FF",X"02",X"02",X"00",
		X"00",X"1F",X"2A",X"7D",X"16",X"22",X"90",X"80",X"3A",X"7F",X"16",X"32",X"92",X"80",X"CD",X"22",
		X"07",X"CD",X"68",X"05",X"3A",X"81",X"16",X"5F",X"16",X"06",X"CD",X"34",X"05",X"3A",X"80",X"16",
		X"47",X"CD",X"D8",X"05",X"C9",X"21",X"90",X"80",X"11",X"7D",X"16",X"CD",X"BB",X"16",X"CD",X"DE",
		X"16",X"AF",X"C9",X"3A",X"92",X"80",X"A9",X"32",X"92",X"80",X"C9",X"3A",X"92",X"80",X"CB",X"47",
		X"28",X"0D",X"35",X"C0",X"1A",X"77",X"06",X"02",X"CD",X"D8",X"05",X"0E",X"01",X"18",X"E4",X"23",
		X"13",X"35",X"C0",X"1A",X"77",X"06",X"08",X"CD",X"D8",X"05",X"0E",X"01",X"18",X"D5",X"16",X"06",
		X"CD",X"0F",X"06",X"3A",X"92",X"80",X"CB",X"4F",X"28",X"0B",X"1C",X"7B",X"FE",X"01",X"0E",X"02",
		X"28",X"C1",X"C3",X"34",X"05",X"1D",X"7B",X"FE",X"15",X"0E",X"02",X"28",X"B6",X"C3",X"34",X"05",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
