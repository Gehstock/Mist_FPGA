library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity spy_hunter_ch_bits is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of spy_hunter_ch_bits is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"3F",X"3F",X"0C",X"0C",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"0C",X"0C",X"3F",X"3F",
		X"00",X"00",X"3F",X"3F",X"0C",X"0C",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"0C",X"0C",X"3F",X"3F",
		X"00",X"00",X"3F",X"FC",X"C0",X"03",X"CC",X"33",X"CC",X"33",X"CF",X"F3",X"C0",X"03",X"3F",X"FC",
		X"33",X"00",X"3F",X"FC",X"00",X"00",X"03",X"FC",X"3F",X"0C",X"33",X"0C",X"3F",X"FC",X"00",X"00",
		X"00",X"0C",X"3F",X"FC",X"00",X"00",X"00",X"0C",X"00",X"0C",X"3F",X"FC",X"00",X"00",X"3F",X"FC",
		X"00",X"00",X"F0",X"00",X"0F",X"C0",X"00",X"3F",X"3C",X"00",X"0F",X"FC",X"3C",X"00",X"00",X"0C",
		X"00",X"00",X"3F",X"FC",X"00",X"00",X"3F",X"FC",X"0C",X"00",X"03",X"00",X"0C",X"00",X"3F",X"FC",
		X"00",X"0C",X"00",X"30",X"00",X"0C",X"3F",X"F0",X"00",X"00",X"0F",X"F0",X"30",X"0C",X"3F",X"FC",
		X"0F",X"FC",X"3C",X"00",X"00",X"00",X"3F",X"FC",X"33",X"00",X"3F",X"FC",X"00",X"00",X"3F",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"00",
		X"15",X"54",X"00",X"00",X"15",X"54",X"10",X"44",X"15",X"44",X"00",X"00",X"15",X"54",X"00",X"00",
		X"00",X"00",X"00",X"00",X"15",X"54",X"11",X"04",X"11",X"04",X"00",X"00",X"15",X"54",X"11",X"04",
		X"00",X"00",X"00",X"00",X"2A",X"A0",X"A0",X"28",X"80",X"08",X"A0",X"28",X"2A",X"A8",X"0A",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"08",X"AA",X"A8",X"2A",X"A8",X"08",X"08",X"00",X"08",
		X"00",X"00",X"00",X"00",X"28",X"08",X"AA",X"08",X"A2",X"88",X"80",X"A8",X"A0",X"A8",X"A0",X"28",
		X"00",X"00",X"00",X"00",X"00",X"A8",X"A8",X"A8",X"82",X"88",X"82",X"08",X"A0",X"28",X"A0",X"28",
		X"00",X"00",X"00",X"00",X"AA",X"A8",X"AA",X"A8",X"02",X"80",X"A2",X"80",X"2A",X"80",X"02",X"80",
		X"00",X"00",X"00",X"00",X"80",X"A8",X"82",X"A8",X"82",X"08",X"82",X"08",X"AA",X"08",X"AA",X"08",
		X"00",X"00",X"00",X"00",X"20",X"A8",X"82",X"88",X"82",X"08",X"A2",X"08",X"2A",X"A8",X"0A",X"A8",
		X"00",X"00",X"00",X"00",X"A8",X"00",X"AA",X"00",X"82",X"80",X"80",X"A0",X"80",X"28",X"A0",X"08",
		X"00",X"00",X"00",X"00",X"28",X"A8",X"AA",X"A8",X"82",X"08",X"AA",X"08",X"2A",X"A8",X"00",X"A8",
		X"00",X"00",X"00",X"00",X"2A",X"A0",X"AA",X"A8",X"82",X"08",X"82",X"80",X"AA",X"80",X"2A",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"FC",X"00",X"FF",X"00",X"0F",X"C0",X"00",X"F0",X"00",X"03",X"00",X"0F",X"00",X"00",
		X"FF",X"FF",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"FF",X"FF",
		X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"FF",X"FF",
		X"FF",X"FF",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"FF",X"FF",
		X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FC",X"00",X"0F",X"C0",X"00",X"FC",X"00",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"3F",X"F0",X"F0",X"3C",X"C0",X"0C",X"F0",X"3C",X"3F",X"FC",X"0F",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"0C",X"FF",X"FC",X"3F",X"FC",X"0C",X"0C",X"00",X"0C",
		X"00",X"00",X"00",X"00",X"3C",X"0C",X"FF",X"0C",X"F3",X"CC",X"C0",X"FC",X"F0",X"FC",X"F0",X"3C",
		X"00",X"00",X"00",X"00",X"00",X"FC",X"FC",X"FC",X"C3",X"CC",X"C3",X"0C",X"F0",X"3C",X"F0",X"3C",
		X"00",X"00",X"00",X"00",X"FF",X"FC",X"FF",X"FC",X"03",X"C0",X"F3",X"C0",X"3F",X"C0",X"03",X"C0",
		X"00",X"00",X"00",X"00",X"C0",X"FC",X"C3",X"FC",X"C3",X"0C",X"C3",X"0C",X"FF",X"0C",X"FF",X"0C",
		X"00",X"00",X"00",X"00",X"30",X"FC",X"C3",X"CC",X"C3",X"0C",X"F3",X"0C",X"3F",X"FC",X"0F",X"FC",
		X"00",X"00",X"00",X"00",X"FC",X"00",X"FF",X"00",X"C3",X"C0",X"C0",X"F0",X"C0",X"3C",X"F0",X"0C",
		X"00",X"00",X"00",X"00",X"3C",X"FC",X"FF",X"FC",X"C3",X"0C",X"FF",X"0C",X"3F",X"FC",X"00",X"FC",
		X"00",X"00",X"00",X"00",X"3F",X"F0",X"FF",X"FC",X"C3",X"0C",X"C3",X"C0",X"FF",X"C0",X"3F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"FF",X"30",X"03",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"F3",X"30",X"03",X"3F",X"FF",
		X"00",X"00",X"00",X"0C",X"3F",X"FC",X"F0",X"C0",X"C0",X"C0",X"FF",X"FC",X"3F",X"FC",X"00",X"0C",
		X"00",X"00",X"00",X"00",X"FC",X"FC",X"FF",X"FC",X"C3",X"0C",X"FF",X"FC",X"FF",X"FC",X"C0",X"0C",
		X"00",X"00",X"00",X"00",X"30",X"3C",X"C0",X"0C",X"C0",X"0C",X"F0",X"3C",X"3F",X"FC",X"0F",X"F0",
		X"00",X"00",X"00",X"00",X"3F",X"F0",X"F0",X"3C",X"C0",X"0C",X"FF",X"FC",X"FF",X"FC",X"C0",X"0C",
		X"00",X"00",X"00",X"00",X"F0",X"3C",X"C0",X"0C",X"CF",X"0C",X"FF",X"FC",X"FF",X"FC",X"C0",X"0C",
		X"00",X"00",X"00",X"00",X"F0",X"00",X"C0",X"00",X"CF",X"0C",X"FF",X"FC",X"FF",X"FC",X"C0",X"0C",
		X"00",X"00",X"00",X"C0",X"30",X"FC",X"C0",X"CC",X"C0",X"0C",X"F0",X"3C",X"3F",X"FC",X"0F",X"F0",
		X"00",X"00",X"C0",X"00",X"FF",X"FC",X"0F",X"00",X"0F",X"00",X"FF",X"FC",X"FF",X"FC",X"C0",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"C0",X"0C",X"FF",X"FC",X"FF",X"FC",X"C0",X"0C",X"00",X"0C",
		X"00",X"00",X"C0",X"00",X"FF",X"FC",X"C0",X"3C",X"C0",X"0C",X"00",X"0C",X"00",X"FC",X"00",X"F0",
		X"00",X"00",X"F0",X"0C",X"FC",X"3C",X"0C",X"F0",X"03",X"00",X"FF",X"FC",X"FF",X"FC",X"C0",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"3C",X"00",X"0C",X"C0",X"0C",X"FF",X"FC",X"FF",X"FC",X"C0",X"00",
		X"00",X"00",X"C0",X"0C",X"FF",X"FC",X"3C",X"00",X"0F",X"00",X"3C",X"00",X"FF",X"FC",X"FF",X"FC",
		X"00",X"00",X"C0",X"00",X"FF",X"FC",X"00",X"F0",X"0F",X"00",X"3C",X"00",X"FF",X"FC",X"FF",X"FC",
		X"00",X"00",X"00",X"00",X"3F",X"F0",X"F0",X"3C",X"C0",X"0C",X"F0",X"3C",X"3F",X"FC",X"0F",X"F0",
		X"00",X"00",X"00",X"00",X"3F",X"C0",X"F3",X"C0",X"C0",X"C0",X"FF",X"FC",X"FF",X"FC",X"C0",X"0C",
		X"00",X"00",X"00",X"00",X"3F",X"CC",X"F0",X"30",X"C0",X"CC",X"F0",X"0C",X"3F",X"FC",X"0F",X"F0",
		X"00",X"00",X"00",X"0C",X"FC",X"3C",X"CF",X"F0",X"C3",X"C0",X"FF",X"FC",X"FF",X"FC",X"C0",X"0C",
		X"00",X"00",X"00",X"00",X"30",X"F0",X"C3",X"FC",X"C3",X"0C",X"FF",X"0C",X"FF",X"3C",X"3C",X"3C",
		X"00",X"00",X"00",X"00",X"F0",X"00",X"C0",X"00",X"FF",X"FC",X"FF",X"FC",X"C0",X"0C",X"F0",X"00",
		X"00",X"00",X"C0",X"00",X"FF",X"FC",X"00",X"0C",X"00",X"0C",X"FF",X"FC",X"FF",X"FC",X"C0",X"00",
		X"00",X"00",X"C0",X"00",X"FC",X"00",X"0F",X"F0",X"00",X"3C",X"0F",X"FC",X"FF",X"C0",X"F0",X"00",
		X"00",X"00",X"F0",X"00",X"3F",X"FC",X"00",X"3C",X"03",X"F0",X"00",X"3C",X"FF",X"FC",X"F0",X"00",
		X"00",X"00",X"C0",X"00",X"F0",X"0C",X"3F",X"3C",X"03",X"C0",X"0F",X"F0",X"FC",X"3C",X"F0",X"0C",
		X"00",X"00",X"C0",X"00",X"FF",X"00",X"03",X"FC",X"03",X"FC",X"FF",X"00",X"FF",X"00",X"F0",X"00",
		X"00",X"00",X"F0",X"00",X"FC",X"0C",X"CF",X"0C",X"C3",X"CC",X"C0",X"FC",X"F0",X"3C",X"00",X"0C",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"08",X"2A",X"A8",X"A0",X"80",X"80",X"80",X"AA",X"A8",X"2A",X"A8",X"00",X"08",
		X"00",X"00",X"00",X"00",X"A8",X"A8",X"AA",X"A8",X"82",X"08",X"AA",X"A8",X"AA",X"A8",X"80",X"08",
		X"00",X"00",X"00",X"00",X"20",X"28",X"80",X"08",X"80",X"08",X"A0",X"28",X"2A",X"A8",X"0A",X"A0",
		X"00",X"00",X"00",X"00",X"2A",X"A0",X"A0",X"28",X"80",X"08",X"AA",X"A8",X"AA",X"A8",X"80",X"08",
		X"00",X"00",X"00",X"00",X"A0",X"28",X"80",X"08",X"8A",X"08",X"AA",X"A8",X"AA",X"A8",X"80",X"08",
		X"00",X"00",X"00",X"00",X"A0",X"00",X"80",X"00",X"8A",X"08",X"AA",X"A8",X"AA",X"A8",X"80",X"08",
		X"00",X"00",X"00",X"80",X"20",X"A8",X"80",X"88",X"80",X"08",X"A0",X"28",X"2A",X"A8",X"0A",X"A0",
		X"00",X"00",X"80",X"00",X"AA",X"A8",X"0A",X"00",X"0A",X"00",X"AA",X"A8",X"AA",X"A8",X"80",X"08",
		X"00",X"00",X"00",X"00",X"00",X"08",X"80",X"08",X"AA",X"A8",X"AA",X"A8",X"80",X"08",X"00",X"08",
		X"00",X"00",X"80",X"00",X"AA",X"A8",X"80",X"28",X"80",X"08",X"00",X"08",X"00",X"A8",X"00",X"A0",
		X"00",X"00",X"A0",X"08",X"A8",X"28",X"08",X"A0",X"02",X"00",X"AA",X"A8",X"AA",X"A8",X"80",X"08",
		X"00",X"00",X"00",X"00",X"00",X"28",X"00",X"08",X"80",X"08",X"AA",X"A8",X"AA",X"A8",X"80",X"00",
		X"00",X"00",X"80",X"08",X"AA",X"A8",X"28",X"00",X"0A",X"00",X"28",X"00",X"AA",X"A8",X"AA",X"A8",
		X"00",X"00",X"80",X"00",X"AA",X"A8",X"00",X"A0",X"0A",X"00",X"28",X"00",X"AA",X"A8",X"AA",X"A8",
		X"00",X"00",X"00",X"00",X"2A",X"A0",X"A0",X"28",X"80",X"08",X"A0",X"28",X"2A",X"A8",X"0A",X"A0",
		X"00",X"00",X"00",X"00",X"2A",X"80",X"A2",X"80",X"80",X"80",X"AA",X"A8",X"AA",X"A8",X"80",X"08",
		X"00",X"00",X"00",X"00",X"2A",X"88",X"A0",X"20",X"80",X"88",X"A0",X"08",X"2A",X"A8",X"0A",X"A0",
		X"00",X"00",X"00",X"08",X"A8",X"28",X"8A",X"A0",X"82",X"80",X"AA",X"A8",X"AA",X"A8",X"80",X"08",
		X"00",X"00",X"00",X"00",X"20",X"A0",X"82",X"A8",X"82",X"08",X"AA",X"08",X"AA",X"28",X"28",X"28",
		X"00",X"00",X"00",X"00",X"A0",X"00",X"80",X"00",X"AA",X"A8",X"AA",X"A8",X"80",X"08",X"A0",X"00",
		X"00",X"00",X"80",X"00",X"AA",X"A8",X"00",X"08",X"00",X"08",X"AA",X"A8",X"AA",X"A8",X"80",X"00",
		X"00",X"00",X"80",X"00",X"A8",X"00",X"0A",X"A0",X"00",X"28",X"0A",X"A8",X"AA",X"80",X"A0",X"00",
		X"00",X"00",X"A0",X"00",X"2A",X"A8",X"00",X"28",X"02",X"A0",X"00",X"28",X"AA",X"A8",X"A0",X"00",
		X"00",X"00",X"80",X"00",X"A0",X"08",X"2A",X"28",X"02",X"80",X"0A",X"A0",X"A8",X"28",X"A0",X"08",
		X"00",X"00",X"80",X"00",X"AA",X"00",X"02",X"A8",X"02",X"A8",X"AA",X"00",X"AA",X"00",X"A0",X"00",
		X"00",X"00",X"A0",X"00",X"A8",X"08",X"8A",X"08",X"82",X"88",X"80",X"A8",X"A0",X"28",X"00",X"08",
		X"00",X"00",X"2A",X"2A",X"08",X"08",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"08",X"08",X"2A",X"2A",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
