library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_PGM_0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_PGM_0 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"DB",X"AF",X"06",X"20",X"09",X"00",X"50",X"5F",X"0B",X"10",X"FC",X"ED",X"56",X"19",X"D9",X"67",
		X"C3",X"C7",X"02",X"3A",X"8E",X"64",X"FE",X"00",X"E0",X"47",X"3E",X"30",X"09",X"35",X"40",X"5F",
		X"2B",X"10",X"FC",X"E1",X"3A",X"8F",X"64",X"FE",X"00",X"E0",X"47",X"3E",X"30",X"09",X"02",X"40",
		X"5F",X"0B",X"10",X"FC",X"E1",X"40",X"00",X"00",X"20",X"F1",X"F5",X"CD",X"FD",X"CD",X"AF",X"1A",
		X"00",X"50",X"2A",X"24",X"64",X"3A",X"26",X"64",X"5F",X"2A",X"27",X"64",X"3A",X"11",X"64",X"5F",
		X"2A",X"14",X"64",X"3A",X"16",X"64",X"5F",X"2A",X"17",X"64",X"3A",X"31",X"64",X"5F",X"2A",X"34",
		X"64",X"3A",X"36",X"64",X"5F",X"2A",X"37",X"64",X"3A",X"09",X"64",X"5F",X"2A",X"0C",X"64",X"3A",
		X"0E",X"64",X"5F",X"2A",X"0F",X"64",X"3A",X"29",X"64",X"5F",X"2A",X"2C",X"64",X"3A",X"2E",X"64",
		X"5F",X"2A",X"2F",X"64",X"3A",X"19",X"64",X"5F",X"2A",X"1C",X"64",X"3A",X"1E",X"64",X"5F",X"2A",
		X"1F",X"64",X"3A",X"39",X"64",X"5F",X"2A",X"3C",X"64",X"3A",X"3E",X"64",X"5F",X"2A",X"3F",X"64",
		X"3A",X"41",X"64",X"5F",X"2A",X"44",X"64",X"3A",X"46",X"64",X"5F",X"2A",X"47",X"64",X"3A",X"61",
		X"64",X"5F",X"2A",X"64",X"64",X"3A",X"66",X"64",X"5F",X"2A",X"67",X"64",X"3A",X"51",X"64",X"5F",
		X"2A",X"54",X"64",X"3A",X"56",X"64",X"5F",X"2A",X"57",X"64",X"3A",X"71",X"64",X"5F",X"09",X"96",
		X"64",X"E3",X"7E",X"28",X"19",X"E3",X"6E",X"08",X"2D",X"06",X"06",X"09",X"4C",X"64",X"11",X"4A",
		X"50",X"3E",X"06",X"26",X"02",X"ED",X"88",X"ED",X"88",X"E5",X"98",X"15",X"10",X"DB",X"06",X"06",
		X"09",X"4E",X"64",X"11",X"DA",X"67",X"3E",X"06",X"26",X"02",X"ED",X"88",X"ED",X"88",X"E5",X"98",
		X"15",X"10",X"DB",X"C3",X"7E",X"01",X"ED",X"73",X"4C",X"64",X"E5",X"60",X"27",X"ED",X"53",X"4A",
		X"50",X"ED",X"73",X"6C",X"64",X"E5",X"60",X"27",X"ED",X"53",X"4C",X"50",X"ED",X"73",X"5C",X"64",
		X"E5",X"60",X"27",X"ED",X"53",X"4E",X"50",X"ED",X"73",X"7C",X"64",X"E5",X"60",X"27",X"ED",X"53",
		X"68",X"50",X"ED",X"73",X"84",X"64",X"E5",X"60",X"27",X"ED",X"53",X"6A",X"50",X"ED",X"73",X"A4",
		X"64",X"E5",X"60",X"27",X"ED",X"53",X"6C",X"50",X"2A",X"4E",X"64",X"E5",X"49",X"27",X"0A",X"DA",
		X"67",X"2A",X"6E",X"64",X"E5",X"49",X"27",X"0A",X"DC",X"67",X"2A",X"5E",X"64",X"E5",X"49",X"27",
		X"0A",X"DE",X"67",X"2A",X"7E",X"64",X"E5",X"49",X"27",X"0A",X"F8",X"67",X"2A",X"86",X"64",X"E5",
		X"49",X"27",X"0A",X"FA",X"67",X"2A",X"A6",X"64",X"E5",X"49",X"27",X"0A",X"FC",X"67",X"2A",X"93",
		X"64",X"0B",X"0A",X"93",X"64",X"7E",X"FE",X"FF",X"08",X"06",X"09",X"8D",X"39",X"0A",X"93",X"64",
		X"09",X"95",X"64",X"E3",X"46",X"08",X"56",X"3A",X"00",X"50",X"E3",X"6F",X"E2",X"2A",X"02",X"E3",
		X"A6",X"E3",X"56",X"08",X"3D",X"3A",X"00",X"50",X"E3",X"7F",X"E2",X"38",X"02",X"3A",X"B0",X"64",
		X"FE",X"06",X"28",X"07",X"3C",X"1A",X"B0",X"64",X"C3",X"3D",X"02",X"AF",X"1A",X"B0",X"64",X"E3",
		X"76",X"08",X"22",X"3A",X"B1",X"64",X"FE",X"00",X"08",X"23",X"C3",X"3D",X"02",X"AF",X"1A",X"07",
		X"50",X"E3",X"B6",X"30",X"68",X"3D",X"1A",X"B1",X"64",X"3E",X"01",X"1A",X"07",X"50",X"E3",X"F6",
		X"30",X"73",X"3A",X"00",X"50",X"E3",X"7F",X"28",X"C4",X"E3",X"96",X"30",X"10",X"3A",X"00",X"50",
		X"E3",X"6F",X"28",X"AD",X"E3",X"86",X"3A",X"B1",X"64",X"3C",X"1A",X"B1",X"64",X"3A",X"B2",X"64",
		X"FE",X"14",X"18",X"32",X"47",X"3A",X"B4",X"64",X"80",X"1A",X"B2",X"64",X"E3",X"3F",X"06",X"00",
		X"80",X"0F",X"1A",X"B5",X"64",X"E5",X"35",X"15",X"E3",X"4E",X"08",X"02",X"E3",X"EE",X"3A",X"05",
		X"65",X"E3",X"C7",X"1A",X"05",X"65",X"E3",X"DE",X"30",X"83",X"E3",X"66",X"08",X"05",X"E3",X"E6",
		X"C3",X"89",X"01",X"E3",X"C6",X"C3",X"B7",X"01",X"E3",X"D6",X"C3",X"AD",X"01",X"00",X"09",X"96",
		X"64",X"E3",X"46",X"28",X"16",X"E5",X"3F",X"16",X"09",X"96",X"64",X"E3",X"7E",X"28",X"04",X"E3",
		X"6E",X"28",X"05",X"E5",X"37",X"16",X"30",X"03",X"E5",X"2F",X"16",X"3A",X"B7",X"64",X"3C",X"1A",
		X"B7",X"64",X"3A",X"B6",X"64",X"3C",X"1A",X"B6",X"64",X"FE",X"3C",X"08",X"23",X"AF",X"1A",X"B6",
		X"64",X"3A",X"88",X"64",X"3C",X"1A",X"88",X"64",X"09",X"95",X"64",X"E3",X"BE",X"3A",X"00",X"50",
		X"E3",X"5F",X"08",X"1D",X"AF",X"1A",X"01",X"50",X"09",X"4A",X"50",X"06",X"24",X"1E",X"00",X"0B",
		X"10",X"FB",X"3E",X"40",X"E5",X"FD",X"14",X"3E",X"21",X"E5",X"25",X"15",X"11",X"D0",X"41",X"09",
		X"92",X"31",X"3E",X"01",X"06",X"04",X"E5",X"D5",X"15",X"06",X"FF",X"09",X"FF",X"FF",X"2B",X"7D",
		X"BC",X"1A",X"C0",X"50",X"08",X"F8",X"10",X"DB",X"5E",X"FB",X"3E",X"01",X"1A",X"00",X"50",X"FD",
		X"C9",X"F5",X"C9",X"F1",X"20",X"ED",X"65",X"3A",X"00",X"50",X"E3",X"4F",X"C2",X"A7",X"05",X"AF",
		X"06",X"20",X"09",X"00",X"50",X"5F",X"0B",X"10",X"FC",X"3E",X"00",X"1A",X"03",X"50",X"19",X"D9",
		X"67",X"E5",X"22",X"16",X"DB",X"20",X"AF",X"20",X"09",X"00",X"40",X"E5",X"16",X"05",X"20",X"E3",
		X"47",X"28",X"02",X"E3",X"D7",X"E3",X"67",X"28",X"02",X"E3",X"F7",X"20",X"09",X"00",X"44",X"E5",
		X"16",X"05",X"20",X"E3",X"47",X"28",X"02",X"E3",X"CF",X"E3",X"67",X"28",X"02",X"E3",X"EF",X"20",
		X"19",X"FD",X"43",X"09",X"00",X"64",X"E5",X"16",X"05",X"20",X"E3",X"47",X"28",X"02",X"E3",X"DF",
		X"E3",X"67",X"28",X"02",X"E3",X"FF",X"20",X"3E",X"01",X"E5",X"25",X"15",X"09",X"00",X"40",X"11",
		X"01",X"40",X"01",X"FE",X"03",X"1E",X"40",X"ED",X"98",X"11",X"4E",X"41",X"09",X"57",X"32",X"3E",
		X"01",X"06",X"23",X"E5",X"D5",X"15",X"11",X"A2",X"40",X"09",X"4A",X"32",X"3E",X"01",X"06",X"30",
		X"E5",X"D5",X"15",X"11",X"EC",X"40",X"09",X"7A",X"32",X"3E",X"01",X"06",X"14",X"E5",X"D5",X"15",
		X"11",X"ED",X"40",X"09",X"A6",X"32",X"3E",X"01",X"06",X"14",X"E5",X"D5",X"15",X"11",X"EE",X"40",
		X"09",X"8A",X"32",X"3E",X"01",X"06",X"14",X"E5",X"D5",X"15",X"11",X"EF",X"40",X"09",X"9E",X"32",
		X"3E",X"01",X"06",X"14",X"E5",X"D5",X"15",X"11",X"93",X"40",X"09",X"46",X"33",X"3E",X"01",X"06",
		X"30",X"E5",X"D5",X"15",X"11",X"DD",X"40",X"09",X"E2",X"32",X"3E",X"01",X"06",X"14",X"E5",X"D5",
		X"15",X"11",X"DE",X"40",X"09",X"F6",X"32",X"3E",X"01",X"06",X"14",X"E5",X"D5",X"15",X"11",X"DF",
		X"40",X"09",X"DA",X"32",X"3E",X"01",X"06",X"14",X"E5",X"D5",X"15",X"11",X"F8",X"40",X"09",X"06",
		X"33",X"3E",X"01",X"06",X"14",X"E5",X"D5",X"15",X"11",X"F9",X"40",X"09",X"32",X"33",X"3E",X"01",
		X"06",X"14",X"E5",X"D5",X"15",X"11",X"FA",X"40",X"09",X"2E",X"33",X"3E",X"01",X"06",X"14",X"E5",
		X"D5",X"15",X"20",X"1A",X"FE",X"64",X"20",X"3A",X"FE",X"64",X"E3",X"57",X"28",X"25",X"11",X"DD",
		X"40",X"09",X"42",X"33",X"3E",X"01",X"06",X"04",X"E5",X"D5",X"15",X"3A",X"FE",X"64",X"E3",X"77",
		X"28",X"25",X"11",X"DE",X"40",X"09",X"42",X"33",X"3E",X"01",X"06",X"04",X"E5",X"D5",X"15",X"3A",
		X"FE",X"64",X"E3",X"4F",X"28",X"25",X"11",X"DF",X"40",X"09",X"42",X"33",X"3E",X"01",X"06",X"04",
		X"E5",X"D5",X"15",X"3A",X"FE",X"64",X"E3",X"6F",X"28",X"25",X"11",X"F8",X"40",X"09",X"42",X"33",
		X"3E",X"01",X"06",X"04",X"E5",X"D5",X"15",X"3A",X"FE",X"64",X"E3",X"5F",X"28",X"25",X"11",X"F9",
		X"40",X"09",X"42",X"33",X"3E",X"01",X"06",X"04",X"E5",X"D5",X"15",X"3A",X"FE",X"64",X"E3",X"7F",
		X"28",X"25",X"11",X"FA",X"40",X"09",X"42",X"33",X"3E",X"01",X"06",X"04",X"E5",X"D5",X"15",X"36",
		X"00",X"09",X"00",X"00",X"E5",X"FD",X"04",X"18",X"02",X"E3",X"C3",X"09",X"00",X"10",X"E5",X"FD",
		X"04",X"18",X"02",X"E3",X"E3",X"09",X"00",X"08",X"E5",X"FD",X"04",X"18",X"02",X"E3",X"D3",X"09",
		X"00",X"18",X"E5",X"FD",X"04",X"18",X"02",X"E3",X"F3",X"3A",X"FE",X"64",X"FE",X"00",X"28",X"02",
		X"3E",X"80",X"9B",X"1A",X"FE",X"64",X"E3",X"47",X"28",X"25",X"11",X"EC",X"40",X"09",X"42",X"33",
		X"3E",X"01",X"06",X"04",X"E5",X"D5",X"15",X"3A",X"FE",X"64",X"E3",X"67",X"28",X"25",X"11",X"ED",
		X"40",X"09",X"42",X"33",X"3E",X"01",X"06",X"04",X"E5",X"D5",X"15",X"3A",X"FE",X"64",X"E3",X"57",
		X"28",X"25",X"11",X"EE",X"40",X"09",X"42",X"33",X"3E",X"01",X"06",X"04",X"E5",X"D5",X"15",X"3A",
		X"FE",X"64",X"E3",X"77",X"28",X"25",X"11",X"EF",X"40",X"09",X"42",X"33",X"3E",X"01",X"06",X"04",
		X"E5",X"D5",X"15",X"3A",X"FE",X"64",X"FE",X"00",X"08",X"26",X"FB",X"3E",X"01",X"1A",X"00",X"50",
		X"3E",X"02",X"E5",X"67",X"15",X"C3",X"F1",X"02",X"1A",X"C0",X"50",X"30",X"FB",X"01",X"00",X"10",
		X"AF",X"1A",X"C0",X"50",X"86",X"0B",X"57",X"23",X"79",X"98",X"7A",X"08",X"DF",X"FE",X"FF",X"28",
		X"02",X"1F",X"E1",X"1F",X"3F",X"E1",X"20",X"CE",X"FC",X"20",X"CD",X"3E",X"11",X"E5",X"1D",X"05",
		X"C9",X"CD",X"3E",X"0A",X"E5",X"1D",X"05",X"C9",X"CD",X"3E",X"44",X"E5",X"1D",X"05",X"C9",X"3E",
		X"A0",X"E5",X"1D",X"05",X"E1",X"1A",X"C0",X"50",X"CD",X"CD",X"D1",X"13",X"01",X"FF",X"03",X"5F",
		X"ED",X"98",X"C9",X"01",X"00",X"04",X"BE",X"C4",X"53",X"05",X"0B",X"77",X"23",X"79",X"98",X"7B",
		X"08",X"DC",X"E1",X"77",X"7E",X"CE",X"27",X"57",X"7B",X"CE",X"27",X"BA",X"28",X"04",X"20",X"E3",
		X"E7",X"20",X"7E",X"CE",X"D8",X"57",X"7B",X"CE",X"D8",X"BA",X"E0",X"20",X"E3",X"C7",X"20",X"7B",
		X"E1",X"65",X"52",X"08",X"54",X"66",X"54",X"2C",X"43",X"67",X"50",X"71",X"52",X"61",X"47",X"60",
		X"54",X"08",X"19",X"39",X"38",X"1B",X"54",X"45",X"64",X"63",X"67",X"08",X"61",X"66",X"43",X"1A",
		X"C0",X"50",X"09",X"00",X"40",X"11",X"01",X"40",X"01",X"FE",X"07",X"1E",X"40",X"ED",X"98",X"1A",
		X"C0",X"50",X"09",X"00",X"64",X"11",X"01",X"64",X"01",X"FE",X"03",X"1E",X"00",X"ED",X"98",X"1A",
		X"C0",X"50",X"09",X"48",X"50",X"11",X"49",X"50",X"01",X"27",X"00",X"1E",X"00",X"ED",X"98",X"1A",
		X"C0",X"50",X"09",X"D8",X"67",X"11",X"D9",X"67",X"01",X"27",X"00",X"1E",X"00",X"ED",X"98",X"1A",
		X"C0",X"50",X"09",X"40",X"50",X"11",X"41",X"50",X"01",X"37",X"00",X"1E",X"00",X"ED",X"98",X"09",
		X"24",X"64",X"11",X"25",X"64",X"01",X"67",X"00",X"1E",X"FF",X"ED",X"98",X"09",X"8D",X"39",X"0A",
		X"93",X"64",X"3A",X"80",X"50",X"47",X"CE",X"03",X"1A",X"B3",X"64",X"09",X"B4",X"33",X"E5",X"98",
		X"15",X"7E",X"1A",X"B4",X"64",X"78",X"CE",X"24",X"E3",X"3F",X"E3",X"3F",X"09",X"89",X"39",X"E5",
		X"98",X"15",X"7E",X"1A",X"8A",X"64",X"78",X"CE",X"18",X"09",X"49",X"39",X"E5",X"98",X"15",X"0A",
		X"8B",X"64",X"78",X"CE",X"18",X"E3",X"3F",X"E3",X"3F",X"E3",X"3F",X"E3",X"3F",X"1A",X"8D",X"64",
		X"78",X"E3",X"5F",X"08",X"05",X"09",X"96",X"64",X"E3",X"FE",X"FB",X"3E",X"01",X"1A",X"00",X"50",
		X"E5",X"04",X"1C",X"09",X"C2",X"43",X"11",X"C3",X"43",X"01",X"3C",X"00",X"1E",X"40",X"ED",X"98",
		X"09",X"C2",X"47",X"11",X"C3",X"47",X"01",X"34",X"00",X"1E",X"05",X"ED",X"98",X"1A",X"C0",X"50",
		X"09",X"CA",X"47",X"11",X"CB",X"47",X"01",X"34",X"00",X"1E",X"21",X"ED",X"98",X"1A",X"C0",X"50",
		X"09",X"A3",X"30",X"11",X"C3",X"43",X"01",X"32",X"00",X"ED",X"98",X"AF",X"1A",X"CC",X"43",X"1A",
		X"ED",X"43",X"1A",X"DE",X"43",X"09",X"BA",X"39",X"11",X"9B",X"64",X"01",X"3C",X"00",X"ED",X"98",
		X"09",X"B8",X"64",X"11",X"DA",X"43",X"E5",X"0E",X"10",X"09",X"02",X"40",X"11",X"03",X"40",X"01",
		X"3C",X"00",X"1E",X"40",X"ED",X"98",X"1A",X"C0",X"50",X"09",X"02",X"44",X"11",X"03",X"44",X"01",
		X"34",X"00",X"1E",X"21",X"ED",X"98",X"09",X"0A",X"44",X"11",X"0B",X"44",X"01",X"34",X"00",X"1E",
		X"11",X"ED",X"98",X"1A",X"C0",X"50",X"09",X"8D",X"30",X"11",X"27",X"40",X"01",X"06",X"00",X"ED",
		X"98",X"AF",X"1A",X"24",X"40",X"3A",X"B3",X"64",X"FE",X"00",X"08",X"23",X"09",X"AB",X"30",X"11",
		X"24",X"40",X"01",X"21",X"00",X"ED",X"98",X"1A",X"C0",X"50",X"09",X"05",X"65",X"11",X"06",X"65",
		X"01",X"FF",X"00",X"1E",X"00",X"ED",X"98",X"09",X"5C",X"1D",X"0A",X"36",X"65",X"0A",X"06",X"65",
		X"09",X"35",X"65",X"0A",X"25",X"65",X"09",X"8A",X"1D",X"0A",X"39",X"65",X"0A",X"09",X"65",X"09",
		X"38",X"65",X"0A",X"28",X"65",X"09",X"B9",X"1D",X"0A",X"54",X"65",X"0A",X"3C",X"65",X"09",X"53",
		X"65",X"0A",X"43",X"65",X"09",X"EB",X"1D",X"0A",X"6F",X"65",X"0A",X"57",X"65",X"09",X"6E",X"65",
		X"0A",X"76",X"65",X"09",X"B0",X"1E",X"0A",X"A2",X"65",X"0A",X"5A",X"65",X"09",X"A1",X"65",X"0A",
		X"79",X"65",X"09",X"E2",X"1E",X"0A",X"8D",X"65",X"0A",X"A5",X"65",X"09",X"8C",X"65",X"0A",X"94",
		X"65",X"09",X"04",X"38",X"0A",X"C0",X"65",X"0A",X"A8",X"65",X"09",X"BF",X"65",X"0A",X"AF",X"65",
		X"09",X"31",X"38",X"0A",X"F3",X"65",X"0A",X"C3",X"65",X"09",X"F2",X"65",X"0A",X"E2",X"65",X"06",
		X"08",X"09",X"40",X"50",X"1E",X"00",X"0B",X"10",X"FB",X"3E",X"00",X"1A",X"03",X"50",X"09",X"96",
		X"64",X"E3",X"EE",X"3A",X"B3",X"64",X"FE",X"00",X"E2",X"39",X"21",X"3A",X"B2",X"64",X"FE",X"00",
		X"C2",X"39",X"21",X"09",X"95",X"64",X"E3",X"8E",X"AF",X"1A",X"01",X"50",X"09",X"96",X"64",X"E3",
		X"86",X"E5",X"22",X"16",X"1A",X"C0",X"50",X"E5",X"D1",X"19",X"3E",X"01",X"E5",X"67",X"15",X"09",
		X"95",X"64",X"E3",X"6E",X"C2",X"39",X"21",X"E5",X"7C",X"10",X"3E",X"07",X"E5",X"67",X"15",X"09",
		X"95",X"64",X"E3",X"6E",X"C2",X"39",X"21",X"3E",X"40",X"E5",X"FD",X"14",X"11",X"44",X"44",X"09",
		X"DE",X"39",X"3E",X"01",X"06",X"34",X"E5",X"EB",X"15",X"11",X"61",X"44",X"09",X"F8",X"39",X"3E",
		X"03",X"06",X"34",X"E5",X"EB",X"15",X"11",X"50",X"44",X"09",X"DF",X"39",X"3E",X"03",X"06",X"34",
		X"E5",X"EB",X"15",X"11",X"70",X"44",X"09",X"F8",X"39",X"3E",X"03",X"06",X"34",X"E5",X"EB",X"15",
		X"11",X"73",X"44",X"09",X"F9",X"39",X"3E",X"03",X"06",X"34",X"E5",X"EB",X"15",X"11",X"C4",X"40",
		X"09",X"96",X"31",X"3E",X"01",X"06",X"14",X"E5",X"D5",X"15",X"11",X"E1",X"40",X"09",X"AB",X"31",
		X"3E",X"01",X"06",X"14",X"E5",X"D5",X"15",X"11",X"A3",X"40",X"09",X"BF",X"31",X"3E",X"01",X"06",
		X"30",X"E5",X"D5",X"15",X"11",X"98",X"40",X"09",X"D7",X"31",X"3E",X"01",X"06",X"16",X"E5",X"D5",
		X"15",X"11",X"52",X"41",X"09",X"ED",X"31",X"3E",X"01",X"06",X"24",X"E5",X"D5",X"15",X"3A",X"B3",
		X"64",X"FE",X"01",X"08",X"27",X"11",X"31",X"41",X"09",X"F9",X"31",X"3E",X"01",X"06",X"27",X"E5",
		X"D5",X"15",X"30",X"08",X"FE",X"02",X"08",X"27",X"11",X"31",X"41",X"09",X"20",X"32",X"3E",X"01",
		X"06",X"27",X"E5",X"D5",X"15",X"30",X"25",X"11",X"31",X"41",X"09",X"17",X"32",X"3E",X"01",X"06",
		X"27",X"E5",X"D5",X"15",X"11",X"B4",X"40",X"09",X"0E",X"32",X"3E",X"01",X"06",X"31",X"E5",X"D5",
		X"15",X"3A",X"8D",X"64",X"FE",X"00",X"08",X"27",X"11",X"7C",X"41",X"09",X"3F",X"32",X"3E",X"01",
		X"06",X"06",X"E5",X"D5",X"15",X"30",X"1B",X"FE",X"01",X"08",X"27",X"11",X"7C",X"41",X"09",X"45",
		X"32",X"3E",X"01",X"06",X"06",X"E5",X"D5",X"15",X"30",X"08",X"FE",X"02",X"08",X"27",X"11",X"7C",
		X"41",X"09",X"63",X"32",X"3E",X"01",X"06",X"06",X"E5",X"D5",X"15",X"30",X"25",X"11",X"7C",X"41",
		X"09",X"51",X"32",X"3E",X"01",X"06",X"06",X"E5",X"D5",X"15",X"3E",X"04",X"E5",X"67",X"15",X"09",
		X"95",X"64",X"E3",X"6E",X"08",X"53",X"E5",X"05",X"1C",X"AF",X"1A",X"FF",X"64",X"1A",X"01",X"65",
		X"1A",X"03",X"65",X"1A",X"00",X"65",X"1A",X"02",X"65",X"1A",X"04",X"65",X"E5",X"07",X"1C",X"E5",
		X"FA",X"26",X"E5",X"14",X"1C",X"E5",X"BC",X"33",X"AF",X"1A",X"08",X"65",X"1A",X"3B",X"65",X"1A",
		X"56",X"65",X"1A",X"59",X"65",X"1A",X"A4",X"65",X"1A",X"8F",X"65",X"1A",X"C2",X"65",X"E5",X"15",
		X"16",X"1A",X"C0",X"50",X"09",X"95",X"64",X"E3",X"6E",X"08",X"26",X"09",X"96",X"64",X"E3",X"66",
		X"08",X"02",X"30",X"E6",X"E3",X"A6",X"C3",X"89",X"07",X"E5",X"22",X"16",X"09",X"95",X"64",X"E3",
		X"CE",X"E3",X"AE",X"09",X"96",X"64",X"E3",X"A6",X"E3",X"96",X"E3",X"B6",X"09",X"97",X"64",X"E3",
		X"96",X"09",X"96",X"64",X"E3",X"C6",X"09",X"24",X"64",X"11",X"25",X"64",X"01",X"67",X"00",X"1E",
		X"FF",X"ED",X"98",X"3E",X"FF",X"1A",X"01",X"50",X"09",X"97",X"64",X"E3",X"56",X"08",X"27",X"3A",
		X"FD",X"64",X"3C",X"1A",X"FD",X"64",X"FE",X"14",X"08",X"04",X"E3",X"D6",X"E3",X"F6",X"00",X"1A",
		X"C0",X"50",X"3E",X"40",X"E5",X"FD",X"14",X"3E",X"03",X"E5",X"25",X"15",X"3A",X"B3",X"64",X"FE",
		X"00",X"E2",X"14",X"22",X"3A",X"B2",X"64",X"FE",X"02",X"18",X"64",X"11",X"58",X"41",X"09",X"9C",
		X"30",X"3E",X"01",X"06",X"23",X"E5",X"D5",X"15",X"3A",X"40",X"50",X"E3",X"6F",X"08",X"5C",X"3A",
		X"B3",X"64",X"FE",X"00",X"28",X"15",X"3A",X"B2",X"64",X"FE",X"02",X"38",X"4E",X"D6",X"02",X"1A",
		X"B2",X"64",X"3A",X"B5",X"64",X"D6",X"01",X"0F",X"1A",X"B5",X"64",X"09",X"96",X"64",X"E3",X"CE",
		X"3A",X"8A",X"64",X"1A",X"8E",X"64",X"E5",X"13",X"00",X"3A",X"B3",X"64",X"FE",X"00",X"E2",X"6F",
		X"22",X"E5",X"35",X"15",X"C3",X"6F",X"22",X"FE",X"04",X"18",X"29",X"11",X"26",X"41",X"09",X"BF",
		X"30",X"3E",X"01",X"06",X"11",X"E5",X"D5",X"15",X"11",X"10",X"42",X"09",X"D0",X"30",X"3E",X"01",
		X"06",X"02",X"E5",X"D5",X"15",X"11",X"5A",X"41",X"09",X"9C",X"30",X"3E",X"01",X"06",X"23",X"E5",
		X"D5",X"15",X"30",X"94",X"11",X"90",X"40",X"09",X"D2",X"30",X"3E",X"01",X"06",X"31",X"E5",X"D5",
		X"15",X"30",X"85",X"3A",X"40",X"50",X"E3",X"5F",X"08",X"1B",X"3A",X"B3",X"64",X"FE",X"00",X"28",
		X"15",X"3A",X"B2",X"64",X"FE",X"04",X"38",X"0D",X"D6",X"04",X"1A",X"B2",X"64",X"3A",X"B5",X"64",
		X"D6",X"02",X"0F",X"1A",X"B5",X"64",X"09",X"96",X"64",X"E3",X"8E",X"3A",X"8A",X"64",X"1A",X"8E",
		X"64",X"1A",X"8F",X"64",X"E5",X"13",X"00",X"E5",X"0C",X"00",X"C3",X"F1",X"21",X"1A",X"C0",X"50",
		X"09",X"95",X"64",X"E3",X"5E",X"08",X"03",X"C3",X"A8",X"21",X"E3",X"9E",X"C3",X"7F",X"21",X"AF",
		X"09",X"A8",X"64",X"11",X"A9",X"64",X"01",X"05",X"00",X"5F",X"ED",X"98",X"1A",X"99",X"64",X"1A",
		X"9A",X"64",X"3E",X"40",X"09",X"CC",X"43",X"11",X"CD",X"43",X"01",X"05",X"00",X"5F",X"ED",X"98",
		X"09",X"DE",X"43",X"11",X"DF",X"43",X"01",X"05",X"00",X"5F",X"ED",X"98",X"AF",X"1A",X"CC",X"43",
		X"1A",X"DE",X"43",X"AF",X"1A",X"FF",X"64",X"1A",X"01",X"65",X"1A",X"03",X"65",X"1A",X"00",X"65",
		X"1A",X"02",X"65",X"1A",X"04",X"65",X"E5",X"06",X"1C",X"E5",X"13",X"1C",X"09",X"97",X"64",X"E3",
		X"E6",X"09",X"96",X"64",X"E3",X"4E",X"28",X"02",X"30",X"32",X"3E",X"00",X"1A",X"03",X"50",X"E5",
		X"44",X"15",X"11",X"50",X"41",X"09",X"EB",X"30",X"3E",X"01",X"06",X"25",X"E5",X"D5",X"15",X"3E",
		X"03",X"E5",X"67",X"15",X"09",X"96",X"64",X"E3",X"EE",X"3A",X"8E",X"64",X"3D",X"1A",X"8E",X"64",
		X"3E",X"40",X"09",X"16",X"40",X"11",X"17",X"40",X"01",X"20",X"00",X"5F",X"ED",X"98",X"E5",X"13",
		X"00",X"3A",X"FF",X"64",X"1A",X"03",X"65",X"3A",X"00",X"65",X"1A",X"04",X"65",X"E5",X"6B",X"1C",
		X"C3",X"B3",X"23",X"09",X"96",X"64",X"E3",X"4E",X"08",X"E2",X"E3",X"6E",X"28",X"AC",X"3A",X"96",
		X"64",X"E3",X"7F",X"08",X"43",X"E5",X"44",X"15",X"11",X"50",X"41",X"09",X"F8",X"30",X"3E",X"01",
		X"06",X"25",X"E5",X"D5",X"15",X"3E",X"03",X"E5",X"67",X"15",X"09",X"96",X"64",X"E3",X"AE",X"3A",
		X"8F",X"64",X"3D",X"1A",X"8F",X"64",X"3E",X"40",X"09",X"02",X"40",X"11",X"03",X"40",X"01",X"20",
		X"00",X"5F",X"ED",X"98",X"E5",X"0C",X"00",X"3A",X"01",X"65",X"1A",X"03",X"65",X"3A",X"02",X"65",
		X"1A",X"04",X"65",X"E5",X"6D",X"1C",X"30",X"1B",X"3E",X"01",X"1A",X"03",X"50",X"30",X"9E",X"E5",
		X"44",X"15",X"09",X"96",X"64",X"E3",X"4E",X"C2",X"E9",X"22",X"11",X"10",X"41",X"09",X"05",X"31",
		X"3E",X"01",X"06",X"11",X"E5",X"D5",X"15",X"09",X"08",X"65",X"E3",X"C6",X"3E",X"01",X"E5",X"67",
		X"15",X"09",X"96",X"64",X"E3",X"6E",X"28",X"8F",X"C3",X"E9",X"22",X"E5",X"FA",X"26",X"09",X"97",
		X"64",X"E3",X"66",X"28",X"13",X"E3",X"A6",X"09",X"C2",X"65",X"E3",X"C6",X"1A",X"C0",X"50",X"3A",
		X"C2",X"65",X"FE",X"00",X"08",X"DE",X"30",X"05",X"3E",X"02",X"E5",X"67",X"15",X"09",X"8F",X"65",
		X"E3",X"C6",X"09",X"59",X"65",X"E3",X"C6",X"E5",X"BC",X"33",X"ED",X"73",X"AE",X"64",X"7B",X"9A",
		X"28",X"21",X"09",X"00",X"00",X"0A",X"AE",X"64",X"E5",X"4E",X"27",X"1A",X"C0",X"50",X"E5",X"15",
		X"16",X"09",X"96",X"64",X"E3",X"66",X"28",X"F7",X"E3",X"A6",X"E5",X"22",X"16",X"09",X"96",X"64",
		X"E3",X"56",X"08",X"27",X"E5",X"59",X"1C",X"E5",X"22",X"16",X"09",X"96",X"64",X"E3",X"76",X"08",
		X"21",X"30",X"4F",X"E3",X"96",X"E5",X"58",X"1C",X"30",X"EA",X"E3",X"B6",X"09",X"97",X"64",X"E3",
		X"E6",X"09",X"96",X"64",X"E3",X"6E",X"08",X"29",X"3A",X"01",X"65",X"3C",X"FE",X"24",X"08",X"02",
		X"3E",X"23",X"1A",X"01",X"65",X"1A",X"03",X"65",X"3A",X"02",X"65",X"3C",X"FE",X"31",X"08",X"02",
		X"3E",X"30",X"1A",X"02",X"65",X"1A",X"04",X"65",X"E5",X"5A",X"1C",X"E5",X"6F",X"1C",X"C3",X"B3",
		X"23",X"3A",X"FF",X"64",X"3C",X"FE",X"24",X"08",X"02",X"3E",X"23",X"1A",X"FF",X"64",X"1A",X"03",
		X"65",X"3A",X"00",X"65",X"3C",X"FE",X"31",X"08",X"02",X"3E",X"30",X"1A",X"00",X"65",X"1A",X"04",
		X"65",X"E5",X"5A",X"1C",X"E5",X"6E",X"1C",X"C3",X"B3",X"23",X"3A",X"98",X"64",X"FE",X"00",X"08",
		X"2E",X"09",X"96",X"64",X"E3",X"6E",X"08",X"2F",X"3A",X"8F",X"64",X"FE",X"00",X"08",X"66",X"E5",
		X"44",X"15",X"11",X"90",X"41",X"09",X"16",X"31",X"3E",X"01",X"06",X"21",X"E5",X"D5",X"15",X"3E",
		X"02",X"E5",X"67",X"15",X"E5",X"EE",X"11",X"09",X"95",X"64",X"E3",X"DE",X"C3",X"79",X"07",X"D6",
		X"01",X"1A",X"98",X"64",X"C3",X"6F",X"23",X"3A",X"8E",X"64",X"FE",X"00",X"08",X"0D",X"09",X"96",
		X"64",X"E3",X"4E",X"08",X"E2",X"E5",X"44",X"15",X"11",X"D8",X"40",X"09",X"37",X"31",X"3E",X"01",
		X"06",X"14",X"E5",X"D5",X"15",X"3E",X"03",X"E5",X"67",X"15",X"C3",X"36",X"23",X"E5",X"6C",X"1C",
		X"C3",X"13",X"23",X"E5",X"6A",X"1C",X"C3",X"13",X"23",X"2A",X"91",X"64",X"EB",X"F5",X"09",X"00",
		X"00",X"F5",X"31",X"F5",X"7E",X"01",X"F5",X"86",X"02",X"47",X"CE",X"27",X"F5",X"5F",X"02",X"E3",
		X"38",X"E3",X"38",X"E3",X"38",X"E3",X"38",X"F5",X"7E",X"00",X"09",X"07",X"25",X"E3",X"0F",X"E5",
		X"98",X"15",X"76",X"0B",X"56",X"EB",X"E9",X"13",X"25",X"13",X"25",X"14",X"25",X"34",X"25",X"0C",
		X"25",X"2C",X"25",X"E1",X"F5",X"7E",X"04",X"90",X"F5",X"5F",X"04",X"E1",X"F5",X"7E",X"04",X"80",
		X"F5",X"5F",X"04",X"E1",X"F5",X"7E",X"03",X"80",X"F5",X"5F",X"03",X"E1",X"F5",X"7E",X"03",X"90",
		X"F5",X"5F",X"03",X"E1",X"2A",X"76",X"64",X"EB",X"F5",X"09",X"00",X"00",X"F5",X"31",X"EB",X"01",
		X"00",X"64",X"1F",X"3F",X"ED",X"42",X"CD",X"F5",X"7E",X"00",X"09",X"57",X"25",X"E3",X"0F",X"E5",
		X"98",X"15",X"76",X"0B",X"56",X"EB",X"E9",X"0F",X"26",X"4B",X"25",X"8E",X"25",X"1E",X"26",X"40",
		X"26",X"53",X"26",X"F5",X"7E",X"03",X"1A",X"74",X"64",X"F5",X"7E",X"04",X"1A",X"75",X"64",X"E5",
		X"BD",X"26",X"F5",X"7E",X"06",X"12",X"3A",X"22",X"64",X"FE",X"00",X"08",X"17",X"3A",X"23",X"64",
		X"FE",X"00",X"08",X"17",X"C1",X"09",X"24",X"64",X"21",X"CD",X"D1",X"13",X"01",X"05",X"00",X"1E",
		X"FF",X"ED",X"98",X"E1",X"F5",X"7E",X"06",X"13",X"12",X"30",X"E9",X"F5",X"7E",X"06",X"09",X"08",
		X"00",X"31",X"EB",X"12",X"30",X"F6",X"E5",X"CD",X"26",X"F5",X"7E",X"03",X"90",X"1A",X"74",X"64",
		X"F5",X"7E",X"04",X"1A",X"75",X"64",X"E5",X"BD",X"26",X"3A",X"22",X"64",X"FE",X"00",X"28",X"1A",
		X"3A",X"22",X"64",X"E3",X"0F",X"F5",X"46",X"05",X"80",X"3D",X"C1",X"FD",X"09",X"24",X"64",X"FD",
		X"21",X"FD",X"5B",X"00",X"FD",X"5A",X"01",X"FD",X"5F",X"02",X"3C",X"13",X"FD",X"5B",X"03",X"FD",
		X"5A",X"04",X"FD",X"5F",X"05",X"3A",X"74",X"64",X"F5",X"5F",X"03",X"3A",X"75",X"64",X"F5",X"5F",
		X"04",X"E1",X"3A",X"23",X"64",X"FE",X"00",X"E2",X"74",X"26",X"3A",X"23",X"64",X"E3",X"0F",X"C6",
		X"27",X"F5",X"46",X"05",X"80",X"C1",X"FD",X"09",X"24",X"64",X"FD",X"21",X"FD",X"5B",X"00",X"FD",
		X"5A",X"01",X"FD",X"5F",X"02",X"3C",X"09",X"08",X"00",X"31",X"EB",X"FD",X"5B",X"03",X"FD",X"5A",
		X"04",X"FD",X"5F",X"05",X"C3",X"CD",X"25",X"F5",X"7E",X"03",X"1A",X"74",X"64",X"F5",X"7E",X"04",
		X"1A",X"75",X"64",X"C3",X"9E",X"25",X"E5",X"CD",X"26",X"F5",X"7E",X"03",X"80",X"C3",X"AD",X"25",
		X"E5",X"CD",X"26",X"F5",X"7E",X"04",X"90",X"1A",X"75",X"64",X"F5",X"7E",X"03",X"1A",X"74",X"64",
		X"C3",X"9E",X"25",X"E5",X"CD",X"26",X"F5",X"7E",X"04",X"80",X"30",X"EB",X"F5",X"7E",X"05",X"C1",
		X"FD",X"09",X"24",X"64",X"FD",X"21",X"FD",X"5B",X"00",X"FD",X"5A",X"01",X"FD",X"5F",X"02",X"3A",
		X"74",X"64",X"F5",X"5F",X"03",X"3A",X"75",X"64",X"F5",X"5F",X"04",X"F5",X"7E",X"00",X"09",X"90",
		X"26",X"E3",X"0F",X"E5",X"98",X"15",X"D5",X"76",X"0B",X"56",X"EB",X"D1",X"F5",X"7E",X"06",X"E9",
		X"B4",X"26",X"B4",X"26",X"B5",X"26",X"A8",X"26",X"AB",X"26",X"9A",X"26",X"E1",X"13",X"FD",X"5B",
		X"03",X"FD",X"5A",X"04",X"FD",X"5F",X"05",X"E1",X"33",X"30",X"DB",X"09",X"08",X"00",X"31",X"EB",
		X"30",X"EC",X"EB",X"11",X"08",X"00",X"1F",X"3F",X"ED",X"52",X"EB",X"30",X"C9",X"3A",X"74",X"64",
		X"CE",X"07",X"1A",X"22",X"64",X"3A",X"75",X"64",X"CE",X"07",X"1A",X"23",X"64",X"3A",X"74",X"64",
		X"E3",X"3F",X"E3",X"3F",X"E3",X"3F",X"57",X"3A",X"75",X"64",X"E3",X"3F",X"E3",X"3F",X"E3",X"3F",
		X"77",X"E5",X"F7",X"14",X"E1",X"F5",X"7E",X"01",X"F5",X"86",X"02",X"47",X"CE",X"27",X"F5",X"5F",
		X"02",X"E3",X"38",X"E3",X"38",X"E3",X"38",X"E3",X"38",X"E1",X"3A",X"03",X"65",X"09",X"20",X"27",
		X"E3",X"0F",X"E3",X"0F",X"E5",X"98",X"15",X"E9",X"E5",X"2B",X"28",X"E1",X"E5",X"4D",X"28",X"E1",
		X"E5",X"B7",X"28",X"E1",X"E5",X"F1",X"28",X"E1",X"E5",X"13",X"29",X"E1",X"E5",X"65",X"29",X"E1",
		X"E5",X"87",X"29",X"E1",X"E5",X"C1",X"29",X"E1",X"E5",X"FB",X"29",X"E1",X"E5",X"1D",X"2A",X"E1",
		X"E5",X"6F",X"2A",X"E1",X"E5",X"A9",X"2A",X"E1",X"E5",X"CB",X"2A",X"E1",X"E5",X"CC",X"2A",X"E1",
		X"E5",X"CD",X"2A",X"E1",X"E5",X"CE",X"2A",X"E1",X"D5",X"1F",X"3F",X"09",X"26",X"01",X"16",X"00",
		X"ED",X"52",X"7D",X"1F",X"3F",X"09",X"10",X"01",X"D1",X"72",X"16",X"00",X"ED",X"52",X"55",X"77",
		X"E1",X"7D",X"EE",X"03",X"6F",X"E1",X"09",X"96",X"64",X"E3",X"46",X"E0",X"E3",X"6E",X"28",X"43",
		X"09",X"A8",X"64",X"7B",X"86",X"0F",X"5F",X"0B",X"7A",X"A6",X"0F",X"5F",X"0B",X"3E",X"00",X"A6",
		X"0F",X"5F",X"38",X"02",X"30",X"1A",X"09",X"96",X"64",X"E3",X"6E",X"28",X"13",X"09",X"DE",X"43",
		X"11",X"DF",X"43",X"01",X"05",X"00",X"1E",X"40",X"ED",X"98",X"AF",X"1A",X"DE",X"43",X"30",X"30",
		X"09",X"CC",X"43",X"11",X"CD",X"43",X"01",X"05",X"00",X"1E",X"40",X"ED",X"98",X"AF",X"1A",X"CC",
		X"43",X"30",X"05",X"09",X"AB",X"64",X"30",X"BB",X"09",X"96",X"64",X"E3",X"6E",X"28",X"74",X"09",
		X"AA",X"64",X"11",X"FB",X"43",X"3A",X"99",X"64",X"DD",X"E5",X"0E",X"10",X"0B",X"0B",X"0B",X"EB",
		X"2A",X"8B",X"64",X"D9",X"FE",X"04",X"D0",X"E3",X"0F",X"E3",X"0F",X"3C",X"3C",X"E5",X"98",X"15",
		X"E5",X"AA",X"11",X"D0",X"3A",X"98",X"64",X"3C",X"1A",X"98",X"64",X"09",X"08",X"65",X"E3",X"C6",
		X"09",X"96",X"64",X"E3",X"6E",X"28",X"12",X"3A",X"99",X"64",X"3C",X"1A",X"99",X"64",X"3A",X"8E",
		X"64",X"3C",X"1A",X"8E",X"64",X"E5",X"13",X"00",X"E1",X"3A",X"9A",X"64",X"3C",X"1A",X"9A",X"64",
		X"3A",X"8F",X"64",X"3C",X"1A",X"8F",X"64",X"E5",X"0C",X"00",X"E1",X"09",X"AD",X"64",X"11",X"E9",
		X"43",X"3A",X"9A",X"64",X"30",X"8A",X"3E",X"03",X"DD",X"7E",X"CE",X"D8",X"E3",X"3F",X"E3",X"3F",
		X"E3",X"3F",X"E3",X"3F",X"47",X"3A",X"96",X"64",X"E3",X"5F",X"28",X"0A",X"78",X"12",X"33",X"7E",
		X"CE",X"27",X"47",X"3A",X"96",X"64",X"E3",X"5F",X"1A",X"96",X"64",X"28",X"08",X"78",X"12",X"2B",
		X"33",X"D9",X"3D",X"08",X"D3",X"3A",X"96",X"64",X"E3",X"9F",X"1A",X"96",X"64",X"E1",X"78",X"FE",
		X"00",X"28",X"F3",X"3A",X"96",X"64",X"E3",X"DF",X"1A",X"96",X"64",X"30",X"E7",X"78",X"FE",X"00",
		X"28",X"F5",X"3A",X"96",X"64",X"E3",X"DF",X"1A",X"96",X"64",X"30",X"D1",X"09",X"97",X"64",X"E3",
		X"76",X"28",X"2C",X"E3",X"B6",X"09",X"40",X"40",X"E5",X"89",X"10",X"FE",X"3A",X"08",X"24",X"09",
		X"40",X"44",X"E5",X"89",X"10",X"FE",X"B4",X"08",X"02",X"30",X"14",X"AF",X"1A",X"B3",X"64",X"30",
		X"26",X"AF",X"11",X"80",X"03",X"86",X"0B",X"33",X"47",X"7A",X"9B",X"78",X"08",X"DF",X"E1",X"00",
		X"3E",X"40",X"E5",X"FD",X"14",X"3E",X"21",X"E5",X"25",X"15",X"11",X"29",X"45",X"09",X"EE",X"10",
		X"3E",X"15",X"06",X"23",X"E5",X"EB",X"15",X"11",X"45",X"41",X"09",X"1B",X"31",X"3E",X"01",X"06",
		X"24",X"E5",X"D5",X"15",X"09",X"77",X"33",X"11",X"E2",X"42",X"01",X"FF",X"21",X"ED",X"88",X"13",
		X"10",X"FB",X"AF",X"12",X"E5",X"02",X"16",X"3E",X"01",X"12",X"E5",X"EF",X"10",X"E1",X"03",X"09",
		X"9B",X"64",X"11",X"6A",X"42",X"E5",X"2F",X"11",X"11",X"6C",X"42",X"E5",X"2F",X"11",X"11",X"6E",
		X"42",X"E5",X"2F",X"11",X"11",X"58",X"42",X"E5",X"2F",X"11",X"11",X"5A",X"42",X"E5",X"2F",X"11",
		X"11",X"5C",X"42",X"E5",X"2F",X"11",X"11",X"5E",X"42",X"E5",X"2F",X"11",X"11",X"78",X"42",X"E5",
		X"2F",X"11",X"11",X"7A",X"42",X"E5",X"2F",X"11",X"11",X"7C",X"42",X"E5",X"2F",X"11",X"E1",X"06",
		X"03",X"26",X"27",X"3E",X"09",X"ED",X"88",X"E5",X"E1",X"15",X"10",X"DF",X"0B",X"0B",X"3E",X"40",
		X"E5",X"E1",X"15",X"E5",X"64",X"11",X"3E",X"04",X"E5",X"98",X"15",X"E1",X"3E",X"03",X"DD",X"7E",
		X"CE",X"D8",X"E3",X"3F",X"E3",X"3F",X"E3",X"3F",X"E3",X"3F",X"47",X"3A",X"96",X"64",X"E3",X"5F",
		X"28",X"2A",X"78",X"12",X"3E",X"08",X"E5",X"E1",X"15",X"7E",X"CE",X"27",X"47",X"3A",X"96",X"64",
		X"E3",X"5F",X"1A",X"96",X"64",X"28",X"0C",X"78",X"12",X"2B",X"3E",X"08",X"E5",X"E1",X"15",X"D9",
		X"3D",X"08",X"E3",X"3A",X"96",X"64",X"E3",X"9F",X"1A",X"96",X"64",X"E1",X"78",X"FE",X"00",X"28",
		X"D3",X"3A",X"96",X"64",X"E3",X"DF",X"1A",X"96",X"64",X"30",X"C7",X"78",X"FE",X"00",X"28",X"F1",
		X"3A",X"96",X"64",X"E3",X"DF",X"1A",X"96",X"64",X"30",X"E5",X"06",X"03",X"32",X"BE",X"38",X"20",
		X"08",X"26",X"2B",X"33",X"10",X"DE",X"30",X"06",X"E5",X"C5",X"11",X"1F",X"3F",X"E1",X"1F",X"E1",
		X"E5",X"C5",X"11",X"1F",X"E1",X"78",X"FE",X"00",X"E0",X"2B",X"33",X"3D",X"08",X"FB",X"E1",X"63",
		X"65",X"52",X"08",X"54",X"66",X"54",X"2C",X"43",X"67",X"50",X"71",X"52",X"61",X"47",X"60",X"54",
		X"08",X"19",X"39",X"38",X"1B",X"54",X"45",X"64",X"63",X"67",X"08",X"61",X"66",X"43",X"09",X"96",
		X"64",X"E3",X"EE",X"09",X"A8",X"64",X"11",X"DD",X"64",X"01",X"03",X"00",X"ED",X"98",X"E5",X"30",
		X"12",X"09",X"96",X"64",X"E3",X"4E",X"C0",X"E3",X"AE",X"09",X"AB",X"64",X"11",X"DD",X"64",X"01",
		X"03",X"00",X"ED",X"98",X"E5",X"30",X"12",X"E1",X"01",X"00",X"22",X"09",X"D9",X"64",X"11",X"DF",
		X"64",X"2B",X"2B",X"2B",X"C5",X"E5",X"AA",X"11",X"C1",X"18",X"22",X"3E",X"06",X"81",X"67",X"10",
		X"ED",X"2B",X"2B",X"30",X"20",X"79",X"FE",X"00",X"E0",X"0B",X"0B",X"0B",X"0B",X"C5",X"CD",X"06",
		X"00",X"09",X"EE",X"64",X"11",X"DC",X"64",X"ED",X"B8",X"3E",X"40",X"E5",X"FD",X"14",X"09",X"96",
		X"64",X"E3",X"6E",X"08",X"33",X"11",X"4A",X"41",X"09",X"FB",X"30",X"3E",X"01",X"06",X"22",X"E5",
		X"D5",X"15",X"09",X"96",X"64",X"E3",X"7E",X"28",X"31",X"3E",X"01",X"1A",X"03",X"50",X"30",X"12",
		X"11",X"4A",X"41",X"09",X"EE",X"30",X"3E",X"01",X"06",X"22",X"E5",X"D5",X"15",X"3E",X"00",X"1A",
		X"03",X"50",X"11",X"40",X"44",X"09",X"F3",X"14",X"3E",X"23",X"06",X"34",X"E5",X"EB",X"15",X"11",
		X"64",X"44",X"09",X"F4",X"14",X"3E",X"03",X"06",X"34",X"E5",X"EB",X"15",X"11",X"51",X"44",X"09",
		X"F5",X"14",X"3E",X"10",X"06",X"34",X"E5",X"EB",X"15",X"11",X"50",X"44",X"09",X"F6",X"14",X"3E",
		X"02",X"06",X"34",X"E5",X"EB",X"15",X"D1",X"D5",X"3E",X"40",X"D5",X"C9",X"13",X"01",X"03",X"00",
		X"5F",X"ED",X"98",X"1E",X"00",X"01",X"02",X"00",X"ED",X"98",X"D1",X"C1",X"D5",X"78",X"09",X"88",
		X"33",X"E3",X"0F",X"E5",X"98",X"15",X"66",X"0B",X"46",X"C5",X"09",X"80",X"04",X"21",X"26",X"01",
		X"06",X"27",X"59",X"3E",X"08",X"E5",X"BF",X"15",X"10",X"F8",X"11",X"C3",X"40",X"09",X"3F",X"31",
		X"3E",X"01",X"06",X"14",X"E5",X"D5",X"15",X"11",X"8D",X"41",X"09",X"53",X"31",X"3E",X"01",X"06",
		X"07",X"E5",X"D5",X"15",X"11",X"8F",X"40",X"09",X"72",X"31",X"3E",X"01",X"06",X"16",X"E5",X"D5",
		X"15",X"11",X"A0",X"40",X"09",X"58",X"31",X"3E",X"01",X"06",X"17",X"E5",X"D5",X"15",X"11",X"69",
		X"42",X"09",X"87",X"31",X"3E",X"01",X"06",X"20",X"E5",X"D5",X"15",X"11",X"64",X"40",X"09",X"A7",
		X"31",X"3E",X"03",X"06",X"01",X"E5",X"D5",X"15",X"11",X"A5",X"40",X"09",X"82",X"33",X"3E",X"01",
		X"06",X"32",X"E5",X"D5",X"15",X"3E",X"01",X"11",X"AD",X"47",X"12",X"AF",X"1A",X"F9",X"64",X"1A",
		X"FA",X"64",X"09",X"AD",X"47",X"0A",X"FB",X"64",X"11",X"59",X"41",X"09",X"1B",X"31",X"3E",X"01",
		X"06",X"24",X"E5",X"D5",X"15",X"09",X"77",X"33",X"11",X"DC",X"42",X"01",X"21",X"00",X"ED",X"98",
		X"AF",X"12",X"E5",X"02",X"16",X"3E",X"01",X"12",X"09",X"9B",X"64",X"11",X"94",X"42",X"E5",X"2F",
		X"11",X"11",X"95",X"42",X"E5",X"2F",X"11",X"11",X"96",X"42",X"E5",X"2F",X"11",X"11",X"97",X"42",
		X"E5",X"2F",X"11",X"11",X"B0",X"42",X"E5",X"2F",X"11",X"11",X"B1",X"42",X"E5",X"2F",X"11",X"11",
		X"B2",X"42",X"E5",X"2F",X"11",X"11",X"B3",X"42",X"E5",X"2F",X"11",X"11",X"B4",X"42",X"E5",X"2F",
		X"11",X"11",X"B5",X"42",X"E5",X"2F",X"11",X"3A",X"F8",X"64",X"E3",X"67",X"E2",X"43",X"14",X"E3",
		X"57",X"E2",X"7B",X"14",X"3A",X"F8",X"64",X"E3",X"4F",X"C2",X"BC",X"14",X"3A",X"F9",X"64",X"FE",
		X"33",X"28",X"37",X"09",X"68",X"33",X"E5",X"98",X"15",X"7E",X"C9",X"D1",X"12",X"13",X"5F",X"3E",
		X"08",X"E5",X"BF",X"15",X"D5",X"CD",X"3A",X"FA",X"64",X"3C",X"1A",X"FA",X"64",X"FE",X"03",X"C2",
		X"E7",X"14",X"09",X"9C",X"33",X"3A",X"FA",X"64",X"E5",X"98",X"15",X"7E",X"C9",X"D1",X"CD",X"E5",
		X"9D",X"15",X"09",X"DD",X"64",X"01",X"03",X"00",X"ED",X"98",X"3A",X"FA",X"64",X"FE",X"00",X"28",
		X"0D",X"09",X"B8",X"33",X"E5",X"98",X"15",X"7E",X"D1",X"E5",X"E1",X"15",X"09",X"DF",X"64",X"E5",
		X"64",X"11",X"09",X"B8",X"64",X"11",X"DA",X"43",X"E5",X"0E",X"10",X"09",X"97",X"64",X"E3",X"86",
		X"3E",X"01",X"E5",X"67",X"15",X"E1",X"D1",X"3E",X"80",X"E5",X"E1",X"15",X"3E",X"08",X"E5",X"E1",
		X"15",X"30",X"F1",X"3A",X"F9",X"64",X"FE",X"00",X"E2",X"C4",X"13",X"3D",X"1A",X"F9",X"64",X"FE",
		X"32",X"28",X"14",X"3E",X"05",X"2A",X"FB",X"64",X"5F",X"3E",X"08",X"E5",X"98",X"15",X"0A",X"FB",
		X"64",X"3E",X"01",X"5F",X"C3",X"C4",X"13",X"3D",X"1A",X"F9",X"64",X"3E",X"05",X"2A",X"FB",X"64",
		X"2B",X"5F",X"0B",X"5F",X"0B",X"5F",X"2B",X"3E",X"40",X"30",X"C8",X"3A",X"F9",X"64",X"FE",X"33",
		X"E2",X"C4",X"13",X"3C",X"1A",X"F9",X"64",X"FE",X"32",X"28",X"14",X"3E",X"05",X"2A",X"FB",X"64",
		X"5F",X"3E",X"08",X"E5",X"BF",X"15",X"0A",X"FB",X"64",X"3E",X"01",X"5F",X"C3",X"C4",X"13",X"3C",
		X"1A",X"F9",X"64",X"3E",X"05",X"2A",X"FB",X"64",X"5F",X"3E",X"40",X"E5",X"BF",X"15",X"0A",X"FB",
		X"64",X"3E",X"01",X"2B",X"5F",X"0B",X"5F",X"0B",X"5F",X"C3",X"C4",X"13",X"3E",X"20",X"E5",X"B3",
		X"15",X"1A",X"C0",X"50",X"06",X"14",X"E5",X"4F",X"15",X"F2",X"DA",X"13",X"C3",X"9F",X"13",X"3A",
		X"F8",X"64",X"E3",X"4F",X"1A",X"C0",X"50",X"28",X"DE",X"30",X"CE",X"21",X"05",X"10",X"01",X"D5",
		X"AF",X"E3",X"0B",X"17",X"E3",X"0B",X"17",X"E3",X"0B",X"17",X"E3",X"0B",X"17",X"E3",X"0B",X"17",
		X"57",X"EB",X"01",X"40",X"40",X"21",X"06",X"00",X"D1",X"62",X"21",X"EB",X"E1",X"09",X"40",X"40",
		X"11",X"41",X"40",X"01",X"7F",X"03",X"5F",X"ED",X"98",X"1A",X"C0",X"50",X"E1",X"09",X"40",X"44",
		X"11",X"41",X"44",X"01",X"7F",X"03",X"5F",X"ED",X"98",X"1A",X"C0",X"50",X"E1",X"3A",X"B3",X"64",
		X"FE",X"00",X"E0",X"3A",X"B5",X"64",X"CE",X"D8",X"E3",X"3F",X"E3",X"3F",X"E3",X"3F",X"E3",X"3F",
		X"FE",X"00",X"28",X"24",X"1A",X"25",X"40",X"3A",X"B5",X"64",X"CE",X"27",X"1A",X"24",X"40",X"E1",
		X"3E",X"40",X"30",X"D8",X"3E",X"21",X"E5",X"25",X"15",X"3E",X"40",X"E5",X"FD",X"14",X"E1",X"47",
		X"AF",X"1A",X"B6",X"64",X"1A",X"88",X"64",X"3A",X"88",X"64",X"B8",X"E0",X"09",X"95",X"64",X"E3",
		X"6E",X"C0",X"1A",X"C0",X"50",X"30",X"D8",X"3A",X"97",X"64",X"E3",X"47",X"28",X"25",X"3A",X"89",
		X"64",X"47",X"3A",X"88",X"64",X"B8",X"18",X"31",X"1F",X"3F",X"E1",X"78",X"1A",X"89",X"64",X"3A",
		X"97",X"64",X"E3",X"C7",X"1A",X"97",X"64",X"AF",X"1A",X"88",X"64",X"1A",X"B6",X"64",X"1F",X"3F",
		X"E1",X"3A",X"97",X"64",X"E3",X"87",X"1A",X"97",X"64",X"1F",X"E1",X"47",X"AF",X"1A",X"B7",X"64",
		X"3A",X"B7",X"64",X"B8",X"E0",X"09",X"95",X"64",X"E3",X"6E",X"C0",X"1A",X"C0",X"50",X"30",X"D8",
		X"85",X"6F",X"D0",X"0C",X"E1",X"83",X"77",X"D0",X"14",X"E1",X"81",X"67",X"D0",X"04",X"E1",X"D5",
		X"16",X"00",X"77",X"1F",X"3F",X"ED",X"52",X"D1",X"E1",X"CD",X"EB",X"16",X"00",X"77",X"1F",X"3F",
		X"ED",X"52",X"EB",X"C9",X"E1",X"1A",X"48",X"64",X"D5",X"3A",X"48",X"64",X"67",X"ED",X"88",X"79",
		X"FE",X"00",X"08",X"F9",X"D1",X"E5",X"02",X"16",X"10",X"EE",X"E1",X"1A",X"48",X"64",X"D5",X"3A",
		X"48",X"64",X"67",X"ED",X"88",X"2B",X"79",X"FE",X"00",X"08",X"F8",X"D1",X"E5",X"02",X"16",X"10",
		X"ED",X"E1",X"CD",X"09",X"08",X"00",X"31",X"EB",X"C9",X"E1",X"09",X"49",X"64",X"06",X"2F",X"1E",
		X"00",X"0B",X"10",X"FB",X"E1",X"09",X"95",X"64",X"E3",X"FE",X"E3",X"7E",X"E0",X"30",X"FB",X"3A",
		X"00",X"50",X"CE",X"27",X"47",X"3A",X"40",X"50",X"CE",X"D8",X"98",X"1A",X"F8",X"64",X"E1",X"3A",
		X"40",X"50",X"47",X"CE",X"27",X"E3",X"78",X"28",X"02",X"E3",X"CF",X"1A",X"F8",X"64",X"E1",X"F5",
		X"09",X"05",X"65",X"F5",X"E3",X"00",X"46",X"C4",X"58",X"17",X"F5",X"E3",X"00",X"56",X"28",X"10",
		X"E5",X"78",X"17",X"FD",X"09",X"51",X"50",X"E5",X"47",X"17",X"F5",X"7E",X"06",X"1A",X"45",X"50",
		X"F5",X"09",X"08",X"65",X"F5",X"E3",X"00",X"46",X"C4",X"58",X"17",X"F5",X"E3",X"00",X"56",X"28",
		X"10",X"E5",X"78",X"17",X"FD",X"09",X"51",X"50",X"E5",X"47",X"17",X"F5",X"7E",X"06",X"1A",X"45",
		X"50",X"F5",X"09",X"3B",X"65",X"F5",X"E3",X"00",X"46",X"C4",X"58",X"17",X"F5",X"E3",X"00",X"56",
		X"28",X"10",X"E5",X"78",X"17",X"FD",X"09",X"51",X"50",X"E5",X"47",X"17",X"F5",X"7E",X"06",X"1A",
		X"45",X"50",X"F5",X"09",X"56",X"65",X"F5",X"E3",X"00",X"46",X"C4",X"58",X"17",X"F5",X"E3",X"00",
		X"56",X"28",X"10",X"E5",X"78",X"17",X"FD",X"09",X"56",X"50",X"E5",X"47",X"17",X"F5",X"7E",X"06",
		X"1A",X"62",X"50",X"F5",X"09",X"59",X"65",X"F5",X"E3",X"00",X"46",X"C4",X"58",X"17",X"F5",X"E3",
		X"00",X"56",X"28",X"10",X"E5",X"78",X"17",X"FD",X"09",X"56",X"50",X"E5",X"47",X"17",X"F5",X"7E",
		X"06",X"1A",X"62",X"50",X"F5",X"09",X"A4",X"65",X"F5",X"E3",X"00",X"46",X"C4",X"58",X"17",X"F5",
		X"E3",X"00",X"56",X"28",X"10",X"E5",X"78",X"17",X"FD",X"09",X"56",X"50",X"E5",X"47",X"17",X"F5",
		X"7E",X"06",X"1A",X"62",X"50",X"F5",X"09",X"8F",X"65",X"F5",X"E3",X"00",X"46",X"C4",X"58",X"17",
		X"F5",X"E3",X"00",X"56",X"28",X"10",X"E5",X"78",X"17",X"FD",X"09",X"73",X"50",X"E5",X"47",X"17",
		X"F5",X"7E",X"06",X"1A",X"67",X"50",X"F5",X"09",X"C2",X"65",X"F5",X"E3",X"00",X"46",X"C4",X"58",
		X"17",X"F5",X"E3",X"00",X"56",X"E0",X"E5",X"78",X"17",X"FD",X"09",X"73",X"50",X"E5",X"47",X"17",
		X"F5",X"7E",X"06",X"1A",X"67",X"50",X"E1",X"F5",X"7E",X"03",X"FD",X"5F",X"00",X"E3",X"3F",X"E3",
		X"3F",X"E3",X"3F",X"E3",X"3F",X"FD",X"5F",X"01",X"F5",X"7E",X"04",X"FD",X"5F",X"02",X"E3",X"3F",
		X"E3",X"3F",X"E3",X"3F",X"E3",X"3F",X"FD",X"5F",X"03",X"F5",X"7E",X"05",X"FD",X"5F",X"04",X"E1",
		X"E5",X"64",X"30",X"F5",X"E3",X"00",X"D6",X"E1",X"F5",X"E3",X"00",X"66",X"C2",X"64",X"30",X"F5",
		X"6E",X"01",X"F5",X"4E",X"02",X"7E",X"E3",X"0F",X"11",X"96",X"17",X"E5",X"9D",X"15",X"0B",X"CD",
		X"32",X"6F",X"13",X"32",X"4F",X"E9",X"98",X"17",X"9C",X"17",X"C2",X"17",X"E3",X"17",X"C9",X"17",
		X"EE",X"17",X"20",X"30",X"09",X"30",X"43",X"30",X"63",X"30",X"6A",X"30",X"5E",X"30",X"82",X"30",
		X"C9",X"C3",X"85",X"17",X"C9",X"7E",X"F5",X"5F",X"03",X"0B",X"7E",X"0B",X"F5",X"5F",X"04",X"C3",
		X"85",X"17",X"C9",X"7E",X"F5",X"5F",X"05",X"0B",X"C3",X"85",X"17",X"C9",X"7E",X"F5",X"46",X"03",
		X"80",X"F5",X"5F",X"03",X"0B",X"7E",X"0B",X"F5",X"46",X"04",X"A0",X"F5",X"5F",X"04",X"C3",X"85",
		X"17",X"C9",X"7E",X"F5",X"46",X"05",X"80",X"F5",X"5F",X"05",X"0B",X"C3",X"85",X"17",X"C9",X"7E",
		X"F5",X"BE",X"07",X"28",X"23",X"F5",X"1C",X"07",X"2B",X"F5",X"5D",X"01",X"F5",X"5C",X"02",X"E1",
		X"F5",X"1E",X"07",X"00",X"0B",X"C3",X"85",X"17",X"F5",X"6E",X"20",X"F5",X"4E",X"21",X"D1",X"D5",
		X"2B",X"5A",X"2B",X"5B",X"2B",X"1E",X"00",X"F5",X"5D",X"20",X"F5",X"5C",X"21",X"C9",X"C3",X"85",
		X"17",X"D1",X"32",X"F5",X"6E",X"20",X"F5",X"4E",X"21",X"BE",X"28",X"21",X"1C",X"0B",X"76",X"0B",
		X"56",X"EB",X"C3",X"85",X"17",X"0B",X"0B",X"0B",X"F5",X"5D",X"20",X"F5",X"5C",X"21",X"13",X"EB",
		X"C3",X"85",X"17",X"C9",X"76",X"0B",X"56",X"EB",X"C3",X"85",X"17",X"C9",X"F5",X"CD",X"F5",X"CD",
		X"C9",X"D1",X"13",X"1E",X"00",X"01",X"30",X"00",X"ED",X"98",X"32",X"F5",X"5F",X"01",X"13",X"32",
		X"F5",X"5F",X"02",X"F5",X"5D",X"20",X"F5",X"5C",X"21",X"E1",X"C9",X"F5",X"5D",X"01",X"F5",X"5C",
		X"02",X"F5",X"1E",X"00",X"00",X"E1",X"C9",X"76",X"0B",X"56",X"EB",X"1E",X"06",X"13",X"EB",X"C3",
		X"85",X"17",X"C9",X"7E",X"F5",X"5F",X"06",X"0B",X"C3",X"85",X"17",X"1A",X"40",X"52",X"45",X"71",
		X"41",X"64",X"50",X"40",X"45",X"52",X"67",X"43",X"53",X"50",X"67",X"54",X"40",X"19",X"40",X"52",
		X"45",X"71",X"41",X"64",X"50",X"54",X"61",X"44",X"45",X"52",X"43",X"71",X"41",X"64",X"50",X"45",
		X"45",X"52",X"46",X"40",X"66",X"61",X"67",X"43",X"40",X"54",X"52",X"45",X"53",X"66",X"61",X"52",
		X"45",X"71",X"41",X"64",X"50",X"40",X"45",X"66",X"67",X"40",X"54",X"43",X"45",X"64",X"45",X"53",
		X"52",X"67",X"53",X"52",X"45",X"71",X"41",X"64",X"50",X"40",X"67",X"57",X"54",X"40",X"52",X"67",
		X"40",X"45",X"66",X"67",X"40",X"54",X"43",X"45",X"64",X"45",X"53",X"50",X"55",X"40",X"45",X"66",
		X"67",X"40",X"52",X"45",X"71",X"41",X"64",X"50",X"50",X"55",X"40",X"67",X"57",X"54",X"40",X"52",
		X"45",X"71",X"41",X"64",X"50",X"66",X"61",X"41",X"47",X"41",X"40",X"52",X"45",X"71",X"41",X"64",
		X"50",X"40",X"45",X"65",X"41",X"53",X"52",X"45",X"56",X"67",X"40",X"45",X"65",X"41",X"47",X"52",
		X"45",X"56",X"67",X"40",X"45",X"65",X"41",X"47",X"40",X"45",X"66",X"67",X"40",X"52",X"45",X"71",
		X"41",X"64",X"50",X"45",X"65",X"41",X"46",X"40",X"46",X"67",X"40",X"64",X"64",X"41",X"60",X"45",
		X"60",X"54",X"40",X"66",X"61",X"40",X"53",X"61",X"40",X"45",X"52",X"67",X"43",X"53",X"40",X"52",
		X"55",X"67",X"71",X"66",X"45",X"54",X"40",X"50",X"67",X"54",X"54",X"43",X"45",X"64",X"45",X"53",
		X"40",X"67",X"54",X"40",X"63",X"43",X"61",X"54",X"53",X"71",X"67",X"62",X"40",X"45",X"53",X"55",
		X"66",X"67",X"54",X"54",X"55",X"42",X"40",X"44",X"45",X"45",X"50",X"53",X"40",X"44",X"66",X"41",
		X"40",X"52",X"45",X"54",X"54",X"45",X"64",X"54",X"66",X"61",X"52",X"50",X"40",X"67",X"54",X"45",
		X"66",X"44",X"65",X"41",X"64",X"53",X"45",X"43",X"66",X"41",X"56",X"44",X"41",X"40",X"45",X"52",
		X"67",X"43",X"53",X"40",X"54",X"66",X"54",X"40",X"52",X"65",X"40",X"45",X"52",X"67",X"43",X"53",
		X"40",X"40",X"53",X"66",X"67",X"61",X"54",X"43",X"45",X"53",X"52",X"45",X"54",X"66",X"61",X"52",
		X"45",X"42",X"65",X"55",X"66",X"40",X"45",X"65",X"41",X"52",X"46",X"40",X"70",X"40",X"53",X"54",
		X"66",X"61",X"67",X"50",X"40",X"18",X"19",X"53",X"66",X"67",X"61",X"54",X"43",X"45",X"53",X"52",
		X"45",X"54",X"66",X"61",X"40",X"40",X"64",X"41",X"61",X"43",X"45",X"50",X"53",X"4C",X"4C",X"4C",
		X"4C",X"40",X"40",X"40",X"45",X"52",X"67",X"43",X"53",X"40",X"71",X"41",X"64",X"50",X"40",X"19",
		X"40",X"53",X"66",X"61",X"67",X"43",X"40",X"1A",X"53",X"71",X"41",X"64",X"50",X"40",X"1A",X"40",
		X"40",X"66",X"61",X"67",X"43",X"40",X"19",X"40",X"71",X"41",X"64",X"50",X"40",X"19",X"40",X"40",
		X"66",X"61",X"67",X"43",X"40",X"19",X"53",X"54",X"66",X"61",X"67",X"50",X"40",X"40",X"40",X"40",
		X"40",X"40",X"40",X"40",X"71",X"52",X"45",X"56",X"45",X"40",X"53",X"55",X"66",X"67",X"42",X"18",
		X"18",X"18",X"18",X"1D",X"19",X"18",X"18",X"18",X"1D",X"1A",X"19",X"18",X"18",X"18",X"18",X"18",
		X"19",X"40",X"18",X"18",X"18",X"1D",X"1F",X"53",X"43",X"61",X"54",X"53",X"67",X"66",X"47",X"41",
		X"61",X"44",X"66",X"67",X"61",X"54",X"61",X"44",X"66",X"67",X"43",X"40",X"40",X"66",X"67",X"61",
		X"54",X"41",X"43",X"67",X"64",X"40",X"40",X"65",X"67",X"52",X"44",X"67",X"67",X"47",X"40",X"40",
		X"40",X"40",X"40",X"40",X"40",X"44",X"1F",X"40",X"40",X"40",X"40",X"40",X"40",X"19",X"44",X"67",
		X"67",X"47",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"46",X"1F",X"40",X"40",X"40",X"40",X"40",
		X"40",X"1A",X"44",X"67",X"67",X"47",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"60",X"1F",X"40",
		X"40",X"40",X"40",X"40",X"40",X"1B",X"44",X"67",X"67",X"47",X"40",X"40",X"40",X"40",X"40",X"40",
		X"40",X"62",X"1F",X"40",X"40",X"40",X"40",X"40",X"40",X"1C",X"44",X"67",X"67",X"47",X"40",X"40",
		X"40",X"40",X"40",X"40",X"40",X"60",X"1C",X"40",X"40",X"40",X"40",X"40",X"40",X"19",X"44",X"67",
		X"67",X"47",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"64",X"1C",X"40",X"40",X"40",X"40",X"40",
		X"40",X"1A",X"44",X"67",X"67",X"47",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"62",X"1C",X"40",
		X"40",X"40",X"40",X"40",X"40",X"1B",X"44",X"67",X"67",X"47",X"40",X"40",X"40",X"40",X"40",X"40",
		X"40",X"65",X"1C",X"40",X"40",X"40",X"40",X"40",X"40",X"1C",X"44",X"67",X"67",X"47",X"40",X"40",
		X"40",X"40",X"40",X"40",X"40",X"63",X"1C",X"40",X"40",X"40",X"40",X"40",X"40",X"1D",X"44",X"67",
		X"67",X"47",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"66",X"1C",X"40",X"40",X"40",X"40",X"40",
		X"40",X"1E",X"44",X"41",X"42",X"40",X"66",X"67",X"61",X"54",X"61",X"44",X"66",X"67",X"43",X"40",
		X"40",X"66",X"67",X"61",X"54",X"41",X"43",X"67",X"64",X"40",X"40",X"65",X"41",X"52",X"00",X"01",
		X"02",X"03",X"04",X"05",X"06",X"07",X"20",X"21",X"41",X"42",X"43",X"44",X"45",X"46",X"47",X"60",
		X"61",X"62",X"63",X"64",X"65",X"66",X"67",X"50",X"51",X"52",X"53",X"54",X"55",X"56",X"57",X"70",
		X"71",X"72",X"72",X"71",X"70",X"57",X"56",X"55",X"54",X"53",X"52",X"51",X"50",X"67",X"66",X"65",
		X"64",X"63",X"62",X"61",X"60",X"47",X"46",X"45",X"44",X"43",X"42",X"41",X"00",X"01",X"04",X"02",
		X"94",X"42",X"95",X"42",X"96",X"42",X"97",X"42",X"B0",X"42",X"B1",X"42",X"B2",X"42",X"B3",X"42",
		X"B4",X"42",X"B5",X"42",X"03",X"02",X"01",X"00",X"00",X"80",X"48",X"40",X"09",X"F5",X"65",X"E3",
		X"46",X"08",X"11",X"E3",X"C6",X"3A",X"2C",X"66",X"2A",X"0F",X"66",X"06",X"10",X"76",X"0B",X"56",
		X"12",X"0B",X"10",X"F9",X"00",X"3E",X"04",X"1A",X"15",X"66",X"3A",X"29",X"66",X"1A",X"16",X"66",
		X"09",X"DA",X"0E",X"11",X"17",X"66",X"01",X"04",X"00",X"ED",X"98",X"FD",X"09",X"A1",X"64",X"FD",
		X"7E",X"07",X"CE",X"C8",X"47",X"3A",X"F8",X"64",X"CE",X"37",X"98",X"FD",X"5F",X"07",X"2A",X"11",
		X"66",X"0A",X"27",X"66",X"09",X"F8",X"65",X"E5",X"3F",X"37",X"09",X"00",X"00",X"0A",X"27",X"66",
		X"3A",X"13",X"66",X"1A",X"15",X"66",X"3A",X"14",X"66",X"1A",X"16",X"66",X"09",X"DE",X"0E",X"11",
		X"17",X"66",X"01",X"04",X"00",X"ED",X"98",X"3A",X"33",X"66",X"FE",X"9D",X"28",X"0D",X"FE",X"3C",
		X"28",X"22",X"FE",X"78",X"28",X"25",X"FE",X"9C",X"28",X"10",X"30",X"13",X"09",X"58",X"64",X"E3",
		X"DE",X"30",X"24",X"09",X"78",X"64",X"E3",X"DE",X"30",X"05",X"09",X"80",X"64",X"E3",X"DE",X"3C",
		X"1A",X"33",X"66",X"00",X"F5",X"09",X"A1",X"64",X"FD",X"09",X"49",X"64",X"E5",X"22",X"0F",X"09",
		X"FB",X"65",X"E5",X"3F",X"37",X"F5",X"09",X"A1",X"64",X"FD",X"09",X"69",X"64",X"E5",X"22",X"0F",
		X"09",X"FE",X"65",X"E5",X"3F",X"37",X"F5",X"09",X"A1",X"64",X"FD",X"09",X"59",X"64",X"E5",X"22",
		X"0F",X"09",X"01",X"66",X"E5",X"3F",X"37",X"F5",X"09",X"A1",X"64",X"FD",X"09",X"79",X"64",X"E5",
		X"22",X"0F",X"09",X"04",X"66",X"E5",X"3F",X"37",X"F5",X"09",X"A1",X"64",X"FD",X"09",X"81",X"64",
		X"E5",X"22",X"0F",X"09",X"07",X"66",X"E5",X"3F",X"37",X"3A",X"2B",X"66",X"3C",X"1A",X"2B",X"66",
		X"FE",X"04",X"08",X"2C",X"AF",X"1A",X"2B",X"66",X"3A",X"2A",X"66",X"47",X"FE",X"02",X"28",X"35",
		X"3C",X"1A",X"2A",X"66",X"3A",X"2C",X"66",X"80",X"67",X"2A",X"0F",X"66",X"06",X"10",X"76",X"0B",
		X"56",X"0B",X"32",X"FE",X"4E",X"38",X"02",X"79",X"12",X"10",X"DB",X"30",X"03",X"AF",X"30",X"C9",
		X"00",X"3A",X"84",X"64",X"FE",X"00",X"28",X"12",X"3A",X"0E",X"66",X"3C",X"1A",X"0E",X"66",X"FE",
		X"1A",X"08",X"07",X"AF",X"1A",X"84",X"64",X"1A",X"0E",X"66",X"3A",X"0A",X"66",X"FE",X"04",X"08",
		X"0A",X"AF",X"1A",X"0A",X"66",X"3A",X"18",X"40",X"47",X"3A",X"2F",X"40",X"67",X"3A",X"0B",X"66",
		X"1A",X"18",X"40",X"3A",X"0C",X"66",X"1A",X"2F",X"40",X"78",X"1A",X"0B",X"66",X"79",X"1A",X"0C",
		X"66",X"30",X"04",X"3C",X"1A",X"0A",X"66",X"3A",X"0D",X"66",X"FE",X"FF",X"E2",X"26",X"36",X"FE",
		X"10",X"C2",X"29",X"36",X"3C",X"1A",X"0D",X"66",X"3A",X"4C",X"64",X"1A",X"2F",X"66",X"3A",X"6C",
		X"64",X"1A",X"18",X"66",X"3A",X"5C",X"64",X"1A",X"19",X"66",X"3A",X"7C",X"64",X"1A",X"1A",X"66",
		X"3A",X"84",X"64",X"1A",X"1B",X"66",X"3A",X"A4",X"64",X"1A",X"1C",X"66",X"AF",X"1A",X"4C",X"64",
		X"1A",X"6C",X"64",X"1A",X"5C",X"64",X"1A",X"7C",X"64",X"1A",X"84",X"64",X"1A",X"A4",X"64",X"06",
		X"34",X"09",X"66",X"40",X"11",X"1D",X"66",X"C5",X"01",X"05",X"00",X"ED",X"98",X"3E",X"33",X"E5",
		X"98",X"15",X"C1",X"10",X"DA",X"3A",X"40",X"44",X"1A",X"C1",X"66",X"11",X"66",X"40",X"09",X"CB",
		X"36",X"3E",X"05",X"06",X"34",X"E5",X"EB",X"15",X"11",X"66",X"44",X"09",X"3E",X"37",X"3E",X"05",
		X"06",X"34",X"E5",X"EB",X"15",X"11",X"6F",X"40",X"09",X"CC",X"36",X"3E",X"01",X"06",X"32",X"E5",
		X"D5",X"15",X"11",X"11",X"41",X"09",X"FE",X"36",X"3E",X"01",X"06",X"10",X"E5",X"D5",X"15",X"3E",
		X"78",X"E5",X"B3",X"15",X"11",X"66",X"44",X"09",X"C1",X"66",X"3E",X"05",X"06",X"34",X"E5",X"EB",
		X"15",X"06",X"34",X"09",X"1D",X"66",X"11",X"66",X"40",X"C5",X"01",X"05",X"00",X"ED",X"98",X"3E",
		X"33",X"E5",X"9D",X"15",X"C1",X"10",X"DA",X"3A",X"2F",X"66",X"1A",X"4C",X"64",X"3A",X"18",X"66",
		X"1A",X"6C",X"64",X"3A",X"19",X"66",X"1A",X"5C",X"64",X"3A",X"1A",X"66",X"1A",X"7C",X"64",X"3A",
		X"1B",X"66",X"1A",X"84",X"64",X"3A",X"1C",X"66",X"1A",X"A4",X"64",X"C3",X"29",X"36",X"AF",X"1A",
		X"4A",X"64",X"1A",X"6A",X"64",X"1A",X"5A",X"64",X"1A",X"7A",X"64",X"1A",X"82",X"64",X"1A",X"A2",
		X"64",X"09",X"59",X"65",X"E3",X"E6",X"C3",X"E0",X"36",X"3A",X"90",X"64",X"E3",X"6F",X"C2",X"CA",
		X"36",X"E3",X"5F",X"08",X"10",X"09",X"96",X"64",X"E3",X"E6",X"3E",X"40",X"1A",X"2F",X"40",X"1A",
		X"18",X"40",X"C3",X"CA",X"36",X"3A",X"68",X"64",X"47",X"3A",X"58",X"64",X"98",X"47",X"3A",X"78",
		X"64",X"98",X"47",X"3A",X"80",X"64",X"98",X"47",X"3A",X"A0",X"64",X"98",X"E3",X"5F",X"C2",X"CA",
		X"36",X"47",X"AF",X"1A",X"A2",X"64",X"09",X"59",X"65",X"E3",X"E6",X"09",X"A4",X"65",X"E3",X"E6",
		X"E3",X"68",X"08",X"6E",X"AF",X"1A",X"A4",X"64",X"3A",X"40",X"44",X"1A",X"C1",X"66",X"11",X"66",
		X"40",X"09",X"CB",X"36",X"3E",X"05",X"06",X"34",X"E5",X"EB",X"15",X"11",X"66",X"44",X"09",X"3E",
		X"37",X"3E",X"05",X"06",X"34",X"E5",X"EB",X"15",X"11",X"2F",X"41",X"09",X"26",X"37",X"3E",X"01",
		X"06",X"27",X"E5",X"D5",X"15",X"11",X"D1",X"40",X"09",X"35",X"37",X"3E",X"01",X"06",X"14",X"E5",
		X"D5",X"15",X"3E",X"78",X"E5",X"B3",X"15",X"11",X"66",X"44",X"09",X"C1",X"66",X"3E",X"05",X"06",
		X"34",X"E5",X"EB",X"15",X"AF",X"1A",X"84",X"64",X"3A",X"84",X"64",X"FE",X"00",X"08",X"13",X"09",
		X"96",X"64",X"E3",X"F6",X"E3",X"E6",X"AF",X"1A",X"33",X"66",X"3E",X"40",X"1A",X"2F",X"40",X"1A",
		X"18",X"40",X"E1",X"40",X"45",X"53",X"55",X"46",X"40",X"71",X"42",X"40",X"44",X"45",X"66",X"52",
		X"55",X"42",X"40",X"54",X"45",X"47",X"52",X"41",X"54",X"40",X"54",X"53",X"41",X"64",X"66",X"55",
		X"52",X"40",X"54",X"53",X"55",X"65",X"40",X"55",X"67",X"71",X"40",X"57",X"67",X"66",X"53",X"66",
		X"67",X"61",X"54",X"41",X"64",X"55",X"54",X"41",X"52",X"47",X"66",X"67",X"43",X"54",X"55",X"67",
		X"40",X"44",X"45",X"66",X"52",X"55",X"42",X"40",X"53",X"45",X"53",X"55",X"46",X"40",X"64",X"64",
		X"41",X"71",X"52",X"52",X"67",X"53",X"44",X"66",X"45",X"40",X"44",X"41",X"45",X"44",X"21",X"F5",
		X"2A",X"DE",X"65",X"FD",X"E3",X"07",X"6E",X"C2",X"5B",X"0B",X"FD",X"E3",X"07",X"5E",X"E0",X"7E",
		X"E3",X"BF",X"E3",X"9F",X"FE",X"03",X"E2",X"0F",X"0B",X"3C",X"47",X"7E",X"CE",X"C0",X"98",X"5F",
		X"3E",X"DB",X"FD",X"46",X"03",X"90",X"1A",X"75",X"64",X"FD",X"7E",X"04",X"D6",X"24",X"1A",X"74",
		X"64",X"CD",X"E5",X"BD",X"26",X"C9",X"3A",X"22",X"64",X"FE",X"00",X"C2",X"20",X"0B",X"3A",X"23",
		X"64",X"FE",X"00",X"C2",X"20",X"0B",X"E3",X"5E",X"C2",X"00",X"0B",X"E3",X"DE",X"32",X"1A",X"22",
		X"66",X"D5",X"33",X"32",X"1A",X"23",X"66",X"13",X"13",X"32",X"1A",X"24",X"66",X"3E",X"09",X"E5",
		X"E1",X"15",X"32",X"1A",X"25",X"66",X"3E",X"40",X"E5",X"9D",X"15",X"32",X"1A",X"26",X"66",X"D1",
		X"E3",X"7E",X"C2",X"B7",X"08",X"3A",X"C2",X"66",X"FE",X"00",X"E2",X"B7",X"08",X"FE",X"01",X"28",
		X"02",X"30",X"56",X"3A",X"90",X"64",X"E3",X"47",X"28",X"07",X"E3",X"77",X"28",X"0F",X"E3",X"9E",
		X"E1",X"FD",X"46",X"00",X"FD",X"1E",X"00",X"02",X"3A",X"30",X"66",X"FD",X"5F",X"05",X"AF",X"1A",
		X"C2",X"66",X"78",X"FE",X"04",X"28",X"07",X"F5",X"7E",X"02",X"12",X"C3",X"6B",X"0A",X"F5",X"7E",
		X"03",X"12",X"C3",X"6B",X"0A",X"FD",X"46",X"00",X"FD",X"1E",X"00",X"03",X"3A",X"17",X"66",X"FD",
		X"5F",X"05",X"AF",X"1A",X"C2",X"66",X"78",X"FE",X"04",X"28",X"07",X"F5",X"7E",X"04",X"12",X"C3",
		X"6B",X"0A",X"F5",X"7E",X"05",X"12",X"C3",X"6B",X"0A",X"3A",X"90",X"64",X"E3",X"67",X"28",X"07",
		X"E3",X"57",X"28",X"0F",X"E3",X"9E",X"E1",X"FD",X"46",X"00",X"FD",X"1E",X"00",X"05",X"3A",X"31",
		X"66",X"FD",X"5F",X"05",X"AF",X"1A",X"C2",X"66",X"78",X"FE",X"02",X"28",X"07",X"F5",X"7E",X"03",
		X"12",X"C3",X"41",X"09",X"F5",X"7E",X"05",X"12",X"C3",X"41",X"09",X"FD",X"46",X"00",X"FD",X"1E",
		X"00",X"04",X"3A",X"32",X"66",X"FD",X"5F",X"05",X"AF",X"1A",X"C2",X"66",X"78",X"FE",X"02",X"28",
		X"07",X"F5",X"7E",X"02",X"12",X"C3",X"41",X"09",X"F5",X"7E",X"04",X"12",X"C3",X"41",X"09",X"FD",
		X"E3",X"07",X"46",X"C0",X"AF",X"1A",X"C2",X"66",X"C3",X"6B",X"0A",X"FD",X"E3",X"07",X"76",X"C0",
		X"AF",X"1A",X"C2",X"66",X"C3",X"6B",X"0A",X"FD",X"E3",X"07",X"56",X"C0",X"AF",X"1A",X"C2",X"66",
		X"C3",X"41",X"09",X"FD",X"E3",X"07",X"66",X"C0",X"AF",X"1A",X"C2",X"66",X"C3",X"41",X"09",X"FD",
		X"7E",X"00",X"FE",X"02",X"E2",X"D6",X"09",X"FE",X"03",X"E2",X"D6",X"09",X"FD",X"E3",X"07",X"46",
		X"08",X"2F",X"3A",X"22",X"66",X"F5",X"BE",X"01",X"E2",X"C3",X"08",X"FE",X"4E",X"F2",X"52",X"09",
		X"E5",X"E1",X"0F",X"E5",X"33",X"28",X"FD",X"7E",X"00",X"FE",X"05",X"28",X"22",X"F5",X"7E",X"03",
		X"1A",X"22",X"66",X"12",X"C3",X"99",X"09",X"F5",X"7E",X"02",X"1A",X"22",X"66",X"12",X"C3",X"99",
		X"09",X"FD",X"E3",X"07",X"76",X"E2",X"06",X"09",X"3A",X"22",X"66",X"F5",X"BE",X"01",X"E2",X"F9",
		X"08",X"FE",X"4E",X"F2",X"52",X"09",X"E5",X"E1",X"0F",X"E5",X"33",X"28",X"F5",X"7E",X"07",X"1A",
		X"22",X"66",X"12",X"C3",X"83",X"09",X"3A",X"22",X"66",X"F5",X"BE",X"01",X"28",X"20",X"FE",X"4E",
		X"F2",X"52",X"09",X"E5",X"E1",X"0F",X"E5",X"33",X"28",X"FD",X"7E",X"00",X"FE",X"05",X"28",X"29",
		X"F5",X"7E",X"05",X"1A",X"22",X"66",X"12",X"3A",X"17",X"66",X"FD",X"5F",X"05",X"FD",X"1E",X"00",
		X"03",X"3A",X"24",X"66",X"F5",X"BE",X"00",X"E2",X"EC",X"0C",X"C3",X"39",X"0D",X"FD",X"E3",X"07",
		X"FE",X"FD",X"0A",X"91",X"64",X"E5",X"F1",X"24",X"E1",X"F5",X"7E",X"04",X"1A",X"22",X"66",X"12",
		X"30",X"D5",X"FD",X"7E",X"00",X"FE",X"05",X"28",X"11",X"3A",X"22",X"66",X"F5",X"BE",X"02",X"08",
		X"13",X"F5",X"7E",X"20",X"1A",X"22",X"66",X"12",X"30",X"BD",X"3A",X"22",X"66",X"F5",X"BE",X"03",
		X"08",X"02",X"30",X"ED",X"3A",X"22",X"66",X"F5",X"BE",X"06",X"08",X"37",X"F5",X"7E",X"20",X"1A",
		X"22",X"66",X"12",X"FD",X"7E",X"00",X"FE",X"05",X"28",X"24",X"3A",X"25",X"66",X"F5",X"BE",X"00",
		X"E2",X"D6",X"0C",X"C3",X"41",X"09",X"3A",X"26",X"66",X"30",X"DA",X"FD",X"7E",X"00",X"FE",X"05",
		X"28",X"0D",X"3A",X"22",X"66",X"F5",X"BE",X"04",X"08",X"0F",X"F5",X"7E",X"20",X"1A",X"22",X"66",
		X"12",X"3A",X"30",X"66",X"FD",X"5F",X"05",X"FD",X"1E",X"00",X"02",X"3A",X"23",X"66",X"F5",X"BE",
		X"00",X"E2",X"8E",X"0C",X"C3",X"34",X"0D",X"3A",X"22",X"66",X"F5",X"BE",X"05",X"08",X"02",X"30",
		X"F1",X"FD",X"E3",X"07",X"EE",X"E1",X"FD",X"E3",X"07",X"56",X"08",X"2F",X"3A",X"22",X"66",X"F5",
		X"BE",X"01",X"E2",X"ED",X"09",X"FE",X"4E",X"F2",X"7C",X"0A",X"E5",X"E1",X"0F",X"E5",X"33",X"28",
		X"FD",X"7E",X"00",X"FE",X"03",X"28",X"22",X"F5",X"7E",X"04",X"1A",X"22",X"66",X"12",X"C3",X"F3",
		X"0A",X"F5",X"7E",X"02",X"1A",X"22",X"66",X"12",X"C3",X"F3",X"0A",X"FD",X"E3",X"07",X"66",X"E2",
		X"18",X"0A",X"3A",X"22",X"66",X"F5",X"BE",X"01",X"E2",X"0B",X"0A",X"FE",X"4E",X"F2",X"7C",X"0A",
		X"E5",X"E1",X"0F",X"E5",X"33",X"28",X"F5",X"7E",X"06",X"1A",X"22",X"66",X"12",X"C3",X"AD",X"0A",
		X"3A",X"22",X"66",X"F5",X"BE",X"01",X"28",X"20",X"FE",X"4E",X"F2",X"7C",X"0A",X"E5",X"E1",X"0F",
		X"E5",X"33",X"28",X"FD",X"7E",X"00",X"FE",X"03",X"28",X"29",X"F5",X"7E",X"05",X"1A",X"22",X"66",
		X"12",X"3A",X"31",X"66",X"FD",X"5F",X"05",X"FD",X"1E",X"00",X"05",X"3A",X"26",X"66",X"F5",X"BE",
		X"00",X"E2",X"B4",X"0D",X"C3",X"E9",X"0D",X"FD",X"E3",X"07",X"FE",X"FD",X"0A",X"91",X"64",X"E5",
		X"F1",X"24",X"E1",X"F5",X"7E",X"03",X"1A",X"22",X"66",X"12",X"30",X"D5",X"FD",X"7E",X"00",X"FE",
		X"03",X"28",X"11",X"3A",X"22",X"66",X"F5",X"BE",X"02",X"08",X"13",X"F5",X"7E",X"20",X"1A",X"22",
		X"66",X"12",X"30",X"BD",X"3A",X"22",X"66",X"F5",X"BE",X"04",X"08",X"02",X"30",X"ED",X"3A",X"22",
		X"66",X"F5",X"BE",X"07",X"08",X"37",X"F5",X"7E",X"20",X"1A",X"22",X"66",X"12",X"FD",X"7E",X"00",
		X"FE",X"03",X"28",X"24",X"3A",X"23",X"66",X"F5",X"BE",X"00",X"E2",X"86",X"0D",X"C3",X"6B",X"0A",
		X"3A",X"24",X"66",X"30",X"DA",X"FD",X"7E",X"00",X"FE",X"03",X"28",X"0D",X"3A",X"22",X"66",X"F5",
		X"BE",X"03",X"08",X"0F",X"F5",X"7E",X"20",X"1A",X"22",X"66",X"12",X"3A",X"32",X"66",X"FD",X"5F",
		X"05",X"FD",X"1E",X"00",X"04",X"3A",X"25",X"66",X"F5",X"BE",X"00",X"E2",X"56",X"0D",X"C3",X"E4",
		X"0D",X"3A",X"22",X"66",X"F5",X"BE",X"05",X"08",X"02",X"30",X"F1",X"FD",X"E3",X"07",X"EE",X"E1",
		X"FD",X"0A",X"91",X"64",X"E5",X"F1",X"24",X"E1",X"E3",X"9E",X"E3",X"7E",X"08",X"DA",X"3A",X"C2",
		X"66",X"FE",X"00",X"28",X"EB",X"FE",X"03",X"E2",X"6F",X"08",X"FE",X"04",X"E2",X"7B",X"08",X"FE",
		X"05",X"E2",X"87",X"08",X"C3",X"93",X"08",X"3E",X"C0",X"8E",X"5F",X"E3",X"7F",X"08",X"36",X"FD",
		X"7E",X"01",X"FE",X"00",X"E0",X"FD",X"E3",X"07",X"4E",X"C2",X"56",X"0B",X"3A",X"15",X"66",X"FD",
		X"46",X"01",X"B8",X"E2",X"48",X"37",X"05",X"FD",X"58",X"01",X"C3",X"48",X"37",X"E5",X"B8",X"0F",
		X"FD",X"E3",X"07",X"7E",X"08",X"11",X"3A",X"16",X"66",X"FD",X"46",X"01",X"B8",X"E2",X"48",X"37",
		X"04",X"FD",X"58",X"01",X"C3",X"48",X"37",X"FD",X"E3",X"07",X"BE",X"3A",X"15",X"66",X"FD",X"5F",
		X"01",X"30",X"CB",X"0B",X"7E",X"FE",X"02",X"08",X"31",X"1E",X"00",X"0B",X"7E",X"FE",X"00",X"28",
		X"13",X"FE",X"27",X"E2",X"CF",X"0E",X"1C",X"09",X"FA",X"0E",X"E5",X"98",X"15",X"7E",X"FD",X"5F",
		X"05",X"E1",X"1C",X"E1",X"1C",X"2B",X"2B",X"FD",X"E3",X"07",X"9E",X"E3",X"7E",X"28",X"26",X"3A",
		X"08",X"65",X"FE",X"00",X"08",X"C9",X"09",X"3B",X"65",X"E3",X"C6",X"30",X"F2",X"09",X"56",X"65",
		X"E3",X"C6",X"09",X"68",X"64",X"E3",X"9E",X"09",X"58",X"64",X"E3",X"9E",X"09",X"78",X"64",X"E3",
		X"9E",X"09",X"80",X"64",X"E3",X"9E",X"09",X"A0",X"64",X"E3",X"9E",X"09",X"90",X"64",X"E3",X"AE",
		X"E3",X"9E",X"3E",X"9D",X"1A",X"33",X"66",X"E5",X"22",X"16",X"3E",X"17",X"E5",X"FD",X"14",X"3E",
		X"14",X"E5",X"25",X"15",X"3E",X"02",X"E5",X"B3",X"15",X"3E",X"14",X"E5",X"FD",X"14",X"3E",X"03",
		X"E5",X"B3",X"15",X"3E",X"17",X"E5",X"FD",X"14",X"3E",X"02",X"E5",X"B3",X"15",X"3E",X"14",X"E5",
		X"FD",X"14",X"3E",X"03",X"E5",X"B3",X"15",X"3E",X"17",X"E5",X"FD",X"14",X"3E",X"02",X"E5",X"B3",
		X"15",X"3E",X"14",X"E5",X"FD",X"14",X"09",X"96",X"64",X"E3",X"46",X"E0",X"3E",X"90",X"E5",X"B3",
		X"15",X"C3",X"78",X"0C",X"09",X"87",X"0E",X"E5",X"19",X"2C",X"3E",X"01",X"E5",X"B3",X"15",X"E5",
		X"81",X"0C",X"3A",X"4C",X"64",X"FE",X"00",X"08",X"D9",X"3A",X"98",X"64",X"FE",X"00",X"08",X"10",
		X"3A",X"8E",X"64",X"FE",X"00",X"08",X"21",X"3A",X"8F",X"64",X"FE",X"00",X"08",X"02",X"30",X"28",
		X"09",X"A4",X"65",X"E3",X"C6",X"3E",X"18",X"E5",X"B3",X"15",X"09",X"9F",X"0E",X"E5",X"19",X"2C",
		X"3E",X"01",X"E5",X"B3",X"15",X"E5",X"81",X"0C",X"09",X"81",X"64",X"0A",X"91",X"64",X"E5",X"F1",
		X"24",X"3A",X"4C",X"64",X"FE",X"EC",X"08",X"E8",X"E5",X"22",X"16",X"09",X"90",X"64",X"E3",X"AE",
		X"E1",X"09",X"49",X"64",X"0A",X"91",X"64",X"E5",X"F1",X"24",X"09",X"69",X"64",X"0A",X"91",X"64",
		X"E5",X"F1",X"24",X"09",X"59",X"64",X"0A",X"91",X"64",X"E5",X"F1",X"24",X"09",X"79",X"64",X"0A",
		X"91",X"64",X"E5",X"F1",X"24",X"E1",X"E3",X"7E",X"C2",X"D1",X"09",X"3A",X"22",X"66",X"F5",X"BE",
		X"20",X"E2",X"39",X"0E",X"F5",X"BE",X"03",X"08",X"11",X"3A",X"32",X"66",X"FD",X"5F",X"05",X"FD",
		X"1E",X"00",X"04",X"F5",X"7E",X"07",X"12",X"C3",X"41",X"09",X"3A",X"31",X"66",X"FD",X"5F",X"05",
		X"FD",X"1E",X"00",X"05",X"30",X"ED",X"E3",X"7E",X"C2",X"D1",X"09",X"3A",X"22",X"66",X"F5",X"BE",
		X"20",X"E2",X"39",X"0E",X"3E",X"01",X"1A",X"C2",X"66",X"E3",X"9E",X"E1",X"E3",X"7E",X"C2",X"D1",
		X"09",X"3A",X"22",X"66",X"F5",X"BE",X"20",X"E2",X"39",X"0E",X"F5",X"BE",X"05",X"08",X"11",X"3A",
		X"32",X"66",X"FD",X"5F",X"05",X"FD",X"1E",X"00",X"04",X"F5",X"7E",X"07",X"12",X"C3",X"41",X"09",
		X"3A",X"31",X"66",X"FD",X"5F",X"05",X"FD",X"1E",X"00",X"05",X"30",X"ED",X"E3",X"7E",X"C2",X"3D",
		X"09",X"3A",X"22",X"66",X"F5",X"BE",X"20",X"C2",X"41",X"09",X"FD",X"E3",X"07",X"46",X"E2",X"41",
		X"09",X"3E",X"03",X"1A",X"C2",X"66",X"C3",X"41",X"09",X"E3",X"7E",X"C2",X"3D",X"09",X"3A",X"22",
		X"66",X"F5",X"BE",X"20",X"C2",X"41",X"09",X"FD",X"E3",X"07",X"76",X"E2",X"41",X"09",X"3E",X"04",
		X"1A",X"C2",X"66",X"C3",X"41",X"09",X"E3",X"7E",X"C2",X"FB",X"0A",X"3A",X"22",X"66",X"F5",X"BE",
		X"20",X"E2",X"39",X"0E",X"F5",X"BE",X"04",X"08",X"11",X"3A",X"30",X"66",X"FD",X"5F",X"05",X"FD",
		X"1E",X"00",X"02",X"F5",X"7E",X"06",X"12",X"C3",X"6B",X"0A",X"3A",X"17",X"66",X"FD",X"5F",X"05",
		X"FD",X"1E",X"00",X"03",X"30",X"ED",X"E3",X"7E",X"C2",X"FB",X"0A",X"3A",X"22",X"66",X"F5",X"BE",
		X"20",X"E2",X"39",X"0E",X"3E",X"02",X"1A",X"C2",X"66",X"E3",X"9E",X"E1",X"E3",X"7E",X"C2",X"FB",
		X"0A",X"3A",X"22",X"66",X"F5",X"BE",X"20",X"E2",X"39",X"0E",X"F5",X"BE",X"05",X"08",X"11",X"3A",
		X"30",X"66",X"FD",X"5F",X"05",X"FD",X"1E",X"00",X"02",X"F5",X"7E",X"06",X"12",X"C3",X"6B",X"0A",
		X"3A",X"17",X"66",X"FD",X"5F",X"05",X"FD",X"1E",X"00",X"03",X"30",X"ED",X"E3",X"7E",X"C2",X"4F",
		X"0A",X"3A",X"22",X"66",X"F5",X"BE",X"20",X"C2",X"6B",X"0A",X"FD",X"E3",X"07",X"56",X"E2",X"6B",
		X"0A",X"3E",X"05",X"1A",X"C2",X"66",X"C3",X"6B",X"0A",X"E3",X"7E",X"C2",X"4F",X"0A",X"3A",X"22",
		X"66",X"F5",X"BE",X"20",X"C2",X"6B",X"0A",X"FD",X"E3",X"07",X"66",X"E2",X"6B",X"0A",X"3E",X"06",
		X"1A",X"C2",X"66",X"C3",X"6B",X"0A",X"FD",X"7E",X"07",X"47",X"FD",X"7E",X"00",X"FE",X"02",X"28",
		X"10",X"FE",X"03",X"28",X"14",X"FE",X"05",X"28",X"30",X"E3",X"60",X"E2",X"3C",X"0B",X"C3",X"56",
		X"0B",X"E3",X"70",X"E2",X"3C",X"0B",X"C3",X"56",X"0B",X"E3",X"40",X"E2",X"3C",X"0B",X"C3",X"56",
		X"0B",X"E3",X"50",X"E2",X"3C",X"0B",X"C3",X"56",X"0B",X"11",X"2E",X"41",X"09",X"CB",X"36",X"3E",
		X"05",X"06",X"26",X"E5",X"EB",X"15",X"11",X"2E",X"45",X"09",X"3E",X"37",X"3E",X"05",X"06",X"26",
		X"E5",X"EB",X"15",X"AF",X"1A",X"4C",X"64",X"1A",X"6C",X"64",X"1A",X"5C",X"64",X"1A",X"7C",X"64",
		X"1A",X"84",X"64",X"11",X"E7",X"41",X"09",X"19",X"37",X"3E",X"01",X"06",X"05",X"E5",X"D5",X"15",
		X"11",X"91",X"41",X"09",X"1E",X"37",X"3E",X"01",X"06",X"20",X"E5",X"D5",X"15",X"3E",X"78",X"E5",
		X"B3",X"15",X"FD",X"E3",X"07",X"EE",X"E1",X"05",X"08",X"00",X"C8",X"58",X"42",X"21",X"00",X"05",
		X"08",X"00",X"D8",X"58",X"3E",X"21",X"00",X"05",X"08",X"00",X"F7",X"48",X"3A",X"21",X"00",X"05",
		X"08",X"00",X"EF",X"48",X"1E",X"21",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"08",X"00",X"02",X"58",X"2E",X"21",X"00",X"04",
		X"08",X"00",X"12",X"58",X"2A",X"21",X"00",X"04",X"08",X"00",X"01",X"48",X"0E",X"21",X"00",X"04",
		X"08",X"00",X"11",X"48",X"0A",X"21",X"00",X"04",X"08",X"00",X"FA",X"80",X"1A",X"21",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1E",X"00",X"FD",X"E3",X"07",X"AE",X"FD",X"1E",X"03",
		X"00",X"E1",X"14",X"10",X"24",X"26",X"30",X"30",X"30",X"30",X"30",X"34",X"30",X"34",X"30",X"34",
		X"30",X"34",X"30",X"34",X"30",X"34",X"30",X"34",X"30",X"34",X"FD",X"E3",X"07",X"5E",X"E0",X"FD",
		X"7E",X"00",X"FE",X"04",X"F2",X"7B",X"0F",X"F5",X"7E",X"03",X"FD",X"BE",X"03",X"F2",X"68",X"0F",
		X"E2",X"7B",X"0F",X"FD",X"7E",X"00",X"FE",X"05",X"E2",X"B2",X"0F",X"FD",X"7E",X"07",X"DE",X"37",
		X"CE",X"FB",X"FD",X"5F",X"07",X"F5",X"7E",X"03",X"FD",X"46",X"03",X"90",X"FE",X"05",X"38",X"05",
		X"FE",X"FB",X"18",X"01",X"E1",X"F5",X"7E",X"04",X"FD",X"46",X"04",X"90",X"FE",X"05",X"38",X"05",
		X"FE",X"FB",X"18",X"01",X"E1",X"F5",X"E3",X"07",X"EE",X"FD",X"E3",X"07",X"EE",X"E1",X"FD",X"7E",
		X"03",X"F5",X"BE",X"03",X"38",X"C5",X"30",X"07",X"FD",X"7E",X"00",X"FE",X"04",X"28",X"2B",X"FD",
		X"7E",X"07",X"DE",X"37",X"CE",X"FD",X"FD",X"5F",X"07",X"30",X"BA",X"F5",X"7E",X"04",X"FD",X"BE",
		X"04",X"38",X"09",X"E2",X"17",X"0F",X"FD",X"7E",X"00",X"FE",X"02",X"28",X"D1",X"FD",X"7E",X"07",
		X"DE",X"37",X"CE",X"DF",X"FD",X"5F",X"07",X"C3",X"1D",X"0F",X"FD",X"7E",X"04",X"F5",X"BE",X"04",
		X"38",X"EB",X"30",X"07",X"FD",X"7E",X"00",X"FE",X"03",X"28",X"9B",X"FD",X"7E",X"07",X"DE",X"37",
		X"CE",X"FE",X"FD",X"5F",X"07",X"C3",X"1D",X"0F",X"FD",X"7E",X"05",X"FE",X"30",X"28",X"05",X"FD",
		X"1E",X"05",X"30",X"E1",X"FD",X"1E",X"05",X"34",X"E1",X"3A",X"0D",X"66",X"3C",X"1A",X"0D",X"66",
		X"E3",X"7E",X"C0",X"2A",X"93",X"64",X"7E",X"09",X"27",X"28",X"E5",X"98",X"15",X"7E",X"1A",X"86",
		X"64",X"3A",X"A4",X"64",X"1A",X"84",X"64",X"3A",X"A5",X"64",X"1A",X"85",X"64",X"D5",X"0B",X"76",
		X"0B",X"56",X"2A",X"AE",X"64",X"31",X"0A",X"AE",X"64",X"D1",X"09",X"8F",X"65",X"E3",X"C6",X"AF",
		X"1A",X"0E",X"66",X"3A",X"0D",X"66",X"FE",X"10",X"C0",X"3E",X"FF",X"1A",X"0D",X"66",X"E1",X"44",
		X"00",X"10",X"60",X"00",X"08",X"64",X"00",X"40",X"50",X"00",X"80",X"D5",X"CD",X"2A",X"27",X"66",
		X"ED",X"73",X"AE",X"64",X"31",X"0A",X"AE",X"64",X"C9",X"D1",X"E1",X"F5",X"09",X"FC",X"2D",X"F5",
		X"0A",X"DE",X"65",X"09",X"6A",X"2F",X"3E",X"32",X"E5",X"C6",X"2B",X"E5",X"9F",X"18",X"3E",X"84",
		X"09",X"06",X"2B",X"E5",X"D5",X"2C",X"09",X"10",X"00",X"0A",X"11",X"66",X"3E",X"02",X"1A",X"13",
		X"66",X"3E",X"05",X"1A",X"14",X"66",X"3E",X"26",X"1A",X"29",X"66",X"09",X"F4",X"2C",X"E5",X"19",
		X"2C",X"E5",X"3A",X"2C",X"E1",X"F5",X"09",X"05",X"2E",X"F5",X"0A",X"DE",X"65",X"09",X"48",X"2E",
		X"3E",X"31",X"E5",X"C6",X"2B",X"E5",X"10",X"19",X"3E",X"87",X"09",X"0E",X"2B",X"E5",X"D5",X"2C",
		X"09",X"08",X"00",X"0A",X"11",X"66",X"3E",X"04",X"1A",X"13",X"66",X"3E",X"07",X"1A",X"14",X"66",
		X"3E",X"26",X"1A",X"29",X"66",X"09",X"24",X"2D",X"E5",X"19",X"2C",X"E5",X"3A",X"2C",X"E1",X"F5",
		X"09",X"05",X"2E",X"F5",X"0A",X"DE",X"65",X"09",X"DF",X"2E",X"3E",X"11",X"E5",X"C6",X"2B",X"E5",
		X"39",X"19",X"3E",X"6C",X"09",X"46",X"2B",X"E5",X"D5",X"2C",X"09",X"18",X"00",X"0A",X"11",X"66",
		X"3E",X"06",X"1A",X"13",X"66",X"3E",X"21",X"1A",X"14",X"66",X"3E",X"26",X"1A",X"29",X"66",X"09",
		X"3C",X"2D",X"E5",X"19",X"2C",X"E5",X"3A",X"2C",X"E1",X"F5",X"09",X"05",X"2E",X"F5",X"0A",X"DE",
		X"65",X"09",X"95",X"18",X"3E",X"26",X"E5",X"C6",X"2B",X"E5",X"86",X"19",X"3E",X"78",X"09",X"4E",
		X"2B",X"E5",X"D5",X"2C",X"09",X"40",X"00",X"0A",X"11",X"66",X"3E",X"20",X"1A",X"13",X"66",X"3E",
		X"24",X"1A",X"14",X"66",X"3E",X"27",X"1A",X"29",X"66",X"09",X"6C",X"2D",X"E5",X"19",X"2C",X"E5",
		X"3A",X"2C",X"E1",X"F5",X"09",X"05",X"2E",X"F5",X"0A",X"DE",X"65",X"09",X"1F",X"18",X"3E",X"37",
		X"E5",X"C6",X"2B",X"E5",X"95",X"19",X"3E",X"5A",X"09",X"86",X"2B",X"E5",X"D5",X"2C",X"09",X"50",
		X"00",X"0A",X"11",X"66",X"3E",X"20",X"1A",X"13",X"66",X"3E",X"24",X"1A",X"14",X"66",X"3E",X"27",
		X"1A",X"29",X"66",X"09",X"B4",X"2D",X"E5",X"19",X"2C",X"E5",X"3A",X"2C",X"E1",X"F5",X"09",X"FC",
		X"2D",X"F5",X"0A",X"DE",X"65",X"09",X"26",X"2E",X"3E",X"32",X"E5",X"C6",X"2B",X"E5",X"9E",X"19",
		X"3E",X"6F",X"09",X"8E",X"2B",X"E5",X"D5",X"2C",X"09",X"48",X"00",X"0A",X"11",X"66",X"3E",X"20",
		X"1A",X"13",X"66",X"3E",X"24",X"1A",X"14",X"66",X"3E",X"27",X"1A",X"29",X"66",X"09",X"E4",X"2D",
		X"E5",X"19",X"2C",X"E5",X"3A",X"2C",X"E1",X"F5",X"09",X"05",X"2E",X"F5",X"0A",X"DE",X"65",X"09",
		X"6A",X"2F",X"3E",X"31",X"E5",X"C6",X"2B",X"E5",X"9F",X"18",X"3E",X"81",X"09",X"06",X"2B",X"E5",
		X"D5",X"2C",X"09",X"58",X"00",X"0A",X"11",X"66",X"3E",X"20",X"1A",X"13",X"66",X"3E",X"24",X"1A",
		X"14",X"66",X"3E",X"27",X"1A",X"29",X"66",X"09",X"F4",X"2C",X"E5",X"19",X"2C",X"E5",X"3A",X"2C",
		X"E1",X"F5",X"09",X"05",X"2E",X"F5",X"0A",X"DE",X"65",X"09",X"48",X"2E",X"3E",X"11",X"E5",X"C6",
		X"2B",X"E5",X"10",X"19",X"3E",X"5D",X"09",X"0E",X"2B",X"E5",X"D5",X"2C",X"09",X"80",X"00",X"0A",
		X"11",X"66",X"3E",X"21",X"1A",X"13",X"66",X"3E",X"25",X"1A",X"14",X"66",X"3E",X"27",X"1A",X"29",
		X"66",X"09",X"24",X"2D",X"E5",X"19",X"2C",X"E5",X"3A",X"2C",X"E1",X"F5",X"09",X"05",X"2E",X"F5",
		X"0A",X"DE",X"65",X"09",X"DF",X"2E",X"3E",X"26",X"E5",X"C6",X"2B",X"E5",X"39",X"19",X"3E",X"69",
		X"09",X"46",X"2B",X"E5",X"D5",X"2C",X"09",X"90",X"00",X"0A",X"11",X"66",X"3E",X"21",X"1A",X"13",
		X"66",X"3E",X"25",X"1A",X"14",X"66",X"3E",X"27",X"1A",X"29",X"66",X"09",X"3C",X"2D",X"E5",X"19",
		X"2C",X"E5",X"3A",X"2C",X"E1",X"F5",X"09",X"05",X"2E",X"F5",X"0A",X"DE",X"65",X"09",X"95",X"18",
		X"3E",X"37",X"E5",X"C6",X"2B",X"E5",X"86",X"19",X"3E",X"7B",X"09",X"4E",X"2B",X"E5",X"D5",X"2C",
		X"09",X"00",X"01",X"0A",X"11",X"66",X"3E",X"22",X"1A",X"13",X"66",X"3E",X"26",X"1A",X"14",X"66",
		X"3E",X"27",X"1A",X"29",X"66",X"09",X"6C",X"2D",X"E5",X"19",X"2C",X"E5",X"3A",X"2C",X"E1",X"F5",
		X"09",X"FC",X"2D",X"F5",X"0A",X"DE",X"65",X"09",X"1F",X"18",X"3E",X"32",X"E5",X"C6",X"2B",X"E5",
		X"95",X"19",X"3E",X"7E",X"09",X"86",X"2B",X"E5",X"D5",X"2C",X"09",X"10",X"01",X"0A",X"11",X"66",
		X"3E",X"24",X"1A",X"13",X"66",X"3E",X"27",X"1A",X"14",X"66",X"3E",X"26",X"1A",X"29",X"66",X"09",
		X"B4",X"2D",X"E5",X"19",X"2C",X"E5",X"3A",X"2C",X"E1",X"F5",X"09",X"05",X"2E",X"F5",X"0A",X"DE",
		X"65",X"09",X"26",X"2E",X"3E",X"31",X"E5",X"C6",X"2B",X"E5",X"9E",X"19",X"3E",X"4E",X"09",X"8E",
		X"2B",X"E5",X"D5",X"2C",X"09",X"08",X"01",X"0A",X"11",X"66",X"3E",X"25",X"1A",X"13",X"66",X"3E",
		X"10",X"1A",X"14",X"66",X"3E",X"26",X"1A",X"29",X"66",X"09",X"E4",X"2D",X"E5",X"19",X"2C",X"E5",
		X"3A",X"2C",X"E1",X"E1",X"E1",X"E1",X"E1",X"27",X"65",X"52",X"08",X"54",X"66",X"54",X"2C",X"43",
		X"67",X"50",X"71",X"52",X"61",X"47",X"60",X"54",X"08",X"19",X"39",X"38",X"1B",X"54",X"45",X"64",
		X"63",X"67",X"08",X"61",X"66",X"43",X"8B",X"40",X"BC",X"40",X"A4",X"41",X"93",X"41",X"6C",X"42",
		X"5B",X"42",X"43",X"43",X"74",X"43",X"A3",X"40",X"94",X"40",X"8C",X"41",X"BB",X"41",X"44",X"42",
		X"73",X"42",X"6B",X"43",X"5C",X"43",X"AC",X"40",X"9B",X"40",X"29",X"41",X"1E",X"41",X"E1",X"42",
		X"D6",X"42",X"64",X"43",X"53",X"43",X"0B",X"41",X"3C",X"41",X"A5",X"41",X"92",X"41",X"6D",X"42",
		X"5A",X"42",X"C3",X"42",X"F4",X"42",X"E5",X"40",X"D2",X"40",X"46",X"41",X"71",X"41",X"8E",X"42",
		X"B9",X"42",X"2D",X"43",X"1A",X"43",X"8B",X"40",X"BC",X"40",X"A2",X"41",X"95",X"41",X"6A",X"42",
		X"5D",X"42",X"43",X"43",X"74",X"43",X"AB",X"40",X"9C",X"40",X"2C",X"41",X"1B",X"41",X"E4",X"42",
		X"D3",X"42",X"63",X"43",X"54",X"43",X"E5",X"41",X"D2",X"41",X"A0",X"41",X"97",X"41",X"68",X"42",
		X"5F",X"42",X"2D",X"42",X"1A",X"42",X"C5",X"40",X"F2",X"40",X"A3",X"41",X"94",X"41",X"6B",X"42",
		X"5C",X"42",X"0D",X"43",X"3A",X"43",X"EC",X"40",X"DB",X"40",X"28",X"41",X"1F",X"41",X"E0",X"42",
		X"D7",X"42",X"24",X"43",X"13",X"43",X"C4",X"40",X"F3",X"40",X"2C",X"41",X"1B",X"41",X"E4",X"42",
		X"D3",X"42",X"0C",X"43",X"3B",X"43",X"A1",X"40",X"96",X"40",X"A8",X"41",X"9F",X"41",X"60",X"42",
		X"57",X"42",X"69",X"43",X"5E",X"43",X"CD",X"E5",X"25",X"15",X"11",X"40",X"40",X"C9",X"D5",X"11",
		X"F7",X"65",X"ED",X"88",X"ED",X"88",X"ED",X"88",X"7E",X"FE",X"27",X"38",X"DD",X"ED",X"88",X"2B",
		X"D1",X"CD",X"09",X"F7",X"65",X"0B",X"46",X"F5",X"7E",X"00",X"12",X"13",X"10",X"FC",X"7E",X"0B",
		X"86",X"2B",X"5F",X"0B",X"0B",X"7E",X"FE",X"D8",X"18",X"30",X"12",X"13",X"0B",X"46",X"F5",X"7E",
		X"01",X"12",X"13",X"10",X"FC",X"7E",X"0B",X"86",X"2B",X"5F",X"0B",X"0B",X"7E",X"12",X"13",X"C3",
		X"CD",X"2B",X"09",X"F7",X"65",X"3A",X"DD",X"65",X"3C",X"1A",X"DD",X"65",X"FE",X"34",X"28",X"23",
		X"7E",X"3D",X"5F",X"FE",X"D9",X"D2",X"CD",X"2B",X"C3",X"E5",X"2B",X"C9",X"AF",X"1A",X"DD",X"65",
		X"E1",X"11",X"49",X"64",X"01",X"18",X"00",X"ED",X"98",X"E1",X"09",X"F8",X"65",X"11",X"F9",X"65",
		X"1E",X"00",X"01",X"11",X"00",X"ED",X"98",X"09",X"FB",X"65",X"E3",X"FE",X"09",X"FE",X"65",X"E3",
		X"FE",X"09",X"01",X"66",X"E3",X"FE",X"09",X"04",X"66",X"E3",X"FE",X"09",X"07",X"66",X"E3",X"FE",
		X"AF",X"1A",X"33",X"66",X"1A",X"0D",X"66",X"1A",X"0E",X"66",X"1A",X"2A",X"66",X"1A",X"2B",X"66",
		X"3A",X"04",X"65",X"17",X"09",X"B5",X"2C",X"E5",X"98",X"15",X"7E",X"1A",X"18",X"40",X"0B",X"7E",
		X"1A",X"2F",X"40",X"3E",X"01",X"1A",X"18",X"44",X"1A",X"2F",X"44",X"3E",X"40",X"1A",X"0B",X"66",
		X"1A",X"0C",X"66",X"09",X"F5",X"65",X"E3",X"86",X"AF",X"1A",X"C2",X"66",X"E1",X"40",X"01",X"40",
		X"02",X"40",X"03",X"40",X"04",X"40",X"05",X"40",X"06",X"40",X"07",X"40",X"20",X"40",X"21",X"01",
		X"00",X"01",X"01",X"01",X"02",X"01",X"03",X"01",X"04",X"01",X"05",X"01",X"06",X"01",X"07",X"01",
		X"20",X"01",X"21",X"02",X"00",X"02",X"01",X"02",X"02",X"02",X"03",X"02",X"04",X"02",X"05",X"02",
		X"06",X"02",X"07",X"02",X"20",X"1A",X"2C",X"66",X"0A",X"0F",X"66",X"E1",X"03",X"02",X"00",X"3B",
		X"14",X"30",X"21",X"77",X"03",X"02",X"00",X"4B",X"14",X"30",X"21",X"37",X"03",X"02",X"00",X"AB",
		X"14",X"30",X"21",X"37",X"03",X"02",X"00",X"D3",X"14",X"30",X"21",X"37",X"00",X"00",X"00",X"00",
		X"00",X"00",X"21",X"00",X"02",X"04",X"00",X"A3",X"CC",X"10",X"21",X"40",X"03",X"02",X"00",X"4B",
		X"14",X"30",X"21",X"77",X"03",X"02",X"00",X"7B",X"14",X"30",X"21",X"37",X"03",X"02",X"00",X"93",
		X"14",X"30",X"21",X"37",X"03",X"02",X"00",X"AB",X"14",X"30",X"21",X"37",X"00",X"00",X"00",X"00",
		X"00",X"00",X"21",X"00",X"02",X"04",X"00",X"A3",X"FC",X"10",X"21",X"40",X"03",X"02",X"00",X"63",
		X"0C",X"30",X"21",X"77",X"03",X"02",X"00",X"5B",X"0C",X"30",X"21",X"37",X"03",X"02",X"00",X"B3",
		X"0C",X"30",X"21",X"37",X"03",X"02",X"00",X"C3",X"0C",X"30",X"21",X"37",X"00",X"00",X"00",X"00",
		X"00",X"00",X"21",X"00",X"02",X"04",X"00",X"A3",X"EC",X"10",X"21",X"40",X"03",X"02",X"00",X"43",
		X"44",X"30",X"21",X"77",X"03",X"02",X"00",X"53",X"1C",X"30",X"21",X"37",X"03",X"02",X"00",X"BB",
		X"1C",X"30",X"21",X"37",X"03",X"02",X"00",X"E3",X"44",X"30",X"21",X"37",X"00",X"00",X"00",X"00",
		X"00",X"00",X"21",X"00",X"02",X"04",X"00",X"A3",X"FC",X"10",X"21",X"40",X"03",X"02",X"00",X"73",
		X"2C",X"30",X"21",X"77",X"03",X"02",X"00",X"5B",X"2C",X"30",X"21",X"37",X"03",X"02",X"00",X"B3",
		X"2C",X"30",X"21",X"37",X"03",X"02",X"00",X"9B",X"2C",X"30",X"21",X"37",X"00",X"00",X"00",X"00",
		X"00",X"00",X"21",X"00",X"02",X"04",X"00",X"A3",X"CC",X"10",X"21",X"40",X"03",X"02",X"00",X"43",
		X"14",X"30",X"21",X"77",X"03",X"02",X"00",X"73",X"14",X"30",X"21",X"37",X"03",X"02",X"00",X"9B",
		X"14",X"30",X"21",X"37",X"03",X"02",X"00",X"E3",X"14",X"30",X"21",X"37",X"00",X"00",X"00",X"00",
		X"00",X"00",X"21",X"00",X"02",X"04",X"00",X"A3",X"F4",X"10",X"21",X"40",X"4D",X"22",X"23",X"24",
		X"25",X"26",X"27",X"10",X"14",X"4D",X"22",X"23",X"24",X"25",X"26",X"27",X"10",X"16",X"D9",X"08",
		X"00",X"DC",X"04",X"FF",X"23",X"06",X"02",X"25",X"20",X"FE",X"23",X"06",X"02",X"25",X"04",X"FF",
		X"DC",X"01",X"00",X"22",X"34",X"00",X"22",X"01",X"00",X"DC",X"01",X"01",X"24",X"34",X"FE",X"26",
		X"01",X"01",X"DA",X"05",X"00",X"22",X"14",X"00",X"22",X"05",X"00",X"DC",X"04",X"FF",X"23",X"16",
		X"02",X"25",X"04",X"FF",X"DC",X"01",X"00",X"22",X"34",X"00",X"22",X"01",X"00",X"DC",X"01",X"01",
		X"24",X"24",X"FE",X"26",X"02",X"02",X"24",X"24",X"FE",X"26",X"01",X"01",X"D9",X"08",X"00",X"FF",
		X"D9",X"08",X"00",X"DB",X"07",X"01",X"24",X"10",X"FE",X"26",X"07",X"01",X"D9",X"22",X"00",X"22",
		X"22",X"00",X"22",X"22",X"00",X"D9",X"21",X"00",X"23",X"24",X"00",X"25",X"21",X"00",X"DA",X"01",
		X"00",X"22",X"02",X"01",X"25",X"03",X"FE",X"23",X"26",X"02",X"25",X"03",X"FE",X"23",X"02",X"01",
		X"22",X"01",X"00",X"DC",X"01",X"00",X"22",X"34",X"00",X"22",X"01",X"00",X"DA",X"01",X"00",X"22",
		X"24",X"FF",X"26",X"02",X"02",X"24",X"24",X"FF",X"22",X"01",X"00",X"DA",X"01",X"00",X"22",X"23",
		X"01",X"25",X"04",X"FE",X"23",X"23",X"01",X"22",X"01",X"00",X"DC",X"01",X"00",X"22",X"34",X"00",
		X"22",X"01",X"00",X"DA",X"01",X"00",X"22",X"03",X"FF",X"26",X"01",X"02",X"24",X"10",X"FE",X"26",
		X"01",X"02",X"24",X"03",X"FF",X"22",X"01",X"00",X"D9",X"21",X"00",X"24",X"24",X"00",X"26",X"21",
		X"00",X"D9",X"22",X"00",X"22",X"22",X"00",X"22",X"22",X"00",X"DB",X"21",X"FF",X"23",X"24",X"02",
		X"25",X"21",X"FF",X"D9",X"08",X"00",X"FF",X"D9",X"08",X"00",X"DC",X"01",X"00",X"22",X"02",X"01",
		X"25",X"20",X"FE",X"23",X"04",X"02",X"25",X"20",X"FE",X"23",X"02",X"01",X"22",X"01",X"00",X"D9",
		X"02",X"00",X"24",X"32",X"00",X"26",X"02",X"00",X"DD",X"03",X"00",X"22",X"30",X"00",X"22",X"03",
		X"00",X"DB",X"03",X"00",X"22",X"22",X"FF",X"26",X"02",X"02",X"24",X"22",X"FF",X"22",X"03",X"00",
		X"DB",X"03",X"00",X"22",X"20",X"01",X"25",X"06",X"FE",X"23",X"20",X"01",X"22",X"03",X"00",X"DD",
		X"03",X"00",X"22",X"30",X"00",X"22",X"03",X"00",X"D9",X"02",X"00",X"23",X"32",X"00",X"25",X"02",
		X"00",X"DC",X"01",X"00",X"22",X"05",X"FF",X"26",X"02",X"02",X"24",X"22",X"FE",X"26",X"02",X"02",
		X"24",X"05",X"FF",X"22",X"01",X"00",X"D9",X"08",X"00",X"FF",X"D9",X"08",X"00",X"DB",X"03",X"FF",
		X"23",X"20",X"02",X"25",X"06",X"FE",X"23",X"20",X"02",X"25",X"03",X"FF",X"D9",X"01",X"00",X"22",
		X"34",X"00",X"22",X"01",X"00",X"DA",X"01",X"00",X"22",X"04",X"FF",X"26",X"02",X"02",X"24",X"24",
		X"FE",X"26",X"02",X"02",X"24",X"04",X"FF",X"22",X"01",X"00",X"DA",X"01",X"00",X"22",X"03",X"01",
		X"25",X"04",X"FE",X"23",X"22",X"02",X"25",X"04",X"FE",X"23",X"03",X"01",X"22",X"01",X"00",X"D9",
		X"01",X"00",X"22",X"34",X"00",X"22",X"01",X"00",X"DA",X"01",X"01",X"24",X"34",X"FE",X"26",X"01",
		X"01",X"DA",X"03",X"01",X"24",X"22",X"FE",X"26",X"02",X"02",X"24",X"22",X"FE",X"26",X"03",X"01",
		X"DA",X"04",X"FF",X"23",X"20",X"02",X"25",X"04",X"FE",X"23",X"20",X"02",X"25",X"04",X"FF",X"DA",
		X"02",X"FF",X"23",X"32",X"02",X"25",X"02",X"FF",X"D9",X"01",X"00",X"22",X"34",X"00",X"22",X"01",
		X"00",X"DA",X"01",X"00",X"22",X"04",X"FF",X"26",X"02",X"02",X"24",X"24",X"FE",X"26",X"02",X"02",
		X"24",X"04",X"FF",X"22",X"01",X"00",X"DA",X"01",X"00",X"22",X"03",X"01",X"25",X"04",X"FE",X"23",
		X"22",X"02",X"25",X"04",X"FE",X"23",X"03",X"01",X"22",X"01",X"00",X"D9",X"01",X"00",X"22",X"34",
		X"00",X"22",X"01",X"00",X"DB",X"01",X"01",X"24",X"24",X"FE",X"26",X"02",X"02",X"24",X"24",X"FE",
		X"26",X"01",X"01",X"D9",X"08",X"00",X"FF",X"D9",X"08",X"00",X"DB",X"05",X"FF",X"23",X"01",X"02",
		X"25",X"06",X"FE",X"23",X"02",X"02",X"25",X"06",X"FE",X"23",X"01",X"02",X"25",X"05",X"FF",X"D9",
		X"02",X"00",X"23",X"32",X"00",X"25",X"02",X"00",X"DB",X"01",X"01",X"24",X"34",X"FE",X"26",X"01",
		X"01",X"FC",X"04",X"00",X"22",X"16",X"00",X"22",X"04",X"00",X"DB",X"03",X"FF",X"23",X"30",X"02",
		X"25",X"03",X"FF",X"D9",X"02",X"00",X"24",X"32",X"00",X"26",X"02",X"00",X"DB",X"03",X"01",X"24",
		X"05",X"FE",X"26",X"02",X"02",X"24",X"06",X"FE",X"26",X"02",X"02",X"24",X"05",X"FE",X"26",X"03",
		X"01",X"D9",X"08",X"00",X"FF",X"D9",X"08",X"00",X"FB",X"23",X"FF",X"23",X"20",X"02",X"25",X"23",
		X"FF",X"DC",X"01",X"00",X"22",X"34",X"00",X"22",X"01",X"00",X"FB",X"01",X"01",X"24",X"34",X"FE",
		X"26",X"01",X"01",X"D9",X"08",X"00",X"FF",X"3E",X"26",X"1A",X"C7",X"40",X"1A",X"D7",X"40",X"1A",
		X"AF",X"41",X"1A",X"87",X"42",X"1A",X"97",X"42",X"1A",X"2F",X"43",X"3E",X"24",X"1A",X"E0",X"40",
		X"1A",X"F0",X"40",X"1A",X"98",X"41",X"1A",X"A0",X"42",X"1A",X"B0",X"42",X"1A",X"18",X"43",X"3E",
		X"25",X"1A",X"E7",X"40",X"1A",X"4F",X"41",X"1A",X"5F",X"41",X"1A",X"67",X"42",X"1A",X"0F",X"43",
		X"1A",X"1F",X"43",X"3E",X"23",X"1A",X"D0",X"40",X"1A",X"68",X"41",X"1A",X"78",X"41",X"1A",X"50",
		X"42",X"1A",X"28",X"43",X"1A",X"38",X"43",X"3E",X"22",X"1A",X"FB",X"41",X"1A",X"33",X"42",X"E1",
		X"3E",X"26",X"1A",X"AF",X"41",X"3E",X"24",X"1A",X"98",X"41",X"3E",X"25",X"1A",X"67",X"42",X"3E",
		X"23",X"1A",X"50",X"42",X"3E",X"24",X"1A",X"C9",X"42",X"3E",X"23",X"1A",X"01",X"41",X"3E",X"25",
		X"1A",X"36",X"41",X"3E",X"26",X"1A",X"FE",X"42",X"E1",X"3E",X"25",X"1A",X"E8",X"40",X"1A",X"DE",
		X"40",X"1A",X"6F",X"42",X"3E",X"23",X"1A",X"E9",X"40",X"1A",X"DF",X"40",X"1A",X"58",X"42",X"3E",
		X"26",X"1A",X"A7",X"41",X"1A",X"20",X"43",X"1A",X"16",X"43",X"3E",X"24",X"1A",X"90",X"41",X"1A",
		X"21",X"43",X"1A",X"17",X"43",X"3E",X"24",X"1A",X"81",X"43",X"1A",X"C1",X"40",X"3E",X"23",X"1A",
		X"09",X"43",X"1A",X"49",X"40",X"3E",X"26",X"1A",X"B6",X"43",X"1A",X"F6",X"40",X"3E",X"25",X"1A",
		X"3E",X"43",X"1A",X"7E",X"40",X"E1",X"3E",X"22",X"1A",X"0D",X"41",X"1A",X"CF",X"40",X"1A",X"C5",
		X"42",X"1A",X"07",X"43",X"E1",X"3E",X"25",X"1A",X"E2",X"40",X"1A",X"D4",X"40",X"3E",X"23",X"1A",
		X"E3",X"40",X"1A",X"D5",X"40",X"3E",X"26",X"1A",X"2A",X"43",X"1A",X"1C",X"43",X"3E",X"24",X"1A",
		X"2B",X"43",X"1A",X"1D",X"43",X"E1",X"3E",X"25",X"1A",X"EF",X"40",X"3E",X"23",X"1A",X"D8",X"40",
		X"1A",X"05",X"42",X"3E",X"24",X"1A",X"CD",X"41",X"1A",X"10",X"43",X"3E",X"26",X"1A",X"27",X"43",
		X"E1",X"3E",X"16",X"E5",X"FD",X"14",X"3E",X"21",X"E5",X"25",X"15",X"11",X"C1",X"44",X"09",X"03",
		X"1C",X"3E",X"05",X"06",X"15",X"E5",X"EB",X"15",X"11",X"7B",X"44",X"09",X"03",X"1C",X"3E",X"05",
		X"06",X"10",X"E5",X"EB",X"15",X"11",X"C1",X"40",X"09",X"39",X"1A",X"3E",X"05",X"06",X"15",X"E5",
		X"D5",X"15",X"11",X"61",X"41",X"09",X"8A",X"1A",X"3E",X"07",X"06",X"11",X"E5",X"D5",X"15",X"3E",
		X"90",X"1A",X"EE",X"40",X"3E",X"A6",X"1A",X"EF",X"40",X"11",X"9A",X"40",X"09",X"31",X"1B",X"3E",
		X"07",X"06",X"16",X"E5",X"D5",X"15",X"11",X"7B",X"40",X"09",X"9B",X"1B",X"3E",X"05",X"06",X"10",
		X"E5",X"D5",X"15",X"3E",X"78",X"E5",X"B3",X"15",X"E1",X"31",X"31",X"31",X"31",X"31",X"31",X"40",
		X"40",X"40",X"31",X"31",X"40",X"53",X"40",X"31",X"31",X"40",X"54",X"40",X"31",X"31",X"40",X"66",
		X"40",X"31",X"31",X"40",X"45",X"40",X"31",X"31",X"40",X"53",X"40",X"31",X"31",X"40",X"45",X"40",
		X"31",X"31",X"40",X"52",X"40",X"31",X"31",X"40",X"50",X"40",X"31",X"31",X"40",X"40",X"40",X"31",
		X"31",X"40",X"40",X"40",X"31",X"31",X"40",X"72",X"40",X"31",X"31",X"40",X"45",X"40",X"31",X"31",
		X"40",X"60",X"40",X"31",X"31",X"40",X"43",X"40",X"31",X"31",X"40",X"66",X"40",X"31",X"31",X"40",
		X"41",X"40",X"31",X"31",X"40",X"53",X"40",X"31",X"31",X"40",X"40",X"40",X"31",X"31",X"31",X"31",
		X"31",X"31",X"16",X"16",X"A5",X"16",X"A2",X"A3",X"A6",X"A3",X"A3",X"A7",X"A4",X"A3",X"A7",X"A6",
		X"A7",X"16",X"16",X"A7",X"16",X"A7",X"A6",X"A7",X"16",X"16",X"A7",X"16",X"16",X"16",X"A7",X"A5",
		X"A5",X"A7",X"A5",X"A5",X"16",X"A7",X"A7",X"A7",X"A7",X"A7",X"A7",X"A6",X"A7",X"16",X"16",X"16",
		X"16",X"A7",X"A6",X"16",X"16",X"16",X"16",X"16",X"A7",X"A6",X"16",X"16",X"16",X"16",X"16",X"16",
		X"16",X"A5",X"16",X"A5",X"A5",X"A5",X"A5",X"16",X"A7",X"A3",X"A7",X"A7",X"A7",X"A7",X"A6",X"A7",
		X"A4",X"16",X"16",X"16",X"A7",X"A6",X"16",X"90",X"A4",X"16",X"16",X"16",X"16",X"16",X"A3",X"91",
		X"16",X"16",X"16",X"16",X"A7",X"91",X"16",X"A5",X"A5",X"A5",X"16",X"A7",X"90",X"A7",X"A7",X"A7",
		X"A7",X"A6",X"16",X"16",X"16",X"16",X"16",X"A7",X"A6",X"A5",X"A5",X"16",X"16",X"16",X"16",X"16",
		X"A7",X"91",X"16",X"16",X"16",X"16",X"16",X"A7",X"A6",X"16",X"A5",X"A5",X"A5",X"16",X"A7",X"A7",
		X"A7",X"A7",X"A7",X"A7",X"A6",X"A7",X"A6",X"16",X"16",X"16",X"16",X"16",X"A7",X"A4",X"16",X"16",
		X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"A5",X"A5",X"A5",X"A5",
		X"16",X"A7",X"90",X"A7",X"A7",X"A7",X"A7",X"A6",X"A7",X"16",X"16",X"A3",X"91",X"16",X"16",X"16",
		X"16",X"A3",X"91",X"A2",X"16",X"16",X"16",X"A3",X"91",X"A2",X"16",X"16",X"16",X"A7",X"91",X"16",
		X"A5",X"A5",X"A5",X"16",X"A7",X"90",X"A7",X"A7",X"A7",X"A7",X"A6",X"16",X"16",X"16",X"16",X"16",
		X"A7",X"A6",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"A5",X"A5",X"16",X"16",X"16",X"16",X"16",
		X"A7",X"91",X"16",X"16",X"16",X"16",X"16",X"A7",X"A6",X"16",X"A5",X"A5",X"A5",X"16",X"A7",X"A7",
		X"A7",X"A7",X"A7",X"A7",X"A6",X"A7",X"A6",X"16",X"16",X"16",X"16",X"16",X"A7",X"A4",X"16",X"16",
		X"16",X"16",X"16",X"31",X"31",X"31",X"31",X"31",X"31",X"40",X"40",X"40",X"31",X"31",X"40",X"67",
		X"40",X"31",X"31",X"40",X"63",X"40",X"31",X"31",X"40",X"64",X"40",X"31",X"31",X"40",X"45",X"40",
		X"31",X"31",X"40",X"54",X"40",X"31",X"31",X"40",X"40",X"40",X"31",X"31",X"40",X"03",X"40",X"31",
		X"31",X"40",X"20",X"40",X"31",X"31",X"40",X"21",X"40",X"31",X"31",X"40",X"01",X"40",X"31",X"31",
		X"40",X"40",X"40",X"31",X"31",X"40",X"32",X"40",X"31",X"31",X"40",X"40",X"40",X"31",X"31",X"31",
		X"31",X"31",X"31",X"05",X"E1",X"E1",X"E1",X"09",X"CC",X"1C",X"0A",X"2D",X"66",X"3E",X"EF",X"1A",
		X"F8",X"64",X"E1",X"E1",X"2A",X"2D",X"66",X"CD",X"09",X"CC",X"1C",X"7D",X"C9",X"BD",X"E4",X"64",
		X"1C",X"7E",X"FE",X"00",X"28",X"26",X"0B",X"46",X"3A",X"A4",X"64",X"B8",X"28",X"14",X"2B",X"0A",
		X"2D",X"66",X"30",X"17",X"0B",X"46",X"3A",X"A5",X"64",X"B8",X"28",X"06",X"2B",X"0A",X"2D",X"66",
		X"30",X"21",X"0B",X"7E",X"1A",X"F8",X"64",X"0B",X"0A",X"2D",X"66",X"E1",X"3E",X"10",X"1A",X"29",
		X"66",X"3E",X"04",X"1A",X"13",X"66",X"3E",X"22",X"1A",X"14",X"66",X"3E",X"07",X"1A",X"4A",X"64",
		X"1A",X"6A",X"64",X"1A",X"5A",X"64",X"1A",X"7A",X"64",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",
		X"E1",X"E1",X"3E",X"40",X"E5",X"FD",X"14",X"3E",X"21",X"E5",X"25",X"15",X"3E",X"31",X"1A",X"34",
		X"66",X"E5",X"92",X"1C",X"3E",X"27",X"E5",X"B3",X"15",X"3E",X"14",X"1A",X"34",X"66",X"E5",X"92",
		X"1C",X"E1",X"09",X"40",X"40",X"0A",X"35",X"66",X"09",X"7F",X"40",X"0A",X"37",X"66",X"3E",X"08",
		X"1A",X"09",X"66",X"E5",X"9D",X"1C",X"3E",X"01",X"E5",X"B3",X"15",X"3A",X"09",X"66",X"3D",X"1A",
		X"09",X"66",X"08",X"EF",X"E1",X"06",X"26",X"ED",X"73",X"35",X"66",X"13",X"ED",X"53",X"35",X"66",
		X"33",X"3A",X"34",X"66",X"12",X"3E",X"40",X"E5",X"9D",X"15",X"10",X"DD",X"06",X"26",X"ED",X"73",
		X"37",X"66",X"33",X"ED",X"53",X"37",X"66",X"13",X"3A",X"34",X"66",X"12",X"3E",X"40",X"E5",X"9D",
		X"15",X"10",X"DD",X"E1",X"00",X"CC",X"FB",X"01",X"B3",X"DF",X"00",X"EC",X"FB",X"01",X"CB",X"FE",
		X"00",X"B4",X"FD",X"01",X"E3",X"FE",X"00",X"4C",X"FB",X"01",X"CB",X"FE",X"00",X"0C",X"FD",X"01",
		X"B3",X"DF",X"00",X"84",X"FB",X"01",X"D3",X"FE",X"00",X"74",X"FD",X"01",X"C3",X"DF",X"00",X"9C",
		X"FB",X"01",X"EB",X"DF",X"00",X"EC",X"FD",X"01",X"CB",X"DF",X"00",X"DC",X"FD",X"01",X"B3",X"FE",
		X"00",X"EC",X"FD",X"01",X"93",X"FE",X"00",X"8C",X"FD",X"01",X"0B",X"DF",X"00",X"EC",X"FB",X"01",
		X"5B",X"FE",X"00",X"A4",X"FD",X"01",X"43",X"FE",X"00",X"4C",X"FD",X"01",X"2B",X"FE",X"00",X"34",
		X"FB",X"01",X"5B",X"DF",X"00",X"74",X"FB",X"01",X"BB",X"DF",X"00",X"A4",X"FB",X"01",X"D3",X"DF",
		X"00",X"C4",X"FB",X"01",X"F3",X"DF",X"00",X"FC",X"FD",X"01",X"AB",X"FE",X"00",X"E4",X"FD",X"01",
		X"7B",X"DF",X"00",X"EC",X"FD",X"01",X"5B",X"DF",X"00",X"DC",X"FD",X"01",X"2B",X"FE",X"00",X"B4",
		X"FB",X"01",X"83",X"DF",X"23",X"08",X"65",X"23",X"3B",X"65",X"24",X"02",X"01",X"43",X"00",X"02",
		X"20",X"05",X"04",X"01",X"54",X"00",X"05",X"04",X"01",X"1A",X"00",X"05",X"04",X"01",X"85",X"00",
		X"05",X"04",X"01",X"8F",X"00",X"05",X"04",X"01",X"4C",X"00",X"05",X"04",X"01",X"23",X"01",X"05",
		X"04",X"21",X"23",X"05",X"65",X"23",X"3B",X"65",X"01",X"D8",X"00",X"24",X"02",X"06",X"02",X"20",
		X"05",X"03",X"02",X"00",X"05",X"03",X"07",X"27",X"21",X"23",X"05",X"65",X"24",X"02",X"01",X"00",
		X"02",X"02",X"05",X"06",X"04",X"05",X"06",X"05",X"01",X"04",X"FF",X"07",X"06",X"07",X"04",X"21",
		X"AE",X"64",X"F8",X"2E",X"46",X"53",X"43",X"67",X"52",X"45",X"08",X"08",X"05",X"00",X"95",X"2B",
		X"A8",X"2B",X"98",X"64",X"DA",X"1C",X"46",X"65",X"45",X"66",X"52",X"23",X"3B",X"65",X"23",X"59",
		X"65",X"23",X"A4",X"65",X"23",X"8F",X"65",X"24",X"02",X"01",X"08",X"00",X"02",X"27",X"06",X"05",
		X"01",X"03",X"18",X"00",X"07",X"14",X"06",X"04",X"FF",X"05",X"04",X"07",X"07",X"01",X"99",X"00",
		X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"04",X"05",X"04",X"01",X"85",X"00",X"02",X"26",
		X"06",X"04",X"FE",X"05",X"02",X"07",X"04",X"05",X"04",X"01",X"7D",X"00",X"02",X"26",X"06",X"04",
		X"FE",X"05",X"02",X"07",X"04",X"05",X"04",X"01",X"5E",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",
		X"02",X"07",X"02",X"05",X"01",X"01",X"69",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",
		X"04",X"05",X"02",X"01",X"70",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"02",X"05",
		X"01",X"01",X"69",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"02",X"05",X"02",X"01",
		X"4C",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"02",X"05",X"01",X"01",X"69",X"00",
		X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"02",X"05",X"02",X"01",X"70",X"00",X"02",X"26",
		X"06",X"04",X"FE",X"05",X"02",X"07",X"06",X"21",X"24",X"01",X"02",X"01",X"06",X"01",X"80",X"00",
		X"06",X"05",X"02",X"03",X"10",X"00",X"07",X"05",X"04",X"02",X"07",X"06",X"20",X"B0",X"1E",X"52",
		X"41",X"65",X"1D",X"08",X"05",X"00",X"95",X"2B",X"A8",X"2B",X"8F",X"65",X"C6",X"1E",X"53",X"67",
		X"55",X"52",X"41",X"65",X"1E",X"08",X"05",X"00",X"95",X"2B",X"24",X"02",X"01",X"99",X"00",X"02",
		X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"02",X"05",X"02",X"01",X"99",X"00",X"02",X"26",X"06",
		X"04",X"FE",X"05",X"02",X"07",X"02",X"05",X"01",X"01",X"99",X"00",X"02",X"26",X"06",X"04",X"FE",
		X"05",X"02",X"07",X"02",X"05",X"01",X"01",X"99",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",
		X"07",X"02",X"05",X"01",X"01",X"99",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"02",
		X"05",X"01",X"01",X"85",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"02",X"05",X"02",
		X"01",X"99",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"02",X"05",X"02",X"01",X"C8",
		X"00",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"02",X"05",X"02",X"01",X"C8",X"00",X"02",
		X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"02",X"05",X"01",X"01",X"C8",X"00",X"02",X"26",X"06",
		X"04",X"FE",X"05",X"02",X"07",X"02",X"05",X"01",X"01",X"C8",X"00",X"02",X"26",X"06",X"04",X"FE",
		X"05",X"02",X"07",X"02",X"05",X"01",X"01",X"C8",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",
		X"07",X"02",X"05",X"01",X"01",X"99",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"02",
		X"05",X"02",X"01",X"C8",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"02",X"05",X"02",
		X"01",X"23",X"01",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"02",X"05",X"02",X"01",X"23",
		X"01",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"02",X"05",X"01",X"01",X"23",X"01",X"02",
		X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"02",X"05",X"01",X"01",X"23",X"01",X"02",X"26",X"06",
		X"04",X"FE",X"05",X"02",X"07",X"02",X"05",X"01",X"01",X"23",X"01",X"02",X"26",X"06",X"04",X"FE",
		X"05",X"02",X"07",X"02",X"05",X"01",X"01",X"C8",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",
		X"07",X"02",X"05",X"02",X"01",X"23",X"01",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"03",
		X"01",X"4C",X"01",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"02",X"06",X"05",X"07",X"04",
		X"FE",X"07",X"04",X"21",X"24",X"01",X"02",X"27",X"06",X"01",X"C0",X"00",X"06",X"05",X"01",X"03",
		X"10",X"00",X"07",X"05",X"04",X"FE",X"07",X"06",X"21",X"23",X"8F",X"65",X"24",X"02",X"01",X"43",
		X"00",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"04",X"05",X"01",X"01",X"70",X"00",X"02",
		X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"04",X"05",X"02",X"01",X"58",X"00",X"02",X"26",X"06",
		X"04",X"FE",X"05",X"02",X"07",X"02",X"01",X"85",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",
		X"07",X"02",X"05",X"01",X"01",X"58",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"04",
		X"01",X"5E",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"04",X"05",X"02",X"01",X"95",
		X"00",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"02",X"01",X"99",X"00",X"02",X"26",X"06",
		X"04",X"FE",X"05",X"02",X"07",X"02",X"05",X"01",X"01",X"95",X"00",X"02",X"26",X"06",X"04",X"FE",
		X"05",X"02",X"07",X"04",X"01",X"85",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"04",
		X"05",X"02",X"01",X"8F",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"02",X"01",X"C7",
		X"00",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"02",X"05",X"01",X"01",X"8F",X"00",X"02",
		X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"04",X"01",X"99",X"00",X"02",X"26",X"06",X"04",X"FE",
		X"05",X"02",X"07",X"02",X"01",X"99",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"02",
		X"01",X"95",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"04",X"01",X"99",X"00",X"02",
		X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"06",X"05",X"02",X"01",X"85",X"00",X"02",X"26",X"06",
		X"04",X"FE",X"05",X"02",X"07",X"04",X"05",X"03",X"01",X"99",X"00",X"02",X"26",X"06",X"04",X"FE",
		X"05",X"02",X"07",X"02",X"01",X"99",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"02",
		X"01",X"99",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"02",X"01",X"A5",X"00",X"02",
		X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"02",X"01",X"95",X"00",X"02",X"26",X"06",X"04",X"FE",
		X"05",X"02",X"07",X"02",X"05",X"01",X"01",X"5E",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",
		X"07",X"06",X"05",X"04",X"01",X"EC",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"06",
		X"21",X"00",X"00",X"15",X"00",X"00",X"00",X"18",X"00",X"00",X"00",X"45",X"00",X"00",X"00",X"48",
		X"00",X"00",X"50",X"12",X"00",X"00",X"00",X"0D",X"00",X"00",X"50",X"1F",X"00",X"00",X"00",X"50",
		X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"18",X"00",X"00",X"00",X"40",
		X"00",X"00",X"50",X"07",X"00",X"00",X"00",X"15",X"00",X"00",X"50",X"0A",X"00",X"00",X"00",X"18",
		X"00",X"05",X"04",X"03",X"02",X"00",X"03",X"06",X"21",X"00",X"03",X"00",X"00",X"06",X"03",X"00",
		X"03",X"00",X"00",X"06",X"03",X"00",X"00",X"21",X"00",X"FF",X"64",X"52",X"53",X"50",X"42",X"03",
		X"65",X"43",X"53",X"48",X"17",X"03",X"62",X"65",X"53",X"08",X"85",X"02",X"42",X"67",X"40",X"90",
		X"5E",X"02",X"62",X"53",X"40",X"50",X"19",X"02",X"62",X"46",X"53",X"90",X"10",X"02",X"46",X"53",
		X"65",X"00",X"05",X"02",X"43",X"53",X"65",X"48",X"01",X"02",X"43",X"44",X"40",X"80",X"B0",X"01",
		X"60",X"44",X"43",X"40",X"86",X"01",X"07",X"10",X"03",X"12",X"97",X"65",X"52",X"08",X"54",X"66",
		X"54",X"2C",X"43",X"67",X"50",X"71",X"52",X"61",X"47",X"60",X"54",X"08",X"19",X"39",X"38",X"1B",
		X"54",X"45",X"64",X"63",X"67",X"08",X"61",X"66",X"43",X"3A",X"2D",X"66",X"63",X"1B",X"41",X"43",
		X"41",X"44",X"44",X"08",X"08",X"08",X"05",X"00",X"8D",X"39",X"B8",X"39",X"CC",X"1C",X"3A",X"2C",
		X"41",X"53",X"54",X"45",X"54",X"41",X"08",X"08",X"61",X"2B",X"77",X"3A",X"03",X"2A",X"66",X"67",
		X"66",X"41",X"65",X"45",X"2A",X"05",X"00",X"00",X"00",X"00",X"00",X"65",X"3A",X"86",X"20",X"9F",
		X"00",X"49",X"39",X"30",X"3A",X"15",X"39",X"54",X"41",X"42",X"64",X"45",X"53",X"08",X"08",X"57",
		X"2B",X"86",X"3A",X"03",X"2A",X"66",X"67",X"66",X"41",X"65",X"45",X"2A",X"06",X"00",X"00",X"00",
		X"00",X"00",X"5C",X"3A",X"86",X"20",X"27",X"00",X"04",X"1C",X"13",X"1C",X"9A",X"1A",X"61",X"66",
		X"61",X"54",X"53",X"08",X"08",X"08",X"4D",X"2B",X"BF",X"3A",X"03",X"2A",X"66",X"67",X"66",X"41",
		X"65",X"45",X"2A",X"07",X"00",X"00",X"00",X"00",X"00",X"CE",X"2E",X"05",X"00",X"D4",X"3A",X"CF",
		X"3A",X"F7",X"65",X"EE",X"2C",X"53",X"42",X"55",X"46",X"46",X"45",X"52",X"08",X"05",X"00",X"D4",
		X"3A",X"CF",X"3A",X"DD",X"65",X"80",X"19",X"64",X"43",X"66",X"54",X"08",X"08",X"08",X"08",X"5B",
		X"2B",X"D4",X"3A",X"03",X"2A",X"66",X"67",X"66",X"41",X"65",X"45",X"2A",X"20",X"00",X"00",X"00",
		X"00",X"00",X"9C",X"2D",X"81",X"2B",X"00",X"00",X"03",X"2A",X"66",X"67",X"66",X"41",X"65",X"45",
		X"2A",X"21",X"00",X"00",X"00",X"00",X"00",X"E9",X"3A",X"86",X"00",X"C2",X"66",X"F5",X"65",X"C2",
		X"66",X"67",X"38",X"50",X"52",X"67",X"52",X"41",X"65",X"08",X"08",X"F5",X"65",X"C2",X"66",X"E9",
		X"3A",X"00",X"00",X"00",X"1E",X"00",X"1F",X"00",X"22",X"3B",X"31",X"3A",X"FF",X"63",X"A7",X"2B",
		X"BC",X"33",X"2A",X"28",X"F8",X"2E",X"31",X"3B",X"00",X"2B",X"28",X"D0",X"19",X"CE",X"2E",X"0A",
		X"3B",X"00",X"D1",X"19",X"03",X"1C",X"9C",X"2D",X"2B",X"3B",X"00",X"04",X"1C",X"13",X"1C",X"5C",
		X"3A",X"1C",X"3B",X"00",X"14",X"1C",X"5B",X"1D",X"BA",X"39",X"3D",X"3B",X"00",X"5C",X"1D",X"48",
		X"39",X"DE",X"1E",X"46",X"3B",X"00",X"49",X"39",X"30",X"3A",X"65",X"3A",X"F0",X"1E",X"00",X"FE",
		X"A5",X"20",X"22",X"07",X"07",X"22",X"29",X"6F",X"21",X"FD",X"04",X"01",X"18",X"23",X"FB",X"85",
		X"20",X"23",X"01",X"58",X"23",X"FA",X"85",X"20",X"24",X"01",X"69",X"02",X"99",X"A0",X"02",X"BA",
		X"6A",X"20",X"25",X"01",X"77",X"02",X"8D",X"4B",X"23",X"29",X"76",X"05",X"2C",X"85",X"01",X"86",
		X"01",X"03",X"05",X"25",X"86",X"20",X"26",X"07",X"07",X"03",X"07",X"06",X"07",X"07",X"02",X"A4",
		X"62",X"20",X"27",X"03",X"22",X"DE",X"84",X"23",X"DD",X"41",X"03",X"25",X"20",X"23",X"FD",X"84",
		X"07",X"01",X"03",X"23",X"FC",X"1D",X"07",X"02",X"03",X"23",X"2B",X"87",X"02",X"DC",X"92",X"3D",
		X"01",X"A2",X"23",X"2D",X"A4",X"02",X"EB",X"A1",X"3D",X"13",X"00",X"07",X"04",X"07",X"20",X"03",
		X"21",X"FC",X"04",X"23",X"F6",X"92",X"09",X"23",X"08",X"81",X"23",X"F9",X"86",X"20",X"07",X"06",
		X"22",X"03",X"02",X"20",X"2C",X"01",X"79",X"23",X"F7",X"A1",X"02",X"C6",X"0C",X"06",X"23",X"03",
		X"01",X"1B",X"23",X"C8",X"C5",X"09",X"23",X"08",X"81",X"23",X"DF",X"88",X"23",X"2C",X"12",X"23",
		X"28",X"27",X"23",X"DE",X"87",X"37",X"07",X"01",X"89",X"01",X"06",X"37",X"F3",X"02",X"8B",X"7A",
		X"23",X"29",X"5F",X"3D",X"07",X"04",X"06",X"01",X"03",X"01",X"13",X"23",X"F9",X"96",X"37",X"06",
		X"23",X"2C",X"4F",X"23",X"28",X"4C",X"23",X"DE",X"49",X"23",X"29",X"76",X"07",X"03",X"06",X"24",
		X"03",X"25",X"20",X"02",X"3C",X"54",X"09",X"01",X"68",X"23",X"C9",X"A9",X"09",X"23",X"28",X"62",
		X"22",X"DE",X"91",X"37",X"D3",X"02",X"6B",X"42",X"23",X"29",X"3F",X"23",X"2C",X"3C",X"23",X"DF",
		X"39",X"01",X"41",X"23",X"29",X"1C",X"23",X"2C",X"19",X"22",X"DF",X"84",X"02",X"13",X"2B",X"09",
		X"01",X"63",X"01",X"0E",X"23",X"CA",X"9A",X"23",X"08",X"81",X"23",X"FA",X"A4",X"23",X"2C",X"5B",
		X"37",X"EB",X"23",X"FE",X"6E",X"06",X"01",X"03",X"23",X"F9",X"A3",X"23",X"2C",X"4D",X"23",X"F9",
		X"4A",X"37",X"20",X"01",X"59",X"23",X"28",X"73",X"23",X"F8",X"70",X"23",X"29",X"55",X"23",X"2C",
		X"52",X"37",X"CB",X"02",X"05",X"75",X"01",X"76",X"23",X"CB",X"A2",X"02",X"15",X"45",X"3D",X"07",
		X"03",X"06",X"25",X"03",X"04",X"00",X"00",X"00",X"00",X"69",X"48",X"66",X"0B",X"46",X"32",X"81",
		X"6F",X"13",X"32",X"A0",X"4F",X"E1",X"EB",X"77",X"16",X"00",X"EB",X"32",X"85",X"6F",X"13",X"32",
		X"A4",X"4F",X"E1",X"EB",X"77",X"16",X"00",X"EB",X"32",X"8D",X"6F",X"13",X"32",X"8C",X"4F",X"E1",
		X"44",X"65",X"09",X"00",X"00",X"3E",X"10",X"DD",X"29",X"EB",X"97",X"29",X"EB",X"A5",X"91",X"6F",
		X"7C",X"B0",X"4F",X"13",X"D2",X"F1",X"3C",X"21",X"33",X"D9",X"3D",X"C2",X"C7",X"3C",X"E1",X"76",
		X"0B",X"56",X"EB",X"29",X"CD",X"29",X"29",X"C1",X"21",X"E1",X"44",X"65",X"09",X"00",X"00",X"3E",
		X"10",X"29",X"EB",X"29",X"EB",X"D2",X"F9",X"3C",X"21",X"3D",X"C2",X"D9",X"3C",X"E1",X"71",X"50",
		X"EB",X"97",X"95",X"6F",X"3E",X"00",X"B4",X"4F",X"E1",X"EB",X"77",X"16",X"00",X"EB",X"32",X"9D",
		X"6F",X"13",X"32",X"9C",X"4F",X"E1",X"77",X"16",X"00",X"7B",X"95",X"6F",X"7A",X"B4",X"4F",X"E1",
		X"67",X"06",X"00",X"7B",X"91",X"6F",X"7A",X"B0",X"4F",X"E1",X"69",X"48",X"66",X"0B",X"46",X"32",
		X"91",X"6F",X"13",X"32",X"B0",X"4F",X"E1",X"6F",X"0E",X"00",X"32",X"95",X"6F",X"13",X"32",X"B4",
		X"4F",X"E1",X"77",X"16",X"00",X"7B",X"96",X"77",X"7A",X"0B",X"B6",X"57",X"EB",X"E1",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"93",X"1B",X"93",X"1B",X"58",X"0E",X"24",X"2A",X"B4",X"03",X"F8",X"29",X"EC",X"2E",X"48",X"2F",
		X"00",X"00",X"F1",X"13",X"9D",X"0C",X"65",X"0E",X"FF",X"7F",X"2F",X"03",X"BA",X"06",X"00",X"04",
		X"FC",X"03",X"F7",X"12",X"8F",X"03",X"D5",X"03",X"F3",X"03",X"A5",X"27",X"EA",X"03",X"DF",X"03",
		X"A2",X"03",X"00",X"12",X"25",X"12",X"32",X"12",X"E7",X"16",X"CA",X"03",X"21",X"13",X"1B",X"13",
		X"F2",X"E7",X"16",X"DA",X"20",X"D2",X"67",X"70",X"A2",X"03",X"F2",X"A8",X"C4",X"52",X"67",X"57",
		X"A5",X"27",X"85",X"C7",X"66",X"61",X"66",X"52",X"41",X"57",X"00",X"12",X"97",X"E5",X"52",X"54",
		X"8D",X"31",X"96",X"10",X"C5",X"64",X"54",X"61",X"54",X"56",X"32",X"A3",X"E5",X"71",X"53",X"AD",
		X"13",X"96",X"40",X"C2",X"55",X"53",X"98",X"14",X"F2",X"90",X"C7",X"66",X"61",X"52",X"54",X"53",
		X"D3",X"31",X"95",X"C5",X"64",X"54",X"61",X"54",X"53",X"06",X"34",X"A4",X"E4",X"52",X"53",X"1C",
		X"12",X"F1",X"38",X"C1",X"52",X"53",X"89",X"14",X"F1",X"28",X"C5",X"43",X"41",X"50",X"53",X"2E",
		X"16",X"A1",X"D0",X"53",X"78",X"00",X"F8",X"18",X"C1",X"64",X"53",X"9A",X"34",X"F1",X"08",X"D2",
		X"60",X"53",X"89",X"12",X"B7",X"E4",X"60",X"53",X"C1",X"12",X"B6",X"D4",X"45",X"53",X"DF",X"34",
		X"F0",X"C0",X"C7",X"45",X"53",X"94",X"00",X"B2",X"E6",X"67",X"61",X"54",X"43",X"45",X"53",X"0F",
		X"12",X"8A",X"00",X"C6",X"43",X"53",X"26",X"35",X"D1",X"1F",X"D2",X"41",X"64",X"41",X"43",X"53",
		X"6B",X"35",X"8F",X"C3",X"42",X"53",X"78",X"30",X"F4",X"B0",X"42",X"D4",X"53",X"52",X"5F",X"15",
		X"F7",X"C4",X"52",X"52",X"D1",X"12",X"D2",X"4F",X"C1",X"43",X"52",X"52",X"B8",X"00",X"D1",X"27",
		X"C3",X"52",X"52",X"59",X"16",X"F1",X"20",X"C1",X"52",X"52",X"C2",X"00",X"D1",X"37",X"D2",X"52",
		X"CD",X"00",X"F1",X"30",X"C4",X"64",X"52",X"F6",X"00",X"D2",X"6F",X"C1",X"43",X"64",X"52",X"4D",
		X"16",X"D1",X"07",X"C3",X"64",X"52",X"49",X"12",X"F1",X"00",X"C1",X"64",X"52",X"DA",X"00",X"D1",
		X"17",X"E4",X"52",X"20",X"01",X"F1",X"10",X"E6",X"54",X"45",X"52",X"D0",X"00",X"D2",X"45",X"E1",
		X"54",X"45",X"52",X"91",X"12",X"D2",X"65",X"D4",X"45",X"52",X"15",X"01",X"D7",X"E1",X"C5",X"65",
		X"55",X"53",X"45",X"52",X"01",X"01",X"8D",X"C5",X"56",X"52",X"45",X"53",X"45",X"52",X"7D",X"16",
		X"8C",X"01",X"D3",X"45",X"52",X"D6",X"00",X"F0",X"80",X"D4",X"41",X"45",X"50",X"45",X"52",X"40",
		X"01",X"A7",X"D2",X"27",X"01",X"DB",X"E0",X"53",X"55",X"50",X"51",X"01",X"F6",X"C5",X"D0",X"67",
		X"50",X"2C",X"01",X"F6",X"C1",X"E7",X"50",X"0D",X"01",X"DA",X"08",X"C5",X"50",X"F9",X"00",X"DA",
		X"28",X"C5",X"47",X"41",X"50",X"26",X"17",X"A0",X"30",X"D0",X"63",X"16",X"DA",X"18",X"E1",X"54",
		X"55",X"67",X"5F",X"01",X"D2",X"8B",X"C4",X"54",X"55",X"67",X"66",X"15",X"D2",X"AB",X"D4",X"55",
		X"67",X"A4",X"01",X"C9",X"41",X"D2",X"61",X"54",X"67",X"71",X"16",X"D2",X"9B",X"D2",X"44",X"54",
		X"67",X"7C",X"01",X"D2",X"BB",X"C7",X"52",X"67",X"E7",X"14",X"81",X"D2",X"67",X"85",X"15",X"F2",
		X"98",X"F2",X"66",X"43",X"12",X"DA",X"00",X"D0",X"67",X"66",X"7F",X"31",X"D1",X"00",X"D4",X"53",
		X"61",X"64",X"67",X"66",X"88",X"00",X"87",X"C7",X"45",X"66",X"45",X"35",X"D2",X"44",X"D2",X"60",
		X"43",X"66",X"8B",X"01",X"B4",X"C3",X"66",X"03",X"33",X"DA",X"10",X"C5",X"65",X"41",X"66",X"D4",
		X"01",X"AB",X"C4",X"67",X"65",X"78",X"34",X"B5",X"C7",X"45",X"65",X"8E",X"17",X"96",X"D8",X"C5",
		X"65",X"38",X"35",X"96",X"FF",X"E7",X"52",X"43",X"41",X"65",X"F5",X"32",X"91",X"E5",X"6F",X"17",
		X"DA",X"38",X"E7",X"64",X"EA",X"32",X"B1",X"D4",X"53",X"61",X"64",X"19",X"15",X"86",X"D2",X"61",
		X"44",X"64",X"A2",X"17",X"D2",X"98",X"E1",X"44",X"64",X"F7",X"14",X"D2",X"88",X"D2",X"44",X"44",
		X"64",X"93",X"17",X"D2",X"B8",X"C4",X"44",X"64",X"06",X"02",X"D2",X"A8",X"C4",X"64",X"14",X"02",
		X"D0",X"E4",X"33",X"02",X"DD",X"05",X"D2",X"62",X"CA",X"15",X"D3",X"30",X"D0",X"62",X"1C",X"02",
		X"D5",X"C3",X"F1",X"61",X"18",X"02",X"FC",X"08",X"F0",X"61",X"81",X"17",X"FD",X"08",X"C5",X"47");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
