`define BUILD_DATE "190908"
`define BUILD_TIME "210120"
