library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity rom_cpu2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of rom_cpu2 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"74",X"06",X"DD",X"75",X"07",X"DD",X"77",X"08",X"08",X"FD",X"72",X"00",X"FD",X"73",X"01",X"FD",
		X"77",X"02",X"C5",X"79",X"87",X"4F",X"87",X"87",X"81",X"5F",X"16",X"00",X"21",X"A3",X"6A",X"19",
		X"11",X"89",X"6A",X"06",X"0A",X"1A",X"4E",X"EB",X"12",X"71",X"EB",X"13",X"23",X"10",X"F6",X"C1",
		X"FD",X"23",X"FD",X"23",X"FD",X"23",X"0C",X"10",X"B3",X"3E",X"04",X"CD",X"A0",X"1B",X"3E",X"24",
		X"21",X"00",X"D3",X"01",X"01",X"60",X"D7",X"DD",X"36",X"01",X"B4",X"DD",X"36",X"03",X"00",X"DD",
		X"36",X"04",X"00",X"DD",X"36",X"05",X"00",X"DD",X"36",X"13",X"FF",X"CD",X"62",X"22",X"CD",X"C0",
		X"21",X"CD",X"E2",X"21",X"CD",X"08",X"22",X"CD",X"27",X"22",X"1E",X"14",X"CD",X"91",X"0F",X"3A",
		X"0B",X"60",X"A7",X"C2",X"8E",X"21",X"CD",X"08",X"22",X"CD",X"53",X"1B",X"06",X"05",X"CD",X"76",
		X"0F",X"CD",X"0C",X"22",X"CD",X"53",X"1B",X"06",X"05",X"CD",X"76",X"0F",X"DD",X"35",X"01",X"CA",
		X"75",X"21",X"3A",X"00",X"60",X"21",X"00",X"90",X"CB",X"6F",X"28",X"03",X"21",X"01",X"90",X"CB",
		X"56",X"28",X"06",X"CB",X"46",X"28",X"1D",X"18",X"47",X"CD",X"E6",X"21",X"DD",X"7E",X"03",X"3C",
		X"FE",X"0E",X"38",X"0B",X"DD",X"7E",X"04",X"FE",X"03",X"30",X"23",X"DD",X"34",X"04",X"AF",X"DD",
		X"77",X"03",X"18",X"1A",X"CD",X"E6",X"21",X"DD",X"7E",X"03",X"A7",X"28",X"03",X"3D",X"18",X"0B",
		X"DD",X"7E",X"04",X"A7",X"28",X"08",X"DD",X"35",X"04",X"3E",X"0D",X"DD",X"77",X"03",X"CD",X"E2",
		X"21",X"1E",X"07",X"21",X"32",X"60",X"34",X"CB",X"46",X"20",X"02",X"1E",X"08",X"CD",X"91",X"0F",
		X"3A",X"00",X"60",X"CB",X"6F",X"20",X"0E",X"3A",X"00",X"90",X"CB",X"5F",X"28",X"19",X"CB",X"4F",
		X"28",X"15",X"C3",X"10",X"21",X"3A",X"01",X"90",X"CB",X"5F",X"28",X"0B",X"CB",X"4F",X"28",X"07",
		X"DD",X"36",X"13",X"FF",X"C3",X"6F",X"20",X"DD",X"7E",X"03",X"DD",X"BE",X"13",X"CA",X"6F",X"20",
		X"DD",X"77",X"13",X"FE",X"0D",X"20",X"25",X"DD",X"7E",X"04",X"FE",X"03",X"CA",X"75",X"21",X"DD",
		X"7E",X"05",X"A7",X"CA",X"6F",X"20",X"CD",X"0C",X"22",X"DD",X"35",X"05",X"CD",X"08",X"22",X"3E",
		X"24",X"CD",X"99",X"21",X"1E",X"03",X"CD",X"91",X"0F",X"C3",X"6F",X"20",X"CD",X"44",X"22",X"B8",
		X"D2",X"6F",X"20",X"DD",X"7E",X"04",X"07",X"07",X"47",X"07",X"80",X"DD",X"86",X"04",X"DD",X"86",
		X"03",X"CD",X"99",X"21",X"CD",X"0C",X"22",X"DD",X"34",X"05",X"CD",X"08",X"22",X"1E",X"09",X"CD",
		X"91",X"0F",X"C3",X"6F",X"20",X"1E",X"0F",X"CD",X"91",X"0F",X"CD",X"5D",X"22",X"0E",X"12",X"3A",
		X"0B",X"60",X"A7",X"C2",X"8E",X"21",X"06",X"0A",X"CD",X"76",X"0F",X"0D",X"20",X"F1",X"CD",X"8C",
		X"3B",X"CD",X"7C",X"1B",X"FD",X"E1",X"DD",X"E1",X"C9",X"DD",X"5E",X"00",X"CB",X"23",X"CB",X"23",
		X"16",X"00",X"21",X"D1",X"22",X"19",X"CF",X"E5",X"F5",X"CD",X"55",X"22",X"4F",X"F1",X"06",X"00",
		X"09",X"77",X"EB",X"CF",X"EB",X"E1",X"CD",X"47",X"22",X"7E",X"12",X"23",X"13",X"10",X"FA",X"C9",
		X"AF",X"21",X"62",X"D2",X"0E",X"04",X"06",X"0D",X"77",X"3C",X"23",X"23",X"10",X"FA",X"11",X"26",
		X"00",X"19",X"0D",X"20",X"F1",X"21",X"E5",X"22",X"06",X"04",X"C5",X"CD",X"39",X"1D",X"C1",X"10",
		X"F9",X"C9",X"0E",X"38",X"18",X"02",X"0E",X"24",X"DD",X"7E",X"04",X"21",X"82",X"D2",X"A7",X"28",
		X"07",X"11",X"40",X"00",X"47",X"19",X"10",X"FD",X"DD",X"7E",X"03",X"87",X"5F",X"16",X"00",X"19",
		X"71",X"CB",X"D4",X"36",X"06",X"CB",X"94",X"C9",X"0E",X"39",X"18",X"02",X"0E",X"24",X"DD",X"7E",
		X"00",X"21",X"31",X"D1",X"A7",X"28",X"07",X"11",X"40",X"00",X"47",X"19",X"10",X"FD",X"CD",X"55",
		X"22",X"5F",X"16",X"00",X"19",X"71",X"C9",X"21",X"1B",X"D1",X"3A",X"02",X"90",X"CB",X"57",X"20",
		X"03",X"21",X"14",X"D1",X"DD",X"7E",X"00",X"A7",X"28",X"07",X"11",X"40",X"00",X"47",X"19",X"10",
		X"FD",X"36",X"28",X"C9",X"DD",X"7E",X"05",X"E5",X"21",X"02",X"90",X"06",X"0A",X"CB",X"56",X"20",
		X"02",X"06",X"03",X"E1",X"C9",X"CD",X"44",X"22",X"B8",X"D8",X"78",X"3D",X"C9",X"3E",X"01",X"CD",
		X"A0",X"1B",X"21",X"B3",X"22",X"06",X"05",X"C5",X"CD",X"39",X"1D",X"C1",X"10",X"F9",X"DD",X"E5",
		X"21",X"0A",X"D1",X"DD",X"21",X"94",X"6A",X"06",X"05",X"11",X"3A",X"00",X"C5",X"06",X"06",X"CD",
		X"95",X"1E",X"19",X"C1",X"10",X"F6",X"DD",X"E1",X"21",X"A3",X"6A",X"11",X"11",X"D1",X"CD",X"AA",
		X"22",X"11",X"51",X"D1",X"CD",X"AA",X"22",X"11",X"91",X"D1",X"CD",X"AA",X"22",X"11",X"D1",X"D1",
		X"CD",X"AA",X"22",X"11",X"11",X"D2",X"CD",X"AA",X"22",X"C9",X"06",X"0A",X"7E",X"12",X"23",X"13",
		X"10",X"FA",X"C9",X"05",X"D1",X"03",X"17",X"18",X"01",X"45",X"D1",X"03",X"17",X"18",X"02",X"85",
		X"D1",X"03",X"17",X"18",X"03",X"C5",X"D1",X"03",X"17",X"18",X"04",X"05",X"D2",X"03",X"17",X"18",
		X"05",X"A3",X"6A",X"11",X"D1",X"AD",X"6A",X"51",X"D1",X"B7",X"6A",X"91",X"D1",X"C1",X"6A",X"D1",
		X"D1",X"CB",X"6A",X"11",X"D2",X"7C",X"D2",X"02",X"34",X"35",X"BC",X"D2",X"02",X"34",X"35",X"FC",
		X"D2",X"02",X"34",X"35",X"3C",X"D3",X"02",X"36",X"37",X"E5",X"2A",X"D8",X"0B",X"ED",X"5B",X"52",
		X"60",X"AF",X"ED",X"52",X"D1",X"19",X"C9",X"21",X"59",X"60",X"34",X"7E",X"FE",X"07",X"38",X"02",
		X"36",X"06",X"CD",X"15",X"0E",X"CD",X"3C",X"0E",X"CD",X"E8",X"0E",X"3A",X"60",X"60",X"CB",X"7F",
		X"28",X"03",X"CD",X"F0",X"0E",X"C9",X"E5",X"21",X"2C",X"60",X"3A",X"00",X"60",X"CB",X"6F",X"28",
		X"03",X"21",X"2E",X"60",X"34",X"7E",X"FE",X"20",X"30",X"07",X"E1",X"1E",X"54",X"16",X"00",X"F7",
		X"C9",X"36",X"00",X"23",X"7E",X"3C",X"27",X"77",X"E1",X"16",X"01",X"5F",X"CB",X"3B",X"CB",X"3B",
		X"CB",X"3B",X"CB",X"3B",X"28",X"0B",X"E5",X"F5",X"7D",X"C6",X"1F",X"E6",X"1F",X"6F",X"F7",X"F1",
		X"E1",X"E6",X"0F",X"5F",X"F7",X"C9",X"21",X"30",X"60",X"3A",X"00",X"60",X"CB",X"6F",X"28",X"03",
		X"21",X"31",X"60",X"3A",X"15",X"60",X"47",X"E6",X"0F",X"CB",X"78",X"20",X"03",X"86",X"18",X"03",
		X"96",X"ED",X"44",X"4F",X"E5",X"3E",X"FC",X"CD",X"31",X"0F",X"C6",X"1C",X"B9",X"30",X"0B",X"3E",
		X"FC",X"CD",X"3C",X"0F",X"D6",X"20",X"B9",X"38",X"01",X"79",X"E1",X"77",X"C9",X"DD",X"E5",X"DD",
		X"21",X"E8",X"61",X"DD",X"36",X"00",X"80",X"DD",X"36",X"02",X"00",X"DD",X"36",X"0E",X"00",X"DD",
		X"E1",X"C9",X"3A",X"60",X"60",X"E6",X"0F",X"FE",X"0F",X"20",X"27",X"21",X"51",X"60",X"7E",X"FE",
		X"04",X"D0",X"34",X"5F",X"16",X"00",X"21",X"43",X"24",X"19",X"5E",X"16",X"05",X"D5",X"21",X"30",
		X"60",X"3A",X"00",X"60",X"CB",X"6F",X"28",X"03",X"21",X"31",X"60",X"7E",X"CD",X"01",X"24",X"D1",
		X"F7",X"C9",X"AF",X"32",X"51",X"60",X"DD",X"34",X"03",X"DD",X"7E",X"03",X"FE",X"03",X"D8",X"DD",
		X"36",X"03",X"00",X"C0",X"3A",X"E8",X"61",X"A7",X"C8",X"CD",X"66",X"23",X"CD",X"01",X"24",X"18",
		X"1A",X"2F",X"E6",X"F8",X"6F",X"26",X"00",X"29",X"29",X"11",X"00",X"D0",X"19",X"3A",X"55",X"60",
		X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"5F",X"16",X"00",X"19",X"C9",X"7E",X"FE",X"24",X"C0",X"3A",
		X"F6",X"61",X"0E",X"00",X"D6",X"05",X"38",X"03",X"0C",X"18",X"F9",X"79",X"FE",X"04",X"38",X"02",
		X"0E",X"03",X"06",X"00",X"E5",X"21",X"3F",X"24",X"09",X"56",X"E1",X"1E",X"53",X"F7",X"C9",X"02",
		X"01",X"06",X"00",X"13",X"1E",X"16",X"19",X"DD",X"7E",X"02",X"21",X"4E",X"24",X"DF",X"56",X"24",
		X"A0",X"24",X"D2",X"25",X"E4",X"25",X"DD",X"7E",X"0E",X"FE",X"14",X"D8",X"3A",X"59",X"60",X"3D",
		X"5F",X"16",X"00",X"21",X"95",X"26",X"19",X"7E",X"DD",X"77",X"0B",X"DD",X"36",X"02",X"01",X"3E",
		X"F8",X"CD",X"31",X"0F",X"47",X"3E",X"F8",X"CD",X"3C",X"0F",X"90",X"CB",X"3F",X"80",X"DD",X"77",
		X"07",X"DD",X"36",X"06",X"00",X"DD",X"36",X"04",X"00",X"DD",X"36",X"05",X"00",X"DD",X"36",X"08",
		X"00",X"DD",X"36",X"09",X"08",X"DD",X"36",X"0A",X"0A",X"DD",X"CB",X"00",X"E6",X"C3",X"CB",X"25",
		X"CD",X"6A",X"0F",X"C3",X"CB",X"25",X"ED",X"5B",X"52",X"60",X"DD",X"6E",X"04",X"DD",X"66",X"05",
		X"AF",X"ED",X"52",X"DD",X"75",X"04",X"DD",X"74",X"05",X"7C",X"FE",X"08",X"30",X"0F",X"DD",X"35",
		X"0B",X"C2",X"6F",X"24",X"DD",X"36",X"0E",X"00",X"DD",X"36",X"02",X"00",X"C9",X"CD",X"46",X"33",
		X"FE",X"08",X"D2",X"AA",X"25",X"CD",X"53",X"33",X"FE",X"08",X"D2",X"AA",X"25",X"DD",X"CB",X"00",
		X"EE",X"21",X"C5",X"69",X"36",X"80",X"3E",X"02",X"32",X"2B",X"62",X"32",X"48",X"62",X"32",X"65",
		X"62",X"32",X"82",X"62",X"32",X"9F",X"62",X"32",X"BC",X"62",X"3A",X"59",X"60",X"3D",X"87",X"47",
		X"87",X"80",X"5F",X"16",X"00",X"21",X"9B",X"26",X"19",X"01",X"06",X"00",X"11",X"F8",X"61",X"ED",
		X"B0",X"DD",X"7E",X"14",X"CB",X"3F",X"DD",X"77",X"14",X"DD",X"77",X"15",X"DD",X"36",X"16",X"00",
		X"CD",X"45",X"3E",X"06",X"02",X"FE",X"02",X"38",X"02",X"06",X"03",X"DD",X"7E",X"17",X"80",X"DD",
		X"77",X"17",X"DD",X"36",X"03",X"02",X"DD",X"36",X"02",X"02",X"21",X"01",X"00",X"22",X"13",X"60",
		X"AF",X"32",X"12",X"60",X"CD",X"C4",X"1E",X"3E",X"0C",X"CD",X"BE",X"0F",X"3E",X"02",X"CD",X"BE",
		X"0F",X"3E",X"02",X"CD",X"BE",X"0F",X"3E",X"11",X"CD",X"BE",X"0F",X"3E",X"10",X"CD",X"86",X"0F",
		X"3E",X"05",X"CD",X"86",X"0F",X"CD",X"50",X"26",X"21",X"E2",X"61",X"CB",X"E6",X"21",X"02",X"62",
		X"36",X"03",X"21",X"D6",X"62",X"11",X"A9",X"63",X"CD",X"95",X"1B",X"DD",X"E5",X"DD",X"21",X"A9",
		X"63",X"DD",X"CB",X"00",X"7E",X"28",X"04",X"DD",X"36",X"02",X"05",X"DD",X"21",X"BE",X"63",X"DD",
		X"CB",X"00",X"7E",X"28",X"04",X"DD",X"36",X"02",X"05",X"DD",X"21",X"D3",X"63",X"DD",X"CB",X"00",
		X"7E",X"28",X"04",X"DD",X"36",X"02",X"05",X"DD",X"E1",X"C9",X"DD",X"35",X"0A",X"20",X"1C",X"DD",
		X"36",X"0A",X"0A",X"DD",X"CB",X"00",X"66",X"28",X"0A",X"DD",X"CB",X"00",X"A6",X"DD",X"36",X"08",
		X"00",X"18",X"08",X"DD",X"CB",X"00",X"E6",X"DD",X"36",X"08",X"01",X"21",X"BF",X"26",X"CD",X"D1",
		X"07",X"C9",X"DD",X"35",X"10",X"C0",X"DD",X"7E",X"11",X"A7",X"28",X"04",X"DD",X"35",X"11",X"C9",
		X"DD",X"36",X"02",X"03",X"DD",X"35",X"15",X"20",X"20",X"DD",X"7E",X"14",X"DD",X"77",X"15",X"DD",
		X"7E",X"03",X"2F",X"E6",X"03",X"DD",X"77",X"03",X"CB",X"47",X"28",X"0A",X"CD",X"7B",X"26",X"3E",
		X"03",X"CD",X"86",X"0F",X"18",X"03",X"CD",X"67",X"26",X"DD",X"35",X"12",X"C0",X"DD",X"7E",X"13",
		X"A7",X"28",X"04",X"DD",X"35",X"13",X"C9",X"21",X"00",X"62",X"CB",X"7E",X"20",X"05",X"DD",X"36",
		X"12",X"01",X"C9",X"CB",X"66",X"20",X"08",X"CD",X"7B",X"26",X"21",X"02",X"62",X"36",X"10",X"CD",
		X"5E",X"29",X"DD",X"CB",X"00",X"AE",X"DD",X"36",X"02",X"00",X"DD",X"36",X"0E",X"00",X"DD",X"36",
		X"17",X"00",X"DD",X"E5",X"DD",X"21",X"C5",X"69",X"06",X"26",X"CD",X"8D",X"1B",X"DD",X"E1",X"C9",
		X"11",X"E0",X"D4",X"21",X"F5",X"67",X"01",X"10",X"01",X"1A",X"ED",X"6F",X"13",X"1A",X"ED",X"6F",
		X"13",X"23",X"0B",X"79",X"B0",X"20",X"F2",X"16",X"07",X"21",X"E0",X"D4",X"01",X"20",X"02",X"7E",
		X"E6",X"F8",X"82",X"77",X"23",X"0B",X"79",X"B0",X"20",X"F5",X"C9",X"11",X"E0",X"D4",X"21",X"F5",
		X"67",X"01",X"10",X"01",X"ED",X"6F",X"12",X"13",X"ED",X"6F",X"12",X"ED",X"6F",X"13",X"23",X"0B",
		X"79",X"B0",X"20",X"F0",X"C9",X"03",X"03",X"02",X"02",X"01",X"01",X"D2",X"00",X"96",X"00",X"1E",
		X"05",X"B4",X"00",X"78",X"00",X"18",X"05",X"A5",X"00",X"69",X"00",X"15",X"05",X"96",X"00",X"5A",
		X"00",X"12",X"05",X"87",X"00",X"4B",X"00",X"0F",X"05",X"78",X"00",X"3C",X"00",X"0C",X"05",X"78",
		X"00",X"7C",X"00",X"DD",X"36",X"09",X"03",X"DD",X"CB",X"00",X"C6",X"DD",X"7E",X"05",X"CD",X"31",
		X"0F",X"C6",X"08",X"DD",X"BE",X"07",X"38",X"0A",X"DD",X"36",X"02",X"02",X"DD",X"36",X"08",X"07",
		X"18",X"22",X"DD",X"36",X"08",X"06",X"DD",X"6E",X"06",X"DD",X"66",X"07",X"11",X"00",X"FC",X"19",
		X"DD",X"75",X"06",X"DD",X"74",X"07",X"CD",X"47",X"27",X"DD",X"7E",X"05",X"FE",X"08",X"38",X"D8",
		X"FE",X"F8",X"30",X"D4",X"C9",X"DD",X"7E",X"05",X"FE",X"08",X"38",X"04",X"FE",X"F8",X"38",X"37",
		X"DD",X"36",X"02",X"00",X"DD",X"CB",X"00",X"86",X"DD",X"CB",X"00",X"9E",X"CD",X"13",X"1F",X"3A",
		X"15",X"60",X"E6",X"3F",X"DD",X"77",X"01",X"DD",X"CB",X"00",X"F6",X"DD",X"36",X"05",X"02",X"3A",
		X"16",X"60",X"E6",X"3F",X"C6",X"B8",X"DD",X"77",X"19",X"E6",X"07",X"5F",X"16",X"00",X"21",X"5C",
		X"27",X"19",X"7E",X"DD",X"77",X"07",X"C9",X"2A",X"52",X"60",X"CD",X"43",X"1F",X"EB",X"DD",X"6E",
		X"04",X"DD",X"66",X"05",X"19",X"DD",X"75",X"04",X"DD",X"74",X"05",X"C9",X"80",X"98",X"7C",X"8C",
		X"78",X"90",X"84",X"88",X"DD",X"7E",X"05",X"FE",X"08",X"D8",X"FE",X"F8",X"D0",X"DD",X"7E",X"03",
		X"FE",X"02",X"C2",X"A2",X"27",X"DD",X"7E",X"05",X"DD",X"CB",X"00",X"5E",X"20",X"04",X"C6",X"08",
		X"18",X"02",X"D6",X"08",X"CD",X"31",X"0F",X"C6",X"10",X"DD",X"BE",X"07",X"DA",X"0E",X"28",X"DD",
		X"34",X"07",X"DD",X"CB",X"00",X"5E",X"C2",X"D1",X"27",X"DD",X"5E",X"11",X"DD",X"56",X"12",X"C3",
		X"C6",X"27",X"DD",X"7E",X"05",X"DD",X"CB",X"00",X"5E",X"20",X"04",X"C6",X"1C",X"18",X"02",X"D6",
		X"04",X"CD",X"31",X"0F",X"C6",X"10",X"DD",X"BE",X"07",X"DA",X"0E",X"28",X"DD",X"CB",X"00",X"5E",
		X"20",X"0F",X"ED",X"5B",X"52",X"60",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"AF",X"ED",X"52",X"18",
		X"0D",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"DD",X"5E",X"11",X"DD",X"56",X"12",X"19",X"DD",X"75",
		X"04",X"DD",X"74",X"05",X"DD",X"34",X"07",X"DD",X"34",X"07",X"DD",X"CB",X"15",X"C6",X"DD",X"CB",
		X"14",X"7E",X"28",X"0F",X"DD",X"6E",X"13",X"DD",X"66",X"14",X"CD",X"43",X"1F",X"DD",X"75",X"13",
		X"DD",X"74",X"14",X"DD",X"36",X"16",X"00",X"DD",X"36",X"17",X"00",X"C3",X"AC",X"28",X"DD",X"7E",
		X"03",X"FE",X"02",X"C2",X"43",X"28",X"DD",X"7E",X"05",X"DD",X"CB",X"00",X"5E",X"20",X"04",X"C6",
		X"08",X"18",X"02",X"D6",X"08",X"CD",X"3C",X"0F",X"D6",X"08",X"DD",X"BE",X"07",X"D2",X"AC",X"28",
		X"DD",X"35",X"07",X"DD",X"CB",X"00",X"5E",X"C2",X"72",X"28",X"DD",X"5E",X"11",X"DD",X"56",X"12",
		X"C3",X"67",X"28",X"DD",X"7E",X"05",X"DD",X"CB",X"00",X"5E",X"20",X"04",X"C6",X"1C",X"18",X"02",
		X"00",X"00",X"CD",X"3C",X"0F",X"D6",X"08",X"DD",X"BE",X"07",X"D2",X"AC",X"28",X"DD",X"CB",X"00",
		X"5E",X"20",X"0F",X"ED",X"5B",X"52",X"60",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"AF",X"ED",X"52",
		X"18",X"0D",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"DD",X"5E",X"11",X"DD",X"56",X"12",X"19",X"DD",
		X"75",X"04",X"DD",X"74",X"05",X"DD",X"35",X"07",X"DD",X"35",X"07",X"DD",X"CB",X"15",X"86",X"DD",
		X"CB",X"14",X"7E",X"20",X"0F",X"DD",X"6E",X"13",X"DD",X"66",X"14",X"CD",X"43",X"1F",X"DD",X"75",
		X"13",X"DD",X"74",X"14",X"DD",X"36",X"16",X"00",X"DD",X"36",X"17",X"00",X"3A",X"00",X"62",X"E6",
		X"30",X"C2",X"09",X"29",X"CD",X"46",X"33",X"FE",X"0A",X"30",X"4E",X"57",X"CD",X"53",X"33",X"FE",
		X"0A",X"30",X"46",X"5F",X"3A",X"E8",X"61",X"CB",X"6F",X"28",X"11",X"21",X"00",X"62",X"CB",X"4E",
		X"C2",X"35",X"29",X"CB",X"CE",X"DD",X"36",X"02",X"04",X"C3",X"35",X"29",X"3A",X"05",X"62",X"DD",
		X"CB",X"00",X"5E",X"20",X"0D",X"DD",X"BE",X"05",X"30",X"15",X"7A",X"FE",X"07",X"38",X"10",X"C3",
		X"09",X"29",X"DD",X"BE",X"05",X"38",X"08",X"7A",X"FE",X"07",X"38",X"03",X"C3",X"09",X"29",X"DD",
		X"36",X"08",X"01",X"CD",X"60",X"33",X"C3",X"35",X"29",X"FD",X"21",X"69",X"63",X"FD",X"CB",X"00",
		X"7E",X"28",X"09",X"CD",X"36",X"29",X"C3",X"1C",X"29",X"C3",X"2C",X"29",X"FD",X"21",X"7B",X"63",
		X"FD",X"CB",X"00",X"7E",X"28",X"0F",X"CD",X"36",X"29",X"C3",X"35",X"29",X"DD",X"36",X"02",X"01",
		X"3E",X"09",X"CD",X"86",X"0F",X"C9",X"FD",X"56",X"05",X"FD",X"5E",X"07",X"CD",X"4E",X"29",X"FE",
		X"14",X"D0",X"CD",X"56",X"29",X"FE",X"14",X"D0",X"E1",X"23",X"23",X"23",X"E5",X"C9",X"DD",X"7E",
		X"05",X"92",X"D0",X"ED",X"44",X"C9",X"DD",X"7E",X"07",X"93",X"D0",X"ED",X"44",X"C9",X"21",X"28",
		X"62",X"11",X"D6",X"62",X"CD",X"95",X"1B",X"DD",X"E5",X"DD",X"21",X"28",X"62",X"DD",X"36",X"00",
		X"C0",X"CD",X"45",X"3E",X"87",X"5F",X"16",X"00",X"21",X"D5",X"29",X"19",X"46",X"23",X"4E",X"DD",
		X"70",X"01",X"DD",X"36",X"03",X"01",X"DD",X"36",X"05",X"02",X"DD",X"36",X"07",X"90",X"DD",X"36",
		X"19",X"D0",X"DD",X"21",X"45",X"62",X"DD",X"36",X"00",X"C0",X"DD",X"71",X"01",X"DD",X"36",X"03",
		X"01",X"DD",X"36",X"05",X"02",X"DD",X"36",X"07",X"80",X"DD",X"36",X"19",X"E0",X"CD",X"45",X"3E",
		X"FE",X"02",X"38",X"1E",X"DD",X"21",X"62",X"62",X"DD",X"36",X"00",X"C0",X"79",X"C6",X"1E",X"DD",
		X"77",X"01",X"DD",X"36",X"03",X"01",X"DD",X"36",X"05",X"02",X"DD",X"36",X"07",X"70",X"DD",X"36",
		X"19",X"D8",X"DD",X"E1",X"C9",X"3C",X"B4",X"28",X"78",X"19",X"50",X"0A",X"28",X"21",X"E8",X"61",
		X"CB",X"7E",X"C8",X"11",X"60",X"28",X"CD",X"0B",X"39",X"01",X"60",X"0A",X"11",X"20",X"00",X"FE",
		X"53",X"28",X"0F",X"79",X"C6",X"08",X"4F",X"AF",X"ED",X"52",X"7E",X"FE",X"53",X"28",X"03",X"10",
		X"F2",X"C9",X"CB",X"D4",X"CB",X"5E",X"CB",X"94",X"20",X"F5",X"CD",X"45",X"3E",X"06",X"04",X"FE",
		X"02",X"38",X"02",X"06",X"03",X"3A",X"FF",X"61",X"B8",X"D0",X"36",X"24",X"5F",X"3C",X"32",X"FF",
		X"61",X"CB",X"23",X"16",X"00",X"21",X"6B",X"2E",X"19",X"CD",X"45",X"3E",X"1E",X"04",X"FE",X"02",
		X"38",X"02",X"1E",X"06",X"16",X"00",X"19",X"CF",X"DD",X"E5",X"E5",X"DD",X"E1",X"DD",X"36",X"00",
		X"80",X"DD",X"36",X"02",X"07",X"DD",X"36",X"03",X"00",X"DD",X"36",X"05",X"28",X"DD",X"71",X"07",
		X"DD",X"36",X"08",X"00",X"DD",X"36",X"09",X"01",X"DD",X"36",X"0C",X"0A",X"3A",X"15",X"60",X"E6",
		X"3F",X"C6",X"B8",X"DD",X"77",X"19",X"DD",X"E1",X"3E",X"06",X"CD",X"86",X"0F",X"C9",X"DD",X"7E",
		X"02",X"21",X"75",X"2A",X"DF",X"EE",X"2A",X"87",X"2C",X"8E",X"2C",X"9B",X"2C",X"A0",X"2C",X"FE",
		X"2C",X"24",X"2D",X"5B",X"2D",X"84",X"2D",X"DD",X"7E",X"00",X"E6",X"03",X"20",X"43",X"CD",X"93",
		X"2A",X"18",X"26",X"DD",X"7E",X"0A",X"A7",X"28",X"05",X"DD",X"35",X"0A",X"18",X"17",X"DD",X"7E",
		X"0B",X"3C",X"FE",X"03",X"38",X"01",X"AF",X"DD",X"77",X"0B",X"5F",X"16",X"00",X"21",X"EB",X"2A",
		X"19",X"7E",X"DD",X"77",X"0A",X"DD",X"7E",X"0B",X"C9",X"DD",X"CB",X"00",X"5E",X"28",X"02",X"C6",
		X"03",X"DD",X"77",X"08",X"21",X"E8",X"2A",X"DD",X"5E",X"03",X"16",X"00",X"19",X"7E",X"DD",X"77",
		X"09",X"21",X"D8",X"2A",X"CD",X"D1",X"07",X"C9",X"90",X"20",X"94",X"20",X"98",X"20",X"90",X"00",
		X"94",X"00",X"98",X"00",X"A8",X"00",X"AC",X"00",X"01",X"0F",X"02",X"05",X"02",X"0A",X"CD",X"6A",
		X"0F",X"C3",X"0B",X"2B",X"3A",X"60",X"60",X"E6",X"0F",X"FE",X"0F",X"20",X"07",X"DD",X"36",X"02",
		X"06",X"C3",X"6E",X"2A",X"DD",X"7E",X"03",X"21",X"16",X"2B",X"DF",X"21",X"E8",X"61",X"CB",X"6E",
		X"CA",X"D1",X"2A",X"C3",X"52",X"2C",X"1C",X"2B",X"65",X"2B",X"C5",X"2B",X"DD",X"CB",X"00",X"6E",
		X"20",X"36",X"DD",X"CB",X"00",X"EE",X"DD",X"CB",X"00",X"9E",X"3A",X"15",X"60",X"CB",X"7F",X"28",
		X"0E",X"DD",X"CB",X"15",X"86",X"DD",X"36",X"13",X"20",X"DD",X"36",X"14",X"FF",X"18",X"0C",X"DD",
		X"CB",X"15",X"C6",X"DD",X"36",X"13",X"E0",X"DD",X"36",X"14",X"00",X"DD",X"36",X"16",X"00",X"DD",
		X"36",X"17",X"00",X"DD",X"36",X"1C",X"20",X"C9",X"CD",X"91",X"2D",X"CD",X"25",X"2E",X"CD",X"64",
		X"27",X"CD",X"87",X"2A",X"C9",X"DD",X"CB",X"00",X"56",X"20",X"2C",X"DD",X"CB",X"00",X"D6",X"DD",
		X"CB",X"00",X"9E",X"DD",X"CB",X"15",X"C6",X"21",X"C0",X"00",X"CD",X"18",X"2E",X"DD",X"75",X"13",
		X"DD",X"74",X"14",X"DD",X"36",X"16",X"00",X"DD",X"36",X"17",X"00",X"CD",X"45",X"3E",X"07",X"07",
		X"07",X"C6",X"28",X"DD",X"77",X"1C",X"C9",X"CD",X"91",X"2D",X"DD",X"CB",X"00",X"5E",X"20",X"1B",
		X"11",X"40",X"00",X"3A",X"07",X"62",X"DD",X"BE",X"07",X"30",X"03",X"11",X"C0",X"FF",X"DD",X"6E",
		X"06",X"DD",X"66",X"07",X"19",X"DD",X"75",X"06",X"DD",X"74",X"07",X"CD",X"25",X"2E",X"CD",X"64",
		X"27",X"CD",X"87",X"2A",X"C9",X"DD",X"CB",X"00",X"66",X"C2",X"EE",X"2B",X"DD",X"CB",X"00",X"E6",
		X"21",X"00",X"02",X"DD",X"CB",X"15",X"46",X"20",X"03",X"21",X"00",X"FE",X"DD",X"75",X"13",X"DD",
		X"74",X"14",X"DD",X"36",X"16",X"00",X"DD",X"36",X"17",X"00",X"DD",X"36",X"1C",X"70",X"11",X"80",
		X"FF",X"DD",X"7E",X"0B",X"FE",X"02",X"20",X"03",X"11",X"80",X"02",X"DD",X"73",X"11",X"DD",X"72",
		X"12",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"DD",X"CB",X"00",X"5E",X"20",X"0C",X"19",X"7C",X"FE",
		X"B8",X"38",X"12",X"DD",X"CB",X"00",X"DE",X"18",X"0C",X"AF",X"ED",X"52",X"7C",X"FE",X"38",X"30",
		X"04",X"DD",X"CB",X"00",X"9E",X"DD",X"75",X"04",X"DD",X"74",X"05",X"11",X"80",X"00",X"3A",X"07",
		X"62",X"DD",X"BE",X"07",X"38",X"03",X"11",X"80",X"FF",X"DD",X"6E",X"06",X"DD",X"66",X"07",X"19",
		X"DD",X"75",X"06",X"DD",X"74",X"07",X"CD",X"25",X"2E",X"CD",X"64",X"27",X"CD",X"93",X"2A",X"DD",
		X"77",X"08",X"3E",X"02",X"21",X"EB",X"61",X"CB",X"46",X"28",X"02",X"3E",X"0F",X"DD",X"77",X"09",
		X"21",X"67",X"2C",X"CD",X"D1",X"07",X"C9",X"A0",X"00",X"A4",X"00",X"9C",X"00",X"A0",X"00",X"A4",
		X"00",X"9C",X"00",X"B0",X"00",X"B4",X"00",X"B8",X"00",X"BC",X"00",X"C0",X"00",X"C4",X"00",X"C8",
		X"00",X"CC",X"00",X"F4",X"00",X"F8",X"00",X"CD",X"C3",X"26",X"CD",X"87",X"2A",X"C9",X"CD",X"6A",
		X"0F",X"C3",X"97",X"2C",X"CD",X"05",X"27",X"CD",X"87",X"2A",X"C9",X"DD",X"36",X"02",X"00",X"C9",
		X"3E",X"04",X"CD",X"86",X"0F",X"21",X"00",X"62",X"CB",X"BE",X"3A",X"05",X"62",X"DD",X"77",X"05",
		X"3A",X"07",X"62",X"DD",X"77",X"07",X"21",X"FE",X"61",X"7E",X"E5",X"87",X"5F",X"16",X"00",X"21",
		X"77",X"2E",X"19",X"56",X"23",X"5E",X"EB",X"22",X"13",X"60",X"AF",X"32",X"12",X"60",X"CD",X"C4",
		X"1E",X"E1",X"7E",X"34",X"DD",X"77",X"08",X"21",X"2A",X"60",X"3A",X"00",X"60",X"CB",X"6F",X"28",
		X"03",X"21",X"2B",X"60",X"7E",X"C6",X"01",X"27",X"77",X"CD",X"EF",X"3A",X"DD",X"36",X"09",X"02",
		X"DD",X"36",X"01",X"0A",X"DD",X"34",X"02",X"21",X"73",X"2C",X"CD",X"D1",X"07",X"C9",X"DD",X"35",
		X"01",X"20",X"F4",X"21",X"00",X"62",X"CB",X"FE",X"06",X"1D",X"CD",X"8D",X"1B",X"21",X"FF",X"61",
		X"35",X"C0",X"DD",X"E5",X"DD",X"21",X"E8",X"61",X"CD",X"17",X"26",X"DD",X"E1",X"C9",X"06",X"1D",
		X"CD",X"8D",X"1B",X"C9",X"3A",X"05",X"62",X"DD",X"BE",X"05",X"30",X"08",X"21",X"80",X"00",X"CD",
		X"F9",X"22",X"18",X"06",X"2A",X"52",X"60",X"CD",X"43",X"1F",X"EB",X"DD",X"6E",X"04",X"DD",X"66",
		X"05",X"19",X"DD",X"75",X"04",X"DD",X"74",X"05",X"7C",X"FE",X"08",X"38",X"04",X"FE",X"F8",X"38",
		X"03",X"C3",X"1E",X"2D",X"CD",X"64",X"27",X"CD",X"87",X"2A",X"C9",X"DD",X"35",X"0C",X"20",X"0B",
		X"DD",X"34",X"02",X"DD",X"36",X"0C",X"0A",X"DD",X"36",X"08",X"01",X"11",X"00",X"01",X"DD",X"6E",
		X"04",X"DD",X"66",X"05",X"AF",X"ED",X"52",X"DD",X"75",X"04",X"DD",X"74",X"05",X"21",X"83",X"2C",
		X"CD",X"D1",X"07",X"C9",X"DD",X"35",X"0C",X"C2",X"6B",X"2D",X"DD",X"36",X"02",X"00",X"C3",X"EE",
		X"2A",X"DD",X"CB",X"00",X"5E",X"20",X"3E",X"21",X"E0",X"FF",X"DD",X"7E",X"0B",X"FE",X"02",X"20",
		X"06",X"21",X"20",X"01",X"CD",X"18",X"2E",X"CD",X"F9",X"22",X"DD",X"75",X"11",X"DD",X"74",X"12",
		X"DD",X"5E",X"04",X"DD",X"56",X"05",X"19",X"DD",X"75",X"04",X"DD",X"74",X"05",X"7C",X"DD",X"BE",
		X"19",X"DA",X"17",X"2E",X"DD",X"CB",X"00",X"DE",X"3A",X"15",X"60",X"E6",X"1F",X"C6",X"0C",X"DD",
		X"77",X"19",X"C3",X"17",X"2E",X"DD",X"7E",X"0B",X"FE",X"02",X"20",X"0E",X"21",X"C0",X"01",X"CD",
		X"18",X"2E",X"E5",X"C1",X"CD",X"60",X"0F",X"EB",X"18",X"03",X"11",X"00",X"00",X"DD",X"73",X"11",
		X"DD",X"72",X"12",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"AF",X"ED",X"52",X"DD",X"75",X"04",X"DD",
		X"74",X"05",X"7C",X"DD",X"BE",X"19",X"D2",X"17",X"2E",X"DD",X"CB",X"00",X"9E",X"3A",X"15",X"60",
		X"E6",X"3F",X"C6",X"B8",X"DD",X"77",X"19",X"C9",X"CD",X"45",X"3E",X"07",X"07",X"07",X"07",X"07",
		X"5F",X"16",X"00",X"19",X"C9",X"DD",X"6E",X"06",X"DD",X"66",X"07",X"DD",X"5E",X"13",X"DD",X"56",
		X"14",X"19",X"DD",X"75",X"06",X"DD",X"74",X"07",X"DD",X"6E",X"16",X"DD",X"66",X"17",X"19",X"DD",
		X"75",X"16",X"DD",X"74",X"17",X"7C",X"CB",X"7F",X"20",X"0B",X"DD",X"BE",X"1C",X"38",X"1B",X"DD",
		X"CB",X"15",X"86",X"18",X"0B",X"ED",X"44",X"DD",X"BE",X"1C",X"38",X"0E",X"DD",X"CB",X"15",X"C6",
		X"EB",X"CD",X"43",X"1F",X"DD",X"75",X"13",X"DD",X"74",X"14",X"C9",X"28",X"62",X"45",X"62",X"62",
		X"62",X"7F",X"62",X"9C",X"62",X"B9",X"62",X"00",X"01",X"50",X"01",X"00",X"02",X"50",X"02",X"00",
		X"03",X"50",X"03",X"B8",X"78",X"E6",X"0A",X"28",X"20",X"21",X"0D",X"32",X"FE",X"02",X"20",X"02",
		X"23",X"23",X"5E",X"23",X"56",X"DD",X"6E",X"0D",X"DD",X"66",X"0E",X"19",X"7C",X"FE",X"08",X"30",
		X"02",X"26",X"08",X"DD",X"75",X"0D",X"DD",X"74",X"0E",X"DD",X"7E",X"05",X"D6",X"04",X"CD",X"31",
		X"0F",X"DD",X"86",X"0E",X"C6",X"08",X"DD",X"77",X"07",X"DD",X"46",X"0D",X"DD",X"70",X"06",X"DD",
		X"7E",X"05",X"C6",X"04",X"CD",X"31",X"0F",X"FE",X"44",X"20",X"10",X"3A",X"60",X"60",X"FE",X"0F",
		X"3E",X"48",X"20",X"07",X"DD",X"36",X"02",X"0A",X"C3",X"D4",X"35",X"57",X"1E",X"00",X"DD",X"6E",
		X"06",X"DD",X"66",X"07",X"AF",X"ED",X"52",X"7C",X"D6",X"08",X"30",X"02",X"3E",X"04",X"DD",X"75",
		X"0B",X"DD",X"77",X"0C",X"C9",X"DD",X"7E",X"05",X"CD",X"31",X"0F",X"C6",X"06",X"DD",X"BE",X"07",
		X"DA",X"0E",X"2F",X"DD",X"36",X"0C",X"08",X"DD",X"36",X"0E",X"08",X"C3",X"4C",X"2F",X"DD",X"7E",
		X"07",X"C6",X"08",X"4F",X"DD",X"7E",X"05",X"CD",X"3C",X"0F",X"B9",X"28",X"01",X"D0",X"FE",X"C8",
		X"38",X"2A",X"DD",X"7E",X"07",X"D6",X"C0",X"4F",X"DD",X"7E",X"07",X"91",X"DD",X"77",X"07",X"DD",
		X"7E",X"0C",X"91",X"DD",X"77",X"0C",X"DD",X"7E",X"0E",X"91",X"DD",X"77",X"0E",X"C9",X"DD",X"36",
		X"02",X"08",X"DD",X"CB",X"00",X"96",X"DD",X"36",X"1D",X"F8",X"18",X"09",X"DD",X"36",X"03",X"04",
		X"E1",X"23",X"23",X"23",X"E5",X"E1",X"23",X"23",X"23",X"E5",X"C9",X"DD",X"5E",X"08",X"16",X"00",
		X"21",X"3B",X"32",X"19",X"7E",X"DD",X"77",X"09",X"21",X"11",X"32",X"CD",X"D1",X"07",X"DD",X"7E",
		X"0E",X"DD",X"CB",X"00",X"DE",X"DD",X"BE",X"0C",X"38",X"07",X"DD",X"CB",X"00",X"9E",X"DD",X"7E",
		X"0C",X"DD",X"36",X"10",X"00",X"47",X"DD",X"56",X"05",X"DD",X"7E",X"07",X"D6",X"10",X"5F",X"78",
		X"D6",X"08",X"30",X"07",X"ED",X"44",X"83",X"5F",X"C3",X"E2",X"2F",X"CD",X"C8",X"32",X"78",X"A7",
		X"28",X"19",X"C5",X"CD",X"40",X"08",X"21",X"95",X"32",X"CD",X"AE",X"08",X"7B",X"D6",X"10",X"5F",
		X"DD",X"7E",X"10",X"C6",X"10",X"DD",X"77",X"10",X"C1",X"10",X"E7",X"79",X"A7",X"28",X"23",X"C5",
		X"DD",X"7E",X"05",X"C6",X"03",X"DD",X"CB",X"00",X"5E",X"28",X"02",X"D6",X"08",X"57",X"CD",X"40",
		X"08",X"C1",X"7B",X"91",X"5F",X"79",X"87",X"81",X"4F",X"06",X"00",X"21",X"98",X"32",X"09",X"CD",
		X"AE",X"08",X"DD",X"7E",X"05",X"C6",X"04",X"DD",X"CB",X"00",X"5E",X"28",X"02",X"D6",X"08",X"57",
		X"7B",X"C6",X"04",X"5F",X"CD",X"76",X"08",X"DD",X"CB",X"00",X"66",X"20",X"1B",X"DD",X"5E",X"1A",
		X"DD",X"56",X"1B",X"2A",X"52",X"60",X"19",X"7C",X"FE",X"06",X"38",X"06",X"21",X"00",X"00",X"DD",
		X"34",X"1C",X"DD",X"75",X"1A",X"DD",X"74",X"1B",X"21",X"50",X"32",X"DD",X"CB",X"1C",X"46",X"28",
		X"03",X"21",X"53",X"32",X"CD",X"AE",X"08",X"DD",X"7E",X"0C",X"DD",X"CB",X"00",X"5E",X"20",X"03",
		X"DD",X"7E",X"0E",X"47",X"D6",X"08",X"30",X"0D",X"ED",X"44",X"DD",X"86",X"07",X"D6",X"10",X"5F",
		X"01",X"00",X"00",X"18",X"12",X"78",X"DD",X"96",X"10",X"D6",X"08",X"CD",X"C8",X"32",X"DD",X"7E",
		X"07",X"DD",X"96",X"10",X"D6",X"10",X"5F",X"DD",X"7E",X"05",X"D6",X"05",X"DD",X"CB",X"00",X"5E",
		X"28",X"02",X"C6",X"08",X"57",X"78",X"A7",X"28",X"11",X"C5",X"CD",X"40",X"08",X"21",X"C5",X"32",
		X"CD",X"AE",X"08",X"7B",X"D6",X"10",X"5F",X"C1",X"10",X"EF",X"79",X"A7",X"28",X"15",X"C5",X"CD",
		X"40",X"08",X"C1",X"7B",X"91",X"5F",X"79",X"87",X"81",X"4F",X"06",X"00",X"21",X"98",X"32",X"09",
		X"CD",X"AE",X"08",X"7B",X"C6",X"04",X"5F",X"14",X"CD",X"76",X"08",X"21",X"50",X"32",X"DD",X"CB",
		X"1C",X"46",X"28",X"03",X"21",X"53",X"32",X"CD",X"AE",X"08",X"C9",X"DD",X"CB",X"00",X"E6",X"DD",
		X"36",X"08",X"13",X"DD",X"E5",X"06",X"04",X"DD",X"7E",X"04",X"DD",X"77",X"13",X"DD",X"23",X"10",
		X"F6",X"DD",X"E1",X"DD",X"36",X"17",X"05",X"DD",X"34",X"02",X"CD",X"8C",X"3B",X"3E",X"0D",X"CD",
		X"86",X"0F",X"DD",X"56",X"14",X"DD",X"5E",X"16",X"21",X"89",X"32",X"CD",X"0C",X"09",X"C3",X"5B",
		X"2F",X"DD",X"35",X"17",X"20",X"EC",X"DD",X"34",X"02",X"DD",X"7E",X"0C",X"DD",X"BE",X"0E",X"38",
		X"03",X"DD",X"7E",X"0E",X"FE",X"09",X"30",X"19",X"DD",X"34",X"02",X"DD",X"36",X"08",X"14",X"DD",
		X"36",X"09",X"03",X"DD",X"36",X"01",X"0F",X"DD",X"7E",X"07",X"D6",X"08",X"DD",X"77",X"07",X"18",
		X"1A",X"DD",X"35",X"0C",X"DD",X"35",X"0C",X"DD",X"35",X"0E",X"DD",X"35",X"0E",X"DD",X"35",X"07",
		X"DD",X"35",X"07",X"C3",X"5B",X"2F",X"DD",X"35",X"01",X"28",X"07",X"21",X"11",X"32",X"CD",X"D1",
		X"07",X"C9",X"3A",X"60",X"60",X"E6",X"0F",X"FE",X"0F",X"20",X"15",X"CD",X"3C",X"39",X"21",X"2A",
		X"60",X"3A",X"00",X"60",X"CB",X"6F",X"28",X"03",X"21",X"2B",X"60",X"36",X"00",X"CD",X"07",X"23",
		X"21",X"28",X"60",X"3A",X"00",X"60",X"CB",X"6F",X"28",X"03",X"21",X"29",X"60",X"36",X"01",X"3A",
		X"D5",X"61",X"CB",X"7F",X"28",X"07",X"3E",X"02",X"32",X"D7",X"61",X"18",X"0A",X"21",X"DD",X"61",
		X"36",X"80",X"21",X"E2",X"61",X"CB",X"A6",X"06",X"78",X"CD",X"76",X"0F",X"C9",X"DD",X"CB",X"00",
		X"56",X"20",X"31",X"DD",X"CB",X"00",X"D6",X"DD",X"7E",X"07",X"DD",X"86",X"1D",X"DD",X"77",X"07",
		X"DD",X"7E",X"0C",X"DD",X"86",X"1D",X"FE",X"F0",X"38",X"02",X"3E",X"08",X"DD",X"77",X"0C",X"DD",
		X"7E",X"0E",X"DD",X"86",X"1D",X"FE",X"F0",X"38",X"02",X"3E",X"08",X"DD",X"77",X"0E",X"DD",X"36",
		X"11",X"0C",X"18",X"2E",X"DD",X"35",X"11",X"20",X"0A",X"DD",X"36",X"02",X"00",X"DD",X"CB",X"00",
		X"96",X"18",X"1F",X"3E",X"04",X"DD",X"CB",X"11",X"46",X"20",X"02",X"ED",X"44",X"47",X"DD",X"86",
		X"07",X"DD",X"77",X"07",X"DD",X"7E",X"0C",X"80",X"DD",X"77",X"0C",X"DD",X"7E",X"0E",X"80",X"DD",
		X"77",X"0E",X"C9",X"06",X"48",X"DD",X"7E",X"07",X"D6",X"08",X"DD",X"96",X"0C",X"B8",X"30",X"06",
		X"DD",X"36",X"02",X"04",X"18",X"10",X"DD",X"6E",X"06",X"DD",X"66",X"07",X"11",X"00",X"FD",X"19",
		X"DD",X"75",X"06",X"DD",X"74",X"07",X"C3",X"5B",X"2F",X"00",X"FD",X"00",X"02",X"00",X"02",X"00",
		X"FE",X"20",X"00",X"24",X"00",X"28",X"00",X"08",X"00",X"0C",X"00",X"00",X"00",X"04",X"00",X"10",
		X"00",X"14",X"00",X"00",X"20",X"04",X"20",X"08",X"20",X"0C",X"20",X"2C",X"20",X"FC",X"20",X"10",
		X"10",X"14",X"10",X"2C",X"00",X"FC",X"00",X"18",X"00",X"1C",X"00",X"00",X"00",X"00",X"0A",X"0A",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"00",X"03",
		X"74",X"00",X"0D",X"75",X"00",X"0D",X"70",X"00",X"00",X"30",X"00",X"00",X"34",X"00",X"00",X"38",
		X"00",X"00",X"3C",X"00",X"00",X"40",X"00",X"00",X"44",X"00",X"00",X"48",X"00",X"00",X"4C",X"00",
		X"00",X"50",X"00",X"00",X"54",X"00",X"00",X"58",X"00",X"00",X"5C",X"00",X"00",X"60",X"00",X"00",
		X"64",X"00",X"00",X"68",X"00",X"00",X"6C",X"00",X"00",X"80",X"00",X"02",X"84",X"00",X"02",X"88",
		X"00",X"02",X"8C",X"00",X"02",X"A0",X"01",X"0C",X"60",X"01",X"0C",X"64",X"01",X"0C",X"68",X"01",
		X"0C",X"6C",X"01",X"0C",X"70",X"01",X"0C",X"74",X"01",X"0C",X"78",X"01",X"0C",X"7C",X"01",X"0C",
		X"80",X"01",X"0C",X"84",X"01",X"0C",X"88",X"01",X"0C",X"8C",X"01",X"0C",X"90",X"01",X"0C",X"94",
		X"01",X"0C",X"98",X"01",X"0C",X"9C",X"01",X"0C",X"01",X"00",X"00",X"D6",X"10",X"38",X"03",X"04",
		X"18",X"F9",X"C6",X"10",X"4F",X"C9",X"DD",X"E5",X"DD",X"21",X"00",X"62",X"06",X"28",X"CD",X"8D",
		X"1B",X"DD",X"36",X"00",X"80",X"DD",X"36",X"05",X"40",X"DD",X"36",X"0E",X"10",X"DD",X"7E",X"05",
		X"D6",X"04",X"CD",X"31",X"0F",X"C6",X"18",X"DD",X"77",X"07",X"DD",X"7E",X"05",X"C6",X"04",X"CD",
		X"31",X"0F",X"47",X"DD",X"7E",X"07",X"D6",X"08",X"90",X"30",X"02",X"3E",X"08",X"DD",X"77",X"0C",
		X"DD",X"7E",X"05",X"C6",X"04",X"CD",X"3C",X"0F",X"D6",X"08",X"DD",X"BE",X"07",X"30",X"18",X"DD",
		X"36",X"0E",X"08",X"DD",X"7E",X"07",X"D6",X"08",X"DD",X"77",X"07",X"DD",X"7E",X"0C",X"D6",X"08",
		X"30",X"02",X"3E",X"08",X"DD",X"77",X"0C",X"DD",X"E1",X"C9",X"DD",X"E5",X"DD",X"21",X"00",X"62",
		X"CD",X"5B",X"2F",X"DD",X"E1",X"C9",X"06",X"00",X"3A",X"05",X"62",X"DD",X"96",X"05",X"D0",X"ED",
		X"44",X"05",X"C9",X"0E",X"00",X"3A",X"07",X"62",X"DD",X"96",X"07",X"D0",X"ED",X"44",X"0D",X"C9",
		X"21",X"00",X"62",X"CB",X"EE",X"21",X"03",X"62",X"36",X"04",X"C9",X"DD",X"7E",X"02",X"21",X"72",
		X"33",X"DF",X"96",X"33",X"17",X"34",X"AB",X"34",X"C1",X"34",X"AC",X"35",X"AF",X"35",X"B2",X"35",
		X"B5",X"35",X"B8",X"35",X"D1",X"35",X"D4",X"35",X"3F",X"36",X"72",X"37",X"3F",X"36",X"77",X"37",
		X"3F",X"36",X"0E",X"35",X"62",X"35",X"DD",X"CB",X"00",X"6E",X"28",X"0E",X"DD",X"7E",X"03",X"DD",
		X"77",X"02",X"21",X"E2",X"61",X"CB",X"E6",X"C3",X"6B",X"33",X"CD",X"B2",X"37",X"CD",X"0E",X"2F",
		X"C3",X"B9",X"33",X"C3",X"F4",X"33",X"C3",X"9C",X"33",X"DD",X"7E",X"0A",X"A7",X"20",X"15",X"CD",
		X"A0",X"38",X"C3",X"F4",X"33",X"DD",X"36",X"0A",X"01",X"DD",X"36",X"08",X"01",X"DD",X"36",X"1E",
		X"03",X"C3",X"13",X"34",X"DD",X"35",X"1E",X"C2",X"13",X"34",X"DD",X"36",X"08",X"02",X"CD",X"E9",
		X"38",X"21",X"F6",X"61",X"34",X"DD",X"36",X"0A",X"00",X"DD",X"36",X"1F",X"00",X"DD",X"36",X"20",
		X"01",X"C3",X"13",X"34",X"DD",X"34",X"1F",X"DD",X"7E",X"1F",X"FE",X"08",X"38",X"07",X"DD",X"36",
		X"1F",X"00",X"DD",X"34",X"20",X"DD",X"36",X"08",X"00",X"DD",X"CB",X"20",X"46",X"28",X"04",X"DD",
		X"36",X"08",X"02",X"CD",X"5B",X"2F",X"C9",X"DD",X"CB",X"00",X"AE",X"DD",X"CB",X"00",X"4E",X"28",
		X"10",X"21",X"E2",X"61",X"CB",X"E6",X"DD",X"36",X"01",X"04",X"DD",X"36",X"02",X"02",X"C3",X"85",
		X"34",X"CD",X"B2",X"37",X"CD",X"82",X"38",X"CD",X"F5",X"2E",X"C3",X"43",X"34",X"C3",X"4C",X"34",
		X"C3",X"9C",X"33",X"CD",X"A0",X"38",X"C3",X"4C",X"34",X"CD",X"E9",X"38",X"DD",X"7E",X"26",X"A7",
		X"28",X"15",X"DD",X"BE",X"27",X"28",X"10",X"DD",X"77",X"27",X"5F",X"16",X"00",X"21",X"9B",X"34",
		X"19",X"7E",X"DD",X"77",X"08",X"18",X"1A",X"DD",X"7E",X"18",X"A7",X"28",X"06",X"DD",X"35",X"18",
		X"C3",X"85",X"34",X"DD",X"CB",X"08",X"46",X"20",X"05",X"DD",X"35",X"08",X"18",X"03",X"DD",X"34",
		X"08",X"DD",X"36",X"18",X"02",X"DD",X"36",X"09",X"0A",X"3A",X"EB",X"61",X"CB",X"47",X"28",X"04",
		X"DD",X"36",X"09",X"00",X"21",X"11",X"32",X"CD",X"D1",X"07",X"C9",X"03",X"0B",X"0F",X"0D",X"03",
		X"03",X"11",X"03",X"07",X"09",X"03",X"03",X"05",X"03",X"03",X"03",X"DD",X"35",X"01",X"C2",X"85",
		X"34",X"21",X"E2",X"61",X"CB",X"A6",X"DD",X"36",X"02",X"01",X"DD",X"CB",X"00",X"8E",X"C3",X"85",
		X"34",X"DD",X"CB",X"00",X"AE",X"11",X"00",X"02",X"DD",X"6E",X"0B",X"DD",X"66",X"0C",X"AF",X"ED",
		X"52",X"7C",X"FE",X"08",X"38",X"1C",X"DD",X"75",X"0B",X"DD",X"74",X"0C",X"DD",X"6E",X"0D",X"DD",
		X"66",X"0E",X"AF",X"ED",X"52",X"7C",X"FE",X"08",X"38",X"08",X"DD",X"75",X"0D",X"DD",X"74",X"0E",
		X"18",X"14",X"21",X"E2",X"61",X"CB",X"A6",X"DD",X"36",X"02",X"01",X"DD",X"36",X"08",X"03",X"DD",
		X"36",X"18",X"02",X"C3",X"85",X"34",X"DD",X"36",X"08",X"02",X"CD",X"5B",X"2F",X"C9",X"3E",X"10",
		X"CD",X"BE",X"0F",X"21",X"E2",X"61",X"CB",X"E6",X"DD",X"34",X"02",X"DD",X"7E",X"05",X"C6",X"04",
		X"CD",X"31",X"0F",X"C6",X"08",X"47",X"DD",X"7E",X"07",X"90",X"38",X"04",X"FE",X"08",X"30",X"02",
		X"3E",X"08",X"DD",X"77",X"12",X"DD",X"7E",X"05",X"D6",X"04",X"CD",X"31",X"0F",X"C6",X"08",X"4F",
		X"DD",X"7E",X"07",X"91",X"38",X"04",X"FE",X"08",X"30",X"02",X"3E",X"08",X"DD",X"77",X"19",X"DD",
		X"36",X"0B",X"00",X"DD",X"36",X"0C",X"08",X"DD",X"36",X"0D",X"00",X"DD",X"36",X"0E",X"08",X"C3",
		X"A4",X"35",X"DD",X"6E",X"0D",X"DD",X"66",X"0E",X"11",X"A0",X"01",X"19",X"DD",X"75",X"0D",X"DD",
		X"74",X"0E",X"7C",X"DD",X"BE",X"19",X"30",X"13",X"DD",X"6E",X"0B",X"DD",X"66",X"0C",X"19",X"DD",
		X"75",X"0B",X"DD",X"74",X"0C",X"7C",X"DD",X"BE",X"12",X"38",X"19",X"DD",X"7E",X"12",X"DD",X"77",
		X"0C",X"DD",X"7E",X"19",X"DD",X"77",X"0E",X"21",X"E2",X"61",X"CB",X"A6",X"DD",X"36",X"02",X"00",
		X"DD",X"36",X"0A",X"00",X"DD",X"36",X"08",X"00",X"CD",X"5B",X"2F",X"C9",X"C3",X"AB",X"30",X"C3",
		X"E1",X"30",X"C3",X"E9",X"30",X"C3",X"26",X"31",X"DD",X"CB",X"00",X"6E",X"C2",X"9C",X"33",X"CD",
		X"7D",X"31",X"CD",X"A9",X"2E",X"CD",X"0E",X"2F",X"C3",X"B9",X"33",X"C3",X"F4",X"33",X"C3",X"9C",
		X"33",X"C3",X"E3",X"31",X"DD",X"CB",X"00",X"6E",X"C2",X"9C",X"33",X"DD",X"CB",X"00",X"46",X"20",
		X"3B",X"DD",X"CB",X"00",X"C6",X"3E",X"0E",X"CD",X"86",X"0F",X"3E",X"10",X"CD",X"BE",X"0F",X"3E",
		X"13",X"CD",X"86",X"0F",X"DD",X"36",X"01",X"0C",X"DD",X"36",X"21",X"00",X"DD",X"36",X"22",X"00",
		X"DD",X"36",X"23",X"05",X"DD",X"36",X"24",X"00",X"DD",X"36",X"07",X"B8",X"DD",X"36",X"0C",X"08",
		X"DD",X"36",X"0E",X"08",X"DD",X"36",X"08",X"02",X"CD",X"5B",X"2F",X"C9",X"DD",X"7E",X"0C",X"FE",
		X"10",X"30",X"06",X"DD",X"34",X"0C",X"DD",X"34",X"0E",X"DD",X"35",X"01",X"20",X"EA",X"DD",X"34",
		X"02",X"DD",X"36",X"08",X"01",X"DD",X"36",X"25",X"01",X"DD",X"CB",X"00",X"86",X"18",X"D9",X"DD",
		X"CB",X"00",X"6E",X"C2",X"9C",X"33",X"DD",X"6E",X"21",X"DD",X"66",X"22",X"DD",X"5E",X"23",X"DD",
		X"56",X"24",X"AF",X"ED",X"52",X"DD",X"75",X"21",X"DD",X"74",X"22",X"EB",X"DD",X"6E",X"06",X"DD",
		X"66",X"07",X"19",X"DD",X"75",X"06",X"DD",X"74",X"07",X"CD",X"43",X"38",X"DD",X"CB",X"25",X"46",
		X"C2",X"97",X"36",X"DD",X"CB",X"22",X"7E",X"20",X"13",X"06",X"00",X"DD",X"35",X"12",X"DD",X"CB",
		X"12",X"56",X"28",X"02",X"06",X"02",X"DD",X"70",X"08",X"C3",X"18",X"36",X"DD",X"CB",X"25",X"C6",
		X"DD",X"36",X"08",X"01",X"C3",X"18",X"36",X"DD",X"7E",X"02",X"FE",X"0B",X"20",X"14",X"DD",X"7E",
		X"05",X"D6",X"04",X"CD",X"31",X"0F",X"DD",X"BE",X"07",X"38",X"07",X"DD",X"36",X"03",X"04",X"C3",
		X"9C",X"33",X"DD",X"7E",X"07",X"FE",X"98",X"30",X"1B",X"06",X"0F",X"FE",X"68",X"30",X"04",X"06",
		X"08",X"18",X"0B",X"4F",X"3E",X"98",X"D6",X"06",X"B9",X"38",X"03",X"05",X"18",X"F8",X"DD",X"70",
		X"0C",X"DD",X"70",X"0E",X"DD",X"7E",X"02",X"FE",X"0F",X"CA",X"3B",X"37",X"DD",X"7E",X"07",X"FE",
		X"68",X"30",X"55",X"FE",X"60",X"38",X"45",X"21",X"8D",X"63",X"CB",X"7E",X"28",X"13",X"3A",X"99",
		X"63",X"D6",X"14",X"DD",X"BE",X"05",X"30",X"09",X"C6",X"28",X"DD",X"BE",X"05",X"38",X"02",X"18",
		X"18",X"21",X"9B",X"63",X"CB",X"7E",X"28",X"30",X"3A",X"A7",X"63",X"D6",X"10",X"DD",X"BE",X"05",
		X"30",X"26",X"C6",X"20",X"DD",X"BE",X"05",X"38",X"1F",X"3E",X"0B",X"CD",X"86",X"0F",X"3E",X"0E",
		X"CD",X"86",X"0F",X"DD",X"36",X"08",X"02",X"DD",X"34",X"02",X"18",X"0C",X"FE",X"58",X"30",X"08",
		X"DD",X"36",X"03",X"04",X"DD",X"CB",X"00",X"EE",X"C3",X"18",X"36",X"DD",X"7E",X"07",X"FE",X"58",
		X"30",X"F6",X"DD",X"56",X"05",X"1E",X"4C",X"CD",X"0B",X"39",X"FE",X"A4",X"FE",X"A4",X"DA",X"AB",
		X"36",X"FE",X"A8",X"D2",X"AB",X"36",X"CD",X"2B",X"39",X"CD",X"07",X"23",X"CD",X"9F",X"3A",X"CD",
		X"EF",X"3A",X"DD",X"36",X"02",X"00",X"CD",X"5E",X"29",X"CD",X"9D",X"23",X"3E",X"14",X"CD",X"86",
		X"0F",X"C9",X"21",X"06",X"00",X"18",X"03",X"21",X"08",X"00",X"DD",X"75",X"23",X"DD",X"74",X"24",
		X"DD",X"6E",X"21",X"DD",X"66",X"22",X"CD",X"43",X"1F",X"DD",X"75",X"21",X"DD",X"74",X"22",X"DD",
		X"CB",X"25",X"86",X"DD",X"7E",X"07",X"C6",X"08",X"DD",X"77",X"07",X"DD",X"36",X"0C",X"10",X"DD",
		X"36",X"0E",X"10",X"DD",X"36",X"08",X"02",X"DD",X"36",X"12",X"00",X"DD",X"34",X"02",X"CD",X"5B",
		X"2F",X"C9",X"3A",X"D5",X"61",X"CB",X"7F",X"28",X"05",X"3A",X"D8",X"61",X"18",X"0F",X"21",X"00",
		X"90",X"3A",X"00",X"60",X"CB",X"6F",X"28",X"03",X"21",X"01",X"90",X"7E",X"2F",X"E6",X"0F",X"DD",
		X"77",X"26",X"47",X"E6",X"05",X"CA",X"37",X"38",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"ED",X"5B",
		X"52",X"60",X"D5",X"FE",X"01",X"20",X"28",X"ED",X"5B",X"09",X"32",X"19",X"7C",X"FE",X"38",X"30",
		X"03",X"21",X"00",X"38",X"DD",X"75",X"04",X"DD",X"74",X"05",X"E1",X"ED",X"5B",X"DE",X"0B",X"19",
		X"ED",X"5B",X"DA",X"0B",X"E5",X"AF",X"ED",X"52",X"E1",X"30",X"01",X"EB",X"C3",X"34",X"38",X"ED",
		X"5B",X"0B",X"32",X"19",X"7C",X"FE",X"B8",X"38",X"03",X"21",X"00",X"B8",X"DD",X"75",X"04",X"DD",
		X"74",X"05",X"E1",X"ED",X"5B",X"DC",X"0B",X"19",X"ED",X"5B",X"D8",X"0B",X"E5",X"AF",X"ED",X"52",
		X"E1",X"38",X"01",X"EB",X"22",X"52",X"60",X"21",X"E8",X"61",X"CB",X"6E",X"C0",X"CD",X"C8",X"0F",
		X"C3",X"84",X"2E",X"21",X"00",X"90",X"3A",X"00",X"60",X"CB",X"6F",X"28",X"03",X"21",X"01",X"90",
		X"7E",X"2F",X"E6",X"05",X"C8",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"FE",X"01",X"20",X"0F",X"ED",
		X"5B",X"09",X"32",X"19",X"7C",X"FE",X"38",X"30",X"12",X"21",X"00",X"38",X"18",X"0D",X"ED",X"5B",
		X"0B",X"32",X"19",X"7C",X"FE",X"B8",X"38",X"03",X"21",X"00",X"B8",X"DD",X"75",X"04",X"DD",X"74",
		X"05",X"C9",X"78",X"E6",X"0A",X"C8",X"21",X"0D",X"32",X"FE",X"02",X"20",X"02",X"23",X"23",X"5E",
		X"23",X"56",X"DD",X"6E",X"06",X"DD",X"66",X"07",X"19",X"DD",X"75",X"06",X"DD",X"74",X"07",X"C9",
		X"DD",X"7E",X"05",X"C6",X"04",X"57",X"DD",X"7E",X"07",X"C6",X"04",X"5F",X"D5",X"CD",X"0B",X"39",
		X"D1",X"FE",X"53",X"28",X"24",X"7B",X"D6",X"08",X"5F",X"D5",X"CD",X"0B",X"39",X"D1",X"FE",X"53",
		X"28",X"17",X"7A",X"D6",X"08",X"57",X"D5",X"CD",X"0B",X"39",X"D1",X"FE",X"53",X"28",X"0A",X"7B",
		X"C6",X"08",X"5F",X"CD",X"0B",X"39",X"FE",X"53",X"C0",X"CB",X"D4",X"CB",X"5E",X"CB",X"94",X"C0",
		X"22",X"33",X"60",X"E1",X"23",X"23",X"23",X"E5",X"C9",X"2A",X"33",X"60",X"36",X"24",X"21",X"00",
		X"20",X"22",X"13",X"60",X"AF",X"32",X"12",X"60",X"CD",X"C4",X"1E",X"21",X"32",X"60",X"34",X"3E",
		X"07",X"CB",X"46",X"20",X"02",X"3E",X"08",X"CD",X"86",X"0F",X"C9",X"3A",X"55",X"60",X"82",X"CB",
		X"3F",X"CB",X"3F",X"CB",X"3F",X"E6",X"1F",X"4F",X"7B",X"ED",X"44",X"E6",X"F8",X"6F",X"26",X"00",
		X"29",X"29",X"11",X"00",X"D0",X"19",X"06",X"00",X"09",X"7E",X"C9",X"21",X"2A",X"60",X"3A",X"00",
		X"60",X"CB",X"6F",X"28",X"03",X"21",X"2B",X"60",X"7E",X"A7",X"20",X"28",X"CD",X"8C",X"3B",X"21",
		X"32",X"D1",X"06",X"08",X"11",X"EC",X"39",X"CD",X"1D",X"3A",X"06",X"B4",X"CD",X"76",X"0F",X"21",
		X"2A",X"60",X"3A",X"00",X"60",X"CB",X"6F",X"28",X"03",X"21",X"2B",X"60",X"36",X"00",X"21",X"32",
		X"D1",X"C3",X"CD",X"39",X"E5",X"21",X"52",X"D1",X"06",X"08",X"11",X"F7",X"39",X"CD",X"1D",X"3A",
		X"CD",X"2C",X"3A",X"CD",X"8C",X"3B",X"E1",X"E5",X"06",X"0A",X"CD",X"76",X"0F",X"E1",X"7E",X"3D",
		X"47",X"E6",X"0F",X"FE",X"0A",X"30",X"03",X"78",X"18",X"07",X"D6",X"06",X"4F",X"78",X"E6",X"F0",
		X"81",X"77",X"E5",X"CD",X"EF",X"3A",X"3A",X"59",X"60",X"3D",X"87",X"5F",X"16",X"00",X"21",X"93",
		X"3A",X"19",X"5E",X"23",X"56",X"EB",X"22",X"13",X"60",X"AF",X"32",X"12",X"60",X"CD",X"C4",X"1E",
		X"3E",X"0F",X"CD",X"86",X"0F",X"E1",X"7E",X"A7",X"20",X"BD",X"06",X"3C",X"CD",X"76",X"0F",X"21",
		X"B5",X"D1",X"06",X"05",X"11",X"02",X"3A",X"CD",X"1D",X"3A",X"21",X"52",X"D1",X"06",X"08",X"11",
		X"02",X"3A",X"CD",X"1D",X"3A",X"CD",X"8C",X"3B",X"3E",X"16",X"CD",X"86",X"0F",X"06",X"01",X"CD",
		X"76",X"0F",X"3A",X"1C",X"6C",X"A7",X"20",X"F5",X"C9",X"72",X"D1",X"08",X"17",X"18",X"24",X"0B",
		X"18",X"17",X"1E",X"1C",X"72",X"D1",X"08",X"24",X"24",X"24",X"0B",X"18",X"17",X"1E",X"1C",X"72",
		X"D1",X"08",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"7D",X"E6",X"E0",X"4F",X"3A",X"55",
		X"60",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"85",X"E6",X"1F",X"81",X"6F",X"C9",X"CD",X"0A",X"3A",
		X"1A",X"77",X"13",X"7D",X"3C",X"E6",X"1F",X"81",X"6F",X"10",X"F5",X"C9",X"21",X"B5",X"D1",X"CD",
		X"0A",X"3A",X"1E",X"52",X"16",X"00",X"F7",X"21",X"B6",X"D1",X"CD",X"0A",X"3A",X"1E",X"21",X"F7",
		X"CD",X"6F",X"3A",X"C5",X"21",X"B7",X"D1",X"CD",X"0A",X"3A",X"C1",X"58",X"F7",X"C5",X"21",X"B8",
		X"D1",X"CD",X"0A",X"3A",X"C1",X"59",X"F7",X"21",X"B9",X"D1",X"CD",X"0A",X"3A",X"1E",X"00",X"F7",
		X"C9",X"21",X"50",X"D3",X"1E",X"21",X"16",X"00",X"F7",X"23",X"CD",X"6F",X"3A",X"18",X"1A",X"3A",
		X"59",X"60",X"3D",X"87",X"4F",X"06",X"00",X"E5",X"21",X"93",X"3A",X"09",X"46",X"23",X"4E",X"CB",
		X"39",X"CB",X"39",X"CB",X"39",X"CB",X"39",X"E1",X"C9",X"58",X"F7",X"23",X"59",X"F7",X"23",X"1E",
		X"00",X"F7",X"C9",X"01",X"00",X"01",X"50",X"02",X"00",X"02",X"50",X"03",X"00",X"03",X"50",X"11",
		X"C2",X"3A",X"0E",X"03",X"21",X"21",X"D3",X"06",X"0F",X"1A",X"13",X"77",X"CB",X"D4",X"36",X"02",
		X"CB",X"94",X"23",X"10",X"F4",X"D5",X"11",X"11",X"00",X"19",X"D1",X"0D",X"20",X"E9",X"CD",X"61",
		X"3A",X"C9",X"40",X"43",X"43",X"43",X"43",X"43",X"43",X"43",X"43",X"43",X"45",X"43",X"43",X"43",
		X"48",X"41",X"1E",X"17",X"12",X"1F",X"0E",X"1B",X"1C",X"0A",X"15",X"46",X"24",X"24",X"24",X"49",
		X"42",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"47",X"44",X"44",X"44",X"4A",X"21",
		X"2A",X"60",X"3A",X"00",X"60",X"CB",X"6F",X"28",X"03",X"21",X"2B",X"60",X"7E",X"E5",X"CB",X"3F",
		X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"21",X"4D",X"D3",X"A7",X"28",X"11",X"16",X"00",X"1E",X"55",
		X"F7",X"23",X"1E",X"56",X"F7",X"2B",X"2B",X"C6",X"56",X"5F",X"F7",X"18",X"09",X"2B",X"36",X"24",
		X"23",X"36",X"24",X"23",X"36",X"24",X"E1",X"7E",X"08",X"7E",X"21",X"42",X"D3",X"0E",X"09",X"E6",
		X"0F",X"47",X"28",X"09",X"16",X"01",X"1E",X"52",X"F7",X"23",X"0D",X"10",X"FB",X"08",X"41",X"E6",
		X"F0",X"28",X"0A",X"78",X"A7",X"28",X"05",X"36",X"24",X"23",X"10",X"FB",X"C9",X"78",X"A7",X"28",
		X"18",X"3E",X"09",X"90",X"5F",X"16",X"00",X"E5",X"21",X"6A",X"3B",X"19",X"EB",X"E1",X"1A",X"13",
		X"D5",X"5F",X"16",X"03",X"F7",X"23",X"D1",X"10",X"F5",X"C9",X"1E",X"17",X"12",X"1F",X"0E",X"1B",
		X"1C",X"0A",X"15",X"21",X"00",X"60",X"3E",X"10",X"CB",X"7E",X"CA",X"86",X"3B",X"3E",X"20",X"CB",
		X"6E",X"CA",X"86",X"3B",X"3E",X"21",X"CD",X"98",X"3B",X"C3",X"0F",X"42",X"21",X"06",X"6C",X"01",
		X"02",X"FA",X"AF",X"D7",X"C3",X"9C",X"43",X"C9",X"C3",X"50",X"59",X"C9",X"E6",X"DD",X"7E",X"02",
		X"21",X"A4",X"3B",X"DF",X"AC",X"3B",X"AA",X"3C",X"98",X"3D",X"0D",X"3E",X"AF",X"21",X"F3",X"69",
		X"01",X"01",X"05",X"D7",X"CD",X"20",X"3E",X"DD",X"36",X"02",X"01",X"21",X"EB",X"69",X"3E",X"01",
		X"06",X"08",X"77",X"23",X"3C",X"10",X"FB",X"21",X"EB",X"69",X"3A",X"05",X"62",X"4F",X"3E",X"54",
		X"06",X"05",X"B9",X"30",X"05",X"C6",X"12",X"23",X"10",X"F8",X"36",X"FF",X"23",X"36",X"FF",X"23",
		X"36",X"FF",X"DD",X"70",X"06",X"21",X"1A",X"60",X"3A",X"00",X"60",X"CB",X"6F",X"28",X"03",X"21",
		X"21",X"60",X"7E",X"FE",X"03",X"38",X"2A",X"23",X"7E",X"FE",X"04",X"38",X"24",X"23",X"01",X"00",
		X"05",X"7E",X"A7",X"28",X"04",X"23",X"0C",X"10",X"F8",X"DD",X"5E",X"06",X"16",X"00",X"21",X"A4",
		X"3C",X"19",X"5E",X"21",X"EB",X"69",X"19",X"36",X"FF",X"06",X"00",X"21",X"F3",X"69",X"09",X"1C",
		X"73",X"06",X"05",X"11",X"F3",X"69",X"1A",X"A7",X"20",X"17",X"C5",X"06",X"00",X"CD",X"13",X"1F",
		X"7C",X"E6",X"07",X"4F",X"21",X"EB",X"69",X"09",X"7E",X"FE",X"FF",X"28",X"F0",X"C1",X"36",X"FF",
		X"12",X"13",X"10",X"E2",X"DD",X"E5",X"11",X"08",X"00",X"DD",X"19",X"FD",X"E5",X"FD",X"21",X"F3",
		X"69",X"01",X"00",X"05",X"FD",X"5E",X"00",X"1D",X"16",X"00",X"21",X"9C",X"3C",X"19",X"7E",X"DD",
		X"77",X"01",X"CD",X"31",X"0F",X"FD",X"77",X"00",X"DD",X"7E",X"01",X"CD",X"3C",X"0F",X"FD",X"96",
		X"00",X"D6",X"16",X"C5",X"57",X"1E",X"00",X"CD",X"13",X"1F",X"4D",X"06",X"00",X"CD",X"4B",X"1F",
		X"C1",X"7C",X"FD",X"86",X"00",X"C6",X"0A",X"DD",X"77",X"03",X"DD",X"71",X"04",X"0C",X"FD",X"23",
		X"11",X"06",X"00",X"DD",X"19",X"10",X"BD",X"FD",X"E1",X"DD",X"E1",X"C9",X"39",X"4B",X"5D",X"6F",
		X"81",X"93",X"A5",X"B7",X"01",X"01",X"00",X"07",X"06",X"06",X"21",X"00",X"62",X"CB",X"7E",X"CA",
		X"6A",X"3D",X"DD",X"35",X"03",X"20",X"08",X"CD",X"20",X"3E",X"DD",X"36",X"02",X"03",X"C9",X"FD",
		X"E5",X"DD",X"E5",X"DD",X"E5",X"FD",X"E1",X"11",X"04",X"00",X"DD",X"19",X"FD",X"36",X"04",X"00",
		X"FD",X"36",X"06",X"05",X"DD",X"7E",X"08",X"FE",X"FF",X"28",X"0E",X"CD",X"46",X"33",X"FE",X"0D",
		X"30",X"07",X"CD",X"53",X"33",X"FE",X"0D",X"38",X"14",X"FD",X"34",X"04",X"11",X"06",X"00",X"DD",
		X"19",X"FD",X"35",X"06",X"20",X"DE",X"DD",X"E1",X"FD",X"E1",X"C3",X"51",X"3D",X"DD",X"36",X"08",
		X"05",X"DD",X"36",X"09",X"08",X"21",X"00",X"62",X"CB",X"BE",X"21",X"E2",X"61",X"CB",X"E6",X"21",
		X"02",X"00",X"22",X"13",X"60",X"AF",X"32",X"12",X"60",X"CD",X"C4",X"1E",X"3E",X"0F",X"CD",X"86",
		X"0F",X"21",X"1C",X"60",X"3A",X"00",X"60",X"CB",X"6F",X"28",X"03",X"21",X"23",X"60",X"E5",X"FD",
		X"5E",X"04",X"16",X"00",X"19",X"7E",X"36",X"FF",X"E1",X"FE",X"FF",X"28",X"02",X"2B",X"34",X"CD",
		X"BA",X"3F",X"DD",X"E1",X"FD",X"E1",X"DD",X"36",X"05",X"0A",X"DD",X"36",X"02",X"02",X"C3",X"6A",
		X"3D",X"3E",X"08",X"DD",X"CB",X"03",X"56",X"28",X"02",X"3E",X"0D",X"DD",X"77",X"0D",X"DD",X"77",
		X"13",X"DD",X"77",X"19",X"DD",X"77",X"1F",X"DD",X"77",X"25",X"DD",X"E5",X"11",X"04",X"00",X"DD",
		X"19",X"06",X"05",X"C5",X"DD",X"7E",X"08",X"FE",X"FF",X"28",X"06",X"21",X"8C",X"3D",X"CD",X"D1",
		X"07",X"11",X"06",X"00",X"DD",X"19",X"C1",X"10",X"EA",X"DD",X"E1",X"C9",X"AC",X"01",X"B0",X"01",
		X"B4",X"01",X"B8",X"01",X"BC",X"01",X"B8",X"00",X"DD",X"35",X"05",X"C2",X"6A",X"3D",X"DD",X"7E",
		X"04",X"87",X"47",X"87",X"80",X"C6",X"08",X"5F",X"16",X"00",X"DD",X"E5",X"DD",X"19",X"DD",X"36",
		X"04",X"FF",X"DD",X"E1",X"3A",X"1B",X"60",X"21",X"00",X"60",X"CB",X"6E",X"28",X"03",X"3A",X"22",
		X"60",X"FE",X"05",X"30",X"11",X"21",X"00",X"62",X"CB",X"FE",X"21",X"E2",X"61",X"CB",X"A6",X"DD",
		X"36",X"02",X"01",X"C3",X"6A",X"3D",X"21",X"1A",X"60",X"3A",X"00",X"60",X"CB",X"6F",X"28",X"03",
		X"21",X"21",X"60",X"34",X"EF",X"DD",X"E5",X"DD",X"21",X"DF",X"61",X"CD",X"8A",X"07",X"EF",X"CD",
		X"8A",X"07",X"DD",X"E1",X"CD",X"4C",X"3E",X"21",X"00",X"62",X"CB",X"FE",X"21",X"E2",X"61",X"CB",
		X"A6",X"DD",X"E5",X"DD",X"21",X"E8",X"61",X"CD",X"17",X"26",X"DD",X"E1",X"C9",X"21",X"00",X"62",
		X"CB",X"7E",X"C8",X"DD",X"35",X"03",X"C0",X"DD",X"36",X"02",X"00",X"DD",X"36",X"03",X"3C",X"C9",
		X"21",X"1A",X"60",X"3A",X"00",X"60",X"CB",X"6F",X"28",X"03",X"21",X"21",X"60",X"7E",X"06",X"15",
		X"A7",X"28",X"08",X"06",X"12",X"FE",X"01",X"28",X"02",X"06",X"0F",X"CD",X"45",X"3E",X"4F",X"78",
		X"91",X"DD",X"77",X"03",X"C9",X"3A",X"02",X"90",X"2F",X"E6",X"03",X"C9",X"21",X"40",X"D1",X"11",
		X"05",X"69",X"CD",X"1D",X"3F",X"21",X"A0",X"D1",X"CD",X"1D",X"3F",X"21",X"00",X"D2",X"CD",X"1D",
		X"3F",X"21",X"48",X"D1",X"11",X"3D",X"3F",X"3E",X"00",X"CD",X"02",X"3F",X"21",X"A6",X"D1",X"CD",
		X"02",X"3F",X"21",X"09",X"D2",X"CD",X"02",X"3F",X"21",X"0F",X"D2",X"3E",X"01",X"CD",X"02",X"3F",
		X"21",X"14",X"D2",X"3E",X"00",X"CD",X"02",X"3F",X"DD",X"36",X"03",X"F0",X"CD",X"EB",X"3E",X"21",
		X"17",X"60",X"3A",X"00",X"60",X"CB",X"6F",X"28",X"03",X"21",X"18",X"60",X"7E",X"C6",X"01",X"27",
		X"77",X"CD",X"51",X"1E",X"3E",X"01",X"CD",X"86",X"0F",X"21",X"00",X"10",X"22",X"12",X"60",X"AF",
		X"32",X"14",X"60",X"CD",X"C4",X"1E",X"DD",X"36",X"03",X"F0",X"CD",X"EB",X"3E",X"21",X"1B",X"60",
		X"3A",X"00",X"60",X"CB",X"6F",X"28",X"03",X"21",X"22",X"60",X"AF",X"01",X"01",X"06",X"D7",X"CD",
		X"74",X"3F",X"CD",X"BA",X"3F",X"21",X"40",X"D1",X"11",X"05",X"69",X"CD",X"2D",X"3F",X"21",X"A0",
		X"D1",X"CD",X"2D",X"3F",X"21",X"00",X"D2",X"CD",X"2D",X"3F",X"C9",X"DD",X"35",X"03",X"C8",X"06",
		X"01",X"CD",X"76",X"0F",X"CD",X"74",X"3F",X"DD",X"CB",X"03",X"56",X"20",X"EE",X"CD",X"BA",X"3F",
		X"18",X"E9",X"08",X"CD",X"0A",X"3A",X"1A",X"47",X"13",X"1A",X"77",X"CB",X"D4",X"08",X"77",X"08",
		X"CB",X"94",X"13",X"7D",X"3C",X"E6",X"1F",X"81",X"6F",X"10",X"EE",X"08",X"C9",X"06",X"20",X"7E",
		X"12",X"13",X"CB",X"D4",X"7E",X"CB",X"94",X"12",X"13",X"23",X"10",X"F3",X"C9",X"06",X"20",X"1A",
		X"77",X"13",X"1A",X"CB",X"D4",X"77",X"CB",X"94",X"13",X"23",X"10",X"F3",X"C9",X"11",X"0C",X"00",
		X"17",X"10",X"1B",X"0A",X"1D",X"1E",X"15",X"0A",X"1D",X"12",X"18",X"17",X"1C",X"24",X"28",X"13",
		X"22",X"00",X"1E",X"24",X"20",X"12",X"17",X"24",X"0A",X"24",X"0E",X"21",X"1D",X"1B",X"0A",X"24",
		X"0C",X"0A",X"1B",X"06",X"0B",X"00",X"17",X"1E",X"1C",X"24",X"05",X"01",X"00",X"00",X"00",X"24",
		X"03",X"19",X"1D",X"1C",X"11",X"94",X"3F",X"0E",X"03",X"21",X"34",X"D3",X"06",X"0B",X"1A",X"13",
		X"77",X"CB",X"D4",X"36",X"03",X"CB",X"94",X"23",X"10",X"F4",X"D5",X"11",X"15",X"00",X"19",X"D1",
		X"0D",X"20",X"E9",X"C9",X"40",X"43",X"45",X"43",X"45",X"43",X"45",X"43",X"45",X"43",X"48",X"41",
		X"24",X"46",X"24",X"46",X"24",X"46",X"24",X"46",X"24",X"49",X"42",X"44",X"47",X"44",X"47",X"44",
		X"47",X"44",X"47",X"44",X"4A",X"0E",X"21",X"1D",X"1B",X"0A",X"11",X"1C",X"60",X"3A",X"00",X"60",
		X"CB",X"6F",X"28",X"03",X"11",X"23",X"60",X"06",X"05",X"21",X"55",X"D3",X"DD",X"E5",X"DD",X"21",
		X"B5",X"3F",X"DD",X"7E",X"00",X"77",X"1A",X"CB",X"D4",X"A7",X"20",X"04",X"36",X"06",X"18",X"02",
		X"36",X"01",X"CB",X"94",X"23",X"23",X"13",X"DD",X"23",X"10",X"E7",X"DD",X"E1",X"C9",X"DD",X"E5",
		X"DD",X"21",X"F8",X"69",X"DD",X"36",X"00",X"30",X"DD",X"36",X"01",X"14",X"3E",X"01",X"21",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
