library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity BASIC10 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of BASIC10 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"4C",X"59",X"EA",X"4C",X"75",X"C4",X"40",X"C9",X"A4",X"C6",X"E3",X"CF",X"E3",X"CF",X"8B",X"CC",
		X"8E",X"CC",X"DF",X"C9",X"C5",X"D9",X"15",X"DA",X"36",X"D9",X"AB",X"D8",X"F9",X"D9",X"15",X"DA",
		X"40",X"C8",X"23",X"C8",X"31",X"C8",X"0B",X"CE",X"09",X"CA",X"C8",X"CC",X"F1",X"D0",X"09",X"CC",
		X"FC",X"CC",X"D1",X"CA",X"B2",X"C9",X"8A",X"C9",X"3D",X"CA",X"1E",X"C9",X"95",X"C9",X"DF",X"C9",
		X"60",X"CA",X"5A",X"E9",X"73",X"E9",X"93",X"E9",X"A8",X"E9",X"BA",X"E9",X"14",X"F4",X"17",X"F4",
		X"1A",X"F4",X"11",X"F4",X"88",X"E8",X"88",X"E8",X"88",X"E8",X"7C",X"E8",X"7C",X"E8",X"7C",X"E8",
		X"7C",X"E8",X"7C",X"E8",X"7C",X"E8",X"7C",X"E8",X"88",X"E8",X"88",X"E8",X"3E",X"C9",X"77",X"CA",
		X"9C",X"D8",X"A9",X"E7",X"DA",X"E7",X"00",X"D4",X"93",X"D8",X"60",X"CB",X"6D",X"C9",X"72",X"C7",
		X"37",X"C7",X"B9",X"CC",X"0C",X"E8",X"88",X"CC",X"18",X"C7",X"12",X"DF",X"A5",X"DF",X"31",X"DF",
		X"21",X"00",X"D6",X"D3",X"FA",X"D3",X"17",X"D9",X"FB",X"02",X"2A",X"E2",X"4B",X"E3",X"79",X"DC",
		X"A6",X"E2",X"87",X"E3",X"8E",X"E3",X"D7",X"E3",X"3B",X"E4",X"7D",X"D8",X"C8",X"D8",X"D0",X"DD",
		X"EB",X"D7",X"D8",X"D4",X"1C",X"D8",X"FA",X"D7",X"5B",X"D7",X"EE",X"D8",X"00",X"DF",X"FC",X"DE",
		X"4F",X"DA",X"B4",X"D9",X"CD",X"E9",X"6F",X"D7",X"9B",X"D7",X"A6",X"D7",X"79",X"99",X"DA",X"79",
		X"82",X"DA",X"7B",X"B9",X"DC",X"7B",X"E2",X"DD",X"7F",X"33",X"E2",X"50",X"59",X"D0",X"46",X"56",
		X"D0",X"7D",X"6C",X"E2",X"5A",X"AF",X"CF",X"64",X"86",X"D0",X"45",X"4E",X"C4",X"45",X"44",X"49",
		X"D4",X"49",X"4E",X"56",X"45",X"52",X"53",X"C5",X"4E",X"4F",X"52",X"4D",X"41",X"CC",X"54",X"52",
		X"4F",X"CE",X"54",X"52",X"4F",X"46",X"C6",X"50",X"4F",X"D0",X"50",X"4C",X"4F",X"D4",X"50",X"55",
		X"4C",X"CC",X"4C",X"4F",X"52",X"45",X"D3",X"44",X"4F",X"4B",X"C5",X"52",X"45",X"50",X"45",X"41",
		X"D4",X"55",X"4E",X"54",X"49",X"CC",X"46",X"4F",X"D2",X"4C",X"4C",X"49",X"53",X"D4",X"4C",X"50",
		X"52",X"49",X"4E",X"D4",X"4E",X"45",X"58",X"D4",X"44",X"41",X"54",X"C1",X"49",X"4E",X"50",X"55",
		X"D4",X"44",X"49",X"CD",X"43",X"4C",X"D3",X"52",X"45",X"41",X"C4",X"4C",X"45",X"D4",X"47",X"4F",
		X"54",X"CF",X"52",X"55",X"CE",X"49",X"C6",X"52",X"45",X"53",X"54",X"4F",X"52",X"C5",X"47",X"4F",
		X"53",X"55",X"C2",X"52",X"45",X"54",X"55",X"52",X"CE",X"52",X"45",X"CD",X"48",X"49",X"4D",X"45",
		X"CD",X"47",X"52",X"41",X"C2",X"52",X"45",X"4C",X"45",X"41",X"53",X"C5",X"54",X"45",X"58",X"D4",
		X"48",X"49",X"52",X"45",X"D3",X"53",X"48",X"4F",X"4F",X"D4",X"45",X"58",X"50",X"4C",X"4F",X"44",
		X"C5",X"5A",X"41",X"D0",X"50",X"49",X"4E",X"C7",X"53",X"4F",X"55",X"4E",X"C4",X"4D",X"55",X"53",
		X"49",X"C3",X"50",X"4C",X"41",X"D9",X"43",X"55",X"52",X"53",X"45",X"D4",X"43",X"55",X"52",X"4D",
		X"4F",X"D6",X"44",X"52",X"41",X"D7",X"43",X"49",X"52",X"43",X"4C",X"C5",X"50",X"41",X"54",X"54",
		X"45",X"52",X"CE",X"46",X"49",X"4C",X"CC",X"43",X"48",X"41",X"D2",X"50",X"41",X"50",X"45",X"D2",
		X"49",X"4E",X"CB",X"53",X"54",X"4F",X"D0",X"4F",X"CE",X"57",X"41",X"49",X"D4",X"43",X"4C",X"4F",
		X"41",X"C4",X"43",X"53",X"41",X"56",X"C5",X"44",X"45",X"C6",X"50",X"4F",X"4B",X"C5",X"50",X"52",
		X"49",X"4E",X"D4",X"43",X"4F",X"4E",X"D4",X"4C",X"49",X"53",X"D4",X"43",X"4C",X"45",X"41",X"D2",
		X"47",X"45",X"D4",X"43",X"41",X"4C",X"CC",X"A1",X"4E",X"45",X"D7",X"54",X"41",X"42",X"A8",X"54",
		X"CF",X"46",X"CE",X"53",X"50",X"43",X"A8",X"C0",X"41",X"55",X"54",X"CF",X"45",X"4C",X"53",X"C5",
		X"54",X"48",X"45",X"CE",X"4E",X"4F",X"D4",X"53",X"54",X"45",X"D0",X"AB",X"AD",X"AA",X"AF",X"DE",
		X"41",X"4E",X"C4",X"4F",X"D2",X"BE",X"BD",X"BC",X"53",X"47",X"CE",X"49",X"4E",X"D4",X"41",X"42",
		X"D3",X"55",X"53",X"D2",X"46",X"52",X"C5",X"50",X"4F",X"D3",X"48",X"45",X"58",X"A4",X"A6",X"53",
		X"51",X"D2",X"52",X"4E",X"C4",X"4C",X"CE",X"45",X"58",X"D0",X"43",X"4F",X"D3",X"53",X"49",X"CE",
		X"54",X"41",X"CE",X"41",X"54",X"CE",X"50",X"45",X"45",X"CB",X"44",X"45",X"45",X"CB",X"4C",X"4F",
		X"C7",X"4C",X"45",X"CE",X"53",X"54",X"52",X"A4",X"56",X"41",X"CC",X"41",X"53",X"C3",X"43",X"48",
		X"52",X"A4",X"50",X"C9",X"54",X"52",X"55",X"C5",X"46",X"41",X"4C",X"53",X"C5",X"4B",X"45",X"59",
		X"A4",X"53",X"43",X"52",X"CE",X"50",X"4F",X"49",X"4E",X"D4",X"4C",X"45",X"46",X"54",X"A4",X"52",
		X"49",X"47",X"48",X"54",X"A4",X"4D",X"49",X"44",X"A4",X"47",X"CF",X"00",X"4E",X"45",X"58",X"54",
		X"20",X"57",X"49",X"54",X"48",X"4F",X"55",X"54",X"20",X"46",X"4F",X"D2",X"53",X"59",X"4E",X"54",
		X"41",X"D8",X"52",X"45",X"54",X"55",X"52",X"4E",X"20",X"57",X"49",X"54",X"48",X"4F",X"55",X"54",
		X"20",X"47",X"4F",X"53",X"55",X"C2",X"4F",X"55",X"54",X"20",X"4F",X"46",X"20",X"44",X"41",X"54",
		X"C1",X"49",X"4C",X"4C",X"45",X"47",X"41",X"4C",X"20",X"51",X"55",X"41",X"4E",X"54",X"49",X"54",
		X"D9",X"4F",X"56",X"45",X"52",X"46",X"4C",X"4F",X"D7",X"4F",X"55",X"54",X"20",X"4F",X"46",X"20",
		X"4D",X"45",X"4D",X"4F",X"52",X"D9",X"55",X"4E",X"44",X"45",X"46",X"27",X"44",X"20",X"53",X"54",
		X"41",X"54",X"45",X"4D",X"45",X"4E",X"D4",X"42",X"41",X"44",X"20",X"53",X"55",X"42",X"53",X"43",
		X"52",X"49",X"50",X"D4",X"52",X"45",X"44",X"49",X"4D",X"27",X"44",X"20",X"41",X"52",X"52",X"41",
		X"D9",X"44",X"49",X"56",X"49",X"53",X"49",X"4F",X"4E",X"20",X"42",X"59",X"20",X"5A",X"45",X"52",
		X"CF",X"49",X"4C",X"4C",X"45",X"47",X"41",X"4C",X"20",X"44",X"49",X"52",X"45",X"43",X"D4",X"44",
		X"49",X"53",X"50",X"20",X"54",X"59",X"50",X"45",X"20",X"4D",X"49",X"53",X"4D",X"41",X"54",X"43",
		X"C8",X"53",X"54",X"52",X"49",X"4E",X"47",X"20",X"54",X"4F",X"4F",X"20",X"4C",X"4F",X"4E",X"C7",
		X"46",X"4F",X"52",X"4D",X"55",X"4C",X"41",X"20",X"54",X"4F",X"4F",X"20",X"43",X"4F",X"4D",X"50",
		X"4C",X"45",X"D8",X"43",X"41",X"4E",X"27",X"54",X"20",X"43",X"4F",X"4E",X"54",X"49",X"4E",X"55",
		X"C5",X"55",X"4E",X"44",X"45",X"46",X"27",X"44",X"20",X"46",X"55",X"4E",X"43",X"54",X"49",X"4F",
		X"CE",X"42",X"41",X"44",X"20",X"55",X"4E",X"54",X"49",X"CC",X"20",X"45",X"52",X"52",X"4F",X"52",
		X"00",X"20",X"49",X"4E",X"20",X"00",X"0D",X"0A",X"52",X"65",X"61",X"64",X"79",X"20",X"0D",X"0A",
		X"00",X"0D",X"0A",X"20",X"42",X"52",X"45",X"41",X"4B",X"00",X"BA",X"E8",X"E8",X"E8",X"E8",X"BD",
		X"01",X"01",X"C9",X"8D",X"D0",X"21",X"A5",X"B9",X"D0",X"0A",X"BD",X"02",X"01",X"85",X"B8",X"BD",
		X"03",X"01",X"85",X"B9",X"DD",X"03",X"01",X"D0",X"07",X"A5",X"B8",X"DD",X"02",X"01",X"F0",X"07",
		X"8A",X"18",X"69",X"12",X"AA",X"D0",X"D8",X"60",X"20",X"48",X"C4",X"85",X"A0",X"84",X"A1",X"38",
		X"A5",X"C9",X"E5",X"CE",X"85",X"91",X"A8",X"A5",X"CA",X"E5",X"CF",X"AA",X"E8",X"98",X"F0",X"23",
		X"A5",X"C9",X"38",X"E5",X"91",X"85",X"C9",X"B0",X"03",X"C6",X"CA",X"38",X"A5",X"C7",X"E5",X"91",
		X"85",X"C7",X"B0",X"08",X"C6",X"C8",X"90",X"04",X"B1",X"C9",X"91",X"C7",X"88",X"D0",X"F9",X"B1",
		X"C9",X"91",X"C7",X"C6",X"CA",X"C6",X"C8",X"CA",X"D0",X"F2",X"60",X"0A",X"69",X"3E",X"B0",X"43",
		X"85",X"91",X"BA",X"E4",X"91",X"90",X"3C",X"60",X"C4",X"A3",X"90",X"28",X"D0",X"04",X"C5",X"A2",
		X"90",X"22",X"48",X"A2",X"09",X"98",X"48",X"B5",X"C6",X"CA",X"10",X"FA",X"20",X"95",X"D5",X"A2",
		X"F7",X"68",X"95",X"D0",X"E8",X"30",X"FA",X"68",X"A8",X"68",X"C4",X"A3",X"90",X"06",X"D0",X"13",
		X"C5",X"A2",X"B0",X"0F",X"60",X"AD",X"C0",X"02",X"29",X"FE",X"8D",X"C0",X"02",X"4E",X"F1",X"02",
		X"4C",X"B5",X"C4",X"A2",X"4D",X"46",X"2E",X"4E",X"F1",X"02",X"4E",X"F2",X"02",X"4E",X"F4",X"02",
		X"20",X"9F",X"CB",X"20",X"10",X"CC",X"BD",X"AC",X"C2",X"48",X"29",X"7F",X"20",X"12",X"CC",X"E8",
		X"68",X"10",X"F3",X"20",X"51",X"C7",X"A9",X"AA",X"A0",X"C3",X"20",X"ED",X"CB",X"A4",X"A9",X"C8",
		X"F0",X"03",X"20",X"B6",X"E0",X"20",X"8F",X"CC",X"46",X"2E",X"4E",X"F1",X"02",X"4E",X"F2",X"02",
		X"A9",X"B6",X"A0",X"C3",X"20",X"1A",X"00",X"4E",X"F1",X"02",X"20",X"A2",X"C5",X"86",X"E9",X"84",
		X"EA",X"20",X"E2",X"00",X"AA",X"F0",X"F0",X"A2",X"FF",X"86",X"A9",X"90",X"06",X"20",X"0A",X"C6",
		X"4C",X"DD",X"C8",X"20",X"98",X"CA",X"20",X"0A",X"C6",X"84",X"26",X"20",X"DE",X"C6",X"90",X"44",
		X"A0",X"01",X"B1",X"CE",X"85",X"92",X"A5",X"9C",X"85",X"91",X"A5",X"CF",X"85",X"94",X"A5",X"CE",
		X"88",X"F1",X"CE",X"18",X"65",X"9C",X"85",X"9C",X"85",X"93",X"A5",X"9D",X"69",X"FF",X"85",X"9D",
		X"E5",X"CF",X"AA",X"38",X"A5",X"CE",X"E5",X"9C",X"A8",X"B0",X"03",X"E8",X"C6",X"94",X"18",X"65",
		X"91",X"90",X"03",X"C6",X"92",X"18",X"B1",X"91",X"91",X"93",X"C8",X"D0",X"F9",X"E6",X"92",X"E6",
		X"94",X"CA",X"D0",X"F2",X"20",X"33",X"C7",X"20",X"6F",X"C5",X"A5",X"35",X"F0",X"89",X"18",X"A5",
		X"9C",X"85",X"C9",X"65",X"26",X"85",X"C7",X"A4",X"9D",X"84",X"CA",X"90",X"01",X"C8",X"84",X"C8",
		X"20",X"F8",X"C3",X"A5",X"A0",X"A4",X"A1",X"85",X"9C",X"84",X"9D",X"A4",X"26",X"88",X"B9",X"31",
		X"00",X"91",X"CE",X"88",X"10",X"F8",X"20",X"33",X"C7",X"20",X"6F",X"C5",X"4C",X"C7",X"C4",X"A5",
		X"9A",X"A4",X"9B",X"85",X"91",X"84",X"92",X"18",X"A0",X"01",X"B1",X"91",X"F0",X"1D",X"A0",X"04",
		X"C8",X"B1",X"91",X"D0",X"FB",X"C8",X"98",X"65",X"91",X"AA",X"A0",X"00",X"91",X"91",X"A5",X"92",
		X"69",X"00",X"C8",X"91",X"91",X"86",X"91",X"85",X"92",X"90",X"DD",X"60",X"CA",X"10",X"05",X"20",
		X"9F",X"CB",X"A2",X"00",X"20",X"F8",X"C5",X"C9",X"01",X"D0",X"0D",X"AC",X"69",X"02",X"B1",X"12",
		X"29",X"7F",X"C9",X"20",X"B0",X"02",X"A9",X"09",X"48",X"20",X"12",X"CC",X"68",X"C9",X"7F",X"F0",
		X"DB",X"C9",X"0D",X"F0",X"30",X"C9",X"03",X"F0",X"28",X"C9",X"18",X"F0",X"0B",X"C9",X"20",X"90",
		X"D3",X"95",X"35",X"E8",X"E0",X"4F",X"90",X"07",X"A9",X"5C",X"20",X"12",X"CC",X"D0",X"C0",X"E0",
		X"4C",X"90",X"C1",X"8A",X"48",X"98",X"48",X"20",X"12",X"F4",X"68",X"A8",X"68",X"AA",X"4C",X"A4",
		X"C5",X"E6",X"17",X"A2",X"00",X"4C",X"99",X"CB",X"20",X"05",X"E9",X"10",X"FB",X"C9",X"0F",X"D0",
		X"08",X"48",X"A5",X"2E",X"49",X"FF",X"85",X"2E",X"68",X"60",X"A6",X"E9",X"A0",X"04",X"84",X"2A",
		X"B5",X"00",X"C9",X"20",X"F0",X"41",X"85",X"25",X"C9",X"22",X"F0",X"5F",X"24",X"2A",X"70",X"37",
		X"C9",X"3F",X"D0",X"04",X"A9",X"BA",X"D0",X"2F",X"C9",X"30",X"90",X"04",X"C9",X"3C",X"90",X"27",
		X"84",X"E0",X"A0",X"00",X"84",X"26",X"A9",X"E9",X"85",X"18",X"A9",X"C0",X"85",X"19",X"86",X"E9",
		X"CA",X"E8",X"E6",X"18",X"D0",X"02",X"E6",X"19",X"B5",X"00",X"38",X"F1",X"18",X"F0",X"F2",X"C9",
		X"80",X"D0",X"2F",X"05",X"26",X"A4",X"E0",X"E8",X"C8",X"99",X"30",X"00",X"B9",X"30",X"00",X"F0",
		X"3C",X"38",X"E9",X"3A",X"F0",X"04",X"C9",X"57",X"D0",X"02",X"85",X"2A",X"38",X"E9",X"63",X"D0",
		X"9F",X"85",X"25",X"B5",X"00",X"F0",X"E0",X"C5",X"25",X"F0",X"DC",X"C8",X"99",X"30",X"00",X"E8",
		X"D0",X"F1",X"A6",X"E9",X"E6",X"26",X"B1",X"18",X"08",X"E6",X"18",X"D0",X"02",X"E6",X"19",X"28",
		X"10",X"F4",X"B1",X"18",X"F0",X"03",X"4C",X"48",X"C6",X"B5",X"00",X"10",X"B8",X"99",X"32",X"00",
		X"A9",X"34",X"85",X"E9",X"60",X"20",X"98",X"CA",X"20",X"DE",X"C6",X"90",X"2E",X"A9",X"80",X"8D",
		X"F2",X"02",X"A9",X"11",X"20",X"12",X"CC",X"AD",X"68",X"02",X"48",X"EA",X"EA",X"EA",X"EA",X"EA",
		X"EA",X"20",X"99",X"C7",X"68",X"8D",X"68",X"02",X"20",X"9F",X"CB",X"EA",X"EA",X"EA",X"A9",X"11",
		X"20",X"12",X"CC",X"4E",X"F2",X"02",X"68",X"68",X"4C",X"C7",X"C4",X"4C",X"F1",X"C9",X"A9",X"00",
		X"85",X"1D",X"85",X"1E",X"A5",X"9A",X"A6",X"9B",X"A0",X"01",X"85",X"CE",X"86",X"CF",X"B1",X"CE",
		X"F0",X"25",X"C8",X"C8",X"E6",X"1D",X"D0",X"02",X"E6",X"1E",X"A5",X"34",X"D1",X"CE",X"90",X"18",
		X"F0",X"03",X"88",X"D0",X"09",X"A5",X"33",X"88",X"D1",X"CE",X"90",X"0C",X"F0",X"0A",X"88",X"B1",
		X"CE",X"AA",X"88",X"B1",X"CE",X"B0",X"D1",X"18",X"60",X"D0",X"FD",X"A9",X"00",X"4E",X"F4",X"02",
		X"A8",X"91",X"9A",X"C8",X"91",X"9A",X"A5",X"9A",X"18",X"69",X"02",X"85",X"9C",X"A5",X"9B",X"69",
		X"00",X"85",X"9D",X"20",X"65",X"C7",X"A9",X"00",X"D0",X"2A",X"A5",X"A6",X"A4",X"A7",X"85",X"A2",
		X"84",X"A3",X"A5",X"9C",X"A4",X"9D",X"85",X"9E",X"84",X"9F",X"85",X"A0",X"84",X"A1",X"20",X"1F",
		X"C9",X"A2",X"88",X"86",X"85",X"68",X"A8",X"68",X"A2",X"FE",X"9A",X"48",X"98",X"48",X"A9",X"00",
		X"85",X"AD",X"85",X"2B",X"60",X"18",X"A5",X"9A",X"69",X"FF",X"85",X"E9",X"A5",X"9B",X"69",X"FF",
		X"85",X"EA",X"60",X"08",X"20",X"98",X"CA",X"20",X"DE",X"C6",X"28",X"F0",X"14",X"20",X"E8",X"00",
		X"F0",X"15",X"C9",X"CD",X"D0",X"92",X"20",X"E2",X"00",X"F0",X"06",X"20",X"98",X"CA",X"F0",X"07",
		X"60",X"A9",X"FF",X"85",X"33",X"85",X"34",X"EA",X"EA",X"A0",X"01",X"B1",X"CE",X"F0",X"47",X"20",
		X"30",X"C9",X"C9",X"20",X"D0",X"08",X"4E",X"DF",X"02",X"20",X"05",X"E9",X"10",X"FB",X"C8",X"B1",
		X"CE",X"AA",X"C8",X"B1",X"CE",X"C5",X"34",X"D0",X"04",X"E4",X"33",X"F0",X"02",X"B0",X"27",X"84",
		X"B8",X"48",X"20",X"9F",X"CB",X"68",X"20",X"C1",X"E0",X"A9",X"20",X"A4",X"B8",X"29",X"7F",X"20",
		X"12",X"CC",X"C8",X"F0",X"11",X"B1",X"CE",X"D0",X"1E",X"A8",X"B1",X"CE",X"AA",X"C8",X"B1",X"CE",
		X"86",X"CE",X"85",X"CF",X"D0",X"B3",X"2C",X"F2",X"02",X"10",X"01",X"60",X"20",X"9F",X"CB",X"4E",
		X"F1",X"02",X"68",X"68",X"4C",X"B5",X"C4",X"10",X"D6",X"38",X"E9",X"7F",X"AA",X"84",X"B8",X"A0",
		X"00",X"A9",X"E9",X"85",X"18",X"A9",X"C0",X"85",X"19",X"CA",X"F0",X"0D",X"E6",X"18",X"D0",X"02",
		X"E6",X"19",X"B1",X"18",X"10",X"F6",X"4C",X"09",X"C8",X"C8",X"B1",X"18",X"30",X"AD",X"20",X"12",
		X"CC",X"4C",X"19",X"C8",X"A9",X"80",X"8D",X"F1",X"02",X"4E",X"F2",X"02",X"20",X"E8",X"00",X"4C",
		X"73",X"C7",X"A9",X"80",X"8D",X"F1",X"02",X"20",X"E8",X"00",X"20",X"61",X"CB",X"4E",X"F1",X"02",
		X"60",X"A9",X"80",X"85",X"2B",X"20",X"D2",X"CA",X"20",X"CA",X"C3",X"D0",X"05",X"8A",X"69",X"0F",
		X"AA",X"9A",X"68",X"68",X"A9",X"09",X"20",X"3B",X"C4",X"20",X"1C",X"CA",X"18",X"98",X"65",X"E9",
		X"48",X"A5",X"EA",X"69",X"00",X"48",X"A5",X"A9",X"48",X"A5",X"A8",X"48",X"A9",X"C3",X"20",X"DB",
		X"CF",X"20",X"7A",X"CE",X"20",X"77",X"CE",X"A5",X"D5",X"09",X"7F",X"25",X"D1",X"85",X"D1",X"A9",
		X"8A",X"A0",X"C8",X"85",X"91",X"84",X"92",X"4C",X"34",X"CF",X"A9",X"4B",X"A0",X"DC",X"20",X"73",
		X"DE",X"20",X"E8",X"00",X"C9",X"CB",X"D0",X"06",X"20",X"E2",X"00",X"20",X"77",X"CE",X"20",X"04",
		X"DF",X"20",X"25",X"CF",X"A5",X"B9",X"48",X"A5",X"B8",X"48",X"A9",X"8D",X"48",X"20",X"30",X"C9",
		X"A5",X"E9",X"A4",X"EA",X"F0",X"06",X"85",X"AC",X"84",X"AD",X"A0",X"00",X"B1",X"E9",X"D0",X"58",
		X"A0",X"02",X"B1",X"E9",X"18",X"D0",X"03",X"4C",X"58",X"C9",X"C8",X"B1",X"E9",X"85",X"A8",X"C8",
		X"B1",X"E9",X"85",X"A9",X"98",X"65",X"E9",X"85",X"E9",X"90",X"02",X"E6",X"EA",X"2C",X"F4",X"02",
		X"10",X"13",X"48",X"A9",X"5B",X"20",X"4D",X"CC",X"A5",X"A9",X"A6",X"A8",X"20",X"C1",X"E0",X"A9",
		X"5D",X"20",X"4D",X"CC",X"68",X"20",X"E2",X"00",X"20",X"FE",X"C8",X"4C",X"AD",X"C8",X"F0",X"2D",
		X"E9",X"80",X"90",X"11",X"C9",X"42",X"B0",X"14",X"0A",X"A8",X"B9",X"07",X"C0",X"48",X"B9",X"06",
		X"C0",X"48",X"4C",X"E2",X"00",X"4C",X"D2",X"CA",X"C9",X"3A",X"F0",X"C1",X"4C",X"E4",X"CF",X"38",
		X"A5",X"9A",X"E9",X"01",X"A4",X"9B",X"B0",X"01",X"88",X"85",X"B0",X"84",X"B1",X"60",X"EA",X"60",
		X"AD",X"DF",X"02",X"10",X"F9",X"29",X"7F",X"A2",X"08",X"C9",X"03",X"D0",X"F1",X"C9",X"03",X"B0",
		X"01",X"18",X"D0",X"43",X"A5",X"E9",X"A4",X"EA",X"F0",X"0C",X"85",X"AC",X"84",X"AD",X"A5",X"A8",
		X"A4",X"A9",X"85",X"AA",X"84",X"AB",X"68",X"68",X"A9",X"C1",X"A0",X"C3",X"A2",X"00",X"8E",X"F1",
		X"02",X"8E",X"DF",X"02",X"86",X"2E",X"90",X"03",X"4C",X"AA",X"C4",X"4C",X"B5",X"C4",X"D0",X"17",
		X"A2",X"D7",X"A4",X"AD",X"D0",X"03",X"4C",X"85",X"C4",X"A5",X"AC",X"85",X"E9",X"84",X"EA",X"A5",
		X"AA",X"A4",X"AB",X"85",X"A8",X"84",X"A9",X"60",X"4C",X"A0",X"D2",X"D0",X"03",X"4C",X"33",X"C7",
		X"20",X"3A",X"C7",X"4C",X"AA",X"C9",X"A9",X"03",X"20",X"3B",X"C4",X"A5",X"EA",X"48",X"A5",X"E9",
		X"48",X"A5",X"A9",X"48",X"A5",X"A8",X"48",X"A9",X"9B",X"48",X"20",X"E8",X"00",X"20",X"B3",X"C9",
		X"4C",X"AD",X"C8",X"20",X"9D",X"E7",X"20",X"1F",X"CA",X"A5",X"A9",X"C5",X"34",X"B0",X"0B",X"98",
		X"38",X"65",X"E9",X"A6",X"EA",X"90",X"07",X"E8",X"B0",X"04",X"A5",X"9A",X"A6",X"9B",X"20",X"E8",
		X"C6",X"90",X"1E",X"A5",X"CE",X"E9",X"01",X"85",X"E9",X"A5",X"CF",X"E9",X"00",X"85",X"EA",X"60",
		X"D0",X"FD",X"A9",X"FF",X"85",X"B9",X"20",X"CA",X"C3",X"9A",X"C9",X"9B",X"F0",X"0B",X"A2",X"16",
		X"2C",X"A2",X"5A",X"4C",X"85",X"C4",X"4C",X"E4",X"CF",X"68",X"68",X"C0",X"0C",X"F0",X"19",X"85",
		X"A8",X"68",X"85",X"A9",X"68",X"85",X"E9",X"68",X"85",X"EA",X"20",X"1C",X"CA",X"98",X"18",X"65",
		X"E9",X"85",X"E9",X"90",X"02",X"E6",X"EA",X"60",X"68",X"68",X"68",X"60",X"A2",X"3A",X"2C",X"A2",
		X"00",X"86",X"24",X"A0",X"00",X"84",X"25",X"A5",X"25",X"A6",X"24",X"85",X"24",X"86",X"25",X"B1",
		X"E9",X"F0",X"E4",X"C5",X"25",X"F0",X"E0",X"C8",X"C9",X"22",X"D0",X"F3",X"F0",X"E9",X"20",X"8B",
		X"CE",X"20",X"E8",X"00",X"C9",X"97",X"F0",X"05",X"A9",X"C9",X"20",X"DB",X"CF",X"A5",X"D0",X"D0",
		X"05",X"20",X"66",X"CA",X"F0",X"B7",X"20",X"E8",X"00",X"B0",X"03",X"4C",X"B3",X"C9",X"4C",X"FE",
		X"C8",X"20",X"1F",X"CA",X"F0",X"A7",X"A0",X"00",X"B1",X"E9",X"F0",X"08",X"C8",X"C9",X"C8",X"D0",
		X"F7",X"4C",X"0D",X"CA",X"60",X"4C",X"E4",X"CF",X"20",X"0D",X"D8",X"48",X"C9",X"9B",X"F0",X"04",
		X"C9",X"97",X"D0",X"F1",X"C6",X"D4",X"D0",X"04",X"68",X"4C",X"00",X"C9",X"20",X"E2",X"00",X"20",
		X"98",X"CA",X"C9",X"2C",X"F0",X"EE",X"68",X"60",X"A2",X"00",X"86",X"33",X"86",X"34",X"B0",X"F7",
		X"E9",X"2F",X"85",X"24",X"A5",X"34",X"85",X"91",X"C9",X"19",X"B0",X"D4",X"A5",X"33",X"0A",X"26",
		X"91",X"0A",X"26",X"91",X"65",X"33",X"85",X"33",X"A5",X"91",X"65",X"34",X"85",X"34",X"06",X"33",
		X"26",X"34",X"A5",X"33",X"65",X"24",X"85",X"33",X"90",X"02",X"E6",X"34",X"20",X"E2",X"00",X"4C",
		X"9E",X"CA",X"20",X"FC",X"D0",X"85",X"B8",X"84",X"B9",X"A9",X"D4",X"20",X"DB",X"CF",X"A5",X"29",
		X"48",X"A5",X"28",X"48",X"20",X"8B",X"CE",X"68",X"2A",X"20",X"7D",X"CE",X"D0",X"18",X"68",X"10",
		X"12",X"20",X"EC",X"DE",X"20",X"17",X"D2",X"A0",X"00",X"A5",X"D3",X"91",X"B8",X"C8",X"A5",X"D4",
		X"91",X"B8",X"60",X"4C",X"A1",X"DE",X"68",X"A0",X"02",X"B1",X"D3",X"C5",X"A3",X"90",X"17",X"D0",
		X"07",X"88",X"B1",X"D3",X"C5",X"A2",X"90",X"0E",X"A4",X"D4",X"C4",X"9D",X"90",X"08",X"D0",X"0D",
		X"A5",X"D3",X"C5",X"9C",X"B0",X"07",X"A5",X"D3",X"A4",X"D4",X"4C",X"43",X"CB",X"A0",X"00",X"B1",
		X"D3",X"20",X"E8",X"D4",X"A5",X"BF",X"A4",X"C0",X"85",X"DE",X"84",X"DF",X"20",X"E9",X"D6",X"A9",
		X"D0",X"A0",X"00",X"85",X"BF",X"84",X"C0",X"20",X"4A",X"D7",X"A0",X"00",X"B1",X"BF",X"91",X"B8",
		X"C8",X"B1",X"BF",X"91",X"B8",X"C8",X"B1",X"BF",X"91",X"B8",X"60",X"20",X"F0",X"CB",X"20",X"E8",
		X"00",X"F0",X"3C",X"F0",X"46",X"C9",X"C2",X"F0",X"61",X"C9",X"C5",X"18",X"F0",X"5C",X"C9",X"2C",
		X"F0",X"3A",X"C9",X"3B",X"F0",X"69",X"20",X"8B",X"CE",X"24",X"28",X"30",X"DE",X"20",X"D1",X"E0",
		X"20",X"FA",X"D4",X"A0",X"00",X"B1",X"D3",X"18",X"65",X"30",X"C5",X"31",X"90",X"03",X"20",X"9F",
		X"CB",X"20",X"F0",X"CB",X"20",X"0D",X"CC",X"D0",X"C5",X"A0",X"00",X"94",X"35",X"A2",X"34",X"A9",
		X"0D",X"85",X"30",X"20",X"12",X"CC",X"A9",X"0A",X"20",X"12",X"CC",X"60",X"EA",X"EA",X"EA",X"EA",
		X"EA",X"EA",X"EA",X"A5",X"30",X"C5",X"32",X"90",X"06",X"20",X"9F",X"CB",X"4C",X"DF",X"CB",X"38",
		X"E9",X"08",X"B0",X"FC",X"49",X"FF",X"69",X"01",X"D0",X"10",X"08",X"20",X"0A",X"D8",X"C9",X"29",
		X"D0",X"18",X"28",X"90",X"06",X"8A",X"E5",X"30",X"90",X"05",X"AA",X"E8",X"CA",X"D0",X"06",X"20",
		X"E2",X"00",X"4C",X"63",X"CB",X"20",X"0D",X"CC",X"D0",X"F2",X"4C",X"E4",X"CF",X"20",X"FA",X"D4",
		X"20",X"15",X"D7",X"AA",X"A0",X"00",X"E8",X"CA",X"F0",X"B1",X"B1",X"91",X"20",X"12",X"CC",X"C8",
		X"C9",X"0D",X"D0",X"F3",X"20",X"AB",X"CB",X"4C",X"F7",X"CB",X"A9",X"0C",X"2C",X"A9",X"20",X"2C",
		X"A9",X"3F",X"24",X"2E",X"30",X"54",X"2C",X"F1",X"02",X"10",X"32",X"48",X"C9",X"20",X"90",X"0B",
		X"A5",X"30",X"C5",X"31",X"D0",X"03",X"20",X"9F",X"CB",X"E6",X"30",X"68",X"85",X"27",X"8A",X"48",
		X"98",X"48",X"A5",X"27",X"20",X"33",X"F4",X"AA",X"10",X"0A",X"A9",X"6D",X"A0",X"CC",X"4E",X"F1",
		X"02",X"20",X"ED",X"CB",X"68",X"A8",X"68",X"AA",X"A5",X"27",X"29",X"FF",X"60",X"85",X"27",X"98",
		X"48",X"8A",X"48",X"A5",X"27",X"C9",X"20",X"90",X"07",X"A8",X"C8",X"30",X"03",X"0D",X"F7",X"02",
		X"AA",X"20",X"09",X"F4",X"68",X"AA",X"68",X"A8",X"A5",X"27",X"29",X"FF",X"60",X"0D",X"0A",X"3F",
		X"50",X"52",X"49",X"4E",X"54",X"45",X"52",X"20",X"45",X"52",X"52",X"4F",X"52",X"0D",X"0A",X"00",
		X"A9",X"80",X"2C",X"A9",X"00",X"8D",X"F7",X"02",X"60",X"6C",X"F5",X"02",X"A9",X"80",X"2C",X"A9",
		X"00",X"8D",X"F4",X"02",X"60",X"A5",X"2C",X"F0",X"11",X"30",X"04",X"A0",X"FF",X"D0",X"04",X"A5",
		X"AE",X"A4",X"AF",X"85",X"A8",X"84",X"A9",X"4C",X"E4",X"CF",X"A9",X"F9",X"A0",X"CD",X"20",X"ED",
		X"CB",X"A5",X"AC",X"A4",X"AD",X"85",X"E9",X"84",X"EA",X"60",X"20",X"19",X"D4",X"A2",X"36",X"A0",
		X"00",X"84",X"36",X"A9",X"40",X"20",X"03",X"CD",X"60",X"46",X"2E",X"C9",X"22",X"D0",X"0B",X"20",
		X"99",X"CF",X"A9",X"3B",X"20",X"DB",X"CF",X"20",X"F0",X"CB",X"20",X"19",X"D4",X"A9",X"2C",X"85",
		X"34",X"A9",X"00",X"85",X"17",X"20",X"F4",X"CC",X"A5",X"35",X"D0",X"16",X"A5",X"17",X"F0",X"F1",
		X"18",X"4C",X"4E",X"C9",X"20",X"10",X"CC",X"20",X"0D",X"CC",X"4C",X"A2",X"C5",X"A6",X"B0",X"A4",
		X"B1",X"A9",X"98",X"85",X"2C",X"86",X"B2",X"84",X"B3",X"20",X"FC",X"D0",X"85",X"B8",X"84",X"B9",
		X"A5",X"E9",X"A4",X"EA",X"85",X"BA",X"84",X"BB",X"A6",X"B2",X"A4",X"B3",X"86",X"E9",X"84",X"EA",
		X"20",X"E8",X"00",X"D0",X"1D",X"24",X"2C",X"50",X"0D",X"20",X"05",X"E9",X"10",X"FB",X"85",X"35",
		X"A2",X"34",X"A0",X"00",X"F0",X"08",X"30",X"71",X"20",X"10",X"CC",X"20",X"F4",X"CC",X"86",X"E9",
		X"84",X"EA",X"20",X"E2",X"00",X"24",X"28",X"10",X"31",X"24",X"2C",X"50",X"09",X"E8",X"86",X"E9",
		X"A9",X"00",X"85",X"24",X"F0",X"0C",X"85",X"24",X"C9",X"22",X"F0",X"07",X"A9",X"3A",X"85",X"24",
		X"A9",X"2C",X"18",X"85",X"25",X"A5",X"E9",X"A4",X"EA",X"69",X"00",X"90",X"01",X"C8",X"20",X"00",
		X"D5",X"20",X"52",X"D8",X"20",X"07",X"CB",X"4C",X"82",X"CD",X"20",X"CF",X"DF",X"A5",X"29",X"20",
		X"EF",X"CA",X"20",X"E8",X"00",X"F0",X"07",X"C9",X"2C",X"F0",X"03",X"4C",X"95",X"CC",X"A5",X"E9",
		X"A4",X"EA",X"85",X"B2",X"84",X"B3",X"A5",X"BA",X"A4",X"BB",X"85",X"E9",X"84",X"EA",X"20",X"E8",
		X"00",X"F0",X"2C",X"20",X"D9",X"CF",X"4C",X"09",X"CD",X"20",X"1C",X"CA",X"C8",X"AA",X"D0",X"12",
		X"A2",X"2A",X"C8",X"B1",X"E9",X"F0",X"69",X"C8",X"B1",X"E9",X"85",X"AE",X"C8",X"B1",X"E9",X"C8",
		X"85",X"AF",X"B1",X"E9",X"AA",X"20",X"0D",X"CA",X"E0",X"91",X"D0",X"DD",X"4C",X"42",X"CD",X"A5",
		X"B2",X"A4",X"B3",X"A6",X"2C",X"10",X"03",X"4C",X"29",X"C9",X"A0",X"00",X"B1",X"B2",X"F0",X"07",
		X"A9",X"E8",X"A0",X"CD",X"4C",X"ED",X"CB",X"60",X"3F",X"45",X"58",X"54",X"52",X"41",X"20",X"49",
		X"47",X"4E",X"4F",X"52",X"45",X"44",X"0D",X"0A",X"00",X"3F",X"52",X"45",X"44",X"4F",X"20",X"46",
		X"52",X"4F",X"4D",X"20",X"53",X"54",X"41",X"52",X"54",X"0D",X"0A",X"00",X"D0",X"04",X"A0",X"00",
		X"F0",X"03",X"20",X"FC",X"D0",X"85",X"B8",X"84",X"B9",X"20",X"CA",X"C3",X"F0",X"04",X"A2",X"00",
		X"F0",X"66",X"9A",X"8A",X"18",X"69",X"04",X"48",X"69",X"06",X"85",X"93",X"68",X"A0",X"01",X"20",
		X"73",X"DE",X"BA",X"BD",X"09",X"01",X"85",X"D5",X"A5",X"B8",X"A4",X"B9",X"20",X"97",X"DA",X"20",
		X"A1",X"DE",X"A0",X"01",X"20",X"36",X"DF",X"BA",X"38",X"FD",X"09",X"01",X"F0",X"17",X"BD",X"0F",
		X"01",X"85",X"A8",X"BD",X"10",X"01",X"85",X"A9",X"BD",X"12",X"01",X"85",X"E9",X"BD",X"11",X"01",
		X"85",X"EA",X"4C",X"AD",X"C8",X"8A",X"69",X"11",X"AA",X"9A",X"20",X"E8",X"00",X"C9",X"2C",X"D0",
		X"F1",X"20",X"E2",X"00",X"20",X"12",X"CE",X"20",X"8B",X"CE",X"18",X"24",X"38",X"24",X"28",X"30",
		X"03",X"B0",X"03",X"60",X"B0",X"FD",X"A2",X"A8",X"4C",X"85",X"C4",X"A6",X"E9",X"D0",X"02",X"C6",
		X"EA",X"C6",X"E9",X"A2",X"00",X"24",X"48",X"8A",X"48",X"A9",X"01",X"20",X"3B",X"C4",X"20",X"74",
		X"CF",X"A9",X"00",X"85",X"BC",X"20",X"E8",X"00",X"38",X"E9",X"D3",X"90",X"17",X"C9",X"03",X"B0",
		X"13",X"C9",X"01",X"2A",X"49",X"01",X"45",X"BC",X"C5",X"BC",X"90",X"61",X"85",X"BC",X"20",X"E2",
		X"00",X"4C",X"A8",X"CE",X"A6",X"BC",X"D0",X"2C",X"B0",X"7F",X"69",X"07",X"90",X"7B",X"65",X"28",
		X"D0",X"03",X"4C",X"AC",X"D6",X"69",X"FF",X"85",X"91",X"0A",X"65",X"91",X"A8",X"68",X"D9",X"CC",
		X"C0",X"B0",X"6B",X"20",X"7A",X"CE",X"48",X"20",X"0D",X"CF",X"68",X"A4",X"BA",X"10",X"17",X"AA",
		X"F0",X"5A",X"D0",X"63",X"46",X"28",X"8A",X"2A",X"A6",X"E9",X"D0",X"02",X"C6",X"EA",X"C6",X"E9",
		X"A0",X"1B",X"85",X"BC",X"D0",X"D7",X"D9",X"CC",X"C0",X"B0",X"4C",X"90",X"D9",X"B9",X"CE",X"C0",
		X"48",X"B9",X"CD",X"C0",X"48",X"20",X"20",X"CF",X"A5",X"BC",X"4C",X"96",X"CE",X"4C",X"E4",X"CF",
		X"A5",X"D5",X"BE",X"CC",X"C0",X"A8",X"68",X"85",X"91",X"68",X"85",X"92",X"E6",X"91",X"D0",X"02",
		X"E6",X"92",X"98",X"48",X"20",X"EC",X"DE",X"A5",X"D4",X"48",X"A5",X"D3",X"48",X"A5",X"D2",X"48",
		X"A5",X"D1",X"48",X"A5",X"D0",X"48",X"6C",X"91",X"00",X"A0",X"FF",X"68",X"F0",X"23",X"C9",X"64",
		X"F0",X"03",X"20",X"7A",X"CE",X"84",X"BA",X"68",X"4A",X"85",X"2D",X"68",X"85",X"D8",X"68",X"85",
		X"D9",X"68",X"85",X"DA",X"68",X"85",X"DB",X"68",X"85",X"DC",X"68",X"85",X"DD",X"45",X"D5",X"85",
		X"DE",X"A5",X"D0",X"60",X"A9",X"00",X"85",X"28",X"20",X"E2",X"00",X"B0",X"03",X"4C",X"CF",X"DF",
		X"20",X"86",X"D1",X"B0",X"6B",X"C9",X"2E",X"F0",X"F4",X"C9",X"23",X"F0",X"F0",X"C9",X"CD",X"F0",
		X"58",X"C9",X"CC",X"F0",X"E3",X"C9",X"22",X"D0",X"0F",X"A5",X"E9",X"A4",X"EA",X"69",X"00",X"90",
		X"01",X"C8",X"20",X"FA",X"D4",X"4C",X"52",X"D8",X"C9",X"CA",X"D0",X"13",X"A0",X"18",X"D0",X"3B",
		X"20",X"17",X"D2",X"A5",X"D4",X"49",X"FF",X"A8",X"A5",X"D3",X"49",X"FF",X"4C",X"ED",X"D3",X"C9",
		X"C4",X"D0",X"03",X"4C",X"67",X"D4",X"C9",X"D6",X"90",X"03",X"4C",X"14",X"D0",X"20",X"D6",X"CF",
		X"20",X"8B",X"CE",X"A9",X"29",X"2C",X"A9",X"28",X"2C",X"A9",X"2C",X"A0",X"00",X"D1",X"E9",X"D0",
		X"03",X"4C",X"E2",X"00",X"A2",X"10",X"4C",X"85",X"C4",X"A0",X"15",X"68",X"68",X"4C",X"E7",X"CE",
		X"20",X"FC",X"D0",X"85",X"D3",X"84",X"D4",X"A6",X"28",X"F0",X"05",X"A2",X"00",X"86",X"DF",X"60",
		X"A6",X"29",X"10",X"0D",X"A0",X"00",X"B1",X"D3",X"AA",X"C8",X"B1",X"D3",X"A8",X"8A",X"4C",X"ED",
		X"D3",X"4C",X"73",X"DE",X"0A",X"48",X"AA",X"20",X"E2",X"00",X"E0",X"DB",X"90",X"24",X"E0",X"E7",
		X"90",X"23",X"20",X"D6",X"CF",X"20",X"8B",X"CE",X"20",X"D9",X"CF",X"20",X"7C",X"CE",X"68",X"AA",
		X"A5",X"D4",X"48",X"A5",X"D3",X"48",X"8A",X"48",X"20",X"0D",X"D8",X"68",X"A8",X"8A",X"48",X"4C",
		X"47",X"D0",X"20",X"CD",X"CF",X"68",X"A8",X"B9",X"DE",X"BF",X"85",X"C4",X"B9",X"DF",X"BF",X"85",
		X"C5",X"20",X"C3",X"00",X"4C",X"7A",X"CE",X"A0",X"FF",X"2C",X"A0",X"00",X"84",X"26",X"20",X"17",
		X"D2",X"A5",X"D3",X"45",X"26",X"85",X"24",X"A5",X"D4",X"45",X"26",X"85",X"25",X"20",X"CD",X"DE",
		X"20",X"17",X"D2",X"A5",X"D4",X"45",X"26",X"25",X"25",X"45",X"26",X"A8",X"A5",X"D3",X"45",X"26",
		X"25",X"24",X"45",X"26",X"4C",X"ED",X"D3",X"20",X"7D",X"CE",X"B0",X"13",X"A5",X"DD",X"09",X"7F",
		X"25",X"D9",X"85",X"D9",X"A9",X"D8",X"A0",X"00",X"20",X"34",X"DF",X"AA",X"4C",X"D2",X"D0",X"A9",
		X"00",X"85",X"28",X"C6",X"BC",X"20",X"15",X"D7",X"85",X"D0",X"86",X"D1",X"84",X"D2",X"A5",X"DB",
		X"A4",X"DC",X"20",X"19",X"D7",X"86",X"DB",X"84",X"DC",X"AA",X"38",X"E5",X"D0",X"F0",X"08",X"A9",
		X"01",X"90",X"04",X"A6",X"D0",X"A9",X"FF",X"85",X"D5",X"A0",X"FF",X"E8",X"C8",X"CA",X"D0",X"07",
		X"A6",X"D5",X"30",X"0F",X"18",X"90",X"0C",X"B1",X"DB",X"D1",X"D1",X"F0",X"EF",X"A2",X"FF",X"B0",
		X"02",X"A2",X"01",X"E8",X"8A",X"2A",X"25",X"2D",X"F0",X"02",X"A9",X"FF",X"4C",X"15",X"DF",X"20",
		X"D9",X"CF",X"AA",X"20",X"01",X"D1",X"20",X"E8",X"00",X"D0",X"F4",X"60",X"A2",X"00",X"20",X"E8",
		X"00",X"86",X"27",X"85",X"B4",X"20",X"E8",X"00",X"20",X"86",X"D1",X"B0",X"03",X"4C",X"E4",X"CF",
		X"A2",X"00",X"86",X"28",X"86",X"29",X"20",X"E2",X"00",X"90",X"05",X"20",X"86",X"D1",X"90",X"0B",
		X"AA",X"20",X"E2",X"00",X"90",X"FB",X"20",X"86",X"D1",X"B0",X"F6",X"C9",X"24",X"D0",X"06",X"A9",
		X"FF",X"85",X"28",X"D0",X"10",X"C9",X"25",X"D0",X"13",X"A5",X"2B",X"D0",X"D0",X"A9",X"80",X"85",
		X"29",X"05",X"B4",X"85",X"B4",X"8A",X"09",X"80",X"AA",X"20",X"E2",X"00",X"86",X"B5",X"38",X"05",
		X"2B",X"E9",X"28",X"D0",X"03",X"4C",X"29",X"D2",X"A9",X"00",X"85",X"2B",X"A5",X"9C",X"A6",X"9D",
		X"A0",X"00",X"86",X"CF",X"85",X"CE",X"E4",X"9F",X"D0",X"04",X"C5",X"9E",X"F0",X"22",X"A5",X"B4",
		X"D1",X"CE",X"D0",X"08",X"A5",X"B5",X"C8",X"D1",X"CE",X"F0",X"6A",X"88",X"18",X"A5",X"CE",X"69",
		X"07",X"90",X"E1",X"E8",X"D0",X"DC",X"C9",X"41",X"90",X"05",X"E9",X"5B",X"38",X"E9",X"A5",X"60",
		X"68",X"48",X"C9",X"F2",X"D0",X"0D",X"BA",X"BD",X"02",X"01",X"C9",X"CF",X"D0",X"05",X"A9",X"03",
		X"A0",X"E2",X"60",X"A5",X"9E",X"A4",X"9F",X"85",X"CE",X"84",X"CF",X"A5",X"A0",X"A4",X"A1",X"85",
		X"C9",X"84",X"CA",X"18",X"69",X"07",X"90",X"01",X"C8",X"85",X"C7",X"84",X"C8",X"20",X"F8",X"C3",
		X"A5",X"C7",X"A4",X"C8",X"C8",X"85",X"9E",X"84",X"9F",X"A0",X"00",X"A5",X"B4",X"91",X"CE",X"C8",
		X"A5",X"B5",X"91",X"CE",X"A9",X"00",X"C8",X"91",X"CE",X"C8",X"91",X"CE",X"C8",X"91",X"CE",X"C8",
		X"91",X"CE",X"C8",X"91",X"CE",X"A5",X"CE",X"18",X"69",X"02",X"A4",X"CF",X"90",X"01",X"C8",X"85",
		X"B6",X"84",X"B7",X"60",X"A5",X"26",X"0A",X"69",X"05",X"65",X"CE",X"A4",X"CF",X"90",X"01",X"C8",
		X"85",X"C7",X"84",X"C8",X"60",X"90",X"80",X"00",X"00",X"00",X"20",X"E2",X"00",X"20",X"8B",X"CE",
		X"20",X"7A",X"CE",X"A5",X"D5",X"30",X"0D",X"A5",X"D0",X"C9",X"90",X"90",X"09",X"A9",X"05",X"A0",
		X"D2",X"20",X"34",X"DF",X"D0",X"7A",X"4C",X"74",X"DF",X"A5",X"27",X"05",X"29",X"48",X"A5",X"28",
		X"48",X"A0",X"00",X"98",X"48",X"A5",X"B5",X"48",X"A5",X"B4",X"48",X"20",X"0A",X"D2",X"68",X"85",
		X"B4",X"68",X"85",X"B5",X"68",X"A8",X"BA",X"BD",X"02",X"01",X"48",X"BD",X"01",X"01",X"48",X"A5",
		X"D3",X"9D",X"02",X"01",X"A5",X"D4",X"9D",X"01",X"01",X"C8",X"20",X"E8",X"00",X"C9",X"2C",X"F0",
		X"D2",X"84",X"26",X"20",X"D3",X"CF",X"68",X"85",X"28",X"68",X"85",X"29",X"29",X"7F",X"85",X"27",
		X"A6",X"9E",X"A5",X"9F",X"86",X"CE",X"85",X"CF",X"C5",X"A1",X"D0",X"04",X"E4",X"A0",X"F0",X"39",
		X"A0",X"00",X"B1",X"CE",X"C8",X"C5",X"B4",X"D0",X"06",X"A5",X"B5",X"D1",X"CE",X"F0",X"16",X"C8",
		X"B1",X"CE",X"18",X"65",X"CE",X"AA",X"C8",X"B1",X"CE",X"65",X"CF",X"90",X"D7",X"A2",X"6B",X"2C",
		X"A2",X"35",X"4C",X"85",X"C4",X"A2",X"78",X"A5",X"27",X"D0",X"F7",X"20",X"F4",X"D1",X"A5",X"26",
		X"A0",X"04",X"D1",X"CE",X"D0",X"E7",X"4C",X"43",X"D3",X"20",X"F4",X"D1",X"20",X"48",X"C4",X"A9",
		X"00",X"A8",X"85",X"E1",X"A2",X"05",X"A5",X"B4",X"91",X"CE",X"10",X"01",X"CA",X"C8",X"A5",X"B5",
		X"91",X"CE",X"10",X"02",X"CA",X"CA",X"86",X"E0",X"A5",X"26",X"C8",X"C8",X"C8",X"91",X"CE",X"A2",
		X"0B",X"A9",X"00",X"24",X"27",X"50",X"08",X"68",X"18",X"69",X"01",X"AA",X"68",X"69",X"00",X"C8",
		X"91",X"CE",X"C8",X"8A",X"91",X"CE",X"20",X"A5",X"D3",X"86",X"E0",X"85",X"E1",X"A4",X"91",X"C6",
		X"26",X"D0",X"DC",X"65",X"C8",X"B0",X"5D",X"85",X"C8",X"A8",X"8A",X"65",X"C7",X"90",X"03",X"C8",
		X"F0",X"52",X"20",X"48",X"C4",X"85",X"A0",X"84",X"A1",X"A9",X"00",X"E6",X"E1",X"A4",X"E0",X"F0",
		X"05",X"88",X"91",X"C7",X"D0",X"FB",X"C6",X"C8",X"C6",X"E1",X"D0",X"F5",X"E6",X"C8",X"38",X"A5",
		X"A0",X"E5",X"CE",X"A0",X"02",X"91",X"CE",X"A5",X"A1",X"C8",X"E5",X"CF",X"91",X"CE",X"A5",X"27",
		X"D0",X"62",X"C8",X"B1",X"CE",X"85",X"26",X"A9",X"00",X"85",X"E0",X"85",X"E1",X"C8",X"68",X"AA",
		X"85",X"D3",X"68",X"85",X"D4",X"D1",X"CE",X"90",X"0E",X"D0",X"06",X"C8",X"8A",X"D1",X"CE",X"90",
		X"07",X"4C",X"9D",X"D2",X"4C",X"83",X"C4",X"C8",X"A5",X"E1",X"05",X"E0",X"18",X"F0",X"0A",X"20",
		X"A5",X"D3",X"8A",X"65",X"D3",X"AA",X"98",X"A4",X"91",X"65",X"D4",X"86",X"E0",X"C6",X"26",X"D0",
		X"CA",X"85",X"E1",X"A2",X"05",X"A5",X"B4",X"10",X"01",X"CA",X"A5",X"B5",X"10",X"02",X"CA",X"CA",
		X"86",X"97",X"A9",X"00",X"20",X"AE",X"D3",X"8A",X"65",X"C7",X"85",X"B6",X"98",X"65",X"C8",X"85",
		X"B7",X"A8",X"A5",X"B6",X"60",X"84",X"91",X"B1",X"CE",X"85",X"97",X"88",X"B1",X"CE",X"85",X"98",
		X"A9",X"10",X"85",X"CC",X"A2",X"00",X"A0",X"00",X"8A",X"0A",X"AA",X"98",X"2A",X"A8",X"B0",X"A4",
		X"06",X"E0",X"26",X"E1",X"90",X"0B",X"18",X"8A",X"65",X"97",X"AA",X"98",X"65",X"98",X"A8",X"B0",
		X"93",X"C6",X"CC",X"D0",X"E3",X"60",X"A5",X"28",X"F0",X"03",X"20",X"15",X"D7",X"20",X"95",X"D5",
		X"38",X"A5",X"A2",X"E5",X"A0",X"A8",X"A5",X"A3",X"E5",X"A1",X"4C",X"D5",X"D8",X"A2",X"00",X"86",
		X"28",X"85",X"D1",X"84",X"D2",X"A2",X"90",X"4C",X"1D",X"DF",X"AC",X"69",X"02",X"A9",X"00",X"F0",
		X"EC",X"C9",X"D9",X"D0",X"21",X"20",X"E2",X"00",X"A9",X"D4",X"20",X"DB",X"CF",X"20",X"9D",X"E7",
		X"A5",X"33",X"A4",X"34",X"85",X"22",X"84",X"23",X"60",X"A6",X"A9",X"E8",X"D0",X"86",X"A2",X"95",
		X"2C",X"A2",X"E5",X"4C",X"85",X"C4",X"20",X"54",X"D4",X"20",X"19",X"D4",X"20",X"D6",X"CF",X"A9",
		X"80",X"85",X"2B",X"20",X"FC",X"D0",X"20",X"7A",X"CE",X"20",X"D3",X"CF",X"A9",X"D4",X"20",X"DB",
		X"CF",X"48",X"A5",X"B7",X"48",X"A5",X"B6",X"48",X"A5",X"EA",X"48",X"A5",X"E9",X"48",X"20",X"0A",
		X"CA",X"4C",X"C2",X"D4",X"A9",X"C4",X"20",X"DB",X"CF",X"09",X"80",X"85",X"2B",X"20",X"03",X"D1",
		X"85",X"BD",X"84",X"BE",X"4C",X"7A",X"CE",X"20",X"54",X"D4",X"A5",X"BE",X"48",X"A5",X"BD",X"48",
		X"20",X"CD",X"CF",X"20",X"7A",X"CE",X"68",X"85",X"BD",X"68",X"85",X"BE",X"A0",X"02",X"B1",X"BD",
		X"85",X"B6",X"AA",X"C8",X"B1",X"BD",X"F0",X"99",X"85",X"B7",X"C8",X"B1",X"B6",X"48",X"88",X"10",
		X"FA",X"A4",X"B7",X"20",X"A5",X"DE",X"A5",X"EA",X"48",X"A5",X"E9",X"48",X"B1",X"BD",X"85",X"E9",
		X"C8",X"B1",X"BD",X"85",X"EA",X"A5",X"B7",X"48",X"A5",X"B6",X"48",X"20",X"77",X"CE",X"68",X"85",
		X"BD",X"68",X"85",X"BE",X"20",X"E8",X"00",X"F0",X"03",X"4C",X"E4",X"CF",X"68",X"85",X"E9",X"68",
		X"85",X"EA",X"A0",X"00",X"68",X"91",X"BD",X"68",X"C8",X"91",X"BD",X"68",X"C8",X"91",X"BD",X"68",
		X"C8",X"91",X"BD",X"68",X"C8",X"91",X"BD",X"60",X"20",X"7A",X"CE",X"A0",X"00",X"20",X"D3",X"E0",
		X"68",X"68",X"A9",X"FF",X"A0",X"00",X"F0",X"12",X"A6",X"D3",X"A4",X"D4",X"86",X"BF",X"84",X"C0",
		X"20",X"63",X"D5",X"86",X"D1",X"84",X"D2",X"85",X"D0",X"60",X"A2",X"22",X"86",X"24",X"86",X"25",
		X"85",X"DE",X"84",X"DF",X"85",X"D1",X"84",X"D2",X"A0",X"FF",X"C8",X"B1",X"DE",X"F0",X"0C",X"C5",
		X"24",X"F0",X"04",X"C5",X"25",X"D0",X"F3",X"C9",X"22",X"F0",X"01",X"18",X"84",X"D0",X"98",X"65",
		X"DE",X"85",X"E0",X"A6",X"DF",X"90",X"01",X"E8",X"86",X"E1",X"A5",X"DF",X"D0",X"0B",X"98",X"20",
		X"E8",X"D4",X"A6",X"DE",X"A4",X"DF",X"20",X"F7",X"D6",X"A6",X"85",X"E0",X"91",X"D0",X"05",X"A2",
		X"C4",X"4C",X"85",X"C4",X"A5",X"D0",X"95",X"00",X"A5",X"D1",X"95",X"01",X"A5",X"D2",X"95",X"02",
		X"A0",X"00",X"86",X"D3",X"84",X"D4",X"84",X"DF",X"88",X"84",X"28",X"86",X"86",X"E8",X"E8",X"E8",
		X"86",X"85",X"60",X"46",X"2A",X"48",X"49",X"FF",X"38",X"65",X"A2",X"A4",X"A3",X"B0",X"01",X"88",
		X"C4",X"A1",X"90",X"11",X"D0",X"04",X"C5",X"A0",X"90",X"0B",X"85",X"A2",X"84",X"A3",X"85",X"A4",
		X"84",X"A5",X"AA",X"68",X"60",X"A2",X"4D",X"A5",X"2A",X"30",X"B6",X"20",X"95",X"D5",X"A9",X"80",
		X"85",X"2A",X"68",X"D0",X"D0",X"A6",X"A6",X"A5",X"A7",X"86",X"A2",X"85",X"A3",X"A0",X"00",X"84",
		X"BE",X"84",X"BD",X"A5",X"A0",X"A6",X"A1",X"85",X"CE",X"86",X"CF",X"A9",X"88",X"A2",X"00",X"85",
		X"91",X"86",X"92",X"C5",X"85",X"F0",X"05",X"20",X"36",X"D6",X"F0",X"F7",X"A9",X"07",X"85",X"C2",
		X"A5",X"9C",X"A6",X"9D",X"85",X"91",X"86",X"92",X"E4",X"9F",X"D0",X"04",X"C5",X"9E",X"F0",X"05",
		X"20",X"2C",X"D6",X"F0",X"F3",X"85",X"C7",X"86",X"C8",X"A9",X"03",X"85",X"C2",X"A5",X"C7",X"A6",
		X"C8",X"E4",X"A1",X"D0",X"07",X"C5",X"A0",X"D0",X"03",X"4C",X"75",X"D6",X"85",X"91",X"86",X"92",
		X"A0",X"00",X"B1",X"91",X"AA",X"C8",X"B1",X"91",X"08",X"C8",X"B1",X"91",X"65",X"C7",X"85",X"C7",
		X"C8",X"B1",X"91",X"65",X"C8",X"85",X"C8",X"28",X"10",X"D3",X"8A",X"30",X"D0",X"C8",X"B1",X"91",
		X"A0",X"00",X"0A",X"69",X"05",X"65",X"91",X"85",X"91",X"90",X"02",X"E6",X"92",X"A6",X"92",X"E4",
		X"C8",X"D0",X"04",X"C5",X"C7",X"F0",X"BA",X"20",X"36",X"D6",X"F0",X"F3",X"B1",X"91",X"30",X"35",
		X"C8",X"B1",X"91",X"10",X"30",X"C8",X"B1",X"91",X"F0",X"2B",X"C8",X"B1",X"91",X"AA",X"C8",X"B1",
		X"91",X"C5",X"A3",X"90",X"06",X"D0",X"1E",X"E4",X"A2",X"B0",X"1A",X"C5",X"CF",X"90",X"16",X"D0",
		X"04",X"E4",X"CE",X"90",X"10",X"86",X"CE",X"85",X"CF",X"A5",X"91",X"A6",X"92",X"85",X"BD",X"86",
		X"BE",X"A5",X"C2",X"85",X"C4",X"A5",X"C2",X"18",X"65",X"91",X"85",X"91",X"90",X"02",X"E6",X"92",
		X"A6",X"92",X"A0",X"00",X"60",X"A5",X"BE",X"05",X"BD",X"F0",X"F5",X"A5",X"C4",X"29",X"04",X"4A",
		X"A8",X"85",X"C4",X"B1",X"BD",X"65",X"CE",X"85",X"C9",X"A5",X"CF",X"69",X"00",X"85",X"CA",X"A5",
		X"A2",X"A6",X"A3",X"85",X"C7",X"86",X"C8",X"20",X"FF",X"C3",X"A4",X"C4",X"C8",X"A5",X"C7",X"91",
		X"BD",X"AA",X"E6",X"C8",X"A5",X"C8",X"C8",X"91",X"BD",X"4C",X"99",X"D5",X"A5",X"D4",X"48",X"A5",
		X"D3",X"48",X"20",X"74",X"CF",X"20",X"7C",X"CE",X"68",X"85",X"DE",X"68",X"85",X"DF",X"A0",X"00",
		X"B1",X"DE",X"18",X"71",X"D3",X"90",X"05",X"A2",X"B5",X"4C",X"85",X"C4",X"20",X"E8",X"D4",X"20",
		X"E9",X"D6",X"A5",X"BF",X"A4",X"C0",X"20",X"19",X"D7",X"20",X"FB",X"D6",X"A5",X"DE",X"A4",X"DF",
		X"20",X"19",X"D7",X"20",X"39",X"D5",X"4C",X"A5",X"CE",X"A0",X"00",X"B1",X"DE",X"48",X"C8",X"B1",
		X"DE",X"AA",X"C8",X"B1",X"DE",X"A8",X"68",X"86",X"91",X"84",X"92",X"A8",X"F0",X"0A",X"48",X"88",
		X"B1",X"91",X"91",X"A4",X"98",X"D0",X"F8",X"68",X"18",X"65",X"A4",X"85",X"A4",X"90",X"02",X"E6",
		X"A5",X"60",X"20",X"7C",X"CE",X"A5",X"D3",X"A4",X"D4",X"85",X"91",X"84",X"92",X"20",X"4A",X"D7",
		X"08",X"A0",X"00",X"B1",X"91",X"48",X"C8",X"B1",X"91",X"AA",X"C8",X"B1",X"91",X"A8",X"68",X"28",
		X"D0",X"13",X"C4",X"A3",X"D0",X"0F",X"E4",X"A2",X"D0",X"0B",X"48",X"18",X"65",X"A2",X"85",X"A2",
		X"90",X"02",X"E6",X"A3",X"68",X"86",X"91",X"84",X"92",X"60",X"C4",X"87",X"D0",X"0C",X"C5",X"86",
		X"D0",X"08",X"85",X"85",X"E9",X"03",X"85",X"86",X"A0",X"00",X"60",X"20",X"10",X"D8",X"8A",X"48",
		X"A9",X"01",X"20",X"F0",X"D4",X"68",X"A0",X"00",X"91",X"D1",X"68",X"68",X"4C",X"39",X"D5",X"20",
		X"D0",X"D7",X"D1",X"BF",X"98",X"90",X"04",X"B1",X"BF",X"AA",X"98",X"48",X"8A",X"48",X"20",X"F0",
		X"D4",X"A5",X"BF",X"A4",X"C0",X"20",X"19",X"D7",X"68",X"A8",X"68",X"18",X"65",X"91",X"85",X"91",
		X"90",X"02",X"E6",X"92",X"98",X"20",X"FB",X"D6",X"4C",X"39",X"D5",X"20",X"D0",X"D7",X"18",X"F1",
		X"BF",X"49",X"FF",X"4C",X"75",X"D7",X"A9",X"FF",X"85",X"D4",X"20",X"E8",X"00",X"C9",X"29",X"F0",
		X"06",X"20",X"D9",X"CF",X"20",X"0D",X"D8",X"20",X"D0",X"D7",X"F0",X"4B",X"CA",X"8A",X"48",X"18",
		X"A2",X"00",X"F1",X"BF",X"B0",X"B6",X"49",X"FF",X"C5",X"D4",X"90",X"B1",X"A5",X"D4",X"B0",X"AD",
		X"20",X"D3",X"CF",X"68",X"A8",X"68",X"85",X"C4",X"68",X"68",X"68",X"AA",X"68",X"85",X"BF",X"68",
		X"85",X"C0",X"A5",X"C4",X"48",X"98",X"48",X"A0",X"00",X"8A",X"60",X"20",X"F1",X"D7",X"4C",X"FD",
		X"D3",X"20",X"12",X"D7",X"A2",X"00",X"86",X"28",X"A8",X"60",X"20",X"F1",X"D7",X"F0",X"08",X"A0",
		X"00",X"B1",X"91",X"A8",X"4C",X"FD",X"D3",X"4C",X"A0",X"D2",X"20",X"E2",X"00",X"20",X"77",X"CE",
		X"20",X"10",X"D2",X"A6",X"D3",X"D0",X"F0",X"A6",X"D4",X"4C",X"E8",X"00",X"20",X"F1",X"D7",X"D0",
		X"03",X"4C",X"27",X"DB",X"A6",X"E9",X"A4",X"EA",X"86",X"E0",X"84",X"E1",X"A6",X"91",X"86",X"E9",
		X"18",X"65",X"91",X"85",X"93",X"A6",X"92",X"86",X"EA",X"90",X"01",X"E8",X"86",X"94",X"A0",X"00",
		X"B1",X"93",X"48",X"A9",X"00",X"91",X"93",X"20",X"E8",X"00",X"20",X"CF",X"DF",X"68",X"A0",X"00",
		X"91",X"93",X"A6",X"E0",X"A4",X"E1",X"86",X"E9",X"84",X"EA",X"60",X"20",X"77",X"CE",X"20",X"67",
		X"D8",X"20",X"D9",X"CF",X"4C",X"0D",X"D8",X"A5",X"D5",X"30",X"9C",X"A5",X"D0",X"C9",X"91",X"B0",
		X"96",X"20",X"74",X"DF",X"A5",X"D3",X"A4",X"D4",X"84",X"33",X"85",X"34",X"60",X"A5",X"34",X"48",
		X"A5",X"33",X"48",X"20",X"67",X"D8",X"A0",X"00",X"B1",X"33",X"A8",X"68",X"85",X"33",X"68",X"85",
		X"34",X"4C",X"FD",X"D3",X"20",X"5B",X"D8",X"8A",X"A0",X"00",X"91",X"33",X"60",X"20",X"77",X"CE",
		X"20",X"67",X"D8",X"A4",X"33",X"A6",X"34",X"A9",X"02",X"4C",X"DC",X"EB",X"20",X"9D",X"E7",X"A5",
		X"33",X"A4",X"34",X"85",X"1D",X"84",X"1E",X"20",X"D9",X"CF",X"20",X"9D",X"E7",X"A0",X"01",X"B9",
		X"33",X"00",X"91",X"1D",X"88",X"10",X"F8",X"60",X"20",X"67",X"D8",X"A0",X"01",X"B1",X"33",X"48",
		X"88",X"B1",X"33",X"A8",X"68",X"20",X"ED",X"D3",X"24",X"D5",X"10",X"07",X"A9",X"E4",X"A0",X"D8",
		X"4C",X"97",X"DA",X"60",X"91",X"00",X"00",X"00",X"00",X"82",X"49",X"0F",X"DA",X"9E",X"A9",X"E9",
		X"A0",X"D8",X"4C",X"73",X"DE",X"48",X"4A",X"4A",X"4A",X"4A",X"20",X"FE",X"D8",X"68",X"29",X"0F",
		X"09",X"30",X"C9",X"3A",X"90",X"02",X"69",X"06",X"C9",X"30",X"D0",X"04",X"A4",X"2F",X"F0",X"06",
		X"85",X"2F",X"9D",X"00",X"01",X"E8",X"60",X"20",X"67",X"D8",X"A2",X"00",X"86",X"2F",X"A9",X"23",
		X"85",X"FF",X"A5",X"34",X"20",X"F5",X"D8",X"A5",X"33",X"20",X"F5",X"D8",X"A9",X"00",X"9D",X"00",
		X"01",X"4C",X"E0",X"D4",X"4C",X"E4",X"CF",X"20",X"A9",X"E9",X"20",X"0D",X"D8",X"8A",X"F0",X"06",
		X"CA",X"D0",X"F1",X"A9",X"09",X"2C",X"A9",X"08",X"A2",X"10",X"8E",X"F8",X"02",X"A2",X"1B",X"48",
		X"8A",X"20",X"65",X"D9",X"AD",X"F8",X"02",X"A0",X"27",X"91",X"1F",X"88",X"D0",X"FB",X"68",X"91",
		X"1F",X"CA",X"D0",X"EB",X"60",X"48",X"A9",X"00",X"85",X"20",X"68",X"85",X"1F",X"0A",X"26",X"20",
		X"0A",X"26",X"20",X"18",X"65",X"1F",X"90",X"02",X"E6",X"20",X"0A",X"26",X"20",X"0A",X"26",X"20",
		X"0A",X"26",X"20",X"85",X"1F",X"18",X"69",X"80",X"48",X"85",X"1F",X"A9",X"BB",X"65",X"20",X"85",
		X"20",X"68",X"60",X"4C",X"07",X"D8",X"20",X"6B",X"DA",X"20",X"0D",X"D8",X"E0",X"27",X"B0",X"F3",
		X"E8",X"8E",X"F8",X"02",X"20",X"D9",X"CF",X"20",X"0D",X"D8",X"E0",X"1B",X"B0",X"E5",X"E8",X"8A",
		X"20",X"65",X"D9",X"60",X"20",X"D6",X"CF",X"20",X"96",X"D9",X"20",X"D3",X"CF",X"AC",X"F8",X"02",
		X"B1",X"1F",X"A8",X"4C",X"FD",X"D3",X"20",X"96",X"D9",X"20",X"D9",X"CF",X"20",X"8B",X"CE",X"24",
		X"28",X"10",X"1D",X"20",X"15",X"D7",X"AA",X"18",X"AD",X"F8",X"02",X"65",X"1F",X"90",X"02",X"E6",
		X"20",X"85",X"1F",X"A0",X"00",X"E8",X"CA",X"F0",X"10",X"B1",X"91",X"91",X"1F",X"C8",X"D0",X"F6",
		X"20",X"10",X"D8",X"8A",X"AC",X"F8",X"02",X"91",X"1F",X"60",X"D0",X"17",X"A9",X"03",X"20",X"3B",
		X"C4",X"A5",X"EA",X"48",X"A5",X"E9",X"48",X"A5",X"A9",X"48",X"A5",X"A8",X"48",X"A9",X"8B",X"48",
		X"4C",X"AD",X"C8",X"4C",X"E4",X"CF",X"A9",X"FF",X"85",X"B9",X"20",X"CA",X"C3",X"9A",X"C9",X"8B",
		X"F0",X"05",X"A2",X"F5",X"4C",X"85",X"C4",X"C0",X"10",X"D0",X"05",X"84",X"D0",X"98",X"D0",X"06",
		X"20",X"E8",X"00",X"20",X"8B",X"CE",X"68",X"A5",X"D0",X"F0",X"05",X"68",X"68",X"68",X"68",X"60",
		X"68",X"85",X"A8",X"68",X"85",X"A9",X"68",X"85",X"E9",X"68",X"85",X"EA",X"4C",X"01",X"DA",X"20",
		X"05",X"E9",X"08",X"48",X"10",X"03",X"A9",X"01",X"2C",X"A9",X"00",X"20",X"F0",X"D4",X"68",X"28",
		X"10",X"04",X"A0",X"00",X"91",X"D1",X"68",X"68",X"4C",X"39",X"D5",X"AD",X"C0",X"02",X"29",X"01",
		X"F0",X"05",X"A2",X"A3",X"4C",X"85",X"C4",X"60",X"60",X"A9",X"01",X"A0",X"E2",X"4C",X"97",X"DA",
		X"20",X"4D",X"DD",X"A5",X"D5",X"49",X"FF",X"85",X"D5",X"45",X"DD",X"85",X"DE",X"A5",X"D0",X"4C",
		X"9A",X"DA",X"20",X"FB",X"DB",X"90",X"3C",X"20",X"4D",X"DD",X"D0",X"03",X"4C",X"CD",X"DE",X"A6",
		X"DF",X"86",X"C5",X"A2",X"D8",X"A5",X"D8",X"A8",X"F0",X"CE",X"38",X"E5",X"D0",X"F0",X"24",X"90",
		X"12",X"84",X"D0",X"A4",X"DD",X"84",X"D5",X"49",X"FF",X"69",X"00",X"A0",X"00",X"84",X"C5",X"A2",
		X"D0",X"D0",X"04",X"A0",X"00",X"84",X"DF",X"C9",X"F9",X"30",X"C7",X"A8",X"A5",X"DF",X"56",X"01",
		X"20",X"14",X"DC",X"24",X"DE",X"10",X"57",X"A0",X"D0",X"E0",X"D8",X"F0",X"02",X"A0",X"D8",X"38",
		X"49",X"FF",X"65",X"C5",X"85",X"DF",X"B9",X"04",X"00",X"F5",X"04",X"85",X"D4",X"B9",X"03",X"00",
		X"F5",X"03",X"85",X"D3",X"B9",X"02",X"00",X"F5",X"02",X"85",X"D2",X"B9",X"01",X"00",X"F5",X"01",
		X"85",X"D1",X"B0",X"03",X"20",X"A9",X"DB",X"A0",X"00",X"98",X"18",X"A6",X"D1",X"D0",X"4A",X"A6",
		X"D2",X"86",X"D1",X"A6",X"D3",X"86",X"D2",X"A6",X"D4",X"86",X"D3",X"A6",X"DF",X"86",X"D4",X"84",
		X"DF",X"69",X"08",X"C9",X"28",X"D0",X"E4",X"A9",X"00",X"85",X"D0",X"85",X"D5",X"60",X"65",X"C5",
		X"85",X"DF",X"A5",X"D4",X"65",X"DC",X"85",X"D4",X"A5",X"D3",X"65",X"DB",X"85",X"D3",X"A5",X"D2",
		X"65",X"DA",X"85",X"D2",X"A5",X"D1",X"65",X"D9",X"85",X"D1",X"4C",X"66",X"DB",X"69",X"01",X"06",
		X"DF",X"26",X"D4",X"26",X"D3",X"26",X"D2",X"26",X"D1",X"10",X"F2",X"38",X"E5",X"D0",X"B0",X"C7",
		X"49",X"FF",X"69",X"01",X"85",X"D0",X"90",X"40",X"E6",X"D0",X"F0",X"74",X"A9",X"00",X"90",X"02",
		X"A9",X"80",X"46",X"D1",X"05",X"D1",X"85",X"D1",X"A9",X"00",X"90",X"02",X"A9",X"80",X"46",X"D2",
		X"05",X"D2",X"85",X"D2",X"A9",X"00",X"90",X"02",X"A9",X"80",X"46",X"D3",X"05",X"D3",X"85",X"D3",
		X"A9",X"00",X"90",X"02",X"A9",X"80",X"46",X"D4",X"05",X"D4",X"85",X"D4",X"A9",X"00",X"90",X"02",
		X"A9",X"80",X"46",X"DF",X"05",X"DF",X"85",X"DF",X"60",X"A5",X"D5",X"49",X"FF",X"85",X"D5",X"A5",
		X"D1",X"49",X"FF",X"85",X"D1",X"A5",X"D2",X"49",X"FF",X"85",X"D2",X"A5",X"D3",X"49",X"FF",X"85",
		X"D3",X"A5",X"D4",X"49",X"FF",X"85",X"D4",X"A5",X"DF",X"49",X"FF",X"85",X"DF",X"E6",X"DF",X"D0",
		X"0E",X"E6",X"D4",X"D0",X"0A",X"E6",X"D3",X"D0",X"06",X"E6",X"D2",X"D0",X"02",X"E6",X"D1",X"60",
		X"A2",X"45",X"4C",X"85",X"C4",X"A2",X"94",X"B4",X"04",X"84",X"DF",X"B4",X"03",X"94",X"04",X"B4",
		X"02",X"94",X"03",X"B4",X"01",X"94",X"02",X"A4",X"D7",X"94",X"01",X"69",X"08",X"30",X"E8",X"F0",
		X"E6",X"E9",X"08",X"A8",X"A5",X"DF",X"B0",X"3C",X"48",X"B5",X"01",X"29",X"80",X"56",X"01",X"15",
		X"01",X"95",X"01",X"24",X"48",X"A9",X"00",X"90",X"02",X"A9",X"80",X"56",X"02",X"15",X"02",X"95",
		X"02",X"A9",X"00",X"90",X"02",X"A9",X"80",X"56",X"03",X"15",X"03",X"95",X"03",X"A9",X"00",X"90",
		X"02",X"A9",X"80",X"56",X"04",X"15",X"04",X"95",X"04",X"68",X"08",X"4A",X"28",X"90",X"02",X"09",
		X"80",X"C8",X"D0",X"C4",X"18",X"60",X"82",X"13",X"5D",X"8D",X"DE",X"81",X"00",X"00",X"00",X"00",
		X"03",X"7F",X"5E",X"56",X"CB",X"79",X"80",X"13",X"9B",X"0B",X"64",X"80",X"76",X"38",X"93",X"16",
		X"82",X"38",X"AA",X"3B",X"20",X"80",X"35",X"04",X"F3",X"34",X"81",X"35",X"04",X"F3",X"34",X"80",
		X"80",X"00",X"00",X"00",X"80",X"31",X"72",X"17",X"F8",X"20",X"04",X"DF",X"F0",X"02",X"10",X"03",
		X"4C",X"A0",X"D2",X"A5",X"D0",X"E9",X"7F",X"48",X"A9",X"80",X"85",X"D0",X"A9",X"65",X"A0",X"DC",
		X"20",X"97",X"DA",X"A9",X"6A",X"A0",X"DC",X"20",X"E0",X"DD",X"A9",X"4B",X"A0",X"DC",X"20",X"80",
		X"DA",X"A9",X"50",X"A0",X"DC",X"20",X"F9",X"E2",X"A9",X"6F",X"A0",X"DC",X"20",X"97",X"DA",X"68",
		X"20",X"72",X"E0",X"A9",X"74",X"A0",X"DC",X"20",X"4D",X"DD",X"D0",X"03",X"4C",X"4C",X"DD",X"20",
		X"78",X"DD",X"A9",X"00",X"85",X"95",X"85",X"96",X"85",X"97",X"85",X"98",X"A5",X"DF",X"20",X"E8",
		X"DC",X"A5",X"D4",X"20",X"E8",X"DC",X"A5",X"D3",X"20",X"E8",X"DC",X"A5",X"D2",X"20",X"E8",X"DC",
		X"A5",X"D1",X"20",X"ED",X"DC",X"4C",X"60",X"DE",X"D0",X"03",X"4C",X"E5",X"DB",X"4A",X"09",X"80",
		X"A8",X"90",X"19",X"18",X"A5",X"98",X"65",X"DC",X"85",X"98",X"A5",X"97",X"65",X"DB",X"85",X"97",
		X"A5",X"96",X"65",X"DA",X"85",X"96",X"A5",X"95",X"65",X"D9",X"85",X"95",X"A9",X"00",X"90",X"02",
		X"A9",X"80",X"46",X"95",X"05",X"95",X"85",X"95",X"A9",X"00",X"90",X"02",X"A9",X"80",X"46",X"96",
		X"05",X"96",X"85",X"96",X"A9",X"00",X"90",X"02",X"A9",X"80",X"46",X"97",X"05",X"97",X"85",X"97",
		X"A9",X"00",X"90",X"02",X"A9",X"80",X"46",X"98",X"05",X"98",X"85",X"98",X"A9",X"00",X"90",X"02",
		X"A9",X"80",X"46",X"DF",X"05",X"DF",X"85",X"DF",X"98",X"4A",X"D0",X"A4",X"60",X"85",X"91",X"84",
		X"92",X"A0",X"04",X"B1",X"91",X"85",X"DC",X"88",X"B1",X"91",X"85",X"DB",X"88",X"B1",X"91",X"85",
		X"DA",X"88",X"B1",X"91",X"85",X"DD",X"45",X"D5",X"85",X"DE",X"A5",X"DD",X"09",X"80",X"85",X"D9",
		X"88",X"B1",X"91",X"85",X"D8",X"A5",X"D0",X"60",X"A5",X"D8",X"F0",X"1F",X"18",X"65",X"D0",X"90",
		X"04",X"30",X"1D",X"18",X"2C",X"10",X"14",X"69",X"80",X"85",X"D0",X"D0",X"03",X"4C",X"2B",X"DB",
		X"A5",X"DE",X"85",X"D5",X"60",X"A5",X"D5",X"49",X"FF",X"30",X"05",X"68",X"68",X"4C",X"27",X"DB",
		X"4C",X"E0",X"DB",X"20",X"DD",X"DE",X"AA",X"F0",X"10",X"18",X"69",X"02",X"B0",X"F2",X"A2",X"00",
		X"86",X"DE",X"20",X"A7",X"DA",X"E6",X"D0",X"F0",X"E7",X"60",X"84",X"20",X"00",X"00",X"00",X"20",
		X"DD",X"DE",X"A9",X"BA",X"A0",X"DD",X"A2",X"00",X"86",X"DE",X"20",X"73",X"DE",X"4C",X"E3",X"DD",
		X"20",X"79",X"DC",X"20",X"DD",X"DE",X"A9",X"46",X"A0",X"DC",X"20",X"73",X"DE",X"4C",X"E3",X"DD",
		X"20",X"4D",X"DD",X"F0",X"76",X"20",X"EC",X"DE",X"A9",X"00",X"38",X"E5",X"D0",X"85",X"D0",X"20",
		X"78",X"DD",X"E6",X"D0",X"F0",X"AA",X"A2",X"FC",X"A9",X"01",X"A4",X"D9",X"C4",X"D1",X"D0",X"10",
		X"A4",X"DA",X"C4",X"D2",X"D0",X"0A",X"A4",X"DB",X"C4",X"D3",X"D0",X"04",X"A4",X"DC",X"C4",X"D4",
		X"08",X"2A",X"90",X"09",X"E8",X"95",X"98",X"F0",X"32",X"10",X"34",X"A9",X"01",X"28",X"B0",X"0E",
		X"06",X"DC",X"26",X"DB",X"26",X"DA",X"26",X"D9",X"B0",X"E6",X"30",X"CE",X"10",X"E2",X"A8",X"A5",
		X"DC",X"E5",X"D4",X"85",X"DC",X"A5",X"DB",X"E5",X"D3",X"85",X"DB",X"A5",X"DA",X"E5",X"D2",X"85",
		X"DA",X"A5",X"D9",X"E5",X"D1",X"85",X"D9",X"98",X"4C",X"20",X"DE",X"A9",X"40",X"D0",X"CE",X"0A",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"85",X"DF",X"28",X"4C",X"60",X"DE",X"A2",X"85",X"4C",X"85",X"C4",
		X"A5",X"95",X"85",X"D1",X"A5",X"96",X"85",X"D2",X"A5",X"97",X"85",X"D3",X"A5",X"98",X"85",X"D4",
		X"4C",X"07",X"DB",X"85",X"91",X"84",X"92",X"A0",X"04",X"B1",X"91",X"85",X"D4",X"88",X"B1",X"91",
		X"85",X"D3",X"88",X"B1",X"91",X"85",X"D2",X"88",X"B1",X"91",X"85",X"D5",X"09",X"80",X"85",X"D1",
		X"88",X"B1",X"91",X"85",X"D0",X"84",X"DF",X"60",X"A2",X"CB",X"2C",X"A2",X"C6",X"A0",X"00",X"F0",
		X"04",X"A6",X"B8",X"A4",X"B9",X"20",X"EC",X"DE",X"86",X"91",X"84",X"92",X"A0",X"04",X"A5",X"D4",
		X"91",X"91",X"88",X"A5",X"D3",X"91",X"91",X"88",X"A5",X"D2",X"91",X"91",X"88",X"A5",X"D5",X"09",
		X"7F",X"25",X"D1",X"91",X"91",X"88",X"A5",X"D0",X"91",X"91",X"84",X"DF",X"60",X"A5",X"DD",X"85",
		X"D5",X"A2",X"05",X"B5",X"D7",X"95",X"CF",X"CA",X"D0",X"F9",X"86",X"DF",X"60",X"20",X"EC",X"DE",
		X"A2",X"06",X"B5",X"CF",X"95",X"D7",X"CA",X"D0",X"F9",X"86",X"DF",X"60",X"A5",X"D0",X"F0",X"FB",
		X"06",X"DF",X"90",X"F7",X"20",X"D1",X"DB",X"D0",X"F2",X"4C",X"68",X"DB",X"A9",X"00",X"F0",X"15",
		X"A9",X"FF",X"30",X"11",X"A5",X"D0",X"F0",X"09",X"A5",X"D5",X"2A",X"A9",X"FF",X"B0",X"02",X"A9",
		X"01",X"60",X"20",X"04",X"DF",X"85",X"D1",X"A9",X"00",X"85",X"D2",X"A2",X"88",X"A5",X"D1",X"49",
		X"FF",X"2A",X"A9",X"00",X"85",X"D4",X"85",X"D3",X"86",X"D0",X"85",X"DF",X"85",X"D5",X"4C",X"02",
		X"DB",X"46",X"D5",X"60",X"85",X"93",X"84",X"94",X"A0",X"00",X"B1",X"93",X"C8",X"AA",X"F0",X"C4",
		X"B1",X"93",X"45",X"D5",X"30",X"C2",X"E4",X"D0",X"D0",X"21",X"B1",X"93",X"09",X"80",X"C5",X"D1",
		X"D0",X"19",X"C8",X"B1",X"93",X"C5",X"D2",X"D0",X"12",X"C8",X"B1",X"93",X"C5",X"D3",X"D0",X"0B",
		X"C8",X"A9",X"7F",X"C5",X"DF",X"B1",X"93",X"E5",X"D4",X"F0",X"28",X"A5",X"D5",X"90",X"02",X"49",
		X"FF",X"4C",X"0A",X"DF",X"A5",X"D0",X"F0",X"4A",X"38",X"E9",X"A0",X"24",X"D5",X"10",X"09",X"AA",
		X"A9",X"FF",X"85",X"D7",X"20",X"AF",X"DB",X"8A",X"A2",X"D0",X"C9",X"F9",X"10",X"06",X"20",X"FB",
		X"DB",X"84",X"D7",X"60",X"A8",X"A5",X"D5",X"29",X"80",X"46",X"D1",X"05",X"D1",X"85",X"D1",X"20",
		X"14",X"DC",X"84",X"D7",X"60",X"A5",X"D0",X"C9",X"A0",X"B0",X"20",X"20",X"74",X"DF",X"84",X"DF",
		X"A5",X"D5",X"84",X"D5",X"49",X"80",X"2A",X"A9",X"A0",X"85",X"D0",X"A5",X"D4",X"85",X"24",X"4C",
		X"02",X"DB",X"85",X"D1",X"85",X"D2",X"85",X"D3",X"85",X"D4",X"A8",X"60",X"4C",X"48",X"E8",X"A0",
		X"00",X"A2",X"0A",X"94",X"CC",X"CA",X"10",X"FB",X"90",X"13",X"C9",X"23",X"F0",X"EE",X"C9",X"2D",
		X"D0",X"04",X"86",X"D6",X"F0",X"04",X"C9",X"2B",X"D0",X"05",X"20",X"E2",X"00",X"90",X"6F",X"C9",
		X"2E",X"F0",X"38",X"C9",X"45",X"D0",X"44",X"20",X"E2",X"00",X"90",X"21",X"C9",X"CD",X"F0",X"0E",
		X"C9",X"2D",X"F0",X"0A",X"C9",X"CC",X"F0",X"12",X"C9",X"2B",X"F0",X"0E",X"D0",X"11",X"A9",X"00",
		X"90",X"02",X"A9",X"80",X"46",X"CF",X"05",X"CF",X"85",X"CF",X"20",X"E2",X"00",X"90",X"66",X"24",
		X"CF",X"10",X"18",X"A9",X"00",X"38",X"E5",X"CD",X"4C",X"3D",X"E0",X"A9",X"00",X"90",X"02",X"A9",
		X"80",X"46",X"CE",X"05",X"CE",X"85",X"CE",X"24",X"CE",X"50",X"AF",X"A5",X"CD",X"38",X"E5",X"CC",
		X"85",X"CD",X"F0",X"12",X"10",X"09",X"20",X"BF",X"DD",X"E6",X"CD",X"D0",X"F9",X"F0",X"07",X"20",
		X"A3",X"DD",X"C6",X"CD",X"D0",X"F9",X"A5",X"D6",X"30",X"01",X"60",X"4C",X"6D",X"E2",X"48",X"24",
		X"CE",X"10",X"02",X"E6",X"CC",X"20",X"A3",X"DD",X"68",X"38",X"E9",X"30",X"20",X"72",X"E0",X"4C",
		X"EA",X"DF",X"48",X"20",X"DD",X"DE",X"68",X"20",X"15",X"DF",X"A5",X"DD",X"45",X"D5",X"85",X"DE",
		X"A6",X"D0",X"4C",X"9A",X"DA",X"A5",X"CD",X"C9",X"0A",X"90",X"09",X"A9",X"64",X"24",X"CF",X"30",
		X"11",X"4C",X"E0",X"DB",X"0A",X"0A",X"18",X"65",X"CD",X"0A",X"18",X"A0",X"00",X"71",X"E9",X"38",
		X"E9",X"30",X"85",X"CD",X"4C",X"1A",X"E0",X"9B",X"3E",X"BC",X"1F",X"FD",X"9E",X"6E",X"6B",X"27",
		X"FD",X"9E",X"6E",X"6B",X"28",X"00",X"A9",X"B1",X"A0",X"C3",X"20",X"CE",X"E0",X"A5",X"A9",X"A6",
		X"A8",X"85",X"D1",X"86",X"D2",X"A2",X"90",X"38",X"20",X"22",X"DF",X"20",X"D1",X"E0",X"4C",X"ED",
		X"CB",X"A0",X"01",X"A9",X"02",X"24",X"D5",X"10",X"02",X"A9",X"2D",X"99",X"FF",X"00",X"85",X"D5",
		X"84",X"E0",X"C8",X"A9",X"30",X"A6",X"D0",X"D0",X"03",X"4C",X"F4",X"E1",X"A9",X"00",X"E0",X"80",
		X"F0",X"02",X"B0",X"09",X"A9",X"B1",X"A0",X"E0",X"20",X"B7",X"DC",X"A9",X"F7",X"85",X"CC",X"A9",
		X"AC",X"A0",X"E0",X"20",X"34",X"DF",X"F0",X"1E",X"10",X"12",X"A9",X"A7",X"A0",X"E0",X"20",X"34",
		X"DF",X"F0",X"02",X"10",X"0E",X"20",X"A3",X"DD",X"C6",X"CC",X"D0",X"EE",X"20",X"BF",X"DD",X"E6",
		X"CC",X"D0",X"DC",X"20",X"79",X"DA",X"20",X"74",X"DF",X"A2",X"01",X"A5",X"CC",X"18",X"69",X"0A",
		X"30",X"09",X"C9",X"0B",X"B0",X"06",X"69",X"FF",X"AA",X"A9",X"02",X"38",X"E9",X"02",X"85",X"CD",
		X"86",X"CC",X"8A",X"F0",X"02",X"10",X"13",X"A4",X"E0",X"A9",X"2E",X"C8",X"99",X"FF",X"00",X"8A",
		X"F0",X"06",X"A9",X"30",X"C8",X"99",X"FF",X"00",X"84",X"E0",X"A0",X"00",X"A2",X"80",X"A5",X"D4",
		X"18",X"79",X"09",X"E2",X"85",X"D4",X"A5",X"D3",X"79",X"08",X"E2",X"85",X"D3",X"A5",X"D2",X"79",
		X"07",X"E2",X"85",X"D2",X"A5",X"D1",X"79",X"06",X"E2",X"85",X"D1",X"E8",X"B0",X"04",X"10",X"DE",
		X"30",X"02",X"30",X"DA",X"8A",X"90",X"04",X"49",X"FF",X"69",X"0A",X"69",X"2F",X"C8",X"C8",X"C8",
		X"C8",X"84",X"B6",X"A4",X"E0",X"C8",X"AA",X"29",X"7F",X"99",X"FF",X"00",X"C6",X"CC",X"D0",X"06",
		X"A9",X"2E",X"C8",X"99",X"FF",X"00",X"84",X"E0",X"A4",X"B6",X"8A",X"49",X"FF",X"29",X"80",X"AA",
		X"C0",X"24",X"D0",X"AA",X"A4",X"E0",X"B9",X"FF",X"00",X"88",X"C9",X"30",X"F0",X"F8",X"C9",X"2E",
		X"F0",X"01",X"C8",X"A9",X"2B",X"A6",X"CD",X"F0",X"2E",X"10",X"08",X"A9",X"00",X"38",X"E5",X"CD",
		X"AA",X"A9",X"2D",X"99",X"01",X"01",X"A9",X"45",X"99",X"00",X"01",X"8A",X"A2",X"2F",X"38",X"E8",
		X"E9",X"0A",X"B0",X"FB",X"69",X"3A",X"99",X"03",X"01",X"8A",X"99",X"02",X"01",X"A9",X"00",X"99",
		X"04",X"01",X"F0",X"08",X"99",X"FF",X"00",X"A9",X"00",X"99",X"00",X"01",X"A9",X"00",X"A0",X"01",
		X"60",X"80",X"00",X"00",X"00",X"00",X"FA",X"0A",X"1F",X"00",X"00",X"98",X"96",X"80",X"FF",X"F0",
		X"BD",X"C0",X"00",X"01",X"86",X"A0",X"FF",X"FF",X"D8",X"F0",X"00",X"00",X"03",X"E8",X"FF",X"FF",
		X"FF",X"9C",X"00",X"00",X"00",X"0A",X"FF",X"FF",X"FF",X"FF",X"20",X"DD",X"DE",X"A9",X"01",X"A0",
		X"E2",X"20",X"73",X"DE",X"F0",X"70",X"A5",X"D8",X"D0",X"03",X"4C",X"29",X"DB",X"A2",X"BD",X"A0",
		X"00",X"20",X"A5",X"DE",X"A5",X"DD",X"10",X"0F",X"20",X"A5",X"DF",X"A9",X"BD",X"A0",X"00",X"20",
		X"34",X"DF",X"D0",X"03",X"98",X"A4",X"24",X"20",X"CF",X"DE",X"98",X"48",X"20",X"79",X"DC",X"A9",
		X"BD",X"A0",X"00",X"20",X"B7",X"DC",X"20",X"A6",X"E2",X"68",X"4A",X"90",X"0A",X"A5",X"D0",X"F0",
		X"06",X"A5",X"D5",X"49",X"FF",X"85",X"D5",X"60",X"81",X"38",X"AA",X"3B",X"29",X"07",X"71",X"34",
		X"58",X"3E",X"56",X"74",X"16",X"7E",X"B3",X"1B",X"77",X"2F",X"EE",X"E3",X"85",X"7A",X"1D",X"84",
		X"1C",X"2A",X"7C",X"63",X"59",X"58",X"0A",X"7E",X"75",X"FD",X"E7",X"C6",X"80",X"31",X"72",X"18",
		X"10",X"81",X"00",X"00",X"00",X"00",X"A9",X"78",X"A0",X"E2",X"20",X"B7",X"DC",X"A5",X"DF",X"69",
		X"50",X"90",X"03",X"20",X"F4",X"DE",X"85",X"C5",X"20",X"E0",X"DE",X"A5",X"D0",X"C9",X"88",X"90",
		X"03",X"20",X"95",X"DD",X"20",X"A5",X"DF",X"A5",X"24",X"18",X"69",X"81",X"F0",X"F3",X"38",X"E9",
		X"01",X"48",X"A2",X"05",X"B5",X"D8",X"B4",X"D0",X"95",X"D0",X"94",X"D8",X"CA",X"10",X"F5",X"A5",
		X"C5",X"85",X"DF",X"20",X"83",X"DA",X"20",X"6D",X"E2",X"A9",X"7D",X"A0",X"E2",X"20",X"0F",X"E3",
		X"A9",X"00",X"85",X"DE",X"68",X"20",X"7A",X"DD",X"60",X"85",X"E0",X"84",X"E1",X"20",X"9B",X"DE",
		X"A9",X"C6",X"20",X"B7",X"DC",X"20",X"13",X"E3",X"A9",X"C6",X"A0",X"00",X"4C",X"B7",X"DC",X"85",
		X"E0",X"84",X"E1",X"20",X"98",X"DE",X"B1",X"E0",X"85",X"D6",X"A4",X"E0",X"C8",X"98",X"D0",X"02",
		X"E6",X"E1",X"85",X"E0",X"A4",X"E1",X"20",X"B7",X"DC",X"A5",X"E0",X"A4",X"E1",X"18",X"69",X"05",
		X"90",X"01",X"C8",X"85",X"E0",X"84",X"E1",X"20",X"97",X"DA",X"A9",X"CB",X"A0",X"00",X"C6",X"D6",
		X"D0",X"E4",X"60",X"98",X"35",X"44",X"7A",X"68",X"28",X"B1",X"46",X"20",X"04",X"DF",X"AA",X"30",
		X"18",X"A9",X"FA",X"A0",X"00",X"20",X"73",X"DE",X"8A",X"F0",X"E7",X"A9",X"43",X"A0",X"E3",X"20",
		X"B7",X"DC",X"A9",X"47",X"A0",X"E3",X"20",X"97",X"DA",X"A6",X"D4",X"A5",X"D1",X"85",X"D4",X"86",
		X"D1",X"A9",X"00",X"85",X"D5",X"A5",X"D0",X"85",X"DF",X"A9",X"80",X"85",X"D0",X"20",X"07",X"DB",
		X"A2",X"FA",X"A0",X"00",X"4C",X"A5",X"DE",X"A9",X"03",X"A0",X"E4",X"20",X"97",X"DA",X"20",X"DD",
		X"DE",X"A9",X"08",X"A0",X"E4",X"A6",X"DD",X"20",X"C8",X"DD",X"20",X"DD",X"DE",X"20",X"A5",X"DF",
		X"A9",X"00",X"85",X"DE",X"20",X"83",X"DA",X"A9",X"0D",X"A0",X"E4",X"20",X"80",X"DA",X"A5",X"D5",
		X"48",X"10",X"0D",X"20",X"79",X"DA",X"A5",X"D5",X"30",X"09",X"A5",X"2D",X"49",X"FF",X"85",X"2D",
		X"20",X"6D",X"E2",X"A9",X"0D",X"A0",X"E4",X"20",X"97",X"DA",X"68",X"10",X"03",X"20",X"6D",X"E2",
		X"A9",X"12",X"A0",X"E4",X"4C",X"F9",X"E2",X"20",X"9B",X"DE",X"A9",X"00",X"85",X"2D",X"20",X"8E",
		X"E3",X"A2",X"BD",X"A0",X"00",X"20",X"84",X"E3",X"A9",X"C6",X"A0",X"00",X"20",X"73",X"DE",X"A9",
		X"00",X"85",X"D5",X"A5",X"2D",X"20",X"FF",X"E3",X"A9",X"BD",X"A0",X"00",X"4C",X"E0",X"DD",X"48",
		X"4C",X"C0",X"E3",X"81",X"49",X"0F",X"DA",X"A2",X"83",X"49",X"0F",X"DA",X"A2",X"7F",X"00",X"00",
		X"00",X"00",X"05",X"84",X"E6",X"1A",X"2D",X"1B",X"86",X"28",X"07",X"FB",X"F8",X"87",X"99",X"68",
		X"89",X"01",X"87",X"23",X"35",X"DF",X"E1",X"86",X"A5",X"5D",X"E7",X"28",X"83",X"49",X"0F",X"DA",
		X"A2",X"A1",X"54",X"46",X"8F",X"13",X"8F",X"52",X"43",X"89",X"CD",X"A5",X"D5",X"48",X"10",X"03",
		X"20",X"6D",X"E2",X"A5",X"D0",X"48",X"C9",X"81",X"90",X"07",X"A9",X"4B",X"A0",X"DC",X"20",X"E0",
		X"DD",X"A9",X"6B",X"A0",X"E4",X"20",X"F9",X"E2",X"68",X"C9",X"81",X"90",X"07",X"A9",X"03",X"A0",
		X"E4",X"20",X"80",X"DA",X"68",X"10",X"03",X"4C",X"6D",X"E2",X"60",X"0B",X"76",X"B3",X"83",X"BD",
		X"D3",X"79",X"1E",X"F4",X"A6",X"F5",X"7B",X"83",X"FC",X"B0",X"10",X"7C",X"0C",X"1F",X"67",X"CA",
		X"7C",X"DE",X"53",X"CB",X"C1",X"7D",X"14",X"64",X"70",X"4C",X"7D",X"B7",X"EA",X"51",X"7A",X"7D",
		X"63",X"30",X"88",X"7E",X"7E",X"92",X"44",X"99",X"3A",X"7E",X"4C",X"CC",X"91",X"C7",X"7F",X"AA",
		X"AA",X"AA",X"13",X"81",X"00",X"00",X"00",X"00",X"20",X"63",X"E5",X"A9",X"03",X"A0",X"E5",X"20",
		X"76",X"E5",X"20",X"96",X"E6",X"20",X"30",X"E6",X"C9",X"24",X"D0",X"F9",X"A2",X"09",X"20",X"30",
		X"E6",X"95",X"5D",X"CA",X"D0",X"F8",X"20",X"30",X"E6",X"F0",X"05",X"95",X"49",X"E8",X"D0",X"F6",
		X"95",X"49",X"20",X"F0",X"E6",X"8A",X"D0",X"D0",X"20",X"63",X"E5",X"A9",X"12",X"A0",X"E5",X"20",
		X"76",X"E5",X"20",X"6E",X"E5",X"EA",X"EA",X"E5",X"EA",X"EA",X"EA",X"A5",X"5F",X"A4",X"60",X"85",
		X"33",X"84",X"34",X"A0",X"00",X"20",X"30",X"E6",X"EA",X"B0",X"43",X"91",X"33",X"20",X"54",X"E5",
		X"90",X"F3",X"60",X"10",X"07",X"53",X"65",X"61",X"72",X"63",X"68",X"69",X"6E",X"67",X"20",X"2E",
		X"2E",X"00",X"10",X"07",X"4C",X"6F",X"61",X"64",X"69",X"6E",X"67",X"20",X"20",X"20",X"2E",X"2E",
		X"00",X"0A",X"0D",X"46",X"49",X"4C",X"45",X"20",X"45",X"52",X"52",X"4F",X"52",X"20",X"2F",X"20",
		X"4C",X"4F",X"41",X"44",X"20",X"41",X"42",X"4F",X"52",X"54",X"45",X"44",X"0D",X"00",X"20",X"63",
		X"E5",X"20",X"19",X"C7",X"20",X"04",X"E8",X"20",X"9F",X"CB",X"A9",X"21",X"A0",X"E5",X"20",X"ED",
		X"CB",X"4C",X"B5",X"C4",X"A5",X"33",X"C5",X"61",X"A5",X"34",X"E5",X"62",X"E6",X"33",X"D0",X"02",
		X"E6",X"34",X"60",X"A2",X"1C",X"A9",X"10",X"9D",X"80",X"BB",X"CA",X"10",X"FA",X"60",X"E8",X"E8",
		X"E8",X"A9",X"35",X"A0",X"00",X"2C",X"A2",X"00",X"4C",X"36",X"F4",X"20",X"BA",X"E6",X"A9",X"24",
		X"20",X"C6",X"E5",X"A2",X"09",X"B5",X"5D",X"20",X"C6",X"E5",X"CA",X"D0",X"F8",X"B5",X"35",X"F0",
		X"06",X"20",X"C6",X"E5",X"E8",X"D0",X"F6",X"20",X"C6",X"E5",X"20",X"63",X"E5",X"A9",X"BC",X"A0",
		X"E5",X"20",X"76",X"E5",X"20",X"6E",X"E5",X"A5",X"5F",X"A4",X"60",X"85",X"33",X"84",X"34",X"A0",
		X"00",X"B1",X"33",X"20",X"C6",X"E5",X"20",X"54",X"E5",X"90",X"F6",X"60",X"10",X"07",X"53",X"61",
		X"76",X"69",X"6E",X"67",X"20",X"00",X"85",X"2F",X"8A",X"48",X"98",X"48",X"20",X"27",X"E6",X"18",
		X"A0",X"09",X"A9",X"00",X"F0",X"06",X"46",X"2F",X"08",X"69",X"00",X"28",X"20",X"F3",X"E5",X"88",
		X"D0",X"F4",X"49",X"01",X"4A",X"A0",X"04",X"20",X"F3",X"E5",X"38",X"88",X"D0",X"F9",X"68",X"A8",
		X"68",X"AA",X"60",X"48",X"08",X"A5",X"67",X"D0",X"0A",X"38",X"20",X"19",X"E6",X"28",X"20",X"19",
		X"E6",X"68",X"60",X"20",X"19",X"E6",X"A2",X"0F",X"28",X"B0",X"02",X"A2",X"07",X"20",X"12",X"E6",
		X"68",X"60",X"20",X"27",X"E6",X"CA",X"D0",X"FA",X"60",X"A9",X"D0",X"A2",X"00",X"B0",X"02",X"0A",
		X"E8",X"8D",X"06",X"03",X"8E",X"07",X"03",X"AD",X"04",X"03",X"2C",X"0D",X"03",X"50",X"FB",X"60",
		X"98",X"48",X"8A",X"48",X"20",X"7D",X"E6",X"20",X"7D",X"E6",X"B0",X"FB",X"20",X"61",X"E6",X"B0",
		X"16",X"A9",X"00",X"A0",X"08",X"20",X"5E",X"E6",X"08",X"66",X"2F",X"28",X"69",X"00",X"88",X"D0",
		X"F4",X"20",X"5E",X"E6",X"69",X"00",X"18",X"68",X"AA",X"68",X"A8",X"A5",X"2F",X"60",X"20",X"7D",
		X"E6",X"A5",X"67",X"F0",X"17",X"48",X"20",X"7D",X"E6",X"A2",X"02",X"90",X"02",X"A2",X"06",X"A9",
		X"00",X"20",X"7D",X"E6",X"69",X"00",X"CA",X"D0",X"F8",X"C9",X"04",X"68",X"60",X"48",X"AD",X"00",
		X"03",X"AD",X"0D",X"03",X"29",X"10",X"F0",X"F9",X"AD",X"09",X"03",X"48",X"A9",X"FF",X"8D",X"09",
		X"03",X"68",X"C9",X"FE",X"68",X"60",X"20",X"5E",X"E6",X"66",X"2F",X"A9",X"16",X"C5",X"2F",X"D0",
		X"F5",X"A5",X"67",X"F0",X"08",X"20",X"7D",X"E6",X"20",X"7D",X"E6",X"B0",X"FB",X"A2",X"03",X"20",
		X"30",X"E6",X"C9",X"16",X"D0",X"E0",X"CA",X"D0",X"F6",X"60",X"A2",X"02",X"A0",X"03",X"A9",X"16",
		X"20",X"C6",X"E5",X"88",X"D0",X"F8",X"CA",X"D0",X"F5",X"60",X"20",X"FD",X"EB",X"A0",X"06",X"78",
		X"BE",X"E2",X"E6",X"B9",X"E9",X"E6",X"9D",X"00",X"03",X"88",X"10",X"F4",X"A9",X"40",X"8D",X"00",
		X"03",X"60",X"05",X"04",X"0B",X"02",X"0C",X"08",X"0E",X"00",X"D0",X"C0",X"FF",X"10",X"F4",X"7F",
		X"A0",X"00",X"A2",X"00",X"A5",X"35",X"F0",X"15",X"B9",X"35",X"00",X"D9",X"49",X"00",X"F0",X"01",
		X"E8",X"99",X"49",X"00",X"C8",X"C0",X"11",X"B0",X"04",X"48",X"68",X"D0",X"EB",X"60",X"20",X"63",
		X"E5",X"A9",X"8D",X"A0",X"EB",X"A2",X"00",X"20",X"76",X"E5",X"20",X"05",X"E9",X"10",X"FB",X"4C",
		X"63",X"E5",X"4C",X"E4",X"CF",X"A9",X"00",X"85",X"67",X"85",X"63",X"85",X"64",X"20",X"8B",X"CE",
		X"24",X"28",X"10",X"EE",X"20",X"15",X"D7",X"AA",X"A0",X"00",X"E8",X"CA",X"F0",X"08",X"B1",X"91",
		X"99",X"35",X"00",X"C8",X"D0",X"F5",X"A9",X"00",X"99",X"35",X"00",X"20",X"E8",X"00",X"F0",X"4C",
		X"C9",X"2C",X"D0",X"CE",X"20",X"E2",X"00",X"F0",X"43",X"C9",X"2C",X"F0",X"F7",X"A0",X"05",X"88",
		X"F0",X"C0",X"D9",X"A5",X"E7",X"D0",X"F8",X"C0",X"04",X"90",X"04",X"84",X"63",X"B0",X"E5",X"C0",
		X"03",X"90",X"04",X"84",X"67",X"B0",X"DD",X"20",X"E2",X"00",X"A2",X"80",X"86",X"64",X"C0",X"02",
		X"90",X"0D",X"20",X"9D",X"E7",X"A5",X"33",X"A4",X"34",X"85",X"5F",X"84",X"60",X"90",X"BC",X"20",
		X"9D",X"E7",X"A5",X"33",X"A4",X"34",X"85",X"61",X"84",X"62",X"90",X"AF",X"60",X"20",X"77",X"CE",
		X"20",X"67",X"D8",X"18",X"60",X"21",X"45",X"41",X"53",X"C7",X"A5",X"9A",X"A4",X"9B",X"85",X"5F",
		X"84",X"60",X"08",X"20",X"25",X"E7",X"20",X"CA",X"E6",X"20",X"A8",X"E4",X"20",X"04",X"E8",X"28",
		X"A6",X"61",X"A5",X"62",X"85",X"9D",X"86",X"9C",X"A5",X"63",X"F0",X"0A",X"A5",X"64",X"F0",X"03",
		X"6C",X"5F",X"00",X"4C",X"8B",X"C9",X"68",X"68",X"4C",X"6B",X"C9",X"A5",X"9A",X"A4",X"9B",X"85",
		X"5F",X"84",X"60",X"A5",X"9C",X"A4",X"9D",X"85",X"61",X"84",X"62",X"08",X"20",X"25",X"E7",X"20",
		X"CA",X"E6",X"20",X"7B",X"E5",X"20",X"04",X"E8",X"28",X"A6",X"A9",X"E8",X"F0",X"01",X"60",X"68",
		X"68",X"4C",X"6B",X"C9",X"20",X"63",X"E5",X"20",X"39",X"F4",X"4C",X"D0",X"EB",X"20",X"9D",X"E7",
		X"6C",X"33",X"00",X"A2",X"00",X"86",X"33",X"86",X"34",X"F0",X"13",X"A2",X"03",X"0A",X"0A",X"0A",
		X"0A",X"0A",X"26",X"33",X"26",X"34",X"90",X"03",X"4C",X"E0",X"DB",X"CA",X"10",X"F3",X"20",X"E2",
		X"00",X"C9",X"80",X"B0",X"0E",X"09",X"80",X"49",X"B0",X"C9",X"0A",X"90",X"DE",X"69",X"88",X"C9",
		X"FA",X"B0",X"D8",X"A5",X"34",X"A4",X"33",X"60",X"20",X"13",X"E8",X"4C",X"D5",X"D8",X"1D",X"F4",
		X"23",X"F4",X"20",X"F4",X"DE",X"EB",X"E1",X"EB",X"E4",X"EB",X"E7",X"EB",X"EA",X"EB",X"F9",X"EB",
		X"ED",X"EB",X"F3",X"EB",X"F6",X"EB",X"03",X"04",X"04",X"03",X"03",X"03",X"02",X"01",X"03",X"03",
		X"01",X"01",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"AD",X"C0",X"02",
		X"29",X"01",X"D0",X"05",X"A2",X"A3",X"4C",X"85",X"C4",X"C0",X"4E",X"B0",X"03",X"4C",X"E4",X"CF",
		X"C0",X"66",X"B0",X"F9",X"98",X"38",X"E9",X"4E",X"A8",X"B9",X"4F",X"E8",X"48",X"B9",X"4E",X"E8",
		X"48",X"98",X"4A",X"A8",X"B9",X"66",X"E8",X"48",X"B9",X"72",X"E8",X"8D",X"C3",X"02",X"A9",X"00",
		X"8D",X"F0",X"02",X"20",X"77",X"CE",X"AD",X"C3",X"02",X"D0",X"06",X"20",X"67",X"D8",X"4C",X"C8",
		X"E8",X"A5",X"D0",X"C9",X"90",X"20",X"6F",X"D8",X"AC",X"F0",X"02",X"A5",X"33",X"99",X"E1",X"02",
		X"A5",X"34",X"99",X"E2",X"02",X"C8",X"C8",X"8C",X"F0",X"02",X"68",X"A8",X"88",X"F0",X"08",X"98",
		X"48",X"20",X"D9",X"CF",X"4C",X"B3",X"E8",X"A9",X"00",X"8D",X"E0",X"02",X"68",X"AA",X"68",X"A8",
		X"A9",X"E8",X"48",X"A9",X"FA",X"48",X"98",X"48",X"8A",X"48",X"60",X"A9",X"01",X"2C",X"E0",X"02",
		X"F0",X"F8",X"4C",X"A0",X"D2",X"AD",X"DF",X"02",X"10",X"0B",X"08",X"29",X"7F",X"48",X"A9",X"00",
		X"8D",X"DF",X"02",X"68",X"28",X"60",X"C4",X"9D",X"B0",X"02",X"38",X"60",X"D0",X"06",X"C5",X"9C",
		X"90",X"F9",X"F0",X"F7",X"20",X"42",X"E9",X"90",X"F2",X"AA",X"AD",X"C0",X"02",X"29",X"02",X"08",
		X"8A",X"28",X"D0",X"E6",X"98",X"48",X"38",X"E9",X"1C",X"A8",X"8A",X"20",X"42",X"E9",X"68",X"A8",
		X"8A",X"60",X"CC",X"C2",X"02",X"90",X"02",X"F0",X"01",X"60",X"CD",X"C1",X"02",X"60",X"AC",X"C2",
		X"02",X"AD",X"C1",X"02",X"D0",X"01",X"88",X"38",X"E9",X"01",X"60",X"20",X"77",X"CE",X"20",X"67",
		X"D8",X"A5",X"33",X"A4",X"34",X"20",X"16",X"E9",X"90",X"03",X"4C",X"83",X"C4",X"85",X"A6",X"84",
		X"A7",X"4C",X"3A",X"C7",X"AD",X"C0",X"02",X"48",X"29",X"01",X"F0",X"05",X"A2",X"A3",X"4C",X"85",
		X"C4",X"68",X"29",X"FD",X"8D",X"C0",X"02",X"20",X"4E",X"E9",X"48",X"98",X"18",X"69",X"1C",X"A8",
		X"68",X"4C",X"6D",X"E9",X"20",X"4E",X"E9",X"20",X"16",X"E9",X"B0",X"CE",X"48",X"AD",X"C0",X"02",
		X"09",X"02",X"8D",X"C0",X"02",X"68",X"4C",X"6D",X"E9",X"AD",X"C0",X"02",X"A8",X"29",X"01",X"F0",
		X"09",X"98",X"29",X"FE",X"8D",X"C0",X"02",X"20",X"27",X"F4",X"60",X"AD",X"C0",X"02",X"48",X"29",
		X"02",X"F0",X"B9",X"68",X"09",X"01",X"8D",X"C0",X"02",X"20",X"2A",X"F4",X"60",X"20",X"D6",X"CF",
		X"20",X"8B",X"CE",X"A5",X"34",X"48",X"A5",X"33",X"48",X"20",X"67",X"D8",X"A5",X"33",X"8D",X"E1",
		X"02",X"A5",X"34",X"8D",X"E2",X"02",X"68",X"85",X"33",X"68",X"85",X"34",X"20",X"D9",X"CF",X"20",
		X"8B",X"CE",X"A5",X"34",X"48",X"A5",X"33",X"48",X"20",X"67",X"D8",X"A5",X"34",X"8D",X"E4",X"02",
		X"A5",X"33",X"8D",X"E3",X"02",X"68",X"85",X"33",X"68",X"85",X"34",X"20",X"F1",X"EB",X"AC",X"E1",
		X"02",X"AD",X"E0",X"02",X"29",X"01",X"D0",X"09",X"AD",X"E2",X"02",X"20",X"ED",X"D3",X"4C",X"D3",
		X"CF",X"4C",X"07",X"D8",X"E6",X"E9",X"D0",X"02",X"E6",X"EA",X"AD",X"60",X"EA",X"C9",X"20",X"F0",
		X"F3",X"20",X"41",X"EA",X"60",X"2C",X"60",X"EA",X"2C",X"60",X"EA",X"60",X"80",X"4F",X"C7",X"52",
		X"58",X"C9",X"C8",X"D0",X"05",X"20",X"61",X"CA",X"D0",X"E0",X"C9",X"27",X"F0",X"F7",X"C9",X"3A",
		X"B0",X"06",X"38",X"E9",X"30",X"38",X"E9",X"D0",X"60",X"D8",X"A2",X"FF",X"86",X"A9",X"9A",X"A9",
		X"59",X"A0",X"EA",X"85",X"1B",X"84",X"1C",X"A9",X"4C",X"85",X"1A",X"85",X"C3",X"85",X"21",X"8D",
		X"FB",X"02",X"A9",X"A0",X"A0",X"D2",X"85",X"22",X"84",X"23",X"8D",X"FC",X"02",X"8C",X"FD",X"02",
		X"8D",X"F5",X"02",X"8C",X"F6",X"02",X"A9",X"50",X"85",X"31",X"A9",X"38",X"85",X"32",X"A2",X"1C",
		X"BD",X"23",X"EA",X"95",X"E1",X"CA",X"D0",X"F8",X"A9",X"03",X"85",X"C2",X"8A",X"85",X"D7",X"85",
		X"87",X"85",X"2F",X"48",X"85",X"2E",X"8D",X"F1",X"02",X"8D",X"F2",X"02",X"20",X"83",X"CC",X"20",
		X"9F",X"CB",X"A2",X"88",X"86",X"85",X"A8",X"AD",X"E1",X"02",X"AC",X"E2",X"02",X"85",X"A6",X"84",
		X"A7",X"A9",X"02",X"8D",X"C0",X"02",X"A9",X"50",X"85",X"31",X"E9",X"0E",X"B0",X"FC",X"49",X"FF",
		X"E9",X"0C",X"18",X"65",X"31",X"85",X"32",X"4E",X"F1",X"02",X"20",X"83",X"CC",X"20",X"0A",X"CC",
		X"A9",X"51",X"A0",X"EB",X"20",X"ED",X"CB",X"20",X"9F",X"CB",X"A2",X"00",X"A0",X"05",X"86",X"9A",
		X"84",X"9B",X"A0",X"00",X"98",X"91",X"9A",X"E6",X"9A",X"D0",X"02",X"E6",X"9B",X"20",X"1B",X"C7",
		X"A5",X"9A",X"A4",X"9B",X"20",X"48",X"C4",X"20",X"9F",X"CB",X"A5",X"A6",X"38",X"E5",X"9A",X"AA",
		X"A5",X"A7",X"E5",X"9B",X"20",X"C1",X"E0",X"A9",X"43",X"A0",X"EB",X"20",X"ED",X"CB",X"38",X"A5",
		X"A6",X"E9",X"FF",X"85",X"A6",X"8D",X"C1",X"02",X"A5",X"A7",X"E9",X"20",X"85",X"A7",X"8D",X"C2",
		X"02",X"A9",X"ED",X"A0",X"CB",X"85",X"1B",X"84",X"1C",X"A9",X"10",X"8D",X"F8",X"02",X"4C",X"B5",
		X"C4",X"00",X"00",X"20",X"42",X"59",X"54",X"45",X"53",X"20",X"46",X"52",X"45",X"45",X"0A",X"0D",
		X"00",X"4F",X"52",X"49",X"43",X"20",X"45",X"58",X"54",X"45",X"4E",X"44",X"45",X"44",X"20",X"42",
		X"41",X"53",X"49",X"43",X"20",X"56",X"31",X"2E",X"30",X"0D",X"0A",X"60",X"20",X"31",X"39",X"38",
		X"33",X"20",X"54",X"41",X"4E",X"47",X"45",X"52",X"49",X"4E",X"45",X"0D",X"0A",X"00",X"0D",X"0A",
		X"54",X"4F",X"4F",X"20",X"4C",X"41",X"52",X"47",X"45",X"0D",X"0A",X"00",X"00",X"53",X"6F",X"66",
		X"74",X"77",X"61",X"72",X"65",X"20",X"62",X"79",X"20",X"50",X"45",X"54",X"45",X"52",X"20",X"48",
		X"41",X"4C",X"46",X"4F",X"52",X"44",X"20",X"41",X"4E",X"44",X"20",X"41",X"4E",X"44",X"59",X"20",
		X"42",X"52",X"4F",X"57",X"4E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"4C",X"C7",X"EC",X"4C",X"8F",X"ED",X"4C",X"81",X"ED",X"4C",X"0C",X"EC",X"4C",X"AD",X"ED",X"4C",
		X"2D",X"F0",X"4C",X"64",X"F0",X"4C",X"79",X"F0",X"4C",X"E5",X"F2",X"4C",X"93",X"F0",X"4C",X"A5",
		X"F0",X"4C",X"41",X"F1",X"4C",X"7F",X"F1",X"4C",X"8B",X"F1",X"4C",X"E5",X"F1",X"4C",X"01",X"ED",
		X"4C",X"BC",X"ED",X"4C",X"09",X"ED",X"4C",X"64",X"F2",X"4C",X"50",X"F2",X"48",X"8A",X"48",X"98",
		X"48",X"A2",X"00",X"A0",X"02",X"20",X"80",X"EC",X"F0",X"60",X"08",X"A0",X"00",X"B0",X"21",X"A0",
		X"04",X"A9",X"00",X"8D",X"06",X"02",X"A9",X"FF",X"8D",X"07",X"02",X"A2",X"06",X"A0",X"04",X"20",
		X"95",X"EC",X"A0",X"06",X"A2",X"00",X"20",X"95",X"EC",X"A2",X"02",X"20",X"95",X"EC",X"A0",X"FF",
		X"AD",X"00",X"02",X"85",X"0C",X"AD",X"01",X"02",X"85",X"0D",X"AD",X"02",X"02",X"85",X"0E",X"AD",
		X"03",X"02",X"85",X"0F",X"A2",X"04",X"20",X"AF",X"EC",X"90",X"1E",X"B1",X"0C",X"91",X"0E",X"28",
		X"08",X"B0",X"0C",X"88",X"C0",X"FF",X"D0",X"EE",X"C6",X"0D",X"C6",X"0F",X"4C",X"56",X"EC",X"C8",
		X"D0",X"E4",X"E6",X"0D",X"E6",X"0F",X"4C",X"56",X"EC",X"28",X"68",X"A8",X"68",X"AA",X"68",X"60",
		X"D8",X"38",X"BD",X"00",X"02",X"F9",X"00",X"02",X"8D",X"06",X"02",X"BD",X"01",X"02",X"F9",X"01",
		X"02",X"0D",X"06",X"02",X"60",X"D8",X"18",X"BD",X"00",X"02",X"79",X"00",X"02",X"9D",X"00",X"02",
		X"48",X"BD",X"01",X"02",X"79",X"01",X"02",X"9D",X"01",X"02",X"68",X"1D",X"00",X"02",X"60",X"D8",
		X"38",X"BD",X"00",X"02",X"E9",X"01",X"9D",X"00",X"02",X"48",X"BD",X"01",X"02",X"E9",X"00",X"9D",
		X"01",X"02",X"68",X"1D",X"00",X"02",X"60",X"48",X"20",X"70",X"ED",X"A9",X"00",X"A2",X"00",X"A0",
		X"03",X"20",X"8F",X"ED",X"A9",X"01",X"A0",X"19",X"20",X"8F",X"ED",X"A9",X"00",X"8D",X"71",X"02",
		X"AD",X"0B",X"03",X"29",X"7F",X"09",X"40",X"8D",X"0B",X"03",X"A9",X"C0",X"8D",X"0E",X"03",X"A9",
		X"10",X"8D",X"06",X"03",X"8D",X"04",X"03",X"A9",X"27",X"8D",X"07",X"03",X"8D",X"05",X"03",X"68",
		X"60",X"48",X"A9",X"40",X"8D",X"0E",X"03",X"68",X"60",X"48",X"AD",X"0D",X"03",X"29",X"40",X"F0",
		X"06",X"8D",X"0D",X"03",X"20",X"1B",X"ED",X"68",X"4C",X"30",X"02",X"48",X"8A",X"48",X"98",X"48",
		X"A0",X"00",X"B9",X"72",X"02",X"38",X"E9",X"01",X"99",X"72",X"02",X"C8",X"B9",X"72",X"02",X"E9",
		X"00",X"99",X"72",X"02",X"C8",X"C0",X"06",X"D0",X"E9",X"A9",X"00",X"20",X"81",X"ED",X"C0",X"00",
		X"D0",X"0D",X"A2",X"00",X"A0",X"03",X"20",X"8F",X"ED",X"4C",X"5E",X"FC",X"8E",X"DF",X"02",X"A9",
		X"01",X"20",X"81",X"ED",X"C0",X"00",X"D0",X"12",X"A2",X"00",X"A0",X"19",X"20",X"8F",X"ED",X"AD",
		X"71",X"02",X"49",X"01",X"8D",X"71",X"02",X"20",X"03",X"F4",X"68",X"A8",X"68",X"AA",X"68",X"60",
		X"48",X"98",X"48",X"A0",X"05",X"A9",X"00",X"99",X"72",X"02",X"88",X"10",X"FA",X"68",X"A8",X"68",
		X"60",X"48",X"0A",X"A8",X"78",X"B9",X"72",X"02",X"BE",X"73",X"02",X"58",X"A8",X"68",X"60",X"48",
		X"8A",X"48",X"98",X"48",X"BA",X"BD",X"03",X"01",X"0A",X"A8",X"68",X"48",X"78",X"99",X"72",X"02",
		X"BD",X"02",X"01",X"99",X"73",X"02",X"58",X"68",X"A8",X"68",X"AA",X"68",X"60",X"20",X"8F",X"ED",
		X"20",X"81",X"ED",X"C0",X"00",X"D0",X"F9",X"E0",X"00",X"D0",X"F5",X"60",X"48",X"8A",X"48",X"98",
		X"48",X"A9",X"00",X"85",X"0C",X"A9",X"BF",X"85",X"0D",X"A2",X"1F",X"A9",X"40",X"A0",X"3F",X"91",
		X"0C",X"88",X"C0",X"FF",X"D0",X"F9",X"C6",X"0D",X"CA",X"E0",X"FF",X"D0",X"F2",X"68",X"A8",X"68",
		X"AA",X"68",X"60",X"0E",X"12",X"02",X"0E",X"12",X"02",X"0E",X"12",X"02",X"0E",X"12",X"02",X"0E",
		X"12",X"02",X"0E",X"12",X"02",X"60",X"48",X"98",X"48",X"20",X"E3",X"ED",X"20",X"A6",X"EF",X"20",
		X"5B",X"EF",X"68",X"A8",X"68",X"60",X"48",X"8A",X"48",X"98",X"48",X"AD",X"13",X"02",X"8D",X"14",
		X"02",X"20",X"E3",X"ED",X"2C",X"03",X"02",X"10",X"0B",X"A9",X"FF",X"4D",X"02",X"02",X"8D",X"02",
		X"02",X"EE",X"02",X"02",X"2C",X"05",X"02",X"10",X"0B",X"A9",X"FF",X"4D",X"04",X"02",X"8D",X"04",
		X"02",X"EE",X"04",X"02",X"AD",X"02",X"02",X"CD",X"04",X"02",X"90",X"2A",X"A9",X"00",X"85",X"0C",
		X"8D",X"01",X"02",X"AD",X"04",X"02",X"85",X"0D",X"AD",X"02",X"02",X"8D",X"00",X"02",X"20",X"FF",
		X"EE",X"20",X"31",X"EF",X"A9",X"00",X"85",X"0E",X"85",X"0F",X"8D",X"00",X"02",X"AE",X"02",X"02",
		X"20",X"BB",X"EE",X"4C",X"8D",X"EE",X"A9",X"00",X"85",X"0C",X"8D",X"01",X"02",X"AD",X"02",X"02",
		X"85",X"0D",X"AD",X"04",X"02",X"8D",X"00",X"02",X"20",X"FF",X"EE",X"20",X"31",X"EF",X"A9",X"00",
		X"85",X"0E",X"85",X"0F",X"8D",X"00",X"02",X"AE",X"04",X"02",X"20",X"93",X"EE",X"68",X"A8",X"68",
		X"AA",X"68",X"60",X"2C",X"05",X"02",X"10",X"06",X"20",X"F5",X"EF",X"4C",X"A1",X"EE",X"20",X"E6",
		X"EF",X"20",X"E3",X"EE",X"F0",X"0E",X"2C",X"03",X"02",X"10",X"06",X"20",X"15",X"F0",X"4C",X"B4",
		X"EE",X"20",X"04",X"F0",X"20",X"4D",X"EF",X"CA",X"D0",X"D9",X"60",X"2C",X"03",X"02",X"10",X"06",
		X"20",X"15",X"F0",X"4C",X"C9",X"EE",X"20",X"04",X"F0",X"20",X"E3",X"EE",X"F0",X"0E",X"2C",X"05",
		X"02",X"10",X"06",X"20",X"F5",X"EF",X"4C",X"DC",X"EE",X"20",X"E6",X"EF",X"20",X"4D",X"EF",X"CA",
		X"D0",X"D9",X"60",X"D8",X"18",X"A5",X"0E",X"65",X"0C",X"85",X"0E",X"A5",X"0F",X"65",X"0D",X"85",
		X"0F",X"24",X"0E",X"10",X"03",X"18",X"69",X"01",X"CD",X"00",X"02",X"8D",X"00",X"02",X"60",X"48",
		X"8A",X"48",X"98",X"48",X"A9",X"00",X"85",X"0E",X"85",X"0F",X"A2",X"10",X"06",X"0C",X"26",X"0D",
		X"26",X"0E",X"26",X"0F",X"A5",X"0E",X"38",X"ED",X"00",X"02",X"A8",X"A5",X"0F",X"ED",X"01",X"02",
		X"90",X"06",X"E6",X"0C",X"84",X"0E",X"85",X"0F",X"CA",X"D0",X"E1",X"68",X"A8",X"68",X"AA",X"68",
		X"60",X"48",X"0E",X"00",X"02",X"2E",X"01",X"02",X"AD",X"00",X"02",X"38",X"E5",X"0E",X"AD",X"01",
		X"02",X"E5",X"0F",X"B0",X"06",X"E6",X"0C",X"D0",X"02",X"E6",X"0D",X"68",X"60",X"2C",X"14",X"02",
		X"18",X"10",X"04",X"20",X"5B",X"EF",X"38",X"2E",X"14",X"02",X"60",X"2C",X"12",X"02",X"30",X"0E",
		X"70",X"06",X"20",X"94",X"EF",X"4C",X"73",X"EF",X"20",X"84",X"EF",X"4C",X"73",X"EF",X"70",X"03",
		X"20",X"74",X"EF",X"60",X"A0",X"00",X"B1",X"10",X"29",X"40",X"F0",X"07",X"B1",X"10",X"4D",X"15",
		X"02",X"91",X"10",X"60",X"A0",X"00",X"B1",X"10",X"29",X"40",X"F0",X"07",X"AD",X"15",X"02",X"11",
		X"10",X"91",X"10",X"60",X"A0",X"00",X"B1",X"10",X"29",X"40",X"F0",X"09",X"AD",X"15",X"02",X"49",
		X"FF",X"31",X"10",X"91",X"10",X"60",X"D8",X"48",X"98",X"48",X"20",X"00",X"F4",X"18",X"69",X"00",
		X"85",X"10",X"98",X"69",X"A0",X"85",X"11",X"A9",X"00",X"85",X"0D",X"8D",X"01",X"02",X"86",X"0C",
		X"A9",X"06",X"8D",X"00",X"02",X"20",X"FF",X"EE",X"18",X"A5",X"0C",X"65",X"10",X"85",X"10",X"A9",
		X"00",X"65",X"11",X"85",X"11",X"A9",X"20",X"A4",X"0E",X"F0",X"04",X"4A",X"88",X"90",X"FA",X"8D",
		X"15",X"02",X"68",X"A8",X"68",X"60",X"D8",X"18",X"A5",X"10",X"69",X"28",X"85",X"10",X"A5",X"11",
		X"69",X"00",X"85",X"11",X"60",X"D8",X"38",X"A5",X"10",X"E9",X"28",X"85",X"10",X"A5",X"11",X"E9",
		X"00",X"85",X"11",X"60",X"4E",X"15",X"02",X"90",X"0B",X"A9",X"20",X"8D",X"15",X"02",X"E6",X"10",
		X"D0",X"02",X"E6",X"11",X"60",X"0E",X"15",X"02",X"2C",X"15",X"02",X"50",X"0F",X"A9",X"01",X"8D",
		X"15",X"02",X"C6",X"10",X"A5",X"10",X"C9",X"FF",X"D0",X"02",X"C6",X"11",X"60",X"A9",X"04",X"A2",
		X"E5",X"20",X"64",X"F2",X"B0",X"2A",X"AD",X"E5",X"02",X"8D",X"12",X"02",X"A9",X"F0",X"A2",X"E1",
		X"20",X"64",X"F2",X"B0",X"1B",X"A9",X"C8",X"A2",X"E3",X"20",X"64",X"F2",X"B0",X"12",X"AE",X"E1",
		X"02",X"8E",X"19",X"02",X"AC",X"E3",X"02",X"8C",X"1A",X"02",X"20",X"F6",X"ED",X"4C",X"63",X"F0",
		X"EE",X"E0",X"02",X"60",X"20",X"76",X"F2",X"B0",X"0C",X"AE",X"19",X"02",X"AC",X"1A",X"02",X"20",
		X"F6",X"ED",X"4C",X"78",X"F0",X"EE",X"E0",X"02",X"60",X"20",X"76",X"F2",X"B0",X"11",X"A2",X"04",
		X"BD",X"E0",X"02",X"9D",X"01",X"02",X"CA",X"D0",X"F7",X"20",X"06",X"EE",X"4C",X"92",X"F0",X"EE",
		X"E0",X"02",X"60",X"AE",X"E2",X"02",X"D0",X"09",X"AE",X"E1",X"02",X"8E",X"13",X"02",X"4C",X"A4",
		X"F0",X"EE",X"E0",X"02",X"60",X"AE",X"E2",X"02",X"D0",X"3D",X"AE",X"E1",X"02",X"E0",X"20",X"90",
		X"36",X"E0",X"80",X"B0",X"32",X"A9",X"02",X"A2",X"E3",X"20",X"64",X"F2",X"B0",X"29",X"A9",X"04",
		X"A2",X"E5",X"20",X"64",X"F2",X"B0",X"20",X"AD",X"19",X"02",X"C9",X"E9",X"B0",X"19",X"AD",X"1A",
		X"02",X"C9",X"C1",X"B0",X"12",X"20",X"EB",X"F0",X"20",X"15",X"F1",X"AE",X"19",X"02",X"AC",X"1A",
		X"02",X"20",X"A6",X"EF",X"4C",X"EA",X"F0",X"EE",X"E0",X"02",X"60",X"D8",X"AD",X"E5",X"02",X"8D",
		X"12",X"02",X"20",X"E3",X"ED",X"AD",X"E1",X"02",X"85",X"0C",X"A9",X"00",X"85",X"0D",X"A2",X"03",
		X"06",X"0C",X"26",X"0D",X"CA",X"D0",X"F9",X"AD",X"E3",X"02",X"0A",X"0A",X"18",X"69",X"98",X"18",
		X"65",X"0D",X"85",X"0D",X"60",X"A0",X"00",X"84",X"0F",X"B1",X"0C",X"85",X"0E",X"20",X"C3",X"F2",
		X"26",X"0E",X"26",X"0E",X"A2",X"06",X"26",X"0E",X"90",X"03",X"20",X"5B",X"EF",X"20",X"04",X"F0",
		X"CA",X"D0",X"F3",X"20",X"D4",X"F2",X"20",X"E6",X"EF",X"A4",X"0F",X"C8",X"C0",X"08",X"D0",X"D7",
		X"60",X"A9",X"F0",X"A2",X"E1",X"20",X"64",X"F2",X"B0",X"31",X"A9",X"C8",X"A2",X"E3",X"20",X"64",
		X"F2",X"B0",X"28",X"AE",X"E1",X"02",X"8E",X"19",X"02",X"AC",X"E3",X"02",X"8C",X"1A",X"02",X"20",
		X"A6",X"EF",X"A0",X"00",X"B1",X"10",X"2D",X"15",X"02",X"F0",X"05",X"A9",X"FF",X"4C",X"72",X"F1",
		X"A9",X"00",X"8D",X"E1",X"02",X"8D",X"E2",X"02",X"4C",X"7E",X"F1",X"EE",X"E0",X"02",X"60",X"A9",
		X"10",X"85",X"0C",X"A9",X"00",X"85",X"0D",X"20",X"97",X"F1",X"60",X"A9",X"00",X"85",X"0C",X"A9",
		X"01",X"85",X"0D",X"20",X"97",X"F1",X"60",X"A9",X"08",X"A2",X"E1",X"20",X"64",X"F2",X"B0",X"41",
		X"20",X"C3",X"F2",X"AD",X"E1",X"02",X"05",X"0C",X"8D",X"02",X"02",X"AE",X"1F",X"02",X"D0",X"12",
		X"A6",X"0D",X"9D",X"6B",X"02",X"A9",X"A8",X"18",X"65",X"0D",X"AA",X"A0",X"BB",X"A9",X"1B",X"4C",
		X"CC",X"F1",X"A9",X"00",X"18",X"65",X"0D",X"AA",X"A0",X"A0",X"A9",X"C8",X"8D",X"00",X"02",X"86",
		X"10",X"84",X"11",X"A9",X"01",X"8D",X"01",X"02",X"20",X"3A",X"F2",X"20",X"D4",X"F2",X"4C",X"E4",
		X"F1",X"EE",X"E0",X"02",X"60",X"D8",X"AD",X"E1",X"02",X"8D",X"00",X"02",X"F0",X"48",X"18",X"6D",
		X"1A",X"02",X"A8",X"AD",X"E2",X"02",X"69",X"00",X"D0",X"3C",X"C0",X"C9",X"B0",X"38",X"AD",X"E3",
		X"02",X"8D",X"01",X"02",X"F0",X"30",X"A0",X"00",X"AD",X"19",X"02",X"38",X"E9",X"06",X"90",X"04",
		X"C8",X"4C",X"0B",X"F2",X"98",X"18",X"6D",X"E3",X"02",X"A8",X"AD",X"E4",X"02",X"69",X"00",X"D0",
		X"15",X"C0",X"29",X"B0",X"11",X"AD",X"E6",X"02",X"D0",X"0C",X"AD",X"E5",X"02",X"8D",X"02",X"02",
		X"20",X"3A",X"F2",X"4C",X"39",X"F2",X"EE",X"E0",X"02",X"60",X"AD",X"02",X"02",X"A0",X"00",X"91",
		X"10",X"C8",X"CC",X"01",X"02",X"D0",X"F8",X"20",X"E6",X"EF",X"CE",X"00",X"02",X"D0",X"EB",X"60",
		X"8D",X"04",X"02",X"BD",X"01",X"02",X"D0",X"0A",X"BD",X"00",X"02",X"F0",X"05",X"CD",X"04",X"02",
		X"90",X"01",X"38",X"60",X"8D",X"04",X"02",X"BD",X"01",X"02",X"D0",X"08",X"BD",X"00",X"02",X"CD",
		X"04",X"02",X"90",X"01",X"38",X"60",X"A9",X"04",X"A2",X"E5",X"20",X"64",X"F2",X"B0",X"43",X"A9",
		X"00",X"8D",X"01",X"02",X"8D",X"03",X"02",X"AD",X"19",X"02",X"8D",X"00",X"02",X"AD",X"1A",X"02",
		X"8D",X"02",X"02",X"A2",X"00",X"A0",X"E1",X"20",X"95",X"EC",X"A9",X"F0",X"20",X"64",X"F2",X"B0",
		X"21",X"A2",X"02",X"A0",X"E3",X"20",X"95",X"EC",X"A9",X"C8",X"20",X"64",X"F2",X"B0",X"13",X"AD",
		X"E5",X"02",X"8D",X"12",X"02",X"AD",X"00",X"02",X"8D",X"19",X"02",X"AD",X"02",X"02",X"8D",X"1A",
		X"02",X"18",X"60",X"A5",X"10",X"8D",X"16",X"02",X"A5",X"11",X"8D",X"17",X"02",X"AD",X"15",X"02",
		X"8D",X"18",X"02",X"60",X"AD",X"16",X"02",X"85",X"10",X"AD",X"17",X"02",X"85",X"11",X"AD",X"18",
		X"02",X"8D",X"15",X"02",X"60",X"AD",X"E2",X"02",X"D0",X"43",X"AD",X"E1",X"02",X"F0",X"3E",X"AD",
		X"19",X"02",X"CD",X"E1",X"02",X"90",X"36",X"18",X"6D",X"E1",X"02",X"C9",X"F0",X"B0",X"2E",X"AD",
		X"1A",X"02",X"CD",X"E1",X"02",X"90",X"26",X"18",X"6D",X"E1",X"02",X"C9",X"C8",X"B0",X"1E",X"A2",
		X"E3",X"A9",X"04",X"20",X"64",X"F2",X"B0",X"15",X"AD",X"E3",X"02",X"8D",X"12",X"02",X"20",X"E3",
		X"ED",X"AD",X"13",X"02",X"8D",X"14",X"02",X"20",X"31",X"F3",X"4C",X"30",X"F3",X"EE",X"E0",X"02",
		X"60",X"20",X"C3",X"F2",X"AD",X"1A",X"02",X"38",X"ED",X"E1",X"02",X"A8",X"AE",X"19",X"02",X"20",
		X"A6",X"EF",X"AD",X"E1",X"02",X"85",X"0F",X"20",X"F0",X"F3",X"A9",X"80",X"8D",X"1B",X"02",X"8D",
		X"1D",X"02",X"A9",X"00",X"8D",X"1C",X"02",X"AD",X"E1",X"02",X"8D",X"1E",X"02",X"A9",X"00",X"85",
		X"0F",X"20",X"7F",X"F3",X"20",X"AF",X"F3",X"A5",X"0F",X"F0",X"03",X"20",X"4D",X"EF",X"AD",X"1C",
		X"02",X"D0",X"EA",X"AD",X"1E",X"02",X"CD",X"E1",X"02",X"D0",X"E2",X"20",X"D4",X"F2",X"60",X"AD",
		X"1D",X"02",X"AE",X"1E",X"02",X"20",X"DF",X"F3",X"A5",X"0C",X"18",X"6D",X"1B",X"02",X"8D",X"1B",
		X"02",X"AD",X"1C",X"02",X"85",X"0C",X"65",X"0D",X"8D",X"1C",X"02",X"C5",X"0C",X"F0",X"0F",X"B0",
		X"06",X"20",X"04",X"F0",X"4C",X"AA",X"F3",X"20",X"15",X"F0",X"A9",X"01",X"85",X"0F",X"60",X"AD",
		X"1B",X"02",X"AE",X"1C",X"02",X"20",X"DF",X"F3",X"38",X"AD",X"1D",X"02",X"E5",X"0C",X"8D",X"1D",
		X"02",X"AD",X"1E",X"02",X"85",X"0C",X"E5",X"0D",X"8D",X"1E",X"02",X"C5",X"0C",X"F0",X"0F",X"B0",
		X"06",X"20",X"E6",X"EF",X"4C",X"DA",X"F3",X"20",X"F5",X"EF",X"A9",X"01",X"85",X"0F",X"60",X"85",
		X"0C",X"86",X"0D",X"A6",X"0E",X"A5",X"0D",X"2A",X"66",X"0D",X"66",X"0C",X"CA",X"D0",X"F6",X"60",
		X"E6",X"0F",X"A9",X"00",X"85",X"0E",X"A9",X"01",X"0A",X"E6",X"0E",X"C5",X"0F",X"90",X"F9",X"60",
		X"4C",X"00",X"F7",X"4C",X"CB",X"F7",X"4C",X"35",X"F5",X"4C",X"3F",X"F7",X"4C",X"E0",X"F7",X"4C",
		X"3C",X"F4",X"4C",X"85",X"FA",X"4C",X"9B",X"FA",X"4C",X"B1",X"FA",X"4C",X"C7",X"FA",X"4C",X"26",
		X"FB",X"4C",X"B6",X"FB",X"4C",X"FE",X"FB",X"4C",X"23",X"F9",X"4C",X"E3",X"F8",X"4C",X"4A",X"F8",
		X"4C",X"82",X"F8",X"4C",X"7B",X"F5",X"4C",X"2F",X"F8",X"4C",X"60",X"F9",X"48",X"08",X"98",X"48",
		X"D8",X"AD",X"08",X"02",X"10",X"1D",X"29",X"87",X"8D",X"10",X"02",X"AE",X"0A",X"02",X"20",X"06",
		X"F5",X"CD",X"10",X"02",X"D0",X"0D",X"CE",X"0E",X"02",X"D0",X"31",X"A9",X"04",X"8D",X"0E",X"02",
		X"4C",X"6B",X"F4",X"A9",X"20",X"8D",X"0E",X"02",X"20",X"C8",X"F4",X"20",X"94",X"F4",X"AA",X"10",
		X"1D",X"48",X"AD",X"6A",X"02",X"29",X"08",X"D0",X"0F",X"68",X"48",X"C9",X"A0",X"90",X"06",X"20",
		X"FA",X"FA",X"4C",X"88",X"F4",X"20",X"10",X"FB",X"68",X"4C",X"8E",X"F4",X"A9",X"00",X"AA",X"68",
		X"A8",X"28",X"68",X"60",X"AD",X"09",X"02",X"A8",X"A9",X"00",X"C0",X"A4",X"F0",X"04",X"C0",X"A7",
		X"D0",X"03",X"18",X"69",X"40",X"18",X"6D",X"08",X"02",X"10",X"1C",X"29",X"7F",X"AA",X"BD",X"70",
		X"FF",X"2D",X"0C",X"02",X"10",X"03",X"38",X"E9",X"20",X"29",X"7F",X"C0",X"A2",X"D0",X"06",X"C9",
		X"40",X"30",X"02",X"29",X"1F",X"09",X"80",X"60",X"A9",X"38",X"8D",X"0D",X"02",X"8D",X"08",X"02",
		X"8D",X"09",X"02",X"A9",X"7F",X"48",X"68",X"48",X"AA",X"A9",X"07",X"20",X"06",X"F5",X"0D",X"0D",
		X"02",X"10",X"12",X"A2",X"00",X"A0",X"20",X"CC",X"0D",X"02",X"D0",X"01",X"E8",X"9D",X"08",X"02",
		X"68",X"48",X"9D",X"0A",X"02",X"38",X"68",X"6A",X"48",X"38",X"AD",X"0D",X"02",X"E9",X"08",X"8D",
		X"0D",X"02",X"10",X"D2",X"68",X"60",X"48",X"A9",X"0E",X"20",X"35",X"F5",X"68",X"29",X"07",X"AA",
		X"8D",X"11",X"02",X"09",X"B8",X"8D",X"00",X"03",X"A0",X"04",X"88",X"D0",X"FD",X"AD",X"00",X"03",
		X"29",X"08",X"D0",X"0D",X"CA",X"8A",X"29",X"07",X"AA",X"CD",X"11",X"02",X"D0",X"E5",X"A9",X"00",
		X"60",X"8A",X"09",X"80",X"60",X"08",X"78",X"8D",X"0F",X"03",X"C9",X"07",X"D0",X"06",X"8A",X"09",
		X"40",X"4C",X"45",X"F5",X"8A",X"48",X"A2",X"0C",X"A0",X"EE",X"A9",X"11",X"20",X"6A",X"F5",X"A0",
		X"CC",X"A9",X"11",X"20",X"6A",X"F5",X"68",X"8D",X"0F",X"03",X"A0",X"EC",X"A9",X"11",X"20",X"6A",
		X"F5",X"A0",X"CC",X"A9",X"11",X"20",X"6A",X"F5",X"28",X"60",X"08",X"78",X"3D",X"00",X"03",X"8D",
		X"0F",X"02",X"98",X"0D",X"0F",X"02",X"9D",X"00",X"03",X"28",X"60",X"8D",X"01",X"03",X"A2",X"00",
		X"A0",X"00",X"A9",X"EF",X"20",X"6A",X"F5",X"A0",X"10",X"A9",X"FF",X"20",X"6A",X"F5",X"A9",X"02",
		X"A2",X"05",X"A0",X"DC",X"20",X"D3",X"EB",X"AD",X"0D",X"03",X"29",X"02",X"D0",X"0F",X"A9",X"02",
		X"20",X"D6",X"EB",X"98",X"D0",X"F1",X"8A",X"D0",X"EE",X"A9",X"FF",X"30",X"05",X"AD",X"0D",X"03",
		X"A9",X"00",X"60",X"6E",X"6E",X"6E",X"6E",X"48",X"6E",X"4B",X"6B",X"00",X"10",X"1D",X"0A",X"32",
		X"23",X"29",X"6E",X"4C",X"4E",X"6E",X"4D",X"58",X"6E",X"6E",X"6E",X"6E",X"6E",X"4A",X"4A",X"6E",
		X"49",X"3F",X"6E",X"29",X"1F",X"AA",X"BD",X"B3",X"F5",X"18",X"69",X"F2",X"8D",X"61",X"02",X"A9",
		X"00",X"69",X"F5",X"8D",X"62",X"02",X"78",X"A9",X"00",X"20",X"CB",X"F7",X"38",X"A9",X"00",X"6C",
		X"61",X"02",X"CE",X"69",X"02",X"10",X"2A",X"A9",X"27",X"8D",X"69",X"02",X"CE",X"68",X"02",X"4C",
		X"7D",X"F6",X"EE",X"69",X"02",X"A2",X"27",X"EC",X"69",X"02",X"10",X"15",X"8D",X"69",X"02",X"EE",
		X"68",X"02",X"4C",X"7D",X"F6",X"8D",X"69",X"02",X"4C",X"CC",X"F6",X"AD",X"68",X"02",X"20",X"D3",
		X"F6",X"4C",X"CC",X"F6",X"AA",X"E8",X"8A",X"20",X"D3",X"F6",X"EC",X"6F",X"02",X"D0",X"F6",X"A9",
		X"00",X"8D",X"69",X"02",X"8D",X"68",X"02",X"F0",X"D6",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",
		X"2A",X"4D",X"6A",X"02",X"8D",X"6A",X"02",X"4C",X"CC",X"F6",X"AD",X"0C",X"02",X"49",X"80",X"8D",
		X"0C",X"02",X"AD",X"1F",X"02",X"D0",X"03",X"20",X"29",X"F7",X"4C",X"CC",X"F6",X"20",X"85",X"FA",
		X"18",X"90",X"69",X"07",X"50",X"52",X"49",X"4E",X"54",X"00",X"07",X"20",X"20",X"20",X"20",X"20",
		X"00",X"07",X"43",X"41",X"50",X"53",X"00",X"07",X"20",X"20",X"20",X"20",X"00",X"AD",X"68",X"02",
		X"20",X"F1",X"F6",X"85",X"12",X"84",X"13",X"AE",X"6F",X"02",X"CA",X"8A",X"20",X"00",X"F7",X"8D",
		X"04",X"02",X"8C",X"05",X"02",X"AE",X"68",X"02",X"F0",X"0F",X"CA",X"EC",X"6F",X"02",X"D0",X"2C",
		X"CE",X"68",X"02",X"A9",X"01",X"A2",X"02",X"D0",X"07",X"EE",X"68",X"02",X"A9",X"02",X"A2",X"01",
		X"20",X"F1",X"F6",X"8D",X"02",X"02",X"8C",X"03",X"02",X"8A",X"20",X"F1",X"F6",X"8D",X"00",X"02",
		X"8C",X"01",X"02",X"20",X"D9",X"EB",X"AD",X"68",X"02",X"20",X"D3",X"F6",X"A9",X"01",X"20",X"CB",
		X"F7",X"58",X"60",X"20",X"F1",X"F6",X"85",X"12",X"84",X"13",X"A0",X"27",X"A9",X"20",X"91",X"12",
		X"88",X"10",X"FB",X"A0",X"00",X"AD",X"6B",X"02",X"91",X"12",X"AD",X"6C",X"02",X"C8",X"91",X"12",
		X"60",X"20",X"00",X"F7",X"18",X"6D",X"6D",X"02",X"48",X"98",X"6D",X"6E",X"02",X"A8",X"68",X"60",
		X"A0",X"00",X"8C",X"63",X"02",X"8D",X"64",X"02",X"0A",X"2E",X"63",X"02",X"0A",X"2E",X"63",X"02",
		X"18",X"6D",X"64",X"02",X"90",X"03",X"EE",X"63",X"02",X"0A",X"2E",X"63",X"02",X"0A",X"2E",X"63",
		X"02",X"0A",X"2E",X"63",X"02",X"AC",X"63",X"02",X"60",X"AD",X"0C",X"02",X"10",X"07",X"A9",X"71",
		X"A0",X"F6",X"4C",X"39",X"F7",X"A9",X"77",X"A0",X"F6",X"A2",X"23",X"20",X"2F",X"F8",X"60",X"48",
		X"08",X"98",X"48",X"8A",X"48",X"D8",X"C9",X"20",X"90",X"4B",X"AD",X"6A",X"02",X"29",X"02",X"F0",
		X"47",X"AD",X"6A",X"02",X"29",X"10",X"F0",X"13",X"8A",X"38",X"E9",X"40",X"30",X"09",X"29",X"1F",
		X"20",X"AC",X"F7",X"A9",X"1B",X"D0",X"2E",X"A9",X"20",X"10",X"F5",X"E0",X"7F",X"F0",X"15",X"20",
		X"9F",X"F7",X"F0",X"08",X"68",X"48",X"20",X"AC",X"F7",X"4C",X"98",X"F7",X"A9",X"09",X"20",X"D3",
		X"F5",X"4C",X"6F",X"F7",X"A9",X"08",X"20",X"D3",X"F5",X"20",X"9F",X"F7",X"F0",X"F6",X"A9",X"20",
		X"20",X"AC",X"F7",X"A9",X"08",X"20",X"D3",X"F5",X"68",X"AA",X"68",X"A8",X"28",X"68",X"60",X"AD",
		X"69",X"02",X"29",X"FE",X"D0",X"05",X"AD",X"6A",X"02",X"29",X"20",X"60",X"48",X"AC",X"69",X"02",
		X"91",X"12",X"AD",X"6A",X"02",X"29",X"40",X"F0",X"0B",X"AD",X"69",X"02",X"18",X"69",X"28",X"A8",
		X"68",X"48",X"91",X"12",X"A9",X"09",X"20",X"D3",X"F5",X"68",X"60",X"2D",X"6A",X"02",X"4A",X"6A",
		X"8D",X"65",X"02",X"AC",X"69",X"02",X"B1",X"12",X"29",X"7F",X"0D",X"65",X"02",X"91",X"12",X"60",
		X"A9",X"00",X"85",X"0C",X"A9",X"B9",X"85",X"0D",X"A9",X"00",X"20",X"F7",X"F7",X"A0",X"BA",X"84",
		X"0D",X"A9",X"20",X"20",X"F7",X"F7",X"60",X"A0",X"00",X"48",X"20",X"1E",X"F8",X"91",X"0C",X"C8",
		X"68",X"48",X"20",X"1C",X"F8",X"68",X"48",X"20",X"1A",X"F8",X"91",X"0C",X"C8",X"C0",X"00",X"F0",
		X"07",X"68",X"18",X"69",X"01",X"4C",X"F9",X"F7",X"68",X"60",X"4A",X"4A",X"4A",X"4A",X"29",X"03",
		X"AA",X"BD",X"2B",X"F8",X"91",X"0C",X"C8",X"91",X"0C",X"C8",X"60",X"00",X"F0",X"0F",X"FF",X"85",
		X"0C",X"84",X"0D",X"A0",X"00",X"B1",X"0C",X"F0",X"07",X"9D",X"80",X"BB",X"E8",X"C8",X"D0",X"F5",
		X"60",X"4C",X"03",X"EC",X"4C",X"30",X"F4",X"01",X"00",X"40",X"A2",X"FF",X"9A",X"58",X"D8",X"A2",
		X"08",X"BD",X"41",X"F8",X"9D",X"28",X"02",X"CA",X"10",X"F7",X"20",X"C0",X"F9",X"08",X"20",X"88",
		X"F8",X"28",X"F0",X"0D",X"A0",X"00",X"BE",X"74",X"F8",X"20",X"3F",X"F7",X"C8",X"C0",X"0E",X"D0",
		X"F5",X"4C",X"00",X"C0",X"4D",X"45",X"4D",X"4F",X"52",X"59",X"20",X"45",X"52",X"52",X"4F",X"52",
		X"0D",X"0A",X"20",X"88",X"F8",X"4C",X"03",X"C0",X"20",X"60",X"F9",X"A9",X"07",X"A2",X"40",X"20",
		X"06",X"F4",X"20",X"D0",X"EB",X"20",X"D1",X"F8",X"20",X"7F",X"F9",X"A2",X"05",X"20",X"3E",X"F9",
		X"20",X"0C",X"F4",X"A9",X"FF",X"8D",X"0C",X"02",X"60",X"48",X"8A",X"48",X"A9",X"00",X"8D",X"69",
		X"02",X"A9",X"01",X"8D",X"1F",X"02",X"8D",X"68",X"02",X"A9",X"40",X"8D",X"6D",X"02",X"A9",X"BF",
		X"8D",X"6E",X"02",X"A9",X"03",X"8D",X"6F",X"02",X"A2",X"0C",X"20",X"09",X"F4",X"68",X"AA",X"68",
		X"60",X"48",X"A9",X"03",X"8D",X"6A",X"02",X"A9",X"00",X"8D",X"6C",X"02",X"A9",X"17",X"8D",X"6B",
		X"02",X"68",X"60",X"48",X"AD",X"1F",X"02",X"D0",X"05",X"A2",X"0B",X"20",X"3E",X"F9",X"A9",X"FE",
		X"2D",X"6A",X"02",X"8D",X"6A",X"02",X"A9",X"1E",X"20",X"B3",X"F9",X"20",X"00",X"EC",X"A9",X"00",
		X"8D",X"19",X"02",X"8D",X"1A",X"02",X"85",X"10",X"A9",X"A0",X"85",X"11",X"A9",X"20",X"8D",X"15",
		X"02",X"A9",X"FF",X"8D",X"13",X"02",X"20",X"A9",X"F8",X"A9",X"01",X"0D",X"6A",X"02",X"8D",X"6A",
		X"02",X"68",X"60",X"48",X"A9",X"FE",X"2D",X"6A",X"02",X"8D",X"6A",X"02",X"A2",X"11",X"20",X"3E",
		X"F9",X"20",X"7F",X"F9",X"A9",X"01",X"0D",X"6A",X"02",X"8D",X"6A",X"02",X"68",X"60",X"A0",X"06",
		X"BD",X"4E",X"F9",X"99",X"FF",X"01",X"CA",X"88",X"D0",X"F6",X"20",X"D9",X"EB",X"60",X"70",X"FC",
		X"00",X"B5",X"00",X"03",X"00",X"B4",X"00",X"98",X"80",X"07",X"00",X"98",X"00",X"B4",X"80",X"07",
		X"A9",X"FF",X"8D",X"03",X"03",X"A9",X"F7",X"8D",X"02",X"03",X"A9",X"B7",X"8D",X"00",X"03",X"A9",
		X"DD",X"8D",X"0C",X"03",X"A9",X"7F",X"8D",X"0E",X"03",X"A9",X"00",X"8D",X"0B",X"03",X"60",X"A9",
		X"1A",X"20",X"B3",X"F9",X"A9",X"20",X"A0",X"28",X"99",X"7F",X"BB",X"88",X"D0",X"FA",X"A9",X"00",
		X"8D",X"1F",X"02",X"8D",X"69",X"02",X"A9",X"01",X"8D",X"68",X"02",X"A9",X"80",X"8D",X"6D",X"02",
		X"A9",X"BB",X"8D",X"6E",X"02",X"A9",X"1B",X"8D",X"6F",X"02",X"A2",X"0C",X"20",X"09",X"F4",X"20",
		X"29",X"F7",X"60",X"8D",X"DF",X"BF",X"A9",X"02",X"A2",X"00",X"A0",X"03",X"20",X"DC",X"EB",X"60",
		X"20",X"DD",X"F9",X"20",X"06",X"FA",X"D0",X"14",X"A9",X"00",X"85",X"0C",X"A9",X"10",X"85",X"0D",
		X"A9",X"00",X"20",X"49",X"FA",X"D0",X"05",X"A9",X"FF",X"20",X"49",X"FA",X"60",X"A9",X"00",X"8D",
		X"00",X"10",X"A9",X"FF",X"8D",X"00",X"50",X"AD",X"00",X"10",X"D0",X"0A",X"A9",X"00",X"8D",X"20",
		X"02",X"A9",X"BF",X"4C",X"FD",X"F9",X"A9",X"01",X"8D",X"20",X"02",X"A9",X"3F",X"8D",X"E2",X"02",
		X"A9",X"FF",X"8D",X"E1",X"02",X"60",X"18",X"AD",X"E1",X"02",X"69",X"01",X"85",X"0E",X"AD",X"E2",
		X"02",X"69",X"00",X"85",X"0F",X"A9",X"00",X"85",X"0C",X"A9",X"04",X"85",X"0D",X"A0",X"00",X"A5",
		X"0E",X"C5",X"0C",X"D0",X"06",X"A5",X"0F",X"C5",X"0D",X"F0",X"1D",X"A9",X"AA",X"91",X"0C",X"B1",
		X"0C",X"C9",X"AA",X"D0",X"13",X"A9",X"55",X"91",X"0C",X"B1",X"0C",X"C9",X"55",X"D0",X"09",X"E6",
		X"0C",X"D0",X"02",X"E6",X"0D",X"4C",X"1F",X"FA",X"60",X"85",X"0E",X"A0",X"00",X"91",X"0C",X"88",
		X"D0",X"FB",X"20",X"61",X"FA",X"A0",X"00",X"B1",X"0C",X"C5",X"0E",X"D0",X"03",X"88",X"D0",X"F7",
		X"60",X"A2",X"06",X"A0",X"00",X"88",X"D0",X"FD",X"CA",X"D0",X"FA",X"60",X"08",X"78",X"86",X"14",
		X"84",X"15",X"A0",X"00",X"B1",X"14",X"AA",X"98",X"48",X"20",X"35",X"F5",X"68",X"A8",X"C8",X"C0",
		X"0E",X"D0",X"F1",X"28",X"60",X"A2",X"8D",X"A0",X"FA",X"20",X"6C",X"FA",X"60",X"18",X"00",X"00",
		X"00",X"00",X"00",X"00",X"3E",X"10",X"00",X"00",X"00",X"0F",X"00",X"A2",X"A3",X"A0",X"FA",X"20",
		X"6C",X"FA",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"07",X"10",X"10",X"10",X"00",X"08",
		X"00",X"A2",X"B9",X"A0",X"FA",X"20",X"6C",X"FA",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",
		X"07",X"10",X"10",X"10",X"00",X"18",X"00",X"A2",X"EC",X"A0",X"FA",X"20",X"6C",X"FA",X"A9",X"00",
		X"AA",X"8A",X"48",X"A9",X"00",X"20",X"35",X"F5",X"A2",X"00",X"CA",X"D0",X"FD",X"68",X"AA",X"E8",
		X"E0",X"70",X"D0",X"ED",X"A9",X"08",X"A2",X"00",X"20",X"35",X"F5",X"60",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"3E",X"0F",X"00",X"00",X"00",X"00",X"00",X"A2",X"02",X"A0",X"FB",X"20",X"6C",
		X"FA",X"60",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"10",X"00",X"00",X"1F",X"00",X"00",
		X"A2",X"18",X"A0",X"FB",X"20",X"6C",X"FA",X"60",X"2F",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",
		X"10",X"00",X"00",X"1F",X"00",X"00",X"AD",X"E1",X"02",X"C9",X"01",X"D0",X"22",X"A9",X"00",X"AE",
		X"E3",X"02",X"20",X"35",X"F5",X"A9",X"01",X"AE",X"E4",X"02",X"20",X"35",X"F5",X"AD",X"E5",X"02",
		X"29",X"0F",X"D0",X"04",X"A2",X"10",X"D0",X"01",X"AA",X"A9",X"08",X"20",X"35",X"F5",X"60",X"C9",
		X"02",X"D0",X"22",X"A9",X"02",X"AE",X"E3",X"02",X"20",X"35",X"F5",X"A9",X"03",X"AE",X"E4",X"02",
		X"20",X"35",X"F5",X"AD",X"E5",X"02",X"29",X"0F",X"D0",X"04",X"A2",X"10",X"D0",X"01",X"AA",X"A9",
		X"09",X"20",X"35",X"F5",X"60",X"C9",X"03",X"D0",X"22",X"A9",X"04",X"AE",X"E3",X"02",X"20",X"35",
		X"F5",X"A9",X"05",X"AE",X"E4",X"02",X"20",X"35",X"F5",X"AD",X"E5",X"02",X"29",X"0F",X"D0",X"04",
		X"A2",X"10",X"D0",X"01",X"AA",X"A9",X"0A",X"20",X"35",X"F5",X"60",X"A9",X"06",X"AE",X"E3",X"02",
		X"20",X"35",X"F5",X"AD",X"E1",X"02",X"C9",X"04",X"F0",X"93",X"C9",X"05",X"F0",X"B5",X"C9",X"06",
		X"F0",X"D7",X"EE",X"E0",X"02",X"60",X"AD",X"E3",X"02",X"0A",X"0A",X"0A",X"0D",X"E1",X"02",X"49",
		X"3F",X"AA",X"A9",X"07",X"20",X"35",X"F5",X"18",X"AD",X"E7",X"02",X"0A",X"8D",X"E7",X"02",X"AD",
		X"E8",X"02",X"2A",X"8D",X"E8",X"02",X"A9",X"0B",X"AE",X"E7",X"02",X"20",X"35",X"F5",X"A9",X"0C",
		X"AE",X"E8",X"02",X"20",X"35",X"F5",X"AD",X"E5",X"02",X"29",X"07",X"A8",X"B9",X"F6",X"FB",X"AA",
		X"A9",X"0D",X"20",X"35",X"F5",X"60",X"00",X"00",X"04",X"08",X"0A",X"0B",X"0C",X"0D",X"A2",X"E1",
		X"A9",X"04",X"20",X"09",X"EC",X"B0",X"39",X"A2",X"E3",X"A9",X"08",X"20",X"06",X"EC",X"B0",X"30",
		X"A2",X"E5",X"A9",X"0D",X"20",X"09",X"EC",X"B0",X"27",X"AC",X"E3",X"02",X"AE",X"E5",X"02",X"BD",
		X"44",X"FC",X"8D",X"E4",X"02",X"BD",X"51",X"FC",X"8D",X"E3",X"02",X"AD",X"E7",X"02",X"8D",X"E5",
		X"02",X"88",X"30",X"09",X"4E",X"E4",X"02",X"6E",X"E3",X"02",X"4C",X"31",X"FC",X"4C",X"26",X"FB",
		X"EE",X"E0",X"02",X"60",X"00",X"07",X"07",X"06",X"06",X"05",X"05",X"05",X"04",X"04",X"04",X"04",
		X"03",X"00",X"77",X"0B",X"A6",X"47",X"EC",X"97",X"47",X"FB",X"B3",X"70",X"30",X"F4",X"20",X"0F",
		X"F4",X"8A",X"10",X"03",X"8E",X"DF",X"02",X"4C",X"4F",X"ED",X"4C",X"67",X"B3",X"4C",X"7B",X"B3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"08",X"08",X"00",X"08",X"00",
		X"14",X"14",X"14",X"00",X"00",X"00",X"00",X"00",X"14",X"14",X"3E",X"14",X"3E",X"14",X"14",X"00",
		X"08",X"1E",X"28",X"1C",X"0A",X"3C",X"08",X"00",X"30",X"32",X"04",X"08",X"10",X"26",X"06",X"00",
		X"10",X"28",X"28",X"10",X"2A",X"24",X"1A",X"00",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",
		X"08",X"10",X"20",X"20",X"20",X"10",X"08",X"00",X"08",X"04",X"02",X"02",X"02",X"04",X"08",X"00",
		X"08",X"2A",X"1C",X"08",X"1C",X"2A",X"08",X"00",X"00",X"08",X"08",X"3E",X"08",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"10",X"00",X"00",X"00",X"3E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"02",X"04",X"08",X"10",X"20",X"00",X"00",
		X"1C",X"22",X"26",X"2A",X"32",X"22",X"1C",X"00",X"08",X"18",X"08",X"08",X"08",X"08",X"1C",X"00",
		X"1C",X"22",X"02",X"04",X"08",X"10",X"3E",X"00",X"3E",X"02",X"04",X"0C",X"02",X"22",X"1C",X"00",
		X"04",X"0C",X"14",X"24",X"3E",X"04",X"04",X"00",X"3E",X"20",X"3C",X"02",X"02",X"22",X"1C",X"00",
		X"0C",X"10",X"20",X"3C",X"22",X"22",X"1C",X"00",X"3E",X"02",X"04",X"08",X"10",X"10",X"10",X"00",
		X"1C",X"22",X"22",X"1C",X"22",X"22",X"1C",X"00",X"1C",X"22",X"22",X"1E",X"02",X"04",X"18",X"00",
		X"00",X"00",X"08",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"08",X"08",X"10",
		X"04",X"08",X"10",X"20",X"10",X"08",X"04",X"00",X"00",X"00",X"3E",X"00",X"3E",X"00",X"00",X"00",
		X"10",X"08",X"04",X"02",X"04",X"08",X"10",X"00",X"1C",X"22",X"04",X"08",X"08",X"00",X"08",X"00",
		X"1C",X"22",X"2A",X"2E",X"2C",X"20",X"1E",X"00",X"08",X"14",X"22",X"22",X"3E",X"22",X"22",X"00",
		X"3C",X"22",X"22",X"3C",X"22",X"22",X"3C",X"00",X"1C",X"22",X"20",X"20",X"20",X"22",X"1C",X"00",
		X"3C",X"22",X"22",X"22",X"22",X"22",X"3C",X"00",X"3E",X"20",X"20",X"3C",X"20",X"20",X"3E",X"00",
		X"3E",X"20",X"20",X"3C",X"20",X"20",X"20",X"00",X"1E",X"20",X"20",X"20",X"26",X"22",X"1E",X"00",
		X"22",X"22",X"22",X"3E",X"22",X"22",X"22",X"00",X"1C",X"08",X"08",X"08",X"08",X"08",X"1C",X"00",
		X"02",X"02",X"02",X"02",X"02",X"22",X"1C",X"00",X"22",X"24",X"28",X"30",X"28",X"24",X"22",X"00",
		X"20",X"20",X"20",X"20",X"20",X"20",X"3E",X"00",X"22",X"36",X"2A",X"2A",X"22",X"22",X"22",X"00",
		X"22",X"22",X"32",X"2A",X"26",X"22",X"22",X"00",X"1C",X"22",X"22",X"22",X"22",X"22",X"1C",X"00",
		X"3C",X"22",X"22",X"3C",X"20",X"20",X"20",X"00",X"1C",X"22",X"22",X"22",X"2A",X"24",X"1A",X"00",
		X"3C",X"22",X"22",X"3C",X"28",X"24",X"22",X"00",X"1C",X"22",X"20",X"1C",X"02",X"22",X"1C",X"00",
		X"3E",X"08",X"08",X"08",X"08",X"08",X"08",X"00",X"22",X"22",X"22",X"22",X"22",X"22",X"1C",X"00",
		X"22",X"22",X"22",X"22",X"22",X"14",X"08",X"00",X"22",X"22",X"22",X"2A",X"2A",X"36",X"22",X"00",
		X"22",X"22",X"14",X"08",X"14",X"22",X"22",X"00",X"22",X"22",X"14",X"08",X"08",X"08",X"08",X"00",
		X"3E",X"02",X"04",X"08",X"10",X"20",X"3E",X"00",X"1E",X"10",X"10",X"10",X"10",X"10",X"1E",X"00",
		X"00",X"20",X"10",X"08",X"04",X"02",X"00",X"00",X"3C",X"04",X"04",X"04",X"04",X"04",X"3C",X"00",
		X"08",X"14",X"2A",X"08",X"08",X"08",X"08",X"00",X"0E",X"10",X"10",X"10",X"3C",X"10",X"3E",X"00",
		X"0C",X"12",X"2D",X"29",X"29",X"2D",X"12",X"0C",X"00",X"00",X"1C",X"02",X"1E",X"22",X"1E",X"00",
		X"20",X"20",X"3C",X"22",X"22",X"22",X"3C",X"00",X"00",X"00",X"1E",X"20",X"20",X"20",X"1E",X"00",
		X"02",X"02",X"1E",X"22",X"22",X"22",X"1E",X"00",X"00",X"00",X"1C",X"22",X"3E",X"20",X"1E",X"00",
		X"0C",X"12",X"10",X"3C",X"10",X"10",X"10",X"00",X"00",X"00",X"1C",X"22",X"22",X"1E",X"02",X"1C",
		X"20",X"20",X"3C",X"22",X"22",X"22",X"22",X"00",X"08",X"00",X"18",X"08",X"08",X"08",X"1C",X"00",
		X"04",X"00",X"0C",X"04",X"04",X"04",X"24",X"18",X"20",X"20",X"22",X"24",X"38",X"24",X"22",X"00",
		X"18",X"08",X"08",X"08",X"08",X"08",X"1C",X"00",X"00",X"00",X"36",X"2A",X"2A",X"2A",X"22",X"00",
		X"00",X"00",X"3C",X"22",X"22",X"22",X"22",X"00",X"00",X"00",X"1C",X"22",X"22",X"22",X"1C",X"00",
		X"00",X"00",X"3C",X"22",X"22",X"3C",X"20",X"20",X"00",X"00",X"1E",X"22",X"22",X"1E",X"02",X"02",
		X"00",X"00",X"2E",X"30",X"20",X"20",X"20",X"00",X"00",X"00",X"1E",X"20",X"1C",X"02",X"3C",X"00",
		X"10",X"10",X"3C",X"10",X"10",X"12",X"0C",X"00",X"00",X"00",X"22",X"22",X"22",X"26",X"1A",X"00",
		X"00",X"00",X"22",X"22",X"22",X"14",X"08",X"00",X"00",X"00",X"22",X"22",X"2A",X"2A",X"36",X"00",
		X"00",X"00",X"22",X"14",X"08",X"14",X"22",X"00",X"00",X"00",X"22",X"22",X"22",X"1E",X"02",X"1C",
		X"00",X"00",X"3E",X"04",X"08",X"10",X"3E",X"00",X"0E",X"18",X"18",X"30",X"18",X"18",X"0E",X"00",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"38",X"0C",X"0C",X"06",X"0C",X"0C",X"38",X"00",
		X"2A",X"15",X"2A",X"15",X"2A",X"15",X"2A",X"15",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"37",X"EA",X"ED",X"EB",X"20",X"F5",X"F9",X"38",X"EE",X"F4",X"36",X"39",X"2C",X"E9",X"E8",X"EC",
		X"35",X"F2",X"E2",X"3B",X"2E",X"EF",X"E7",X"30",X"F6",X"E6",X"34",X"2D",X"0B",X"F0",X"E5",X"2F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"31",X"1B",X"FA",X"00",X"08",X"7F",X"E1",X"0D",
		X"F8",X"F1",X"32",X"5C",X"0A",X"5D",X"F3",X"00",X"33",X"E4",X"E3",X"27",X"09",X"5B",X"F7",X"3D",
		X"26",X"4A",X"4D",X"4B",X"20",X"55",X"59",X"2A",X"4E",X"54",X"5E",X"28",X"3C",X"49",X"48",X"4C",
		X"25",X"52",X"42",X"3A",X"3E",X"4F",X"47",X"29",X"56",X"46",X"24",X"5F",X"0B",X"50",X"45",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"1B",X"5A",X"00",X"08",X"7F",X"41",X"0D",
		X"58",X"51",X"40",X"7C",X"0A",X"7D",X"53",X"00",X"23",X"44",X"43",X"22",X"09",X"7B",X"57",X"2B",
		X"A0",X"E8",X"B7",X"B7",X"BA",X"A4",X"A3",X"A0",X"B0",X"C4",X"2B",X"02",X"2D",X"F4",X"28",X"02");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
