library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity col1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(7 downto 0);
	data : out std_logic_vector(3 downto 0)
);
end entity;

architecture prom of col1 is
	type rom is array(0 to  255) of std_logic_vector(3 downto 0);
	signal rom_data: rom := (
		"1111","0110","1110","0001","1111","0000","0001","0000","1111","0000","0001","1111","1111","1111","0001","1110",
		"1111","0001","0000","0001","1111","0000","0001","0000","1111","0001","1111","1110","1111","0101","0000","0000",
		"1111","0101","0000","0001","1111","0000","0001","0001","1111","1111","0000","0001","1111","1111","0001","0000",
		"1111","0000","1110","1111","1111","0001","0000","0001","1111","0010","0000","1111","1111","0000","0001","1111",
		"1111","0110","1110","0001","1111","0000","0001","0000","1111","0000","0001","1111","1111","0001","0000","0000",
		"1111","0001","0000","0000","1111","0001","0000","0000","1111","0001","0000","0000","1111","0101","0000","0000",
		"1111","0101","0000","0001","1111","0000","0001","0001","1111","1111","0000","0001","1111","1111","0001","0000",
		"1111","0000","1110","1111","1111","0001","0000","0001","1111","0010","0000","1111","1111","0000","0001","1111",
		"1111","0110","1110","0001","1111","0000","0001","0000","1111","0000","0001","1111","1111","0001","0111","1110",
		"1111","0001","0111","1110","1111","0001","0111","1110","1111","0001","0111","1110","1111","0101","0000","0000",
		"1111","0101","0000","0001","1111","0000","0001","0001","1111","1111","0000","0001","1111","1111","0001","0000",
		"1111","0000","1110","1111","1111","0001","0000","0001","1111","0010","0000","1111","1111","0000","0001","1111",
		"1111","0110","1110","0001","1111","0000","0001","0000","1111","0000","0001","1111","1111","1111","1110","0000",
		"1111","1111","1110","0000","1111","1111","1110","0000","1111","1111","1110","0000","1111","0101","0000","0000",
		"1111","0101","0000","0001","1111","0000","0001","0001","1111","1111","0000","0001","1111","1111","0001","0000",
		"1111","0000","1110","1111","1111","0001","0000","0001","1111","0010","0000","1111","1111","0000","0001","1111");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
