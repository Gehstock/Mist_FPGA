library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity GALAXIAN_1H is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of GALAXIAN_1H is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"22",X"3E",X"00",X"3E",X"2A",X"2A",X"2A",X"00",X"00",X"3E",X"22",X"22",X"3E",X"00",X"3E",X"22",
		X"22",X"3E",X"00",X"02",X"3E",X"22",X"00",X"00",X"00",X"3E",X"22",X"22",X"3E",X"00",X"3E",X"22",
		X"C0",X"E0",X"E0",X"F0",X"70",X"70",X"78",X"78",X"03",X"07",X"07",X"0F",X"0E",X"0E",X"1E",X"1E",
		X"3C",X"3C",X"3E",X"1F",X"1F",X"0F",X"07",X"03",X"3C",X"3C",X"7C",X"F8",X"F8",X"F0",X"E0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"43",X"12",X"06",X"0C",X"38",X"7A",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"01",X"00",X"00",X"00",X"60",X"E0",X"F0",X"F0",X"FC",
		X"03",X"07",X"0F",X"0E",X"00",X"00",X"00",X"00",X"E0",X"E0",X"30",X"18",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"40",X"E0",X"F0",X"E0",
		X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"06",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"8F",X"FF",X"7F",X"3F",X"7F",X"FF",X"FF",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"08",X"18",X"7D",X"00",X"00",X"00",X"00",X"00",X"40",X"C0",X"80",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"C0",X"F0",X"F0",X"E0",X"C0",X"C0",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"7F",X"3F",X"3F",X"3F",X"7F",X"FF",X"EF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"E7",X"00",X"00",X"80",X"80",X"80",X"80",X"C0",X"E0",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"00",X"00",X"01",X"03",X"07",X"07",X"07",X"9F",X"80",X"80",X"C0",X"E0",X"F0",X"F0",X"FF",X"FF",
		X"9F",X"07",X"07",X"07",X"03",X"01",X"00",X"00",X"FF",X"FF",X"F0",X"F0",X"E0",X"C0",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"60",X"60",X"02",X"02",X"63",X"00",X"00",X"00",X"01",X"03",X"07",X"03",X"03",
		X"63",X"03",X"03",X"63",X"63",X"03",X"03",X"63",X"03",X"03",X"03",X"33",X"33",X"32",X"30",X"20",
		X"63",X"03",X"03",X"63",X"63",X"03",X"03",X"63",X"20",X"30",X"32",X"33",X"33",X"03",X"03",X"03",
		X"63",X"02",X"02",X"60",X"60",X"00",X"00",X"00",X"03",X"03",X"07",X"03",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"3F",X"00",X"00",X"00",X"00",X"F8",X"F9",X"6F",X"0F",
		X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"67",X"F9",X"F8",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"1F",X"1F",X"7F",X"FF",X"F0",X"FF",X"FF",X"E0",X"E0",X"E0",X"C0",X"80",X"80",X"F0",X"F0",
		X"FF",X"F0",X"FF",X"7F",X"1F",X"1F",X"1F",X"00",X"F0",X"80",X"80",X"C0",X"E0",X"E0",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"3F",X"00",X"00",X"00",X"00",X"F8",X"69",X"0F",X"6F",
		X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"0F",X"69",X"F9",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"1F",X"1F",X"7F",X"FF",X"F0",X"FF",X"FF",X"E0",X"E0",X"E0",X"C0",X"80",X"80",X"F0",X"F0",
		X"FF",X"F0",X"FF",X"7F",X"1F",X"1F",X"1F",X"00",X"F0",X"80",X"80",X"C0",X"E0",X"E0",X"E0",X"00",
		X"71",X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",X"1F",X"87",X"CF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"1F",X"1F",X"7F",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"79",X"F0",X"F0",X"F0",X"E0",X"80",
		X"00",X"18",X"B8",X"FC",X"FF",X"FF",X"FF",X"FF",X"1F",X"3F",X"7E",X"F8",X"F0",X"F0",X"C0",X"80",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"FF",X"FF",X"E0",X"E0",X"E0",X"E0",X"E0",X"F0",X"F0",X"F8",
		X"1F",X"1F",X"1F",X"3F",X"7F",X"FF",X"FF",X"E7",X"00",X"80",X"CB",X"CF",X"FF",X"FF",X"FF",X"FF",
		X"E3",X"C7",X"CF",X"1F",X"3C",X"78",X"F0",X"80",X"FF",X"FF",X"FF",X"FF",X"7F",X"7E",X"3C",X"10",
		X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"FC",X"FF",X"FF",X"FE",X"E0",X"E0",X"E0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"0F",X"06",X"F0",X"F0",X"F8",X"FC",X"FE",X"C7",X"83",X"00",
		X"3C",X"18",X"81",X"C3",X"C3",X"81",X"18",X"3C",X"82",X"C6",X"6E",X"3C",X"18",X"FE",X"FE",X"00",
		X"3C",X"18",X"BD",X"FF",X"FF",X"BD",X"18",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",X"00",X"02",X"02",X"FE",X"FE",X"42",X"02",X"00",X"00",
		X"62",X"F2",X"BA",X"9A",X"9E",X"CE",X"46",X"00",X"8C",X"DE",X"F2",X"B2",X"92",X"86",X"04",X"00",
		X"08",X"FE",X"FE",X"C8",X"68",X"38",X"18",X"00",X"1C",X"BE",X"A2",X"A2",X"A2",X"E6",X"E4",X"00",
		X"0C",X"9E",X"92",X"92",X"D2",X"7E",X"3C",X"00",X"C0",X"E0",X"B0",X"9E",X"8E",X"C0",X"C0",X"00",
		X"0C",X"6E",X"9A",X"9A",X"B2",X"F2",X"6C",X"00",X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",X"00",
		X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",X"44",X"C6",X"82",X"82",X"C6",X"7C",X"38",X"00",
		X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",X"82",X"92",X"92",X"92",X"FE",X"FE",X"00",X"00",
		X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",X"82",X"82",X"FE",X"FE",X"82",X"82",X"00",X"00",
		X"02",X"02",X"02",X"02",X"FE",X"FE",X"00",X"00",X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",
		X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",X"00",X"70",X"F8",X"88",X"88",X"88",X"FE",X"FE",X"00",
		X"72",X"F6",X"9E",X"8C",X"88",X"FE",X"FE",X"00",X"0C",X"5E",X"D2",X"92",X"92",X"F6",X"64",X"00",
		X"80",X"80",X"FE",X"FE",X"80",X"80",X"00",X"00",X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",
		X"C0",X"F0",X"1E",X"1E",X"F0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"FF",X"F0",X"F0",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FC",X"FF",X"07",X"07",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"80",X"80",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"F8",X"FC",X"3C",X"3C",X"FC",X"FC",X"FC",X"FC",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"1F",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"F0",X"F8",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"3F",X"7F",X"FE",X"FE",X"FE",X"FE",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"7F",X"FF",X"F0",X"F0",X"FF",X"7F",X"3F",
		X"FF",X"FF",X"FF",X"03",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C0",X"C0",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"80",X"80",X"80",X"00",X"00",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"FF",X"7F",X"3F",X"1F",X"00",X"00",X"1F",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",
		X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"F0",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"1F",X"3F",X"7F",X"FF",X"F0",
		X"FF",X"00",X"00",X"E0",X"E0",X"E0",X"E0",X"00",X"FF",X"00",X"00",X"7F",X"7F",X"7F",X"7F",X"00",
		X"00",X"00",X"00",X"80",X"C0",X"E0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"C3",X"E7",X"FF",X"3C",X"3C",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"07",X"07",X"07",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"81",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"07",X"07",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"F0",X"F0",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"3F",X"3C",X"3C",X"3F",X"1F",X"0F",X"07",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FF",X"0F",X"0F",X"FF",X"FE",X"FC",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"07",X"07",X"07",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"07",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"F8",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"3C",X"3C",X"3C",X"3C",X"3C",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",
		X"03",X"07",X"0F",X"1F",X"1F",X"3E",X"3C",X"3C",X"C0",X"E0",X"F0",X"F8",X"F8",X"7C",X"3C",X"3C",
		X"78",X"78",X"70",X"70",X"F0",X"E0",X"E0",X"C0",X"1E",X"1E",X"0E",X"0E",X"0F",X"07",X"07",X"03",
		X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"3F",X"00",X"00",X"00",X"00",X"F8",X"69",X"0F",X"0F",
		X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"0F",X"69",X"F8",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"1F",X"1F",X"7F",X"FF",X"F0",X"FF",X"FF",X"E0",X"E0",X"E0",X"C0",X"80",X"80",X"F0",X"F0",
		X"FF",X"F0",X"FF",X"7F",X"1F",X"1F",X"1F",X"00",X"F0",X"80",X"80",X"C0",X"E0",X"E0",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"C1",X"00",X"00",X"00",X"00",X"00",X"01",X"57",X"50",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F7",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"2F",X"00",X"7F",X"FF",X"FF",X"FF",X"01",X"00",X"C0",X"00",X"C0",X"80",X"80",X"F0",X"F0",
		X"FF",X"FF",X"FF",X"7F",X"00",X"2F",X"00",X"00",X"F0",X"80",X"80",X"C0",X"00",X"C0",X"00",X"00",
		X"7F",X"7F",X"3F",X"1F",X"0F",X"07",X"03",X"01",X"07",X"07",X"03",X"03",X"01",X"01",X"00",X"00",
		X"3F",X"3F",X"1F",X"1F",X"1F",X"0F",X"0F",X"0F",X"FF",X"7F",X"7F",X"7F",X"7F",X"7F",X"3F",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"3F",X"7F",X"7F",X"7F",X"7F",X"7F",X"FF",
		X"0F",X"0F",X"0F",X"1F",X"1F",X"1F",X"3F",X"3F",X"00",X"00",X"01",X"01",X"03",X"03",X"07",X"07",
		X"01",X"03",X"07",X"0F",X"1F",X"3F",X"7F",X"7F",X"C0",X"7A",X"38",X"0C",X"06",X"12",X"43",X"01",
		X"01",X"43",X"12",X"06",X"0C",X"38",X"7A",X"C0",X"18",X"9A",X"28",X"1C",X"49",X"18",X"08",X"18",
		X"9E",X"9E",X"92",X"82",X"C6",X"7C",X"38",X"00",X"FC",X"FE",X"02",X"02",X"02",X"FE",X"FC",X"00",
		X"80",X"90",X"90",X"90",X"FE",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
