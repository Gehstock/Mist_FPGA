library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity prog is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of prog is
	type rom is array(0 to  32767) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"F3",X"ED",X"56",X"31",X"00",X"F0",X"21",X"00",X"E0",X"11",X"01",X"E0",X"01",X"FF",X"0F",X"36",
		X"00",X"ED",X"B0",X"21",X"25",X"EB",X"22",X"03",X"EB",X"DB",X"04",X"CB",X"7F",X"CA",X"66",X"76",
		X"CD",X"8F",X"05",X"21",X"CC",X"05",X"11",X"06",X"EA",X"01",X"78",X"00",X"ED",X"B0",X"2A",X"3F",
		X"06",X"7D",X"6C",X"67",X"18",X"4C",X"C7",X"C7",X"08",X"D9",X"2A",X"03",X"EB",X"11",X"20",X"C0",
		X"01",X"C0",X"00",X"ED",X"B0",X"3A",X"02",X"E9",X"32",X"00",X"A0",X"3A",X"03",X"E9",X"32",X"00",
		X"B0",X"FD",X"E5",X"DD",X"E5",X"C3",X"8D",X"00",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"ED",X"45",X"63",X"AD",X"9C",X"52",X"72",X"CF",X"87",X"41",
		X"54",X"37",X"A7",X"43",X"91",X"51",X"A7",X"43",X"91",X"51",X"9F",X"B8",X"E5",X"D6",X"85",X"56",
		X"35",X"23",X"22",X"80",X"E9",X"21",X"17",X"E9",X"34",X"FB",X"C3",X"7E",X"48",X"3A",X"00",X"E0",
		X"A7",X"FA",X"F8",X"01",X"DB",X"04",X"CB",X"67",X"20",X"1D",X"21",X"05",X"E0",X"CB",X"7E",X"20",
		X"16",X"CB",X"46",X"DB",X"00",X"20",X"09",X"E6",X"02",X"20",X"0C",X"CB",X"C6",X"C3",X"F0",X"01",
		X"E6",X"01",X"C2",X"F0",X"01",X"CB",X"86",X"DB",X"04",X"CB",X"5F",X"20",X"10",X"21",X"04",X"E9",
		X"CB",X"4E",X"28",X"09",X"21",X"0E",X"E8",X"35",X"F2",X"F0",X"01",X"36",X"08",X"3A",X"00",X"E0",
		X"FE",X"06",X"3E",X"47",X"28",X"02",X"ED",X"5F",X"21",X"10",X"E0",X"86",X"77",X"23",X"86",X"77",
		X"21",X"14",X"E0",X"34",X"7E",X"E6",X"03",X"16",X"00",X"5F",X"3A",X"00",X"E0",X"21",X"7E",X"00",
		X"FE",X"06",X"28",X"13",X"21",X"6E",X"00",X"3A",X"80",X"E0",X"E6",X"38",X"FE",X"20",X"38",X"02",
		X"3E",X"18",X"0F",X"4F",X"06",X"00",X"09",X"19",X"7E",X"21",X"15",X"E0",X"86",X"77",X"23",X"86",
		X"77",X"23",X"86",X"77",X"CD",X"05",X"0D",X"CD",X"48",X"0D",X"CD",X"2F",X"48",X"CD",X"E5",X"0D",
		X"3A",X"01",X"E0",X"A7",X"20",X"07",X"3A",X"13",X"E9",X"A7",X"C2",X"17",X"02",X"CD",X"F8",X"03",
		X"3A",X"00",X"E0",X"FE",X"0B",X"D2",X"DD",X"01",X"3E",X"18",X"32",X"00",X"EB",X"21",X"25",X"EB",
		X"22",X"03",X"EB",X"22",X"01",X"EB",X"3A",X"00",X"E0",X"87",X"5F",X"16",X"00",X"21",X"56",X"01",
		X"19",X"5E",X"23",X"56",X"EB",X"E9",X"C4",X"01",X"C4",X"01",X"BE",X"01",X"68",X"01",X"68",X"01",
		X"B4",X"01",X"68",X"01",X"B9",X"01",X"BE",X"01",X"CD",X"3F",X"41",X"CD",X"2C",X"40",X"3A",X"80",
		X"E0",X"E6",X"07",X"FE",X"04",X"28",X"08",X"CD",X"E5",X"40",X"CD",X"B3",X"1C",X"18",X"06",X"CD",
		X"B3",X"1C",X"CD",X"E5",X"40",X"CD",X"B6",X"47",X"3A",X"00",X"E1",X"A7",X"28",X"0E",X"FE",X"0A",
		X"38",X"05",X"CD",X"DE",X"37",X"18",X"08",X"CD",X"95",X"35",X"18",X"03",X"CD",X"AC",X"12",X"CD",
		X"C7",X"2F",X"3A",X"3F",X"E3",X"A7",X"C4",X"C1",X"2E",X"CD",X"C0",X"39",X"CD",X"72",X"2D",X"CD",
		X"06",X"2F",X"18",X"10",X"CD",X"24",X"4D",X"18",X"0B",X"CD",X"36",X"54",X"18",X"06",X"CD",X"00",
		X"40",X"CD",X"E5",X"40",X"3A",X"00",X"EB",X"A7",X"28",X"13",X"47",X"FD",X"2A",X"01",X"EB",X"AF",
		X"11",X"08",X"00",X"FD",X"77",X"04",X"FD",X"77",X"05",X"FD",X"19",X"10",X"F6",X"3A",X"00",X"E0",
		X"FE",X"06",X"3E",X"37",X"28",X"02",X"ED",X"5F",X"21",X"12",X"E0",X"86",X"77",X"23",X"86",X"77",
		X"DD",X"E1",X"FD",X"E1",X"D9",X"08",X"FB",X"C9",X"F5",X"3E",X"18",X"32",X"00",X"EB",X"21",X"25",
		X"EB",X"22",X"03",X"EB",X"22",X"01",X"EB",X"F1",X"3C",X"C4",X"AE",X"7A",X"CD",X"F8",X"03",X"CD",
		X"05",X"0D",X"CD",X"E5",X"0D",X"18",X"AD",X"31",X"00",X"F0",X"3E",X"01",X"32",X"01",X"E0",X"AF",
		X"32",X"00",X"E0",X"FB",X"CD",X"78",X"51",X"3E",X"FF",X"32",X"06",X"E0",X"21",X"80",X"E0",X"11",
		X"81",X"E0",X"01",X"1F",X"00",X"36",X"00",X"ED",X"B0",X"DB",X"03",X"E6",X"01",X"20",X"08",X"3E",
		X"08",X"32",X"80",X"E0",X"32",X"90",X"E0",X"CD",X"6F",X"05",X"32",X"84",X"E0",X"32",X"94",X"E0",
		X"21",X"05",X"E0",X"CB",X"BE",X"AF",X"32",X"00",X"E0",X"DB",X"04",X"E6",X"02",X"21",X"10",X"E9",
		X"28",X"0B",X"3A",X"02",X"E0",X"E6",X"01",X"28",X"04",X"CB",X"C6",X"18",X"02",X"CB",X"86",X"21",
		X"85",X"E0",X"CB",X"4E",X"20",X"0F",X"CB",X"CE",X"CD",X"0D",X"52",X"3E",X"E1",X"CD",X"0F",X"57",
		X"3E",X"70",X"CD",X"0F",X"57",X"CD",X"57",X"11",X"AF",X"32",X"07",X"E0",X"32",X"08",X"E0",X"CD",
		X"49",X"04",X"3E",X"04",X"32",X"00",X"E0",X"3E",X"24",X"CD",X"FE",X"0D",X"DB",X"04",X"CB",X"67",
		X"28",X"0C",X"CB",X"6F",X"20",X"08",X"21",X"04",X"E9",X"CB",X"46",X"C2",X"9C",X"03",X"3A",X"00",
		X"E0",X"FE",X"0B",X"CA",X"3A",X"03",X"FE",X"0C",X"CA",X"C0",X"02",X"CD",X"B8",X"0F",X"18",X"DC",
		X"3E",X"00",X"CD",X"FE",X"0D",X"3E",X"22",X"CD",X"FE",X"0D",X"3E",X"E1",X"CD",X"82",X"05",X"3E",
		X"38",X"CD",X"82",X"05",X"3E",X"01",X"CD",X"82",X"05",X"21",X"09",X"E7",X"7E",X"A7",X"FA",X"EA",
		X"02",X"35",X"CD",X"97",X"2F",X"CD",X"5F",X"05",X"18",X"EA",X"11",X"00",X"00",X"D5",X"3E",X"03",
		X"CD",X"82",X"05",X"D1",X"2A",X"03",X"E0",X"7D",X"B4",X"28",X"22",X"7B",X"C6",X"01",X"27",X"5F",
		X"ED",X"52",X"19",X"30",X"02",X"5D",X"54",X"7D",X"93",X"27",X"6F",X"7C",X"9A",X"27",X"67",X"22",
		X"03",X"E0",X"D5",X"CD",X"9A",X"2F",X"3E",X"16",X"CD",X"FE",X"0D",X"18",X"D1",X"3E",X"38",X"CD",
		X"82",X"05",X"3A",X"80",X"E0",X"E6",X"01",X"C4",X"C2",X"53",X"3A",X"80",X"E0",X"E6",X"07",X"FE",
		X"04",X"CC",X"E9",X"4F",X"CD",X"32",X"04",X"CD",X"50",X"02",X"3E",X"2D",X"CD",X"0F",X"57",X"2A",
		X"03",X"E0",X"7D",X"B4",X"CC",X"B5",X"56",X"21",X"84",X"E0",X"35",X"28",X"10",X"3A",X"07",X"E0",
		X"A7",X"28",X"0D",X"CD",X"FE",X"0D",X"3E",X"A9",X"CD",X"0F",X"57",X"18",X"03",X"CD",X"F4",X"54",
		X"21",X"02",X"E0",X"CB",X"4E",X"28",X"1B",X"3A",X"94",X"E0",X"A7",X"28",X"15",X"7E",X"EE",X"01",
		X"77",X"06",X"10",X"21",X"80",X"E0",X"11",X"90",X"E0",X"4E",X"1A",X"EB",X"71",X"12",X"23",X"13",
		X"10",X"F7",X"3A",X"84",X"E0",X"A7",X"C2",X"50",X"02",X"21",X"10",X"E9",X"CB",X"86",X"AF",X"32",
		X"06",X"E0",X"3A",X"13",X"E9",X"A7",X"C2",X"17",X"02",X"C3",X"7E",X"48",X"21",X"05",X"E0",X"CB",
		X"FE",X"3E",X"00",X"CD",X"FE",X"0D",X"AF",X"32",X"00",X"E0",X"CD",X"57",X"11",X"21",X"00",X"00",
		X"22",X"02",X"E9",X"CD",X"0D",X"57",X"21",X"5B",X"59",X"CD",X"1C",X"11",X"0E",X"14",X"11",X"A7",
		X"D3",X"3A",X"80",X"E0",X"E6",X"F8",X"0F",X"0F",X"0F",X"CD",X"5B",X"05",X"11",X"27",X"D4",X"CD",
		X"56",X"05",X"3A",X"06",X"E9",X"E6",X"A0",X"20",X"F9",X"21",X"04",X"E9",X"CB",X"4E",X"C2",X"50",
		X"02",X"21",X"06",X"E9",X"CB",X"7E",X"20",X"06",X"CB",X"6E",X"20",X"07",X"18",X"EB",X"CD",X"1B",
		X"04",X"18",X"C9",X"CD",X"32",X"04",X"18",X"C4",X"21",X"80",X"E8",X"35",X"23",X"7E",X"A7",X"28",
		X"01",X"35",X"23",X"7E",X"A7",X"28",X"01",X"35",X"23",X"7E",X"A7",X"28",X"01",X"35",X"23",X"7E",
		X"A7",X"28",X"01",X"35",X"23",X"7E",X"A7",X"28",X"01",X"35",X"C9",X"21",X"80",X"E0",X"35",X"7E",
		X"E6",X"07",X"FE",X"07",X"C0",X"7E",X"E6",X"F8",X"FE",X"F8",X"20",X"02",X"3E",X"28",X"F6",X"04",
		X"77",X"C9",X"21",X"80",X"E0",X"34",X"7E",X"E6",X"07",X"FE",X"05",X"C0",X"7E",X"E6",X"F8",X"C6",
		X"08",X"FE",X"30",X"20",X"02",X"3E",X"28",X"77",X"C9",X"32",X"1C",X"E8",X"3E",X"01",X"32",X"00",
		X"E0",X"CD",X"44",X"06",X"3A",X"80",X"E0",X"E6",X"01",X"21",X"21",X"00",X"20",X"03",X"21",X"E0",
		X"BF",X"E5",X"22",X"17",X"E8",X"CD",X"9B",X"0E",X"AF",X"32",X"15",X"E9",X"CD",X"56",X"57",X"3A",
		X"1C",X"E8",X"A7",X"CC",X"E5",X"04",X"3E",X"02",X"32",X"00",X"E0",X"3E",X"27",X"CD",X"0F",X"57",
		X"21",X"07",X"00",X"22",X"17",X"E8",X"21",X"15",X"E9",X"34",X"21",X"A1",X"5A",X"CD",X"BF",X"04",
		X"3E",X"0B",X"CD",X"0F",X"57",X"21",X"15",X"E9",X"34",X"21",X"F0",X"5A",X"CD",X"BF",X"04",X"3A",
		X"1C",X"E8",X"A7",X"21",X"3F",X"05",X"CC",X"1C",X"11",X"3E",X"54",X"CD",X"0F",X"57",X"E1",X"22",
		X"17",X"E8",X"CD",X"56",X"57",X"21",X"00",X"00",X"22",X"14",X"E0",X"22",X"16",X"E0",X"C9",X"3A",
		X"80",X"E0",X"E6",X"07",X"C8",X"E6",X"01",X"CA",X"1C",X"11",X"CD",X"56",X"57",X"3A",X"15",X"E9",
		X"FE",X"02",X"C0",X"21",X"D9",X"04",X"C3",X"1C",X"11",X"FD",X"67",X"D6",X"FE",X"92",X"81",X"7F",
		X"FD",X"A7",X"D6",X"83",X"FF",X"21",X"FD",X"04",X"CD",X"1C",X"11",X"3A",X"02",X"E0",X"E6",X"01",
		X"3C",X"CD",X"08",X"11",X"CD",X"1C",X"11",X"CD",X"56",X"05",X"C3",X"1C",X"11",X"FD",X"67",X"D3",
		X"FE",X"DB",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"FD",X"A7",X"D3",X"20",X"FF",X"2D",X"50",X"4C",X"41",X"59",X"45",X"52",
		X"20",X"FF",X"2D",X"46",X"4C",X"4F",X"4F",X"52",X"20",X"FD",X"E7",X"D3",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"FF",X"FE",
		X"DB",X"FD",X"2C",X"D4",X"20",X"52",X"45",X"41",X"44",X"59",X"20",X"FD",X"6C",X"D4",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"FF",X"3A",X"80",X"E0",X"E6",X"07",X"3C",X"C3",X"08",X"11",X"3A",
		X"83",X"E8",X"A7",X"C0",X"3E",X"03",X"32",X"83",X"E8",X"3E",X"16",X"CD",X"FE",X"0D",X"C9",X"DB",
		X"03",X"2F",X"E6",X"0C",X"0F",X"0F",X"C6",X"02",X"FE",X"04",X"D0",X"3C",X"FE",X"03",X"C8",X"3E",
		X"02",X"C9",X"32",X"82",X"E8",X"CD",X"E3",X"0F",X"3A",X"82",X"E8",X"A7",X"20",X"F7",X"C9",X"DB",
		X"03",X"2F",X"1F",X"1F",X"1F",X"1F",X"47",X"21",X"0A",X"E9",X"DB",X"04",X"CB",X"57",X"20",X"11",
		X"78",X"3C",X"E6",X"03",X"77",X"23",X"78",X"1F",X"1F",X"E6",X"03",X"FE",X"02",X"DE",X"F5",X"77",
		X"C9",X"78",X"3C",X"E6",X"0F",X"FE",X"07",X"38",X"0A",X"FE",X"09",X"38",X"04",X"FE",X"0E",X"38",
		X"02",X"3E",X"01",X"CB",X"5F",X"28",X"01",X"3C",X"77",X"23",X"77",X"C9",X"00",X"14",X"95",X"54",
		X"41",X"2E",X"00",X"15",X"38",X"41",X"41",X"41",X"00",X"15",X"72",X"4E",X"4E",X"49",X"00",X"16",
		X"52",X"41",X"41",X"41",X"00",X"18",X"21",X"49",X"4B",X"4F",X"00",X"19",X"85",X"41",X"49",X"2E",
		X"00",X"20",X"07",X"41",X"4E",X"4F",X"00",X"21",X"01",X"4D",X"2E",X"4B",X"00",X"25",X"51",X"49",
		X"49",X"41",X"00",X"25",X"70",X"48",X"41",X"54",X"00",X"26",X"35",X"41",X"2E",X"54",X"00",X"28",
		X"11",X"59",X"45",X"2E",X"00",X"30",X"21",X"53",X"41",X"49",X"00",X"35",X"50",X"49",X"48",X"4D",
		X"00",X"38",X"10",X"41",X"4E",X"49",X"00",X"39",X"18",X"54",X"53",X"49",X"00",X"39",X"75",X"42",
		X"41",X"48",X"00",X"40",X"10",X"54",X"2E",X"4B",X"00",X"43",X"15",X"53",X"55",X"49",X"00",X"48",
		X"52",X"4E",X"2E",X"41",X"21",X"80",X"00",X"22",X"02",X"E9",X"21",X"25",X"EB",X"11",X"26",X"EB",
		X"01",X"BF",X"00",X"36",X"00",X"ED",X"B0",X"CD",X"4D",X"07",X"CD",X"BE",X"06",X"21",X"80",X"E3",
		X"11",X"81",X"E3",X"01",X"31",X"01",X"36",X"00",X"ED",X"B0",X"CD",X"66",X"08",X"21",X"8A",X"08",
		X"09",X"7E",X"32",X"00",X"E1",X"A7",X"28",X"11",X"21",X"B0",X"08",X"11",X"60",X"E3",X"01",X"18",
		X"00",X"CD",X"B2",X"06",X"3E",X"01",X"32",X"80",X"E3",X"21",X"20",X"E5",X"11",X"21",X"E5",X"01",
		X"43",X"01",X"36",X"00",X"ED",X"B0",X"CD",X"66",X"08",X"21",X"9E",X"08",X"09",X"7E",X"A7",X"C8",
		X"32",X"00",X"E1",X"21",X"20",X"09",X"11",X"00",X"E5",X"01",X"11",X"00",X"CD",X"B2",X"06",X"C3",
		X"53",X"3D",X"87",X"C5",X"4F",X"09",X"C1",X"7E",X"23",X"66",X"6F",X"ED",X"B0",X"C9",X"21",X"00",
		X"E7",X"11",X"01",X"E7",X"01",X"23",X"00",X"36",X"00",X"ED",X"B0",X"3A",X"80",X"E0",X"E6",X"07",
		X"87",X"4F",X"21",X"80",X"08",X"09",X"7E",X"23",X"66",X"6F",X"22",X"03",X"E0",X"3E",X"3F",X"32",
		X"09",X"E7",X"21",X"00",X"50",X"22",X"10",X"E7",X"3A",X"80",X"E0",X"E6",X"01",X"32",X"01",X"E1",
		X"28",X"2B",X"21",X"00",X"E7",X"36",X"20",X"23",X"36",X"40",X"21",X"40",X"CE",X"22",X"02",X"E1",
		X"21",X"00",X"09",X"22",X"12",X"E7",X"21",X"00",X"10",X"22",X"07",X"E7",X"21",X"00",X"CD",X"22",
		X"06",X"E1",X"21",X"C0",X"02",X"22",X"04",X"E1",X"3E",X"01",X"C3",X"49",X"07",X"3A",X"80",X"E0",
		X"E6",X"07",X"21",X"E0",X"10",X"FE",X"04",X"20",X"03",X"21",X"00",X"10",X"22",X"02",X"E1",X"21",
		X"60",X"D5",X"22",X"12",X"E7",X"21",X"00",X"D0",X"22",X"07",X"E7",X"21",X"40",X"DC",X"22",X"06",
		X"E1",X"21",X"C0",X"11",X"22",X"04",X"E1",X"3E",X"DF",X"32",X"14",X"E7",X"C9",X"21",X"00",X"E2",
		X"11",X"01",X"E2",X"01",X"52",X"01",X"36",X"00",X"ED",X"B0",X"3A",X"80",X"E0",X"E6",X"07",X"FE",
		X"04",X"20",X"2E",X"21",X"00",X"06",X"22",X"42",X"E3",X"21",X"80",X"07",X"22",X"4E",X"E3",X"21",
		X"00",X"50",X"22",X"44",X"E3",X"22",X"50",X"E3",X"3E",X"04",X"32",X"46",X"E3",X"3E",X"07",X"32",
		X"52",X"E3",X"3E",X"40",X"32",X"4C",X"E3",X"3E",X"50",X"32",X"40",X"E3",X"3E",X"05",X"32",X"47",
		X"E3",X"DD",X"21",X"D8",X"E2",X"DD",X"36",X"0A",X"3F",X"DD",X"36",X"07",X"07",X"21",X"00",X"50",
		X"22",X"DC",X"E2",X"3A",X"80",X"E0",X"E6",X"01",X"21",X"00",X"15",X"11",X"00",X"31",X"28",X"06",
		X"21",X"00",X"CC",X"11",X"00",X"B0",X"22",X"DA",X"E2",X"ED",X"53",X"D3",X"E2",X"CD",X"66",X"08",
		X"C5",X"CB",X"21",X"C5",X"C5",X"21",X"B0",X"09",X"09",X"7E",X"23",X"66",X"6F",X"11",X"9C",X"E1",
		X"01",X"1D",X"00",X"ED",X"B0",X"21",X"80",X"09",X"C1",X"09",X"7E",X"23",X"66",X"6F",X"B4",X"28",
		X"05",X"01",X"08",X"00",X"ED",X"B0",X"C1",X"21",X"E0",X"0B",X"09",X"11",X"96",X"E1",X"ED",X"A0",
		X"ED",X"A0",X"AF",X"12",X"C1",X"21",X"18",X"0B",X"09",X"7E",X"32",X"C1",X"E1",X"21",X"08",X"0C",
		X"09",X"7E",X"32",X"99",X"E1",X"32",X"9A",X"E1",X"32",X"9B",X"E1",X"FD",X"21",X"00",X"00",X"21",
		X"2E",X"0C",X"09",X"09",X"5E",X"23",X"56",X"FD",X"19",X"DD",X"21",X"0A",X"E1",X"11",X"1C",X"0C",
		X"06",X"23",X"CD",X"45",X"08",X"FD",X"23",X"10",X"F9",X"21",X"FF",X"E1",X"22",X"08",X"E1",X"CD",
		X"66",X"08",X"50",X"59",X"21",X"2C",X"0B",X"19",X"EB",X"29",X"29",X"29",X"19",X"11",X"F0",X"E1",
		X"0E",X"09",X"ED",X"B0",X"C9",X"FD",X"7E",X"00",X"F5",X"0F",X"0F",X"0F",X"0F",X"CD",X"51",X"08",
		X"F1",X"E6",X"0F",X"87",X"26",X"00",X"6F",X"19",X"7E",X"DD",X"77",X"00",X"23",X"7E",X"DD",X"77",
		X"01",X"DD",X"23",X"DD",X"23",X"C9",X"3A",X"80",X"E0",X"6F",X"E6",X"07",X"67",X"7D",X"E6",X"38",
		X"FE",X"20",X"38",X"02",X"3E",X"18",X"0F",X"6F",X"0F",X"0F",X"85",X"84",X"4F",X"06",X"00",X"C9",
		X"00",X"20",X"00",X"20",X"00",X"20",X"00",X"20",X"00",X"20",X"00",X"01",X"00",X"02",X"00",X"00",
		X"03",X"00",X"02",X"00",X"00",X"04",X"00",X"02",X"00",X"00",X"05",X"00",X"02",X"00",X"00",X"00",
		X"00",X"0A",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",
		X"0D",X"00",X"BC",X"08",X"1C",X"09",X"D4",X"08",X"EC",X"08",X"04",X"09",X"00",X"00",X"70",X"00",
		X"0D",X"54",X"A8",X"43",X"5A",X"70",X"66",X"CC",X"00",X"00",X"36",X"00",X"16",X"A9",X"B6",X"01",
		X"4B",X"01",X"7C",X"00",X"00",X"00",X"70",X"00",X"0D",X"54",X"A8",X"2D",X"43",X"5A",X"66",X"CC",
		X"00",X"00",X"36",X"00",X"16",X"A9",X"B6",X"01",X"4B",X"01",X"7C",X"00",X"00",X"00",X"70",X"00",
		X"0D",X"54",X"A8",X"1C",X"38",X"43",X"66",X"CC",X"00",X"00",X"36",X"00",X"16",X"A9",X"B6",X"01",
		X"4B",X"01",X"7C",X"00",X"00",X"00",X"70",X"00",X"0D",X"54",X"A8",X"1C",X"2D",X"38",X"66",X"CC",
		X"00",X"00",X"36",X"00",X"16",X"A9",X"B6",X"01",X"4B",X"01",X"7C",X"00",X"00",X"00",X"00",X"36",
		X"00",X"30",X"49",X"00",X"00",X"00",X"61",X"00",X"A4",X"00",X"36",X"00",X"16",X"00",X"52",X"00",
		X"49",X"00",X"2D",X"00",X"3C",X"09",X"4D",X"09",X"5E",X"09",X"6F",X"09",X"20",X"00",X"32",X"00",
		X"28",X"00",X"33",X"00",X"23",X"00",X"6B",X"07",X"7F",X"3F",X"3F",X"38",X"70",X"32",X"00",X"3B",
		X"00",X"3F",X"00",X"50",X"00",X"38",X"00",X"6B",X"07",X"B2",X"3F",X"66",X"38",X"70",X"32",X"00",
		X"3B",X"00",X"3F",X"00",X"50",X"00",X"38",X"00",X"38",X"04",X"7F",X"66",X"66",X"1C",X"38",X"3B",
		X"00",X"44",X"00",X"4A",X"00",X"5F",X"00",X"44",X"00",X"38",X"04",X"B2",X"66",X"7F",X"1C",X"38",
		X"00",X"00",X"A8",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A8",X"09",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"A8",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A8",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"B3",X"FF",X"07",X"00",X"2E",X"00",X"D7",X"00",
		X"D8",X"09",X"E1",X"09",X"EF",X"09",X"FD",X"09",X"0B",X"0A",X"28",X"0A",X"31",X"0A",X"3F",X"0A",
		X"4D",X"0A",X"5B",X"0A",X"78",X"0A",X"81",X"0A",X"8F",X"0A",X"9D",X"0A",X"AB",X"0A",X"C8",X"0A",
		X"D1",X"0A",X"DF",X"0A",X"ED",X"0A",X"FB",X"0A",X"99",X"E5",X"66",X"99",X"54",X"A8",X"21",X"16",
		X"0B",X"66",X"7F",X"CC",X"03",X"54",X"A8",X"2D",X"5A",X"70",X"54",X"A8",X"1C",X"2D",X"38",X"CC",
		X"E5",X"A8",X"FC",X"54",X"A8",X"2D",X"5A",X"70",X"00",X"00",X"00",X"00",X"16",X"54",X"A8",X"99",
		X"B7",X"7F",X"FC",X"70",X"A9",X"A9",X"54",X"54",X"38",X"70",X"A9",X"66",X"CC",X"54",X"A8",X"54",
		X"A8",X"0B",X"16",X"21",X"54",X"A8",X"05",X"08",X"0B",X"03",X"80",X"00",X"99",X"7F",X"66",X"7F",
		X"CC",X"66",X"4C",X"7F",X"99",X"7F",X"7F",X"4C",X"7F",X"BF",X"33",X"66",X"54",X"A8",X"1F",X"15",
		X"0B",X"4C",X"66",X"B2",X"03",X"54",X"A8",X"2D",X"5A",X"70",X"54",X"A8",X"1C",X"2D",X"38",X"B2",
		X"E5",X"A8",X"FC",X"54",X"A8",X"21",X"38",X"5A",X"00",X"00",X"00",X"00",X"10",X"54",X"A8",X"7F",
		X"B2",X"7F",X"FC",X"70",X"A9",X"A9",X"54",X"54",X"1C",X"38",X"70",X"66",X"CC",X"54",X"A8",X"54",
		X"A8",X"0B",X"16",X"21",X"54",X"A8",X"05",X"08",X"0B",X"03",X"80",X"00",X"99",X"7F",X"7F",X"7F",
		X"CC",X"7F",X"66",X"7F",X"99",X"7F",X"7F",X"7F",X"4C",X"B2",X"33",X"66",X"54",X"A8",X"1C",X"13",
		X"0B",X"33",X"7F",X"CC",X"03",X"54",X"A8",X"2D",X"5A",X"70",X"54",X"A8",X"10",X"1C",X"2D",X"99",
		X"E5",X"7F",X"FC",X"54",X"A8",X"16",X"2D",X"43",X"00",X"00",X"00",X"00",X"0B",X"54",X"A8",X"66",
		X"B2",X"7F",X"FC",X"70",X"A9",X"A9",X"54",X"54",X"1C",X"38",X"70",X"66",X"CC",X"54",X"A8",X"54",
		X"A8",X"0B",X"16",X"21",X"54",X"A8",X"05",X"08",X"0B",X"03",X"80",X"00",X"CC",X"CC",X"7F",X"CC",
		X"CC",X"7F",X"4C",X"7F",X"CC",X"CC",X"CC",X"4C",X"4C",X"99",X"33",X"66",X"54",X"A8",X"19",X"13",
		X"0B",X"19",X"7F",X"E5",X"03",X"54",X"A8",X"2D",X"5A",X"70",X"54",X"A8",X"10",X"1C",X"2D",X"7F",
		X"CC",X"54",X"FC",X"54",X"A8",X"16",X"2D",X"43",X"00",X"00",X"00",X"00",X"0B",X"54",X"A8",X"54",
		X"A8",X"7F",X"FC",X"70",X"A9",X"A9",X"54",X"54",X"1C",X"1C",X"70",X"66",X"CC",X"54",X"A8",X"54",
		X"A8",X"0B",X"16",X"21",X"54",X"A8",X"05",X"08",X"0B",X"03",X"80",X"00",X"E5",X"CC",X"7F",X"CC",
		X"E5",X"99",X"7F",X"7F",X"E5",X"CC",X"CC",X"7F",X"00",X"00",X"26",X"33",X"4C",X"00",X"19",X"26",
		X"33",X"4C",X"00",X"19",X"33",X"4C",X"66",X"00",X"19",X"4C",X"66",X"7F",X"04",X"3F",X"5A",X"B4",
		X"E1",X"1A",X"01",X"49",X"00",X"04",X"3F",X"5A",X"B4",X"E1",X"1A",X"01",X"49",X"00",X"04",X"55",
		X"5A",X"B4",X"E1",X"1A",X"01",X"49",X"00",X"04",X"55",X"5A",X"B4",X"E1",X"1A",X"01",X"49",X"00",
		X"04",X"66",X"5A",X"B4",X"E1",X"1A",X"01",X"49",X"00",X"04",X"66",X"5A",X"B4",X"E1",X"E1",X"00",
		X"52",X"00",X"04",X"66",X"5A",X"B4",X"E1",X"E1",X"00",X"52",X"00",X"04",X"66",X"5A",X"B4",X"E1",
		X"E1",X"00",X"52",X"00",X"04",X"66",X"5A",X"B4",X"E1",X"E1",X"00",X"52",X"00",X"04",X"66",X"5A",
		X"B4",X"E1",X"E1",X"00",X"52",X"00",X"04",X"7F",X"5A",X"B4",X"E1",X"A9",X"00",X"5B",X"00",X"04",
		X"7F",X"5A",X"B4",X"E1",X"A9",X"00",X"5B",X"00",X"04",X"7F",X"5A",X"B4",X"E1",X"A9",X"00",X"5B",
		X"00",X"04",X"7F",X"5A",X"B4",X"E1",X"A9",X"00",X"5B",X"00",X"04",X"7F",X"5A",X"B4",X"E1",X"A9",
		X"00",X"5B",X"00",X"04",X"7F",X"5A",X"B4",X"E1",X"A9",X"00",X"5B",X"00",X"04",X"7F",X"5A",X"B4",
		X"E1",X"A9",X"00",X"5B",X"00",X"04",X"7F",X"5A",X"B4",X"E1",X"A9",X"00",X"5B",X"00",X"04",X"7F",
		X"5A",X"B4",X"E1",X"A9",X"00",X"5B",X"00",X"04",X"7F",X"5A",X"B4",X"E1",X"A9",X"00",X"5B",X"00",
		X"03",X"03",X"04",X"03",X"05",X"03",X"05",X"03",X"05",X"03",X"05",X"03",X"05",X"03",X"05",X"03",
		X"05",X"03",X"05",X"03",X"05",X"03",X"05",X"03",X"05",X"03",X"05",X"04",X"05",X"04",X"05",X"03",
		X"05",X"03",X"05",X"03",X"05",X"05",X"05",X"05",X"0D",X"0C",X"0B",X"0A",X"09",X"0B",X"0A",X"09",
		X"08",X"08",X"0A",X"09",X"09",X"08",X"07",X"09",X"08",X"08",X"07",X"07",X"80",X"00",X"00",X"1C",
		X"00",X"38",X"00",X"70",X"00",X"E1",X"04",X"1C",X"04",X"38",X"04",X"70",X"04",X"E1",X"56",X"0C",
		X"79",X"0C",X"9C",X"0C",X"BF",X"0C",X"E2",X"0C",X"56",X"0C",X"79",X"0C",X"9C",X"0C",X"BF",X"0C",
		X"E2",X"0C",X"56",X"0C",X"79",X"0C",X"9C",X"0C",X"BF",X"0C",X"E2",X"0C",X"56",X"0C",X"79",X"0C",
		X"9C",X"0C",X"BF",X"0C",X"E2",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"00",X"04",X"42",X"43",X"43",X"42",X"44",X"23",X"34",X"43",X"43",X"43",X"33",X"34",
		X"34",X"43",X"43",X"33",X"43",X"34",X"43",X"30",X"00",X"00",X"61",X"03",X"22",X"00",X"30",X"32",
		X"40",X"27",X"23",X"00",X"23",X"12",X"73",X"32",X"03",X"27",X"20",X"73",X"32",X"71",X"03",X"02",
		X"52",X"32",X"75",X"21",X"63",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"34",X"45",X"13",X"17",X"17",X"73",X"21",
		X"37",X"27",X"32",X"63",X"37",X"34",X"32",X"43",X"22",X"32",X"42",X"23",X"23",X"20",X"00",X"01",
		X"23",X"03",X"25",X"00",X"70",X"16",X"31",X"06",X"31",X"00",X"25",X"13",X"54",X"23",X"00",X"07",
		X"12",X"63",X"61",X"61",X"27",X"12",X"56",X"72",X"16",X"21",X"52",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"03",
		X"31",X"21",X"23",X"17",X"63",X"61",X"32",X"25",X"72",X"53",X"27",X"32",X"15",X"31",X"06",X"21",
		X"73",X"16",X"13",X"50",X"00",X"3A",X"10",X"E9",X"E6",X"01",X"DB",X"01",X"28",X"02",X"DB",X"02",
		X"2A",X"06",X"E9",X"CD",X"3B",X"0D",X"22",X"06",X"E9",X"21",X"08",X"E9",X"17",X"CB",X"16",X"17",
		X"17",X"CB",X"16",X"17",X"17",X"CB",X"16",X"DB",X"00",X"E6",X"0F",X"47",X"DB",X"02",X"E6",X"10",
		X"B0",X"2A",X"04",X"E9",X"CD",X"3B",X"0D",X"22",X"04",X"E9",X"C9",X"2F",X"47",X"AC",X"4F",X"A5",
		X"6F",X"79",X"2F",X"A4",X"B5",X"6F",X"60",X"C9",X"0F",X"0F",X"0F",X"47",X"3A",X"11",X"E9",X"17",
		X"4F",X"E6",X"49",X"FE",X"49",X"20",X"0A",X"21",X"14",X"E9",X"34",X"7E",X"E6",X"0F",X"CC",X"D6",
		X"0D",X"21",X"0C",X"E9",X"11",X"0A",X"E9",X"CD",X"B1",X"0D",X"21",X"0E",X"E9",X"13",X"CD",X"B1",
		X"0D",X"21",X"11",X"E9",X"71",X"2B",X"4E",X"2B",X"06",X"04",X"CD",X"A2",X"0D",X"21",X"0D",X"E9",
		X"06",X"02",X"CD",X"A2",X"0D",X"79",X"32",X"10",X"E9",X"D3",X"01",X"DB",X"04",X"2F",X"A9",X"E6",
		X"01",X"28",X"01",X"3C",X"32",X"16",X"E9",X"3A",X"0A",X"E9",X"A7",X"C0",X"3E",X"02",X"32",X"13",
		X"E9",X"C9",X"35",X"F0",X"36",X"0C",X"2B",X"7E",X"A7",X"C8",X"78",X"A9",X"4F",X"A0",X"C0",X"35",
		X"C9",X"CB",X"08",X"CB",X"11",X"79",X"E6",X"49",X"FE",X"01",X"C0",X"34",X"3A",X"06",X"E0",X"A7",
		X"3E",X"01",X"CC",X"FE",X"0D",X"1A",X"FE",X"01",X"28",X"10",X"FE",X"08",X"30",X"0A",X"21",X"12",
		X"E9",X"34",X"BE",X"C0",X"36",X"00",X"3E",X"09",X"D6",X"08",X"21",X"13",X"E9",X"86",X"27",X"30",
		X"02",X"3E",X"99",X"77",X"C9",X"21",X"17",X"E9",X"7E",X"A7",X"C8",X"35",X"23",X"7E",X"D3",X"00",
		X"F6",X"80",X"D3",X"00",X"23",X"11",X"18",X"E9",X"01",X"0F",X"00",X"ED",X"B0",X"C9",X"E5",X"D5",
		X"57",X"CB",X"7A",X"28",X"08",X"3A",X"06",X"E0",X"A7",X"28",X"12",X"CB",X"BA",X"21",X"17",X"E9",
		X"7E",X"FE",X"10",X"30",X"08",X"34",X"23",X"5F",X"7A",X"16",X"00",X"19",X"77",X"D1",X"E1",X"C9",
		X"E5",X"4F",X"3A",X"00",X"EB",X"47",X"FD",X"2A",X"01",X"EB",X"CB",X"71",X"21",X"20",X"00",X"20",
		X"03",X"21",X"D0",X"FF",X"19",X"22",X"05",X"E8",X"E1",X"05",X"04",X"C8",X"7E",X"3C",X"28",X"52",
		X"3A",X"05",X"E8",X"CB",X"71",X"20",X"0B",X"86",X"FD",X"77",X"06",X"3A",X"06",X"E8",X"CE",X"00",
		X"18",X"09",X"96",X"FD",X"77",X"06",X"3A",X"06",X"E8",X"DE",X"00",X"FD",X"77",X"07",X"23",X"3A",
		X"16",X"E9",X"5F",X"7E",X"93",X"5F",X"3A",X"07",X"E8",X"83",X"FD",X"77",X"02",X"3A",X"08",X"E8",
		X"CE",X"00",X"FD",X"77",X"03",X"23",X"7E",X"E6",X"1F",X"FD",X"77",X"00",X"7E",X"07",X"07",X"E6",
		X"03",X"B1",X"FD",X"77",X"05",X"23",X"7E",X"FD",X"77",X"04",X"11",X"08",X"00",X"FD",X"19",X"23",
		X"10",X"AA",X"FD",X"22",X"01",X"EB",X"78",X"32",X"00",X"EB",X"C9",X"21",X"A7",X"59",X"CD",X"1C",
		X"11",X"CD",X"A5",X"10",X"CD",X"AB",X"10",X"CD",X"CF",X"10",X"CD",X"D9",X"10",X"CD",X"E6",X"10",
		X"3A",X"1C",X"E8",X"A7",X"CC",X"1A",X"0F",X"3E",X"03",X"32",X"81",X"E8",X"3A",X"09",X"E7",X"32",
		X"1A",X"E8",X"3A",X"E2",X"E2",X"32",X"19",X"E8",X"CD",X"78",X"0F",X"CD",X"6B",X"0F",X"11",X"A0",
		X"D0",X"01",X"94",X"05",X"3E",X"A1",X"CD",X"10",X"11",X"3C",X"13",X"10",X"F9",X"3A",X"80",X"E0",
		X"E6",X"07",X"3C",X"67",X"3E",X"A6",X"11",X"E0",X"D0",X"CD",X"0A",X"0F",X"3C",X"11",X"20",X"D1",
		X"CD",X"0A",X"0F",X"11",X"E1",X"D0",X"0E",X"94",X"3E",X"A8",X"CD",X"01",X"0F",X"11",X"21",X"D1",
		X"3C",X"06",X"04",X"CD",X"10",X"11",X"13",X"10",X"FA",X"C9",X"6C",X"06",X"05",X"0E",X"94",X"CD",
		X"10",X"11",X"13",X"2D",X"20",X"01",X"0C",X"10",X"F6",X"C9",X"3A",X"80",X"E0",X"E6",X"F8",X"0F",
		X"0F",X"0F",X"47",X"DB",X"03",X"E6",X"01",X"20",X"01",X"05",X"78",X"A7",X"C8",X"FE",X"03",X"38",
		X"02",X"3E",X"03",X"47",X"0E",X"80",X"11",X"29",X"D1",X"CD",X"3F",X"0F",X"10",X"FB",X"C9",X"3E",
		X"B8",X"CD",X"4F",X"0F",X"D5",X"21",X"3E",X"00",X"19",X"EB",X"CD",X"4F",X"0F",X"D1",X"C9",X"CD",
		X"10",X"11",X"3C",X"CD",X"10",X"11",X"3C",X"C9",X"11",X"29",X"D1",X"AF",X"4F",X"CD",X"63",X"0F",
		X"11",X"69",X"D1",X"06",X"06",X"CD",X"10",X"11",X"10",X"FB",X"C9",X"11",X"16",X"D1",X"21",X"19",
		X"E8",X"3A",X"E2",X"E2",X"0E",X"15",X"18",X"0B",X"11",X"96",X"D0",X"21",X"1A",X"E8",X"3A",X"09",
		X"E7",X"0E",X"14",X"96",X"FA",X"8F",X"0F",X"FE",X"03",X"38",X"0A",X"3E",X"03",X"18",X"06",X"FE",
		X"FD",X"30",X"02",X"3E",X"FD",X"86",X"77",X"06",X"08",X"D6",X"08",X"6F",X"38",X"05",X"FA",X"AD",
		X"0F",X"3E",X"8A",X"C6",X"78",X"FE",X"77",X"20",X"08",X"3E",X"02",X"18",X"04",X"2E",X"FF",X"3E",
		X"03",X"CD",X"10",X"11",X"7D",X"10",X"E2",X"C9",X"3A",X"00",X"E0",X"FE",X"03",X"28",X"24",X"2A",
		X"03",X"E0",X"11",X"CD",X"FC",X"19",X"38",X"1B",X"21",X"08",X"E0",X"7E",X"A7",X"20",X"06",X"3E",
		X"00",X"CD",X"FE",X"0D",X"34",X"21",X"85",X"E8",X"7E",X"A7",X"20",X"07",X"36",X"38",X"3E",X"97",
		X"CD",X"FE",X"0D",X"21",X"1B",X"E8",X"3A",X"80",X"E8",X"BE",X"28",X"4E",X"77",X"CD",X"78",X"0F",
		X"CD",X"6B",X"0F",X"21",X"E0",X"D0",X"3A",X"80",X"E0",X"E6",X"07",X"87",X"5F",X"16",X"00",X"19",
		X"3A",X"80",X"E8",X"CB",X"DC",X"3A",X"80",X"E8",X"E6",X"18",X"3E",X"95",X"28",X"01",X"3D",X"77",
		X"11",X"40",X"00",X"19",X"77",X"3A",X"1C",X"E8",X"A7",X"20",X"3F",X"47",X"DB",X"03",X"E6",X"01",
		X"3A",X"80",X"E0",X"20",X"02",X"D6",X"08",X"FE",X"20",X"38",X"0F",X"3A",X"80",X"E8",X"E6",X"18",
		X"28",X"05",X"CD",X"1A",X"0F",X"18",X"03",X"CD",X"58",X"0F",X"3A",X"85",X"E0",X"E6",X"01",X"20",
		X"19",X"2A",X"81",X"E0",X"11",X"00",X"50",X"ED",X"52",X"38",X"0F",X"21",X"85",X"E0",X"CB",X"C6",
		X"2B",X"34",X"3E",X"98",X"CD",X"FE",X"0D",X"CD",X"E6",X"10",X"3A",X"00",X"E0",X"FE",X"03",X"28",
		X"1F",X"FE",X"0C",X"28",X"1B",X"21",X"81",X"E8",X"7E",X"A7",X"20",X"14",X"36",X"03",X"2A",X"03",
		X"E0",X"7D",X"D6",X"01",X"27",X"6F",X"7C",X"DE",X"00",X"27",X"67",X"38",X"03",X"22",X"03",X"E0",
		X"CD",X"D9",X"10",X"3A",X"83",X"E0",X"4F",X"ED",X"5B",X"81",X"E0",X"3A",X"82",X"E9",X"2A",X"80",
		X"E9",X"91",X"38",X"06",X"20",X"0F",X"ED",X"52",X"30",X"0B",X"79",X"32",X"82",X"E9",X"ED",X"53",
		X"80",X"E9",X"CD",X"CF",X"10",X"AF",X"11",X"83",X"E0",X"18",X"05",X"3E",X"01",X"11",X"93",X"E0",
		X"21",X"02",X"E0",X"AE",X"EB",X"E6",X"01",X"11",X"29",X"D0",X"20",X"03",X"11",X"14",X"D0",X"0E",
		X"15",X"7E",X"2B",X"CD",X"08",X"11",X"CD",X"FD",X"10",X"CD",X"FD",X"10",X"AF",X"18",X"39",X"21",
		X"82",X"E9",X"11",X"1F",X"D0",X"0E",X"00",X"18",X"E8",X"0E",X"14",X"21",X"04",X"E0",X"11",X"EA",
		X"D0",X"CD",X"FD",X"10",X"18",X"17",X"3A",X"84",X"E0",X"11",X"62",X"D1",X"6F",X"06",X"07",X"0E",
		X"03",X"3E",X"FE",X"2D",X"20",X"01",X"AF",X"CD",X"10",X"11",X"10",X"F7",X"C9",X"7E",X"2B",X"F5",
		X"0F",X"0F",X"0F",X"0F",X"CD",X"08",X"11",X"F1",X"E6",X"0F",X"C6",X"90",X"27",X"CE",X"40",X"27",
		X"EB",X"77",X"CB",X"DC",X"71",X"CB",X"9C",X"23",X"EB",X"C9",X"4E",X"23",X"7E",X"23",X"3C",X"C8",
		X"3C",X"28",X"F7",X"3C",X"28",X"07",X"D6",X"03",X"CD",X"10",X"11",X"18",X"EF",X"5E",X"23",X"56",
		X"18",X"E9",X"4E",X"23",X"7E",X"23",X"3C",X"C8",X"3C",X"28",X"F7",X"3C",X"28",X"10",X"D6",X"03",
		X"CD",X"10",X"11",X"FE",X"20",X"20",X"ED",X"3E",X"0B",X"CD",X"0F",X"57",X"18",X"E6",X"5E",X"23",
		X"56",X"18",X"E0",X"16",X"01",X"18",X"02",X"16",X"DB",X"1E",X"20",X"01",X"00",X"08",X"21",X"00",
		X"D0",X"FD",X"21",X"00",X"D8",X"73",X"FD",X"72",X"00",X"23",X"FD",X"23",X"0B",X"78",X"B1",X"20",
		X"F4",X"C9",X"AF",X"29",X"17",X"6C",X"67",X"D5",X"11",X"10",X"00",X"19",X"D1",X"22",X"15",X"E8",
		X"19",X"22",X"13",X"E8",X"3A",X"06",X"E7",X"87",X"5F",X"16",X"00",X"21",X"4D",X"66",X"19",X"5E",
		X"23",X"56",X"FD",X"21",X"00",X"00",X"FD",X"19",X"2A",X"17",X"E7",X"FD",X"7E",X"00",X"FE",X"FF",
		X"C8",X"5F",X"16",X"00",X"19",X"ED",X"5B",X"13",X"E8",X"ED",X"52",X"30",X"54",X"2A",X"17",X"E7",
		X"FD",X"5E",X"01",X"16",X"00",X"19",X"ED",X"5B",X"15",X"E8",X"ED",X"52",X"38",X"43",X"2A",X"12",
		X"E7",X"3A",X"01",X"E7",X"E6",X"40",X"28",X"0A",X"FD",X"5E",X"04",X"FD",X"56",X"05",X"ED",X"52",
		X"18",X"07",X"FD",X"5E",X"02",X"FD",X"56",X"03",X"19",X"A7",X"ED",X"5B",X"0F",X"E8",X"ED",X"52",
		X"38",X"1F",X"2A",X"12",X"E7",X"A7",X"28",X"0A",X"FD",X"5E",X"02",X"FD",X"56",X"03",X"ED",X"52",
		X"18",X"07",X"FD",X"5E",X"04",X"FD",X"56",X"05",X"19",X"A7",X"ED",X"5B",X"11",X"E8",X"ED",X"52",
		X"D8",X"11",X"06",X"00",X"FD",X"19",X"18",X"90",X"3A",X"00",X"E0",X"FE",X"06",X"C8",X"DB",X"04",
		X"2F",X"CB",X"77",X"C9",X"BE",X"38",X"05",X"23",X"BE",X"38",X"01",X"23",X"23",X"23",X"7E",X"C9",
		X"22",X"05",X"E8",X"3A",X"06",X"E7",X"21",X"6E",X"12",X"16",X"00",X"5F",X"19",X"7E",X"A7",X"C8",
		X"FD",X"21",X"90",X"12",X"87",X"87",X"5F",X"FD",X"19",X"2A",X"10",X"E7",X"FD",X"5E",X"02",X"FD",
		X"56",X"03",X"19",X"E5",X"FD",X"5E",X"00",X"FD",X"56",X"01",X"2A",X"12",X"E7",X"3A",X"01",X"E7",
		X"E6",X"40",X"28",X"03",X"19",X"18",X"02",X"ED",X"52",X"DD",X"5E",X"02",X"DD",X"56",X"03",X"ED",
		X"52",X"ED",X"5B",X"05",X"E8",X"38",X"04",X"ED",X"52",X"18",X"01",X"19",X"D1",X"C9",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"01",X"01",X"00",X"03",X"00",X"02",X"02",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"01",X"05",X"05",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"80",X"18",X"00",X"02",X"80",X"13",X"80",X"03",X"00",X"04",
		X"80",X"03",X"80",X"18",X"A0",X"02",X"00",X"18",X"20",X"03",X"80",X"0F",X"21",X"00",X"E7",X"CB",
		X"4E",X"20",X"12",X"21",X"00",X"E2",X"CD",X"CB",X"12",X"CD",X"FE",X"12",X"CD",X"8F",X"13",X"CD",
		X"EE",X"13",X"CD",X"3F",X"14",X"CD",X"3D",X"15",X"C9",X"23",X"23",X"7E",X"A7",X"C8",X"35",X"C2",
		X"C9",X"12",X"23",X"4E",X"06",X"00",X"EB",X"21",X"0A",X"E1",X"09",X"09",X"CB",X"BE",X"2A",X"08",
		X"E1",X"ED",X"A8",X"ED",X"A8",X"22",X"08",X"E1",X"23",X"36",X"00",X"EB",X"C3",X"CA",X"12",X"00",
		X"00",X"00",X"01",X"01",X"01",X"02",X"02",X"02",X"03",X"03",X"03",X"04",X"04",X"04",X"3A",X"01",
		X"E7",X"E6",X"80",X"0E",X"E4",X"28",X"02",X"0E",X"1C",X"3A",X"13",X"E7",X"81",X"FE",X"E0",X"D0",
		X"32",X"09",X"E8",X"5F",X"E6",X"0F",X"3D",X"F8",X"21",X"EF",X"12",X"06",X"00",X"4F",X"09",X"4E",
		X"7B",X"E6",X"F0",X"0F",X"0F",X"5F",X"0F",X"0F",X"83",X"81",X"4F",X"DD",X"21",X"0A",X"E1",X"DD",
		X"09",X"DD",X"09",X"DD",X"CB",X"00",X"7E",X"C0",X"2A",X"08",X"E1",X"11",X"13",X"E2",X"ED",X"52",
		X"C8",X"47",X"3A",X"01",X"E7",X"E6",X"80",X"21",X"35",X"E2",X"11",X"9A",X"E1",X"28",X"04",X"21",
		X"15",X"E2",X"13",X"7E",X"A7",X"C0",X"23",X"7E",X"FE",X"0A",X"D0",X"E5",X"D5",X"34",X"23",X"5F",
		X"87",X"83",X"16",X"00",X"5F",X"19",X"72",X"23",X"3A",X"09",X"E8",X"77",X"23",X"DD",X"7E",X"00",
		X"77",X"DD",X"7E",X"01",X"2A",X"08",X"E1",X"23",X"77",X"23",X"71",X"22",X"08",X"E1",X"DD",X"CB",
		X"00",X"FE",X"E1",X"D1",X"35",X"C0",X"3A",X"99",X"E1",X"77",X"EB",X"2B",X"36",X"01",X"C9",X"21",
		X"36",X"E2",X"7E",X"A7",X"C8",X"47",X"16",X"00",X"23",X"7E",X"C6",X"36",X"77",X"23",X"7E",X"8A",
		X"D2",X"A4",X"13",X"3D",X"77",X"23",X"23",X"10",X"F0",X"2A",X"37",X"E2",X"7C",X"FE",X"BE",X"30",
		X"0B",X"01",X"00",X"12",X"09",X"ED",X"4B",X"12",X"E7",X"ED",X"42",X"D8",X"21",X"55",X"E2",X"7E",
		X"FE",X"0A",X"D0",X"34",X"5F",X"21",X"56",X"E2",X"19",X"3A",X"39",X"E2",X"F6",X"58",X"77",X"EB",
		X"21",X"36",X"E2",X"35",X"28",X"10",X"7E",X"11",X"37",X"E2",X"21",X"3A",X"E2",X"4F",X"87",X"81",
		X"4F",X"06",X"00",X"ED",X"B0",X"C9",X"2B",X"7E",X"A7",X"C8",X"EB",X"CB",X"C6",X"C9",X"21",X"16",
		X"E2",X"7E",X"A7",X"C8",X"47",X"16",X"00",X"23",X"7E",X"D6",X"36",X"77",X"23",X"7E",X"9A",X"D2",
		X"03",X"14",X"3C",X"77",X"23",X"23",X"10",X"F0",X"2A",X"17",X"E2",X"7C",X"FE",X"22",X"38",X"0C",
		X"01",X"00",X"12",X"ED",X"42",X"ED",X"4B",X"12",X"E7",X"ED",X"42",X"D0",X"21",X"55",X"E2",X"7E",
		X"FE",X"0A",X"D0",X"34",X"5F",X"21",X"56",X"E2",X"19",X"3A",X"19",X"E2",X"F6",X"30",X"77",X"EB",
		X"21",X"16",X"E2",X"35",X"28",X"B0",X"7E",X"11",X"17",X"E2",X"21",X"1A",X"E2",X"18",X"9E",X"3A",
		X"60",X"E2",X"47",X"EE",X"28",X"C8",X"3A",X"D8",X"E2",X"E6",X"10",X"3A",X"96",X"E1",X"28",X"03",
		X"3A",X"97",X"E1",X"A7",X"28",X"06",X"4F",X"3A",X"61",X"E2",X"B9",X"D0",X"21",X"55",X"E2",X"7E",
		X"A7",X"C8",X"4F",X"23",X"CB",X"76",X"20",X"0D",X"CB",X"68",X"28",X"53",X"0D",X"C8",X"23",X"CB",
		X"76",X"28",X"F9",X"18",X"04",X"CB",X"58",X"20",X"3F",X"CD",X"24",X"15",X"F5",X"2A",X"12",X"E7",
		X"11",X"00",X"12",X"ED",X"52",X"11",X"00",X"BE",X"ED",X"52",X"30",X"02",X"19",X"EB",X"3A",X"D8",
		X"E2",X"6F",X"CB",X"65",X"28",X"1B",X"3A",X"97",X"E1",X"A7",X"28",X"0B",X"CB",X"75",X"28",X"11",
		X"2A",X"DA",X"E2",X"ED",X"52",X"38",X"0A",X"21",X"35",X"E2",X"F1",X"E6",X"01",X"C8",X"36",X"00",
		X"C9",X"21",X"60",X"E2",X"CB",X"DE",X"18",X"3E",X"0D",X"C8",X"23",X"CB",X"76",X"20",X"F9",X"CD",
		X"24",X"15",X"F5",X"2A",X"12",X"E7",X"11",X"00",X"12",X"19",X"11",X"00",X"22",X"ED",X"52",X"38",
		X"02",X"19",X"EB",X"3A",X"D8",X"E2",X"6F",X"CB",X"65",X"28",X"16",X"3A",X"97",X"E1",X"A7",X"28",
		X"0B",X"CB",X"75",X"20",X"0C",X"2A",X"DA",X"E2",X"ED",X"52",X"30",X"05",X"21",X"15",X"E2",X"18",
		X"B9",X"21",X"60",X"E2",X"CB",X"EE",X"21",X"61",X"E2",X"34",X"23",X"01",X"10",X"00",X"7E",X"A7",
		X"28",X"03",X"09",X"18",X"F9",X"F1",X"77",X"AF",X"23",X"36",X"00",X"23",X"73",X"23",X"72",X"23",
		X"36",X"00",X"23",X"36",X"50",X"23",X"77",X"23",X"36",X"07",X"23",X"77",X"23",X"77",X"23",X"36",
		X"02",X"23",X"77",X"C9",X"7E",X"0D",X"28",X"07",X"54",X"5D",X"23",X"06",X"00",X"ED",X"B0",X"21",
		X"55",X"E2",X"35",X"C9",X"C1",X"11",X"10",X"00",X"DD",X"19",X"10",X"1A",X"C9",X"3A",X"01",X"E7",
		X"E6",X"03",X"20",X"03",X"32",X"D2",X"E2",X"21",X"01",X"01",X"22",X"1B",X"E7",X"22",X"1D",X"E7",
		X"DD",X"21",X"62",X"E2",X"06",X"05",X"C5",X"21",X"34",X"15",X"E5",X"DD",X"4E",X"00",X"CB",X"61",
		X"C8",X"CB",X"69",X"C4",X"26",X"1C",X"CB",X"59",X"C4",X"3D",X"1C",X"CB",X"41",X"DD",X"7E",X"01",
		X"C2",X"6E",X"18",X"CB",X"51",X"C2",X"8A",X"16",X"21",X"2F",X"16",X"E5",X"21",X"00",X"E7",X"CB",
		X"4E",X"C2",X"E2",X"1B",X"FE",X"01",X"CA",X"AA",X"1B",X"38",X"47",X"FE",X"09",X"CA",X"DD",X"15",
		X"30",X"16",X"CD",X"EF",X"1B",X"11",X"00",X"EF",X"19",X"D0",X"CD",X"7A",X"1B",X"79",X"E6",X"28",
		X"2F",X"21",X"60",X"E2",X"A6",X"77",X"E1",X"C9",X"CD",X"E7",X"1B",X"DD",X"7E",X"06",X"FE",X"0A",
		X"30",X"04",X"DD",X"36",X"06",X"0D",X"CD",X"3E",X"16",X"D8",X"11",X"00",X"FF",X"2A",X"0C",X"E8",
		X"19",X"D2",X"20",X"1B",X"C9",X"3E",X"0A",X"DD",X"86",X"06",X"DD",X"77",X"06",X"DD",X"36",X"01",
		X"0A",X"C9",X"CD",X"E7",X"1B",X"11",X"00",X"F8",X"19",X"D2",X"C5",X"15",X"C9",X"CD",X"54",X"1B",
		X"CD",X"61",X"1C",X"DD",X"BE",X"0F",X"28",X"0A",X"DD",X"35",X"0B",X"28",X"39",X"DD",X"77",X"0F",
		X"18",X"09",X"DD",X"35",X"0E",X"20",X"08",X"DD",X"36",X"0B",X"06",X"DD",X"36",X"0E",X"05",X"DD",
		X"35",X"07",X"C0",X"3A",X"1C",X"E8",X"A7",X"3E",X"02",X"20",X"0A",X"DB",X"03",X"E6",X"02",X"3E",
		X"04",X"20",X"02",X"3E",X"03",X"DD",X"77",X"07",X"21",X"09",X"E7",X"7E",X"A7",X"F8",X"35",X"F0",
		X"21",X"1F",X"E7",X"CB",X"CE",X"C9",X"21",X"1A",X"E7",X"35",X"3E",X"09",X"C3",X"90",X"1B",X"21",
		X"7B",X"6A",X"DD",X"7E",X"01",X"FE",X"05",X"C2",X"7D",X"1A",X"79",X"C3",X"80",X"1A",X"11",X"80",
		X"16",X"CD",X"D2",X"1A",X"D0",X"F5",X"3E",X"91",X"CD",X"FE",X"0D",X"F1",X"FA",X"53",X"16",X"3E",
		X"80",X"18",X"24",X"21",X"D2",X"E2",X"34",X"CD",X"C9",X"1A",X"7E",X"20",X"0E",X"FE",X"02",X"3E",
		X"80",X"38",X"14",X"3E",X"82",X"28",X"10",X"3E",X"85",X"18",X"0C",X"FE",X"02",X"3E",X"8C",X"38",
		X"06",X"3E",X"80",X"28",X"02",X"3E",X"82",X"21",X"D2",X"00",X"EB",X"CD",X"60",X"2F",X"37",X"C9",
		X"F2",X"F0",X"F2",X"F2",X"F2",X"02",X"01",X"FF",X"FF",X"FF",X"21",X"22",X"18",X"E5",X"21",X"00",
		X"E7",X"CB",X"4E",X"C2",X"E2",X"1B",X"FE",X"09",X"CA",X"DD",X"15",X"D2",X"0B",X"17",X"FE",X"01",
		X"CA",X"AA",X"1B",X"D2",X"92",X"15",X"CD",X"E7",X"1B",X"CD",X"28",X"18",X"D8",X"2A",X"0C",X"E8",
		X"11",X"00",X"E1",X"19",X"DA",X"7A",X"1B",X"DD",X"CB",X"0B",X"46",X"20",X"26",X"2A",X"0C",X"E8",
		X"11",X"00",X"FA",X"19",X"38",X"1D",X"DD",X"CB",X"0B",X"C6",X"3A",X"02",X"E7",X"FE",X"03",X"28",
		X"08",X"FE",X"06",X"28",X"04",X"FE",X"07",X"20",X"0A",X"3A",X"13",X"E0",X"21",X"C1",X"E1",X"BE",
		X"DA",X"E5",X"17",X"2A",X"10",X"E7",X"11",X"80",X"A1",X"19",X"D8",X"2A",X"0A",X"E8",X"11",X"C0",
		X"00",X"CB",X"71",X"28",X"03",X"19",X"18",X"02",X"ED",X"52",X"DA",X"20",X"1B",X"C9",X"DD",X"36",
		X"01",X"00",X"DD",X"36",X"06",X"00",X"DD",X"36",X"07",X"07",X"C9",X"DD",X"5E",X"0E",X"DD",X"56",
		X"0F",X"DD",X"7E",X"06",X"FE",X"0A",X"F5",X"C4",X"70",X"1C",X"CD",X"E2",X"1B",X"F1",X"28",X"1D",
		X"11",X"D6",X"FF",X"CD",X"AC",X"1C",X"19",X"CD",X"A5",X"1C",X"EB",X"CD",X"9E",X"1C",X"19",X"11",
		X"00",X"50",X"ED",X"52",X"19",X"30",X"01",X"EB",X"CD",X"97",X"1C",X"38",X"C1",X"DD",X"CB",X"0B",
		X"4E",X"20",X"1C",X"CD",X"8A",X"1C",X"11",X"60",X"FF",X"19",X"22",X"0F",X"E8",X"11",X"40",X"01",
		X"19",X"22",X"11",X"E8",X"CD",X"9E",X"1C",X"11",X"14",X"00",X"CD",X"72",X"11",X"38",X"28",X"DD",
		X"35",X"07",X"20",X"18",X"DD",X"7E",X"0A",X"3C",X"DD",X"77",X"0A",X"87",X"5F",X"16",X"00",X"21",
		X"FC",X"17",X"19",X"7E",X"DD",X"77",X"07",X"23",X"7E",X"DD",X"77",X"06",X"DD",X"7E",X"06",X"FE",
		X"0F",X"D8",X"79",X"EE",X"C0",X"4F",X"C9",X"3A",X"02",X"E7",X"FE",X"03",X"28",X"08",X"FE",X"06",
		X"28",X"04",X"FE",X"07",X"20",X"24",X"CD",X"9E",X"1C",X"11",X"0C",X"01",X"3E",X"91",X"CD",X"FE",
		X"0D",X"CD",X"E2",X"2E",X"3E",X"07",X"F5",X"CD",X"AC",X"1C",X"EB",X"21",X"00",X"00",X"ED",X"52",
		X"CD",X"A5",X"1C",X"DD",X"CB",X"0B",X"CE",X"F1",X"18",X"AE",X"DD",X"36",X"06",X"09",X"CD",X"9E",
		X"1C",X"11",X"00",X"0A",X"19",X"AF",X"29",X"07",X"6C",X"67",X"EB",X"CD",X"8A",X"1C",X"CD",X"C9",
		X"1A",X"3E",X"80",X"20",X"02",X"3E",X"82",X"CD",X"60",X"2F",X"3E",X"91",X"CD",X"FE",X"0D",X"21",
		X"5B",X"1C",X"C3",X"96",X"1B",X"DD",X"36",X"01",X"0A",X"21",X"A0",X"03",X"CD",X"A5",X"1C",X"21",
		X"28",X"00",X"DD",X"75",X"0E",X"DD",X"74",X"0F",X"AF",X"C3",X"68",X"17",X"03",X"0A",X"07",X"0C",
		X"07",X"0D",X"07",X"0E",X"07",X"0F",X"07",X"10",X"FF",X"0B",X"03",X"0A",X"07",X"0D",X"07",X"0E",
		X"07",X"0F",X"07",X"10",X"FF",X"0B",X"03",X"0A",X"07",X"10",X"07",X"0F",X"07",X"0E",X"07",X"0D",
		X"FF",X"0B",X"21",X"2F",X"6B",X"C3",X"32",X"16",X"11",X"64",X"18",X"CD",X"D2",X"1A",X"D0",X"F5",
		X"3A",X"0B",X"E8",X"E6",X"80",X"CB",X"B1",X"28",X"02",X"CB",X"F1",X"DD",X"71",X"00",X"3E",X"91",
		X"CD",X"FE",X"0D",X"F1",X"FA",X"4B",X"18",X"3E",X"81",X"18",X"13",X"21",X"D2",X"E2",X"34",X"7E",
		X"FE",X"02",X"3E",X"80",X"DA",X"77",X"16",X"3E",X"81",X"CA",X"77",X"16",X"3E",X"84",X"21",X"BE",
		X"00",X"C3",X"7A",X"16",X"FF",X"F0",X"FF",X"FF",X"FF",X"FF",X"01",X"FF",X"FF",X"FF",X"21",X"72",
		X"1A",X"E5",X"21",X"00",X"E7",X"CB",X"4E",X"20",X"2A",X"DD",X"6E",X"08",X"DD",X"66",X"09",X"2B",
		X"CB",X"7C",X"20",X"06",X"DD",X"75",X"08",X"DD",X"74",X"09",X"87",X"16",X"00",X"5F",X"21",X"97",
		X"18",X"19",X"7E",X"23",X"66",X"6F",X"E9",X"28",X"1A",X"AA",X"1B",X"6C",X"19",X"C2",X"19",X"AE",
		X"18",X"99",X"19",X"F5",X"CD",X"E2",X"1B",X"F1",X"FE",X"05",X"CA",X"BD",X"19",X"C9",X"CD",X"E2",
		X"1B",X"CD",X"49",X"1A",X"30",X"20",X"DD",X"35",X"0A",X"F5",X"3E",X"91",X"CD",X"FE",X"0D",X"F1",
		X"28",X"04",X"DD",X"34",X"01",X"C9",X"CD",X"77",X"16",X"21",X"15",X"E2",X"CB",X"71",X"28",X"03",
		X"21",X"35",X"E2",X"36",X"00",X"C9",X"11",X"00",X"FF",X"2A",X"0C",X"E8",X"19",X"38",X"0B",X"3E",
		X"05",X"21",X"5A",X"00",X"DD",X"36",X"06",X"02",X"18",X"65",X"DD",X"7E",X"08",X"A7",X"CA",X"FD",
		X"19",X"DD",X"7E",X"06",X"FE",X"02",X"28",X"65",X"DD",X"35",X"07",X"C0",X"DD",X"7E",X"0E",X"A7",
		X"C2",X"42",X"19",X"21",X"2B",X"E3",X"7E",X"FE",X"03",X"DD",X"34",X"07",X"D0",X"87",X"86",X"34",
		X"23",X"16",X"00",X"5F",X"19",X"E5",X"CD",X"8A",X"1C",X"11",X"C0",X"00",X"79",X"E6",X"40",X"28",
		X"03",X"19",X"18",X"02",X"ED",X"52",X"EB",X"E1",X"47",X"DD",X"7E",X"06",X"D6",X"09",X"B0",X"77",
		X"23",X"73",X"23",X"72",X"CD",X"BF",X"1D",X"DD",X"35",X"0E",X"DD",X"36",X"07",X"10",X"DD",X"34",
		X"06",X"C9",X"DD",X"36",X"06",X"02",X"DD",X"35",X"0B",X"C0",X"2A",X"F5",X"E1",X"3E",X"03",X"DD",
		X"75",X"08",X"DD",X"74",X"09",X"DD",X"77",X"01",X"DD",X"36",X"07",X"02",X"C9",X"2A",X"0C",X"E8",
		X"11",X"A0",X"F5",X"19",X"21",X"5A",X"00",X"3E",X"00",X"38",X"E4",X"C9",X"CD",X"E2",X"1B",X"3E",
		X"02",X"DD",X"BE",X"06",X"28",X"0C",X"DD",X"35",X"07",X"C0",X"DD",X"77",X"06",X"DD",X"36",X"07",
		X"03",X"C9",X"CD",X"49",X"1A",X"DA",X"B6",X"18",X"DD",X"35",X"07",X"C0",X"DD",X"36",X"08",X"04",
		X"DD",X"36",X"09",X"00",X"DD",X"36",X"01",X"03",X"C9",X"CD",X"EF",X"1B",X"CD",X"49",X"1A",X"DA",
		X"B6",X"18",X"DD",X"7E",X"08",X"A7",X"20",X"06",X"DD",X"7E",X"09",X"A7",X"28",X"45",X"11",X"00",
		X"F6",X"2A",X"0C",X"E8",X"19",X"DA",X"3C",X"1A",X"CD",X"B8",X"1A",X"38",X"7F",X"79",X"EE",X"40",
		X"4F",X"C9",X"CD",X"E2",X"1B",X"CD",X"49",X"1A",X"DA",X"B6",X"18",X"DD",X"7E",X"08",X"A7",X"20",
		X"06",X"DD",X"7E",X"09",X"A7",X"28",X"1C",X"11",X"00",X"F7",X"2A",X"0C",X"E8",X"19",X"30",X"0A",
		X"11",X"00",X"FE",X"19",X"D0",X"DD",X"36",X"01",X"00",X"C9",X"CD",X"B8",X"1A",X"D8",X"DD",X"36",
		X"01",X"05",X"C9",X"DD",X"36",X"01",X"04",X"3A",X"F0",X"E1",X"DD",X"77",X"0B",X"21",X"F1",X"E1",
		X"3A",X"10",X"E0",X"BE",X"3E",X"09",X"38",X"02",X"3E",X"0B",X"DD",X"77",X"06",X"23",X"3A",X"11",
		X"E0",X"FE",X"55",X"38",X"06",X"23",X"FE",X"AA",X"38",X"01",X"23",X"7E",X"DD",X"77",X"08",X"DD",
		X"36",X"0E",X"00",X"DD",X"36",X"07",X"0B",X"C9",X"CD",X"E7",X"1B",X"11",X"00",X"F6",X"19",X"D8",
		X"DD",X"7E",X"08",X"A7",X"20",X"06",X"DD",X"7E",X"09",X"A7",X"28",X"B7",X"DD",X"36",X"01",X"03",
		X"DD",X"36",X"06",X"02",X"DD",X"36",X"07",X"02",X"C9",X"3A",X"01",X"E7",X"E6",X"03",X"20",X"04",
		X"DD",X"CB",X"00",X"96",X"DD",X"CB",X"00",X"56",X"C0",X"11",X"80",X"16",X"CD",X"D2",X"1A",X"D0",
		X"DD",X"CB",X"00",X"D6",X"3E",X"85",X"F0",X"CD",X"C9",X"1A",X"3E",X"83",X"20",X"02",X"3E",X"87",
		X"37",X"C9",X"2A",X"0C",X"E8",X"11",X"00",X"E4",X"19",X"D8",X"21",X"E7",X"6B",X"79",X"EE",X"40",
		X"E6",X"C0",X"DD",X"CB",X"00",X"66",X"C8",X"EB",X"CD",X"9E",X"1C",X"29",X"6C",X"26",X"00",X"CB",
		X"14",X"22",X"07",X"E8",X"2A",X"0A",X"E8",X"DD",X"4E",X"06",X"D5",X"06",X"00",X"16",X"FF",X"29",
		X"38",X"01",X"50",X"29",X"29",X"5C",X"2A",X"15",X"E7",X"19",X"22",X"03",X"E8",X"EB",X"E1",X"09",
		X"09",X"4E",X"23",X"66",X"69",X"C3",X"20",X"0E",X"CD",X"91",X"1C",X"2A",X"06",X"E1",X"CB",X"71",
		X"28",X"04",X"2A",X"04",X"E1",X"EB",X"ED",X"52",X"C9",X"3A",X"02",X"E7",X"FE",X"08",X"C8",X"FE",
		X"09",X"C9",X"D5",X"CD",X"E7",X"1A",X"E1",X"D0",X"CD",X"18",X"1B",X"D0",X"F5",X"E6",X"0F",X"CD",
		X"8E",X"1B",X"CD",X"91",X"1C",X"F1",X"C9",X"3A",X"0B",X"E8",X"47",X"3A",X"01",X"E7",X"07",X"A8",
		X"E6",X"80",X"C8",X"3A",X"01",X"E7",X"E6",X"03",X"C8",X"E6",X"02",X"11",X"C0",X"02",X"06",X"05",
		X"20",X"04",X"11",X"00",X"04",X"47",X"ED",X"52",X"D0",X"3A",X"02",X"E7",X"FE",X"06",X"D8",X"04",
		X"D6",X"08",X"D8",X"04",X"80",X"47",X"37",X"C9",X"58",X"16",X"00",X"19",X"7E",X"FE",X"FF",X"C9",
		X"CD",X"08",X"12",X"20",X"55",X"3A",X"1C",X"E8",X"A7",X"3E",X"02",X"20",X"0A",X"DB",X"03",X"E6",
		X"02",X"3E",X"04",X"20",X"02",X"3E",X"03",X"DD",X"77",X"07",X"DD",X"36",X"06",X"09",X"DD",X"36",
		X"01",X"09",X"21",X"1A",X"E7",X"34",X"CD",X"61",X"1C",X"DD",X"77",X"0F",X"DD",X"36",X"0B",X"06",
		X"DD",X"36",X"0E",X"05",X"DD",X"CB",X"00",X"56",X"21",X"1B",X"E7",X"28",X"02",X"23",X"23",X"DD",
		X"CB",X"00",X"76",X"11",X"80",X"FF",X"20",X"04",X"23",X"11",X"80",X"00",X"34",X"46",X"2A",X"12",
		X"E7",X"19",X"10",X"FD",X"CD",X"83",X"1C",X"C3",X"E2",X"1B",X"DD",X"CB",X"00",X"4E",X"20",X"09",
		X"DD",X"36",X"00",X"00",X"21",X"61",X"E2",X"35",X"C9",X"DD",X"CB",X"00",X"A6",X"C9",X"C6",X"04",
		X"DD",X"77",X"06",X"21",X"55",X"1C",X"DD",X"36",X"01",X"01",X"7E",X"23",X"DD",X"77",X"07",X"CD",
		X"A5",X"1C",X"AF",X"DD",X"77",X"0E",X"DD",X"77",X"0F",X"C9",X"DD",X"35",X"07",X"C2",X"C4",X"1B",
		X"CD",X"AC",X"1C",X"7E",X"A7",X"FA",X"7A",X"1B",X"23",X"DD",X"77",X"06",X"7E",X"23",X"DD",X"77",
		X"07",X"CD",X"A5",X"1C",X"DD",X"5E",X"0E",X"DD",X"56",X"0F",X"21",X"16",X"00",X"19",X"DD",X"75",
		X"0E",X"DD",X"74",X"0F",X"CD",X"9E",X"1C",X"ED",X"52",X"CD",X"97",X"1C",X"11",X"39",X"00",X"CD",
		X"7A",X"1C",X"CD",X"8A",X"1C",X"18",X"21",X"11",X"36",X"00",X"CD",X"70",X"1C",X"18",X"06",X"11",
		X"36",X"00",X"CD",X"7A",X"1C",X"DD",X"35",X"07",X"20",X"0E",X"DD",X"36",X"07",X"07",X"DD",X"35",
		X"06",X"F2",X"08",X"1C",X"DD",X"36",X"06",X"03",X"ED",X"5B",X"12",X"E7",X"7B",X"E6",X"E0",X"5F",
		X"7D",X"E6",X"E0",X"6F",X"ED",X"52",X"22",X"0A",X"E8",X"30",X"06",X"11",X"01",X"00",X"EB",X"ED",
		X"52",X"22",X"0C",X"E8",X"A7",X"C9",X"2A",X"12",X"E7",X"11",X"00",X"10",X"19",X"CD",X"91",X"1C",
		X"ED",X"52",X"D8",X"DD",X"CB",X"00",X"AE",X"21",X"60",X"E2",X"CB",X"AE",X"C9",X"CD",X"8A",X"1C",
		X"11",X"00",X"10",X"19",X"ED",X"5B",X"12",X"E7",X"ED",X"52",X"D8",X"DD",X"CB",X"00",X"9E",X"21",
		X"60",X"E2",X"CB",X"9E",X"C9",X"05",X"07",X"07",X"08",X"11",X"FF",X"05",X"07",X"0A",X"08",X"17",
		X"FF",X"3A",X"00",X"E0",X"FE",X"06",X"3A",X"09",X"E9",X"C8",X"3A",X"07",X"E9",X"E6",X"0F",X"C9",
		X"CD",X"8A",X"1C",X"CB",X"71",X"28",X"0A",X"19",X"18",X"09",X"CD",X"8A",X"1C",X"CB",X"71",X"28",
		X"F6",X"ED",X"52",X"DD",X"75",X"02",X"DD",X"74",X"03",X"C9",X"DD",X"6E",X"02",X"DD",X"66",X"03",
		X"C9",X"EB",X"CD",X"8A",X"1C",X"EB",X"C9",X"DD",X"75",X"04",X"DD",X"74",X"05",X"C9",X"DD",X"6E",
		X"04",X"DD",X"66",X"05",X"C9",X"DD",X"75",X"0C",X"DD",X"74",X"0D",X"C9",X"DD",X"6E",X"0C",X"DD",
		X"66",X"0D",X"C9",X"CD",X"4A",X"1E",X"CD",X"FD",X"1D",X"DD",X"21",X"FB",X"E2",X"CD",X"C4",X"1C",
		X"DD",X"21",X"0B",X"E3",X"DD",X"7E",X"00",X"4F",X"E6",X"10",X"C8",X"3A",X"00",X"E7",X"E6",X"02",
		X"C2",X"A7",X"1D",X"DD",X"7E",X"01",X"FE",X"01",X"DA",X"4B",X"1D",X"28",X"26",X"CD",X"E9",X"1D",
		X"3A",X"D9",X"E2",X"FE",X"01",X"28",X"07",X"3A",X"D8",X"E2",X"E6",X"10",X"20",X"6D",X"ED",X"5B",
		X"12",X"E7",X"ED",X"52",X"DA",X"5B",X"1D",X"11",X"00",X"EC",X"19",X"30",X"5E",X"DD",X"36",X"00",
		X"00",X"18",X"58",X"DD",X"7E",X"0B",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"CB",X"47",X"28",X"0C",
		X"ED",X"5B",X"BF",X"E1",X"FE",X"03",X"28",X"08",X"ED",X"52",X"18",X"05",X"ED",X"5B",X"BD",X"E1",
		X"19",X"DD",X"75",X"04",X"DD",X"74",X"05",X"DD",X"6E",X"0C",X"DD",X"66",X"0D",X"ED",X"5B",X"BB",
		X"E1",X"19",X"DD",X"75",X"0C",X"DD",X"74",X"0D",X"CD",X"EF",X"1D",X"DD",X"5E",X"0E",X"DD",X"56",
		X"0F",X"ED",X"52",X"38",X"16",X"DD",X"CB",X"00",X"AE",X"18",X"0D",X"CD",X"E9",X"1D",X"DD",X"5E",
		X"0E",X"DD",X"56",X"0F",X"ED",X"52",X"30",X"03",X"DD",X"34",X"01",X"DD",X"CB",X"00",X"6E",X"20",
		X"2E",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"11",X"40",X"FF",X"19",X"22",X"0F",X"E8",X"11",X"80",
		X"01",X"19",X"22",X"11",X"E8",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"11",X"08",X"00",X"E5",X"CD",
		X"72",X"11",X"E1",X"30",X"0A",X"11",X"18",X"01",X"CD",X"9A",X"2C",X"DD",X"CB",X"00",X"EE",X"DD",
		X"35",X"07",X"20",X"13",X"DD",X"36",X"07",X"02",X"DD",X"7E",X"06",X"3C",X"FE",X"06",X"38",X"04",
		X"CD",X"BF",X"1D",X"AF",X"DD",X"77",X"06",X"CD",X"E2",X"1B",X"11",X"00",X"E8",X"19",X"D8",X"DD",
		X"7E",X"06",X"FE",X"03",X"3E",X"40",X"38",X"01",X"AF",X"21",X"A5",X"75",X"C3",X"7E",X"1A",X"E5",
		X"D5",X"2A",X"03",X"E0",X"11",X"CD",X"FC",X"19",X"3E",X"95",X"38",X"02",X"3E",X"99",X"CD",X"FE",
		X"0D",X"D1",X"E1",X"C9",X"E5",X"D5",X"2A",X"03",X"E0",X"11",X"CD",X"FC",X"19",X"3E",X"92",X"38",
		X"02",X"3E",X"9A",X"CD",X"FE",X"0D",X"D1",X"E1",X"C9",X"DD",X"6E",X"0C",X"DD",X"66",X"0D",X"DD",
		X"5E",X"02",X"DD",X"56",X"03",X"19",X"DD",X"75",X"02",X"DD",X"74",X"03",X"C9",X"DD",X"21",X"1B",
		X"E3",X"DD",X"4E",X"00",X"CB",X"61",X"C8",X"DD",X"35",X"07",X"20",X"14",X"DD",X"36",X"07",X"05",
		X"DD",X"34",X"06",X"3A",X"21",X"E3",X"FE",X"04",X"38",X"06",X"20",X"29",X"DD",X"CB",X"00",X"FE",
		X"11",X"72",X"00",X"CD",X"7A",X"1C",X"CD",X"E2",X"1B",X"2A",X"27",X"E3",X"11",X"1B",X"00",X"19",
		X"22",X"27",X"E3",X"EB",X"2A",X"1F",X"E3",X"ED",X"52",X"22",X"1F",X"E3",X"21",X"D2",X"73",X"3A",
		X"1B",X"E3",X"C3",X"7E",X"1A",X"DD",X"36",X"00",X"00",X"C9",X"3A",X"D8",X"E2",X"4F",X"A7",X"28",
		X"3D",X"E6",X"10",X"C8",X"2A",X"E0",X"E2",X"2B",X"CB",X"7C",X"20",X"03",X"22",X"E0",X"E2",X"DD",
		X"21",X"D8",X"E2",X"3A",X"E2",X"E2",X"21",X"FA",X"E2",X"A7",X"FA",X"77",X"1E",X"FE",X"3F",X"28",
		X"06",X"35",X"20",X"05",X"DD",X"34",X"0A",X"36",X"70",X"3A",X"80",X"E0",X"E6",X"07",X"21",X"84",
		X"1E",X"C3",X"26",X"1F",X"19",X"1F",X"98",X"22",X"3E",X"21",X"F0",X"24",X"F2",X"28",X"3A",X"80",
		X"E0",X"E6",X"07",X"2A",X"D3",X"E2",X"ED",X"5B",X"12",X"E7",X"ED",X"52",X"CB",X"47",X"28",X"01",
		X"3F",X"D8",X"FE",X"03",X"20",X"06",X"21",X"4F",X"03",X"22",X"F8",X"E2",X"CB",X"47",X"4F",X"3E",
		X"12",X"20",X"02",X"3E",X"52",X"32",X"D8",X"E2",X"3E",X"70",X"32",X"FA",X"E2",X"3A",X"61",X"E2",
		X"21",X"97",X"E1",X"96",X"D8",X"C8",X"06",X"05",X"DD",X"21",X"62",X"E2",X"DD",X"CB",X"00",X"46",
		X"20",X"31",X"2A",X"12",X"E7",X"DD",X"5E",X"02",X"DD",X"56",X"03",X"CB",X"41",X"28",X"0C",X"DD",
		X"CB",X"00",X"76",X"28",X"1E",X"ED",X"52",X"38",X"1A",X"18",X"0A",X"DD",X"CB",X"00",X"76",X"20",
		X"12",X"ED",X"52",X"30",X"0E",X"6F",X"DD",X"7E",X"01",X"A7",X"7D",X"20",X"06",X"DD",X"36",X"01",
		X"05",X"3D",X"C8",X"11",X"10",X"00",X"DD",X"19",X"10",X"C2",X"C9",X"30",X"1F",X"F9",X"1F",X"11",
		X"20",X"45",X"1F",X"59",X"1F",X"64",X"20",X"1B",X"20",X"CD",X"6F",X"2C",X"21",X"96",X"20",X"E5",
		X"21",X"0B",X"1F",X"DD",X"7E",X"01",X"87",X"16",X"00",X"5F",X"19",X"7E",X"23",X"66",X"6F",X"E9",
		X"CD",X"0D",X"2D",X"11",X"00",X"FA",X"19",X"D2",X"CF",X"1F",X"11",X"00",X"C0",X"2A",X"DA",X"E2",
		X"19",X"DA",X"50",X"1F",X"C9",X"CD",X"E2",X"1B",X"11",X"00",X"FA",X"19",X"D2",X"CF",X"1F",X"C9",
		X"DD",X"36",X"01",X"03",X"DD",X"36",X"06",X"00",X"C9",X"CD",X"E2",X"1B",X"CD",X"E3",X"20",X"DA",
		X"36",X"20",X"DD",X"35",X"07",X"C0",X"DD",X"35",X"0E",X"FA",X"85",X"20",X"28",X"54",X"DD",X"34",
		X"06",X"DD",X"36",X"07",X"05",X"3A",X"E6",X"E2",X"FE",X"02",X"C0",X"CD",X"D4",X"1D",X"ED",X"5B",
		X"0C",X"E8",X"21",X"60",X"FA",X"19",X"D8",X"21",X"00",X"FE",X"19",X"D0",X"2A",X"DA",X"E2",X"11",
		X"00",X"02",X"19",X"22",X"0F",X"E8",X"11",X"C0",X"02",X"19",X"22",X"11",X"E8",X"3A",X"DE",X"E2",
		X"FE",X"0B",X"38",X"0C",X"28",X"05",X"21",X"00",X"69",X"18",X"08",X"21",X"80",X"61",X"18",X"03",
		X"21",X"80",X"59",X"11",X"05",X"00",X"E5",X"CD",X"72",X"11",X"E1",X"D0",X"11",X"10",X"01",X"C3",
		X"95",X"2C",X"DD",X"35",X"0B",X"20",X"0B",X"DD",X"34",X"06",X"DD",X"36",X"07",X"05",X"C9",X"CD",
		X"E8",X"2C",X"3A",X"11",X"E0",X"21",X"9E",X"E1",X"06",X"04",X"BE",X"38",X"08",X"23",X"06",X"09",
		X"BE",X"38",X"02",X"06",X"0E",X"DD",X"70",X"06",X"DD",X"36",X"0E",X"04",X"3A",X"12",X"E0",X"21",
		X"A0",X"E1",X"CD",X"14",X"12",X"32",X"DF",X"E2",X"C9",X"CD",X"AA",X"1B",X"DD",X"CB",X"00",X"66",
		X"C0",X"E1",X"21",X"D8",X"E2",X"CB",X"A6",X"21",X"E8",X"E2",X"CB",X"A6",X"C9",X"DD",X"36",X"01",
		X"02",X"CD",X"E2",X"1B",X"DD",X"35",X"07",X"CA",X"CF",X"1F",X"C9",X"ED",X"5B",X"04",X"E1",X"DD",
		X"6E",X"02",X"DD",X"66",X"03",X"ED",X"52",X"38",X"E4",X"11",X"55",X"00",X"CD",X"7A",X"1C",X"18",
		X"E0",X"DD",X"36",X"01",X"06",X"C9",X"C6",X"13",X"32",X"DE",X"E2",X"FE",X"16",X"21",X"26",X"21",
		X"38",X"03",X"21",X"2C",X"21",X"CD",X"96",X"1B",X"21",X"67",X"2D",X"11",X"D8",X"00",X"CD",X"19",
		X"2D",X"3E",X"08",X"DA",X"7A",X"24",X"DD",X"7E",X"FE",X"DD",X"36",X"FE",X"1C",X"A7",X"20",X"D1",
		X"DD",X"34",X"01",X"C9",X"CD",X"13",X"2D",X"CD",X"E3",X"20",X"DA",X"36",X"20",X"ED",X"5B",X"04",
		X"E1",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"ED",X"52",X"38",X"05",X"DD",X"7E",X"08",X"A7",X"C0",
		X"DD",X"36",X"01",X"00",X"C9",X"DD",X"36",X"06",X"00",X"DD",X"36",X"07",X"07",X"DD",X"36",X"01",
		X"05",X"DD",X"36",X"08",X"25",X"C9",X"CD",X"B9",X"2C",X"CD",X"78",X"2C",X"21",X"8D",X"6C",X"11",
		X"A0",X"FE",X"3A",X"01",X"E7",X"E6",X"03",X"20",X"04",X"DD",X"CB",X"00",X"AE",X"E5",X"DD",X"7E",
		X"01",X"FE",X"01",X"28",X"1D",X"2A",X"0C",X"E8",X"19",X"21",X"01",X"E7",X"DD",X"CB",X"00",X"76",
		X"28",X"0A",X"38",X"04",X"CB",X"E6",X"18",X"11",X"CB",X"A6",X"18",X"0D",X"38",X"09",X"CB",X"EE",
		X"18",X"07",X"21",X"01",X"E7",X"CB",X"A6",X"CB",X"AE",X"E1",X"CD",X"01",X"2D",X"DD",X"7E",X"00",
		X"C3",X"7E",X"1A",X"CD",X"09",X"21",X"D0",X"2A",X"0C",X"E8",X"11",X"60",X"FE",X"19",X"D0",X"3A",
		X"DE",X"E2",X"FE",X"04",X"38",X"07",X"FE",X"09",X"21",X"12",X"21",X"38",X"03",X"21",X"1C",X"21",
		X"CD",X"18",X"1B",X"D0",X"DD",X"CB",X"00",X"EE",X"C9",X"DD",X"7E",X"00",X"E6",X"20",X"C0",X"C3",
		X"E7",X"1A",X"04",X"03",X"FF",X"FF",X"FF",X"FF",X"04",X"FF",X"FF",X"FF",X"02",X"00",X"02",X"02",
		X"02",X"02",X"01",X"FF",X"FF",X"FF",X"06",X"18",X"08",X"19",X"11",X"FF",X"06",X"1A",X"08",X"1B",
		X"11",X"FF",X"48",X"21",X"F9",X"1F",X"00",X"22",X"5D",X"21",X"67",X"21",X"17",X"22",X"21",X"39",
		X"22",X"E5",X"21",X"32",X"21",X"C3",X"23",X"1F",X"CD",X"0D",X"2D",X"11",X"00",X"FB",X"19",X"D2",
		X"DC",X"21",X"11",X"00",X"C0",X"2A",X"DA",X"E2",X"19",X"DA",X"50",X"1F",X"C9",X"CD",X"E2",X"1B",
		X"11",X"00",X"FB",X"19",X"30",X"76",X"C9",X"CD",X"E2",X"1B",X"CD",X"4B",X"22",X"DA",X"0A",X"22",
		X"DD",X"35",X"07",X"C0",X"DD",X"35",X"0E",X"28",X"5B",X"DD",X"34",X"06",X"DD",X"36",X"07",X"0B",
		X"3A",X"E6",X"E2",X"FE",X"02",X"C0",X"CD",X"D4",X"1D",X"2A",X"DA",X"E2",X"3A",X"DE",X"E2",X"FE",
		X"07",X"38",X"16",X"11",X"E0",X"01",X"19",X"22",X"0F",X"E8",X"11",X"20",X"02",X"19",X"22",X"11",
		X"E8",X"21",X"00",X"5E",X"11",X"11",X"00",X"18",X"14",X"11",X"40",X"02",X"19",X"22",X"0F",X"E8",
		X"11",X"E0",X"01",X"19",X"22",X"11",X"E8",X"21",X"00",X"6A",X"11",X"0A",X"00",X"CD",X"72",X"11",
		X"D0",X"3A",X"DE",X"E2",X"FE",X"07",X"21",X"80",X"6C",X"38",X"03",X"21",X"80",X"60",X"11",X"18",
		X"00",X"C3",X"95",X"2C",X"DD",X"35",X"0B",X"20",X"06",X"C3",X"20",X"22",X"CD",X"E8",X"2C",X"3A",
		X"11",X"E0",X"21",X"9E",X"E1",X"06",X"04",X"BE",X"38",X"02",X"06",X"07",X"DD",X"70",X"06",X"3A",
		X"12",X"E0",X"21",X"A5",X"E1",X"CD",X"14",X"12",X"32",X"DF",X"E2",X"DD",X"36",X"0E",X"03",X"C9",
		X"CD",X"E2",X"1B",X"DD",X"35",X"07",X"CA",X"50",X"1F",X"C9",X"DD",X"36",X"06",X"00",X"DD",X"36",
		X"07",X"0B",X"DD",X"36",X"01",X"02",X"C9",X"CD",X"13",X"2D",X"CD",X"4B",X"22",X"C3",X"6D",X"20",
		X"DD",X"36",X"06",X"00",X"DD",X"36",X"07",X"07",X"DD",X"36",X"01",X"05",X"3A",X"13",X"E0",X"21",
		X"A0",X"E1",X"CD",X"14",X"12",X"DD",X"77",X"08",X"C9",X"CD",X"B9",X"2C",X"CD",X"78",X"2C",X"21",
		X"65",X"6E",X"11",X"20",X"FE",X"CD",X"A2",X"20",X"C3",X"70",X"2E",X"3A",X"D8",X"E2",X"E6",X"20",
		X"C0",X"21",X"E0",X"00",X"CD",X"20",X"12",X"D0",X"DD",X"CB",X"00",X"EE",X"D5",X"21",X"05",X"00",
		X"CD",X"5C",X"2E",X"21",X"6A",X"2D",X"CD",X"19",X"2D",X"D1",X"38",X"05",X"21",X"00",X"90",X"19",
		X"C9",X"F1",X"11",X"EE",X"00",X"3E",X"09",X"CD",X"7A",X"24",X"DD",X"36",X"06",X"00",X"21",X"84",
		X"22",X"C3",X"96",X"1B",X"06",X"0A",X"08",X"0B",X"13",X"FF",X"A5",X"22",X"F9",X"1F",X"09",X"24",
		X"C7",X"22",X"D2",X"22",X"80",X"24",X"32",X"24",X"CD",X"6F",X"2C",X"21",X"9F",X"24",X"E5",X"21",
		X"8A",X"22",X"C3",X"23",X"1F",X"CD",X"0D",X"2D",X"11",X"00",X"F6",X"19",X"D2",X"C6",X"23",X"11",
		X"00",X"5F",X"2A",X"DA",X"E2",X"19",X"D2",X"50",X"1F",X"C9",X"DD",X"36",X"01",X"00",X"DD",X"36",
		X"06",X"00",X"DD",X"36",X"07",X"02",X"C9",X"CD",X"E2",X"1B",X"11",X"00",X"F6",X"19",X"D2",X"C6",
		X"23",X"C9",X"CD",X"E2",X"1B",X"CD",X"B0",X"24",X"DA",X"48",X"24",X"DD",X"35",X"07",X"C0",X"DD",
		X"35",X"0E",X"28",X"60",X"FA",X"B4",X"23",X"DD",X"34",X"06",X"DD",X"36",X"07",X"0B",X"FD",X"21",
		X"FB",X"E2",X"FD",X"CB",X"00",X"66",X"28",X"04",X"FD",X"21",X"0B",X"E3",X"3A",X"E7",X"E2",X"FE",
		X"02",X"21",X"00",X"69",X"38",X"03",X"21",X"80",X"56",X"FD",X"75",X"04",X"FD",X"74",X"05",X"FD",
		X"77",X"0B",X"2A",X"DA",X"E2",X"11",X"00",X"FF",X"19",X"FD",X"75",X"02",X"FD",X"74",X"03",X"11",
		X"00",X"ED",X"19",X"FD",X"75",X"0E",X"FD",X"74",X"0F",X"2A",X"B9",X"E1",X"FD",X"75",X"0C",X"FD",
		X"74",X"0D",X"3E",X"50",X"FD",X"77",X"00",X"AF",X"FD",X"77",X"01",X"FD",X"77",X"06",X"3E",X"02",
		X"FD",X"77",X"07",X"C9",X"DD",X"34",X"0E",X"DD",X"34",X"07",X"FD",X"21",X"FB",X"E2",X"FD",X"CB",
		X"00",X"66",X"28",X"14",X"FD",X"CB",X"0D",X"7E",X"C0",X"DD",X"CB",X"FF",X"46",X"28",X"12",X"FD",
		X"CB",X"10",X"66",X"20",X"0C",X"C3",X"D3",X"23",X"FD",X"21",X"0B",X"E3",X"FD",X"CB",X"0D",X"7E",
		X"C0",X"FD",X"7E",X"0B",X"A7",X"28",X"08",X"FE",X"03",X"28",X"04",X"3E",X"0A",X"18",X"02",X"3E",
		X"0C",X"DD",X"77",X"06",X"2A",X"DA",X"E2",X"11",X"C0",X"FE",X"19",X"FD",X"5E",X"02",X"FD",X"56",
		X"03",X"ED",X"52",X"D0",X"FD",X"36",X"00",X"00",X"DD",X"35",X"06",X"3A",X"0B",X"E3",X"E6",X"10",
		X"3E",X"0B",X"20",X"0C",X"DD",X"35",X"0E",X"3A",X"11",X"E0",X"21",X"A5",X"E1",X"CD",X"14",X"12",
		X"32",X"DF",X"E2",X"C9",X"2A",X"0C",X"E8",X"11",X"00",X"F5",X"19",X"DA",X"BA",X"22",X"DD",X"35",
		X"0B",X"20",X"09",X"C3",X"20",X"22",X"3A",X"9F",X"E1",X"32",X"E3",X"E2",X"ED",X"5F",X"E6",X"01",
		X"DD",X"77",X"FF",X"DD",X"36",X"01",X"04",X"3A",X"10",X"E0",X"21",X"9C",X"E1",X"06",X"00",X"BE",
		X"38",X"0B",X"23",X"04",X"BE",X"38",X"06",X"23",X"04",X"BE",X"38",X"01",X"04",X"DD",X"70",X"0F",
		X"78",X"06",X"09",X"FE",X"02",X"30",X"02",X"06",X"0B",X"DD",X"70",X"06",X"DD",X"36",X"07",X"0B",
		X"DD",X"36",X"0E",X"02",X"C9",X"DD",X"36",X"01",X"02",X"CD",X"E2",X"1B",X"DD",X"35",X"07",X"C0",
		X"DD",X"34",X"07",X"3A",X"0B",X"E3",X"E6",X"10",X"20",X"0D",X"3A",X"FB",X"E2",X"E6",X"10",X"28",
		X"A5",X"DD",X"CB",X"FF",X"46",X"20",X"AC",X"3A",X"E4",X"E2",X"32",X"DE",X"E2",X"DD",X"36",X"01",
		X"04",X"C9",X"ED",X"5B",X"06",X"E1",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"ED",X"52",X"30",X"C5",
		X"11",X"55",X"00",X"CD",X"7A",X"1C",X"18",X"C1",X"DD",X"46",X"06",X"C6",X"04",X"32",X"DE",X"E2",
		X"21",X"6D",X"2D",X"CD",X"19",X"2D",X"38",X"17",X"DD",X"70",X"0C",X"DD",X"36",X"07",X"06",X"DD",
		X"7E",X"FE",X"DD",X"36",X"FE",X"1C",X"A7",X"C2",X"31",X"20",X"DD",X"36",X"01",X"02",X"C9",X"21",
		X"CC",X"24",X"CD",X"96",X"1B",X"11",X"DC",X"00",X"3E",X"09",X"2A",X"DA",X"E2",X"C3",X"60",X"2F",
		X"CD",X"13",X"2D",X"CD",X"B0",X"24",X"38",X"C0",X"ED",X"5B",X"06",X"E1",X"DD",X"6E",X"02",X"DD",
		X"66",X"03",X"ED",X"52",X"D2",X"80",X"20",X"DD",X"7E",X"08",X"A7",X"CA",X"80",X"20",X"C9",X"21",
		X"00",X"E7",X"CB",X"F6",X"CD",X"B9",X"2C",X"CD",X"78",X"2C",X"21",X"4E",X"6F",X"C3",X"9F",X"20",
		X"CD",X"09",X"21",X"D0",X"2A",X"0C",X"E8",X"11",X"60",X"FE",X"19",X"D0",X"21",X"C2",X"24",X"C3",
		X"00",X"21",X"02",X"00",X"02",X"02",X"02",X"02",X"01",X"FF",X"FF",X"FF",X"06",X"07",X"08",X"08",
		X"11",X"FF",X"18",X"25",X"F9",X"1F",X"C3",X"25",X"35",X"25",X"40",X"25",X"1B",X"27",X"7F",X"26",
		X"D6",X"26",X"E2",X"1B",X"03",X"28",X"BA",X"27",X"37",X"27",X"84",X"27",X"E3",X"25",X"2F",X"26",
		X"2A",X"F8",X"E2",X"7D",X"B4",X"28",X"04",X"2B",X"22",X"F8",X"E2",X"21",X"D6",X"E2",X"7E",X"A7",
		X"28",X"01",X"35",X"CD",X"0F",X"25",X"DD",X"21",X"E8",X"E2",X"DD",X"CB",X"00",X"66",X"C8",X"21",
		X"D2",X"24",X"CD",X"23",X"1F",X"C3",X"93",X"28",X"CD",X"0D",X"2D",X"11",X"00",X"F8",X"19",X"D2",
		X"89",X"25",X"DD",X"CB",X"00",X"76",X"C0",X"11",X"00",X"5F",X"DD",X"6E",X"02",X"DD",X"66",X"03",
		X"19",X"D2",X"50",X"1F",X"C9",X"CD",X"E2",X"1B",X"11",X"00",X"F8",X"19",X"D2",X"89",X"25",X"C9",
		X"CD",X"E2",X"1B",X"CD",X"BA",X"28",X"DA",X"4B",X"26",X"DD",X"7E",X"0E",X"A7",X"FC",X"AF",X"25",
		X"DD",X"35",X"07",X"C0",X"A7",X"28",X"15",X"FA",X"8C",X"25",X"DD",X"86",X"06",X"DD",X"77",X"06",
		X"CD",X"DD",X"34",X"DD",X"36",X"07",X"0B",X"DD",X"36",X"0E",X"00",X"C9",X"DD",X"35",X"0B",X"CA",
		X"20",X"22",X"CD",X"AF",X"25",X"DD",X"36",X"06",X"00",X"DD",X"35",X"0E",X"3A",X"11",X"E0",X"21",
		X"A5",X"E1",X"CD",X"14",X"12",X"DD",X"77",X"07",X"C9",X"CD",X"E8",X"2C",X"CD",X"D4",X"2C",X"CA",
		X"DF",X"27",X"3A",X"12",X"E0",X"21",X"9E",X"E1",X"06",X"01",X"BE",X"38",X"06",X"04",X"23",X"BE",
		X"38",X"01",X"04",X"DD",X"70",X"0E",X"DD",X"36",X"06",X"04",X"DD",X"36",X"07",X"0B",X"C9",X"2A",
		X"0C",X"E8",X"11",X"80",X"F3",X"19",X"D0",X"F1",X"DD",X"36",X"06",X"00",X"DD",X"36",X"07",X"07",
		X"C3",X"80",X"20",X"CD",X"E2",X"1B",X"DD",X"35",X"07",X"C0",X"3A",X"D7",X"E2",X"A7",X"CA",X"50",
		X"1F",X"DD",X"36",X"01",X"0D",X"DD",X"36",X"06",X"1A",X"DD",X"36",X"07",X"08",X"21",X"00",X"E7",
		X"CB",X"C6",X"C9",X"CD",X"E2",X"1B",X"DD",X"35",X"07",X"C0",X"DD",X"36",X"07",X"08",X"DD",X"34",
		X"06",X"DD",X"7E",X"06",X"FE",X"22",X"C0",X"DD",X"34",X"01",X"DD",X"36",X"06",X"1E",X"DD",X"6E",
		X"02",X"DD",X"66",X"03",X"DD",X"CB",X"00",X"76",X"28",X"0E",X"11",X"00",X"A1",X"ED",X"52",X"19",
		X"38",X"14",X"11",X"80",X"FD",X"19",X"18",X"0E",X"11",X"80",X"02",X"19",X"ED",X"5B",X"06",X"E1",
		X"ED",X"52",X"19",X"38",X"01",X"EB",X"DD",X"75",X"02",X"DD",X"74",X"03",X"C3",X"E2",X"1B",X"CD",
		X"E2",X"1B",X"DD",X"35",X"07",X"C0",X"DD",X"36",X"07",X"08",X"DD",X"34",X"06",X"DD",X"7E",X"06",
		X"FE",X"26",X"C0",X"21",X"00",X"E7",X"CB",X"86",X"C3",X"50",X"1F",X"A7",X"28",X"4A",X"DD",X"36",
		X"06",X"08",X"21",X"70",X"2D",X"CD",X"19",X"2D",X"21",X"D6",X"28",X"38",X"11",X"7E",X"DD",X"77",
		X"07",X"DD",X"36",X"01",X"02",X"21",X"D6",X"E2",X"7E",X"36",X"1C",X"23",X"77",X"C9",X"CD",X"96",
		X"1B",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"11",X"D7",X"00",X"3E",X"0A",X"C3",X"60",X"2F",X"CD",
		X"E2",X"1B",X"DD",X"35",X"07",X"C0",X"DD",X"7E",X"06",X"3C",X"FE",X"13",X"38",X"40",X"20",X"5D",
		X"DD",X"36",X"07",X"1C",X"3E",X"26",X"18",X"3A",X"3E",X"91",X"CD",X"FE",X"0D",X"DD",X"6E",X"02",
		X"DD",X"66",X"03",X"22",X"1D",X"E3",X"DD",X"7E",X"00",X"E6",X"50",X"32",X"1B",X"E3",X"21",X"00",
		X"65",X"22",X"1F",X"E3",X"21",X"5B",X"00",X"22",X"27",X"E3",X"3E",X"05",X"32",X"22",X"E3",X"AF",
		X"32",X"21",X"E3",X"21",X"00",X"E7",X"CB",X"C6",X"DD",X"36",X"01",X"06",X"3E",X"0B",X"DD",X"36",
		X"07",X"08",X"DD",X"77",X"06",X"C9",X"CD",X"E2",X"1B",X"DD",X"35",X"07",X"C0",X"DD",X"7E",X"06",
		X"3C",X"FE",X"1A",X"38",X"E9",X"21",X"00",X"E7",X"CB",X"86",X"C3",X"89",X"25",X"DD",X"34",X"01",
		X"DD",X"6E",X"02",X"DD",X"66",X"03",X"11",X"80",X"02",X"DD",X"CB",X"00",X"76",X"20",X"0D",X"19",
		X"EB",X"2A",X"06",X"E1",X"ED",X"52",X"19",X"38",X"05",X"EB",X"18",X"02",X"ED",X"52",X"DD",X"75",
		X"02",X"DD",X"74",X"03",X"CD",X"E2",X"1B",X"3E",X"0F",X"18",X"B3",X"CD",X"13",X"2D",X"CD",X"BA",
		X"28",X"DA",X"4B",X"26",X"CD",X"D4",X"2C",X"CA",X"80",X"20",X"DD",X"CB",X"00",X"76",X"CA",X"88",
		X"24",X"11",X"00",X"A1",X"C3",X"71",X"20",X"DD",X"35",X"07",X"20",X"16",X"DD",X"34",X"07",X"CD",
		X"87",X"28",X"20",X"6C",X"DD",X"36",X"07",X"07",X"DD",X"35",X"06",X"F2",X"52",X"27",X"DD",X"36",
		X"06",X"03",X"2A",X"12",X"E7",X"DD",X"5E",X"0C",X"DD",X"56",X"0D",X"ED",X"52",X"EB",X"DD",X"CB",
		X"00",X"76",X"20",X"0D",X"2A",X"06",X"E1",X"ED",X"52",X"30",X"04",X"ED",X"5B",X"06",X"E1",X"18",
		X"0A",X"21",X"80",X"85",X"ED",X"52",X"38",X"03",X"11",X"80",X"85",X"DD",X"73",X"02",X"DD",X"72",
		X"03",X"C3",X"E2",X"1B",X"CD",X"E2",X"1B",X"CD",X"87",X"28",X"28",X"17",X"DD",X"35",X"07",X"C0",
		X"DD",X"7E",X"0E",X"A7",X"CA",X"75",X"25",X"FA",X"92",X"25",X"DD",X"86",X"06",X"DD",X"77",X"06",
		X"C3",X"63",X"25",X"DD",X"36",X"06",X"00",X"DD",X"36",X"07",X"02",X"DD",X"36",X"01",X"0B",X"C9",
		X"DD",X"36",X"01",X"0C",X"CD",X"92",X"25",X"C3",X"E2",X"1B",X"CD",X"E2",X"1B",X"DD",X"35",X"07",
		X"C0",X"DD",X"36",X"07",X"08",X"DD",X"34",X"06",X"DD",X"7E",X"06",X"FE",X"22",X"C0",X"21",X"8B",
		X"01",X"22",X"F8",X"E2",X"DD",X"36",X"00",X"00",X"21",X"01",X"E7",X"CB",X"A6",X"18",X"5E",X"21",
		X"00",X"E7",X"CB",X"C6",X"3A",X"E8",X"E2",X"E6",X"10",X"28",X"64",X"DD",X"E5",X"DD",X"21",X"D8",
		X"E2",X"CD",X"7E",X"28",X"DD",X"36",X"17",X"08",X"DD",X"36",X"16",X"1A",X"DD",X"36",X"11",X"0A",
		X"DD",X"E1",X"C9",X"CD",X"E2",X"1B",X"DD",X"35",X"07",X"C0",X"DD",X"36",X"07",X"08",X"DD",X"34",
		X"06",X"DD",X"7E",X"06",X"FE",X"26",X"C0",X"21",X"1A",X"01",X"22",X"F8",X"E2",X"CD",X"A3",X"27",
		X"CD",X"3D",X"28",X"ED",X"5F",X"E6",X"01",X"C8",X"DD",X"36",X"F1",X"0B",X"DD",X"36",X"01",X"00",
		X"21",X"00",X"00",X"ED",X"5B",X"F4",X"E2",X"ED",X"52",X"22",X"E4",X"E2",X"C9",X"DD",X"36",X"F6",
		X"00",X"DD",X"36",X"F7",X"02",X"DD",X"36",X"F1",X"00",X"21",X"00",X"E7",X"CB",X"86",X"C9",X"ED",
		X"5B",X"0A",X"E8",X"21",X"60",X"FD",X"19",X"38",X"03",X"11",X"A0",X"02",X"2A",X"12",X"E7",X"ED",
		X"53",X"F4",X"E2",X"ED",X"52",X"22",X"EA",X"E2",X"21",X"00",X"50",X"22",X"EC",X"E2",X"DD",X"36",
		X"10",X"50",X"DD",X"36",X"17",X"08",X"DD",X"36",X"16",X"1E",X"DD",X"36",X"11",X"09",X"DD",X"36",
		X"01",X"08",X"DD",X"36",X"06",X"1A",X"C9",X"3A",X"02",X"E7",X"FE",X"01",X"C8",X"FE",X"09",X"C8",
		X"FE",X"0A",X"C9",X"2A",X"0C",X"E8",X"11",X"00",X"E8",X"19",X"21",X"97",X"E1",X"11",X"98",X"E1",
		X"30",X"08",X"3A",X"E8",X"E2",X"E6",X"10",X"20",X"01",X"EB",X"7E",X"A7",X"28",X"03",X"12",X"36",
		X"00",X"21",X"47",X"70",X"11",X"00",X"FE",X"C3",X"AD",X"20",X"CD",X"E7",X"1A",X"D0",X"2A",X"0C",
		X"E8",X"11",X"60",X"FE",X"19",X"D0",X"21",X"CC",X"28",X"C3",X"18",X"1B",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"01",X"FF",X"FF",X"FF",X"06",X"09",X"08",X"0A",X"13",X"FF",X"FC",X"28",X"F9",X"1F",
		X"EE",X"2A",X"56",X"29",X"CC",X"29",X"8C",X"2A",X"14",X"29",X"8F",X"29",X"C8",X"2A",X"28",X"2B",
		X"32",X"2B",X"21",X"5A",X"2C",X"E5",X"21",X"DC",X"28",X"C3",X"23",X"1F",X"CD",X"0D",X"2D",X"11",
		X"60",X"F7",X"19",X"30",X"2A",X"18",X"1C",X"DD",X"36",X"07",X"07",X"DD",X"36",X"01",X"00",X"DD",
		X"36",X"06",X"00",X"C9",X"CD",X"3C",X"29",X"CD",X"70",X"1C",X"CD",X"E2",X"1B",X"11",X"60",X"F7",
		X"19",X"38",X"E4",X"11",X"00",X"C0",X"2A",X"DA",X"E2",X"19",X"DA",X"50",X"1F",X"18",X"36",X"DD",
		X"36",X"07",X"09",X"DD",X"36",X"06",X"04",X"DD",X"36",X"01",X"06",X"C9",X"DD",X"35",X"07",X"20",
		X"11",X"DD",X"36",X"07",X"09",X"DD",X"7E",X"06",X"3C",X"FE",X"05",X"28",X"02",X"3E",X"04",X"DD",
		X"77",X"06",X"11",X"12",X"00",X"C9",X"CD",X"E2",X"1B",X"11",X"60",X"F7",X"19",X"3E",X"04",X"30",
		X"01",X"AF",X"DD",X"77",X"06",X"CD",X"A0",X"2B",X"2A",X"0C",X"E8",X"11",X"80",X"FB",X"19",X"D8",
		X"DD",X"7E",X"08",X"A7",X"C2",X"E9",X"2A",X"DD",X"36",X"06",X"04",X"2A",X"0C",X"E8",X"11",X"00",
		X"FD",X"19",X"30",X"1C",X"3A",X"AA",X"E1",X"DD",X"77",X"07",X"DD",X"36",X"01",X"07",X"C9",X"ED",
		X"5B",X"AB",X"E1",X"CD",X"70",X"1C",X"CD",X"E2",X"1B",X"CD",X"A0",X"2B",X"DD",X"35",X"07",X"C0",
		X"CD",X"E8",X"2C",X"2A",X"0C",X"E8",X"11",X"80",X"FC",X"19",X"DA",X"55",X"2A",X"3A",X"11",X"E0",
		X"21",X"9E",X"E1",X"06",X"06",X"BE",X"38",X"08",X"23",X"06",X"0B",X"BE",X"38",X"02",X"06",X"10",
		X"DD",X"70",X"06",X"DD",X"36",X"07",X"05",X"DD",X"36",X"0E",X"05",X"C9",X"CD",X"E2",X"1B",X"CD",
		X"A0",X"2B",X"DD",X"35",X"07",X"C0",X"DD",X"35",X"0E",X"28",X"62",X"FA",X"A3",X"29",X"DD",X"7E",
		X"0E",X"FE",X"03",X"20",X"47",X"DD",X"7E",X"06",X"FE",X"0C",X"21",X"73",X"2A",X"38",X"08",X"21",
		X"7A",X"2A",X"28",X"03",X"21",X"81",X"2A",X"DD",X"7E",X"02",X"86",X"23",X"5F",X"DD",X"7E",X"03",
		X"8E",X"23",X"57",X"ED",X"53",X"0F",X"E8",X"7B",X"86",X"23",X"5F",X"7A",X"8E",X"23",X"57",X"ED",
		X"53",X"11",X"E8",X"5E",X"23",X"56",X"23",X"6E",X"26",X"00",X"EB",X"E5",X"CD",X"72",X"11",X"E1",
		X"30",X"0A",X"11",X"00",X"04",X"19",X"11",X"18",X"00",X"CD",X"95",X"2C",X"DD",X"34",X"06",X"DD",
		X"5E",X"0E",X"16",X"00",X"21",X"87",X"2A",X"19",X"7E",X"DD",X"77",X"07",X"C9",X"DD",X"35",X"0B",
		X"28",X"13",X"3A",X"12",X"E0",X"21",X"A5",X"E1",X"CD",X"14",X"12",X"DD",X"77",X"07",X"C9",X"21",
		X"00",X"50",X"22",X"DC",X"E2",X"DD",X"36",X"06",X"04",X"2A",X"DA",X"E2",X"11",X"00",X"FE",X"19",
		X"ED",X"5B",X"04",X"E1",X"ED",X"52",X"38",X"71",X"DD",X"36",X"01",X"08",X"3A",X"AA",X"E1",X"DD",
		X"77",X"07",X"C9",X"20",X"01",X"60",X"01",X"80",X"67",X"07",X"40",X"01",X"20",X"02",X"00",X"66",
		X"0E",X"80",X"01",X"00",X"02",X"00",X"50",X"0A",X"01",X"10",X"0B",X"10",X"CD",X"3C",X"29",X"CD",
		X"7A",X"1C",X"CD",X"B6",X"2A",X"CD",X"A0",X"2B",X"DD",X"7E",X"08",X"A7",X"CA",X"77",X"29",X"2A",
		X"0C",X"E8",X"11",X"00",X"FB",X"19",X"DA",X"37",X"29",X"2A",X"DA",X"E2",X"ED",X"5B",X"04",X"E1",
		X"ED",X"52",X"DA",X"77",X"29",X"C9",X"2A",X"DA",X"E2",X"ED",X"5B",X"04",X"E1",X"ED",X"52",X"30",
		X"04",X"ED",X"53",X"DA",X"E2",X"C3",X"E2",X"1B",X"ED",X"5B",X"AB",X"E1",X"CD",X"7A",X"1C",X"CD",
		X"B6",X"2A",X"CD",X"A0",X"2B",X"DD",X"35",X"07",X"C0",X"3A",X"12",X"E0",X"21",X"A0",X"E1",X"CD",
		X"14",X"12",X"DD",X"77",X"08",X"DD",X"36",X"07",X"09",X"DD",X"36",X"01",X"05",X"C9",X"CD",X"E2",
		X"1B",X"DD",X"35",X"07",X"CA",X"4F",X"2A",X"C9",X"E1",X"78",X"FE",X"02",X"3E",X"1B",X"38",X"04",
		X"28",X"01",X"3D",X"3D",X"DD",X"77",X"06",X"78",X"FE",X"03",X"28",X"04",X"AF",X"32",X"D6",X"E2",
		X"21",X"69",X"2C",X"CD",X"96",X"1B",X"21",X"67",X"2D",X"11",X"DE",X"00",X"CD",X"19",X"2D",X"3E",
		X"0B",X"DA",X"7A",X"24",X"DD",X"34",X"01",X"C9",X"CD",X"E2",X"1B",X"DD",X"35",X"07",X"CA",X"55",
		X"2A",X"C9",X"CD",X"E2",X"1B",X"21",X"D7",X"E2",X"7E",X"A7",X"20",X"12",X"3A",X"DE",X"E2",X"FE",
		X"1E",X"20",X"0B",X"36",X"01",X"21",X"00",X"60",X"11",X"18",X"00",X"CD",X"95",X"2C",X"2A",X"E4",
		X"E2",X"DD",X"35",X"07",X"20",X"14",X"23",X"23",X"7E",X"FE",X"FF",X"CA",X"4F",X"2A",X"DD",X"77",
		X"06",X"23",X"7E",X"DD",X"77",X"07",X"23",X"22",X"E4",X"E2",X"7E",X"DD",X"86",X"04",X"DD",X"77",
		X"04",X"23",X"7E",X"DD",X"8E",X"05",X"DD",X"77",X"05",X"C9",X"20",X"01",X"18",X"03",X"AA",X"00",
		X"18",X"02",X"00",X"00",X"18",X"03",X"56",X"FF",X"17",X"04",X"E0",X"FE",X"FF",X"20",X"01",X"1E",
		X"03",X"AA",X"00",X"1E",X"02",X"00",X"00",X"1E",X"03",X"56",X"FF",X"17",X"04",X"E0",X"FE",X"FF",
		X"CD",X"E7",X"1A",X"D0",X"21",X"36",X"2C",X"CD",X"18",X"1B",X"D0",X"47",X"DD",X"5E",X"06",X"16",
		X"00",X"21",X"40",X"2C",X"19",X"7E",X"FE",X"FF",X"C8",X"21",X"D6",X"E2",X"34",X"FE",X"FE",X"28",
		X"1C",X"FE",X"08",X"38",X"0B",X"5F",X"78",X"FE",X"02",X"38",X"62",X"7B",X"FE",X"09",X"28",X"0D",
		X"80",X"5F",X"21",X"AD",X"E1",X"19",X"3A",X"13",X"E0",X"BE",X"D2",X"F8",X"2A",X"E1",X"78",X"FE",
		X"02",X"28",X"38",X"38",X"32",X"DD",X"36",X"07",X"05",X"DD",X"36",X"01",X"0A",X"DD",X"36",X"06",
		X"17",X"3A",X"80",X"E0",X"0F",X"0F",X"0F",X"E6",X"03",X"5F",X"16",X"00",X"21",X"32",X"2C",X"19",
		X"3A",X"D6",X"E2",X"BE",X"21",X"7A",X"2B",X"38",X"0A",X"21",X"8D",X"2B",X"AF",X"32",X"D7",X"E2",
		X"32",X"D6",X"E2",X"22",X"E4",X"E2",X"C9",X"3E",X"15",X"18",X"02",X"3E",X"16",X"DD",X"77",X"06",
		X"DD",X"36",X"01",X"09",X"DD",X"36",X"07",X"0B",X"3E",X"91",X"CD",X"FE",X"0D",X"AF",X"32",X"D6",
		X"E2",X"C9",X"04",X"03",X"02",X"02",X"00",X"03",X"00",X"00",X"00",X"01",X"02",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"00",X"00",X"00",X"FE",X"FE",X"04",X"04",X"04",X"FE",
		X"09",X"08",X"08",X"08",X"09",X"FF",X"FF",X"FF",X"FF",X"FF",X"CD",X"B9",X"2C",X"CD",X"7E",X"2C",
		X"11",X"00",X"FE",X"21",X"FA",X"71",X"C3",X"AD",X"20",X"0B",X"1C",X"08",X"1D",X"13",X"FF",X"DD",
		X"7E",X"FE",X"A7",X"C8",X"DD",X"35",X"FE",X"C9",X"3A",X"80",X"E0",X"E6",X"FC",X"C0",X"2A",X"0C",
		X"E8",X"11",X"00",X"E8",X"19",X"21",X"98",X"E1",X"11",X"97",X"E1",X"38",X"01",X"EB",X"7E",X"A7",
		X"C8",X"12",X"36",X"00",X"C9",X"3E",X"91",X"CD",X"FE",X"0D",X"3A",X"09",X"E7",X"93",X"F2",X"B6",
		X"2C",X"CD",X"08",X"12",X"20",X"10",X"3A",X"80",X"E0",X"E6",X"07",X"FE",X"02",X"3E",X"04",X"20",
		X"02",X"3E",X"05",X"32",X"07",X"E0",X"C3",X"E2",X"2E",X"2A",X"0C",X"E8",X"11",X"60",X"F7",X"19",
		X"21",X"00",X"E7",X"CB",X"A6",X"D8",X"DD",X"7E",X"01",X"FE",X"01",X"C8",X"3A",X"61",X"E2",X"A7",
		X"C0",X"CB",X"E6",X"C9",X"2A",X"F8",X"E2",X"7D",X"B4",X"C0",X"3A",X"02",X"E7",X"FE",X"09",X"28",
		X"05",X"FE",X"0A",X"28",X"01",X"7C",X"A7",X"C9",X"3A",X"10",X"E0",X"21",X"9C",X"E1",X"06",X"01",
		X"BE",X"38",X"06",X"23",X"04",X"BE",X"38",X"01",X"04",X"DD",X"70",X"0B",X"DD",X"36",X"01",X"04",
		X"C9",X"E5",X"2A",X"0C",X"E8",X"11",X"00",X"EE",X"19",X"E1",X"D0",X"F1",X"C9",X"11",X"1B",X"00",
		X"C3",X"EA",X"1B",X"11",X"1B",X"00",X"C3",X"F2",X"1B",X"3E",X"83",X"CD",X"FE",X"0D",X"3E",X"91",
		X"CD",X"FE",X"0D",X"D5",X"3A",X"06",X"E7",X"E5",X"21",X"42",X"2D",X"5F",X"16",X"00",X"19",X"5E",
		X"E1",X"19",X"3A",X"E2",X"E2",X"96",X"32",X"E2",X"E2",X"D1",X"D0",X"3E",X"87",X"CD",X"FE",X"0D",
		X"37",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"01",X"01",X"00",X"02",X"00",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"03",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"0C",X"20",X"0C",X"08",X"18",X"10",X"10",
		X"20",X"10",X"21",X"2B",X"E3",X"7E",X"A7",X"C8",X"47",X"23",X"C5",X"4E",X"11",X"B4",X"00",X"CB",
		X"49",X"28",X"03",X"11",X"D2",X"00",X"CB",X"61",X"28",X"07",X"E5",X"21",X"18",X"00",X"19",X"EB",
		X"E1",X"ED",X"53",X"07",X"E8",X"23",X"5E",X"E5",X"23",X"56",X"3A",X"00",X"E7",X"2A",X"F7",X"E1",
		X"CB",X"71",X"28",X"1A",X"EB",X"CB",X"4F",X"20",X"01",X"19",X"E5",X"ED",X"5B",X"12",X"E7",X"ED",
		X"52",X"22",X"0A",X"E8",X"38",X"26",X"11",X"00",X"F0",X"19",X"38",X"5E",X"18",X"1B",X"EB",X"CB",
		X"4F",X"20",X"02",X"ED",X"52",X"E5",X"38",X"52",X"ED",X"5B",X"12",X"E7",X"ED",X"52",X"22",X"0A",
		X"E8",X"30",X"09",X"11",X"00",X"10",X"19",X"30",X"41",X"2A",X"0A",X"E8",X"CB",X"4F",X"20",X"10",
		X"CB",X"61",X"20",X"0C",X"11",X"60",X"00",X"19",X"11",X"C0",X"00",X"ED",X"52",X"DC",X"31",X"2E",
		X"2A",X"0A",X"E8",X"16",X"FF",X"29",X"38",X"02",X"16",X"00",X"29",X"29",X"5C",X"2A",X"15",X"E7",
		X"19",X"EB",X"21",X"A0",X"75",X"79",X"EE",X"40",X"E6",X"40",X"CD",X"20",X"0E",X"D1",X"E1",X"73",
		X"23",X"72",X"23",X"C1",X"05",X"C2",X"7A",X"2D",X"C9",X"E1",X"21",X"2B",X"E3",X"7E",X"35",X"87",
		X"86",X"23",X"16",X"00",X"5F",X"19",X"D1",X"D1",X"13",X"01",X"03",X"00",X"ED",X"B8",X"EB",X"18",
		X"E1",X"CB",X"49",X"20",X"0D",X"2A",X"10",X"E7",X"11",X"00",X"A6",X"19",X"D8",X"21",X"00",X"5A",
		X"18",X"12",X"3A",X"02",X"E7",X"FE",X"06",X"C8",X"FE",X"07",X"C8",X"3A",X"06",X"E7",X"FE",X"05",
		X"C8",X"21",X"00",X"69",X"11",X"18",X"01",X"CD",X"E2",X"2E",X"18",X"BD",X"22",X"38",X"E3",X"EB",
		X"29",X"6C",X"26",X"00",X"30",X"01",X"24",X"22",X"36",X"E3",X"3E",X"07",X"32",X"35",X"E3",X"C9",
		X"21",X"35",X"E3",X"7E",X"A7",X"C8",X"35",X"C8",X"2A",X"36",X"E3",X"C5",X"22",X"07",X"E8",X"2A",
		X"38",X"E3",X"ED",X"5B",X"03",X"E8",X"19",X"EB",X"AF",X"21",X"84",X"74",X"CD",X"20",X"0E",X"C1",
		X"C9",X"3A",X"20",X"E7",X"FE",X"03",X"3E",X"01",X"28",X"01",X"AF",X"32",X"3F",X"E3",X"3A",X"01",
		X"E7",X"CB",X"77",X"21",X"FE",X"FF",X"28",X"03",X"21",X"02",X"00",X"22",X"3D",X"E3",X"2A",X"22",
		X"E7",X"29",X"6C",X"26",X"00",X"30",X"01",X"24",X"22",X"3B",X"E3",X"3E",X"0E",X"32",X"3A",X"E3",
		X"C9",X"21",X"3A",X"E3",X"7E",X"A7",X"C8",X"35",X"C8",X"2A",X"3B",X"E3",X"C5",X"22",X"07",X"E8",
		X"2A",X"3D",X"E3",X"ED",X"5B",X"15",X"E7",X"19",X"EB",X"AF",X"21",X"89",X"74",X"CD",X"20",X"0E",
		X"C1",X"C9",X"3A",X"1F",X"E7",X"E6",X"01",X"20",X"12",X"22",X"22",X"E7",X"21",X"1F",X"E7",X"CB",
		X"C6",X"23",X"72",X"23",X"73",X"3E",X"83",X"CD",X"FE",X"0D",X"C9",X"3A",X"09",X"E7",X"93",X"30",
		X"01",X"AF",X"32",X"09",X"E7",X"C9",X"21",X"4C",X"E6",X"06",X"04",X"7E",X"A7",X"C8",X"35",X"28",
		X"35",X"C5",X"23",X"5E",X"23",X"56",X"ED",X"53",X"07",X"E8",X"23",X"5E",X"23",X"56",X"23",X"4E",
		X"23",X"E5",X"2A",X"12",X"E7",X"7D",X"E6",X"E0",X"6F",X"EB",X"ED",X"52",X"E5",X"11",X"00",X"1C",
		X"38",X"04",X"ED",X"52",X"18",X"01",X"19",X"E1",X"30",X"07",X"11",X"F7",X"75",X"AF",X"CD",X"9A",
		X"1A",X"E1",X"C1",X"10",X"C6",X"C9",X"05",X"28",X"14",X"C5",X"E5",X"EB",X"21",X"06",X"00",X"19",
		X"78",X"87",X"80",X"87",X"4F",X"06",X"00",X"ED",X"B0",X"AF",X"12",X"18",X"E4",X"36",X"00",X"C9",
		X"C5",X"D5",X"E5",X"11",X"63",X"E6",X"21",X"5D",X"E6",X"01",X"12",X"00",X"ED",X"B8",X"57",X"E6",
		X"7F",X"5F",X"32",X"51",X"E6",X"E1",X"22",X"4F",X"E6",X"E1",X"22",X"4D",X"E6",X"3E",X"A9",X"CB",
		X"7A",X"28",X"02",X"3E",X"0B",X"32",X"4C",X"E6",X"16",X"00",X"21",X"AD",X"2F",X"19",X"19",X"5E",
		X"23",X"56",X"CD",X"9A",X"2F",X"C1",X"C9",X"11",X"10",X"00",X"21",X"81",X"E0",X"7E",X"83",X"27",
		X"77",X"23",X"7E",X"8A",X"27",X"77",X"23",X"7E",X"CE",X"00",X"27",X"77",X"C9",X"20",X"00",X"30",
		X"00",X"40",X"00",X"50",X"00",X"60",X"00",X"80",X"00",X"90",X"00",X"00",X"01",X"00",X"02",X"00",
		X"03",X"00",X"05",X"00",X"10",X"10",X"00",X"3A",X"81",X"E3",X"A7",X"C8",X"DD",X"21",X"82",X"E3",
		X"06",X"10",X"C5",X"DD",X"4E",X"00",X"CB",X"61",X"C4",X"E4",X"2F",X"C1",X"11",X"13",X"00",X"DD",
		X"19",X"10",X"EF",X"C9",X"21",X"E7",X"36",X"E5",X"21",X"F7",X"2F",X"DD",X"5E",X"01",X"16",X"00",
		X"19",X"19",X"7E",X"23",X"66",X"6F",X"E9",X"7F",X"33",X"D4",X"31",X"19",X"30",X"98",X"33",X"D4",
		X"33",X"C8",X"32",X"49",X"30",X"EE",X"31",X"25",X"32",X"8B",X"32",X"54",X"31",X"5D",X"31",X"66",
		X"31",X"44",X"34",X"78",X"34",X"84",X"34",X"37",X"35",X"CD",X"E2",X"1B",X"21",X"00",X"70",X"CD",
		X"1D",X"37",X"DA",X"CD",X"30",X"CD",X"73",X"37",X"DA",X"1E",X"33",X"CD",X"46",X"37",X"3E",X"91",
		X"DA",X"27",X"33",X"DD",X"35",X"07",X"C0",X"DD",X"36",X"07",X"03",X"DD",X"7E",X"06",X"3C",X"FE",
		X"04",X"20",X"02",X"3E",X"02",X"DD",X"77",X"06",X"C9",X"CD",X"E2",X"1B",X"DD",X"35",X"08",X"CA",
		X"06",X"31",X"DD",X"6E",X"0E",X"DD",X"66",X"0F",X"11",X"20",X"00",X"DD",X"CB",X"00",X"56",X"28",
		X"0D",X"ED",X"52",X"30",X"16",X"DD",X"CB",X"00",X"96",X"21",X"00",X"00",X"18",X"0D",X"19",X"E5",
		X"11",X"80",X"FF",X"19",X"E1",X"30",X"04",X"DD",X"CB",X"00",X"D6",X"DD",X"75",X"0E",X"DD",X"74",
		X"0F",X"DD",X"5E",X"0A",X"DD",X"56",X"0B",X"19",X"DD",X"75",X"02",X"DD",X"74",X"03",X"DD",X"6E",
		X"10",X"DD",X"66",X"11",X"11",X"49",X"00",X"DD",X"CB",X"00",X"46",X"28",X"0D",X"ED",X"52",X"30",
		X"16",X"DD",X"CB",X"00",X"86",X"21",X"00",X"00",X"18",X"0D",X"19",X"E5",X"11",X"00",X"FE",X"19",
		X"E1",X"30",X"04",X"DD",X"CB",X"00",X"C6",X"DD",X"75",X"10",X"DD",X"74",X"11",X"DD",X"5E",X"0C",
		X"DD",X"56",X"0D",X"19",X"DD",X"75",X"04",X"DD",X"74",X"05",X"C3",X"25",X"30",X"DD",X"36",X"01",
		X"06",X"3A",X"71",X"E3",X"DD",X"77",X"08",X"11",X"40",X"00",X"DD",X"6E",X"02",X"DD",X"66",X"03",
		X"ED",X"52",X"DD",X"75",X"0A",X"DD",X"74",X"0B",X"DD",X"73",X"0E",X"DD",X"72",X"0F",X"11",X"00",
		X"01",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"ED",X"52",X"DD",X"75",X"0C",X"DD",X"74",X"0D",X"DD",
		X"73",X"10",X"DD",X"72",X"11",X"C9",X"CD",X"3A",X"33",X"3E",X"86",X"CD",X"FE",X"0D",X"FD",X"21",
		X"82",X"E3",X"06",X"10",X"0E",X"0A",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"FD",X"CB",X"00",X"66",
		X"20",X"2A",X"FD",X"CB",X"00",X"E6",X"FD",X"36",X"07",X"07",X"FD",X"36",X"06",X"14",X"FD",X"75",
		X"02",X"FD",X"74",X"03",X"11",X"00",X"74",X"FD",X"73",X"04",X"FD",X"72",X"05",X"FD",X"71",X"01",
		X"3A",X"81",X"E3",X"3C",X"32",X"81",X"E3",X"79",X"0C",X"FE",X"0C",X"C8",X"11",X"13",X"00",X"FD",
		X"19",X"10",X"C9",X"C9",X"ED",X"5B",X"76",X"E3",X"CD",X"70",X"1C",X"18",X"10",X"CD",X"E2",X"1B",
		X"ED",X"5B",X"72",X"E3",X"18",X"0E",X"ED",X"5B",X"76",X"E3",X"CD",X"7A",X"1C",X"CD",X"E2",X"1B",
		X"ED",X"5B",X"74",X"E3",X"21",X"00",X"50",X"CD",X"32",X"37",X"DA",X"13",X"37",X"2A",X"0C",X"E8",
		X"11",X"00",X"03",X"ED",X"52",X"30",X"23",X"DD",X"5E",X"02",X"DD",X"56",X"03",X"21",X"E0",X"FF",
		X"19",X"22",X"0F",X"E8",X"21",X"20",X"00",X"19",X"22",X"11",X"E8",X"DD",X"6E",X"04",X"DD",X"66",
		X"05",X"11",X"01",X"00",X"CD",X"72",X"11",X"DA",X"C0",X"31",X"DD",X"35",X"07",X"C0",X"DD",X"36",
		X"07",X"03",X"DD",X"7E",X"06",X"3C",X"FE",X"16",X"20",X"02",X"3E",X"14",X"DD",X"77",X"06",X"C9",
		X"DD",X"6E",X"04",X"DD",X"66",X"05",X"11",X"20",X"01",X"3E",X"91",X"CD",X"FE",X"0D",X"CD",X"E2",
		X"2E",X"C3",X"13",X"37",X"CD",X"E2",X"1B",X"CD",X"73",X"37",X"DA",X"ED",X"32",X"CD",X"46",X"37",
		X"3E",X"91",X"DA",X"27",X"33",X"21",X"00",X"50",X"CD",X"1D",X"37",X"38",X"26",X"C9",X"CD",X"E2",
		X"1B",X"DD",X"35",X"07",X"C0",X"DD",X"34",X"06",X"DD",X"7E",X"06",X"FE",X"10",X"20",X"21",X"DD",
		X"34",X"01",X"3A",X"0B",X"E8",X"CB",X"7F",X"DD",X"CB",X"00",X"F6",X"20",X"13",X"DD",X"CB",X"00",
		X"B6",X"18",X"0D",X"3E",X"86",X"CD",X"FE",X"0D",X"DD",X"36",X"01",X"07",X"DD",X"36",X"06",X"0D",
		X"DD",X"36",X"07",X"07",X"C9",X"CD",X"E2",X"1B",X"21",X"40",X"01",X"CD",X"20",X"12",X"3A",X"02",
		X"E7",X"30",X"0A",X"FE",X"04",X"CA",X"A8",X"32",X"FE",X"05",X"CA",X"A8",X"32",X"FE",X"06",X"28",
		X"34",X"FE",X"07",X"28",X"30",X"3A",X"06",X"E7",X"FE",X"05",X"28",X"29",X"CB",X"69",X"20",X"25",
		X"DD",X"7E",X"06",X"FE",X"12",X"20",X"1E",X"2A",X"0A",X"E8",X"11",X"80",X"06",X"CB",X"71",X"20",
		X"04",X"ED",X"52",X"18",X"01",X"19",X"30",X"0D",X"21",X"00",X"6B",X"11",X"20",X"01",X"CD",X"CA",
		X"36",X"DD",X"CB",X"00",X"EE",X"DD",X"35",X"07",X"C0",X"DD",X"7E",X"06",X"FE",X"13",X"CA",X"A2",
		X"32",X"DD",X"34",X"06",X"3A",X"70",X"E3",X"DD",X"77",X"07",X"C9",X"CD",X"E2",X"1B",X"DD",X"35",
		X"07",X"C0",X"DD",X"7E",X"06",X"FE",X"18",X"CA",X"13",X"37",X"DD",X"34",X"06",X"DD",X"36",X"07",
		X"07",X"C9",X"DD",X"36",X"06",X"17",X"18",X"17",X"3E",X"86",X"CD",X"FE",X"0D",X"DD",X"6E",X"02",
		X"DD",X"66",X"03",X"11",X"DC",X"00",X"3E",X"88",X"CD",X"60",X"2F",X"DD",X"36",X"06",X"16",X"DD",
		X"36",X"01",X"09",X"DD",X"36",X"07",X"07",X"C9",X"CD",X"E2",X"1B",X"DD",X"35",X"07",X"C0",X"DD",
		X"7E",X"06",X"DD",X"34",X"06",X"DD",X"36",X"07",X"07",X"FE",X"0C",X"C0",X"DD",X"7E",X"0E",X"A7",
		X"FC",X"BA",X"3C",X"C3",X"13",X"37",X"3E",X"93",X"CD",X"FE",X"0D",X"18",X"05",X"3E",X"86",X"CD",
		X"FE",X"0D",X"3A",X"01",X"E7",X"E6",X"01",X"20",X"07",X"06",X"84",X"11",X"81",X"80",X"18",X"05",
		X"06",X"82",X"11",X"80",X"8C",X"ED",X"5F",X"E6",X"7F",X"FE",X"2A",X"38",X"2F",X"43",X"FE",X"55",
		X"38",X"2A",X"42",X"18",X"27",X"06",X"88",X"3E",X"86",X"CD",X"FE",X"0D",X"18",X"1E",X"06",X"87",
		X"3E",X"86",X"CD",X"FE",X"0D",X"18",X"15",X"CD",X"FE",X"0D",X"DD",X"6E",X"04",X"DD",X"66",X"05",
		X"11",X"80",X"02",X"19",X"11",X"20",X"01",X"CD",X"CA",X"36",X"06",X"00",X"DD",X"70",X"0E",X"DD",
		X"36",X"07",X"07",X"DD",X"36",X"01",X"05",X"DD",X"36",X"06",X"0A",X"C9",X"3E",X"86",X"CD",X"FE",
		X"0D",X"18",X"E7",X"CD",X"F6",X"36",X"DD",X"7E",X"02",X"FD",X"77",X"02",X"DD",X"7E",X"03",X"FD",
		X"77",X"03",X"DD",X"7E",X"04",X"FD",X"77",X"04",X"DD",X"7E",X"05",X"FD",X"77",X"05",X"FD",X"CB",
		X"00",X"E6",X"FD",X"36",X"07",X"07",X"FD",X"36",X"01",X"05",X"FD",X"36",X"06",X"0A",X"C9",X"CD",
		X"E2",X"1B",X"CD",X"73",X"37",X"DA",X"E6",X"32",X"CD",X"46",X"37",X"3E",X"93",X"38",X"98",X"21",
		X"00",X"50",X"CD",X"1D",X"37",X"38",X"2B",X"C9",X"CD",X"E2",X"1B",X"CD",X"73",X"37",X"DA",X"F2",
		X"32",X"DD",X"35",X"07",X"C0",X"DD",X"36",X"07",X"05",X"DD",X"34",X"06",X"DD",X"7E",X"06",X"FE",
		X"07",X"20",X"7F",X"3A",X"0B",X"E8",X"CB",X"7F",X"DD",X"CB",X"00",X"F6",X"C8",X"DD",X"CB",X"00",
		X"B6",X"C9",X"DD",X"36",X"01",X"03",X"DD",X"36",X"07",X"05",X"DD",X"36",X"06",X"04",X"3E",X"93",
		X"CD",X"FE",X"0D",X"C9",X"ED",X"5B",X"6E",X"E3",X"CD",X"7A",X"1C",X"CD",X"E2",X"1B",X"11",X"00",
		X"E4",X"19",X"DA",X"13",X"37",X"CB",X"69",X"20",X"33",X"3A",X"02",X"E7",X"FE",X"0C",X"28",X"2C",
		X"2A",X"0A",X"E8",X"11",X"E0",X"00",X"CB",X"71",X"28",X"04",X"ED",X"52",X"18",X"01",X"19",X"30",
		X"1B",X"2A",X"10",X"E7",X"11",X"00",X"AD",X"19",X"38",X"12",X"21",X"00",X"56",X"11",X"20",X"03",
		X"3E",X"94",X"CD",X"FE",X"0D",X"CD",X"CA",X"36",X"DD",X"CB",X"00",X"EE",X"DD",X"35",X"07",X"C0",
		X"DD",X"36",X"07",X"09",X"DD",X"7E",X"06",X"3C",X"FE",X"0A",X"20",X"02",X"3E",X"08",X"DD",X"77",
		X"06",X"C9",X"FE",X"08",X"C0",X"DD",X"36",X"01",X"04",X"DD",X"36",X"06",X"08",X"DD",X"36",X"07",
		X"09",X"C3",X"B3",X"33",X"ED",X"5B",X"72",X"E3",X"CD",X"7A",X"1C",X"CD",X"E2",X"1B",X"CD",X"BF",
		X"37",X"DA",X"15",X"33",X"CD",X"92",X"37",X"3E",X"91",X"DA",X"27",X"33",X"DD",X"35",X"08",X"CA",
		X"6B",X"35",X"DD",X"35",X"07",X"C8",X"DD",X"36",X"07",X"0B",X"DD",X"7E",X"06",X"3C",X"FE",X"1B",
		X"38",X"02",X"3E",X"19",X"DD",X"77",X"06",X"C9",X"ED",X"5B",X"74",X"E3",X"CD",X"7A",X"1C",X"2A",
		X"6A",X"E3",X"18",X"0A",X"ED",X"5B",X"76",X"E3",X"CD",X"7A",X"1C",X"2A",X"6C",X"E3",X"22",X"00",
		X"E8",X"CD",X"E2",X"1B",X"CD",X"BF",X"37",X"DA",X"15",X"33",X"CD",X"92",X"37",X"3E",X"91",X"DA",
		X"27",X"33",X"ED",X"5B",X"00",X"E8",X"21",X"00",X"50",X"CD",X"32",X"37",X"38",X"16",X"DD",X"35",
		X"07",X"C8",X"DD",X"36",X"07",X"0B",X"DD",X"7E",X"06",X"3C",X"FE",X"1D",X"38",X"02",X"3E",X"1B",
		X"DD",X"77",X"06",X"C9",X"3E",X"86",X"CD",X"FE",X"0D",X"ED",X"5F",X"E6",X"03",X"CA",X"18",X"32",
		X"F5",X"CD",X"53",X"33",X"F1",X"FE",X"01",X"CA",X"35",X"34",X"C3",X"13",X"37",X"CD",X"F6",X"36",
		X"DD",X"6E",X"02",X"DD",X"66",X"03",X"11",X"00",X"02",X"DD",X"7E",X"00",X"E6",X"40",X"28",X"03",
		X"19",X"18",X"02",X"ED",X"52",X"FD",X"75",X"02",X"FD",X"74",X"03",X"EE",X"50",X"FD",X"77",X"00",
		X"DD",X"7E",X"0E",X"C6",X"0C",X"FD",X"77",X"01",X"87",X"5F",X"16",X"00",X"21",X"17",X"35",X"19",
		X"5E",X"FD",X"73",X"04",X"23",X"5E",X"FD",X"73",X"05",X"FD",X"36",X"07",X"0B",X"FE",X"1A",X"20",
		X"0B",X"FD",X"36",X"06",X"19",X"3A",X"65",X"E3",X"FD",X"77",X"08",X"C9",X"FD",X"36",X"06",X"1B",
		X"C9",X"00",X"66",X"00",X"5F",X"00",X"5A",X"ED",X"5B",X"63",X"E3",X"CD",X"7A",X"1C",X"CD",X"E2",
		X"1B",X"CD",X"73",X"37",X"DA",X"15",X"33",X"CD",X"46",X"37",X"3E",X"94",X"DA",X"27",X"33",X"DD",
		X"35",X"08",X"CA",X"4C",X"33",X"DD",X"35",X"07",X"C0",X"DD",X"36",X"07",X"0B",X"DD",X"7E",X"06",
		X"3C",X"FE",X"1F",X"38",X"02",X"3E",X"1D",X"DD",X"77",X"06",X"C9",X"CD",X"53",X"33",X"3E",X"86",
		X"CD",X"FE",X"0D",X"ED",X"5F",X"E6",X"01",X"CA",X"13",X"37",X"3E",X"40",X"DD",X"AE",X"00",X"DD",
		X"77",X"00",X"DD",X"36",X"01",X"10",X"DD",X"36",X"06",X"1D",X"DD",X"36",X"07",X"0B",X"3A",X"66",
		X"E3",X"DD",X"77",X"08",X"C9",X"3A",X"60",X"E3",X"ED",X"5B",X"12",X"E7",X"2A",X"61",X"E3",X"ED",
		X"52",X"38",X"0B",X"2A",X"63",X"E3",X"ED",X"52",X"38",X"0B",X"FE",X"01",X"18",X"01",X"A7",X"C0",
		X"AF",X"32",X"00",X"E1",X"C9",X"21",X"80",X"E3",X"35",X"C0",X"34",X"23",X"7E",X"FE",X"10",X"D0",
		X"3A",X"17",X"E0",X"21",X"6A",X"E3",X"1E",X"00",X"BE",X"38",X"1D",X"23",X"1C",X"BE",X"38",X"18",
		X"1C",X"3A",X"16",X"E0",X"FE",X"7F",X"3E",X"F8",X"38",X"02",X"3E",X"06",X"21",X"01",X"E7",X"CB",
		X"76",X"20",X"02",X"ED",X"44",X"57",X"18",X"23",X"3A",X"16",X"E0",X"16",X"F7",X"FE",X"2A",X"38",
		X"1A",X"16",X"FA",X"FE",X"55",X"38",X"14",X"16",X"FD",X"FE",X"7F",X"38",X"0E",X"16",X"03",X"FE",
		X"AA",X"38",X"08",X"16",X"06",X"FE",X"D4",X"38",X"02",X"16",X"09",X"3A",X"02",X"E7",X"FE",X"01",
		X"28",X"06",X"FE",X"09",X"3E",X"03",X"20",X"02",X"3E",X"06",X"21",X"01",X"E7",X"CB",X"76",X"28",
		X"02",X"ED",X"44",X"BA",X"20",X"02",X"16",X"00",X"3A",X"02",X"E7",X"FE",X"01",X"28",X"06",X"FE",
		X"09",X"3E",X"03",X"20",X"02",X"3E",X"09",X"CB",X"76",X"20",X"02",X"ED",X"44",X"82",X"57",X"3A",
		X"13",X"E7",X"82",X"57",X"CB",X"C2",X"EB",X"DD",X"21",X"6F",X"E3",X"11",X"13",X"00",X"06",X"10",
		X"DD",X"19",X"DD",X"CB",X"00",X"66",X"28",X"14",X"DD",X"7E",X"01",X"FE",X"03",X"38",X"08",X"FE",
		X"06",X"38",X"09",X"FE",X"09",X"30",X"05",X"DD",X"7E",X"12",X"BC",X"C8",X"10",X"E2",X"EB",X"3A",
		X"15",X"E0",X"21",X"65",X"E3",X"CD",X"14",X"12",X"21",X"80",X"E3",X"77",X"23",X"34",X"DD",X"21",
		X"6F",X"E3",X"01",X"13",X"00",X"DD",X"09",X"DD",X"CB",X"00",X"66",X"20",X"F8",X"ED",X"5F",X"E6",
		X"40",X"F6",X"10",X"DD",X"77",X"00",X"DD",X"73",X"01",X"DD",X"73",X"06",X"DD",X"72",X"12",X"DD",
		X"72",X"03",X"DD",X"36",X"02",X"00",X"21",X"00",X"90",X"DD",X"75",X"04",X"DD",X"74",X"05",X"DD",
		X"36",X"07",X"03",X"21",X"0A",X"00",X"11",X"7D",X"00",X"DD",X"75",X"0A",X"DD",X"74",X"0B",X"2A",
		X"6C",X"E3",X"19",X"DD",X"75",X"0C",X"DD",X"74",X"0D",X"C9",X"3A",X"80",X"E0",X"E6",X"07",X"FE",
		X"03",X"20",X"11",X"3A",X"09",X"E7",X"93",X"F2",X"E4",X"36",X"CD",X"08",X"12",X"20",X"05",X"3E",
		X"05",X"32",X"07",X"E0",X"C3",X"E2",X"2E",X"2A",X"0C",X"E8",X"11",X"00",X"E4",X"19",X"D8",X"21",
		X"8E",X"74",X"79",X"C3",X"7E",X"1A",X"3A",X"81",X"E3",X"FE",X"10",X"30",X"14",X"3C",X"32",X"81",
		X"E3",X"FD",X"21",X"6F",X"E3",X"11",X"13",X"00",X"FD",X"19",X"FD",X"CB",X"00",X"66",X"20",X"F8",
		X"C9",X"F1",X"C9",X"DD",X"36",X"00",X"00",X"21",X"81",X"E3",X"35",X"F1",X"C9",X"E5",X"DD",X"6E",
		X"0A",X"DD",X"66",X"0B",X"DD",X"5E",X"0C",X"DD",X"56",X"0D",X"19",X"DD",X"75",X"0C",X"DD",X"74",
		X"0D",X"E1",X"E5",X"A7",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"ED",X"52",X"DD",X"75",X"04",X"DD",
		X"74",X"05",X"D1",X"ED",X"52",X"C9",X"2A",X"0C",X"E8",X"11",X"00",X"03",X"ED",X"52",X"D0",X"DD",
		X"5E",X"02",X"DD",X"56",X"03",X"21",X"80",X"FF",X"19",X"22",X"0F",X"E8",X"21",X"80",X"00",X"19",
		X"22",X"11",X"E8",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"11",X"80",X"00",X"19",X"11",X"08",X"00",
		X"C3",X"72",X"11",X"21",X"40",X"01",X"CD",X"20",X"12",X"D0",X"A7",X"DD",X"6E",X"04",X"DD",X"66",
		X"05",X"ED",X"52",X"D0",X"21",X"00",X"F8",X"19",X"DD",X"5E",X"04",X"DD",X"56",X"05",X"A7",X"ED",
		X"52",X"C9",X"2A",X"0C",X"E8",X"11",X"00",X"03",X"ED",X"52",X"D0",X"DD",X"5E",X"02",X"DD",X"56",
		X"03",X"21",X"C0",X"FF",X"19",X"22",X"0F",X"E8",X"21",X"40",X"00",X"19",X"22",X"11",X"E8",X"DD",
		X"6E",X"04",X"DD",X"66",X"05",X"11",X"80",X"00",X"19",X"11",X"04",X"00",X"C3",X"72",X"11",X"21",
		X"E0",X"00",X"CD",X"20",X"12",X"D0",X"A7",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"ED",X"52",X"D0",
		X"21",X"80",X"FB",X"19",X"DD",X"5E",X"04",X"DD",X"56",X"05",X"A7",X"ED",X"52",X"C9",X"2A",X"12",
		X"E7",X"11",X"00",X"80",X"19",X"38",X"0A",X"CD",X"F6",X"37",X"CD",X"FF",X"38",X"CD",X"60",X"39",
		X"C9",X"AF",X"32",X"00",X"E1",X"C9",X"06",X"04",X"21",X"72",X"E5",X"7E",X"A7",X"28",X"05",X"35",
		X"23",X"10",X"F8",X"C9",X"C5",X"E5",X"3A",X"80",X"E0",X"FE",X"10",X"21",X"DB",X"38",X"38",X"03",
		X"21",X"EB",X"38",X"16",X"00",X"58",X"CB",X"03",X"CB",X"03",X"19",X"5E",X"23",X"56",X"E5",X"ED",
		X"4B",X"12",X"E7",X"21",X"40",X"0F",X"09",X"ED",X"52",X"DA",X"D9",X"38",X"21",X"C0",X"F0",X"09",
		X"ED",X"52",X"D2",X"D9",X"38",X"21",X"76",X"E5",X"3A",X"0B",X"E5",X"BE",X"DA",X"D9",X"38",X"34",
		X"FD",X"21",X"62",X"E5",X"01",X"15",X"00",X"FD",X"09",X"FD",X"CB",X"00",X"66",X"20",X"F8",X"FD",
		X"73",X"02",X"FD",X"72",X"03",X"2A",X"12",X"E7",X"3E",X"10",X"ED",X"52",X"38",X"02",X"3E",X"50",
		X"FD",X"77",X"00",X"CD",X"C5",X"3D",X"D5",X"3A",X"12",X"E0",X"21",X"0D",X"E5",X"BE",X"30",X"0F",
		X"FD",X"CB",X"14",X"CE",X"E6",X"02",X"3E",X"38",X"28",X"02",X"3E",X"A9",X"FD",X"77",X"13",X"3A",
		X"13",X"E0",X"21",X"0E",X"E5",X"BE",X"30",X"0E",X"FD",X"CB",X"14",X"C6",X"E6",X"02",X"23",X"28",
		X"01",X"23",X"7E",X"FD",X"77",X"12",X"D1",X"E1",X"23",X"7E",X"23",X"66",X"6F",X"FD",X"75",X"04",
		X"FD",X"74",X"05",X"ED",X"52",X"FD",X"75",X"0C",X"FD",X"74",X"0D",X"F5",X"FD",X"7E",X"01",X"C6",
		X"04",X"FD",X"77",X"01",X"FE",X"04",X"28",X"09",X"F1",X"ED",X"5F",X"CB",X"47",X"28",X"05",X"18",
		X"07",X"F1",X"38",X"04",X"FD",X"CB",X"00",X"DE",X"FD",X"36",X"06",X"06",X"FD",X"36",X"07",X"10",
		X"3A",X"0A",X"E5",X"E1",X"77",X"C1",X"C3",X"00",X"38",X"E1",X"E1",X"C1",X"C3",X"00",X"38",X"00",
		X"71",X"00",X"80",X"00",X"5B",X"00",X"54",X"00",X"3D",X"00",X"70",X"00",X"23",X"00",X"80",X"00",
		X"71",X"00",X"80",X"00",X"5B",X"00",X"70",X"00",X"3D",X"00",X"70",X"00",X"23",X"00",X"80",X"3A",
		X"20",X"E5",X"A7",X"C8",X"47",X"DD",X"21",X"21",X"E5",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"11",
		X"29",X"00",X"ED",X"52",X"EB",X"21",X"00",X"08",X"ED",X"52",X"38",X"05",X"CD",X"0E",X"3D",X"18",
		X"24",X"DD",X"73",X"00",X"DD",X"72",X"01",X"2A",X"12",X"E7",X"ED",X"52",X"38",X"0A",X"11",X"00",
		X"F0",X"19",X"38",X"25",X"0E",X"FF",X"18",X"08",X"11",X"00",X"10",X"19",X"30",X"1B",X"0E",X"00",
		X"C5",X"CD",X"55",X"3D",X"C1",X"21",X"20",X"E5",X"35",X"C8",X"05",X"C8",X"7E",X"23",X"07",X"16",
		X"00",X"5F",X"19",X"7E",X"23",X"66",X"6F",X"18",X"B6",X"DD",X"23",X"DD",X"23",X"10",X"AA",X"C9",
		X"3A",X"49",X"E5",X"A7",X"C8",X"47",X"DD",X"21",X"4A",X"E5",X"DD",X"6E",X"00",X"DD",X"66",X"01",
		X"11",X"29",X"00",X"19",X"EB",X"21",X"00",X"80",X"ED",X"52",X"30",X"05",X"CD",X"09",X"3D",X"18",
		X"24",X"DD",X"73",X"00",X"DD",X"72",X"01",X"2A",X"12",X"E7",X"ED",X"52",X"38",X"0A",X"11",X"00",
		X"F0",X"19",X"38",X"25",X"0E",X"FF",X"18",X"08",X"11",X"00",X"10",X"19",X"30",X"1B",X"0E",X"00",
		X"C5",X"CD",X"59",X"3D",X"C1",X"21",X"49",X"E5",X"35",X"C8",X"05",X"C8",X"7E",X"23",X"07",X"16",
		X"00",X"5F",X"19",X"7E",X"23",X"66",X"6F",X"18",X"B7",X"DD",X"23",X"DD",X"23",X"10",X"AB",X"C9",
		X"3A",X"76",X"E5",X"A7",X"C8",X"DD",X"21",X"77",X"E5",X"3A",X"0B",X"E5",X"47",X"C5",X"DD",X"4E",
		X"00",X"CB",X"61",X"C4",X"DF",X"39",X"C1",X"11",X"15",X"00",X"DD",X"19",X"10",X"EF",X"C9",X"DD",
		X"7E",X"01",X"FE",X"04",X"38",X"0B",X"FE",X"07",X"DA",X"3B",X"3C",X"CA",X"E9",X"3B",X"C3",X"1F",
		X"3B",X"DD",X"35",X"07",X"20",X"0D",X"DD",X"36",X"07",X"05",X"DD",X"35",X"06",X"28",X"04",X"DD",
		X"36",X"06",X"01",X"DD",X"CB",X"14",X"4E",X"28",X"1D",X"DD",X"35",X"13",X"20",X"18",X"DD",X"CB",
		X"14",X"56",X"20",X"0A",X"DD",X"CB",X"14",X"D6",X"DD",X"36",X"13",X"A9",X"18",X"08",X"DD",X"CB",
		X"14",X"96",X"DD",X"CB",X"14",X"8E",X"DD",X"CB",X"14",X"46",X"28",X"06",X"DD",X"35",X"12",X"CA",
		X"92",X"3B",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"DD",X"5E",X"10",X"DD",X"56",X"11",X"DD",X"CB",
		X"14",X"56",X"28",X"03",X"11",X"00",X"00",X"CB",X"71",X"20",X"13",X"ED",X"52",X"EB",X"21",X"00",
		X"F4",X"19",X"38",X"1C",X"DD",X"CB",X"00",X"F6",X"21",X"AB",X"3E",X"C3",X"AA",X"3B",X"19",X"EB",
		X"21",X"00",X"84",X"19",X"30",X"0A",X"DD",X"CB",X"00",X"B6",X"21",X"7F",X"3E",X"C3",X"AA",X"3B",
		X"DD",X"73",X"02",X"DD",X"72",X"03",X"D5",X"2A",X"12",X"E7",X"ED",X"52",X"11",X"00",X"11",X"38",
		X"08",X"ED",X"52",X"D1",X"38",X"0E",X"C3",X"FB",X"3C",X"19",X"D1",X"38",X"07",X"21",X"00",X"DF",
		X"19",X"DA",X"FB",X"3C",X"FE",X"03",X"28",X"5C",X"CD",X"22",X"3D",X"3D",X"FA",X"E4",X"3A",X"D5",
		X"DD",X"6E",X"0C",X"DD",X"66",X"0D",X"28",X"06",X"ED",X"5B",X"04",X"E5",X"18",X"04",X"ED",X"5B",
		X"06",X"E5",X"CB",X"59",X"28",X"0D",X"ED",X"52",X"EB",X"CB",X"7A",X"28",X"1E",X"DD",X"CB",X"00",
		X"9E",X"18",X"18",X"19",X"EB",X"CB",X"7A",X"20",X"12",X"A7",X"28",X"05",X"21",X"00",X"EC",X"18",
		X"03",X"21",X"00",X"F0",X"19",X"30",X"04",X"DD",X"CB",X"00",X"DE",X"DD",X"73",X"0C",X"DD",X"72",
		X"0D",X"E1",X"19",X"EB",X"DD",X"6E",X"08",X"DD",X"66",X"09",X"19",X"DD",X"75",X"04",X"DD",X"74",
		X"05",X"C3",X"7A",X"3C",X"CD",X"22",X"3D",X"D5",X"ED",X"5B",X"04",X"E5",X"DD",X"6E",X"0C",X"DD",
		X"66",X"0D",X"CB",X"59",X"28",X"04",X"ED",X"52",X"18",X"01",X"19",X"30",X"07",X"DD",X"36",X"01",
		X"00",X"21",X"00",X"00",X"DD",X"75",X"0C",X"DD",X"74",X"0D",X"D1",X"19",X"EB",X"18",X"C5",X"DD",
		X"6E",X"0E",X"DD",X"66",X"0F",X"DD",X"35",X"07",X"20",X"09",X"11",X"05",X"00",X"19",X"CD",X"D5",
		X"3B",X"28",X"24",X"7E",X"DD",X"86",X"02",X"DD",X"77",X"02",X"23",X"7E",X"DD",X"8E",X"03",X"DD",
		X"77",X"03",X"23",X"7E",X"DD",X"86",X"04",X"DD",X"77",X"04",X"23",X"7E",X"DD",X"8E",X"05",X"DD",
		X"77",X"05",X"23",X"4E",X"C3",X"7A",X"3C",X"DD",X"36",X"0A",X"00",X"DD",X"36",X"06",X"00",X"DD",
		X"36",X"07",X"05",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"DD",X"5E",X"08",X"DD",X"56",X"09",X"ED",
		X"52",X"DD",X"75",X"0C",X"DD",X"74",X"0D",X"DD",X"7E",X"01",X"D6",X"08",X"20",X"0E",X"3E",X"03",
		X"DD",X"CB",X"00",X"9E",X"CB",X"7C",X"20",X"04",X"DD",X"CB",X"00",X"DE",X"DD",X"77",X"01",X"C3",
		X"7A",X"3C",X"DD",X"CB",X"14",X"86",X"DD",X"CB",X"00",X"76",X"21",X"7F",X"3E",X"DD",X"CB",X"00",
		X"B6",X"20",X"07",X"DD",X"CB",X"00",X"F6",X"21",X"AB",X"3E",X"E5",X"DD",X"6E",X"04",X"DD",X"66",
		X"05",X"11",X"00",X"98",X"19",X"E1",X"30",X"04",X"11",X"16",X"00",X"19",X"CD",X"D5",X"3B",X"11",
		X"04",X"00",X"19",X"4E",X"DD",X"7E",X"01",X"C6",X"08",X"FE",X"0B",X"20",X"02",X"3E",X"08",X"DD",
		X"77",X"01",X"C3",X"7A",X"3C",X"7E",X"FE",X"FF",X"C8",X"DD",X"77",X"07",X"23",X"7E",X"DD",X"77",
		X"06",X"23",X"DD",X"75",X"0E",X"DD",X"74",X"0F",X"C9",X"DD",X"35",X"07",X"C2",X"A9",X"3C",X"DD",
		X"7E",X"06",X"FE",X"09",X"28",X"0A",X"DD",X"36",X"07",X"05",X"DD",X"34",X"06",X"C3",X"A9",X"3C",
		X"DD",X"7E",X"0E",X"A7",X"CA",X"F2",X"3C",X"CD",X"BA",X"3C",X"C3",X"F2",X"3C",X"3E",X"86",X"CD",
		X"FE",X"0D",X"3A",X"01",X"E7",X"E6",X"01",X"3E",X"83",X"20",X"0F",X"3C",X"18",X"0C",X"11",X"15",
		X"01",X"CD",X"E2",X"2E",X"3E",X"94",X"CD",X"FE",X"0D",X"AF",X"DD",X"77",X"0E",X"DD",X"36",X"07",
		X"05",X"DD",X"36",X"06",X"07",X"DD",X"36",X"01",X"07",X"18",X"6E",X"DD",X"35",X"07",X"28",X"26",
		X"3A",X"00",X"EB",X"F5",X"3E",X"01",X"32",X"00",X"EB",X"2A",X"01",X"EB",X"E5",X"2A",X"03",X"EB",
		X"11",X"F8",X"FF",X"19",X"22",X"01",X"EB",X"22",X"03",X"EB",X"CD",X"A9",X"3C",X"E1",X"22",X"01",
		X"EB",X"F1",X"32",X"00",X"EB",X"C9",X"DD",X"36",X"06",X"00",X"DD",X"36",X"07",X"05",X"DD",X"7E",
		X"01",X"D6",X"04",X"20",X"02",X"3E",X"03",X"DD",X"77",X"01",X"CD",X"CF",X"3C",X"DA",X"0D",X"3C",
		X"DD",X"5E",X"02",X"DD",X"56",X"03",X"21",X"C0",X"FF",X"19",X"22",X"0F",X"E8",X"21",X"80",X"00",
		X"19",X"22",X"11",X"E8",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"11",X"00",X"02",X"19",X"11",X"06",
		X"00",X"E5",X"CD",X"72",X"11",X"E1",X"DA",X"1E",X"3C",X"CD",X"E2",X"1B",X"11",X"00",X"E4",X"19",
		X"D8",X"21",X"C0",X"75",X"79",X"EE",X"40",X"C3",X"80",X"1A",X"DD",X"6E",X"04",X"DD",X"66",X"05",
		X"29",X"16",X"00",X"CB",X"12",X"5C",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"C3",X"60",X"2F",X"21",
		X"40",X"01",X"CD",X"20",X"12",X"D0",X"21",X"80",X"01",X"19",X"EB",X"DD",X"6E",X"04",X"DD",X"66",
		X"05",X"ED",X"52",X"D0",X"21",X"80",X"F3",X"19",X"DD",X"5E",X"04",X"DD",X"56",X"05",X"A7",X"ED",
		X"52",X"C9",X"21",X"76",X"E5",X"35",X"DD",X"36",X"00",X"00",X"C9",X"21",X"76",X"E5",X"35",X"DD",
		X"CB",X"00",X"76",X"DD",X"36",X"00",X"00",X"20",X"05",X"21",X"20",X"E5",X"18",X"03",X"21",X"49",
		X"E5",X"7E",X"FE",X"14",X"C8",X"34",X"23",X"C5",X"07",X"06",X"00",X"4F",X"09",X"73",X"23",X"72",
		X"C1",X"C9",X"DD",X"6E",X"0A",X"DD",X"66",X"0B",X"ED",X"5B",X"08",X"E5",X"DD",X"CB",X"00",X"56",
		X"28",X"0E",X"ED",X"52",X"EB",X"30",X"15",X"DD",X"CB",X"00",X"96",X"11",X"00",X"00",X"18",X"0C",
		X"19",X"EB",X"21",X"00",X"FC",X"19",X"30",X"04",X"DD",X"CB",X"00",X"D6",X"DD",X"73",X"0A",X"DD",
		X"72",X"0B",X"C9",X"0E",X"00",X"06",X"10",X"18",X"02",X"06",X"50",X"21",X"76",X"E5",X"3A",X"0B",
		X"E5",X"BE",X"D8",X"34",X"FD",X"21",X"62",X"E5",X"11",X"15",X"00",X"FD",X"19",X"FD",X"CB",X"00",
		X"66",X"20",X"F8",X"ED",X"5F",X"E6",X"0C",X"B0",X"FD",X"77",X"00",X"2A",X"12",X"E7",X"11",X"80",
		X"10",X"CB",X"41",X"28",X"04",X"ED",X"52",X"18",X"0A",X"19",X"11",X"80",X"20",X"ED",X"52",X"19",
		X"30",X"01",X"EB",X"FD",X"75",X"02",X"FD",X"74",X"03",X"FD",X"36",X"07",X"05",X"FD",X"36",X"06",
		X"00",X"CD",X"C5",X"3D",X"FD",X"7E",X"01",X"FE",X"01",X"D8",X"21",X"5F",X"3E",X"28",X"03",X"21",
		X"6F",X"3E",X"3A",X"10",X"E0",X"E6",X"0E",X"16",X"00",X"5F",X"19",X"7E",X"FD",X"77",X"0C",X"23",
		X"7E",X"FD",X"77",X"0D",X"C9",X"21",X"49",X"E6",X"7E",X"A7",X"20",X"0F",X"36",X"03",X"ED",X"5F",
		X"E6",X"1C",X"21",X"1F",X"3E",X"16",X"00",X"5F",X"19",X"18",X"04",X"35",X"2A",X"4A",X"E6",X"7E",
		X"23",X"22",X"4A",X"E6",X"FD",X"77",X"01",X"FD",X"36",X"14",X"00",X"21",X"3F",X"3E",X"A7",X"28",
		X"03",X"21",X"4F",X"3E",X"ED",X"5F",X"E6",X"0E",X"16",X"00",X"5F",X"19",X"5E",X"23",X"56",X"FD",
		X"73",X"08",X"FD",X"72",X"09",X"FD",X"36",X"0B",X"02",X"3A",X"11",X"E0",X"21",X"0C",X"E5",X"BE",
		X"2A",X"00",X"E5",X"38",X"03",X"2A",X"02",X"E5",X"FD",X"75",X"10",X"FD",X"74",X"11",X"C9",X"02",
		X"00",X"01",X"00",X"01",X"02",X"00",X"00",X"00",X"00",X"02",X"01",X"00",X"01",X"00",X"02",X"02",
		X"00",X"00",X"01",X"00",X"02",X"01",X"00",X"00",X"01",X"02",X"00",X"01",X"00",X"00",X"02",X"00",
		X"50",X"80",X"54",X"00",X"59",X"80",X"5D",X"00",X"62",X"80",X"66",X"00",X"6B",X"80",X"6F",X"00",
		X"4E",X"80",X"51",X"00",X"55",X"80",X"58",X"00",X"5C",X"80",X"5F",X"00",X"63",X"80",X"66",X"00",
		X"00",X"80",X"02",X"00",X"05",X"00",X"07",X"80",X"09",X"80",X"0B",X"00",X"0E",X"00",X"10",X"00",
		X"00",X"00",X"03",X"00",X"06",X"80",X"08",X"80",X"0B",X"00",X"0E",X"00",X"0C",X"00",X"14",X"12",
		X"02",X"2A",X"00",X"47",X"00",X"40",X"12",X"03",X"00",X"00",X"8E",X"00",X"40",X"12",X"02",X"D6",
		X"FF",X"47",X"00",X"00",X"FF",X"12",X"04",X"2A",X"00",X"B9",X"FF",X"C0",X"12",X"05",X"00",X"00",
		X"72",X"FF",X"C0",X"12",X"04",X"D6",X"FF",X"B9",X"FF",X"80",X"FF",X"12",X"02",X"D6",X"FF",X"47",
		X"00",X"00",X"12",X"03",X"00",X"00",X"8E",X"00",X"00",X"12",X"02",X"2A",X"00",X"47",X"00",X"40",
		X"FF",X"12",X"04",X"D6",X"FF",X"B9",X"FF",X"80",X"12",X"05",X"00",X"00",X"72",X"FF",X"80",X"12",
		X"04",X"2A",X"00",X"B9",X"FF",X"C0",X"FF",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"2A",X"12",X"E7",X"ED",X"5B",X"07",X"E7",X"3A",X"80",X"E0",X"E6",X"01",X"28",X"01",X"EB",X"ED",
		X"52",X"3E",X"01",X"30",X"02",X"3E",X"00",X"32",X"02",X"E7",X"38",X"10",X"21",X"03",X"E7",X"7E",
		X"35",X"A7",X"20",X"08",X"CD",X"3F",X"43",X"3E",X"90",X"CD",X"FE",X"0D",X"2A",X"12",X"E7",X"3A",
		X"1A",X"E7",X"A7",X"C2",X"AD",X"40",X"3A",X"00",X"E0",X"FE",X"03",X"28",X"70",X"3A",X"02",X"E7",
		X"FE",X"0B",X"28",X"69",X"30",X"3A",X"FE",X"09",X"30",X"0B",X"FE",X"01",X"20",X"5F",X"3A",X"06",
		X"E7",X"FE",X"04",X"28",X"58",X"3A",X"00",X"E7",X"CB",X"6F",X"3A",X"01",X"E7",X"11",X"29",X"00",
		X"28",X"27",X"E6",X"20",X"20",X"47",X"19",X"11",X"00",X"DB",X"ED",X"52",X"19",X"38",X"01",X"EB",
		X"E5",X"7C",X"D6",X"0F",X"21",X"14",X"E7",X"BE",X"20",X"2F",X"34",X"7E",X"C6",X"1F",X"18",X"26",
		X"3A",X"00",X"E7",X"E6",X"20",X"20",X"11",X"18",X"E7",X"E6",X"10",X"20",X"20",X"ED",X"52",X"11",
		X"00",X"04",X"ED",X"52",X"19",X"30",X"01",X"EB",X"E5",X"3E",X"10",X"84",X"21",X"14",X"E7",X"BE",
		X"20",X"07",X"35",X"7E",X"C6",X"E0",X"CD",X"65",X"57",X"E1",X"22",X"12",X"E7",X"AF",X"29",X"17",
		X"29",X"17",X"29",X"17",X"6C",X"67",X"11",X"80",X"00",X"ED",X"52",X"38",X"11",X"19",X"11",X"80",
		X"06",X"ED",X"52",X"30",X"09",X"19",X"22",X"00",X"E9",X"21",X"00",X"01",X"18",X"08",X"ED",X"53",
		X"00",X"E9",X"11",X"00",X"01",X"19",X"22",X"15",X"E7",X"AF",X"2A",X"10",X"E7",X"29",X"17",X"6C",
		X"67",X"22",X"17",X"E7",X"C9",X"2A",X"17",X"E7",X"22",X"07",X"E8",X"3A",X"06",X"E7",X"87",X"21",
		X"FF",X"65",X"06",X"00",X"4F",X"09",X"7E",X"23",X"66",X"6F",X"3A",X"01",X"E7",X"E6",X"40",X"ED",
		X"5B",X"15",X"E7",X"CD",X"20",X"0E",X"3A",X"00",X"E0",X"FE",X"05",X"C8",X"FE",X"07",X"C8",X"FE",
		X"03",X"2A",X"00",X"E9",X"20",X"1E",X"EB",X"2A",X"02",X"E9",X"3A",X"01",X"E1",X"01",X"02",X"00",
		X"A7",X"20",X"08",X"ED",X"42",X"ED",X"52",X"30",X"07",X"18",X"08",X"09",X"ED",X"52",X"30",X"03",
		X"19",X"18",X"01",X"EB",X"22",X"02",X"E9",X"3A",X"3F",X"E3",X"A7",X"CC",X"C1",X"2E",X"C9",X"CD",
		X"08",X"12",X"20",X"0C",X"2A",X"03",X"E0",X"7C",X"B5",X"20",X"05",X"21",X"1F",X"E7",X"CB",X"CE",
		X"CD",X"74",X"41",X"21",X"00",X"E7",X"CB",X"66",X"28",X"0E",X"CB",X"6E",X"28",X"05",X"CB",X"76",
		X"20",X"0E",X"C9",X"CB",X"76",X"28",X"05",X"C9",X"CB",X"6E",X"20",X"04",X"23",X"CB",X"B6",X"C9",
		X"23",X"CB",X"F6",X"C9",X"21",X"19",X"E7",X"35",X"C2",X"9A",X"41",X"3A",X"80",X"E0",X"E6",X"18",
		X"FE",X"08",X"16",X"00",X"38",X"0C",X"16",X"A9",X"28",X"08",X"FE",X"10",X"16",X"70",X"28",X"02",
		X"16",X"38",X"72",X"21",X"01",X"E7",X"7E",X"EE",X"80",X"77",X"3A",X"00",X"E0",X"FE",X"03",X"CA",
		X"A0",X"46",X"CD",X"04",X"47",X"21",X"02",X"E7",X"7E",X"FE",X"0D",X"CA",X"F6",X"45",X"FE",X"04",
		X"DA",X"89",X"42",X"FE",X"0B",X"CA",X"DE",X"44",X"D2",X"02",X"45",X"FE",X"08",X"D2",X"06",X"44",
		X"3A",X"1F",X"E7",X"E6",X"01",X"C2",X"51",X"45",X"3A",X"09",X"E9",X"57",X"7E",X"FE",X"06",X"30",
		X"05",X"CB",X"52",X"C2",X"87",X"43",X"CB",X"5A",X"C2",X"B5",X"43",X"21",X"00",X"E7",X"CB",X"4A",
		X"28",X"02",X"CB",X"AE",X"CB",X"42",X"28",X"02",X"CB",X"EE",X"21",X"03",X"E7",X"35",X"20",X"39",
		X"3A",X"04",X"E7",X"3C",X"28",X"4A",X"3D",X"20",X"19",X"3C",X"32",X"04",X"E7",X"2A",X"0A",X"E7",
		X"7E",X"32",X"03",X"E7",X"23",X"3A",X"01",X"E7",X"A6",X"32",X"01",X"E7",X"23",X"7E",X"32",X"06",
		X"E7",X"C9",X"21",X"02",X"E7",X"7E",X"FE",X"06",X"01",X"00",X"04",X"38",X"03",X"01",X"03",X"05",
		X"71",X"78",X"32",X"06",X"E7",X"23",X"36",X"05",X"C9",X"3A",X"04",X"E7",X"3D",X"C0",X"2A",X"0A",
		X"E7",X"23",X"CB",X"4E",X"28",X"05",X"CB",X"6A",X"20",X"0A",X"C9",X"CB",X"62",X"20",X"05",X"C9",
		X"AF",X"32",X"05",X"E7",X"AF",X"32",X"04",X"E7",X"57",X"3A",X"02",X"E7",X"D6",X"04",X"87",X"5F",
		X"87",X"83",X"5F",X"21",X"8D",X"65",X"19",X"7E",X"32",X"03",X"E7",X"23",X"3A",X"01",X"E7",X"B6",
		X"32",X"01",X"E7",X"23",X"CB",X"4F",X"7E",X"23",X"22",X"0A",X"E7",X"21",X"05",X"E7",X"28",X"05",
		X"CB",X"46",X"28",X"01",X"3C",X"32",X"06",X"E7",X"34",X"3A",X"84",X"E8",X"A7",X"C0",X"3E",X"0B",
		X"32",X"84",X"E8",X"3E",X"82",X"CD",X"FE",X"0D",X"C9",X"3A",X"1F",X"E7",X"CB",X"4F",X"C2",X"36",
		X"46",X"CB",X"47",X"C2",X"5A",X"45",X"3A",X"03",X"E7",X"3D",X"FA",X"A0",X"42",X"32",X"03",X"E7",
		X"3A",X"09",X"E9",X"CB",X"6F",X"C2",X"65",X"43",X"CB",X"67",X"C2",X"52",X"43",X"CB",X"5F",X"C2",
		X"BD",X"43",X"CB",X"57",X"C2",X"87",X"43",X"CB",X"4F",X"20",X"4C",X"CB",X"47",X"20",X"20",X"21",
		X"02",X"E7",X"7E",X"FE",X"02",X"36",X"00",X"D2",X"47",X"43",X"FE",X"00",X"3A",X"05",X"E7",X"28",
		X"02",X"3E",X"05",X"3D",X"32",X"05",X"E7",X"C0",X"2A",X"12",X"E7",X"22",X"07",X"E7",X"C9",X"2A",
		X"12",X"E7",X"11",X"00",X"DB",X"ED",X"52",X"28",X"D6",X"21",X"01",X"E7",X"CB",X"6E",X"2B",X"20",
		X"08",X"CB",X"6E",X"20",X"3C",X"CB",X"EE",X"18",X"26",X"CB",X"EE",X"18",X"02",X"CB",X"AE",X"2A",
		X"12",X"E7",X"22",X"07",X"E7",X"18",X"B8",X"2A",X"12",X"E7",X"11",X"00",X"04",X"ED",X"52",X"28",
		X"AE",X"21",X"01",X"E7",X"CB",X"66",X"2B",X"20",X"E4",X"CB",X"6E",X"28",X"14",X"CB",X"AE",X"3A",
		X"02",X"E7",X"FE",X"04",X"20",X"05",X"3E",X"05",X"32",X"03",X"E7",X"2A",X"12",X"E7",X"22",X"07",
		X"E7",X"21",X"02",X"E7",X"3E",X"01",X"BE",X"77",X"38",X"0D",X"3A",X"03",X"E7",X"A7",X"C0",X"3A",
		X"06",X"E7",X"3C",X"FE",X"04",X"38",X"02",X"3E",X"00",X"32",X"06",X"E7",X"3E",X"05",X"32",X"03",
		X"E7",X"C9",X"7E",X"FE",X"03",X"3E",X"05",X"20",X"02",X"3E",X"07",X"77",X"2A",X"12",X"E7",X"22",
		X"07",X"E7",X"C3",X"40",X"42",X"3E",X"01",X"32",X"03",X"E7",X"7E",X"FE",X"03",X"0E",X"04",X"3E",
		X"06",X"20",X"04",X"0E",X"06",X"3E",X"0B",X"71",X"32",X"06",X"E7",X"3E",X"FF",X"32",X"04",X"E7",
		X"2A",X"12",X"E7",X"22",X"07",X"E7",X"C9",X"7E",X"FE",X"02",X"28",X"19",X"FE",X"03",X"C8",X"36",
		X"02",X"2A",X"12",X"E7",X"22",X"07",X"E7",X"3E",X"02",X"32",X"03",X"E7",X"3A",X"01",X"E7",X"E6",
		X"FC",X"32",X"01",X"E7",X"C9",X"3A",X"03",X"E7",X"A7",X"C0",X"3E",X"03",X"32",X"02",X"E7",X"3E",
		X"05",X"32",X"06",X"E7",X"C9",X"3A",X"01",X"E7",X"E6",X"FC",X"32",X"01",X"E7",X"2A",X"12",X"E7",
		X"ED",X"5B",X"07",X"E7",X"3A",X"00",X"E7",X"E6",X"20",X"20",X"01",X"EB",X"ED",X"52",X"3E",X"08",
		X"11",X"00",X"04",X"ED",X"52",X"38",X"01",X"3C",X"32",X"02",X"E7",X"D6",X"08",X"87",X"06",X"00",
		X"4F",X"11",X"03",X"E7",X"21",X"A5",X"65",X"09",X"7E",X"23",X"66",X"6F",X"ED",X"A0",X"03",X"22",
		X"0C",X"E7",X"21",X"A9",X"65",X"09",X"7E",X"23",X"66",X"6F",X"ED",X"A0",X"22",X"0E",X"E7",X"AF",
		X"12",X"7E",X"32",X"06",X"E7",X"C9",X"21",X"1F",X"E7",X"CB",X"46",X"C2",X"4B",X"46",X"3A",X"1A",
		X"E7",X"A7",X"C2",X"56",X"46",X"2A",X"0C",X"E7",X"5E",X"23",X"56",X"E5",X"2A",X"10",X"E7",X"19",
		X"22",X"10",X"E7",X"E1",X"3A",X"03",X"E7",X"3D",X"20",X"06",X"23",X"7E",X"23",X"22",X"0C",X"E7",
		X"32",X"03",X"E7",X"2A",X"0E",X"E7",X"3A",X"04",X"E7",X"3D",X"20",X"09",X"23",X"7E",X"A7",X"28",
		X"2D",X"23",X"22",X"0E",X"E7",X"32",X"04",X"E7",X"4E",X"3A",X"05",X"E7",X"A7",X"28",X"58",X"2A",
		X"0A",X"E7",X"3A",X"05",X"E7",X"3D",X"20",X"2E",X"CB",X"7E",X"28",X"04",X"CB",X"79",X"20",X"29",
		X"23",X"7E",X"32",X"05",X"E7",X"23",X"A7",X"28",X"21",X"22",X"0A",X"E7",X"18",X"1B",X"21",X"00",
		X"05",X"22",X"02",X"E7",X"3E",X"04",X"32",X"06",X"E7",X"21",X"00",X"50",X"22",X"10",X"E7",X"2A",
		X"12",X"E7",X"22",X"07",X"E7",X"C9",X"32",X"05",X"E7",X"4E",X"3A",X"01",X"E7",X"CB",X"CF",X"CB",
		X"71",X"20",X"0A",X"CB",X"8F",X"CB",X"C7",X"CB",X"69",X"20",X"02",X"CB",X"87",X"32",X"01",X"E7",
		X"79",X"E6",X"1F",X"32",X"06",X"E7",X"C9",X"CB",X"79",X"28",X"F5",X"3A",X"09",X"E9",X"E6",X"30",
		X"28",X"EE",X"06",X"F8",X"CB",X"67",X"20",X"09",X"06",X"FB",X"3E",X"81",X"CD",X"FE",X"0D",X"18",
		X"03",X"CD",X"79",X"42",X"3A",X"02",X"E7",X"80",X"87",X"16",X"00",X"5F",X"21",X"AD",X"65",X"19",
		X"7E",X"23",X"66",X"6F",X"7E",X"32",X"05",X"E7",X"23",X"22",X"0A",X"E7",X"18",X"AB",X"3A",X"1F",
		X"E7",X"E6",X"01",X"20",X"75",X"21",X"03",X"E7",X"35",X"C0",X"21",X"02",X"E7",X"3A",X"06",X"E7",
		X"FE",X"05",X"36",X"03",X"C8",X"36",X"00",X"3E",X"00",X"32",X"06",X"E7",X"3E",X"05",X"32",X"03",
		X"E7",X"C9",X"21",X"03",X"E7",X"35",X"20",X"19",X"2A",X"0A",X"E7",X"7E",X"FE",X"FF",X"28",X"3B",
		X"32",X"06",X"E7",X"23",X"7E",X"23",X"32",X"03",X"E7",X"22",X"0A",X"E7",X"21",X"00",X"E7",X"CB",
		X"CE",X"ED",X"5B",X"0E",X"E7",X"2A",X"07",X"E7",X"19",X"22",X"0E",X"E7",X"2A",X"10",X"E7",X"ED",
		X"52",X"22",X"10",X"E7",X"2A",X"12",X"E7",X"ED",X"5B",X"0C",X"E7",X"3A",X"00",X"E7",X"E6",X"20",
		X"28",X"04",X"ED",X"52",X"18",X"01",X"19",X"22",X"12",X"E7",X"C9",X"3E",X"0B",X"32",X"00",X"E0",
		X"C9",X"7E",X"FE",X"06",X"3E",X"05",X"30",X"0C",X"18",X"07",X"3A",X"06",X"E7",X"FE",X"05",X"28",
		X"06",X"CD",X"8E",X"46",X"32",X"06",X"E7",X"CD",X"91",X"2E",X"2A",X"12",X"E7",X"22",X"07",X"E7",
		X"3A",X"01",X"E7",X"E6",X"FC",X"32",X"01",X"E7",X"21",X"1F",X"E7",X"CB",X"86",X"3E",X"08",X"32",
		X"03",X"E7",X"21",X"21",X"E7",X"3A",X"09",X"E7",X"A7",X"37",X"FA",X"91",X"45",X"96",X"32",X"09",
		X"E7",X"21",X"02",X"E7",X"36",X"0B",X"D0",X"CD",X"08",X"12",X"C0",X"34",X"3A",X"20",X"E7",X"A7",
		X"F5",X"3E",X"00",X"CD",X"FE",X"0D",X"3E",X"87",X"CD",X"FE",X"0D",X"F1",X"21",X"EC",X"45",X"11",
		X"0C",X"00",X"01",X"12",X"00",X"20",X"23",X"2A",X"12",X"E7",X"ED",X"5B",X"DA",X"E2",X"ED",X"52",
		X"21",X"01",X"E7",X"38",X"07",X"CB",X"B6",X"2B",X"CB",X"AE",X"18",X"05",X"CB",X"F6",X"2B",X"CB",
		X"EE",X"21",X"F1",X"45",X"11",X"39",X"00",X"01",X"1B",X"00",X"22",X"0A",X"E7",X"ED",X"53",X"0C",
		X"E7",X"ED",X"43",X"07",X"E7",X"21",X"00",X"00",X"22",X"0E",X"E7",X"C9",X"22",X"0A",X"23",X"18",
		X"FF",X"24",X"08",X"25",X"16",X"FF",X"21",X"1F",X"E7",X"CB",X"46",X"28",X"0C",X"CD",X"91",X"2E",
		X"CD",X"75",X"46",X"CD",X"8E",X"46",X"32",X"06",X"E7",X"ED",X"5B",X"0E",X"E7",X"21",X"12",X"00",
		X"19",X"22",X"0E",X"E7",X"2A",X"10",X"E7",X"ED",X"52",X"EB",X"21",X"00",X"B0",X"19",X"30",X"05",
		X"ED",X"53",X"10",X"E7",X"C9",X"21",X"00",X"50",X"21",X"1F",X"E7",X"CB",X"4E",X"28",X"14",X"CB",
		X"8E",X"CD",X"08",X"12",X"20",X"0D",X"3E",X"0C",X"32",X"02",X"E7",X"3E",X"05",X"32",X"03",X"E7",
		X"C3",X"9F",X"45",X"21",X"02",X"E7",X"36",X"00",X"C3",X"47",X"43",X"CD",X"91",X"2E",X"CD",X"75",
		X"46",X"CD",X"8E",X"46",X"18",X"02",X"3E",X"10",X"32",X"06",X"E7",X"3E",X"0D",X"32",X"02",X"E7",
		X"21",X"80",X"00",X"22",X"0E",X"E7",X"2A",X"12",X"E7",X"22",X"07",X"E7",X"3A",X"01",X"E7",X"E6",
		X"FC",X"32",X"01",X"E7",X"C9",X"21",X"21",X"E7",X"3A",X"09",X"E7",X"A7",X"FA",X"84",X"46",X"96",
		X"0E",X"00",X"30",X"02",X"0E",X"02",X"32",X"09",X"E7",X"21",X"1F",X"E7",X"71",X"C9",X"2A",X"10",
		X"E7",X"11",X"00",X"18",X"19",X"ED",X"5B",X"22",X"E7",X"ED",X"52",X"3E",X"20",X"D8",X"3C",X"C9",
		X"CD",X"03",X"59",X"FE",X"04",X"28",X"4D",X"21",X"03",X"E7",X"35",X"C0",X"36",X"08",X"21",X"05",
		X"E7",X"35",X"20",X"24",X"36",X"02",X"2B",X"35",X"28",X"34",X"2A",X"12",X"E7",X"11",X"00",X"01",
		X"3A",X"01",X"E1",X"A7",X"28",X"03",X"19",X"18",X"02",X"ED",X"52",X"22",X"12",X"E7",X"2A",X"10",
		X"E7",X"11",X"00",X"06",X"19",X"22",X"10",X"E7",X"3A",X"06",X"E7",X"3C",X"FE",X"20",X"20",X"02",
		X"3E",X"1C",X"32",X"06",X"E7",X"E6",X"01",X"C0",X"3E",X"90",X"CD",X"FE",X"0D",X"C9",X"3E",X"0C",
		X"32",X"00",X"E0",X"C9",X"3A",X"06",X"E7",X"FE",X"26",X"C0",X"3E",X"0C",X"32",X"00",X"E0",X"AF",
		X"32",X"40",X"E3",X"C9",X"2A",X"02",X"E1",X"ED",X"5B",X"12",X"E7",X"CD",X"03",X"59",X"FE",X"04",
		X"28",X"72",X"3A",X"01",X"E1",X"FE",X"01",X"FD",X"21",X"00",X"50",X"38",X"06",X"C0",X"FD",X"21",
		X"00",X"52",X"EB",X"A7",X"ED",X"52",X"D8",X"E5",X"2A",X"10",X"E7",X"11",X"00",X"50",X"ED",X"52",
		X"38",X"50",X"29",X"7C",X"E1",X"06",X"0C",X"D6",X"0C",X"38",X"0E",X"11",X"00",X"01",X"ED",X"52",
		X"D8",X"11",X"00",X"06",X"FD",X"19",X"05",X"18",X"EE",X"FD",X"22",X"10",X"E7",X"3E",X"00",X"CD",
		X"FE",X"0D",X"3E",X"03",X"32",X"00",X"E0",X"EB",X"2A",X"12",X"E7",X"3A",X"01",X"E1",X"A7",X"28",
		X"05",X"ED",X"52",X"11",X"00",X"01",X"19",X"22",X"12",X"E7",X"21",X"00",X"E7",X"CB",X"CE",X"3E",
		X"1C",X"32",X"06",X"E7",X"3E",X"08",X"32",X"03",X"E7",X"3E",X"01",X"32",X"05",X"E7",X"78",X"32",
		X"04",X"E7",X"F1",X"C9",X"ED",X"52",X"D8",X"3A",X"02",X"E7",X"FE",X"02",X"D0",X"21",X"41",X"E3",
		X"34",X"3E",X"05",X"32",X"46",X"E3",X"3E",X"05",X"32",X"47",X"E3",X"3E",X"03",X"21",X"01",X"E7",
		X"CB",X"B6",X"2B",X"CB",X"AE",X"CB",X"CE",X"32",X"00",X"E0",X"3E",X"00",X"CD",X"FE",X"0D",X"F1",
		X"3E",X"03",X"32",X"06",X"E7",X"C9",X"DD",X"21",X"4C",X"E3",X"DD",X"CB",X"00",X"66",X"C4",X"21",
		X"48",X"DD",X"21",X"40",X"E3",X"DD",X"4E",X"00",X"CB",X"61",X"C8",X"DD",X"7E",X"01",X"FE",X"01",
		X"38",X"39",X"28",X"13",X"11",X"1B",X"00",X"CD",X"EA",X"1B",X"11",X"20",X"FF",X"19",X"38",X"41",
		X"3E",X"26",X"32",X"06",X"E7",X"18",X"3A",X"DD",X"35",X"07",X"20",X"35",X"DD",X"36",X"07",X"0B",
		X"DD",X"34",X"06",X"DD",X"7E",X"06",X"FE",X"07",X"38",X"27",X"DD",X"36",X"07",X"07",X"DD",X"34",
		X"01",X"DD",X"36",X"06",X"01",X"DD",X"CB",X"0C",X"E6",X"18",X"16",X"DD",X"35",X"07",X"20",X"11",
		X"DD",X"36",X"07",X"08",X"DD",X"7E",X"06",X"3C",X"FE",X"05",X"28",X"02",X"3E",X"04",X"DD",X"77",
		X"06",X"CD",X"E2",X"1B",X"11",X"00",X"EE",X"19",X"D8",X"21",X"F0",X"73",X"C3",X"7D",X"1A",X"3A",
		X"00",X"E0",X"FE",X"06",X"20",X"17",X"21",X"22",X"E0",X"35",X"C0",X"EB",X"2A",X"23",X"E0",X"7E",
		X"FE",X"FF",X"28",X"34",X"23",X"12",X"7E",X"23",X"22",X"23",X"E0",X"18",X"27",X"3A",X"06",X"E9",
		X"E6",X"04",X"21",X"00",X"E7",X"CB",X"46",X"20",X"1B",X"3A",X"06",X"E9",X"E6",X"07",X"4F",X"3A",
		X"1A",X"E7",X"A7",X"79",X"20",X"0E",X"3A",X"08",X"E9",X"2F",X"47",X"2F",X"07",X"07",X"07",X"A0",
		X"E6",X"38",X"47",X"B1",X"32",X"09",X"E9",X"C9",X"3E",X"0B",X"32",X"00",X"E0",X"C9",X"F3",X"31",
		X"00",X"F0",X"AF",X"32",X"01",X"E0",X"32",X"20",X"E0",X"32",X"21",X"E0",X"32",X"80",X"E0",X"FB",
		X"CD",X"00",X"57",X"CD",X"4A",X"06",X"21",X"6D",X"4B",X"CD",X"1C",X"11",X"21",X"01",X"4F",X"22",
		X"0E",X"E7",X"3E",X"9C",X"32",X"05",X"E7",X"21",X"A0",X"30",X"22",X"12",X"E7",X"21",X"00",X"5C",
		X"22",X"10",X"E7",X"22",X"44",X"E3",X"21",X"A0",X"34",X"22",X"42",X"E3",X"3E",X"10",X"32",X"40",
		X"E3",X"3E",X"05",X"32",X"47",X"E3",X"DD",X"21",X"62",X"E2",X"01",X"50",X"07",X"21",X"00",X"0F",
		X"06",X"07",X"DD",X"36",X"04",X"00",X"DD",X"36",X"05",X"5C",X"DD",X"36",X"07",X"07",X"DD",X"36",
		X"0E",X"38",X"DD",X"70",X"0F",X"DD",X"71",X"00",X"DD",X"75",X"02",X"DD",X"74",X"03",X"78",X"FE",
		X"07",X"28",X"08",X"FE",X"04",X"38",X"04",X"DD",X"36",X"06",X"0A",X"FE",X"05",X"30",X"05",X"21",
		X"00",X"31",X"0E",X"10",X"11",X"10",X"00",X"DD",X"19",X"10",X"C7",X"3E",X"05",X"32",X"00",X"E0",
		X"11",X"52",X"D1",X"0E",X"0B",X"21",X"86",X"4B",X"CD",X"34",X"11",X"3A",X"20",X"E0",X"FE",X"08",
		X"20",X"F9",X"CD",X"1C",X"11",X"3A",X"20",X"E0",X"FE",X"0B",X"20",X"F9",X"CD",X"AE",X"49",X"21",
		X"0E",X"4C",X"CD",X"34",X"11",X"3E",X"E1",X"CD",X"0F",X"57",X"CD",X"AE",X"49",X"21",X"71",X"4C",
		X"CD",X"1C",X"11",X"CD",X"C0",X"49",X"3A",X"00",X"E0",X"FE",X"0B",X"20",X"F6",X"AF",X"21",X"00",
		X"00",X"32",X"81",X"E0",X"22",X"82",X"E0",X"3C",X"32",X"84",X"E0",X"32",X"22",X"E0",X"21",X"25",
		X"E0",X"7E",X"36",X"09",X"11",X"55",X"4A",X"A7",X"28",X"05",X"11",X"0A",X"4B",X"36",X"00",X"32",
		X"80",X"E0",X"ED",X"53",X"23",X"E0",X"CD",X"57",X"11",X"3E",X"01",X"CD",X"49",X"04",X"F3",X"3E",
		X"06",X"32",X"00",X"E0",X"21",X"00",X"00",X"22",X"81",X"E0",X"22",X"82",X"E0",X"22",X"10",X"E0",
		X"22",X"12",X"E0",X"FB",X"CD",X"B8",X"0F",X"3A",X"00",X"E0",X"FE",X"0B",X"20",X"F6",X"3E",X"38",
		X"CD",X"0F",X"57",X"CD",X"20",X"56",X"3E",X"E1",X"CD",X"0F",X"57",X"C3",X"7E",X"48",X"11",X"50",
		X"D1",X"06",X"04",X"D5",X"CD",X"2A",X"57",X"E1",X"11",X"80",X"00",X"19",X"EB",X"10",X"F4",X"C9",
		X"11",X"16",X"D3",X"01",X"0B",X"19",X"3A",X"80",X"E8",X"E6",X"30",X"CA",X"1F",X"57",X"2A",X"0A",
		X"E9",X"7D",X"AC",X"20",X"14",X"13",X"CD",X"F7",X"49",X"CB",X"5D",X"C0",X"11",X"97",X"D3",X"7D",
		X"87",X"27",X"CD",X"10",X"4A",X"3E",X"02",X"18",X"21",X"3E",X"41",X"CD",X"F4",X"49",X"6C",X"11",
		X"96",X"D3",X"3E",X"42",X"CD",X"2C",X"4A",X"CB",X"5D",X"3E",X"01",X"20",X"01",X"7D",X"CD",X"10",
		X"4A",X"CB",X"5D",X"3E",X"01",X"28",X"03",X"7D",X"E6",X"07",X"E5",X"21",X"39",X"4A",X"18",X"04",
		X"E5",X"21",X"34",X"4A",X"F5",X"C5",X"48",X"CD",X"F7",X"56",X"C1",X"13",X"CD",X"1C",X"11",X"F1",
		X"D5",X"FE",X"01",X"3E",X"53",X"C4",X"10",X"11",X"D1",X"13",X"E1",X"C9",X"CD",X"10",X"11",X"3E",
		X"2D",X"C3",X"10",X"11",X"43",X"4F",X"49",X"4E",X"FF",X"50",X"4C",X"41",X"59",X"45",X"52",X"FF",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"FF",X"42",X"02",X"01",X"20",X"28",X"02",X"02",X"10",X"18",X"02",X"03",
		X"10",X"18",X"02",X"02",X"10",X"24",X"02",X"02",X"20",X"38",X"02",X"10",X"04",X"02",X"20",X"1E",
		X"02",X"10",X"08",X"02",X"20",X"2C",X"01",X"04",X"20",X"28",X"02",X"08",X"01",X"02",X"10",X"28",
		X"01",X"10",X"08",X"18",X"20",X"08",X"01",X"40",X"02",X"08",X"08",X"08",X"20",X"48",X"02",X"03",
		X"01",X"03",X"02",X"03",X"01",X"03",X"06",X"03",X"05",X"03",X"06",X"03",X"01",X"03",X"02",X"03",
		X"01",X"03",X"01",X"03",X"02",X"03",X"01",X"03",X"06",X"03",X"05",X"03",X"06",X"03",X"01",X"03",
		X"02",X"03",X"01",X"03",X"02",X"03",X"01",X"03",X"06",X"03",X"05",X"03",X"06",X"03",X"01",X"18",
		X"02",X"02",X"08",X"48",X"02",X"02",X"10",X"18",X"00",X"02",X"10",X"18",X"00",X"0A",X"01",X"0A",
		X"04",X"02",X"10",X"18",X"04",X"02",X"20",X"18",X"04",X"02",X"10",X"10",X"04",X"28",X"01",X"03",
		X"20",X"20",X"01",X"03",X"20",X"18",X"01",X"03",X"20",X"08",X"00",X"28",X"02",X"08",X"04",X"03",
		X"20",X"10",X"10",X"34",X"02",X"04",X"08",X"10",X"20",X"28",X"02",X"05",X"01",X"05",X"02",X"05",
		X"01",X"05",X"06",X"05",X"05",X"05",X"06",X"80",X"00",X"FF",X"1C",X"01",X"04",X"00",X"01",X"10",
		X"44",X"01",X"10",X"00",X"28",X"01",X"02",X"20",X"10",X"02",X"20",X"01",X"02",X"08",X"50",X"01",
		X"02",X"08",X"36",X"01",X"0A",X"02",X"30",X"00",X"10",X"10",X"20",X"00",X"1B",X"02",X"02",X"08",
		X"10",X"10",X"48",X"02",X"02",X"08",X"10",X"20",X"28",X"04",X"02",X"20",X"20",X"04",X"68",X"01",
		X"0A",X"00",X"04",X"20",X"10",X"02",X"10",X"00",X"28",X"01",X"01",X"02",X"60",X"04",X"38",X"01",
		X"02",X"08",X"10",X"10",X"30",X"00",X"50",X"01",X"20",X"02",X"02",X"08",X"10",X"20",X"20",X"00",
		X"18",X"02",X"10",X"08",X"10",X"20",X"10",X"00",X"40",X"01",X"A0",X"04",X"FF",X"FE",X"1D",X"FD",
		X"D8",X"D6",X"40",X"20",X"31",X"39",X"38",X"34",X"20",X"FE",X"DA",X"49",X"52",X"45",X"4D",X"20",
		X"43",X"4F",X"52",X"50",X"2E",X"FF",X"41",X"20",X"4B",X"55",X"4E",X"47",X"2D",X"46",X"55",X"20",
		X"4D",X"41",X"53",X"54",X"45",X"52",X"2C",X"FE",X"1A",X"54",X"48",X"4F",X"4D",X"41",X"53",X"FE",
		X"0B",X"20",X"41",X"4E",X"44",X"20",X"FD",X"D2",X"D1",X"FE",X"1A",X"53",X"49",X"4C",X"56",X"49",
		X"41",X"FE",X"0B",X"20",X"57",X"45",X"52",X"45",X"20",X"53",X"55",X"44",X"44",X"45",X"4E",X"4C",
		X"59",X"20",X"41",X"54",X"54",X"41",X"43",X"4B",X"45",X"44",X"20",X"FD",X"52",X"D2",X"42",X"59",
		X"20",X"53",X"45",X"56",X"45",X"52",X"41",X"4C",X"20",X"55",X"4E",X"4B",X"4E",X"4F",X"57",X"4E",
		X"20",X"47",X"55",X"59",X"53",X"2E",X"FF",X"FD",X"D0",X"D2",X"28",X"FE",X"1A",X"53",X"49",X"4C",
		X"56",X"49",X"41",X"FE",X"0B",X"20",X"57",X"41",X"53",X"20",X"4B",X"49",X"44",X"4E",X"41",X"50",
		X"50",X"45",X"44",X"20",X"42",X"59",X"20",X"54",X"48",X"45",X"4D",X"2E",X"29",X"FF",X"FD",X"53",
		X"D1",X"4C",X"41",X"54",X"45",X"52",X"20",X"FE",X"1A",X"54",X"48",X"4F",X"4D",X"41",X"53",X"FE",
		X"0B",X"20",X"46",X"4F",X"55",X"4E",X"44",X"20",X"41",X"20",X"4C",X"45",X"54",X"54",X"45",X"52",
		X"20",X"FD",X"D3",X"D1",X"46",X"52",X"4F",X"4D",X"20",X"FE",X"1A",X"58",X"FE",X"0B",X"2E",X"20",
		X"FD",X"53",X"D2",X"48",X"45",X"20",X"49",X"53",X"20",X"41",X"4E",X"20",X"49",X"4E",X"48",X"41",
		X"42",X"49",X"54",X"41",X"4E",X"54",X"20",X"4F",X"46",X"20",X"54",X"48",X"45",X"20",X"FD",X"D3",
		X"D2",X"44",X"45",X"56",X"49",X"4C",X"27",X"53",X"20",X"54",X"45",X"4D",X"50",X"4C",X"45",X"2E",
		X"FF",X"FE",X"DA",X"FD",X"DA",X"D0",X"80",X"81",X"82",X"83",X"84",X"85",X"86",X"87",X"88",X"89",
		X"8A",X"FD",X"1A",X"D1",X"8B",X"8C",X"8D",X"8E",X"8F",X"90",X"91",X"92",X"93",X"94",X"95",X"FD",
		X"57",X"D1",X"96",X"97",X"98",X"99",X"9A",X"9B",X"9C",X"9D",X"9E",X"9F",X"A0",X"A1",X"A2",X"A3",
		X"A4",X"A5",X"A4",X"A6",X"FD",X"96",X"D1",X"A7",X"A8",X"A9",X"AA",X"AB",X"AC",X"AD",X"AE",X"AF",
		X"B0",X"B1",X"B2",X"B3",X"B4",X"B5",X"B6",X"B7",X"B3",X"B8",X"B9",X"FD",X"D6",X"D1",X"BA",X"BB",
		X"BC",X"BD",X"BE",X"BF",X"C0",X"C1",X"C2",X"C3",X"C4",X"C5",X"C6",X"C7",X"C8",X"C9",X"CA",X"CB",
		X"CC",X"CD",X"FD",X"15",X"D2",X"CE",X"CF",X"D0",X"D1",X"D2",X"D3",X"D4",X"D5",X"D6",X"D7",X"D8",
		X"D9",X"06",X"DA",X"DB",X"DC",X"DD",X"DE",X"DF",X"E0",X"E1",X"FD",X"55",X"D2",X"E2",X"E3",X"E4",
		X"E5",X"E6",X"E7",X"E8",X"E9",X"EA",X"EB",X"EC",X"ED",X"06",X"EE",X"EF",X"F0",X"F1",X"06",X"F2",
		X"F3",X"F4",X"F5",X"FD",X"95",X"D2",X"F6",X"F7",X"F8",X"F9",X"FA",X"FB",X"70",X"71",X"72",X"73",
		X"74",X"75",X"06",X"76",X"77",X"78",X"79",X"7A",X"7B",X"7C",X"7D",X"7E",X"FF",X"3E",X"0B",X"32",
		X"00",X"E0",X"18",X"30",X"21",X"03",X"E7",X"7E",X"A7",X"28",X"01",X"35",X"21",X"05",X"E7",X"35",
		X"20",X"4D",X"ED",X"5B",X"0E",X"E7",X"1A",X"A7",X"FA",X"1D",X"4D",X"CB",X"77",X"28",X"04",X"21",
		X"20",X"E0",X"34",X"CB",X"6F",X"28",X"0D",X"F5",X"21",X"B7",X"65",X"7E",X"23",X"22",X"0C",X"E7",
		X"32",X"03",X"E7",X"F1",X"6F",X"CB",X"65",X"28",X"05",X"3E",X"02",X"32",X"03",X"E7",X"CB",X"5D",
		X"28",X"08",X"3A",X"01",X"E7",X"EE",X"40",X"32",X"01",X"E7",X"7D",X"E6",X"03",X"32",X"21",X"E0",
		X"13",X"1A",X"32",X"05",X"E7",X"13",X"1A",X"32",X"06",X"E7",X"13",X"ED",X"53",X"0E",X"E7",X"3A",
		X"21",X"E0",X"21",X"BC",X"4D",X"CD",X"26",X"1F",X"3A",X"20",X"E0",X"DD",X"21",X"40",X"E3",X"DD",
		X"4E",X"00",X"FE",X"0A",X"28",X"0A",X"30",X"11",X"A7",X"20",X"0B",X"CD",X"D4",X"47",X"18",X"09",
		X"11",X"36",X"00",X"CD",X"7A",X"1C",X"CD",X"21",X"48",X"3A",X"20",X"E0",X"DD",X"21",X"62",X"E2",
		X"DD",X"4E",X"00",X"21",X"C2",X"4D",X"CD",X"26",X"1F",X"C3",X"72",X"2D",X"FA",X"4D",X"12",X"4E",
		X"DA",X"4D",X"24",X"4E",X"25",X"4E",X"3A",X"4E",X"71",X"4E",X"AF",X"4E",X"A8",X"4E",X"A1",X"4E",
		X"9A",X"4E",X"93",X"4E",X"8C",X"4E",X"7F",X"4E",X"24",X"4E",X"2A",X"0C",X"E7",X"5E",X"23",X"56",
		X"E5",X"2A",X"10",X"E7",X"19",X"22",X"10",X"E7",X"E1",X"3A",X"03",X"E7",X"A7",X"20",X"23",X"23",
		X"7E",X"23",X"22",X"0C",X"E7",X"32",X"03",X"E7",X"18",X"18",X"CD",X"1F",X"43",X"2A",X"12",X"E7",
		X"11",X"E5",X"FF",X"3A",X"01",X"E7",X"E6",X"40",X"20",X"03",X"19",X"18",X"02",X"ED",X"52",X"22",
		X"12",X"E7",X"2A",X"12",X"E7",X"AF",X"29",X"17",X"29",X"17",X"29",X"17",X"6C",X"67",X"CD",X"D6",
		X"40",X"CD",X"E5",X"40",X"C9",X"CD",X"E7",X"1B",X"2A",X"64",X"E2",X"11",X"00",X"E7",X"19",X"30",
		X"3A",X"21",X"20",X"E0",X"34",X"21",X"E5",X"4E",X"18",X"09",X"21",X"69",X"E2",X"35",X"20",X"28",
		X"2A",X"6E",X"E2",X"7E",X"FE",X"FF",X"28",X"2E",X"32",X"68",X"E2",X"23",X"7E",X"32",X"69",X"E2",
		X"23",X"7E",X"A7",X"28",X"0F",X"E5",X"21",X"2B",X"E3",X"36",X"01",X"23",X"77",X"23",X"36",X"40",
		X"23",X"36",X"1A",X"E1",X"23",X"22",X"6E",X"E2",X"CD",X"E2",X"1B",X"CB",X"61",X"C2",X"72",X"1A",
		X"C9",X"CD",X"DF",X"4E",X"18",X"F5",X"21",X"20",X"E0",X"34",X"CD",X"DF",X"17",X"18",X"E9",X"21",
		X"A2",X"E2",X"11",X"10",X"00",X"06",X"03",X"CB",X"F6",X"19",X"10",X"FB",X"DD",X"21",X"C2",X"E2",
		X"CD",X"D7",X"4E",X"DD",X"21",X"B2",X"E2",X"CD",X"D7",X"4E",X"DD",X"21",X"A2",X"E2",X"CD",X"D7",
		X"4E",X"DD",X"21",X"82",X"E2",X"CD",X"B3",X"4E",X"DD",X"21",X"92",X"E2",X"CD",X"B3",X"4E",X"DD",
		X"21",X"72",X"E2",X"DD",X"4E",X"00",X"21",X"D1",X"4E",X"E5",X"DD",X"7E",X"01",X"FE",X"01",X"28",
		X"1E",X"CD",X"A8",X"15",X"DD",X"35",X"0E",X"C0",X"DD",X"7E",X"0F",X"DD",X"77",X"06",X"C3",X"DF",
		X"17",X"CB",X"61",X"C8",X"C3",X"2F",X"16",X"DD",X"4E",X"00",X"CD",X"E7",X"1B",X"18",X"F2",X"CB",
		X"61",X"C2",X"AA",X"1B",X"C9",X"0B",X"0B",X"00",X"0C",X"38",X"52",X"00",X"0B",X"00",X"09",X"0B",
		X"00",X"0A",X"38",X"50",X"00",X"2B",X"00",X"06",X"0A",X"00",X"00",X"18",X"00",X"06",X"01",X"00",
		X"FF",X"41",X"16",X"00",X"01",X"32",X"04",X"01",X"1C",X"05",X"01",X"2D",X"04",X"22",X"04",X"10",
		X"02",X"06",X"12",X"02",X"10",X"13",X"02",X"06",X"14",X"02",X"04",X"10",X"10",X"21",X"00",X"01",
		X"0B",X"04",X"22",X"04",X"10",X"02",X"06",X"12",X"02",X"10",X"18",X"02",X"06",X"14",X"02",X"04",
		X"10",X"01",X"08",X"06",X"01",X"08",X"07",X"01",X"08",X"06",X"01",X"13",X"04",X"41",X"21",X"04",
		X"41",X"0E",X"04",X"01",X"08",X"08",X"01",X"08",X"09",X"01",X"02",X"08",X"41",X"05",X"08",X"41",
		X"08",X"05",X"41",X"08",X"0B",X"41",X"08",X"0C",X"01",X"08",X"0B",X"01",X"08",X"05",X"01",X"08",
		X"0D",X"01",X"08",X"0E",X"01",X"09",X"0D",X"41",X"08",X"05",X"01",X"1C",X"04",X"09",X"10",X"00",
		X"10",X"27",X"00",X"41",X"E1",X"03",X"01",X"A9",X"03",X"01",X"16",X"04",X"01",X"08",X"06",X"01",
		X"08",X"07",X"01",X"08",X"06",X"01",X"08",X"04",X"01",X"08",X"08",X"01",X"08",X"09",X"01",X"08",
		X"08",X"09",X"08",X"04",X"01",X"08",X"06",X"01",X"08",X"07",X"01",X"08",X"06",X"01",X"08",X"04",
		X"01",X"08",X"05",X"01",X"08",X"0B",X"01",X"08",X"0C",X"01",X"08",X"0B",X"01",X"08",X"05",X"01",
		X"08",X"04",X"01",X"08",X"08",X"01",X"08",X"09",X"01",X"08",X"08",X"09",X"08",X"05",X"01",X"08",
		X"0B",X"01",X"08",X"0C",X"01",X"08",X"0B",X"01",X"08",X"05",X"22",X"04",X"10",X"02",X"06",X"12",
		X"02",X"10",X"18",X"02",X"06",X"14",X"02",X"04",X"10",X"09",X"08",X"04",X"01",X"08",X"06",X"01",
		X"08",X"07",X"01",X"08",X"06",X"01",X"A9",X"04",X"FF",X"3E",X"23",X"CD",X"FE",X"0D",X"AF",X"32",
		X"02",X"E7",X"32",X"20",X"E0",X"32",X"83",X"E8",X"3E",X"08",X"32",X"00",X"E0",X"CD",X"95",X"50",
		X"0E",X"D9",X"21",X"32",X"51",X"CD",X"1C",X"11",X"21",X"47",X"51",X"CD",X"1C",X"11",X"21",X"57",
		X"51",X"CD",X"1C",X"11",X"21",X"62",X"51",X"CD",X"1C",X"11",X"21",X"6D",X"51",X"CD",X"1C",X"11",
		X"21",X"A7",X"50",X"CD",X"79",X"50",X"3E",X"F8",X"CD",X"38",X"50",X"CD",X"91",X"50",X"21",X"FF",
		X"50",X"0E",X"D9",X"CD",X"79",X"50",X"3E",X"F8",X"E5",X"C5",X"D5",X"32",X"82",X"E8",X"0E",X"D9",
		X"21",X"83",X"E8",X"7E",X"A7",X"20",X"1A",X"36",X"0B",X"21",X"20",X"E0",X"35",X"35",X"F2",X"53",
		X"50",X"36",X"08",X"5E",X"16",X"00",X"21",X"6B",X"50",X"19",X"7E",X"23",X"66",X"6F",X"CD",X"1C",
		X"11",X"3A",X"82",X"E8",X"A7",X"20",X"D9",X"D1",X"C1",X"E1",X"C9",X"5D",X"51",X"68",X"51",X"4D",
		X"51",X"2D",X"51",X"3D",X"51",X"5E",X"23",X"56",X"23",X"7E",X"23",X"3C",X"C8",X"3C",X"3C",X"28",
		X"F4",X"D6",X"03",X"CD",X"10",X"11",X"FE",X"20",X"20",X"EF",X"3E",X"0B",X"CD",X"38",X"50",X"18",
		X"E8",X"06",X"08",X"18",X"02",X"06",X"19",X"0E",X"0B",X"11",X"9F",X"D1",X"CD",X"1A",X"57",X"21",
		X"1F",X"00",X"19",X"EB",X"10",X"F6",X"C9",X"FD",X"63",X"D2",X"41",X"20",X"4B",X"55",X"4E",X"47",
		X"2D",X"46",X"55",X"20",X"4D",X"41",X"53",X"54",X"45",X"52",X"2C",X"54",X"48",X"4F",X"4D",X"41",
		X"53",X"20",X"41",X"4E",X"44",X"20",X"FD",X"E3",X"D2",X"53",X"49",X"4C",X"56",X"49",X"41",X"20",
		X"45",X"4E",X"4A",X"4F",X"59",X"45",X"44",X"20",X"48",X"41",X"50",X"50",X"49",X"4E",X"45",X"53",
		X"53",X"20",X"FD",X"63",X"D3",X"41",X"47",X"41",X"49",X"4E",X"20",X"46",X"4F",X"52",X"20",X"41",
		X"20",X"4C",X"49",X"54",X"54",X"4C",X"45",X"20",X"57",X"48",X"49",X"4C",X"45",X"2E",X"FF",X"FD",
		X"A6",X"D2",X"42",X"55",X"54",X"20",X"54",X"48",X"45",X"49",X"52",X"20",X"48",X"41",X"50",X"50",
		X"59",X"20",X"44",X"41",X"59",X"53",X"20",X"FD",X"28",X"D3",X"44",X"49",X"44",X"20",X"4E",X"4F",
		X"54",X"20",X"4C",X"41",X"53",X"54",X"20",X"4C",X"4F",X"4E",X"47",X"2E",X"FF",X"FD",X"2E",X"D4",
		X"00",X"00",X"FD",X"AC",X"D4",X"60",X"61",X"FD",X"EC",X"D4",X"62",X"63",X"FF",X"FD",X"AC",X"D4",
		X"00",X"00",X"FD",X"EC",X"D4",X"00",X"00",X"FD",X"6D",X"D4",X"64",X"65",X"FF",X"FD",X"B0",X"D4",
		X"00",X"00",X"FD",X"F0",X"D4",X"00",X"00",X"FD",X"2E",X"D4",X"66",X"67",X"FF",X"FD",X"6D",X"D4",
		X"00",X"00",X"FD",X"6F",X"D4",X"68",X"69",X"FF",X"FD",X"6F",X"D4",X"00",X"00",X"FD",X"B0",X"D4",
		X"6A",X"6B",X"FD",X"F0",X"D4",X"6C",X"6D",X"FF",X"21",X"05",X"E0",X"CB",X"FE",X"CD",X"57",X"11",
		X"CD",X"03",X"57",X"11",X"5A",X"D2",X"0E",X"14",X"3A",X"80",X"E8",X"E6",X"18",X"28",X"08",X"21",
		X"D8",X"51",X"CD",X"1C",X"11",X"18",X"03",X"CD",X"25",X"57",X"11",X"19",X"D3",X"3A",X"13",X"E9",
		X"F5",X"FE",X"01",X"21",X"E5",X"51",X"28",X"03",X"21",X"F3",X"51",X"CD",X"1C",X"11",X"21",X"02",
		X"52",X"CD",X"1C",X"11",X"F1",X"CD",X"FF",X"10",X"3A",X"04",X"E9",X"E6",X"03",X"28",X"C4",X"E6",
		X"02",X"32",X"02",X"E0",X"06",X"01",X"28",X"01",X"04",X"21",X"13",X"E9",X"7E",X"90",X"38",X"B3",
		X"27",X"77",X"21",X"05",X"E0",X"CB",X"BE",X"C9",X"50",X"55",X"53",X"48",X"20",X"20",X"42",X"55",
		X"54",X"54",X"4F",X"4E",X"FF",X"4F",X"4E",X"4C",X"59",X"20",X"31",X"20",X"50",X"4C",X"41",X"59",
		X"45",X"52",X"FF",X"31",X"20",X"4F",X"52",X"20",X"32",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",
		X"53",X"FF",X"FD",X"E1",X"D5",X"43",X"52",X"45",X"44",X"49",X"54",X"20",X"FF",X"CD",X"57",X"11",
		X"CD",X"03",X"57",X"3E",X"20",X"CD",X"FE",X"0D",X"0E",X"1B",X"11",X"53",X"D1",X"06",X"17",X"CD",
		X"25",X"57",X"21",X"26",X"00",X"19",X"EB",X"10",X"F6",X"21",X"32",X"52",X"CD",X"39",X"57",X"C3",
		X"1C",X"11",X"FD",X"55",X"D1",X"CC",X"FD",X"60",X"D1",X"CC",X"FD",X"67",X"D1",X"CC",X"FD",X"92",
		X"D3",X"E3",X"FD",X"D1",X"D3",X"D9",X"D8",X"00",X"D0",X"D1",X"CD",X"FD",X"10",X"D4",X"E0",X"DB",
		X"DA",X"00",X"D2",X"D3",X"CF",X"FD",X"50",X"D4",X"E2",X"07",X"DC",X"DD",X"D4",X"D5",X"FD",X"90",
		X"D4",X"E4",X"07",X"DE",X"DF",X"D6",X"D7",X"FD",X"D0",X"D4",X"E6",X"07",X"07",X"07",X"E5",X"FD",
		X"10",X"D5",X"E1",X"07",X"E8",X"E9",X"E7",X"FD",X"50",X"D5",X"07",X"07",X"EA",X"EB",X"FD",X"90",
		X"D5",X"07",X"07",X"EC",X"ED",X"FD",X"D0",X"D5",X"07",X"EF",X"EE",X"FD",X"10",X"D6",X"07",X"F1",
		X"FD",X"50",X"D6",X"F0",X"F3",X"FD",X"90",X"D6",X"F2",X"FD",X"D0",X"D6",X"F4",X"FD",X"D6",X"D6",
		X"CE",X"FD",X"E4",X"D6",X"CE",X"FE",X"FD",X"AD",X"D3",X"E3",X"FD",X"E9",X"D3",X"CD",X"D1",X"D0",
		X"00",X"D8",X"D9",X"FD",X"29",X"D4",X"CF",X"D3",X"D2",X"00",X"DA",X"DB",X"E0",X"FD",X"6A",X"D4",
		X"D5",X"D4",X"DD",X"DC",X"07",X"E2",X"FD",X"AA",X"D4",X"D7",X"D6",X"DF",X"DE",X"07",X"E4",X"FD",
		X"EB",X"D4",X"E5",X"07",X"07",X"07",X"E6",X"FD",X"2B",X"D5",X"E7",X"E9",X"E8",X"07",X"E1",X"FD",
		X"6C",X"D5",X"EB",X"EA",X"07",X"07",X"FD",X"AC",X"D5",X"ED",X"EC",X"07",X"07",X"FD",X"ED",X"D5",
		X"EE",X"EF",X"07",X"FD",X"2E",X"D6",X"F1",X"07",X"FD",X"6E",X"D6",X"F3",X"F0",X"FD",X"AF",X"D6",
		X"F2",X"FD",X"EF",X"D6",X"F4",X"FF",X"FE",X"1B",X"FD",X"17",X"D2",X"59",X"4F",X"55",X"52",X"20",
		X"4C",X"4F",X"56",X"45",X"20",X"FE",X"1F",X"53",X"49",X"4C",X"56",X"49",X"41",X"FE",X"1B",X"FD",
		X"97",X"D2",X"49",X"53",X"20",X"49",X"4E",X"20",X"43",X"55",X"53",X"54",X"4F",X"44",X"59",X"20",
		X"4E",X"4F",X"57",X"2E",X"FD",X"16",X"D3",X"49",X"46",X"20",X"59",X"4F",X"55",X"20",X"57",X"41",
		X"4E",X"54",X"20",X"54",X"4F",X"20",X"53",X"41",X"56",X"45",X"FD",X"97",X"D3",X"59",X"4F",X"55",
		X"52",X"20",X"44",X"45",X"41",X"52",X"20",X"FE",X"1F",X"53",X"49",X"4C",X"56",X"49",X"41",X"27",
		X"53",X"FD",X"19",X"D4",X"FE",X"1F",X"4C",X"49",X"46",X"45",X"FE",X"1B",X"2C",X"20",X"43",X"4F",
		X"4D",X"45",X"20",X"54",X"4F",X"FD",X"97",X"D4",X"54",X"48",X"45",X"20",X"44",X"45",X"56",X"49",
		X"4C",X"27",X"53",X"20",X"54",X"45",X"4D",X"50",X"4C",X"45",X"FD",X"17",X"D5",X"41",X"54",X"20",
		X"4F",X"4E",X"43",X"45",X"2E",X"FD",X"96",X"D5",X"35",X"20",X"53",X"4F",X"4E",X"53",X"20",X"4F",
		X"46",X"20",X"54",X"48",X"45",X"20",X"44",X"45",X"56",X"49",X"4C",X"FD",X"17",X"D6",X"57",X"49",
		X"4C",X"4C",X"20",X"45",X"4E",X"54",X"45",X"52",X"54",X"41",X"49",X"4E",X"20",X"59",X"4F",X"55",
		X"2E",X"FF",X"CD",X"00",X"57",X"3E",X"05",X"CD",X"FE",X"0D",X"3A",X"80",X"E0",X"F5",X"3E",X"04",
		X"32",X"80",X"E0",X"CD",X"4A",X"06",X"21",X"00",X"54",X"22",X"10",X"E7",X"22",X"44",X"E3",X"21",
		X"00",X"27",X"22",X"12",X"E7",X"21",X"00",X"1A",X"22",X"42",X"E3",X"F1",X"32",X"80",X"E0",X"21",
		X"47",X"54",X"CD",X"1C",X"11",X"3E",X"07",X"32",X"00",X"E0",X"3E",X"70",X"CD",X"16",X"54",X"21",
		X"AB",X"54",X"CD",X"1C",X"11",X"3E",X"05",X"CD",X"FE",X"0D",X"3E",X"70",X"CD",X"16",X"54",X"3E",
		X"05",X"CD",X"FE",X"0D",X"3E",X"C0",X"32",X"82",X"E8",X"3A",X"80",X"E8",X"11",X"95",X"D2",X"0E",
		X"D9",X"21",X"85",X"54",X"E6",X"18",X"20",X"03",X"21",X"98",X"54",X"CD",X"1C",X"11",X"21",X"82",
		X"E8",X"7E",X"A7",X"20",X"E4",X"C9",X"21",X"03",X"E7",X"7E",X"A7",X"28",X"01",X"35",X"CD",X"1F",
		X"43",X"CD",X"12",X"4E",X"C3",X"B6",X"47",X"FE",X"96",X"FD",X"18",X"D5",X"B7",X"FD",X"57",X"D5",
		X"AA",X"AB",X"FD",X"97",X"D5",X"AC",X"AD",X"FD",X"D7",X"D5",X"F6",X"F5",X"FC",X"FD",X"17",X"D6",
		X"F8",X"F9",X"F7",X"FD",X"57",X"D6",X"FA",X"FB",X"FE",X"D6",X"18",X"FD",X"56",X"D1",X"FE",X"D7",
		X"4C",X"45",X"54",X"27",X"53",X"20",X"54",X"52",X"59",X"20",X"4E",X"45",X"58",X"54",X"20",X"46",
		X"4C",X"4F",X"4F",X"52",X"FF",X"48",X"45",X"4C",X"50",X"20",X"4D",X"45",X"2C",X"FD",X"15",X"D3",
		X"54",X"48",X"4F",X"4D",X"41",X"53",X"21",X"FF",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"FD",X"15",X"D3",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"FF",X"FE",X"DA",X"FD",X"A3",X"D2",
		X"49",X"27",X"4D",X"20",X"43",X"4F",X"4D",X"49",X"4E",X"47",X"FD",X"23",X"D3",X"52",X"49",X"47",
		X"48",X"54",X"20",X"41",X"57",X"41",X"59",X"2C",X"FD",X"A5",X"D3",X"53",X"49",X"4C",X"56",X"49",
		X"41",X"21",X"FF",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"47",
		X"41",X"4D",X"45",X"20",X"4F",X"56",X"45",X"52",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"3E",X"21",X"CD",X"FE",X"0D",X"11",X"40",X"D3",X"0E",X"DB",X"DD",X"21",
		X"D3",X"54",X"CD",X"C3",X"56",X"3E",X"E1",X"CD",X"0F",X"57",X"3E",X"38",X"CD",X"0F",X"57",X"AF",
		X"32",X"00",X"E7",X"32",X"1A",X"E7",X"11",X"83",X"E0",X"21",X"00",X"EA",X"06",X"03",X"1A",X"77",
		X"23",X"1B",X"10",X"FA",X"06",X"03",X"36",X"20",X"23",X"10",X"FB",X"0E",X"14",X"11",X"00",X"EA",
		X"06",X"03",X"1A",X"BE",X"38",X"1C",X"20",X"06",X"13",X"23",X"10",X"F6",X"18",X"14",X"78",X"C6",
		X"03",X"47",X"7E",X"F5",X"1A",X"77",X"F1",X"12",X"23",X"13",X"10",X"F6",X"0D",X"20",X"E1",X"13",
		X"13",X"13",X"79",X"FE",X"14",X"C8",X"04",X"05",X"28",X"03",X"13",X"10",X"FD",X"D5",X"F5",X"3E",
		X"24",X"CD",X"FE",X"0D",X"CD",X"20",X"56",X"21",X"8A",X"56",X"CD",X"1C",X"11",X"F1",X"11",X"11",
		X"DA",X"FE",X"0A",X"38",X"05",X"D6",X"0A",X"11",X"21",X"DA",X"2E",X"00",X"CB",X"3F",X"CB",X"1D",
		X"67",X"19",X"D1",X"06",X"0D",X"36",X"00",X"23",X"10",X"FB",X"01",X"FD",X"F7",X"09",X"06",X"03",
		X"3E",X"41",X"77",X"12",X"3E",X"20",X"32",X"26",X"E0",X"D5",X"11",X"60",X"D1",X"0E",X"00",X"CD",
		X"FF",X"10",X"D1",X"3E",X"38",X"32",X"81",X"E8",X"CD",X"0D",X"57",X"3A",X"04",X"E9",X"E6",X"03",
		X"20",X"69",X"3A",X"06",X"E9",X"E6",X"03",X"28",X"25",X"3A",X"83",X"E8",X"A7",X"20",X"23",X"3E",
		X"0B",X"32",X"83",X"E8",X"3A",X"06",X"E9",X"CB",X"47",X"7E",X"20",X"09",X"3D",X"FE",X"41",X"30",
		X"24",X"3E",X"5C",X"18",X"20",X"3C",X"FE",X"5D",X"38",X"1B",X"3E",X"41",X"18",X"17",X"AF",X"32",
		X"83",X"E8",X"3A",X"09",X"E9",X"E6",X"30",X"28",X"0E",X"7E",X"FE",X"5C",X"28",X"2D",X"13",X"23",
		X"05",X"28",X"1A",X"3E",X"41",X"77",X"12",X"3A",X"81",X"E8",X"A7",X"20",X"AB",X"3A",X"26",X"E0",
		X"D6",X"01",X"27",X"20",X"91",X"11",X"60",X"D1",X"0E",X"00",X"CD",X"FF",X"10",X"CD",X"2C",X"56",
		X"3E",X"1C",X"CD",X"0F",X"57",X"3E",X"00",X"CD",X"FE",X"0D",X"C9",X"3E",X"20",X"12",X"18",X"ED",
		X"CD",X"57",X"11",X"CD",X"03",X"57",X"21",X"75",X"56",X"CD",X"1C",X"11",X"21",X"06",X"EA",X"11",
		X"A1",X"D6",X"3E",X"20",X"F5",X"0E",X"D8",X"CD",X"F7",X"56",X"0E",X"15",X"13",X"7E",X"23",X"A7",
		X"D5",X"C4",X"08",X"11",X"D1",X"13",X"06",X"02",X"7E",X"23",X"CD",X"FF",X"10",X"10",X"F9",X"3E",
		X"30",X"CD",X"10",X"11",X"0E",X"00",X"13",X"06",X"03",X"7E",X"23",X"CD",X"10",X"11",X"10",X"F9",
		X"F1",X"D6",X"01",X"27",X"C8",X"E5",X"21",X"73",X"FF",X"19",X"EB",X"E1",X"FE",X"10",X"20",X"C4",
		X"11",X"91",X"D6",X"18",X"BF",X"FE",X"DB",X"FD",X"D8",X"D0",X"42",X"45",X"53",X"54",X"20",X"32",
		X"30",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"53",X"FF",X"FD",X"5A",X"D1",X"FE",X"14",X"54",
		X"49",X"4D",X"45",X"FF",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"54",X"49",X"4D",X"45",X"20",X"4F",X"56",X"45",X"52",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"0E",X"D8",X"DD",X"21",X"94",X"56",X"CD",X"C3",X"56",X"3E",X"70",
		X"C3",X"0F",X"57",X"2A",X"02",X"E9",X"11",X"04",X"00",X"19",X"29",X"29",X"29",X"29",X"29",X"7C",
		X"C6",X"1A",X"11",X"40",X"D3",X"6F",X"26",X"03",X"E5",X"06",X"0B",X"D5",X"7D",X"2C",X"E6",X"3F",
		X"B3",X"5F",X"DD",X"7E",X"00",X"DD",X"23",X"CD",X"10",X"11",X"D1",X"10",X"EE",X"21",X"40",X"00",
		X"19",X"EB",X"E1",X"25",X"20",X"E2",X"C9",X"FE",X"10",X"D2",X"FF",X"10",X"13",X"C3",X"08",X"11",
		X"CD",X"53",X"11",X"AF",X"32",X"00",X"E0",X"21",X"00",X"00",X"22",X"02",X"E9",X"3E",X"01",X"E5",
		X"21",X"82",X"E8",X"77",X"7E",X"A7",X"20",X"FC",X"E1",X"C9",X"C5",X"06",X"21",X"18",X"0E",X"CD",
		X"25",X"57",X"11",X"96",X"D3",X"C5",X"06",X"1A",X"18",X"03",X"C5",X"06",X"20",X"AF",X"CD",X"10",
		X"11",X"10",X"FB",X"C1",X"C9",X"5E",X"23",X"56",X"23",X"7E",X"23",X"3C",X"C8",X"3C",X"20",X"04",
		X"CB",X"E9",X"18",X"F5",X"3C",X"28",X"EE",X"D6",X"03",X"CB",X"B9",X"FE",X"08",X"38",X"02",X"CB",
		X"F9",X"CD",X"10",X"11",X"18",X"E3",X"2A",X"17",X"E8",X"7C",X"E5",X"CD",X"65",X"57",X"E1",X"24",
		X"7C",X"BD",X"20",X"F6",X"C9",X"FE",X"E0",X"D0",X"32",X"02",X"E8",X"C6",X"20",X"E6",X"3F",X"21",
		X"80",X"D1",X"B5",X"6F",X"3A",X"02",X"E8",X"CD",X"00",X"58",X"3A",X"80",X"E0",X"E6",X"01",X"20",
		X"05",X"CD",X"5F",X"58",X"18",X"03",X"CD",X"35",X"58",X"CD",X"03",X"59",X"20",X"05",X"CD",X"D3",
		X"58",X"18",X"03",X"CD",X"F1",X"58",X"CD",X"D4",X"57",X"CD",X"03",X"59",X"FE",X"03",X"C0",X"3A",
		X"02",X"E8",X"01",X"08",X"00",X"21",X"30",X"5A",X"ED",X"B9",X"C0",X"CB",X"01",X"CB",X"01",X"3A",
		X"80",X"E0",X"FE",X"10",X"21",X"31",X"5A",X"38",X"03",X"21",X"51",X"5A",X"09",X"5E",X"23",X"56",
		X"23",X"EB",X"0E",X"11",X"1A",X"13",X"77",X"CB",X"DC",X"71",X"1A",X"11",X"40",X"F8",X"19",X"77",
		X"CB",X"DC",X"71",X"C9",X"3A",X"80",X"E0",X"E6",X"01",X"21",X"7C",X"5A",X"20",X"03",X"21",X"88",
		X"5A",X"3A",X"02",X"E8",X"01",X"0C",X"00",X"ED",X"B9",X"C0",X"21",X"89",X"5A",X"09",X"09",X"3A",
		X"02",X"E8",X"EB",X"C6",X"20",X"E6",X"3F",X"21",X"80",X"D3",X"B5",X"6F",X"0E",X"8B",X"18",X"C4",
		X"11",X"E7",X"61",X"FE",X"DA",X"D2",X"18",X"59",X"D6",X"D5",X"38",X"0C",X"E5",X"21",X"DB",X"59",
		X"5F",X"16",X"00",X"19",X"7E",X"E1",X"18",X"04",X"E6",X"01",X"C6",X"52",X"0E",X"5C",X"CD",X"09",
		X"59",X"3A",X"02",X"E8",X"E6",X"07",X"E5",X"21",X"E1",X"59",X"4F",X"09",X"7E",X"E1",X"77",X"CB",
		X"DC",X"36",X"5E",X"19",X"C9",X"3A",X"02",X"E8",X"FE",X"DD",X"D0",X"FE",X"0D",X"38",X"0A",X"FE",
		X"CF",X"38",X"2A",X"11",X"83",X"5F",X"C3",X"C5",X"58",X"47",X"3A",X"15",X"E9",X"FE",X"01",X"78",
		X"11",X"48",X"5D",X"28",X"70",X"11",X"18",X"5E",X"30",X"6B",X"11",X"8E",X"5C",X"18",X"66",X"3A",
		X"02",X"E8",X"FE",X"DD",X"D0",X"FE",X"13",X"38",X"36",X"FE",X"D3",X"30",X"19",X"E6",X"1F",X"F5",
		X"E5",X"87",X"4F",X"21",X"E9",X"59",X"09",X"7E",X"23",X"4E",X"E1",X"77",X"CB",X"DC",X"71",X"19",
		X"F1",X"11",X"6A",X"5B",X"18",X"3F",X"47",X"11",X"CB",X"61",X"CD",X"03",X"59",X"28",X"0D",X"3A",
		X"15",X"E9",X"FE",X"01",X"11",X"76",X"61",X"30",X"03",X"11",X"F5",X"60",X"78",X"18",X"26",X"5F",
		X"CD",X"03",X"59",X"FE",X"04",X"7B",X"11",X"B3",X"60",X"28",X"1A",X"11",X"A9",X"5E",X"CD",X"18",
		X"59",X"CD",X"03",X"59",X"3A",X"02",X"E8",X"20",X"05",X"FE",X"03",X"30",X"0B",X"C9",X"FE",X"02",
		X"30",X"06",X"11",X"54",X"65",X"CD",X"18",X"59",X"36",X"05",X"CB",X"DC",X"36",X"01",X"11",X"40",
		X"F8",X"19",X"C9",X"0E",X"4F",X"3A",X"02",X"E8",X"FE",X"C0",X"30",X"10",X"FE",X"20",X"38",X"07",
		X"E6",X"1F",X"11",X"0C",X"65",X"18",X"31",X"11",X"02",X"64",X"18",X"2C",X"11",X"F8",X"62",X"18",
		X"27",X"3A",X"02",X"E8",X"11",X"A7",X"63",X"FE",X"DC",X"30",X"1D",X"E6",X"01",X"C6",X"24",X"0E",
		X"42",X"18",X"06",X"3A",X"80",X"E0",X"E6",X"07",X"C9",X"06",X"03",X"11",X"40",X"F8",X"77",X"CB",
		X"DC",X"71",X"19",X"C6",X"02",X"10",X"F7",X"C9",X"EB",X"C5",X"06",X"00",X"4F",X"09",X"09",X"C1",
		X"7E",X"23",X"66",X"6F",X"EB",X"06",X"01",X"1A",X"13",X"3C",X"28",X"13",X"3C",X"28",X"17",X"C6",
		X"FE",X"77",X"CB",X"DC",X"71",X"3E",X"40",X"85",X"6F",X"3E",X"F8",X"8C",X"67",X"18",X"E8",X"05",
		X"C8",X"D1",X"13",X"13",X"18",X"E1",X"1A",X"13",X"FE",X"FC",X"38",X"0C",X"28",X"02",X"D5",X"04",
		X"EB",X"7E",X"23",X"66",X"6F",X"EB",X"18",X"CF",X"4F",X"18",X"CC",X"FE",X"15",X"FD",X"D8",X"D2",
		X"53",X"45",X"4C",X"45",X"43",X"54",X"20",X"47",X"41",X"4D",X"45",X"20",X"46",X"4C",X"4F",X"4F",
		X"52",X"FD",X"9A",X"D3",X"48",X"4F",X"55",X"53",X"45",X"20",X"4E",X"55",X"4D",X"42",X"45",X"52",
		X"2D",X"FD",X"1A",X"D4",X"46",X"4C",X"4F",X"4F",X"52",X"20",X"4E",X"55",X"4D",X"42",X"45",X"52",
		X"2D",X"FD",X"98",X"D4",X"50",X"55",X"4E",X"43",X"48",X"2D",X"55",X"50",X"20",X"4B",X"49",X"43",
		X"4B",X"2D",X"44",X"4F",X"57",X"4E",X"FF",X"FE",X"15",X"FD",X"11",X"D0",X"31",X"50",X"2D",X"FD",
		X"26",X"D0",X"32",X"50",X"2D",X"FE",X"00",X"FD",X"1B",X"D0",X"54",X"4F",X"50",X"2D",X"FE",X"14",
		X"FD",X"AA",X"D0",X"54",X"49",X"4D",X"45",X"FE",X"94",X"FD",X"91",X"D0",X"98",X"99",X"9A",X"9B",
		X"9C",X"FE",X"95",X"FD",X"11",X"D1",X"9D",X"9E",X"9F",X"A0",X"FF",X"58",X"59",X"60",X"61",X"68",
		X"69",X"67",X"6E",X"5E",X"5E",X"5E",X"5E",X"5F",X"66",X"F1",X"08",X"06",X"01",X"06",X"01",X"06",
		X"01",X"06",X"01",X"14",X"41",X"15",X"41",X"EE",X"08",X"EF",X"08",X"06",X"01",X"06",X"01",X"18",
		X"41",X"19",X"41",X"06",X"01",X"06",X"01",X"EE",X"08",X"EF",X"08",X"06",X"01",X"06",X"01",X"14",
		X"41",X"15",X"41",X"06",X"01",X"06",X"01",X"EE",X"08",X"EF",X"08",X"18",X"41",X"19",X"41",X"06",
		X"01",X"06",X"01",X"06",X"01",X"06",X"01",X"F0",X"08",X"22",X"23",X"3C",X"3D",X"5A",X"5B",X"70",
		X"71",X"02",X"D3",X"7C",X"7E",X"03",X"D3",X"01",X"7F",X"1C",X"D4",X"7C",X"7E",X"1D",X"D4",X"01",
		X"7F",X"FA",X"D5",X"7C",X"7E",X"FB",X"D5",X"01",X"7F",X"10",X"D3",X"7C",X"7E",X"11",X"D3",X"01",
		X"7F",X"02",X"D3",X"7C",X"7E",X"03",X"D3",X"01",X"7F",X"1C",X"D4",X"7C",X"7E",X"1D",X"D4",X"01",
		X"7F",X"3A",X"D4",X"7C",X"7E",X"3B",X"D4",X"01",X"7F",X"10",X"D3",X"7C",X"7E",X"11",X"D3",X"01",
		X"7F",X"1F",X"20",X"3F",X"40",X"5F",X"60",X"7F",X"80",X"9F",X"A0",X"BF",X"C0",X"BF",X"C0",X"9F",
		X"A0",X"7F",X"80",X"5F",X"60",X"3F",X"40",X"1F",X"20",X"04",X"06",X"05",X"7D",X"7E",X"96",X"95",
		X"97",X"BC",X"BE",X"BD",X"BF",X"C0",X"C2",X"C1",X"C3",X"C4",X"C6",X"C5",X"C7",X"C8",X"CA",X"C9",
		X"CB",X"FD",X"FB",X"D4",X"FE",X"41",X"22",X"FD",X"3A",X"D5",X"80",X"FE",X"91",X"1F",X"94",X"FD",
		X"79",X"D5",X"26",X"FE",X"11",X"00",X"00",X"00",X"FD",X"B8",X"D5",X"FE",X"91",X"27",X"28",X"29",
		X"FE",X"11",X"00",X"00",X"FD",X"F8",X"D5",X"FE",X"91",X"30",X"2A",X"FE",X"11",X"03",X"FE",X"91",
		X"20",X"21",X"FD",X"38",X"D6",X"31",X"2C",X"2D",X"FE",X"11",X"03",X"FE",X"91",X"23",X"FD",X"79",
		X"D6",X"2E",X"2F",X"22",X"FE",X"11",X"03",X"FD",X"BA",X"D6",X"FE",X"91",X"2B",X"24",X"25",X"FF",
		X"FD",X"FC",X"D4",X"FE",X"41",X"22",X"FD",X"3B",X"D5",X"80",X"80",X"FD",X"79",X"D5",X"80",X"FD",
		X"B8",X"D5",X"80",X"80",X"80",X"FD",X"F8",X"D5",X"80",X"80",X"80",X"80",X"80",X"FD",X"38",X"D6",
		X"86",X"86",X"86",X"86",X"86",X"FD",X"77",X"D6",X"FE",X"91",X"36",X"37",X"32",X"32",X"32",X"33",
		X"FD",X"B6",X"D6",X"38",X"39",X"34",X"34",X"34",X"34",X"35",X"FF",X"FE",X"01",X"06",X"FE",X"FD",
		X"39",X"5B",X"80",X"80",X"86",X"FF",X"FE",X"01",X"06",X"FE",X"01",X"FE",X"FD",X"52",X"5B",X"FE",
		X"41",X"22",X"80",X"80",X"FF",X"FE",X"09",X"FE",X"FD",X"53",X"5B",X"FE",X"FC",X"53",X"5B",X"FE",
		X"01",X"06",X"F9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FE",X"01",X"03",X"03",X"03",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"FF",X"AA",X"5B",X"B3",X"5B",X"C4",X"5B",
		X"CE",X"5B",X"C4",X"5B",X"D5",X"5B",X"E8",X"5B",X"FB",X"5B",X"10",X"5C",X"25",X"5C",X"3A",X"5C",
		X"4F",X"5C",X"62",X"5C",X"CE",X"5B",X"C4",X"5B",X"CE",X"5B",X"C4",X"5B",X"CE",X"5B",X"C4",X"5B",
		X"D5",X"5B",X"E8",X"5B",X"FB",X"5B",X"10",X"5C",X"25",X"5C",X"3A",X"5C",X"4F",X"5C",X"62",X"5C",
		X"CE",X"5B",X"C4",X"5B",X"CE",X"5B",X"75",X"5C",X"83",X"5C",X"FE",X"FD",X"5B",X"5B",X"F2",X"F4",
		X"F6",X"04",X"FF",X"FE",X"FD",X"39",X"5B",X"FE",X"01",X"F7",X"F3",X"F5",X"FE",X"41",X"84",X"7C",
		X"FF",X"FE",X"01",X"06",X"FE",X"FD",X"2E",X"5B",X"7C",X"84",X"FF",X"FE",X"01",X"06",X"FE",X"FD",
		X"2E",X"5B",X"84",X"7C",X"FF",X"FE",X"41",X"16",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"1E",
		X"80",X"80",X"80",X"80",X"14",X"84",X"7C",X"FF",X"FE",X"41",X"17",X"88",X"1C",X"88",X"88",X"88",
		X"88",X"88",X"1F",X"88",X"88",X"88",X"88",X"15",X"7C",X"84",X"FF",X"FE",X"01",X"F9",X"FE",X"41",
		X"80",X"89",X"00",X"02",X"04",X"06",X"10",X"22",X"80",X"80",X"80",X"80",X"86",X"84",X"7C",X"FF",
		X"FE",X"01",X"F9",X"FE",X"41",X"80",X"89",X"01",X"03",X"05",X"07",X"11",X"22",X"80",X"80",X"80",
		X"80",X"86",X"7C",X"84",X"FF",X"FE",X"01",X"F9",X"FE",X"41",X"80",X"89",X"08",X"0A",X"0C",X"0E",
		X"12",X"22",X"80",X"80",X"80",X"80",X"86",X"84",X"7C",X"FF",X"FE",X"01",X"F9",X"FE",X"41",X"80",
		X"89",X"09",X"0B",X"0D",X"0F",X"13",X"22",X"80",X"80",X"80",X"80",X"86",X"7C",X"84",X"FF",X"FE",
		X"41",X"1A",X"23",X"1D",X"23",X"23",X"23",X"23",X"23",X"20",X"23",X"23",X"23",X"23",X"18",X"84",
		X"7C",X"FF",X"FE",X"41",X"1B",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"21",X"80",X"80",X"80",
		X"80",X"19",X"7C",X"84",X"FF",X"FE",X"FD",X"39",X"5B",X"FE",X"01",X"F8",X"FA",X"FC",X"FE",X"41",
		X"7C",X"84",X"FF",X"FE",X"FD",X"5B",X"5B",X"FB",X"FD",X"FE",X"41",X"7B",X"7C",X"FF",X"A8",X"5C",
		X"C2",X"5C",X"DD",X"5C",X"F3",X"5C",X"08",X"5D",X"20",X"5D",X"33",X"5D",X"3C",X"5D",X"0A",X"5E",
		X"CB",X"5B",X"C1",X"5B",X"CB",X"5B",X"C1",X"5B",X"FE",X"03",X"EF",X"FE",X"09",X"00",X"00",X"00",
		X"00",X"FE",X"92",X"3A",X"3C",X"3E",X"8E",X"FE",X"09",X"FE",X"FD",X"54",X"5B",X"CC",X"FE",X"01",
		X"ED",X"FF",X"FE",X"09",X"FE",X"FD",X"55",X"5B",X"FE",X"92",X"3B",X"3D",X"46",X"44",X"46",X"FE",
		X"09",X"00",X"00",X"00",X"00",X"FE",X"92",X"49",X"FE",X"93",X"4B",X"4D",X"FF",X"FE",X"41",X"15",
		X"17",X"88",X"88",X"88",X"88",X"FE",X"93",X"3F",X"40",X"42",X"47",X"45",X"48",X"4A",X"4C",X"4E",
		X"5C",X"5E",X"FF",X"FE",X"01",X"06",X"F9",X"FE",X"FD",X"55",X"5B",X"FE",X"93",X"41",X"43",X"52",
		X"54",X"56",X"58",X"5A",X"86",X"5D",X"5F",X"FF",X"FE",X"01",X"06",X"F9",X"FE",X"FD",X"54",X"5B",
		X"FE",X"93",X"51",X"53",X"55",X"57",X"59",X"5B",X"FE",X"01",X"06",X"FE",X"93",X"63",X"5F",X"FF",
		X"FE",X"FD",X"4F",X"5B",X"FE",X"93",X"4F",X"50",X"FE",X"13",X"00",X"00",X"00",X"06",X"FE",X"93",
		X"63",X"5F",X"FF",X"FE",X"FD",X"2B",X"5B",X"FE",X"93",X"63",X"5F",X"FF",X"FE",X"08",X"EE",X"FE",
		X"FD",X"2E",X"5B",X"FE",X"93",X"60",X"62",X"FF",X"62",X"5D",X"7D",X"5D",X"98",X"5D",X"B2",X"5D",
		X"CA",X"5D",X"D6",X"5D",X"E2",X"5D",X"F7",X"5D",X"0A",X"5E",X"CB",X"5B",X"C1",X"5B",X"CB",X"5B",
		X"C1",X"5B",X"FE",X"03",X"EF",X"FE",X"09",X"00",X"00",X"00",X"00",X"FE",X"92",X"87",X"8A",X"8C",
		X"8E",X"FE",X"09",X"FE",X"FD",X"55",X"5B",X"00",X"CC",X"FE",X"01",X"ED",X"FF",X"FE",X"09",X"FE",
		X"FD",X"55",X"5B",X"FE",X"92",X"88",X"8B",X"8D",X"8F",X"92",X"FE",X"09",X"00",X"00",X"00",X"00",
		X"CD",X"FE",X"01",X"ED",X"FE",X"92",X"74",X"FF",X"FE",X"41",X"15",X"17",X"88",X"88",X"88",X"88",
		X"88",X"FE",X"93",X"89",X"90",X"93",X"65",X"FE",X"41",X"88",X"88",X"88",X"15",X"FE",X"93",X"73",
		X"75",X"FF",X"FE",X"01",X"06",X"F9",X"FE",X"FD",X"54",X"5B",X"FE",X"93",X"91",X"64",X"FE",X"41",
		X"80",X"80",X"80",X"80",X"FE",X"93",X"6E",X"70",X"72",X"FF",X"FE",X"FD",X"36",X"5B",X"80",X"FE",
		X"93",X"6D",X"6F",X"71",X"5F",X"FF",X"FE",X"FD",X"36",X"5B",X"FE",X"93",X"68",X"6A",X"6C",X"63",
		X"5F",X"FF",X"FE",X"FD",X"4F",X"5B",X"FE",X"41",X"22",X"80",X"FE",X"93",X"66",X"69",X"6B",X"FE",
		X"13",X"02",X"FE",X"93",X"63",X"5F",X"FF",X"FE",X"08",X"EE",X"FE",X"FD",X"39",X"5B",X"FE",X"93",
		X"67",X"FE",X"41",X"80",X"86",X"FE",X"93",X"60",X"62",X"FF",X"FE",X"08",X"EF",X"FE",X"FD",X"2E",
		X"5B",X"FE",X"93",X"61",X"FE",X"41",X"84",X"FF",X"32",X"5E",X"4C",X"5E",X"74",X"5E",X"7D",X"5E",
		X"7D",X"5E",X"7D",X"5E",X"86",X"5E",X"8F",X"5E",X"9B",X"5E",X"CB",X"5B",X"C1",X"5B",X"CB",X"5B",
		X"C1",X"5B",X"FE",X"03",X"EF",X"FE",X"09",X"00",X"00",X"00",X"00",X"FE",X"92",X"76",X"3C",X"79",
		X"FE",X"09",X"FE",X"FD",X"54",X"5B",X"00",X"CC",X"FE",X"01",X"ED",X"FF",X"FE",X"09",X"FE",X"FD",
		X"55",X"5B",X"FE",X"92",X"77",X"78",X"FE",X"09",X"FE",X"FD",X"53",X"5B",X"CD",X"FE",X"92",X"7A",
		X"7C",X"FF",X"FE",X"41",X"15",X"17",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"1F",X"88",X"88",
		X"88",X"88",X"15",X"FF",X"FE",X"FD",X"62",X"5E",X"FE",X"92",X"7B",X"34",X"FF",X"FE",X"FD",X"2B",
		X"5B",X"FE",X"91",X"32",X"34",X"FF",X"FE",X"FD",X"2B",X"5B",X"FE",X"91",X"80",X"82",X"FF",X"FE",
		X"08",X"EE",X"FE",X"FD",X"2E",X"5B",X"FE",X"91",X"81",X"83",X"FF",X"FE",X"08",X"EF",X"FE",X"FD",
		X"2E",X"5B",X"FE",X"91",X"7F",X"FE",X"41",X"84",X"FF",X"CF",X"5E",X"E2",X"5E",X"F4",X"5E",X"0C",
		X"5F",X"21",X"5F",X"39",X"5F",X"53",X"5F",X"6D",X"5F",X"8B",X"5F",X"A7",X"5F",X"C3",X"5F",X"DF",
		X"5F",X"FD",X"5F",X"18",X"60",X"2B",X"60",X"47",X"60",X"65",X"60",X"83",X"60",X"9B",X"60",X"FE",
		X"03",X"EF",X"FE",X"09",X"00",X"00",X"00",X"C4",X"C6",X"C8",X"C8",X"C8",X"C9",X"CB",X"00",X"00",
		X"00",X"FF",X"FE",X"09",X"00",X"00",X"00",X"00",X"C5",X"C7",X"C7",X"C7",X"C7",X"CA",X"00",X"00",
		X"00",X"00",X"CD",X"FF",X"FE",X"09",X"C3",X"FE",X"41",X"17",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"1F",X"88",X"88",X"88",X"88",X"15",X"FE",X"07",X"80",X"82",X"FF",X"FE",X"06",X"A7",X"A8",
		X"FE",X"FD",X"53",X"5B",X"FE",X"41",X"22",X"80",X"80",X"80",X"80",X"86",X"FE",X"07",X"81",X"83",
		X"FF",X"FE",X"45",X"8A",X"FE",X"06",X"04",X"A9",X"AA",X"AB",X"AB",X"AB",X"AB",X"AB",X"BD",X"AB",
		X"AB",X"AB",X"AB",X"C0",X"FE",X"0A",X"D6",X"D4",X"FF",X"FE",X"06",X"A1",X"A2",X"FE",X"05",X"8C",
		X"FE",X"06",X"AC",X"AD",X"AE",X"AE",X"AE",X"AE",X"BE",X"AE",X"AE",X"AE",X"AE",X"C1",X"FE",X"4A",
		X"7D",X"7E",X"FF",X"FE",X"06",X"9E",X"A3",X"A6",X"FE",X"05",X"8F",X"FE",X"06",X"04",X"AF",X"B0",
		X"B1",X"B1",X"BF",X"B1",X"B1",X"B1",X"B1",X"C2",X"FE",X"4A",X"7F",X"83",X"FF",X"FE",X"08",X"EC",
		X"FE",X"06",X"A4",X"94",X"96",X"99",X"FE",X"05",X"8C",X"FE",X"06",X"B2",X"B3",X"00",X"FE",X"41",
		X"22",X"80",X"80",X"80",X"FE",X"04",X"84",X"86",X"88",X"8A",X"FF",X"FE",X"08",X"EF",X"FE",X"06",
		X"A5",X"95",X"97",X"9A",X"93",X"FE",X"05",X"8E",X"FE",X"06",X"04",X"B4",X"B5",X"00",X"00",X"00",
		X"FE",X"04",X"85",X"87",X"89",X"8B",X"FF",X"FE",X"01",X"06",X"F9",X"00",X"FE",X"06",X"98",X"9B",
		X"94",X"96",X"99",X"FE",X"05",X"8C",X"FE",X"06",X"B6",X"B7",X"AB",X"AB",X"AB",X"C0",X"FE",X"0A",
		X"D4",X"D6",X"FF",X"FE",X"01",X"06",X"F9",X"00",X"00",X"FE",X"06",X"9C",X"95",X"97",X"9A",X"93",
		X"FE",X"05",X"8E",X"FE",X"06",X"04",X"B8",X"B9",X"AE",X"C1",X"FE",X"0A",X"D5",X"D7",X"FF",X"FE",
		X"01",X"06",X"F9",X"00",X"00",X"00",X"00",X"FE",X"06",X"98",X"9B",X"94",X"9D",X"A0",X"FE",X"05",
		X"8C",X"FE",X"06",X"BA",X"BB",X"C2",X"FE",X"0A",X"D8",X"FE",X"41",X"7C",X"FF",X"FE",X"01",X"06",
		X"F9",X"FE",X"FD",X"55",X"5B",X"FE",X"06",X"9C",X"95",X"9E",X"9A",X"93",X"FE",X"05",X"8E",X"FE",
		X"06",X"04",X"BC",X"FE",X"0A",X"D3",X"03",X"FF",X"FE",X"FD",X"4F",X"5B",X"FE",X"06",X"9F",X"9B",
		X"94",X"96",X"99",X"FE",X"05",X"8C",X"FE",X"0A",X"D1",X"D2",X"FF",X"FE",X"01",X"06",X"F9",X"FE",
		X"0B",X"D9",X"DC",X"DC",X"DC",X"DC",X"DE",X"FE",X"41",X"80",X"22",X"FE",X"06",X"9C",X"95",X"97",
		X"9A",X"90",X"FE",X"05",X"8D",X"07",X"FF",X"FE",X"08",X"EE",X"FE",X"01",X"F9",X"FE",X"0B",X"DA",
		X"07",X"DB",X"DD",X"DF",X"E9",X"FE",X"41",X"80",X"22",X"80",X"80",X"FE",X"06",X"98",X"9B",X"91",
		X"FE",X"0A",X"CF",X"D0",X"FF",X"FE",X"08",X"EF",X"FE",X"01",X"F9",X"FE",X"0B",X"DA",X"E0",X"E2",
		X"E4",X"E6",X"E9",X"FE",X"41",X"80",X"22",X"80",X"80",X"80",X"FE",X"06",X"9C",X"92",X"FE",X"0A",
		X"CE",X"03",X"FF",X"FE",X"01",X"06",X"F9",X"FE",X"0B",X"DA",X"E1",X"E3",X"E5",X"E7",X"E9",X"FE",
		X"41",X"80",X"22",X"80",X"80",X"80",X"80",X"86",X"84",X"7C",X"FF",X"FE",X"01",X"06",X"F9",X"FE",
		X"0B",X"EB",X"E8",X"E8",X"E8",X"E8",X"EA",X"FE",X"41",X"80",X"22",X"80",X"80",X"80",X"80",X"86",
		X"7C",X"84",X"FF",X"15",X"61",X"09",X"61",X"02",X"61",X"F6",X"60",X"E5",X"60",X"D9",X"60",X"37",
		X"63",X"85",X"63",X"90",X"63",X"30",X"63",X"37",X"63",X"30",X"63",X"37",X"63",X"30",X"63",X"37",
		X"63",X"85",X"63",X"90",X"63",X"30",X"63",X"37",X"63",X"FE",X"FD",X"36",X"5B",X"80",X"80",X"FE",
		X"96",X"B4",X"B6",X"B5",X"FF",X"FE",X"FD",X"4F",X"5B",X"FE",X"41",X"22",X"80",X"FE",X"96",X"B7",
		X"AB",X"AD",X"AF",X"B1",X"B3",X"FF",X"FE",X"FD",X"36",X"5B",X"FE",X"96",X"AA",X"AC",X"AE",X"B0",
		X"B2",X"FF",X"FE",X"FD",X"62",X"5E",X"84",X"84",X"FF",X"FE",X"FD",X"45",X"5B",X"FE",X"92",X"49",
		X"FE",X"01",X"ED",X"04",X"FF",X"FE",X"03",X"EF",X"FE",X"FD",X"45",X"5B",X"CC",X"FE",X"01",X"ED",
		X"FF",X"3D",X"61",X"59",X"61",X"7B",X"61",X"9B",X"61",X"BB",X"61",X"D5",X"61",X"EB",X"61",X"03",
		X"62",X"1B",X"62",X"37",X"62",X"53",X"62",X"69",X"62",X"7D",X"62",X"91",X"62",X"FE",X"08",X"EE",
		X"FE",X"01",X"F9",X"FE",X"0B",X"D9",X"DC",X"DC",X"DC",X"DC",X"DE",X"04",X"FE",X"41",X"22",X"80",
		X"80",X"80",X"80",X"86",X"FE",X"4A",X"4E",X"81",X"FF",X"FE",X"08",X"EF",X"FE",X"01",X"F9",X"FE",
		X"0B",X"DA",X"FE",X"4B",X"87",X"8D",X"90",X"FE",X"0B",X"07",X"E9",X"04",X"FE",X"41",X"22",X"80",
		X"80",X"80",X"80",X"FE",X"46",X"4B",X"FE",X"4C",X"9B",X"A9",X"FF",X"FE",X"01",X"06",X"F9",X"FE",
		X"0B",X"DA",X"FE",X"4B",X"87",X"8E",X"91",X"FE",X"0B",X"07",X"E9",X"04",X"FE",X"41",X"22",X"80",
		X"80",X"FE",X"46",X"4C",X"FE",X"4C",X"83",X"9F",X"A7",X"87",X"FF",X"FE",X"01",X"06",X"F9",X"FE",
		X"0B",X"DA",X"FE",X"4B",X"8C",X"8F",X"92",X"FE",X"0B",X"07",X"E9",X"04",X"FE",X"41",X"22",X"80",
		X"FE",X"46",X"4B",X"FE",X"4C",X"9B",X"9C",X"49",X"A8",X"87",X"FF",X"FE",X"01",X"06",X"F9",X"FE",
		X"0B",X"EB",X"E8",X"E8",X"E8",X"E8",X"EA",X"04",X"FE",X"46",X"4D",X"FE",X"4C",X"83",X"9F",X"A0",
		X"A1",X"85",X"87",X"87",X"FF",X"FE",X"01",X"06",X"F9",X"FE",X"FD",X"54",X"5B",X"FE",X"46",X"4B",
		X"FE",X"4C",X"9B",X"A5",X"A6",X"9A",X"9A",X"42",X"43",X"44",X"FF",X"FE",X"01",X"06",X"F9",X"00",
		X"00",X"00",X"00",X"FE",X"46",X"4C",X"FE",X"4C",X"83",X"9F",X"A3",X"A4",X"3E",X"3E",X"3E",X"45",
		X"48",X"87",X"FF",X"FE",X"01",X"06",X"F9",X"00",X"00",X"00",X"FE",X"46",X"4B",X"FE",X"4C",X"9B",
		X"9C",X"A2",X"40",X"3D",X"3D",X"3D",X"3D",X"46",X"47",X"87",X"FF",X"FE",X"08",X"EE",X"FE",X"01",
		X"F9",X"00",X"FE",X"46",X"4C",X"FE",X"4C",X"83",X"9F",X"A0",X"A1",X"80",X"FE",X"41",X"22",X"80",
		X"80",X"80",X"80",X"86",X"84",X"84",X"FF",X"FE",X"08",X"EF",X"FE",X"01",X"F9",X"FE",X"46",X"4B",
		X"FE",X"4C",X"9B",X"9C",X"9D",X"9E",X"80",X"80",X"FE",X"41",X"22",X"80",X"80",X"80",X"80",X"86",
		X"84",X"84",X"FF",X"FE",X"46",X"4A",X"FE",X"4C",X"83",X"98",X"99",X"9A",X"9A",X"9A",X"9A",X"9A",
		X"41",X"9A",X"9A",X"9A",X"9A",X"42",X"43",X"44",X"FF",X"FE",X"4C",X"9B",X"95",X"96",X"97",X"3E",
		X"3E",X"3E",X"3E",X"3E",X"3F",X"3E",X"3E",X"3E",X"3E",X"45",X"48",X"87",X"FF",X"FE",X"4C",X"93",
		X"94",X"3D",X"3D",X"3D",X"3D",X"3D",X"3D",X"3D",X"40",X"3D",X"3D",X"3D",X"3D",X"46",X"47",X"87",
		X"FF",X"FE",X"4C",X"3C",X"FE",X"FD",X"2E",X"5B",X"84",X"84",X"FF",X"30",X"63",X"37",X"63",X"30",
		X"63",X"AF",X"62",X"B8",X"62",X"C4",X"62",X"D0",X"62",X"E5",X"62",X"F6",X"62",X"09",X"63",X"FE",
		X"FD",X"2B",X"5B",X"7C",X"FE",X"91",X"1C",X"FF",X"FE",X"08",X"EE",X"FE",X"FD",X"2E",X"5B",X"FE",
		X"91",X"18",X"1E",X"FF",X"FE",X"08",X"EF",X"FE",X"FD",X"2E",X"5B",X"FE",X"91",X"14",X"16",X"FF",
		X"FE",X"FD",X"4F",X"5B",X"FE",X"41",X"22",X"80",X"FE",X"91",X"1A",X"FE",X"41",X"80",X"80",X"86",
		X"FE",X"91",X"14",X"16",X"FF",X"FE",X"FD",X"4F",X"5B",X"FE",X"41",X"22",X"FE",X"91",X"19",X"1B",
		X"1D",X"10",X"12",X"14",X"16",X"FF",X"FE",X"FD",X"4F",X"5B",X"FE",X"91",X"08",X"0A",X"0C",X"FE",
		X"11",X"03",X"FE",X"91",X"11",X"13",X"15",X"17",X"FF",X"FE",X"FD",X"4F",X"5B",X"FE",X"91",X"09",
		X"0B",X"0D",X"0F",X"FE",X"11",X"03",X"03",X"FE",X"91",X"07",X"0E",X"FF",X"30",X"63",X"37",X"63",
		X"30",X"63",X"3E",X"63",X"47",X"63",X"53",X"63",X"5F",X"63",X"5F",X"63",X"5F",X"63",X"68",X"63",
		X"FE",X"FD",X"2B",X"5B",X"84",X"7C",X"FF",X"FE",X"FD",X"2B",X"5B",X"7C",X"84",X"FF",X"FE",X"FD",
		X"2B",X"5B",X"7C",X"FE",X"91",X"38",X"FF",X"FE",X"08",X"EE",X"FE",X"FD",X"2E",X"5B",X"FE",X"91",
		X"36",X"39",X"FF",X"FE",X"08",X"EF",X"FE",X"FD",X"2E",X"5B",X"FE",X"91",X"37",X"34",X"FF",X"FE",
		X"FD",X"2B",X"5B",X"FE",X"91",X"32",X"34",X"FF",X"FE",X"FD",X"2B",X"5B",X"FE",X"91",X"33",X"35",
		X"FF",X"30",X"63",X"37",X"63",X"30",X"63",X"37",X"63",X"85",X"63",X"90",X"63",X"30",X"63",X"37",
		X"63",X"30",X"63",X"37",X"63",X"FE",X"08",X"EE",X"FE",X"FD",X"2E",X"5B",X"FE",X"FC",X"34",X"63",
		X"FE",X"08",X"EF",X"FE",X"FD",X"2E",X"5B",X"FE",X"FC",X"3B",X"63",X"A7",X"63",X"B0",X"63",X"B9",
		X"63",X"C2",X"63",X"CF",X"63",X"E9",X"63",X"FE",X"5C",X"69",X"6B",X"6D",X"FE",X"5E",X"8B",X"FF",
		X"FE",X"5C",X"70",X"72",X"FE",X"5E",X"78",X"84",X"FF",X"FE",X"5C",X"71",X"73",X"FE",X"5E",X"79",
		X"84",X"FF",X"FE",X"5C",X"74",X"76",X"FE",X"5D",X"4F",X"87",X"87",X"FE",X"FC",X"D8",X"63",X"FE",
		X"5C",X"75",X"77",X"FE",X"5D",X"50",X"FE",X"5F",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",
		X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"FF",X"FE",X"5C",X"6F",X"7A",X"FE",X"5D",X"51",
		X"FE",X"5F",X"87",X"87",X"87",X"87",X"87",X"37",X"38",X"39",X"39",X"3A",X"3B",X"87",X"87",X"87",
		X"87",X"FF",X"42",X"64",X"4E",X"64",X"5D",X"64",X"BC",X"64",X"C0",X"64",X"64",X"64",X"68",X"64",
		X"D8",X"64",X"E8",X"64",X"74",X"64",X"6C",X"64",X"70",X"64",X"D8",X"64",X"E8",X"64",X"D8",X"64",
		X"E8",X"64",X"D8",X"64",X"DC",X"64",X"E0",X"64",X"E4",X"64",X"E8",X"64",X"D8",X"64",X"DC",X"64",
		X"E0",X"64",X"E4",X"64",X"E8",X"64",X"D8",X"64",X"E8",X"64",X"C8",X"64",X"CC",X"64",X"D0",X"64",
		X"D4",X"64",X"FE",X"4D",X"FA",X"FC",X"FE",X"70",X"AF",X"B1",X"B3",X"B5",X"B7",X"FF",X"FE",X"4D",
		X"FD",X"FE",X"8D",X"85",X"FE",X"8E",X"84",X"FE",X"50",X"B2",X"B4",X"B6",X"FF",X"FE",X"8E",X"00",
		X"01",X"02",X"03",X"FF",X"F4",X"F6",X"D8",X"FF",X"F5",X"F7",X"80",X"FF",X"F0",X"F2",X"D8",X"FF",
		X"F1",X"F3",X"80",X"FF",X"F8",X"D5",X"D7",X"FF",X"D8",X"64",X"E8",X"64",X"B8",X"64",X"BC",X"64",
		X"C0",X"64",X"C4",X"64",X"D8",X"64",X"E8",X"64",X"C8",X"64",X"CC",X"64",X"D0",X"64",X"D4",X"64",
		X"D8",X"64",X"E8",X"64",X"D8",X"64",X"E8",X"64",X"D8",X"64",X"E8",X"64",X"D8",X"64",X"DC",X"64",
		X"E0",X"64",X"E4",X"64",X"E8",X"64",X"D8",X"64",X"DC",X"64",X"E0",X"64",X"E4",X"64",X"E8",X"64",
		X"EC",X"64",X"F2",X"64",X"F9",X"64",X"02",X"65",X"C6",X"C2",X"80",X"FF",X"C7",X"C2",X"80",X"FF",
		X"CE",X"D5",X"D7",X"FF",X"CF",X"D6",X"D8",X"FF",X"C8",X"CA",X"80",X"FF",X"C9",X"CB",X"CD",X"FF",
		X"D0",X"D2",X"D4",X"FF",X"D1",X"D3",X"80",X"FF",X"AA",X"C2",X"80",X"FF",X"B8",X"C2",X"C4",X"FF",
		X"C1",X"C3",X"C5",X"FF",X"AA",X"C0",X"CC",X"FF",X"B8",X"C2",X"80",X"FF",X"BA",X"BC",X"FE",X"50",
		X"BE",X"FF",X"FE",X"50",X"B9",X"BB",X"BD",X"BF",X"FF",X"FE",X"50",X"AC",X"AE",X"B0",X"B2",X"B4",
		X"B6",X"FF",X"FE",X"50",X"AB",X"AD",X"AF",X"B1",X"B3",X"B5",X"B7",X"FF",X"4C",X"65",X"D8",X"64",
		X"E8",X"64",X"50",X"65",X"E0",X"64",X"E4",X"64",X"E8",X"64",X"D8",X"64",X"DC",X"64",X"E0",X"64",
		X"E4",X"64",X"E8",X"64",X"D8",X"64",X"E8",X"64",X"D8",X"64",X"E8",X"64",X"D8",X"64",X"DC",X"64",
		X"E0",X"64",X"E4",X"64",X"E8",X"64",X"D8",X"64",X"DC",X"64",X"E0",X"64",X"E4",X"64",X"E8",X"64",
		X"D8",X"64",X"E8",X"64",X"C8",X"64",X"CC",X"64",X"D0",X"64",X"D4",X"64",X"E3",X"E5",X"80",X"FF",
		X"E4",X"E6",X"C4",X"FF",X"46",X"5E",X"58",X"65",X"FE",X"01",X"ED",X"FE",X"41",X"7C",X"FF",X"67",
		X"65",X"6D",X"65",X"76",X"65",X"81",X"65",X"FE",X"42",X"24",X"26",X"30",X"FF",X"FE",X"5D",X"87",
		X"FE",X"42",X"2A",X"2C",X"2E",X"FF",X"FE",X"5F",X"87",X"87",X"35",X"FE",X"42",X"2B",X"2D",X"2F",
		X"FF",X"FE",X"5F",X"87",X"87",X"36",X"FE",X"42",X"31",X"32",X"33",X"34",X"FF",X"05",X"01",X"07",
		X"0B",X"FE",X"06",X"05",X"02",X"09",X"0B",X"FD",X"08",X"05",X"01",X"0C",X"0B",X"FE",X"0B",X"05",
		X"02",X"0E",X"0B",X"FD",X"0D",X"B7",X"65",X"B7",X"65",X"D5",X"65",X"E0",X"65",X"EB",X"65",X"F1",
		X"65",X"00",X"00",X"F7",X"65",X"FB",X"65",X"02",X"00",X"00",X"02",X"00",X"03",X"05",X"19",X"01",
		X"05",X"B3",X"00",X"05",X"00",X"00",X"05",X"4D",X"FF",X"05",X"E7",X"FE",X"02",X"00",X"FD",X"02",
		X"00",X"00",X"FF",X"00",X"00",X"04",X"10",X"06",X"12",X"10",X"93",X"06",X"14",X"04",X"10",X"00",
		X"04",X"11",X"06",X"12",X"10",X"93",X"06",X"14",X"04",X"10",X"00",X"05",X"55",X"01",X"88",X"00",
		X"00",X"05",X"56",X"01",X"88",X"00",X"00",X"05",X"B8",X"00",X"00",X"05",X"B9",X"00",X"00",X"9B",
		X"66",X"BF",X"66",X"D9",X"66",X"FD",X"66",X"1D",X"67",X"45",X"67",X"93",X"68",X"BD",X"68",X"47",
		X"68",X"6B",X"68",X"1F",X"68",X"77",X"69",X"A1",X"69",X"2B",X"69",X"4F",X"69",X"03",X"69",X"9F",
		X"67",X"C9",X"69",X"B9",X"67",X"D9",X"67",X"FF",X"67",X"6B",X"68",X"6B",X"68",X"6B",X"68",X"E5",
		X"68",X"E5",X"68",X"00",X"00",X"00",X"00",X"63",X"67",X"74",X"67",X"81",X"67",X"92",X"67",X"F3",
		X"69",X"07",X"6A",X"27",X"6A",X"3C",X"6A",X"51",X"6A",X"66",X"6A",X"66",X"74",X"AC",X"66",X"CC",
		X"66",X"EA",X"66",X"0A",X"67",X"32",X"67",X"56",X"67",X"A4",X"68",X"D2",X"68",X"58",X"68",X"80",
		X"68",X"34",X"68",X"88",X"69",X"B6",X"69",X"3C",X"69",X"64",X"69",X"18",X"69",X"AC",X"67",X"DA",
		X"69",X"C6",X"67",X"E6",X"67",X"0C",X"68",X"80",X"68",X"80",X"68",X"80",X"68",X"F6",X"68",X"F6",
		X"68",X"00",X"00",X"00",X"00",X"BE",X"66",X"BE",X"66",X"BE",X"66",X"BE",X"66",X"00",X"6A",X"14",
		X"6A",X"BE",X"66",X"BE",X"66",X"BE",X"66",X"BE",X"66",X"BE",X"66",X"27",X"10",X"02",X"80",X"2D",
		X"10",X"02",X"82",X"23",X"2C",X"00",X"84",X"28",X"30",X"01",X"02",X"FF",X"3D",X"4A",X"A0",X"FF",
		X"20",X"FF",X"0F",X"3F",X"40",X"00",X"40",X"FF",X"0F",X"38",X"A0",X"00",X"00",X"00",X"FF",X"29",
		X"10",X"02",X"86",X"28",X"30",X"01",X"03",X"28",X"40",X"00",X"04",X"FF",X"42",X"4B",X"C0",X"FF",
		X"40",X"FF",X"0F",X"42",X"60",X"00",X"60",X"FF",X"FF",X"26",X"10",X"02",X"8E",X"2D",X"10",X"02",
		X"90",X"22",X"2C",X"00",X"92",X"28",X"2F",X"01",X"0B",X"FF",X"30",X"49",X"C0",X"FF",X"40",X"FF",
		X"0F",X"3E",X"A0",X"00",X"C0",X"FF",X"0F",X"28",X"00",X"00",X"00",X"FF",X"FF",X"27",X"3F",X"00",
		X"04",X"28",X"10",X"02",X"94",X"28",X"30",X"01",X"0D",X"FF",X"40",X"4B",X"C0",X"FF",X"20",X"FF",
		X"0F",X"41",X"40",X"00",X"60",X"FF",X"0F",X"1C",X"A0",X"00",X"00",X"00",X"FF",X"2A",X"3B",X"00",
		X"2A",X"22",X"10",X"02",X"88",X"2A",X"10",X"02",X"8A",X"22",X"30",X"01",X"05",X"29",X"2D",X"01",
		X"06",X"FF",X"0F",X"45",X"40",X"00",X"E0",X"FF",X"0F",X"3A",X"E0",X"00",X"A0",X"FF",X"0F",X"26",
		X"00",X"00",X"40",X"FF",X"FF",X"25",X"10",X"02",X"8C",X"2E",X"10",X"02",X"08",X"28",X"20",X"01",
		X"09",X"27",X"2D",X"00",X"0A",X"FF",X"0F",X"35",X"A0",X"FF",X"20",X"FF",X"0F",X"2C",X"80",X"00",
		X"A0",X"FF",X"FF",X"1F",X"1D",X"02",X"9A",X"24",X"12",X"02",X"9C",X"25",X"32",X"01",X"17",X"25",
		X"42",X"00",X"16",X"FF",X"2A",X"10",X"02",X"9E",X"2A",X"30",X"01",X"19",X"28",X"40",X"00",X"1C",
		X"FF",X"20",X"1D",X"02",X"A0",X"25",X"12",X"02",X"A2",X"25",X"32",X"01",X"1B",X"24",X"42",X"00",
		X"1A",X"FF",X"2A",X"10",X"02",X"A4",X"2A",X"30",X"01",X"1D",X"28",X"40",X"00",X"1C",X"FF",X"2A",
		X"3C",X"00",X"21",X"28",X"10",X"02",X"A6",X"28",X"2E",X"01",X"1F",X"FF",X"0F",X"46",X"00",X"00",
		X"80",X"FF",X"0F",X"37",X"A0",X"00",X"00",X"00",X"FF",X"29",X"49",X"00",X"21",X"28",X"10",X"02",
		X"A8",X"28",X"2B",X"01",X"AA",X"FF",X"46",X"50",X"E0",X"FF",X"60",X"FF",X"39",X"46",X"60",X"00",
		X"A0",X"FF",X"14",X"39",X"60",X"00",X"C0",X"FF",X"FF",X"28",X"17",X"02",X"AC",X"29",X"31",X"01",
		X"22",X"28",X"41",X"00",X"21",X"FF",X"36",X"4A",X"C0",X"FF",X"40",X"FF",X"2B",X"3F",X"C0",X"00",
		X"E0",X"FF",X"1E",X"2C",X"20",X"00",X"40",X"FF",X"1A",X"1E",X"40",X"00",X"00",X"00",X"FF",X"28",
		X"49",X"00",X"21",X"28",X"10",X"02",X"A8",X"29",X"2B",X"01",X"AE",X"FF",X"48",X"53",X"C0",X"FF",
		X"40",X"FF",X"2F",X"48",X"60",X"00",X"A0",X"FF",X"14",X"2F",X"40",X"00",X"C0",X"FF",X"FF",X"25",
		X"10",X"02",X"B0",X"2A",X"10",X"02",X"B2",X"1C",X"38",X"01",X"24",X"2A",X"30",X"01",X"25",X"2C",
		X"40",X"00",X"26",X"FF",X"0F",X"4B",X"40",X"01",X"C0",X"FF",X"0F",X"29",X"80",X"01",X"00",X"FF",
		X"0F",X"2F",X"80",X"01",X"A0",X"FF",X"FF",X"25",X"10",X"02",X"B0",X"2A",X"10",X"02",X"B2",X"29",
		X"30",X"01",X"28",X"29",X"40",X"00",X"27",X"FF",X"0F",X"4B",X"40",X"00",X"C0",X"FF",X"0F",X"2A",
		X"80",X"00",X"00",X"FF",X"32",X"40",X"A0",X"00",X"20",X"00",X"FF",X"25",X"10",X"02",X"B0",X"2A",
		X"10",X"02",X"B2",X"1C",X"38",X"01",X"29",X"28",X"30",X"01",X"2B",X"28",X"40",X"00",X"2A",X"FF",
		X"0F",X"4A",X"40",X"00",X"A0",X"FF",X"0F",X"29",X"80",X"00",X"00",X"FF",X"29",X"3F",X"80",X"00",
		X"C0",X"FF",X"FF",X"1D",X"24",X"02",X"B4",X"2D",X"10",X"02",X"B8",X"2D",X"30",X"01",X"B6",X"2D",
		X"40",X"00",X"2C",X"FF",X"27",X"4B",X"80",X"00",X"00",X"00",X"0F",X"27",X"C0",X"00",X"40",X"00",
		X"30",X"3F",X"E0",X"00",X"A0",X"00",X"2F",X"37",X"00",X"00",X"40",X"FF",X"FF",X"0E",X"38",X"02",
		X"2D",X"1E",X"30",X"02",X"32",X"28",X"10",X"02",X"C4",X"2E",X"30",X"01",X"34",X"2E",X"40",X"00",
		X"33",X"FF",X"37",X"4A",X"A0",X"00",X"20",X"00",X"35",X"3F",X"20",X"01",X"20",X"FF",X"13",X"38",
		X"40",X"00",X"A0",X"FF",X"FF",X"27",X"46",X"00",X"27",X"28",X"10",X"02",X"C6",X"28",X"28",X"01",
		X"CA",X"18",X"37",X"02",X"C8",X"FF",X"13",X"51",X"00",X"00",X"80",X"FF",X"31",X"47",X"80",X"00",
		X"00",X"00",X"FF",X"25",X"10",X"02",X"96",X"35",X"10",X"02",X"98",X"1E",X"28",X"01",X"11",X"2E",
		X"23",X"01",X"0F",X"2D",X"33",X"00",X"0E",X"FF",X"0F",X"3A",X"60",X"00",X"E0",X"FF",X"0F",X"31",
		X"C0",X"00",X"00",X"00",X"0F",X"22",X"40",X"00",X"20",X"FF",X"FF",X"25",X"10",X"02",X"96",X"35",
		X"10",X"02",X"98",X"2A",X"23",X"01",X"13",X"2A",X"33",X"00",X"12",X"FF",X"0F",X"3A",X"60",X"00",
		X"E0",X"FF",X"0F",X"32",X"C0",X"00",X"20",X"00",X"0F",X"22",X"20",X"00",X"20",X"FF",X"FF",X"25",
		X"10",X"02",X"96",X"35",X"10",X"02",X"98",X"1F",X"28",X"01",X"10",X"28",X"23",X"01",X"15",X"28",
		X"33",X"00",X"14",X"FF",X"0F",X"3A",X"40",X"00",X"C0",X"FF",X"0F",X"30",X"C0",X"00",X"E0",X"FF",
		X"0F",X"22",X"E0",X"FF",X"00",X"FF",X"FF",X"20",X"10",X"02",X"CC",X"28",X"20",X"00",X"CE",X"30",
		X"10",X"02",X"37",X"30",X"20",X"01",X"36",X"FF",X"1D",X"38",X"80",X"00",X"00",X"00",X"0F",X"2C",
		X"40",X"01",X"A0",X"00",X"1F",X"2B",X"00",X"00",X"40",X"FF",X"0F",X"1F",X"40",X"FF",X"C0",X"FE",
		X"FF",X"0F",X"10",X"02",X"3B",X"1F",X"10",X"02",X"D4",X"26",X"1A",X"00",X"D8",X"30",X"10",X"02",
		X"D6",X"2D",X"23",X"01",X"3C",X"FF",X"1A",X"38",X"20",X"00",X"A0",X"FF",X"19",X"2D",X"00",X"01",
		X"E0",X"FE",X"0F",X"1F",X"C0",X"01",X"E0",X"00",X"FF",X"18",X"39",X"00",X"21",X"12",X"1B",X"02",
		X"2E",X"22",X"10",X"02",X"C2",X"1B",X"2B",X"01",X"31",X"FF",X"39",X"42",X"C0",X"FD",X"40",X"FD",
		X"2A",X"39",X"A0",X"FE",X"C0",X"FD",X"1F",X"2F",X"40",X"FF",X"40",X"FE",X"0F",X"20",X"A0",X"FF",
		X"00",X"FF",X"FF",X"29",X"40",X"00",X"3E",X"29",X"30",X"01",X"3F",X"29",X"10",X"02",X"42",X"FF",
		X"0F",X"4B",X"20",X"00",X"A0",X"FF",X"FF",X"25",X"3F",X"00",X"07",X"2B",X"2F",X"01",X"35",X"2C",
		X"10",X"02",X"44",X"FF",X"40",X"48",X"A0",X"FF",X"20",X"FF",X"34",X"3F",X"60",X"00",X"C0",X"FF",
		X"0F",X"3A",X"C0",X"00",X"20",X"00",X"FF",X"2A",X"40",X"00",X"3D",X"20",X"30",X"41",X"2B",X"30",
		X"30",X"41",X"3E",X"20",X"10",X"02",X"46",X"30",X"10",X"02",X"48",X"FF",X"26",X"33",X"41",X"3F",
		X"36",X"31",X"80",X"EA",X"1C",X"14",X"02",X"4A",X"2C",X"13",X"02",X"4C",X"3C",X"19",X"00",X"4E",
		X"FF",X"2E",X"40",X"80",X"EB",X"1E",X"30",X"81",X"EC",X"2E",X"30",X"81",X"ED",X"1E",X"10",X"02",
		X"50",X"2E",X"10",X"02",X"52",X"FF",X"27",X"36",X"81",X"EE",X"37",X"2C",X"80",X"EF",X"17",X"10",
		X"02",X"54",X"27",X"16",X"01",X"56",X"37",X"10",X"01",X"58",X"FF",X"97",X"6A",X"A4",X"6A",X"B1",
		X"6A",X"A4",X"6A",X"D8",X"6A",X"CB",X"6A",X"BE",X"6A",X"E5",X"6A",X"F2",X"6A",X"FF",X"6A",X"22",
		X"6B",X"19",X"6B",X"0C",X"6B",X"19",X"6B",X"2D",X"40",X"45",X"00",X"27",X"10",X"44",X"80",X"2D",
		X"10",X"44",X"40",X"FF",X"2D",X"40",X"45",X"00",X"29",X"30",X"44",X"01",X"29",X"10",X"44",X"42",
		X"FF",X"2D",X"40",X"45",X"00",X"28",X"10",X"44",X"84",X"31",X"10",X"44",X"44",X"FF",X"27",X"3C",
		X"45",X"02",X"21",X"20",X"44",X"46",X"2C",X"10",X"44",X"48",X"FF",X"24",X"28",X"44",X"4A",X"28",
		X"2B",X"45",X"4C",X"28",X"10",X"44",X"4E",X"FF",X"2C",X"0C",X"45",X"98",X"25",X"20",X"44",X"56",
		X"25",X"10",X"44",X"04",X"FF",X"19",X"0D",X"45",X"88",X"1F",X"1A",X"44",X"50",X"2F",X"0D",X"44",
		X"8C",X"FF",X"1C",X"0D",X"45",X"90",X"2C",X"17",X"44",X"52",X"35",X"0D",X"44",X"54",X"FF",X"28",
		X"3F",X"45",X"00",X"26",X"10",X"44",X"94",X"36",X"30",X"44",X"03",X"FF",X"29",X"40",X"85",X"00",
		X"26",X"10",X"44",X"F6",X"36",X"10",X"84",X"DA",X"FF",X"2A",X"40",X"85",X"00",X"2A",X"10",X"44",
		X"FC",X"FF",X"2A",X"40",X"85",X"00",X"26",X"10",X"44",X"FA",X"36",X"10",X"C4",X"F2",X"FF",X"51",
		X"6B",X"5E",X"6B",X"6B",X"6B",X"5E",X"6B",X"85",X"6B",X"78",X"6B",X"00",X"00",X"92",X"6B",X"9B",
		X"6B",X"A4",X"6B",X"B1",X"6B",X"B1",X"6B",X"BA",X"6B",X"C3",X"6B",X"CC",X"6B",X"D5",X"6B",X"DE",
		X"6B",X"28",X"30",X"91",X"10",X"28",X"20",X"91",X"11",X"28",X"10",X"92",X"82",X"FF",X"28",X"30",
		X"91",X"10",X"28",X"20",X"91",X"12",X"28",X"10",X"92",X"84",X"FF",X"27",X"30",X"91",X"10",X"28",
		X"20",X"91",X"13",X"28",X"10",X"92",X"86",X"FF",X"28",X"20",X"91",X"88",X"28",X"10",X"92",X"8A",
		X"2B",X"2E",X"47",X"0C",X"FF",X"28",X"20",X"91",X"92",X"28",X"10",X"92",X"94",X"2C",X"0C",X"47",
		X"0C",X"FF",X"22",X"18",X"91",X"96",X"2D",X"10",X"92",X"98",X"FF",X"1E",X"12",X"91",X"8C",X"2E",
		X"12",X"92",X"8E",X"FF",X"27",X"2D",X"91",X"10",X"29",X"10",X"92",X"90",X"2C",X"20",X"91",X"14",
		X"FF",X"2A",X"18",X"D1",X"F4",X"2A",X"10",X"D2",X"F6",X"FF",X"2C",X"1E",X"D1",X"F8",X"2A",X"0A",
		X"D2",X"FA",X"FF",X"29",X"0D",X"D1",X"FC",X"26",X"12",X"92",X"FB",X"FF",X"27",X"0D",X"D1",X"FE",
		X"20",X"16",X"92",X"FC",X"FF",X"27",X"0D",X"D1",X"FC",X"24",X"18",X"92",X"FB",X"FF",X"28",X"0A",
		X"D1",X"FE",X"21",X"11",X"92",X"FC",X"FF",X"01",X"6C",X"0E",X"6C",X"17",X"6C",X"0E",X"6C",X"2D",
		X"6C",X"3A",X"6C",X"24",X"6C",X"47",X"6C",X"54",X"6C",X"77",X"6C",X"84",X"6C",X"61",X"6C",X"6A",
		X"6C",X"25",X"30",X"06",X"BE",X"25",X"10",X"06",X"C0",X"2A",X"10",X"46",X"58",X"FF",X"25",X"30",
		X"06",X"BA",X"25",X"10",X"06",X"BC",X"FF",X"25",X"30",X"06",X"D0",X"25",X"10",X"06",X"D2",X"2B",
		X"10",X"46",X"5A",X"FF",X"27",X"10",X"46",X"A0",X"2D",X"3E",X"47",X"05",X"FF",X"20",X"29",X"46",
		X"06",X"26",X"0C",X"46",X"AC",X"30",X"0C",X"47",X"07",X"FF",X"20",X"10",X"46",X"D0",X"2A",X"2D",
		X"47",X"0C",X"30",X"10",X"46",X"D4",X"FF",X"17",X"25",X"46",X"5C",X"27",X"0E",X"46",X"B0",X"37",
		X"10",X"46",X"5E",X"FF",X"17",X"0A",X"46",X"B4",X"27",X"0A",X"46",X"B8",X"37",X"0A",X"46",X"60",
		X"FF",X"27",X"10",X"46",X"BC",X"27",X"48",X"47",X"08",X"FF",X"26",X"10",X"46",X"C0",X"36",X"37",
		X"46",X"09",X"36",X"10",X"46",X"0A",X"FF",X"17",X"30",X"46",X"0B",X"17",X"10",X"46",X"62",X"27",
		X"10",X"46",X"C4",X"FF",X"1F",X"10",X"46",X"C8",X"2F",X"10",X"46",X"CC",X"FF",X"C5",X"6C",X"D6",
		X"6C",X"E7",X"6C",X"D6",X"6C",X"26",X"6D",X"50",X"6D",X"93",X"6D",X"50",X"6D",X"26",X"6D",X"0D",
		X"6D",X"3B",X"6D",X"7E",X"6D",X"3B",X"6D",X"0D",X"6D",X"F8",X"6C",X"3B",X"6D",X"65",X"6D",X"3B",
		X"6D",X"F8",X"6C",X"DA",X"6D",X"C5",X"6D",X"AC",X"6D",X"0C",X"6E",X"F3",X"6D",X"25",X"6E",X"36",
		X"6E",X"43",X"6E",X"58",X"6E",X"20",X"10",X"48",X"64",X"30",X"10",X"49",X"66",X"24",X"30",X"49",
		X"68",X"34",X"30",X"49",X"0D",X"FF",X"26",X"10",X"48",X"0E",X"26",X"20",X"49",X"6A",X"26",X"40",
		X"49",X"0F",X"36",X"28",X"49",X"10",X"FF",X"20",X"10",X"49",X"6C",X"27",X"30",X"49",X"6E",X"30",
		X"10",X"48",X"70",X"38",X"29",X"49",X"10",X"FF",X"21",X"10",X"48",X"72",X"31",X"10",X"48",X"74",
		X"18",X"2D",X"49",X"76",X"28",X"20",X"49",X"D8",X"18",X"4C",X"48",X"11",X"FF",X"25",X"40",X"49",
		X"0F",X"08",X"30",X"49",X"78",X"18",X"36",X"49",X"12",X"21",X"10",X"48",X"72",X"30",X"10",X"48",
		X"74",X"28",X"2B",X"49",X"7A",X"FF",X"20",X"10",X"48",X"25",X"30",X"10",X"49",X"26",X"14",X"28",
		X"09",X"FC",X"1A",X"20",X"49",X"27",X"2A",X"20",X"49",X"7C",X"FF",X"29",X"3C",X"49",X"0F",X"1D",
		X"10",X"48",X"7E",X"2D",X"10",X"08",X"DA",X"1D",X"40",X"49",X"13",X"25",X"2A",X"09",X"DC",X"FF",
		X"2B",X"2B",X"49",X"0F",X"1C",X"10",X"48",X"14",X"2C",X"10",X"49",X"15",X"1C",X"2C",X"49",X"16",
		X"28",X"20",X"09",X"DE",X"FF",X"27",X"40",X"49",X"0F",X"23",X"10",X"08",X"E0",X"33",X"10",X"09",
		X"E2",X"25",X"30",X"09",X"E4",X"35",X"38",X"49",X"17",X"45",X"38",X"49",X"18",X"FF",X"1C",X"08",
		X"08",X"E6",X"1C",X"28",X"49",X"19",X"2C",X"10",X"49",X"DC",X"3C",X"30",X"49",X"1A",X"4B",X"30",
		X"49",X"1B",X"FF",X"2A",X"2B",X"49",X"0F",X"1F",X"10",X"48",X"1C",X"2F",X"10",X"09",X"E8",X"26",
		X"20",X"49",X"1D",X"3E",X"20",X"49",X"1E",X"4E",X"20",X"49",X"1F",X"FF",X"18",X"38",X"09",X"EA",
		X"18",X"30",X"48",X"20",X"25",X"10",X"08",X"EC",X"28",X"28",X"09",X"EE",X"28",X"48",X"49",X"21",
		X"2B",X"3C",X"47",X"0C",X"FF",X"0F",X"48",X"09",X"F0",X"17",X"38",X"49",X"22",X"27",X"10",X"08",
		X"F2",X"27",X"2E",X"09",X"F4",X"2D",X"2B",X"47",X"07",X"FF",X"12",X"3F",X"09",X"F6",X"16",X"38",
		X"49",X"23",X"26",X"30",X"09",X"F8",X"28",X"28",X"49",X"24",X"25",X"10",X"08",X"FA",X"2C",X"0E",
		X"47",X"0C",X"FF",X"20",X"10",X"48",X"25",X"30",X"10",X"49",X"26",X"14",X"28",X"09",X"FC",X"1A",
		X"20",X"49",X"27",X"28",X"20",X"09",X"FE",X"2D",X"2B",X"47",X"0C",X"FF",X"20",X"10",X"48",X"25",
		X"30",X"10",X"49",X"26",X"14",X"28",X"09",X"FC",X"1A",X"20",X"49",X"27",X"2A",X"20",X"09",X"60",
		X"33",X"0D",X"47",X"0C",X"FF",X"26",X"10",X"09",X"62",X"30",X"18",X"09",X"64",X"20",X"30",X"08",
		X"66",X"2C",X"38",X"09",X"68",X"FF",X"17",X"28",X"09",X"6A",X"1F",X"18",X"49",X"E0",X"2F",X"10",
		X"49",X"E4",X"FF",X"20",X"11",X"08",X"6C",X"1F",X"31",X"49",X"28",X"22",X"41",X"49",X"29",X"2F",
		X"15",X"09",X"6E",X"2F",X"35",X"49",X"2A",X"FF",X"17",X"22",X"09",X"6A",X"1F",X"12",X"49",X"E0",
		X"2F",X"0A",X"49",X"E4",X"FF",X"7D",X"6E",X"92",X"6E",X"A3",X"6E",X"92",X"6E",X"B8",X"6E",X"CD",
		X"6E",X"7D",X"6E",X"EA",X"6E",X"FF",X"6E",X"7D",X"6E",X"18",X"6F",X"31",X"6F",X"28",X"48",X"8E",
		X"20",X"29",X"30",X"8F",X"22",X"2B",X"38",X"8E",X"01",X"21",X"10",X"8F",X"24",X"31",X"10",X"8F",
		X"26",X"FF",X"28",X"48",X"8E",X"28",X"28",X"30",X"90",X"2A",X"28",X"10",X"8F",X"2C",X"18",X"10",
		X"8F",X"02",X"FF",X"28",X"48",X"8E",X"2E",X"28",X"38",X"8E",X"03",X"2B",X"30",X"8F",X"04",X"21",
		X"10",X"8F",X"30",X"31",X"10",X"8F",X"32",X"FF",X"2C",X"40",X"8E",X"34",X"26",X"30",X"8E",X"36",
		X"28",X"30",X"8F",X"05",X"1D",X"10",X"8F",X"38",X"2D",X"10",X"8F",X"3A",X"FF",X"2B",X"50",X"8E",
		X"06",X"23",X"30",X"8E",X"3C",X"32",X"40",X"8E",X"07",X"3F",X"40",X"8E",X"08",X"29",X"30",X"8F",
		X"0A",X"1B",X"10",X"8F",X"3E",X"2B",X"10",X"8F",X"40",X"FF",X"29",X"40",X"8E",X"42",X"24",X"30",
		X"8E",X"44",X"27",X"30",X"8F",X"09",X"1C",X"10",X"8F",X"46",X"2C",X"10",X"8F",X"48",X"FF",X"29",
		X"40",X"8E",X"4A",X"23",X"30",X"8E",X"4C",X"21",X"10",X"8F",X"4E",X"29",X"20",X"8F",X"50",X"39",
		X"30",X"8F",X"0B",X"49",X"31",X"8F",X"0C",X"FF",X"2B",X"45",X"8E",X"52",X"23",X"33",X"90",X"54",
		X"2C",X"2E",X"90",X"56",X"25",X"2D",X"8F",X"0D",X"2C",X"0E",X"8F",X"58",X"3C",X"15",X"8F",X"5A",
		X"FF",X"2B",X"3C",X"8E",X"5C",X"29",X"1D",X"8F",X"5E",X"1B",X"1C",X"4E",X"A6",X"39",X"0C",X"4F",
		X"AA",X"47",X"1C",X"8F",X"80",X"2B",X"4C",X"8F",X"0F",X"29",X"2D",X"8E",X"0E",X"FF",X"68",X"6F",
		X"7D",X"6F",X"92",X"6F",X"7D",X"6F",X"FB",X"6F",X"0C",X"70",X"EE",X"6F",X"1D",X"70",X"32",X"70",
		X"C0",X"6F",X"D9",X"6F",X"92",X"6F",X"AB",X"6F",X"1D",X"48",X"83",X"E8",X"28",X"40",X"87",X"15",
		X"21",X"10",X"53",X"9C",X"31",X"20",X"93",X"9A",X"31",X"10",X"94",X"9C",X"FF",X"1D",X"48",X"83",
		X"E8",X"28",X"40",X"87",X"15",X"1F",X"30",X"93",X"9E",X"2F",X"20",X"93",X"A0",X"27",X"10",X"94",
		X"A2",X"FF",X"1D",X"48",X"83",X"E8",X"28",X"40",X"87",X"15",X"21",X"30",X"93",X"A4",X"31",X"20",
		X"93",X"A6",X"26",X"10",X"94",X"A8",X"36",X"10",X"94",X"16",X"FF",X"29",X"3F",X"87",X"15",X"24",
		X"30",X"93",X"18",X"33",X"31",X"93",X"17",X"24",X"10",X"94",X"AA",X"34",X"10",X"94",X"AC",X"FF",
		X"13",X"28",X"83",X"E9",X"2A",X"37",X"87",X"15",X"20",X"29",X"93",X"19",X"30",X"19",X"93",X"AE",
		X"25",X"10",X"94",X"B0",X"35",X"10",X"94",X"1A",X"FF",X"2A",X"37",X"87",X"15",X"24",X"28",X"93",
		X"1B",X"34",X"18",X"93",X"B2",X"23",X"10",X"94",X"B4",X"33",X"10",X"94",X"B6",X"FF",X"28",X"2B",
		X"93",X"B8",X"28",X"28",X"93",X"1C",X"28",X"10",X"94",X"BA",X"FF",X"28",X"3E",X"87",X"1D",X"24",
		X"1E",X"93",X"BC",X"28",X"10",X"94",X"BE",X"31",X"0B",X"93",X"1E",X"FF",X"2B",X"3B",X"87",X"1F",
		X"21",X"28",X"93",X"C0",X"31",X"2B",X"93",X"C2",X"24",X"10",X"94",X"C4",X"FF",X"26",X"35",X"87",
		X"E0",X"20",X"19",X"93",X"C6",X"30",X"29",X"93",X"E1",X"2B",X"13",X"94",X"C8",X"3B",X"10",X"94",
		X"CA",X"FF",X"18",X"2A",X"87",X"E2",X"20",X"14",X"93",X"CC",X"2C",X"31",X"93",X"CE",X"2C",X"13",
		X"94",X"D0",X"3C",X"10",X"94",X"D2",X"FF",X"BB",X"70",X"AA",X"70",X"95",X"70",X"AA",X"70",X"D0",
		X"70",X"E9",X"70",X"02",X"71",X"1B",X"71",X"BB",X"71",X"D0",X"71",X"E5",X"71",X"8B",X"71",X"70",
		X"71",X"79",X"71",X"82",X"71",X"0D",X"75",X"12",X"75",X"1B",X"75",X"2D",X"75",X"82",X"71",X"79",
		X"71",X"70",X"71",X"8B",X"71",X"94",X"71",X"A1",X"71",X"AE",X"71",X"34",X"71",X"49",X"71",X"56",
		X"71",X"63",X"71",X"0D",X"75",X"12",X"75",X"1B",X"75",X"2D",X"75",X"63",X"71",X"56",X"71",X"49",
		X"71",X"34",X"71",X"BE",X"66",X"26",X"38",X"D6",X"00",X"1E",X"20",X"D7",X"20",X"2E",X"20",X"D7",
		X"22",X"1E",X"10",X"D6",X"02",X"2E",X"10",X"D6",X"03",X"FF",X"26",X"38",X"D6",X"00",X"1D",X"20",
		X"D7",X"24",X"2D",X"20",X"D7",X"26",X"21",X"10",X"D6",X"01",X"FF",X"26",X"38",X"D6",X"00",X"1E",
		X"20",X"D7",X"20",X"2E",X"20",X"D7",X"22",X"1E",X"10",X"D6",X"28",X"2E",X"10",X"D6",X"2A",X"FF",
		X"2C",X"38",X"D6",X"00",X"24",X"20",X"D7",X"2C",X"2B",X"30",X"D6",X"2E",X"34",X"20",X"D6",X"05",
		X"1C",X"10",X"D6",X"0A",X"2C",X"10",X"D6",X"07",X"FF",X"2E",X"38",X"D6",X"00",X"23",X"20",X"D7",
		X"30",X"2F",X"20",X"D7",X"32",X"3F",X"30",X"D6",X"09",X"1C",X"10",X"D6",X"0A",X"2C",X"10",X"D6",
		X"07",X"FF",X"2E",X"38",X"D6",X"00",X"23",X"20",X"D7",X"30",X"2F",X"20",X"D7",X"34",X"3F",X"28",
		X"D6",X"09",X"1C",X"10",X"D6",X"0A",X"2C",X"10",X"D6",X"07",X"FF",X"2E",X"38",X"D6",X"00",X"23",
		X"20",X"D7",X"30",X"2F",X"20",X"D7",X"36",X"3F",X"20",X"D6",X"0C",X"1C",X"10",X"D6",X"0A",X"2C",
		X"10",X"D6",X"07",X"FF",X"28",X"38",X"D6",X"00",X"22",X"20",X"D7",X"38",X"2E",X"32",X"D6",X"14",
		X"2E",X"22",X"D7",X"15",X"26",X"10",X"D6",X"13",X"FF",X"1E",X"28",X"D8",X"3A",X"2E",X"28",X"D8",
		X"3C",X"24",X"10",X"D8",X"3E",X"FF",X"1E",X"28",X"D8",X"40",X"2E",X"28",X"D8",X"42",X"24",X"10",
		X"D8",X"44",X"FF",X"1E",X"28",X"D8",X"46",X"2E",X"28",X"D8",X"48",X"24",X"10",X"D8",X"4A",X"FF",
		X"22",X"30",X"D8",X"16",X"22",X"10",X"D8",X"4C",X"FF",X"22",X"30",X"D8",X"17",X"22",X"10",X"D8",
		X"4E",X"FF",X"22",X"30",X"D8",X"18",X"22",X"10",X"D8",X"50",X"FF",X"22",X"20",X"D7",X"52",X"22",
		X"10",X"D6",X"19",X"FF",X"25",X"31",X"D6",X"1A",X"22",X"20",X"D7",X"52",X"22",X"10",X"D6",X"19",
		X"FF",X"27",X"34",X"D6",X"00",X"22",X"20",X"D7",X"52",X"22",X"10",X"D6",X"19",X"FF",X"28",X"38",
		X"D6",X"00",X"22",X"20",X"D7",X"52",X"22",X"10",X"D6",X"19",X"FF",X"27",X"38",X"D6",X"1B",X"23",
		X"20",X"D7",X"54",X"33",X"20",X"D7",X"1C",X"29",X"10",X"D6",X"1D",X"2A",X"27",X"D8",X"1E",X"FF",
		X"23",X"30",X"D6",X"1F",X"1C",X"18",X"D7",X"56",X"29",X"15",X"D7",X"58",X"39",X"10",X"D6",X"5A",
		X"39",X"28",X"D6",X"60",X"FF",X"1E",X"27",X"D6",X"61",X"20",X"16",X"D7",X"5C",X"30",X"13",X"D7",
		X"5E",X"3E",X"10",X"D6",X"80",X"2E",X"30",X"D6",X"62",X"FF",X"38",X"72",X"4D",X"72",X"5A",X"72",
		X"4D",X"72",X"6B",X"72",X"80",X"72",X"6B",X"72",X"C3",X"72",X"D8",X"72",X"C3",X"72",X"6B",X"72",
		X"6B",X"72",X"95",X"72",X"AA",X"72",X"95",X"72",X"6B",X"72",X"ED",X"72",X"FE",X"72",X"13",X"73",
		X"FE",X"72",X"ED",X"72",X"46",X"73",X"57",X"73",X"2C",X"73",X"39",X"73",X"8A",X"73",X"68",X"73",
		X"75",X"73",X"9B",X"73",X"AC",X"73",X"BD",X"73",X"26",X"47",X"D9",X"68",X"24",X"30",X"D9",X"82",
		X"2C",X"27",X"D9",X"69",X"20",X"10",X"DA",X"84",X"30",X"10",X"DA",X"86",X"FF",X"26",X"48",X"D9",
		X"04",X"26",X"28",X"D9",X"88",X"26",X"10",X"DA",X"8A",X"FF",X"26",X"47",X"D9",X"04",X"26",X"27",
		X"D9",X"8C",X"1D",X"10",X"DA",X"8E",X"2D",X"10",X"DA",X"90",X"FF",X"25",X"45",X"D9",X"06",X"24",
		X"26",X"D9",X"92",X"34",X"30",X"D9",X"94",X"21",X"10",X"DA",X"96",X"31",X"10",X"DA",X"98",X"FF",
		X"25",X"47",X"D9",X"06",X"24",X"28",X"D9",X"9A",X"24",X"10",X"DA",X"9E",X"34",X"10",X"DA",X"0B",
		X"34",X"3A",X"D9",X"9C",X"FF",X"23",X"47",X"D9",X"04",X"22",X"27",X"D9",X"A0",X"32",X"36",X"D9",
		X"67",X"1C",X"10",X"DA",X"A2",X"2C",X"1E",X"DA",X"A4",X"FF",X"1D",X"48",X"D9",X"06",X"1C",X"28",
		X"D9",X"A6",X"2C",X"28",X"D9",X"A8",X"3A",X"3C",X"DA",X"6A",X"4A",X"3C",X"DA",X"6B",X"1F",X"10",
		X"DA",X"AA",X"FF",X"25",X"46",X"D9",X"04",X"24",X"26",X"D9",X"AC",X"34",X"38",X"D9",X"6C",X"25",
		X"10",X"DA",X"AE",X"35",X"10",X"DA",X"6D",X"FF",X"28",X"47",X"D9",X"04",X"26",X"27",X"D9",X"B0",
		X"36",X"38",X"D9",X"6E",X"21",X"10",X"DA",X"B2",X"31",X"10",X"DA",X"B4",X"FF",X"1C",X"20",X"D9",
		X"B6",X"2C",X"20",X"D9",X"B8",X"1C",X"10",X"DA",X"6F",X"2C",X"10",X"DA",X"70",X"FF",X"2A",X"30",
		X"D9",X"71",X"20",X"1C",X"D9",X"BA",X"30",X"1A",X"D9",X"BC",X"1F",X"10",X"DA",X"72",X"33",X"10",
		X"DA",X"73",X"FF",X"25",X"2C",X"D9",X"74",X"1F",X"10",X"D9",X"BE",X"2F",X"10",X"D9",X"C0",X"1D",
		X"10",X"DA",X"75",X"3D",X"10",X"DA",X"76",X"4D",X"10",X"DA",X"6D",X"FF",X"29",X"50",X"D9",X"68",
		X"25",X"30",X"D9",X"C2",X"25",X"10",X"DA",X"C4",X"FF",X"28",X"44",X"D9",X"77",X"22",X"24",X"D9",
		X"C6",X"24",X"14",X"DA",X"C8",X"FF",X"26",X"30",X"D9",X"CA",X"2D",X"33",X"D9",X"CC",X"1F",X"10",
		X"DA",X"CE",X"2F",X"10",X"DA",X"D0",X"FF",X"26",X"31",X"D9",X"D2",X"25",X"28",X"D9",X"78",X"1D",
		X"10",X"DA",X"79",X"27",X"10",X"DA",X"D4",X"FF",X"29",X"30",X"D9",X"D6",X"19",X"27",X"D9",X"D8",
		X"26",X"10",X"DA",X"DA",X"FF",X"23",X"33",X"D9",X"DC",X"23",X"23",X"D9",X"7A",X"27",X"10",X"DA",
		X"DE",X"37",X"10",X"DA",X"7C",X"33",X"3E",X"DA",X"7B",X"FF",X"2B",X"30",X"D9",X"E0",X"20",X"28",
		X"D9",X"E2",X"25",X"10",X"DA",X"E4",X"31",X"0C",X"DA",X"7D",X"FF",X"28",X"29",X"D9",X"E6",X"23",
		X"23",X"D9",X"E8",X"2E",X"10",X"DA",X"EA",X"3E",X"10",X"DA",X"7E",X"FF",X"1D",X"1B",X"D9",X"EC",
		X"18",X"10",X"D9",X"7F",X"28",X"10",X"D9",X"EE",X"38",X"11",X"DA",X"F0",X"FF",X"24",X"3A",X"99",
		X"66",X"22",X"28",X"99",X"68",X"26",X"0F",X"9A",X"6A",X"32",X"2F",X"9A",X"6E",X"42",X"2F",X"9A",
		X"70",X"FF",X"DC",X"73",X"E1",X"73",X"E6",X"73",X"EB",X"73",X"DC",X"73",X"28",X"10",X"D6",X"63",
		X"FF",X"28",X"10",X"D6",X"64",X"FF",X"28",X"10",X"D6",X"65",X"FF",X"28",X"10",X"D6",X"66",X"FF",
		X"00",X"74",X"0D",X"74",X"1A",X"74",X"0D",X"74",X"27",X"74",X"38",X"74",X"4D",X"74",X"7F",X"74",
		X"28",X"3B",X"1B",X"39",X"27",X"2B",X"1C",X"3A",X"28",X"10",X"9C",X"60",X"FF",X"28",X"3C",X"1B",
		X"39",X"28",X"2C",X"9C",X"FA",X"28",X"10",X"9C",X"62",X"FF",X"28",X"3C",X"9B",X"FD",X"29",X"2C",
		X"9C",X"FE",X"27",X"10",X"9C",X"64",X"FF",X"1F",X"32",X"1B",X"2F",X"1E",X"1A",X"1C",X"5E",X"25",
		X"0E",X"9C",X"DC",X"1E",X"26",X"1D",X"20",X"FF",X"23",X"32",X"1B",X"38",X"1F",X"1A",X"9C",X"DE",
		X"25",X"0E",X"1C",X"5A",X"23",X"2E",X"9D",X"F9",X"1C",X"23",X"1D",X"1E",X"FF",X"23",X"32",X"1B",
		X"38",X"1F",X"1A",X"9C",X"DE",X"25",X"0E",X"1C",X"5A",X"17",X"20",X"1D",X"0C",X"27",X"20",X"1D",
		X"18",X"29",X"2B",X"9D",X"FF",X"FF",X"23",X"38",X"1B",X"23",X"25",X"30",X"1C",X"30",X"1E",X"10",
		X"9C",X"74",X"25",X"40",X"80",X"76",X"25",X"30",X"81",X"78",X"2B",X"10",X"82",X"7A",X"FF",X"28",
		X"04",X"9D",X"6C",X"FF",X"2B",X"0A",X"47",X"0C",X"FF",X"2B",X"0A",X"4B",X"0C",X"FF",X"CC",X"74",
		X"D1",X"74",X"D6",X"74",X"DB",X"74",X"CC",X"74",X"E0",X"74",X"E9",X"74",X"F2",X"74",X"FF",X"74",
		X"04",X"75",X"61",X"75",X"6A",X"75",X"73",X"75",X"0D",X"75",X"12",X"75",X"1B",X"75",X"20",X"75",
		X"43",X"75",X"4C",X"75",X"43",X"75",X"78",X"75",X"7D",X"75",X"32",X"75",X"20",X"75",X"2D",X"75",
		X"82",X"75",X"87",X"75",X"8C",X"75",X"91",X"75",X"96",X"75",X"9B",X"75",X"28",X"10",X"0A",X"70",
		X"FF",X"28",X"10",X"4D",X"35",X"FF",X"28",X"10",X"4B",X"3A",X"FF",X"28",X"10",X"4B",X"3C",X"FF",
		X"20",X"10",X"4A",X"2C",X"30",X"10",X"4A",X"2D",X"FF",X"20",X"10",X"4A",X"2E",X"30",X"10",X"4A",
		X"2F",X"FF",X"28",X"10",X"4B",X"32",X"20",X"10",X"4A",X"30",X"30",X"10",X"4A",X"31",X"FF",X"28",
		X"10",X"4B",X"32",X"FF",X"21",X"10",X"4B",X"33",X"31",X"10",X"4B",X"34",X"FF",X"28",X"10",X"0C",
		X"72",X"FF",X"28",X"10",X"0C",X"74",X"28",X"30",X"4C",X"36",X"FF",X"28",X"10",X"4C",X"EC",X"FF",
		X"26",X"17",X"4C",X"F0",X"36",X"2F",X"0C",X"76",X"28",X"0F",X"4C",X"E8",X"FF",X"28",X"0F",X"4C",
		X"E8",X"FF",X"26",X"17",X"4C",X"F0",X"36",X"2F",X"0C",X"76",X"21",X"35",X"0C",X"78",X"31",X"35",
		X"0C",X"7A",X"FF",X"26",X"17",X"4C",X"F0",X"36",X"2F",X"0C",X"76",X"FF",X"26",X"17",X"4C",X"F0",
		X"36",X"2F",X"0C",X"76",X"38",X"3F",X"4C",X"37",X"48",X"3F",X"4C",X"38",X"58",X"3F",X"4C",X"39",
		X"FF",X"20",X"08",X"0C",X"78",X"30",X"08",X"0C",X"7A",X"FF",X"20",X"08",X"0C",X"7C",X"30",X"08",
		X"0C",X"7E",X"FF",X"28",X"08",X"0C",X"40",X"FF",X"2B",X"0D",X"4B",X"3B",X"FF",X"2B",X"0D",X"4B",
		X"3D",X"FF",X"2C",X"0E",X"D8",X"0D",X"FF",X"2C",X"0E",X"D8",X"0E",X"FF",X"2C",X"0D",X"D8",X"0F",
		X"FF",X"2C",X"0D",X"D8",X"10",X"FF",X"28",X"10",X"D8",X"11",X"FF",X"28",X"10",X"D8",X"12",X"FF",
		X"24",X"09",X"01",X"01",X"FF",X"B1",X"75",X"B6",X"75",X"BB",X"75",X"B6",X"75",X"B1",X"75",X"BB",
		X"75",X"28",X"10",X"83",X"E3",X"FF",X"28",X"10",X"83",X"E4",X"FF",X"28",X"10",X"83",X"E5",X"FF",
		X"D4",X"75",X"D9",X"75",X"DE",X"75",X"E3",X"75",X"E8",X"75",X"ED",X"75",X"F2",X"75",X"61",X"75",
		X"6A",X"75",X"73",X"75",X"28",X"10",X"95",X"D4",X"FF",X"28",X"10",X"95",X"E6",X"FF",X"28",X"10",
		X"95",X"D6",X"FF",X"28",X"10",X"95",X"D8",X"FF",X"28",X"03",X"95",X"D6",X"FF",X"28",X"03",X"95",
		X"D8",X"FF",X"28",X"10",X"95",X"E7",X"FF",X"11",X"76",X"16",X"76",X"1B",X"76",X"20",X"76",X"25",
		X"76",X"2A",X"76",X"2F",X"76",X"34",X"76",X"3D",X"76",X"46",X"76",X"4F",X"76",X"58",X"76",X"61",
		X"76",X"28",X"10",X"8C",X"F0",X"FF",X"28",X"10",X"8C",X"F1",X"FF",X"27",X"10",X"8C",X"F2",X"FF",
		X"28",X"10",X"8C",X"F3",X"FF",X"28",X"10",X"8C",X"F4",X"FF",X"28",X"10",X"8C",X"F5",X"FF",X"28",
		X"10",X"8C",X"F6",X"FF",X"24",X"10",X"8C",X"F8",X"2A",X"10",X"8C",X"F7",X"FF",X"25",X"10",X"8C",
		X"F0",X"2A",X"10",X"8C",X"F7",X"FF",X"25",X"10",X"8C",X"F1",X"2A",X"10",X"8C",X"F7",X"FF",X"25",
		X"10",X"8C",X"F3",X"2A",X"10",X"8C",X"F7",X"FF",X"21",X"10",X"8C",X"F8",X"2C",X"10",X"8C",X"F7",
		X"FF",X"28",X"10",X"8C",X"F8",X"FF",X"3E",X"FF",X"32",X"00",X"E0",X"FB",X"CD",X"0D",X"57",X"CD",
		X"57",X"11",X"F3",X"DD",X"21",X"00",X"00",X"06",X"00",X"3E",X"00",X"5F",X"16",X"0D",X"0E",X"10",
		X"21",X"00",X"E0",X"77",X"23",X"3C",X"15",X"20",X"03",X"16",X"0D",X"3C",X"10",X"F5",X"0D",X"20",
		X"F2",X"7B",X"21",X"00",X"E0",X"16",X"0D",X"0E",X"10",X"BE",X"C2",X"F6",X"77",X"23",X"3C",X"15",
		X"20",X"03",X"16",X"0D",X"3C",X"10",X"F2",X"0D",X"20",X"EF",X"7B",X"3C",X"FE",X"14",X"20",X"CB",
		X"3E",X"00",X"5F",X"16",X"0D",X"0E",X"10",X"21",X"00",X"D0",X"77",X"23",X"3C",X"15",X"20",X"03",
		X"16",X"0D",X"3C",X"10",X"F5",X"0D",X"20",X"F2",X"7B",X"21",X"00",X"D0",X"16",X"0D",X"0E",X"10",
		X"BE",X"C2",X"BD",X"77",X"23",X"3C",X"15",X"20",X"03",X"16",X"0D",X"3C",X"10",X"F2",X"0D",X"20",
		X"EF",X"7B",X"3C",X"FE",X"14",X"20",X"CB",X"CD",X"57",X"11",X"21",X"00",X"E0",X"11",X"01",X"E0",
		X"01",X"FF",X"0F",X"36",X"00",X"ED",X"B0",X"21",X"25",X"EB",X"22",X"03",X"EB",X"3E",X"FF",X"32",
		X"00",X"E0",X"11",X"00",X"00",X"CD",X"10",X"7C",X"ED",X"4B",X"6A",X"00",X"AF",X"ED",X"42",X"28",
		X"01",X"3C",X"CD",X"10",X"7C",X"ED",X"4B",X"6C",X"00",X"ED",X"42",X"28",X"02",X"CB",X"CF",X"F5",
		X"47",X"0E",X"14",X"11",X"D5",X"D1",X"3E",X"31",X"CD",X"F7",X"7B",X"11",X"55",X"D2",X"3E",X"32",
		X"CD",X"F7",X"7B",X"DD",X"E5",X"E1",X"7D",X"B4",X"11",X"55",X"D1",X"21",X"89",X"78",X"20",X"03",
		X"21",X"91",X"78",X"CD",X"1C",X"11",X"FB",X"3E",X"70",X"CD",X"0F",X"57",X"78",X"A7",X"C4",X"E8",
		X"7B",X"CD",X"57",X"11",X"21",X"F7",X"7C",X"CD",X"1C",X"11",X"AF",X"32",X"82",X"E8",X"3A",X"1D",
		X"E8",X"32",X"1D",X"E8",X"0E",X"00",X"CD",X"D7",X"7B",X"3A",X"06",X"E9",X"E6",X"03",X"21",X"82",
		X"E8",X"28",X"25",X"47",X"7E",X"A7",X"20",X"22",X"36",X"10",X"0E",X"14",X"3A",X"1D",X"E8",X"F5",
		X"CD",X"D7",X"7B",X"F1",X"CB",X"48",X"20",X"08",X"3D",X"F2",X"61",X"77",X"3E",X"05",X"18",X"D1",
		X"3C",X"FE",X"06",X"38",X"CC",X"AF",X"18",X"C9",X"36",X"00",X"3A",X"04",X"E9",X"CB",X"47",X"28",
		X"C8",X"CD",X"57",X"11",X"21",X"51",X"77",X"E5",X"3A",X"1D",X"E8",X"21",X"B1",X"77",X"C3",X"26",
		X"1F",X"99",X"78",X"3E",X"79",X"BA",X"79",X"8B",X"7A",X"10",X"7B",X"78",X"7B",X"08",X"D9",X"11",
		X"00",X"E0",X"21",X"55",X"D1",X"01",X"20",X"00",X"ED",X"B0",X"11",X"20",X"E0",X"21",X"55",X"D9",
		X"01",X"20",X"00",X"ED",X"B0",X"DD",X"21",X"DB",X"77",X"18",X"21",X"D9",X"21",X"00",X"E0",X"11",
		X"55",X"D1",X"01",X"20",X"00",X"ED",X"B0",X"21",X"20",X"E0",X"11",X"55",X"D9",X"01",X"20",X"00",
		X"ED",X"B0",X"D9",X"C3",X"D4",X"76",X"DD",X"21",X"9D",X"76",X"08",X"D9",X"21",X"55",X"D1",X"11",
		X"89",X"78",X"06",X"07",X"1A",X"13",X"FD",X"21",X"0C",X"78",X"18",X"73",X"10",X"F6",X"3E",X"3A",
		X"FD",X"21",X"16",X"78",X"18",X"69",X"D9",X"7C",X"D9",X"FD",X"21",X"1F",X"78",X"18",X"42",X"D9",
		X"7D",X"D9",X"FD",X"21",X"28",X"78",X"18",X"39",X"3E",X"3A",X"FD",X"21",X"30",X"78",X"18",X"4F",
		X"08",X"5F",X"08",X"7B",X"FD",X"21",X"3A",X"78",X"18",X"27",X"23",X"D9",X"7E",X"D9",X"FD",X"21",
		X"44",X"78",X"18",X"1D",X"DB",X"00",X"CB",X"47",X"CA",X"E7",X"76",X"CB",X"4F",X"20",X"F5",X"01",
		X"00",X"10",X"0B",X"79",X"B0",X"20",X"FB",X"DB",X"00",X"CB",X"4F",X"28",X"FA",X"D9",X"08",X"DD",
		X"E9",X"5F",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"C6",X"90",X"27",X"CE",X"40",X"27",X"77",X"CB",
		X"DC",X"36",X"14",X"CB",X"9C",X"23",X"7B",X"E6",X"0F",X"C6",X"90",X"27",X"CE",X"40",X"27",X"77",
		X"CB",X"DC",X"36",X"14",X"CB",X"9C",X"23",X"FD",X"E9",X"52",X"41",X"4D",X"20",X"20",X"4E",X"47",
		X"FF",X"52",X"41",X"4D",X"20",X"20",X"4F",X"4B",X"FF",X"21",X"30",X"7C",X"CD",X"1C",X"11",X"CD",
		X"C1",X"7B",X"CD",X"1C",X"11",X"11",X"99",X"D1",X"DB",X"03",X"CD",X"B2",X"7B",X"11",X"D9",X"D1",
		X"DB",X"04",X"CD",X"B2",X"7B",X"DB",X"04",X"CB",X"4F",X"21",X"96",X"7C",X"20",X"03",X"21",X"9E",
		X"7C",X"11",X"5D",X"D3",X"CD",X"1C",X"11",X"DB",X"03",X"E6",X"01",X"21",X"A6",X"7C",X"20",X"03",
		X"21",X"B0",X"7C",X"11",X"9E",X"D3",X"CD",X"1C",X"11",X"DB",X"03",X"E6",X"02",X"21",X"BA",X"7C",
		X"20",X"03",X"21",X"BF",X"7C",X"11",X"DE",X"D3",X"CD",X"1C",X"11",X"CD",X"6F",X"05",X"11",X"1F",
		X"D4",X"CD",X"08",X"11",X"CD",X"8F",X"05",X"41",X"11",X"9A",X"D2",X"2A",X"0A",X"E9",X"7D",X"A7",
		X"28",X"28",X"BC",X"F5",X"3E",X"20",X"28",X"02",X"3E",X"41",X"CD",X"10",X"11",X"CD",X"F7",X"49",
		X"F1",X"11",X"D0",X"D2",X"28",X"1D",X"E5",X"21",X"8C",X"7C",X"CD",X"1C",X"11",X"13",X"3E",X"42",
		X"CD",X"10",X"11",X"E1",X"6C",X"CD",X"F7",X"49",X"18",X"0C",X"21",X"C4",X"7C",X"CD",X"1C",X"11",
		X"11",X"D0",X"D2",X"CD",X"1A",X"57",X"DB",X"00",X"CB",X"4F",X"C2",X"A5",X"78",X"C9",X"01",X"14",
		X"03",X"11",X"55",X"D4",X"C5",X"21",X"D8",X"7C",X"CD",X"1C",X"11",X"E5",X"13",X"78",X"CD",X"08",
		X"11",X"CD",X"C1",X"7B",X"21",X"2C",X"00",X"19",X"EB",X"E1",X"CD",X"1C",X"11",X"21",X"B6",X"FE",
		X"19",X"EB",X"C1",X"10",X"DF",X"21",X"EC",X"7C",X"CD",X"1C",X"11",X"21",X"99",X"99",X"22",X"03",
		X"E0",X"3E",X"38",X"32",X"82",X"E8",X"21",X"03",X"E0",X"7E",X"C6",X"01",X"27",X"77",X"23",X"7E",
		X"CE",X"00",X"27",X"77",X"11",X"62",X"D5",X"CD",X"FD",X"10",X"CD",X"FD",X"10",X"DB",X"00",X"11",
		X"A2",X"D2",X"CD",X"B2",X"7B",X"DB",X"01",X"11",X"A2",X"D3",X"CD",X"B2",X"7B",X"DB",X"02",X"11",
		X"A2",X"D4",X"CD",X"B2",X"7B",X"3A",X"82",X"E8",X"A7",X"28",X"C6",X"3A",X"04",X"E9",X"CB",X"4F",
		X"28",X"DB",X"3A",X"06",X"E9",X"CB",X"4F",X"28",X"D4",X"C9",X"AF",X"32",X"82",X"E8",X"F5",X"21",
		X"61",X"7A",X"5F",X"16",X"00",X"19",X"19",X"3A",X"04",X"E9",X"CB",X"47",X"20",X"F9",X"7E",X"32",
		X"83",X"E8",X"32",X"1F",X"E8",X"23",X"3E",X"00",X"CD",X"FE",X"0D",X"7E",X"CD",X"FE",X"0D",X"21",
		X"56",X"7D",X"CD",X"1C",X"11",X"F1",X"32",X"1E",X"E8",X"0E",X"00",X"CD",X"CE",X"7B",X"3A",X"06",
		X"E9",X"E6",X"03",X"21",X"82",X"E8",X"28",X"2E",X"47",X"7E",X"A7",X"20",X"F1",X"3E",X"00",X"CD",
		X"FE",X"0D",X"AF",X"32",X"1F",X"E8",X"36",X"10",X"0E",X"14",X"3A",X"1E",X"E8",X"F5",X"CD",X"CE",
		X"7B",X"F1",X"CB",X"48",X"20",X"08",X"3D",X"F2",X"E6",X"79",X"3E",X"14",X"18",X"C8",X"3C",X"FE",
		X"15",X"38",X"C3",X"AF",X"18",X"C0",X"36",X"00",X"3A",X"1F",X"E8",X"A7",X"28",X"12",X"47",X"3A",
		X"83",X"E8",X"A7",X"28",X"11",X"3A",X"04",X"E9",X"E6",X"03",X"28",X"B2",X"CB",X"4F",X"20",X"1B",
		X"3A",X"1E",X"E8",X"C3",X"BE",X"79",X"78",X"FE",X"BA",X"32",X"83",X"E8",X"3E",X"01",X"32",X"1F",
		X"E8",X"30",X"9B",X"3A",X"1E",X"E8",X"3C",X"FE",X"15",X"38",X"E8",X"3E",X"00",X"CD",X"FE",X"0D",
		X"C9",X"2D",X"01",X"2D",X"02",X"2D",X"03",X"B4",X"05",X"9E",X"04",X"2D",X"06",X"2D",X"07",X"2D",
		X"10",X"2D",X"11",X"2D",X"12",X"2D",X"13",X"2D",X"14",X"2D",X"15",X"2D",X"16",X"BA",X"20",X"FF",
		X"24",X"BA",X"22",X"FF",X"23",X"BA",X"21",X"2D",X"17",X"2D",X"18",X"CD",X"53",X"11",X"21",X"00",
		X"E0",X"36",X"FE",X"3A",X"06",X"E9",X"E6",X"03",X"28",X"0A",X"CB",X"4F",X"28",X"04",X"36",X"FD",
		X"18",X"02",X"36",X"FE",X"3A",X"04",X"E9",X"CB",X"4F",X"28",X"E8",X"36",X"FF",X"C9",X"0E",X"00",
		X"3C",X"20",X"32",X"21",X"10",X"01",X"11",X"E0",X"00",X"3E",X"00",X"CD",X"DC",X"7A",X"21",X"10",
		X"01",X"11",X"20",X"01",X"3E",X"40",X"CD",X"DC",X"7A",X"21",X"D0",X"00",X"11",X"E0",X"00",X"3E",
		X"80",X"CD",X"DC",X"7A",X"21",X"D0",X"00",X"11",X"20",X"01",X"3E",X"C0",X"22",X"07",X"E8",X"21",
		X"DE",X"75",X"C3",X"20",X"0E",X"21",X"C0",X"00",X"22",X"07",X"E8",X"11",X"D0",X"00",X"21",X"9B",
		X"66",X"CD",X"0C",X"7B",X"11",X"F0",X"00",X"21",X"6A",X"6C",X"CD",X"0C",X"7B",X"11",X"10",X"01",
		X"21",X"7D",X"6E",X"CD",X"0C",X"7B",X"11",X"30",X"01",X"21",X"6B",X"72",X"AF",X"C3",X"20",X"0E",
		X"11",X"D0",X"D1",X"0E",X"14",X"3E",X"41",X"06",X"1A",X"CD",X"C7",X"7B",X"11",X"10",X"D2",X"3E",
		X"30",X"06",X"0A",X"CD",X"C7",X"7B",X"CD",X"E8",X"7B",X"3E",X"04",X"11",X"04",X"00",X"CD",X"5B",
		X"11",X"CD",X"E8",X"7B",X"1E",X"01",X"CD",X"5B",X"11",X"CD",X"E8",X"7B",X"1E",X"02",X"CD",X"5B",
		X"11",X"CD",X"E8",X"7B",X"01",X"00",X"02",X"1E",X"06",X"CD",X"5E",X"11",X"01",X"00",X"04",X"1E",
		X"00",X"CD",X"65",X"11",X"01",X"00",X"02",X"1E",X"07",X"CD",X"65",X"11",X"21",X"10",X"D4",X"0E",
		X"08",X"3E",X"00",X"06",X"04",X"77",X"23",X"10",X"FC",X"3C",X"E6",X"07",X"20",X"F5",X"11",X"20",
		X"00",X"19",X"0D",X"20",X"EC",X"C3",X"E8",X"7B",X"0E",X"00",X"11",X"10",X"D0",X"3E",X"0B",X"2E",
		X"20",X"E5",X"06",X"10",X"CD",X"10",X"11",X"3D",X"CD",X"10",X"11",X"3C",X"10",X"F6",X"21",X"20",
		X"00",X"19",X"EB",X"FE",X"0B",X"3E",X"0B",X"20",X"02",X"3E",X"09",X"E1",X"2D",X"20",X"E2",X"21",
		X"DF",X"D3",X"36",X"0C",X"23",X"36",X"0D",X"21",X"1F",X"D4",X"36",X"0E",X"23",X"36",X"0F",X"C3",
		X"E8",X"7B",X"2F",X"6F",X"06",X"08",X"AF",X"CB",X"0D",X"CB",X"17",X"CD",X"08",X"11",X"10",X"F6",
		X"C9",X"13",X"13",X"3E",X"31",X"06",X"08",X"CD",X"10",X"11",X"3C",X"10",X"FA",X"C9",X"FE",X"06",
		X"38",X"01",X"3C",X"A7",X"28",X"01",X"3C",X"6F",X"26",X"00",X"29",X"29",X"29",X"29",X"29",X"29",
		X"11",X"50",X"D9",X"19",X"71",X"23",X"71",X"C9",X"3A",X"04",X"E9",X"CB",X"4F",X"28",X"F9",X"3A",
		X"04",X"E9",X"CB",X"4F",X"20",X"F9",X"C9",X"F5",X"21",X"2C",X"7C",X"CD",X"1C",X"11",X"F1",X"CD",
		X"10",X"11",X"13",X"21",X"29",X"7C",X"CB",X"08",X"38",X"03",X"21",X"26",X"7C",X"C3",X"1C",X"11",
		X"F5",X"01",X"00",X"40",X"21",X"00",X"00",X"1A",X"85",X"6F",X"3E",X"00",X"8C",X"67",X"13",X"0B",
		X"79",X"B0",X"20",X"F3",X"F1",X"C9",X"4F",X"4B",X"FF",X"4E",X"47",X"FF",X"52",X"4F",X"4D",X"FF",
		X"FE",X"14",X"FD",X"50",X"D1",X"44",X"49",X"50",X"20",X"53",X"57",X"20",X"FF",X"FD",X"94",X"D1",
		X"44",X"53",X"57",X"31",X"FD",X"D4",X"D1",X"44",X"53",X"57",X"32",X"FD",X"A3",X"D1",X"31",X"2E",
		X"4F",X"4E",X"FD",X"E3",X"D1",X"30",X"2E",X"4F",X"46",X"46",X"FD",X"50",X"D3",X"42",X"4F",X"44",
		X"59",X"20",X"54",X"59",X"50",X"45",X"FD",X"90",X"D3",X"44",X"49",X"46",X"46",X"49",X"43",X"55",
		X"4C",X"54",X"59",X"FD",X"D0",X"D3",X"44",X"45",X"43",X"52",X"45",X"41",X"53",X"45",X"FD",X"10",
		X"D4",X"46",X"49",X"47",X"48",X"54",X"45",X"52",X"53",X"FD",X"90",X"D2",X"43",X"4F",X"49",X"4E",
		X"20",X"4D",X"4F",X"44",X"45",X"FF",X"54",X"41",X"42",X"4C",X"45",X"20",X"20",X"FF",X"55",X"50",
		X"52",X"49",X"47",X"48",X"54",X"FF",X"45",X"41",X"53",X"59",X"20",X"20",X"20",X"20",X"20",X"FF",
		X"44",X"49",X"46",X"46",X"49",X"43",X"55",X"4C",X"54",X"FF",X"53",X"4C",X"4F",X"57",X"FF",X"46",
		X"41",X"53",X"54",X"FF",X"20",X"20",X"20",X"20",X"20",X"46",X"52",X"45",X"45",X"20",X"20",X"20",
		X"50",X"4C",X"41",X"59",X"20",X"20",X"20",X"FF",X"49",X"4E",X"54",X"45",X"52",X"46",X"41",X"43",
		X"45",X"FF",X"52",X"45",X"41",X"44",X"20",X"44",X"41",X"54",X"41",X"FF",X"FD",X"57",X"D5",X"54",
		X"49",X"4D",X"4D",X"49",X"4E",X"47",X"FF",X"FE",X"14",X"FD",X"50",X"D1",X"30",X"31",X"20",X"44",
		X"49",X"50",X"20",X"53",X"57",X"49",X"54",X"43",X"48",X"FD",X"90",X"D1",X"30",X"32",X"20",X"49",
		X"2F",X"4F",X"20",X"50",X"4F",X"52",X"54",X"FD",X"D0",X"D1",X"30",X"33",X"20",X"53",X"4F",X"55",
		X"4E",X"44",X"FD",X"10",X"D2",X"30",X"34",X"20",X"43",X"48",X"41",X"52",X"41",X"43",X"54",X"45",
		X"52",X"FD",X"50",X"D2",X"30",X"35",X"20",X"43",X"4F",X"4C",X"4F",X"52",X"FD",X"90",X"D2",X"30",
		X"36",X"20",X"43",X"52",X"4F",X"53",X"53",X"20",X"48",X"41",X"54",X"43",X"48",X"20",X"50",X"41",
		X"54",X"54",X"45",X"52",X"4E",X"FF",X"FE",X"14",X"FD",X"15",X"D1",X"53",X"4F",X"55",X"4E",X"44",
		X"FD",X"50",X"D1",X"30",X"31",X"20",X"59",X"45",X"4C",X"4C",X"20",X"4F",X"46",X"20",X"50",X"4C",
		X"41",X"59",X"45",X"52",X"28",X"4A",X"55",X"4D",X"50",X"2D",X"4B",X"49",X"43",X"4B",X"53",X"29",
		X"FD",X"93",X"D1",X"43",X"52",X"45",X"44",X"49",X"54",X"20",X"41",X"44",X"44",X"49",X"4E",X"47",
		X"20",X"53",X"4F",X"55",X"4E",X"44",X"FD",X"D0",X"D1",X"30",X"32",X"20",X"59",X"45",X"4C",X"4C",
		X"20",X"4F",X"46",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"28",X"50",X"55",X"4E",X"43",X"48",
		X"45",X"53",X"2C",X"4B",X"49",X"43",X"4B",X"53",X"29",X"FD",X"10",X"D2",X"30",X"33",X"20",X"47",
		X"52",X"4F",X"41",X"4E",X"20",X"4F",X"46",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"4F",
		X"52",X"20",X"45",X"4E",X"45",X"4D",X"59",X"FD",X"50",X"D2",X"30",X"34",X"20",X"4C",X"41",X"55",
		X"47",X"48",X"49",X"4E",X"47",X"20",X"56",X"4F",X"49",X"43",X"45",X"20",X"4F",X"46",X"20",X"45",
		X"4E",X"45",X"4D",X"49",X"45",X"53",X"2D",X"31",X"FD",X"90",X"D2",X"30",X"35",X"20",X"4C",X"41",
		X"55",X"47",X"48",X"49",X"4E",X"47",X"20",X"56",X"4F",X"49",X"43",X"45",X"20",X"4F",X"46",X"20",
		X"45",X"4E",X"45",X"4D",X"49",X"45",X"53",X"2D",X"32",X"FD",X"D0",X"D2",X"30",X"36",X"20",X"42",
		X"55",X"52",X"53",X"54",X"49",X"4E",X"47",X"20",X"4F",X"46",X"20",X"50",X"41",X"50",X"45",X"52",
		X"20",X"42",X"41",X"4C",X"4C",X"FD",X"13",X"D3",X"42",X"55",X"52",X"53",X"54",X"49",X"4E",X"47",
		X"20",X"4F",X"46",X"20",X"44",X"52",X"41",X"47",X"4F",X"4E",X"27",X"53",X"20",X"45",X"47",X"47",
		X"FD",X"50",X"D3",X"30",X"37",X"20",X"53",X"48",X"52",X"49",X"45",X"4B",X"20",X"4F",X"46",X"20",
		X"50",X"4C",X"41",X"59",X"45",X"52",X"FD",X"90",X"D3",X"30",X"38",X"20",X"50",X"4C",X"41",X"59",
		X"45",X"52",X"20",X"52",X"55",X"4E",X"4E",X"49",X"4E",X"47",X"FD",X"D0",X"D3",X"30",X"39",X"20",
		X"48",X"49",X"54",X"54",X"49",X"4E",X"47",X"20",X"53",X"4F",X"55",X"4E",X"44",X"FD",X"10",X"D4",
		X"31",X"30",X"20",X"53",X"57",X"49",X"53",X"48",X"49",X"4E",X"47",X"20",X"53",X"4F",X"55",X"4E",
		X"44",X"FD",X"50",X"D4",X"31",X"31",X"20",X"42",X"55",X"52",X"53",X"54",X"49",X"4E",X"47",X"20",
		X"4F",X"46",X"20",X"53",X"4E",X"41",X"4B",X"45",X"20",X"50",X"4F",X"54",X"FD",X"90",X"D4",X"31",
		X"32",X"20",X"42",X"49",X"54",X"49",X"4E",X"47",X"20",X"53",X"4F",X"55",X"4E",X"44",X"FD",X"D0",
		X"D4",X"31",X"33",X"20",X"53",X"4F",X"55",X"4E",X"44",X"20",X"4F",X"46",X"20",X"4B",X"4E",X"49",
		X"56",X"45",X"53",X"2C",X"42",X"4F",X"4F",X"4D",X"45",X"52",X"41",X"4E",X"47",X"53",X"FD",X"10",
		X"D5",X"31",X"34",X"20",X"43",X"4F",X"55",X"4E",X"54",X"49",X"4E",X"47",X"20",X"50",X"4F",X"49",
		X"4E",X"54",X"53",X"FD",X"50",X"D5",X"31",X"35",X"20",X"47",X"41",X"4D",X"45",X"20",X"53",X"54",
		X"41",X"52",X"54",X"FD",X"90",X"D5",X"31",X"36",X"20",X"42",X"47",X"4D",X"FD",X"D0",X"D5",X"31",
		X"37",X"20",X"43",X"4F",X"4D",X"50",X"4C",X"45",X"54",X"49",X"4F",X"4E",X"20",X"4F",X"46",X"20",
		X"45",X"41",X"43",X"48",X"20",X"50",X"41",X"54",X"54",X"45",X"52",X"4E",X"FD",X"10",X"D6",X"31",
		X"38",X"20",X"43",X"4F",X"4D",X"50",X"4C",X"45",X"54",X"49",X"4F",X"4E",X"20",X"4F",X"46",X"20",
		X"47",X"41",X"4D",X"45",X"FD",X"50",X"D6",X"31",X"39",X"20",X"47",X"41",X"4D",X"45",X"20",X"4F",
		X"56",X"45",X"52",X"FD",X"90",X"D6",X"32",X"30",X"20",X"54",X"49",X"4D",X"45",X"20",X"55",X"50",
		X"20",X"57",X"41",X"52",X"4E",X"49",X"4E",X"47",X"FD",X"D0",X"D6",X"32",X"31",X"20",X"41",X"44",
		X"44",X"49",X"54",X"49",X"4F",X"4E",X"41",X"4C",X"20",X"46",X"49",X"47",X"48",X"54",X"45",X"52",
		X"FD",X"16",X"D7",X"4D",X"55",X"53",X"49",X"43",X"20",X"45",X"4E",X"44",X"FF",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
