library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity twotiger_sp_bits_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of twotiger_sp_bits_1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"0E",X"FF",X"EE",X"00",X"EE",X"FF",X"FF",X"00",X"EE",X"FF",X"FF",X"00",X"EE",X"EE",X"FF",
		X"00",X"55",X"55",X"EE",X"00",X"55",X"55",X"55",X"00",X"55",X"5E",X"F5",X"00",X"6F",X"E1",X"E5",
		X"00",X"EE",X"EF",X"0E",X"00",X"00",X"0E",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"EF",X"00",X"00",X"F0",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"0E",X"FF",X"00",X"00",X"EE",X"FF",X"00",X"00",X"EE",X"FF",X"EE",X"00",X"E5",X"55",X"FF",
		X"00",X"E5",X"5E",X"FF",X"00",X"FF",X"55",X"FE",X"00",X"EE",X"EE",X"EE",X"00",X"00",X"1F",X"55",
		X"00",X"0E",X"EE",X"55",X"00",X"0E",X"00",X"55",X"00",X"EF",X"00",X"5E",X"00",X"EF",X"00",X"5E",
		X"00",X"FF",X"00",X"5E",X"00",X"EE",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"EF",X"00",X"00",X"00",X"EF",X"00",X"00",X"EE",X"FF",X"00",
		X"00",X"5E",X"FF",X"00",X"00",X"5F",X"FF",X"00",X"00",X"6E",X"FF",X"00",X"00",X"F6",X"EF",X"00",
		X"00",X"EE",X"EE",X"00",X"00",X"EE",X"E5",X"EE",X"00",X"F0",X"1E",X"5F",X"00",X"E0",X"F1",X"FF",
		X"00",X"00",X"EE",X"5F",X"00",X"00",X"FE",X"55",X"00",X"00",X"FE",X"55",X"00",X"00",X"E0",X"55",
		X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"0E",X"00",X"00",X"0E",X"EF",X"00",X"00",X"0E",X"EF",X"00",X"00",X"EF",X"FF",X"00",
		X"00",X"E5",X"FF",X"00",X"00",X"E5",X"FF",X"00",X"00",X"E5",X"FF",X"EE",X"00",X"65",X"55",X"FF",
		X"00",X"EF",X"55",X"FF",X"00",X"EE",X"55",X"FF",X"00",X"00",X"EE",X"FF",X"00",X"00",X"16",X"FF",
		X"00",X"00",X"EE",X"EE",X"00",X"00",X"E0",X"55",X"00",X"0E",X"00",X"55",X"00",X"0E",X"00",X"55",
		X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"EE",X"EF",X"00",X"00",X"55",X"FF",X"00",
		X"00",X"55",X"FF",X"00",X"00",X"5E",X"FF",X"00",X"00",X"6F",X"FF",X"00",X"00",X"FE",X"E5",X"E0",
		X"00",X"E0",X"55",X"FE",X"00",X"00",X"E5",X"FE",X"00",X"00",X"1E",X"FE",X"00",X"00",X"F1",X"E0",
		X"00",X"00",X"EE",X"E0",X"00",X"0E",X"00",X"5E",X"00",X"EF",X"00",X"5E",X"00",X"EF",X"00",X"5E",
		X"00",X"0E",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"0E",X"00",X"00",X"EE",X"EF",X"00",X"00",X"55",X"FF",X"00",
		X"00",X"5F",X"FF",X"00",X"00",X"6E",X"FF",X"00",X"00",X"6E",X"FF",X"00",X"00",X"EE",X"FF",X"EE",
		X"00",X"E0",X"EF",X"FE",X"00",X"00",X"5E",X"FE",X"00",X"00",X"E5",X"FE",X"00",X"00",X"FE",X"FE",
		X"00",X"00",X"EE",X"E5",X"00",X"00",X"FE",X"55",X"00",X"00",X"E0",X"55",X"00",X"00",X"00",X"55",
		X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"E5",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"E5",X"EE",X"00",X"00",X"F5",X"EF",X"00",
		X"00",X"E6",X"FF",X"00",X"00",X"0E",X"FF",X"00",X"00",X"0E",X"FF",X"00",X"00",X"0F",X"FF",X"00",
		X"00",X"EE",X"EF",X"EE",X"00",X"F0",X"55",X"EF",X"00",X"00",X"EE",X"FF",X"00",X"00",X"F1",X"FF",
		X"00",X"00",X"EE",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FE",X"EE",X"00",X"00",X"E0",X"55",
		X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"5E",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"0E",X"00",X"00",X"F5",X"EF",X"00",
		X"00",X"FE",X"FF",X"00",X"00",X"EF",X"FF",X"00",X"00",X"FE",X"FF",X"00",X"00",X"0E",X"FF",X"00",
		X"00",X"00",X"EF",X"00",X"00",X"00",X"55",X"EE",X"00",X"00",X"E5",X"FE",X"00",X"00",X"1E",X"FE",
		X"00",X"00",X"E1",X"FE",X"00",X"00",X"FE",X"EE",X"00",X"00",X"E0",X"5E",X"00",X"00",X"00",X"5E",
		X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"F5",X"E0",X"00",X"00",X"EF",X"5E",X"00",X"00",X"EE",X"5E",X"00",
		X"00",X"0E",X"EF",X"00",X"00",X"F0",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"EF",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"1E",X"E0",
		X"00",X"00",X"EE",X"FE",X"00",X"00",X"EE",X"FE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",
		X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"0E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"F5",X"E0",X"00",X"00",X"EF",X"EE",X"00",X"00",X"EE",X"5E",X"00",X"00",X"0F",X"5E",X"00",
		X"00",X"E0",X"EE",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"5F",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"E5",X"00",X"00",X"0E",X"E5",X"00",
		X"00",X"0E",X"15",X"00",X"00",X"0E",X"65",X"E0",X"00",X"0E",X"EF",X"E0",X"00",X"00",X"0E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"0E",X"E0",X"00",X"00",X"0E",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"E0",X"00",X"00",X"E5",X"00",X"00",X"00",X"EF",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"0E",X"E0",X"00",X"00",X"00",X"5E",X"00",X"00",X"0F",X"5E",X"00",
		X"00",X"EE",X"5E",X"00",X"00",X"F0",X"EF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"EF",X"00",X"00",X"00",X"5F",X"00",X"00",X"0E",X"5E",X"00",X"00",X"0E",X"E5",X"00",
		X"00",X"0E",X"E5",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"E6",X"E0",X"00",X"00",X"0E",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"5E",X"00",X"00",X"0E",X"55",X"00",X"00",X"FE",X"55",X"E0",
		X"00",X"00",X"5E",X"E0",X"00",X"00",X"5F",X"E0",X"00",X"00",X"5F",X"00",X"00",X"00",X"5F",X"00",
		X"00",X"00",X"5F",X"00",X"00",X"00",X"55",X"00",X"00",X"0E",X"E5",X"00",X"00",X"0E",X"E5",X"00",
		X"00",X"0E",X"E5",X"00",X"00",X"0E",X"65",X"00",X"00",X"00",X"E6",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"E5",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"FE",X"00",X"00",X"0E",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"0E",X"5E",X"00",X"00",X"EF",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"5E",X"00",X"00",X"00",X"EF",X"E0",X"00",X"00",X"FF",X"E0",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"EF",X"00",X"00",X"0E",X"5E",X"00",X"00",X"EE",X"55",X"00",
		X"00",X"0E",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"E5",X"00",
		X"00",X"00",X"E5",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"0E",X"5E",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"E5",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"EF",X"E0",X"00",X"00",X"FF",X"E0",
		X"00",X"0E",X"FF",X"E0",X"00",X"EE",X"5F",X"E0",X"00",X"EF",X"5E",X"00",X"00",X"EF",X"55",X"00",
		X"00",X"EE",X"5E",X"00",X"00",X"0E",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"5E",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"0E",X"5E",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"E0",
		X"00",X"0E",X"FF",X"E0",X"00",X"EF",X"EF",X"E0",X"00",X"EF",X"EF",X"00",X"00",X"0F",X"EF",X"00",
		X"00",X"00",X"5E",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"5E",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"5F",X"00",X"00",X"00",X"EF",X"00",
		X"00",X"00",X"5E",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"5E",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"2E",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"5E",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"EF",X"00",X"00",X"00",X"EF",X"00",
		X"00",X"00",X"EF",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",
		X"EE",X"00",X"E0",X"00",X"E9",X"00",X"E0",X"00",X"E9",X"00",X"E0",X"00",X"E9",X"00",X"1E",X"00",
		X"E9",X"00",X"99",X"E0",X"99",X"00",X"99",X"EE",X"99",X"EE",X"EE",X"3E",X"99",X"BE",X"EB",X"9E",
		X"99",X"BB",X"BB",X"E2",X"9E",X"BB",X"BB",X"2E",X"EE",X"BB",X"EB",X"EE",X"0E",X"BB",X"EB",X"EB",
		X"0E",X"BB",X"EB",X"E9",X"0E",X"EE",X"EE",X"E9",X"0E",X"00",X"19",X"EE",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",
		X"EE",X"00",X"E0",X"00",X"E9",X"00",X"E0",X"00",X"E9",X"00",X"E0",X"00",X"E9",X"00",X"1E",X"00",
		X"E9",X"00",X"99",X"E0",X"9E",X"00",X"BB",X"EF",X"9E",X"EE",X"EE",X"FF",X"9E",X"AA",X"EA",X"EE",
		X"9E",X"AA",X"BE",X"BB",X"9E",X"EE",X"EE",X"BB",X"EE",X"BB",X"BB",X"BB",X"0E",X"BB",X"BB",X"BB",
		X"0E",X"EE",X"BB",X"BB",X"0E",X"F3",X"EE",X"BB",X"0E",X"3F",X"99",X"BB",X"0E",X"EE",X"B9",X"EE",
		X"0E",X"00",X"BB",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"3E",X"00",X"00",X"00",X"F1",X"00",
		X"00",X"00",X"F3",X"00",X"00",X"00",X"F3",X"00",X"00",X"00",X"1E",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"E0",X"00",
		X"EE",X"0E",X"E0",X"00",X"E9",X"EE",X"E0",X"00",X"E9",X"3E",X"FE",X"00",X"E9",X"EE",X"EE",X"00",
		X"E9",X"E1",X"EE",X"E0",X"99",X"11",X"E1",X"EE",X"99",X"E1",X"11",X"3E",X"99",X"EE",X"33",X"EE",
		X"99",X"EE",X"31",X"E2",X"9E",X"EE",X"11",X"2E",X"EE",X"EE",X"1E",X"EE",X"0E",X"11",X"1E",X"E2",
		X"0E",X"11",X"1E",X"E2",X"0E",X"13",X"11",X"E2",X"0E",X"11",X"11",X"EE",X"00",X"11",X"31",X"00",
		X"00",X"1E",X"EE",X"00",X"00",X"1E",X"EE",X"00",X"00",X"1E",X"EE",X"00",X"00",X"EE",X"E0",X"00",
		X"00",X"E0",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"F0",X"00",X"33",X"11",X"00",
		X"EE",X"3E",X"11",X"00",X"E9",X"E3",X"11",X"30",X"E9",X"31",X"FE",X"10",X"E9",X"E1",X"EE",X"00",
		X"E9",X"E1",X"EE",X"E0",X"99",X"EE",X"EE",X"EE",X"99",X"EE",X"EE",X"3E",X"99",X"EE",X"EE",X"EE",
		X"99",X"33",X"EE",X"E2",X"9E",X"11",X"EE",X"2E",X"EE",X"1E",X"EE",X"EE",X"0E",X"1E",X"EE",X"E2",
		X"0E",X"EE",X"EE",X"E2",X"0E",X"EE",X"EE",X"E2",X"0E",X"EE",X"EE",X"EE",X"00",X"EE",X"EE",X"00",
		X"00",X"EE",X"EE",X"33",X"00",X"EE",X"EE",X"11",X"00",X"EE",X"1E",X"10",X"00",X"EE",X"11",X"00",
		X"00",X"E3",X"E1",X"00",X"00",X"01",X"E1",X"00",X"00",X"11",X"E0",X"00",X"00",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"AA",X"AE",X"00",X"00",X"EA",X"AE",X"00",X"00",X"EA",X"AA",X"00",X"00",X"EA",X"AA",X"00",
		X"00",X"AE",X"AA",X"00",X"00",X"AA",X"1A",X"EE",X"00",X"2E",X"1A",X"EE",X"00",X"2E",X"EE",X"AE",
		X"00",X"BE",X"EE",X"BB",X"00",X"EE",X"32",X"1B",X"00",X"EE",X"AA",X"EE",X"00",X"EE",X"AA",X"EB",
		X"00",X"01",X"AA",X"BE",X"00",X"EE",X"EA",X"B9",X"00",X"EB",X"EA",X"B9",X"00",X"BB",X"9E",X"99",
		X"00",X"BB",X"EE",X"EE",X"00",X"B2",X"EA",X"00",X"00",X"B9",X"EA",X"00",X"00",X"99",X"EA",X"00",
		X"00",X"9E",X"EA",X"00",X"00",X"E0",X"EA",X"00",X"00",X"00",X"EA",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"00",X"3A",X"00",X"00",X"00",X"EA",X"00",X"00",X"00",X"EA",X"00",X"00",X"00",X"AA",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"EA",X"00",X"00",X"AE",X"AA",X"00",X"00",X"E0",X"EE",X"00",X"00",X"0E",X"2E",X"00",
		X"00",X"EE",X"2A",X"00",X"00",X"AE",X"EA",X"00",X"00",X"AE",X"EE",X"00",X"00",X"AA",X"AE",X"00",
		X"00",X"E2",X"AA",X"00",X"00",X"E2",X"EE",X"00",X"00",X"EA",X"EE",X"00",X"00",X"AA",X"AE",X"00",
		X"00",X"AA",X"EA",X"00",X"00",X"EE",X"AE",X"00",X"00",X"2E",X"EE",X"00",X"00",X"12",X"EE",X"00",
		X"00",X"EE",X"12",X"00",X"00",X"EE",X"EE",X"00",X"00",X"AE",X"1E",X"00",X"00",X"AE",X"2E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"0E",X"00",X"00",X"0A",X"EE",X"00",X"00",X"0E",X"EE",X"00",X"00",
		X"00",X"EF",X"EE",X"E0",X"00",X"BF",X"EE",X"EE",X"00",X"BE",X"EE",X"EE",X"0E",X"EE",X"EA",X"EE",
		X"00",X"AE",X"EE",X"E5",X"00",X"AA",X"EE",X"7E",X"00",X"EE",X"1E",X"BE",X"00",X"BB",X"EE",X"EE",
		X"00",X"BB",X"EE",X"E9",X"00",X"BB",X"99",X"99",X"00",X"EB",X"BB",X"BB",X"00",X"E2",X"92",X"22",
		X"00",X"02",X"20",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"E0",X"00",X"0F",X"01",X"E0",X"00",
		X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"E0",X"10",X"E0",X"00",X"00",X"10",X"00",
		X"00",X"10",X"11",X"11",X"00",X"00",X"10",X"00",X"0F",X"E0",X"10",X"E0",X"0F",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"0F",X"01",X"E0",X"00",X"0F",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"0E",X"EE",X"00",X"11",X"EE",X"99",X"00",X"01",X"99",X"AA",X"00",X"00",X"99",X"AA",
		X"00",X"F0",X"92",X"EE",X"00",X"EE",X"22",X"00",X"00",X"1E",X"EE",X"E3",X"00",X"11",X"EE",X"EE",
		X"00",X"E1",X"1E",X"E3",X"00",X"EE",X"1E",X"EE",X"00",X"EE",X"3F",X"EE",X"00",X"EE",X"EE",X"EE",
		X"00",X"EE",X"3E",X"EE",X"00",X"FF",X"3F",X"FE",X"00",X"EF",X"3F",X"EE",X"00",X"EE",X"FF",X"EF",
		X"00",X"EE",X"11",X"EF",X"00",X"0E",X"EE",X"EE",X"00",X"EF",X"FE",X"FE",X"00",X"EE",X"11",X"EE",
		X"00",X"13",X"11",X"E3",X"00",X"11",X"EE",X"EE",X"00",X"11",X"EE",X"03",X"00",X"EE",X"22",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"2E",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"EF",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"21",X"00",X"10",X"00",X"92",X"EE",X"10",X"00",X"AA",X"99",X"11",X"00",X"A1",X"99",X"11",
		X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"E1",X"00",X"11",X"11",X"EE",X"01",X"1E",X"1E",X"EE",
		X"01",X"EE",X"EE",X"E0",X"01",X"1E",X"EE",X"30",X"01",X"1E",X"EE",X"30",X"00",X"11",X"EE",X"30",
		X"00",X"11",X"EE",X"E3",X"00",X"EE",X"EE",X"E3",X"0E",X"EE",X"EE",X"33",X"0E",X"EE",X"EE",X"33",
		X"0E",X"EE",X"EE",X"EE",X"00",X"1E",X"EE",X"EE",X"00",X"EE",X"EE",X"EE",X"00",X"11",X"EE",X"3E",
		X"00",X"11",X"EE",X"31",X"00",X"33",X"E1",X"3E",X"00",X"13",X"E1",X"1E",X"00",X"33",X"11",X"13",
		X"00",X"31",X"11",X"1E",X"00",X"01",X"11",X"EE",X"00",X"11",X"13",X"E1",X"00",X"11",X"13",X"13",
		X"00",X"11",X"10",X"11",X"00",X"EE",X"11",X"00",X"00",X"EE",X"11",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"60",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"62",X"F0",X"00",X"06",X"00",X"00",
		X"00",X"26",X"20",X"02",X"00",X"02",X"06",X"00",X"00",X"66",X"66",X"00",X"00",X"0F",X"66",X"06",
		X"0F",X"02",X"F6",X"F0",X"00",X"22",X"F6",X"20",X"00",X"20",X"62",X"00",X"00",X"20",X"62",X"00",
		X"00",X"22",X"22",X"00",X"00",X"02",X"2F",X"02",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",
		X"0F",X"F2",X"02",X"20",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"20",X"22",X"00",
		X"00",X"20",X"22",X"00",X"00",X"20",X"22",X"00",X"00",X"20",X"22",X"00",X"00",X"20",X"22",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",
		X"00",X"02",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",
		X"00",X"20",X"06",X"00",X"00",X"22",X"06",X"00",X"00",X"02",X"26",X"06",X"00",X"00",X"26",X"60",
		X"00",X"00",X"2F",X"60",X"00",X"20",X"22",X"00",X"00",X"22",X"22",X"60",X"00",X"00",X"22",X"26",
		X"00",X"02",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"27",X"00",X"00",X"00",X"27",X"00",
		X"00",X"00",X"27",X"00",X"00",X"00",X"27",X"00",X"00",X"00",X"27",X"00",X"00",X"00",X"27",X"00",
		X"00",X"00",X"27",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E8",
		X"00",X"00",X"00",X"86",X"00",X"00",X"00",X"6C",X"00",X"00",X"00",X"42",X"00",X"00",X"00",X"4C",
		X"00",X"00",X"00",X"E2",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"7F",X"00",X"00",X"00",X"7F",X"70",
		X"00",X"70",X"00",X"0F",X"00",X"EF",X"00",X"07",X"00",X"70",X"70",X"00",X"F0",X"FF",X"FF",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"66",X"EE",X"00",X"00",X"66",X"E5",X"00",X"00",X"E6",X"FE",X"00",
		X"00",X"E6",X"FF",X"00",X"00",X"EA",X"FF",X"00",X"00",X"EA",X"FF",X"0E",X"00",X"EF",X"EE",X"EF",
		X"00",X"EE",X"EF",X"FF",X"00",X"66",X"66",X"66",X"00",X"AA",X"EE",X"E2",X"00",X"FF",X"FF",X"EE",
		X"00",X"FF",X"EE",X"BB",X"00",X"FF",X"EE",X"BB",X"00",X"FF",X"EE",X"EE",X"00",X"EE",X"EE",X"00",
		X"0E",X"AA",X"00",X"00",X"0E",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"E1",X"00",X"00",
		X"00",X"11",X"E0",X"00",X"00",X"EE",X"9E",X"00",X"00",X"0E",X"D9",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"DE",X"00",X"00",X"00",X"EF",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"BB",X"E0",X"00",X"00",X"BB",X"EE",
		X"00",X"00",X"BB",X"BE",X"00",X"00",X"EB",X"BB",X"00",X"00",X"EB",X"BB",X"00",X"00",X"EB",X"BB",
		X"00",X"00",X"EB",X"BB",X"00",X"00",X"EB",X"EE",X"00",X"00",X"EE",X"F7",X"0F",X"7F",X"F7",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"0E",X"EE",
		X"00",X"00",X"EB",X"AA",X"0E",X"00",X"BE",X"AA",X"EB",X"00",X"BE",X"EE",X"BB",X"00",X"BB",X"CC",
		X"EE",X"00",X"EB",X"EF",X"77",X"F7",X"EB",X"EF",X"77",X"10",X"71",X"E7",X"00",X"70",X"00",X"00",
		X"00",X"01",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"FC",
		X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"EE",X"00",X"00",X"07",X"EE",X"9A",X"E0",X"00",X"EE",
		X"BB",X"E7",X"7E",X"BB",X"77",X"E7",X"EE",X"E7",X"77",X"00",X"7E",X"E7",X"00",X"70",X"00",X"06",
		X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"E0",X"00",
		X"0E",X"00",X"2E",X"00",X"0E",X"00",X"21",X"00",X"0E",X"00",X"EE",X"EE",X"0E",X"EE",X"E2",X"2E",
		X"0E",X"22",X"22",X"E1",X"00",X"22",X"22",X"FE",X"E0",X"22",X"E2",X"EE",X"00",X"22",X"E2",X"22",
		X"00",X"EE",X"EE",X"22",X"00",X"00",X"EE",X"EE",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",
		X"00",X"00",X"22",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"E0",X"00",
		X"E0",X"0E",X"E0",X"00",X"00",X"EE",X"E0",X"00",X"0E",X"2E",X"5E",X"00",X"0E",X"EE",X"EE",X"00",
		X"0E",X"E7",X"2E",X"E0",X"0E",X"77",X"22",X"EE",X"0E",X"E7",X"22",X"6E",X"00",X"26",X"22",X"EE",
		X"00",X"26",X"22",X"E2",X"00",X"26",X"22",X"2E",X"00",X"26",X"E2",X"EE",X"00",X"66",X"E2",X"E2",
		X"0E",X"62",X"22",X"E2",X"0E",X"22",X"26",X"E2",X"0E",X"22",X"77",X"EE",X"0E",X"22",X"26",X"00",
		X"0E",X"6E",X"66",X"00",X"00",X"6E",X"EE",X"00",X"00",X"6E",X"EE",X"00",X"00",X"EE",X"E0",X"00",
		X"00",X"E0",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"05",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"0E",X"DD",X"EE",X"00",X"EE",X"DD",X"DD",X"00",X"EE",X"DD",X"DD",X"00",X"EE",X"EE",X"DD",
		X"00",X"CC",X"CC",X"EE",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CE",X"BC",X"00",X"BB",X"E2",X"EC",
		X"00",X"EE",X"EF",X"0E",X"00",X"00",X"0E",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"ED",X"00",X"00",X"F0",X"DD",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"0E",X"DD",X"00",X"00",X"EE",X"DD",X"00",X"00",X"EE",X"DD",X"EE",X"00",X"EC",X"CC",X"DD",
		X"00",X"EC",X"CE",X"DD",X"00",X"BB",X"CC",X"DE",X"00",X"EE",X"EE",X"DE",X"00",X"00",X"1B",X"CC",
		X"00",X"0E",X"EE",X"CC",X"00",X"0E",X"00",X"CC",X"00",X"ED",X"00",X"CE",X"00",X"ED",X"00",X"CE",
		X"00",X"DD",X"00",X"CE",X"00",X"EE",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"ED",X"00",X"00",X"00",X"ED",X"00",X"00",X"EE",X"DD",X"00",
		X"00",X"CE",X"DD",X"00",X"00",X"CF",X"DD",X"00",X"00",X"CC",X"DD",X"00",X"00",X"B6",X"ED",X"00",
		X"00",X"EE",X"EE",X"00",X"00",X"EE",X"EC",X"EE",X"00",X"F0",X"2E",X"CD",X"00",X"E0",X"F2",X"DD",
		X"00",X"00",X"EE",X"CD",X"00",X"00",X"DE",X"CC",X"00",X"00",X"DE",X"CC",X"00",X"00",X"E0",X"CC",
		X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"0E",X"00",X"00",X"0E",X"ED",X"00",X"00",X"0E",X"ED",X"00",X"00",X"EF",X"DD",X"00",
		X"00",X"EC",X"DD",X"00",X"00",X"EC",X"DD",X"00",X"00",X"EC",X"DD",X"EE",X"00",X"FC",X"CC",X"DD",
		X"00",X"EB",X"CC",X"DD",X"00",X"EE",X"CC",X"DD",X"00",X"00",X"EE",X"DD",X"00",X"00",X"2F",X"DD",
		X"00",X"00",X"EE",X"EE",X"00",X"00",X"E0",X"CC",X"00",X"0E",X"00",X"CC",X"00",X"0E",X"00",X"CC",
		X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"EE",X"ED",X"00",X"00",X"CC",X"DD",X"00",
		X"00",X"CC",X"DD",X"00",X"00",X"CE",X"DD",X"00",X"00",X"BB",X"DD",X"00",X"00",X"FE",X"EC",X"E0",
		X"00",X"E0",X"CC",X"DE",X"00",X"00",X"EC",X"DE",X"00",X"00",X"2E",X"DE",X"00",X"00",X"B2",X"E0",
		X"00",X"00",X"EE",X"E0",X"00",X"0E",X"00",X"CE",X"00",X"ED",X"00",X"CE",X"00",X"ED",X"00",X"CE",
		X"00",X"0E",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"0E",X"00",X"00",X"EE",X"ED",X"00",X"00",X"CC",X"DD",X"00",
		X"00",X"CF",X"DD",X"00",X"00",X"BE",X"DD",X"00",X"00",X"BE",X"DD",X"00",X"00",X"EE",X"DD",X"EE",
		X"00",X"E0",X"EE",X"DE",X"00",X"00",X"CE",X"DE",X"00",X"00",X"EC",X"DE",X"00",X"00",X"FE",X"DE",
		X"00",X"00",X"EE",X"EC",X"00",X"00",X"DE",X"CC",X"00",X"00",X"E0",X"CC",X"00",X"00",X"00",X"CC",
		X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"EC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"EC",X"EE",X"00",X"00",X"BC",X"ED",X"00",
		X"00",X"EB",X"DD",X"00",X"00",X"0E",X"DD",X"00",X"00",X"0E",X"DD",X"00",X"00",X"0F",X"DD",X"00",
		X"00",X"EE",X"CE",X"EE",X"00",X"F0",X"CC",X"ED",X"00",X"00",X"EE",X"DD",X"00",X"00",X"B2",X"DD",
		X"00",X"00",X"EE",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DE",X"EE",X"00",X"00",X"E0",X"CC",
		X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"CE",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"0E",X"00",X"00",X"BC",X"ED",X"00",
		X"00",X"FE",X"DD",X"00",X"00",X"EB",X"DD",X"00",X"00",X"FE",X"DD",X"00",X"00",X"0E",X"DD",X"00",
		X"00",X"00",X"DD",X"00",X"00",X"00",X"CC",X"EE",X"00",X"00",X"EC",X"DE",X"00",X"00",X"2E",X"DE",
		X"00",X"00",X"E2",X"DE",X"00",X"00",X"DE",X"EE",X"00",X"00",X"E0",X"CE",X"00",X"00",X"00",X"CE",
		X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"BC",X"E0",X"00",X"00",X"EB",X"CE",X"00",X"00",X"EE",X"CE",X"00",
		X"00",X"0E",X"ED",X"00",X"00",X"F0",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"DD",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"2E",X"E0",
		X"00",X"00",X"EE",X"DE",X"00",X"00",X"EE",X"DE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",
		X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"0E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"BC",X"E0",X"00",X"00",X"EB",X"EE",X"00",X"00",X"EE",X"CE",X"00",X"00",X"0F",X"CE",X"00",
		X"00",X"E0",X"EE",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"CD",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"EC",X"00",X"00",X"0E",X"EC",X"00",
		X"00",X"0E",X"2C",X"00",X"00",X"0E",X"BC",X"E0",X"00",X"0E",X"EB",X"E0",X"00",X"00",X"0E",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"0E",X"E0",X"00",X"00",X"0E",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"E0",X"00",X"00",X"EC",X"00",X"00",X"00",X"EB",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"0E",X"E0",X"00",X"00",X"00",X"CE",X"00",X"00",X"0F",X"CE",X"00",
		X"00",X"EE",X"CE",X"00",X"00",X"F0",X"ED",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"DD",X"00",X"00",X"00",X"CD",X"00",X"00",X"0E",X"CE",X"00",X"00",X"0E",X"EC",X"00",
		X"00",X"0E",X"EC",X"00",X"00",X"00",X"BC",X"00",X"00",X"00",X"EB",X"E0",X"00",X"00",X"0E",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"CE",X"00",X"00",X"0E",X"CC",X"00",X"00",X"FE",X"CC",X"E0",
		X"00",X"00",X"CE",X"E0",X"00",X"00",X"CD",X"E0",X"00",X"00",X"CD",X"00",X"00",X"00",X"CD",X"00",
		X"00",X"00",X"CD",X"00",X"00",X"00",X"CC",X"00",X"00",X"0E",X"EC",X"00",X"00",X"0E",X"EC",X"00",
		X"00",X"0E",X"EC",X"00",X"00",X"0E",X"BC",X"00",X"00",X"00",X"EB",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"EC",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"FE",X"00",X"00",X"0E",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"0E",X"CE",X"00",X"00",X"EF",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CE",X"00",X"00",X"00",X"ED",X"E0",X"00",X"00",X"DD",X"E0",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"DD",X"00",X"00",X"00",X"ED",X"00",X"00",X"0E",X"CE",X"00",X"00",X"EE",X"CC",X"00",
		X"00",X"0E",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"EC",X"00",
		X"00",X"00",X"EC",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"0E",X"CE",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"EC",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"ED",X"E0",X"00",X"00",X"DD",X"E0",
		X"00",X"0E",X"DD",X"E0",X"00",X"EE",X"CD",X"E0",X"00",X"ED",X"CE",X"00",X"00",X"ED",X"CC",X"00",
		X"00",X"EE",X"CE",X"00",X"00",X"0E",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CE",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"0E",X"CE",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"E0",
		X"00",X"0E",X"DD",X"E0",X"00",X"ED",X"ED",X"E0",X"00",X"ED",X"ED",X"00",X"00",X"0D",X"ED",X"00",
		X"00",X"00",X"CE",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CE",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CD",X"00",X"00",X"00",X"ED",X"00",
		X"00",X"00",X"CE",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"CE",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"2E",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"CE",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CE",X"00",X"00",X"00",X"ED",X"00",X"00",X"00",X"ED",X"00",X"00",X"00",X"ED",X"00",
		X"00",X"00",X"CE",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",X"EE",
		X"00",X"00",X"EE",X"3E",X"00",X"00",X"2E",X"E0",X"00",X"E0",X"22",X"EE",X"00",X"3E",X"22",X"2E",
		X"00",X"E3",X"22",X"2E",X"00",X"EE",X"22",X"E3",X"00",X"E2",X"22",X"3E",X"00",X"22",X"22",X"EE",
		X"00",X"22",X"32",X"EE",X"00",X"22",X"32",X"22",X"00",X"22",X"E2",X"22",X"00",X"3E",X"22",X"22",
		X"00",X"E2",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",
		X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"E2",X"22",X"22",X"00",X"E2",X"22",X"22",
		X"00",X"EE",X"22",X"22",X"00",X"E3",X"22",X"22",X"00",X"3E",X"22",X"2E",X"00",X"07",X"77",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"E0",X"00",X"00",X"F5",X"FE",
		X"00",X"00",X"55",X"5F",X"00",X"00",X"55",X"55",X"00",X"00",X"5E",X"55",X"00",X"00",X"EF",X"E5",
		X"00",X"06",X"EF",X"EF",X"00",X"00",X"EE",X"EF",X"00",X"00",X"00",X"FF",X"00",X"60",X"00",X"FF",
		X"00",X"00",X"00",X"F5",X"00",X"EE",X"00",X"55",X"00",X"EE",X"00",X"55",X"00",X"EE",X"00",X"55",
		X"00",X"EE",X"06",X"E5",X"00",X"EE",X"00",X"E5",X"00",X"5E",X"00",X"E5",X"00",X"55",X"00",X"EE",
		X"AE",X"55",X"E6",X"E0",X"AE",X"55",X"00",X"00",X"0D",X"55",X"00",X"00",X"0E",X"EE",X"00",X"00",
		X"00",X"5E",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"E0",X"00",X"00",X"FC",X"FE",
		X"00",X"00",X"CC",X"CF",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CE",X"CC",X"00",X"00",X"EF",X"EC",
		X"00",X"06",X"EF",X"EF",X"00",X"00",X"EE",X"EF",X"00",X"00",X"00",X"FF",X"00",X"60",X"00",X"FF",
		X"00",X"00",X"00",X"FC",X"00",X"EE",X"00",X"CC",X"00",X"EE",X"00",X"CC",X"00",X"EE",X"00",X"CC",
		X"00",X"EE",X"06",X"EC",X"00",X"EE",X"00",X"EC",X"00",X"BE",X"00",X"EC",X"00",X"CB",X"00",X"EE",
		X"AE",X"CB",X"E6",X"E0",X"AE",X"CC",X"00",X"00",X"0D",X"CC",X"00",X"00",X"0E",X"EE",X"00",X"00",
		X"00",X"BE",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"00",
		X"00",X"55",X"55",X"00",X"0E",X"55",X"5E",X"00",X"0E",X"BB",X"BB",X"E0",X"0E",X"BB",X"BB",X"E0",
		X"0E",X"BB",X"BB",X"E0",X"E9",X"BB",X"BB",X"E0",X"E9",X"BB",X"BB",X"E0",X"E9",X"BB",X"BB",X"E0",
		X"E9",X"BB",X"BB",X"EE",X"7B",X"BB",X"BB",X"BE",X"E7",X"BB",X"BB",X"BE",X"00",X"BB",X"7B",X"7E",
		X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"0F",X"00",X"00",X"00",X"30",X"0F",X"00",X"30",X"00",X"30",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",X"03",X"00",X"00",X"F0",X"F0",X"F0",
		X"00",X"01",X"20",X"00",X"00",X"11",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"0E",X"E0",X"00",X"00",X"0E",X"E0",X"00",X"00",X"E6",X"20",X"00",
		X"00",X"E6",X"00",X"00",X"00",X"E6",X"00",X"00",X"00",X"EE",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"10",X"E1",X"00",X"00",X"1E",X"66",X"00",X"00",X"E6",X"E6",X"00",X"00",X"66",X"E6",X"00",
		X"00",X"16",X"66",X"00",X"00",X"66",X"E6",X"00",X"00",X"66",X"BE",X"00",X"00",X"66",X"BE",X"00",
		X"00",X"EE",X"BE",X"00",X"00",X"00",X"BE",X"00",X"00",X"00",X"5B",X"00",X"00",X"00",X"5B",X"00",
		X"00",X"00",X"5B",X"00",X"00",X"00",X"5B",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"5E",X"00",
		X"00",X"01",X"20",X"00",X"00",X"11",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"0E",X"E0",X"00",X"00",X"0E",X"E0",X"00",X"00",X"ED",X"20",X"00",
		X"00",X"ED",X"00",X"00",X"00",X"ED",X"00",X"00",X"00",X"EE",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"E1",X"00",X"00",X"0E",X"DD",X"00",X"00",X"ED",X"ED",X"00",X"00",X"DD",X"ED",X"00",
		X"00",X"3D",X"DD",X"00",X"00",X"DD",X"ED",X"00",X"00",X"DD",X"BE",X"00",X"00",X"DD",X"BE",X"00",
		X"00",X"EE",X"BE",X"00",X"00",X"00",X"BE",X"00",X"00",X"00",X"CB",X"00",X"00",X"00",X"CB",X"00",
		X"00",X"00",X"CB",X"00",X"00",X"00",X"CB",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"CE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
