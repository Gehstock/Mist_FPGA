library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity bg is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(18 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of bg is
	type rom is array(0 to  262623) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FE",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"02",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FE",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"01",X"00",X"FF",X"FF",X"01",X"00",X"FE",X"FF",X"02",X"00",X"FF",X"FF",X"01",X"00",X"FE",X"FF",
		X"03",X"00",X"F9",X"FF",X"34",X"00",X"25",X"01",X"DD",X"01",X"55",X"02",X"A3",X"02",X"D6",X"02",
		X"F1",X"02",X"FD",X"02",X"FE",X"02",X"F6",X"02",X"E6",X"02",X"D5",X"02",X"BE",X"02",X"A3",X"02",
		X"89",X"02",X"69",X"02",X"4A",X"02",X"2B",X"02",X"09",X"02",X"E5",X"01",X"C3",X"01",X"9E",X"01",
		X"7A",X"01",X"53",X"01",X"30",X"01",X"09",X"01",X"E5",X"00",X"BB",X"00",X"A6",X"00",X"DC",X"00",
		X"50",X"01",X"EA",X"01",X"9E",X"02",X"5D",X"03",X"27",X"04",X"F3",X"04",X"BF",X"05",X"88",X"06",
		X"4E",X"07",X"0D",X"08",X"CB",X"08",X"81",X"09",X"33",X"0A",X"E0",X"0A",X"87",X"0B",X"29",X"0C",
		X"C6",X"0C",X"5A",X"0D",X"EE",X"0D",X"7C",X"0E",X"02",X"0F",X"86",X"0F",X"04",X"10",X"7F",X"10",
		X"F5",X"10",X"69",X"11",X"AC",X"11",X"9A",X"11",X"54",X"11",X"EB",X"10",X"6D",X"10",X"DD",X"0F",
		X"47",X"0F",X"AD",X"0E",X"0F",X"0E",X"74",X"0D",X"D9",X"0C",X"3E",X"0C",X"A9",X"0B",X"18",X"0B",
		X"88",X"0A",X"FD",X"09",X"74",X"09",X"F0",X"08",X"6E",X"08",X"F0",X"07",X"76",X"07",X"00",X"07",
		X"8C",X"06",X"1B",X"06",X"AC",X"05",X"44",X"05",X"DB",X"04",X"7F",X"04",X"6E",X"04",X"A5",X"04",
		X"04",X"05",X"81",X"05",X"0D",X"06",X"A7",X"06",X"44",X"07",X"E6",X"07",X"86",X"08",X"26",X"09",
		X"C2",X"09",X"5A",X"0A",X"F1",X"0A",X"82",X"0B",X"10",X"0C",X"9A",X"0C",X"20",X"0D",X"A2",X"0D",
		X"1E",X"0E",X"98",X"0E",X"0F",X"0F",X"81",X"0F",X"EE",X"0F",X"5A",X"10",X"C2",X"10",X"26",X"11",
		X"89",X"11",X"C5",X"11",X"AA",X"11",X"5D",X"11",X"E7",X"10",X"5C",X"10",X"C3",X"0F",X"1F",X"0F",
		X"7A",X"0E",X"D2",X"0D",X"29",X"0D",X"83",X"0C",X"E1",X"0B",X"41",X"0B",X"A4",X"0A",X"0D",X"0A",
		X"77",X"09",X"E8",X"08",X"5A",X"08",X"D2",X"07",X"4C",X"07",X"CC",X"06",X"4D",X"06",X"D5",X"05",
		X"5E",X"05",X"EB",X"04",X"7B",X"04",X"0F",X"04",X"A9",X"03",X"8A",X"03",X"B5",X"03",X"0C",X"04",
		X"81",X"04",X"09",X"05",X"9E",X"05",X"38",X"06",X"D7",X"06",X"75",X"07",X"11",X"08",X"AC",X"08",
		X"43",X"09",X"D6",X"09",X"67",X"0A",X"F3",X"0A",X"7B",X"0B",X"FE",X"0B",X"80",X"0C",X"FC",X"0C",
		X"75",X"0D",X"EA",X"0D",X"5B",X"0E",X"C9",X"0E",X"34",X"0F",X"9C",X"0F",X"FE",X"0F",X"62",X"10",
		X"A4",X"10",X"93",X"10",X"49",X"10",X"D9",X"0F",X"4F",X"0F",X"B5",X"0E",X"12",X"0E",X"6D",X"0D",
		X"C4",X"0C",X"1C",X"0C",X"77",X"0B",X"D2",X"0A",X"30",X"0A",X"94",X"09",X"FC",X"08",X"65",X"08",
		X"D5",X"07",X"48",X"07",X"BE",X"06",X"39",X"06",X"B8",X"05",X"3A",X"05",X"BF",X"04",X"48",X"04",
		X"D6",X"03",X"64",X"03",X"F9",X"02",X"90",X"02",X"65",X"02",X"88",X"02",X"DB",X"02",X"4F",X"03",
		X"D5",X"03",X"68",X"04",X"02",X"05",X"A1",X"05",X"3F",X"06",X"DB",X"06",X"75",X"07",X"0D",X"08",
		X"A3",X"08",X"35",X"09",X"C1",X"09",X"4A",X"0A",X"D0",X"0A",X"50",X"0B",X"CE",X"0B",X"46",X"0C",
		X"BE",X"0C",X"2F",X"0D",X"9F",X"0D",X"0A",X"0E",X"71",X"0E",X"D6",X"0E",X"39",X"0F",X"85",X"0F",
		X"7E",X"0F",X"3B",X"0F",X"CE",X"0E",X"47",X"0E",X"AF",X"0D",X"10",X"0D",X"69",X"0C",X"C1",X"0B",
		X"19",X"0B",X"73",X"0A",X"CF",X"09",X"2F",X"09",X"92",X"08",X"F8",X"07",X"63",X"07",X"D2",X"06",
		X"44",X"06",X"BB",X"05",X"37",X"05",X"B4",X"04",X"36",X"04",X"BC",X"03",X"45",X"03",X"D1",X"02",
		X"61",X"02",X"F5",X"01",X"8C",X"01",X"25",X"01",X"C1",X"00",X"61",X"00",X"03",X"00",X"AA",X"FF",
		X"51",X"FF",X"FB",X"FE",X"A9",X"FE",X"58",X"FE",X"09",X"FE",X"BF",X"FD",X"74",X"FD",X"2C",X"FD",
		X"E8",X"FC",X"A5",X"FC",X"63",X"FC",X"24",X"FC",X"E6",X"FB",X"AB",X"FB",X"71",X"FB",X"42",X"FB",
		X"42",X"FB",X"43",X"FB",X"46",X"FB",X"4A",X"FB",X"4D",X"FB",X"4D",X"FB",X"50",X"FB",X"50",X"FB",
		X"58",X"FB",X"50",X"FB",X"BE",X"FB",X"89",X"FC",X"4B",X"FD",X"1C",X"FE",X"E6",X"FE",X"B6",X"FF",
		X"7D",X"00",X"46",X"01",X"05",X"02",X"C3",X"02",X"7B",X"03",X"2F",X"04",X"DC",X"04",X"87",X"05",
		X"2A",X"06",X"CA",X"06",X"64",X"07",X"FB",X"07",X"8C",X"08",X"19",X"09",X"A3",X"09",X"27",X"0A",
		X"A7",X"0A",X"24",X"0B",X"9C",X"0B",X"11",X"0C",X"83",X"0C",X"F0",X"0C",X"5B",X"0D",X"C1",X"0D",
		X"25",X"0E",X"85",X"0E",X"E2",X"0E",X"3D",X"0F",X"94",X"0F",X"E8",X"0F",X"3A",X"10",X"8A",X"10",
		X"D5",X"10",X"21",X"11",X"68",X"11",X"AE",X"11",X"EF",X"11",X"30",X"12",X"6E",X"12",X"AB",X"12",
		X"E5",X"12",X"1B",X"13",X"54",X"13",X"86",X"13",X"BC",X"13",X"CD",X"13",X"89",X"13",X"11",X"13",
		X"75",X"12",X"C2",X"11",X"01",X"11",X"39",X"10",X"6E",X"0F",X"A3",X"0E",X"D8",X"0D",X"10",X"0D",
		X"4E",X"0C",X"8D",X"0B",X"D1",X"0A",X"1C",X"0A",X"6B",X"09",X"BD",X"08",X"17",X"08",X"72",X"07",
		X"D3",X"06",X"39",X"06",X"A4",X"05",X"12",X"05",X"85",X"04",X"FB",X"03",X"76",X"03",X"F4",X"02",
		X"77",X"02",X"FE",X"01",X"86",X"01",X"14",X"01",X"A4",X"00",X"39",X"00",X"CF",X"FF",X"6B",X"FF",
		X"08",X"FF",X"A8",X"FE",X"4B",X"FE",X"F0",X"FD",X"98",X"FD",X"44",X"FD",X"F1",X"FC",X"A2",X"FC",
		X"53",X"FC",X"09",X"FC",X"C1",X"FB",X"79",X"FB",X"35",X"FB",X"F2",X"FA",X"B1",X"FA",X"73",X"FA",
		X"36",X"FA",X"FD",X"F9",X"C1",X"F9",X"94",X"F9",X"90",X"F9",X"A3",X"F9",X"0E",X"FA",X"A3",X"FA",
		X"4E",X"FB",X"09",X"FC",X"CC",X"FC",X"91",X"FD",X"58",X"FE",X"1D",X"FF",X"E0",X"FF",X"9E",X"00",
		X"59",X"01",X"0E",X"02",X"BF",X"02",X"6B",X"03",X"13",X"04",X"B7",X"04",X"54",X"05",X"EF",X"05",
		X"82",X"06",X"14",X"07",X"A0",X"07",X"28",X"08",X"AC",X"08",X"2C",X"09",X"A7",X"09",X"1E",X"0A",
		X"91",X"0A",X"03",X"0B",X"71",X"0B",X"DB",X"0B",X"40",X"0C",X"A2",X"0C",X"03",X"0D",X"61",X"0D",
		X"BA",X"0D",X"12",X"0E",X"65",X"0E",X"B7",X"0E",X"06",X"0F",X"52",X"0F",X"9C",X"0F",X"E2",X"0F",
		X"28",X"10",X"6A",X"10",X"AA",X"10",X"E8",X"10",X"25",X"11",X"5F",X"11",X"97",X"11",X"CE",X"11",
		X"02",X"12",X"33",X"12",X"66",X"12",X"84",X"12",X"53",X"12",X"E5",X"11",X"4E",X"11",X"9E",X"10",
		X"DE",X"0F",X"17",X"0F",X"48",X"0E",X"7C",X"0D",X"B0",X"0C",X"E5",X"0B",X"1E",X"0B",X"5D",X"0A",
		X"9F",X"09",X"E8",X"08",X"33",X"08",X"84",X"07",X"DA",X"06",X"34",X"06",X"93",X"05",X"F8",X"04",
		X"5F",X"04",X"CC",X"03",X"3C",X"03",X"B2",X"02",X"2A",X"02",X"A8",X"01",X"29",X"01",X"AF",X"00",
		X"35",X"00",X"C3",X"FF",X"52",X"FF",X"E4",X"FE",X"7B",X"FE",X"13",X"FE",X"AF",X"FD",X"4E",X"FD",
		X"F0",X"FC",X"93",X"FC",X"3B",X"FC",X"E5",X"FB",X"93",X"FB",X"43",X"FB",X"F5",X"FA",X"A7",X"FA",
		X"5D",X"FA",X"17",X"FA",X"D2",X"F9",X"8E",X"F9",X"4D",X"F9",X"0E",X"F9",X"D2",X"F8",X"96",X"F8",
		X"5D",X"F8",X"25",X"F8",X"07",X"F8",X"1D",X"F8",X"7A",X"F8",X"09",X"F9",X"AE",X"F9",X"65",X"FA",
		X"27",X"FB",X"ED",X"FB",X"B4",X"FC",X"79",X"FD",X"3D",X"FE",X"FD",X"FE",X"B9",X"FF",X"70",X"00",
		X"23",X"01",X"D0",X"01",X"7B",X"02",X"1F",X"03",X"BE",X"03",X"58",X"04",X"EF",X"04",X"81",X"05",
		X"0F",X"06",X"98",X"06",X"1D",X"07",X"9E",X"07",X"1A",X"08",X"94",X"08",X"0B",X"09",X"7B",X"09",
		X"E9",X"09",X"53",X"0A",X"BC",X"0A",X"20",X"0B",X"81",X"0B",X"DF",X"0B",X"3A",X"0C",X"92",X"0C",
		X"E8",X"0C",X"3B",X"0D",X"8A",X"0D",X"D8",X"0D",X"23",X"0E",X"6B",X"0E",X"B1",X"0E",X"F4",X"0E",
		X"37",X"0F",X"76",X"0F",X"B4",X"0F",X"EE",X"0F",X"26",X"10",X"5D",X"10",X"91",X"10",X"C7",X"10",
		X"F7",X"10",X"22",X"11",X"08",X"11",X"A4",X"10",X"17",X"10",X"6E",X"0F",X"B1",X"0E",X"EB",X"0D",
		X"20",X"0D",X"53",X"0C",X"87",X"0B",X"BC",X"0A",X"F5",X"09",X"33",X"09",X"76",X"08",X"BC",X"07",
		X"07",X"07",X"58",X"06",X"AC",X"05",X"06",X"05",X"66",X"04",X"C7",X"03",X"2F",X"03",X"9C",X"02",
		X"0B",X"02",X"80",X"01",X"FA",X"00",X"74",X"00",X"F6",X"FF",X"7C",X"FF",X"02",X"FF",X"8E",X"FE",
		X"1E",X"FE",X"AF",X"FD",X"45",X"FD",X"DF",X"FC",X"7A",X"FC",X"19",X"FC",X"BB",X"FB",X"5F",X"FB",
		X"06",X"FB",X"B0",X"FA",X"5C",X"FA",X"0C",X"FA",X"BD",X"F9",X"71",X"F9",X"27",X"F9",X"E2",X"F8",
		X"9A",X"F8",X"58",X"F8",X"17",X"F8",X"D8",X"F7",X"9B",X"F7",X"5F",X"F7",X"29",X"F7",X"EE",X"F6",
		X"C6",X"F6",X"CE",X"F6",X"1B",X"F7",X"A1",X"F7",X"41",X"F8",X"F8",X"F8",X"B5",X"F9",X"7C",X"FA",
		X"43",X"FB",X"0A",X"FC",X"CE",X"FC",X"90",X"FD",X"4D",X"FE",X"07",X"FF",X"BC",X"FF",X"6B",X"00",
		X"16",X"01",X"BB",X"01",X"5E",X"02",X"FA",X"02",X"92",X"03",X"26",X"04",X"B5",X"04",X"40",X"05",
		X"C7",X"05",X"48",X"06",X"C8",X"06",X"43",X"07",X"B9",X"07",X"2B",X"08",X"9B",X"08",X"08",X"09",
		X"71",X"09",X"D6",X"09",X"3A",X"0A",X"98",X"0A",X"F4",X"0A",X"4F",X"0B",X"A4",X"0B",X"F8",X"0B",
		X"48",X"0C",X"97",X"0C",X"E4",X"0C",X"2C",X"0D",X"74",X"0D",X"BB",X"0D",X"FC",X"0D",X"3D",X"0E",
		X"79",X"0E",X"B7",X"0E",X"F0",X"0E",X"29",X"0F",X"5D",X"0F",X"93",X"0F",X"C4",X"0F",X"F8",X"0F",
		X"F2",X"0F",X"9C",X"0F",X"1A",X"0F",X"75",X"0E",X"BF",X"0D",X"FA",X"0C",X"31",X"0C",X"65",X"0B",
		X"99",X"0A",X"CE",X"09",X"08",X"09",X"45",X"08",X"86",X"07",X"CC",X"06",X"17",X"06",X"64",X"05",
		X"BB",X"04",X"13",X"04",X"72",X"03",X"D3",X"02",X"3A",X"02",X"A4",X"01",X"17",X"01",X"89",X"00",
		X"02",X"00",X"7F",X"FF",X"FF",X"FE",X"82",X"FE",X"0B",X"FE",X"96",X"FD",X"25",X"FD",X"B5",X"FC",
		X"4C",X"FC",X"E5",X"FB",X"7E",X"FB",X"1D",X"FB",X"BF",X"FA",X"63",X"FA",X"0A",X"FA",X"B3",X"F9",
		X"61",X"F9",X"0E",X"F9",X"C0",X"F8",X"75",X"F8",X"2C",X"F8",X"E5",X"F7",X"9F",X"F7",X"5B",X"F7",
		X"1B",X"F7",X"DC",X"F6",X"9F",X"F6",X"63",X"F6",X"2B",X"F6",X"F3",X"F5",X"C3",X"F5",X"BF",X"F5",
		X"C4",X"F5",X"C8",X"F5",X"CC",X"F5",X"D2",X"F5",X"D6",X"F5",X"DB",X"F5",X"DE",X"F5",X"E3",X"F5",
		X"E8",X"F5",X"EC",X"F5",X"F2",X"F5",X"F4",X"F5",X"F9",X"F5",X"FE",X"F5",X"03",X"F6",X"08",X"F6",
		X"0A",X"F6",X"11",X"F6",X"16",X"F6",X"19",X"F6",X"1E",X"F6",X"22",X"F6",X"27",X"F6",X"2B",X"F6",
		X"30",X"F6",X"33",X"F6",X"39",X"F6",X"3D",X"F6",X"40",X"F6",X"45",X"F6",X"49",X"F6",X"4E",X"F6",
		X"52",X"F6",X"56",X"F6",X"5A",X"F6",X"60",X"F6",X"62",X"F6",X"67",X"F6",X"6C",X"F6",X"70",X"F6",
		X"74",X"F6",X"78",X"F6",X"7C",X"F6",X"80",X"F6",X"84",X"F6",X"89",X"F6",X"8E",X"F6",X"92",X"F6",
		X"97",X"F6",X"9B",X"F6",X"9F",X"F6",X"A4",X"F6",X"A7",X"F6",X"AC",X"F6",X"B0",X"F6",X"B5",X"F6",
		X"B7",X"F6",X"BC",X"F6",X"C0",X"F6",X"C4",X"F6",X"C8",X"F6",X"CD",X"F6",X"D0",X"F6",X"D5",X"F6",
		X"D9",X"F6",X"DE",X"F6",X"E1",X"F6",X"E5",X"F6",X"EB",X"F6",X"EE",X"F6",X"F1",X"F6",X"F6",X"F6",
		X"F9",X"F6",X"FD",X"F6",X"02",X"F7",X"06",X"F7",X"09",X"F7",X"0E",X"F7",X"12",X"F7",X"14",X"F7",
		X"1A",X"F7",X"1E",X"F7",X"21",X"F7",X"25",X"F7",X"2A",X"F7",X"2C",X"F7",X"32",X"F7",X"36",X"F7",
		X"39",X"F7",X"3F",X"F7",X"41",X"F7",X"47",X"F7",X"4A",X"F7",X"4E",X"F7",X"52",X"F7",X"55",X"F7",
		X"59",X"F7",X"5C",X"F7",X"61",X"F7",X"65",X"F7",X"69",X"F7",X"6C",X"F7",X"71",X"F7",X"75",X"F7",
		X"7A",X"F7",X"7B",X"F7",X"81",X"F7",X"83",X"F7",X"88",X"F7",X"8B",X"F7",X"8F",X"F7",X"93",X"F7",
		X"96",X"F7",X"9A",X"F7",X"9D",X"F7",X"A3",X"F7",X"A6",X"F7",X"AA",X"F7",X"AE",X"F7",X"B1",X"F7",
		X"B4",X"F7",X"B7",X"F7",X"BD",X"F7",X"C0",X"F7",X"C4",X"F7",X"C7",X"F7",X"CC",X"F7",X"CF",X"F7",
		X"D3",X"F7",X"D7",X"F7",X"DB",X"F7",X"DE",X"F7",X"E2",X"F7",X"E4",X"F7",X"E8",X"F7",X"EC",X"F7",
		X"F0",X"F7",X"F5",X"F7",X"F8",X"F7",X"F9",X"F7",X"FF",X"F7",X"01",X"F8",X"07",X"F8",X"07",X"F8",
		X"11",X"F8",X"0A",X"F8",X"87",X"F8",X"7C",X"F9",X"5D",X"FA",X"41",X"FB",X"19",X"FC",X"F1",X"FC",
		X"BE",X"FD",X"89",X"FE",X"4B",X"FF",X"08",X"00",X"BF",X"00",X"72",X"01",X"1E",X"02",X"C7",X"02",
		X"69",X"03",X"08",X"04",X"A1",X"04",X"37",X"05",X"C6",X"05",X"53",X"06",X"D9",X"06",X"5D",X"07",
		X"DC",X"07",X"58",X"08",X"D1",X"08",X"45",X"09",X"B5",X"09",X"22",X"0A",X"8C",X"0A",X"F1",X"0A",
		X"55",X"0B",X"B5",X"0B",X"12",X"0C",X"6B",X"0C",X"C2",X"0C",X"18",X"0D",X"67",X"0D",X"B6",X"0D",
		X"03",X"0E",X"4E",X"0E",X"94",X"0E",X"DA",X"0E",X"1E",X"0F",X"5D",X"0F",X"9C",X"0F",X"CC",X"0F",
		X"B3",X"0F",X"54",X"0F",X"CD",X"0E",X"2C",X"0E",X"79",X"0D",X"BC",X"0C",X"FC",X"0B",X"39",X"0B",
		X"76",X"0A",X"B5",X"09",X"FA",X"08",X"40",X"08",X"8C",X"07",X"DC",X"06",X"31",X"06",X"88",X"05",
		X"E6",X"04",X"4A",X"04",X"AF",X"03",X"1B",X"03",X"8A",X"02",X"FE",X"01",X"75",X"01",X"F0",X"00",
		X"70",X"00",X"F3",X"FF",X"7C",X"FF",X"05",X"FF",X"94",X"FE",X"24",X"FE",X"B9",X"FD",X"51",X"FD",
		X"ED",X"FC",X"8C",X"FC",X"2C",X"FC",X"D0",X"FB",X"77",X"FB",X"1E",X"FB",X"CC",X"FA",X"7A",X"FA",
		X"2C",X"FA",X"DE",X"F9",X"94",X"F9",X"4B",X"F9",X"06",X"F9",X"C4",X"F8",X"83",X"F8",X"42",X"F8",
		X"04",X"F8",X"C8",X"F7",X"8F",X"F7",X"58",X"F7",X"24",X"F7",X"15",X"F7",X"1E",X"F7",X"1E",X"F7",
		X"3C",X"F7",X"C4",X"F7",X"6D",X"F8",X"26",X"F9",X"E8",X"F9",X"B0",X"FA",X"7A",X"FB",X"42",X"FC",
		X"08",X"FD",X"CD",X"FD",X"8B",X"FE",X"46",X"FF",X"FB",X"FF",X"AB",X"00",X"56",X"01",X"FD",X"01",
		X"A0",X"02",X"3E",X"03",X"D6",X"03",X"6C",X"04",X"FB",X"04",X"87",X"05",X"0D",X"06",X"90",X"06",
		X"0E",X"07",X"8D",X"07",X"E8",X"07",X"ED",X"07",X"BB",X"07",X"60",X"07",X"ED",X"06",X"6A",X"06",
		X"E0",X"05",X"4D",X"05",X"BB",X"04",X"28",X"04",X"96",X"03",X"07",X"03",X"79",X"02",X"EF",X"01",
		X"68",X"01",X"E5",X"00",X"68",X"00",X"EB",X"FF",X"74",X"FF",X"00",X"FF",X"8E",X"FE",X"1E",X"FE",
		X"B3",X"FD",X"4C",X"FD",X"E8",X"FC",X"85",X"FC",X"28",X"FC",X"CD",X"FB",X"B4",X"FB",X"E8",X"FB",
		X"48",X"FC",X"C9",X"FC",X"5D",X"FD",X"FD",X"FD",X"A3",X"FE",X"4B",X"FF",X"F3",X"FF",X"9C",X"00",
		X"41",X"01",X"E3",X"01",X"82",X"02",X"1B",X"03",X"B3",X"03",X"44",X"04",X"D3",X"04",X"5E",X"05",
		X"E3",X"05",X"66",X"06",X"E4",X"06",X"5E",X"07",X"D4",X"07",X"47",X"08",X"B8",X"08",X"22",X"09",
		X"8F",X"09",X"DF",X"09",X"DB",X"09",X"9D",X"09",X"36",X"09",X"B5",X"08",X"24",X"08",X"89",X"07",
		X"E9",X"06",X"49",X"06",X"A6",X"05",X"05",X"05",X"68",X"04",X"CF",X"03",X"38",X"03",X"A3",X"02",
		X"14",X"02",X"88",X"01",X"02",X"01",X"7F",X"00",X"FF",X"FF",X"82",X"FF",X"09",X"FF",X"95",X"FE",
		X"23",X"FE",X"B4",X"FD",X"48",X"FD",X"E2",X"FC",X"7D",X"FC",X"51",X"FC",X"73",X"FC",X"C6",X"FC",
		X"3F",X"FD",X"C6",X"FD",X"5E",X"FE",X"FD",X"FE",X"A0",X"FF",X"40",X"00",X"E2",X"00",X"82",X"01",
		X"1F",X"02",X"B8",X"02",X"4D",X"03",X"DF",X"03",X"6D",X"04",X"F6",X"04",X"7B",X"05",X"FD",X"05",
		X"7B",X"06",X"F5",X"06",X"6D",X"07",X"DE",X"07",X"4E",X"08",X"B9",X"08",X"21",X"09",X"89",X"09",
		X"DD",X"09",X"E0",X"09",X"A5",X"09",X"3D",X"09",X"BC",X"08",X"2A",X"08",X"8C",X"07",X"EB",X"06",
		X"46",X"06",X"A1",X"05",X"FE",X"04",X"5E",X"04",X"C0",X"03",X"26",X"03",X"90",X"02",X"FF",X"01",
		X"70",X"01",X"E6",X"00",X"5E",X"00",X"DC",X"FF",X"5E",X"FF",X"E2",X"FE",X"6C",X"FE",X"F8",X"FD",
		X"88",X"FD",X"1A",X"FD",X"B0",X"FC",X"48",X"FC",X"E6",X"FB",X"83",X"FB",X"27",X"FB",X"CA",X"FA",
		X"71",X"FA",X"1E",X"FA",X"CA",X"F9",X"7A",X"F9",X"2D",X"F9",X"E0",X"F8",X"96",X"F8",X"4F",X"F8",
		X"0C",X"F8",X"CA",X"F7",X"8A",X"F7",X"4A",X"F7",X"0B",X"F7",X"D2",X"F6",X"99",X"F6",X"61",X"F6",
		X"33",X"F6",X"30",X"F6",X"37",X"F6",X"3C",X"F6",X"3F",X"F6",X"44",X"F6",X"47",X"F6",X"4F",X"F6",
		X"4E",X"F6",X"59",X"F6",X"55",X"F6",X"BB",X"F6",X"85",X"F7",X"4B",X"F8",X"20",X"F9",X"EC",X"F9",
		X"BE",X"FA",X"89",X"FB",X"54",X"FC",X"15",X"FD",X"D8",X"FD",X"8F",X"FE",X"49",X"FF",X"F8",X"FF",
		X"A5",X"00",X"4B",X"01",X"EE",X"01",X"8A",X"02",X"24",X"03",X"B6",X"03",X"48",X"04",X"D2",X"04",
		X"5B",X"05",X"DC",X"05",X"60",X"06",X"B8",X"06",X"BD",X"06",X"8C",X"06",X"33",X"06",X"C2",X"05",
		X"43",X"05",X"B9",X"04",X"2C",X"04",X"9D",X"03",X"0C",X"03",X"7E",X"02",X"F2",X"01",X"67",X"01",
		X"E0",X"00",X"5E",X"00",X"E0",X"FF",X"62",X"FF",X"EA",X"FE",X"75",X"FE",X"01",X"FE",X"92",X"FD",
		X"27",X"FD",X"BE",X"FC",X"58",X"FC",X"F7",X"FB",X"99",X"FB",X"3B",X"FB",X"E4",X"FA",X"D4",X"FA",
		X"0C",X"FB",X"72",X"FB",X"F4",X"FB",X"8C",X"FC",X"2D",X"FD",X"D7",X"FD",X"81",X"FE",X"2B",X"FF",
		X"D4",X"FF",X"7B",X"00",X"1D",X"01",X"BE",X"01",X"59",X"02",X"F0",X"02",X"83",X"03",X"14",X"04",
		X"9F",X"04",X"27",X"05",X"AB",X"05",X"28",X"06",X"A4",X"06",X"1B",X"07",X"91",X"07",X"00",X"08",
		X"6E",X"08",X"D6",X"08",X"FE",X"08",X"D9",X"08",X"89",X"08",X"14",X"08",X"8D",X"07",X"F8",X"06",
		X"5C",X"06",X"BC",X"05",X"20",X"05",X"7E",X"04",X"E3",X"03",X"48",X"03",X"B3",X"02",X"1F",X"02",
		X"90",X"01",X"03",X"01",X"7B",X"00",X"F8",X"FF",X"79",X"FF",X"FB",X"FE",X"83",X"FE",X"0E",X"FE",
		X"9C",X"FD",X"2D",X"FD",X"C2",X"FC",X"5A",X"FC",X"F6",X"FB",X"93",X"FB",X"35",X"FB",X"D8",X"FA",
		X"7E",X"FA",X"29",X"FA",X"D5",X"F9",X"84",X"F9",X"35",X"F9",X"E7",X"F8",X"9D",X"F8",X"55",X"F8",
		X"10",X"F8",X"CC",X"F7",X"8B",X"F7",X"4B",X"F7",X"0E",X"F7",X"D4",X"F6",X"9A",X"F6",X"64",X"F6",
		X"2A",X"F6",X"17",X"F6",X"1F",X"F6",X"21",X"F6",X"27",X"F6",X"2B",X"F6",X"31",X"F6",X"33",X"F6",
		X"37",X"F6",X"3B",X"F6",X"41",X"F6",X"42",X"F6",X"5B",X"F6",X"05",X"F7",X"D2",X"F7",X"9D",X"F8",
		X"70",X"F9",X"41",X"FA",X"10",X"FB",X"DA",X"FB",X"A2",X"FC",X"65",X"FD",X"23",X"FE",X"DA",X"FE",
		X"90",X"FF",X"3E",X"00",X"E8",X"00",X"8C",X"01",X"2B",X"02",X"C8",X"02",X"5E",X"03",X"F1",X"03",
		X"7E",X"04",X"08",X"05",X"8D",X"05",X"0D",X"06",X"8B",X"06",X"05",X"07",X"7A",X"07",X"ED",X"07",
		X"5C",X"08",X"C7",X"08",X"2E",X"09",X"92",X"09",X"F5",X"09",X"52",X"0A",X"AD",X"0A",X"06",X"0B",
		X"5D",X"0B",X"AE",X"0B",X"01",X"0C",X"4E",X"0C",X"98",X"0C",X"E2",X"0C",X"29",X"0D",X"6C",X"0D",
		X"AE",X"0D",X"EF",X"0D",X"2C",X"0E",X"67",X"0E",X"A0",X"0E",X"DA",X"0E",X"0D",X"0F",X"44",X"0F",
		X"4E",X"0F",X"05",X"0F",X"8A",X"0E",X"ED",X"0D",X"3B",X"0D",X"7B",X"0C",X"B3",X"0B",X"E9",X"0A",
		X"20",X"0A",X"57",X"09",X"93",X"08",X"D2",X"07",X"13",X"07",X"5B",X"06",X"A7",X"05",X"F7",X"04",
		X"4C",X"04",X"A7",X"03",X"06",X"03",X"69",X"02",X"D1",X"01",X"3E",X"01",X"B0",X"00",X"25",X"00",
		X"9E",X"FF",X"1C",X"FF",X"9D",X"FE",X"23",X"FE",X"AA",X"FD",X"35",X"FD",X"C6",X"FC",X"56",X"FC",
		X"EE",X"FB",X"86",X"FB",X"23",X"FB",X"C3",X"FA",X"65",X"FA",X"0B",X"FA",X"B3",X"F9",X"5D",X"F9",
		X"09",X"F9",X"B9",X"F8",X"6B",X"F8",X"21",X"F8",X"D7",X"F7",X"91",X"F7",X"4C",X"F7",X"0A",X"F7",
		X"CA",X"F6",X"8B",X"F6",X"4F",X"F6",X"15",X"F6",X"DC",X"F5",X"A4",X"F5",X"73",X"F5",X"6D",X"F5",
		X"73",X"F5",X"78",X"F5",X"7D",X"F5",X"80",X"F5",X"87",X"F5",X"8A",X"F5",X"91",X"F5",X"93",X"F5",
		X"9B",X"F5",X"9E",X"F5",X"A3",X"F5",X"A7",X"F5",X"AC",X"F5",X"B1",X"F5",X"B5",X"F5",X"BB",X"F5",
		X"BF",X"F5",X"C5",X"F5",X"C9",X"F5",X"CD",X"F5",X"D2",X"F5",X"D8",X"F5",X"DC",X"F5",X"E0",X"F5",
		X"E6",X"F5",X"EA",X"F5",X"EF",X"F5",X"F5",X"F5",X"F7",X"F5",X"FB",X"F5",X"02",X"F6",X"07",X"F6",
		X"0A",X"F6",X"0F",X"F6",X"14",X"F6",X"19",X"F6",X"1D",X"F6",X"21",X"F6",X"26",X"F6",X"2A",X"F6",
		X"30",X"F6",X"32",X"F6",X"37",X"F6",X"3D",X"F6",X"41",X"F6",X"45",X"F6",X"4A",X"F6",X"4E",X"F6",
		X"52",X"F6",X"57",X"F6",X"5D",X"F6",X"61",X"F6",X"67",X"F6",X"6A",X"F6",X"6E",X"F6",X"72",X"F6",
		X"76",X"F6",X"7B",X"F6",X"7F",X"F6",X"83",X"F6",X"87",X"F6",X"8B",X"F6",X"A1",X"F6",X"5F",X"F7",
		X"4F",X"F8",X"2F",X"F9",X"11",X"FA",X"E6",X"FA",X"BB",X"FB",X"88",X"FC",X"50",X"FD",X"10",X"FE",
		X"CF",X"FE",X"84",X"FF",X"36",X"00",X"E1",X"00",X"89",X"01",X"2B",X"02",X"C9",X"02",X"61",X"03",
		X"F5",X"03",X"84",X"04",X"0F",X"05",X"96",X"05",X"1A",X"06",X"9A",X"06",X"16",X"07",X"8D",X"07",
		X"00",X"08",X"70",X"08",X"DC",X"08",X"46",X"09",X"AC",X"09",X"0F",X"0A",X"6F",X"0A",X"CB",X"0A",
		X"25",X"0B",X"7D",X"0B",X"D0",X"0B",X"23",X"0C",X"71",X"0C",X"BC",X"0C",X"08",X"0D",X"4F",X"0D",
		X"94",X"0D",X"D7",X"0D",X"17",X"0E",X"55",X"0E",X"94",X"0E",X"BF",X"0E",X"9B",X"0E",X"37",X"0E",
		X"AC",X"0D",X"07",X"0D",X"52",X"0C",X"92",X"0B",X"CF",X"0A",X"0C",X"0A",X"48",X"09",X"88",X"08",
		X"CA",X"07",X"11",X"07",X"5B",X"06",X"AA",X"05",X"00",X"05",X"57",X"04",X"B5",X"03",X"16",X"03",
		X"7C",X"02",X"E8",X"01",X"56",X"01",X"C9",X"00",X"40",X"00",X"BD",X"FF",X"3B",X"FF",X"C0",X"FE",
		X"44",X"FE",X"FC",X"FD",X"09",X"FE",X"43",X"FE",X"A5",X"FE",X"1C",X"FF",X"A1",X"FF",X"2E",X"00",
		X"BE",X"00",X"52",X"01",X"E5",X"01",X"77",X"02",X"07",X"03",X"92",X"03",X"1B",X"04",X"9E",X"04",
		X"21",X"05",X"9E",X"05",X"18",X"06",X"8F",X"06",X"02",X"07",X"70",X"07",X"DD",X"07",X"47",X"08",
		X"AB",X"08",X"10",X"09",X"6E",X"09",X"CB",X"09",X"1C",X"0A",X"1F",X"0A",X"E0",X"09",X"75",X"09",
		X"EF",X"08",X"55",X"08",X"B2",X"07",X"09",X"07",X"5E",X"06",X"B3",X"05",X"0A",X"05",X"62",X"04",
		X"BE",X"03",X"1D",X"03",X"82",X"02",X"EA",X"01",X"55",X"01",X"C3",X"00",X"38",X"00",X"B2",X"FF",
		X"2C",X"FF",X"AC",X"FE",X"30",X"FE",X"B6",X"FD",X"43",X"FD",X"CF",X"FC",X"62",X"FC",X"F5",X"FB",
		X"B0",X"FB",X"C0",X"FB",X"05",X"FC",X"6F",X"FC",X"F2",X"FC",X"82",X"FD",X"1B",X"FE",X"B8",X"FE",
		X"56",X"FF",X"F4",X"FF",X"8F",X"00",X"29",X"01",X"BF",X"01",X"52",X"02",X"E0",X"02",X"6D",X"03",
		X"F3",X"03",X"78",X"04",X"F7",X"04",X"74",X"05",X"EA",X"05",X"5F",X"06",X"D0",X"06",X"3E",X"07",
		X"A8",X"07",X"0F",X"08",X"72",X"08",X"CF",X"08",X"E5",X"08",X"B2",X"08",X"53",X"08",X"D4",X"07",
		X"42",X"07",X"A7",X"06",X"03",X"06",X"5D",X"05",X"B7",X"04",X"12",X"04",X"70",X"03",X"D0",X"02",
		X"34",X"02",X"9C",X"01",X"08",X"01",X"76",X"00",X"EB",X"FF",X"63",X"FF",X"DE",X"FE",X"5D",X"FE",
		X"E2",X"FD",X"68",X"FD",X"F1",X"FC",X"80",X"FC",X"11",X"FC",X"A5",X"FB",X"3D",X"FB",X"D9",X"FA",
		X"75",X"FA",X"17",X"FA",X"BB",X"F9",X"62",X"F9",X"0A",X"F9",X"B6",X"F8",X"66",X"F8",X"16",X"F8",
		X"CA",X"F7",X"7F",X"F7",X"39",X"F7",X"F4",X"F6",X"AF",X"F6",X"6E",X"F6",X"30",X"F6",X"F2",X"F5",
		X"B6",X"F5",X"7D",X"F5",X"47",X"F5",X"0E",X"F5",X"EB",X"F4",X"EF",X"F4",X"F5",X"F4",X"FA",X"F4",
		X"FF",X"F4",X"04",X"F5",X"08",X"F5",X"0F",X"F5",X"14",X"F5",X"18",X"F5",X"1E",X"F5",X"24",X"F5",
		X"28",X"F5",X"2E",X"F5",X"32",X"F5",X"36",X"F5",X"3B",X"F5",X"41",X"F5",X"45",X"F5",X"4A",X"F5",
		X"51",X"F5",X"54",X"F5",X"59",X"F5",X"60",X"F5",X"64",X"F5",X"6A",X"F5",X"6E",X"F5",X"73",X"F5",
		X"76",X"F5",X"7D",X"F5",X"81",X"F5",X"88",X"F5",X"8B",X"F5",X"90",X"F5",X"94",X"F5",X"99",X"F5",
		X"9F",X"F5",X"A4",X"F5",X"A8",X"F5",X"AD",X"F5",X"B0",X"F5",X"B7",X"F5",X"BB",X"F5",X"C1",X"F5",
		X"C7",X"F5",X"CA",X"F5",X"CE",X"F5",X"D4",X"F5",X"DA",X"F5",X"DC",X"F5",X"E4",X"F5",X"E7",X"F5",
		X"EC",X"F5",X"EF",X"F5",X"F5",X"F5",X"F8",X"F5",X"FE",X"F5",X"02",X"F6",X"0A",X"F6",X"0B",X"F6",
		X"11",X"F6",X"15",X"F6",X"1B",X"F6",X"1E",X"F6",X"26",X"F6",X"26",X"F6",X"2F",X"F6",X"2E",X"F6",
		X"3A",X"F6",X"31",X"F6",X"B2",X"F6",X"AB",X"F7",X"89",X"F8",X"6F",X"F9",X"46",X"FA",X"20",X"FB",
		X"ED",X"FB",X"B8",X"FC",X"7B",X"FD",X"3A",X"FE",X"F3",X"FE",X"A8",X"FF",X"54",X"00",X"FF",X"00",
		X"A0",X"01",X"41",X"02",X"DC",X"02",X"73",X"03",X"04",X"04",X"90",X"04",X"19",X"05",X"9F",X"05",
		X"20",X"06",X"9D",X"06",X"15",X"07",X"8B",X"07",X"FB",X"07",X"6B",X"08",X"D5",X"08",X"3B",X"09",
		X"A0",X"09",X"01",X"0A",X"5F",X"0A",X"BB",X"0A",X"12",X"0B",X"68",X"0B",X"B9",X"0B",X"0A",X"0C",
		X"58",X"0C",X"A2",X"0C",X"EC",X"0C",X"32",X"0D",X"76",X"0D",X"B6",X"0D",X"F8",X"0D",X"33",X"0E",
		X"70",X"0E",X"A8",X"0E",X"DF",X"0E",X"16",X"0F",X"49",X"0F",X"7A",X"0F",X"AA",X"0F",X"DA",X"0F",
		X"05",X"10",X"31",X"10",X"5B",X"10",X"82",X"10",X"AA",X"10",X"CF",X"10",X"F3",X"10",X"17",X"11",
		X"36",X"11",X"58",X"11",X"76",X"11",X"95",X"11",X"B0",X"11",X"CD",X"11",X"E7",X"11",X"FF",X"11",
		X"19",X"12",X"2F",X"12",X"45",X"12",X"5D",X"12",X"52",X"12",X"F2",X"11",X"60",X"11",X"AA",X"10",
		X"DF",X"0F",X"04",X"0F",X"26",X"0E",X"44",X"0D",X"64",X"0C",X"82",X"0B",X"A6",X"0A",X"CF",X"09",
		X"FB",X"08",X"2D",X"08",X"65",X"07",X"A2",X"06",X"E2",X"05",X"2C",X"05",X"79",X"04",X"C8",X"03",
		X"20",X"03",X"7C",X"02",X"DB",X"01",X"41",X"01",X"AA",X"00",X"19",X"00",X"8D",X"FF",X"03",X"FF",
		X"7E",X"FE",X"FD",X"FD",X"7E",X"FD",X"04",X"FD",X"90",X"FC",X"1D",X"FC",X"AE",X"FB",X"42",X"FB",
		X"D9",X"FA",X"75",X"FA",X"13",X"FA",X"B3",X"F9",X"57",X"F9",X"FC",X"F8",X"A5",X"F8",X"51",X"F8",
		X"FF",X"F7",X"B1",X"F7",X"64",X"F7",X"1A",X"F7",X"D2",X"F6",X"8D",X"F6",X"48",X"F6",X"08",X"F6",
		X"C8",X"F5",X"8B",X"F5",X"4E",X"F5",X"2B",X"F5",X"5D",X"F5",X"C7",X"F5",X"57",X"F6",X"00",X"F7",
		X"B8",X"F7",X"77",X"F8",X"39",X"F9",X"FE",X"F9",X"BF",X"FA",X"81",X"FB",X"3C",X"FC",X"F6",X"FC",
		X"AA",X"FD",X"58",X"FE",X"03",X"FF",X"AA",X"FF",X"49",X"00",X"E7",X"00",X"7E",X"01",X"13",X"02",
		X"A2",X"02",X"2B",X"03",X"B3",X"03",X"35",X"04",X"B5",X"04",X"30",X"05",X"A5",X"05",X"1A",X"06",
		X"8A",X"06",X"F7",X"06",X"60",X"07",X"C6",X"07",X"28",X"08",X"89",X"08",X"E5",X"08",X"40",X"09",
		X"98",X"09",X"EC",X"09",X"3B",X"0A",X"8C",X"0A",X"D7",X"0A",X"24",X"0B",X"6A",X"0B",X"B0",X"0B",
		X"F3",X"0B",X"33",X"0C",X"72",X"0C",X"AF",X"0C",X"EA",X"0C",X"23",X"0D",X"59",X"0D",X"8E",X"0D",
		X"C1",X"0D",X"F3",X"0D",X"14",X"0E",X"E4",X"0D",X"75",X"0D",X"DF",X"0C",X"31",X"0C",X"72",X"0B",
		X"AB",X"0A",X"E0",X"09",X"12",X"09",X"49",X"08",X"7F",X"07",X"BB",X"06",X"F9",X"05",X"3F",X"05",
		X"89",X"04",X"D4",X"03",X"27",X"03",X"7E",X"02",X"DA",X"01",X"3A",X"01",X"9F",X"00",X"09",X"00",
		X"77",X"FF",X"EB",X"FE",X"62",X"FE",X"DA",X"FD",X"5B",X"FD",X"DB",X"FC",X"90",X"FC",X"98",X"FC",
		X"D1",X"FC",X"31",X"FD",X"A4",X"FD",X"25",X"FE",X"B0",X"FE",X"3E",X"FF",X"CD",X"FF",X"5C",X"00",
		X"EB",X"00",X"77",X"01",X"00",X"02",X"86",X"02",X"07",X"03",X"88",X"03",X"02",X"04",X"7B",X"04",
		X"EF",X"04",X"60",X"05",X"CD",X"05",X"37",X"06",X"9E",X"06",X"02",X"07",X"62",X"07",X"BF",X"07",
		X"1C",X"08",X"6A",X"08",X"6C",X"08",X"29",X"08",X"BB",X"07",X"33",X"07",X"98",X"06",X"F4",X"05",
		X"4A",X"05",X"9D",X"04",X"F1",X"03",X"46",X"03",X"9F",X"02",X"FA",X"01",X"58",X"01",X"BD",X"00",
		X"23",X"00",X"90",X"FF",X"FF",X"FE",X"72",X"FE",X"E9",X"FD",X"65",X"FD",X"E6",X"FC",X"67",X"FC",
		X"EF",X"FB",X"79",X"FB",X"06",X"FB",X"98",X"FA",X"2D",X"FA",X"C7",X"F9",X"60",X"F9",X"FF",X"F8",
		X"A0",X"F8",X"44",X"F8",X"EB",X"F7",X"95",X"F7",X"41",X"F7",X"EF",X"F6",X"A2",X"F6",X"55",X"F6",
		X"0B",X"F6",X"C5",X"F5",X"80",X"F5",X"3C",X"F5",X"FA",X"F4",X"BD",X"F4",X"7F",X"F4",X"46",X"F4",
		X"0C",X"F4",X"D5",X"F3",X"9E",X"F3",X"74",X"F3",X"78",X"F3",X"7D",X"F3",X"82",X"F3",X"88",X"F3",
		X"8E",X"F3",X"95",X"F3",X"99",X"F3",X"AF",X"F3",X"48",X"F4",X"0B",X"F5",X"D3",X"F5",X"A2",X"F6",
		X"70",X"F7",X"3F",X"F8",X"0A",X"F9",X"D5",X"F9",X"98",X"FA",X"59",X"FB",X"15",X"FC",X"CA",X"FC",
		X"7C",X"FD",X"29",X"FE",X"D1",X"FE",X"74",X"FF",X"0F",X"00",X"A9",X"00",X"3D",X"01",X"CF",X"01",
		X"59",X"02",X"E1",X"02",X"64",X"03",X"E5",X"03",X"60",X"04",X"D8",X"04",X"4B",X"05",X"BC",X"05",
		X"2B",X"06",X"96",X"06",X"FB",X"06",X"5F",X"07",X"BF",X"07",X"1E",X"08",X"78",X"08",X"D0",X"08",
		X"24",X"09",X"77",X"09",X"C6",X"09",X"15",X"0A",X"5E",X"0A",X"A6",X"0A",X"ED",X"0A",X"30",X"0B",
		X"72",X"0B",X"B2",X"0B",X"EF",X"0B",X"2B",X"0C",X"64",X"0C",X"9A",X"0C",X"D1",X"0C",X"04",X"0D",
		X"37",X"0D",X"66",X"0D",X"95",X"0D",X"C3",X"0D",X"EE",X"0D",X"19",X"0E",X"3F",X"0E",X"67",X"0E",
		X"8D",X"0E",X"B0",X"0E",X"D6",X"0E",X"F6",X"0E",X"16",X"0F",X"35",X"0F",X"54",X"0F",X"71",X"0F",
		X"8D",X"0F",X"A7",X"0F",X"C2",X"0F",X"DA",X"0F",X"F3",X"0F",X"09",X"10",X"1E",X"10",X"34",X"10",
		X"47",X"10",X"59",X"10",X"6F",X"10",X"6D",X"10",X"1A",X"10",X"8C",X"0F",X"D9",X"0E",X"0E",X"0E",
		X"34",X"0D",X"54",X"0C",X"6F",X"0B",X"8A",X"0A",X"A9",X"09",X"C9",X"08",X"EF",X"07",X"19",X"07",
		X"48",X"06",X"7E",X"05",X"B7",X"04",X"F7",X"03",X"3D",X"03",X"88",X"02",X"D6",X"01",X"2B",X"01",
		X"85",X"00",X"E4",X"FF",X"47",X"FF",X"AF",X"FE",X"1B",X"FE",X"8E",X"FD",X"02",X"FD",X"7B",X"FC",
		X"F8",X"FB",X"78",X"FB",X"FE",X"FA",X"85",X"FA",X"13",X"FA",X"A3",X"F9",X"36",X"F9",X"CC",X"F8",
		X"66",X"F8",X"01",X"F8",X"A2",X"F7",X"44",X"F7",X"EB",X"F6",X"93",X"F6",X"3E",X"F6",X"EB",X"F5",
		X"9D",X"F5",X"4F",X"F5",X"04",X"F5",X"BB",X"F4",X"76",X"F4",X"32",X"F4",X"F1",X"F3",X"AF",X"F3",
		X"75",X"F3",X"36",X"F3",X"27",X"F3",X"6C",X"F3",X"E0",X"F3",X"79",X"F4",X"25",X"F5",X"DF",X"F5",
		X"9F",X"F6",X"62",X"F7",X"27",X"F8",X"E8",X"F8",X"A8",X"F9",X"63",X"FA",X"19",X"FB",X"CD",X"FB",
		X"79",X"FC",X"23",X"FD",X"C8",X"FD",X"68",X"FE",X"04",X"FF",X"9A",X"FF",X"2B",X"00",X"B9",X"00",
		X"43",X"01",X"C9",X"01",X"4C",X"02",X"C9",X"02",X"44",X"03",X"B3",X"03",X"D5",X"03",X"B0",X"03",
		X"62",X"03",X"F2",X"02",X"75",X"02",X"EB",X"01",X"5A",X"01",X"C3",X"00",X"31",X"00",X"9C",X"FF",
		X"0B",X"FF",X"7B",X"FE",X"F2",X"FD",X"68",X"FD",X"E3",X"FC",X"61",X"FC",X"E4",X"FB",X"68",X"FB",
		X"F2",X"FA",X"7F",X"FA",X"10",X"FA",X"A3",X"F9",X"39",X"F9",X"D4",X"F8",X"72",X"F8",X"11",X"F8",
		X"B3",X"F7",X"5A",X"F7",X"03",X"F7",X"AE",X"F6",X"5A",X"F6",X"0B",X"F6",X"C0",X"F5",X"74",X"F5",
		X"2D",X"F5",X"E7",X"F4",X"A2",X"F4",X"62",X"F4",X"22",X"F4",X"E4",X"F3",X"A8",X"F3",X"70",X"F3",
		X"36",X"F3",X"02",X"F3",X"CB",X"F2",X"BA",X"F2",X"C2",X"F2",X"C8",X"F2",X"CE",X"F2",X"D3",X"F2",
		X"DB",X"F2",X"E1",X"F2",X"E7",X"F2",X"ED",X"F2",X"F3",X"F2",X"FA",X"F2",X"00",X"F3",X"06",X"F3",
		X"13",X"F3",X"AF",X"F3",X"83",X"F4",X"55",X"F5",X"2C",X"F6",X"FD",X"F6",X"D0",X"F7",X"9C",X"F8",
		X"67",X"F9",X"2D",X"FA",X"EE",X"FA",X"A7",X"FB",X"5E",X"FC",X"0E",X"FD",X"BA",X"FD",X"60",X"FE",
		X"03",X"FF",X"9F",X"FF",X"39",X"00",X"CD",X"00",X"5A",X"01",X"E6",X"01",X"6B",X"02",X"F2",X"02",
		X"58",X"03",X"69",X"03",X"41",X"03",X"F0",X"02",X"85",X"02",X"09",X"02",X"84",X"01",X"FB",X"00",
		X"6D",X"00",X"E1",X"FF",X"55",X"FF",X"CB",X"FE",X"45",X"FE",X"C0",X"FD",X"40",X"FD",X"C1",X"FC",
		X"48",X"FC",X"D1",X"FB",X"5E",X"FB",X"EC",X"FA",X"81",X"FA",X"16",X"FA",X"B0",X"F9",X"4C",X"F9",
		X"ED",X"F8",X"8F",X"F8",X"35",X"F8",X"DF",X"F7",X"C4",X"F7",X"F9",X"F7",X"5B",X"F8",X"DE",X"F8",
		X"74",X"F9",X"17",X"FA",X"C2",X"FA",X"6E",X"FB",X"1A",X"FC",X"C6",X"FC",X"71",X"FD",X"17",X"FE",
		X"B9",X"FE",X"59",X"FF",X"F1",X"FF",X"86",X"00",X"19",X"01",X"A6",X"01",X"31",X"02",X"B5",X"02",
		X"37",X"03",X"B6",X"03",X"2F",X"04",X"A6",X"04",X"19",X"05",X"87",X"05",X"F4",X"05",X"5C",X"06",
		X"C0",X"06",X"23",X"07",X"83",X"07",X"DF",X"07",X"39",X"08",X"90",X"08",X"E3",X"08",X"35",X"09",
		X"82",X"09",X"D0",X"09",X"18",X"0A",X"61",X"0A",X"A6",X"0A",X"E8",X"0A",X"29",X"0B",X"68",X"0B",
		X"A4",X"0B",X"E0",X"0B",X"18",X"0C",X"4E",X"0C",X"82",X"0C",X"B6",X"0C",X"E8",X"0C",X"18",X"0D",
		X"46",X"0D",X"71",X"0D",X"9C",X"0D",X"C7",X"0D",X"EF",X"0D",X"14",X"0E",X"3B",X"0E",X"5E",X"0E",
		X"81",X"0E",X"A2",X"0E",X"C2",X"0E",X"E0",X"0E",X"01",X"0F",X"1C",X"0F",X"37",X"0F",X"51",X"0F",
		X"6C",X"0F",X"84",X"0F",X"9C",X"0F",X"B3",X"0F",X"C6",X"0F",X"DB",X"0F",X"F1",X"0F",X"03",X"10",
		X"16",X"10",X"27",X"10",X"37",X"10",X"46",X"10",X"56",X"10",X"5E",X"10",X"54",X"10",X"4C",X"10",
		X"43",X"10",X"39",X"10",X"2F",X"10",X"27",X"10",X"1C",X"10",X"14",X"10",X"0A",X"10",X"02",X"10",
		X"F8",X"0F",X"EF",X"0F",X"E7",X"0F",X"DC",X"0F",X"D3",X"0F",X"CC",X"0F",X"C2",X"0F",X"B8",X"0F",
		X"AF",X"0F",X"A6",X"0F",X"9D",X"0F",X"93",X"0F",X"8C",X"0F",X"82",X"0F",X"78",X"0F",X"71",X"0F",
		X"67",X"0F",X"5E",X"0F",X"56",X"0F",X"4C",X"0F",X"44",X"0F",X"3C",X"0F",X"32",X"0F",X"2A",X"0F",
		X"20",X"0F",X"17",X"0F",X"0E",X"0F",X"06",X"0F",X"FC",X"0E",X"F4",X"0E",X"EA",X"0E",X"E2",X"0E",
		X"DA",X"0E",X"D1",X"0E",X"C9",X"0E",X"C0",X"0E",X"B8",X"0E",X"AE",X"0E",X"A6",X"0E",X"9F",X"0E",
		X"96",X"0E",X"8C",X"0E",X"84",X"0E",X"7B",X"0E",X"73",X"0E",X"6A",X"0E",X"63",X"0E",X"59",X"0E",
		X"52",X"0E",X"48",X"0E",X"41",X"0E",X"37",X"0E",X"30",X"0E",X"27",X"0E",X"1F",X"0E",X"16",X"0E",
		X"0E",X"0E",X"05",X"0E",X"FD",X"0D",X"F5",X"0D",X"ED",X"0D",X"E5",X"0D",X"DB",X"0D",X"D3",X"0D",
		X"CC",X"0D",X"C4",X"0D",X"BC",X"0D",X"B3",X"0D",X"AC",X"0D",X"A4",X"0D",X"9B",X"0D",X"94",X"0D",
		X"8B",X"0D",X"82",X"0D",X"7B",X"0D",X"72",X"0D",X"6A",X"0D",X"62",X"0D",X"5A",X"0D",X"52",X"0D",
		X"4A",X"0D",X"43",X"0D",X"3B",X"0D",X"32",X"0D",X"2B",X"0D",X"22",X"0D",X"1A",X"0D",X"11",X"0D",
		X"0A",X"0D",X"03",X"0D",X"FB",X"0C",X"F3",X"0C",X"EC",X"0C",X"E2",X"0C",X"DC",X"0C",X"D3",X"0C",
		X"CC",X"0C",X"C3",X"0C",X"BD",X"0C",X"B4",X"0C",X"AD",X"0C",X"A5",X"0C",X"9F",X"0C",X"93",X"0C",
		X"92",X"0C",X"60",X"0C",X"7D",X"0B",X"82",X"0A",X"8A",X"09",X"92",X"08",X"9E",X"07",X"AF",X"06",
		X"C6",X"05",X"E2",X"04",X"02",X"04",X"29",X"03",X"58",X"02",X"8A",X"01",X"C3",X"00",X"03",X"00",
		X"48",X"FF",X"91",X"FE",X"E1",X"FD",X"35",X"FD",X"8F",X"FC",X"EC",X"FB",X"50",X"FB",X"B8",X"FA",
		X"25",X"FA",X"95",X"F9",X"0B",X"F9",X"85",X"F8",X"03",X"F8",X"84",X"F7",X"09",X"F7",X"92",X"F6",
		X"1E",X"F6",X"AF",X"F5",X"43",X"F5",X"D9",X"F4",X"74",X"F4",X"11",X"F4",X"B2",X"F3",X"55",X"F3",
		X"FC",X"F2",X"A5",X"F2",X"50",X"F2",X"FF",X"F1",X"B1",X"F1",X"66",X"F1",X"1B",X"F1",X"D4",X"F0",
		X"8E",X"F0",X"4C",X"F0",X"0C",X"F0",X"CD",X"EF",X"8F",X"EF",X"54",X"EF",X"1D",X"EF",X"E5",X"EE",
		X"B2",X"EE",X"7C",X"EE",X"59",X"EE",X"60",X"EE",X"69",X"EE",X"71",X"EE",X"7A",X"EE",X"81",X"EE",
		X"88",X"EE",X"93",X"EE",X"99",X"EE",X"A3",X"EE",X"AA",X"EE",X"B2",X"EE",X"BA",X"EE",X"C3",X"EE",
		X"CB",X"EE",X"D4",X"EE",X"DA",X"EE",X"E2",X"EE",X"E9",X"EE",X"F3",X"EE",X"FA",X"EE",X"04",X"EF",
		X"09",X"EF",X"14",X"EF",X"17",X"EF",X"26",X"EF",X"23",X"EF",X"69",X"EF",X"4B",X"F0",X"29",X"F1",
		X"0A",X"F2",X"E6",X"F2",X"BF",X"F3",X"90",X"F4",X"60",X"F5",X"27",X"F6",X"ED",X"F6",X"AA",X"F7",
		X"65",X"F8",X"18",X"F9",X"C7",X"F9",X"71",X"FA",X"15",X"FB",X"B5",X"FB",X"51",X"FC",X"E7",X"FC",
		X"78",X"FD",X"08",X"FE",X"90",X"FE",X"17",X"FF",X"99",X"FF",X"16",X"00",X"8F",X"00",X"05",X"01",
		X"78",X"01",X"E8",X"01",X"53",X"02",X"BD",X"02",X"22",X"03",X"84",X"03",X"E3",X"03",X"41",X"04",
		X"9A",X"04",X"F1",X"04",X"45",X"05",X"98",X"05",X"E6",X"05",X"33",X"06",X"7D",X"06",X"C6",X"06",
		X"0C",X"07",X"4F",X"07",X"90",X"07",X"CF",X"07",X"0C",X"08",X"48",X"08",X"81",X"08",X"B8",X"08",
		X"EF",X"08",X"23",X"09",X"55",X"09",X"86",X"09",X"B3",X"09",X"E2",X"09",X"0E",X"0A",X"39",X"0A",
		X"61",X"0A",X"89",X"0A",X"B0",X"0A",X"D6",X"0A",X"F7",X"0A",X"1A",X"0B",X"3B",X"0B",X"5A",X"0B",
		X"7A",X"0B",X"97",X"0B",X"B5",X"0B",X"D1",X"0B",X"EC",X"0B",X"05",X"0C",X"1D",X"0C",X"36",X"0C",
		X"4B",X"0C",X"5D",X"0C",X"2B",X"0C",X"B0",X"0B",X"0C",X"0B",X"4B",X"0A",X"79",X"09",X"9E",X"08",
		X"BF",X"07",X"DE",X"06",X"FF",X"05",X"22",X"05",X"49",X"04",X"75",X"03",X"A7",X"02",X"DC",X"01",
		X"17",X"01",X"59",X"00",X"A1",X"FF",X"ED",X"FE",X"3C",X"FE",X"94",X"FD",X"ED",X"FC",X"4E",X"FC",
		X"B3",X"FB",X"1D",X"FB",X"8A",X"FA",X"FD",X"F9",X"72",X"F9",X"ED",X"F8",X"6D",X"F8",X"EE",X"F7",
		X"75",X"F7",X"FE",X"F6",X"8D",X"F6",X"1D",X"F6",X"B2",X"F5",X"49",X"F5",X"E5",X"F4",X"83",X"F4",
		X"26",X"F4",X"C7",X"F3",X"70",X"F3",X"1A",X"F3",X"C6",X"F2",X"76",X"F2",X"27",X"F2",X"DD",X"F1",
		X"94",X"F1",X"4B",X"F1",X"08",X"F1",X"C5",X"F0",X"84",X"F0",X"46",X"F0",X"0A",X"F0",X"D0",X"EF",
		X"98",X"EF",X"60",X"EF",X"2D",X"EF",X"FA",X"EE",X"E7",X"EE",X"F2",X"EE",X"F7",X"EE",X"00",X"EF",
		X"08",X"EF",X"10",X"EF",X"18",X"EF",X"20",X"EF",X"29",X"EF",X"30",X"EF",X"38",X"EF",X"40",X"EF",
		X"48",X"EF",X"50",X"EF",X"59",X"EF",X"60",X"EF",X"68",X"EF",X"70",X"EF",X"78",X"EF",X"7E",X"EF",
		X"86",X"EF",X"8E",X"EF",X"96",X"EF",X"9C",X"EF",X"A6",X"EF",X"AB",X"EF",X"B5",X"EF",X"BC",X"EF",
		X"C5",X"EF",X"CB",X"EF",X"E2",X"EF",X"AA",X"F0",X"93",X"F1",X"71",X"F2",X"51",X"F3",X"28",X"F4",
		X"FE",X"F4",X"CD",X"F5",X"98",X"F6",X"5B",X"F7",X"1D",X"F8",X"D6",X"F8",X"8D",X"F9",X"3B",X"FA",
		X"E6",X"FA",X"8C",X"FB",X"2E",X"FC",X"CA",X"FC",X"62",X"FD",X"F4",X"FD",X"84",X"FE",X"0E",X"FF",
		X"62",X"FF",X"64",X"FF",X"35",X"FF",X"E1",X"FE",X"79",X"FE",X"00",X"FE",X"82",X"FD",X"FD",X"FC",
		X"77",X"FC",X"F1",X"FB",X"6D",X"FB",X"E9",X"FA",X"6C",X"FA",X"EF",X"F9",X"76",X"F9",X"FE",X"F8",
		X"8B",X"F8",X"1A",X"F8",X"AE",X"F7",X"45",X"F7",X"DF",X"F6",X"7D",X"F6",X"1D",X"F6",X"BF",X"F5",
		X"65",X"F5",X"0D",X"F5",X"B7",X"F4",X"73",X"F4",X"7A",X"F4",X"C5",X"F4",X"38",X"F5",X"C7",X"F5",
		X"67",X"F6",X"11",X"F7",X"C0",X"F7",X"71",X"F8",X"23",X"F9",X"D1",X"F9",X"7D",X"FA",X"25",X"FB",
		X"CA",X"FB",X"69",X"FC",X"09",X"FD",X"A0",X"FD",X"33",X"FE",X"C3",X"FE",X"4E",X"FF",X"D7",X"FF",
		X"59",X"00",X"D9",X"00",X"55",X"01",X"CC",X"01",X"41",X"02",X"B4",X"02",X"20",X"03",X"8C",X"03",
		X"F2",X"03",X"56",X"04",X"B8",X"04",X"15",X"05",X"70",X"05",X"C9",X"05",X"1D",X"06",X"72",X"06",
		X"C2",X"06",X"0F",X"07",X"5B",X"07",X"A3",X"07",X"EA",X"07",X"2F",X"08",X"71",X"08",X"B1",X"08",
		X"EF",X"08",X"2B",X"09",X"66",X"09",X"9E",X"09",X"D4",X"09",X"09",X"0A",X"3C",X"0A",X"6F",X"0A",
		X"9D",X"0A",X"CD",X"0A",X"F9",X"0A",X"23",X"0B",X"4D",X"0B",X"74",X"0B",X"9B",X"0B",X"C1",X"0B",
		X"E5",X"0B",X"07",X"0C",X"28",X"0C",X"49",X"0C",X"68",X"0C",X"87",X"0C",X"A4",X"0C",X"BF",X"0C",
		X"DA",X"0C",X"F4",X"0C",X"0D",X"0D",X"26",X"0D",X"3C",X"0D",X"52",X"0D",X"66",X"0D",X"7C",X"0D",
		X"8F",X"0D",X"A2",X"0D",X"B3",X"0D",X"C5",X"0D",X"D4",X"0D",X"E6",X"0D",X"D6",X"0D",X"76",X"0D",
		X"DF",X"0C",X"26",X"0C",X"53",X"0B",X"78",X"0A",X"94",X"09",X"AE",X"08",X"C8",X"07",X"E4",X"06",
		X"05",X"06",X"2A",X"05",X"55",X"04",X"83",X"03",X"B8",X"02",X"F1",X"01",X"31",X"01",X"76",X"00",
		X"C1",X"FF",X"12",X"FF",X"66",X"FE",X"C0",X"FD",X"1F",X"FD",X"82",X"FC",X"EA",X"FB",X"56",X"FB",
		X"C8",X"FA",X"40",X"FA",X"FC",X"F9",X"05",X"FA",X"3C",X"FA",X"92",X"FA",X"FE",X"FA",X"77",X"FB",
		X"F7",X"FB",X"7C",X"FC",X"01",X"FD",X"88",X"FD",X"0B",X"FE",X"8E",X"FE",X"0C",X"FF",X"88",X"FF",
		X"01",X"00",X"77",X"00",X"E9",X"00",X"5A",X"01",X"C5",X"01",X"2E",X"02",X"94",X"02",X"F7",X"02",
		X"57",X"03",X"B2",X"03",X"0F",X"04",X"64",X"04",X"BC",X"04",X"F9",X"04",X"E0",X"04",X"8E",X"04",
		X"15",X"04",X"82",X"03",X"E1",X"02",X"37",X"02",X"89",X"01",X"D8",X"00",X"28",X"00",X"7D",X"FF",
		X"D1",X"FE",X"2A",X"FE",X"88",X"FD",X"E9",X"FC",X"4D",X"FC",X"B6",X"FB",X"26",X"FB",X"97",X"FA",
		X"0E",X"FA",X"88",X"F9",X"06",X"F9",X"88",X"F8",X"0F",X"F8",X"99",X"F7",X"25",X"F7",X"B6",X"F6",
		X"4A",X"F6",X"1B",X"F6",X"38",X"F6",X"88",X"F6",X"F7",X"F6",X"7B",X"F7",X"0F",X"F8",X"A9",X"F8",
		X"45",X"F9",X"E2",X"F9",X"82",X"FA",X"1A",X"FB",X"B3",X"FB",X"48",X"FC",X"DB",X"FC",X"6A",X"FD",
		X"F3",X"FD",X"7A",X"FE",X"FC",X"FE",X"7C",X"FF",X"F8",X"FF",X"6E",X"00",X"E1",X"00",X"52",X"01",
		X"C0",X"01",X"29",X"02",X"8F",X"02",X"F4",X"02",X"55",X"03",X"B3",X"03",X"0D",X"04",X"66",X"04",
		X"BB",X"04",X"0C",X"05",X"5E",X"05",X"AC",X"05",X"F6",X"05",X"40",X"06",X"87",X"06",X"CA",X"06",
		X"0E",X"07",X"4E",X"07",X"8C",X"07",X"C7",X"07",X"02",X"08",X"3B",X"08",X"71",X"08",X"A6",X"08",
		X"D9",X"08",X"0A",X"09",X"3A",X"09",X"6A",X"09",X"95",X"09",X"C2",X"09",X"EA",X"09",X"15",X"0A",
		X"0F",X"0A",X"B7",X"09",X"2F",X"09",X"85",X"08",X"C9",X"07",X"FD",X"06",X"2E",X"06",X"5B",X"05",
		X"8B",X"04",X"BA",X"03",X"EF",X"02",X"24",X"02",X"62",X"01",X"A1",X"00",X"E8",X"FF",X"33",X"FF",
		X"83",X"FE",X"D9",X"FD",X"32",X"FD",X"91",X"FC",X"F5",X"FB",X"5D",X"FB",X"C9",X"FA",X"3B",X"FA",
		X"B0",X"F9",X"2A",X"F9",X"A8",X"F8",X"29",X"F8",X"AF",X"F7",X"36",X"F7",X"C5",X"F6",X"54",X"F6",
		X"E8",X"F5",X"80",X"F5",X"18",X"F5",X"B9",X"F4",X"58",X"F4",X"FC",X"F3",X"A3",X"F3",X"4A",X"F3",
		X"F6",X"F2",X"A6",X"F2",X"56",X"F2",X"0A",X"F2",X"C1",X"F1",X"79",X"F1",X"34",X"F1",X"F1",X"F0",
		X"B1",X"F0",X"73",X"F0",X"36",X"F0",X"FB",X"EF",X"C3",X"EF",X"8C",X"EF",X"5C",X"EF",X"72",X"EF",
		X"CF",X"EF",X"5A",X"F0",X"FF",X"F0",X"B6",X"F1",X"79",X"F2",X"3F",X"F3",X"08",X"F4",X"D1",X"F4",
		X"96",X"F5",X"59",X"F6",X"17",X"F7",X"D1",X"F7",X"86",X"F8",X"37",X"F9",X"E4",X"F9",X"8C",X"FA",
		X"2F",X"FB",X"CC",X"FB",X"65",X"FC",X"FA",X"FC",X"8A",X"FD",X"17",X"FE",X"9E",X"FE",X"24",X"FF",
		X"A4",X"FF",X"22",X"00",X"7E",X"00",X"86",X"00",X"54",X"00",X"FC",X"FF",X"8C",X"FF",X"0A",X"FF",
		X"81",X"FE",X"F1",X"FD",X"61",X"FD",X"CF",X"FC",X"3E",X"FC",X"B1",X"FB",X"26",X"FB",X"9D",X"FA",
		X"1A",X"FA",X"99",X"F9",X"1C",X"F9",X"A1",X"F8",X"2B",X"F8",X"B6",X"F7",X"4A",X"F7",X"DD",X"F6",
		X"74",X"F6",X"0E",X"F6",X"AB",X"F5",X"4D",X"F5",X"F2",X"F4",X"99",X"F4",X"82",X"F4",X"B4",X"F4",
		X"18",X"F5",X"9D",X"F5",X"32",X"F6",X"D4",X"F6",X"7B",X"F7",X"26",X"F8",X"D2",X"F8",X"7E",X"F9",
		X"25",X"FA",X"C9",X"FA",X"6C",X"FB",X"0A",X"FC",X"A3",X"FC",X"38",X"FD",X"CA",X"FD",X"56",X"FE",
		X"DF",X"FE",X"64",X"FF",X"E6",X"FF",X"64",X"00",X"DC",X"00",X"52",X"01",X"C5",X"01",X"33",X"02",
		X"A2",X"02",X"F7",X"02",X"F8",X"02",X"BD",X"02",X"58",X"02",X"DB",X"01",X"4F",X"01",X"B6",X"00",
		X"1B",X"00",X"7D",X"FF",X"DC",X"FE",X"41",X"FE",X"A5",X"FD",X"0E",X"FD",X"7A",X"FC",X"EB",X"FB",
		X"5E",X"FB",X"D7",X"FA",X"51",X"FA",X"D0",X"F9",X"52",X"F9",X"DA",X"F8",X"64",X"F8",X"F1",X"F7",
		X"83",X"F7",X"17",X"F7",X"AF",X"F6",X"4B",X"F6",X"EA",X"F5",X"8C",X"F5",X"2F",X"F5",X"D7",X"F4",
		X"7F",X"F4",X"2D",X"F4",X"DB",X"F3",X"8D",X"F3",X"41",X"F3",X"F8",X"F2",X"B1",X"F2",X"6D",X"F2",
		X"2A",X"F2",X"E9",X"F1",X"AC",X"F1",X"70",X"F1",X"34",X"F1",X"FD",X"F0",X"C7",X"F0",X"92",X"F0",
		X"60",X"F0",X"55",X"F0",X"60",X"F0",X"67",X"F0",X"6F",X"F0",X"75",X"F0",X"7F",X"F0",X"85",X"F0",
		X"8C",X"F0",X"92",X"F0",X"9A",X"F0",X"A2",X"F0",X"AA",X"F0",X"B1",X"F0",X"B9",X"F0",X"BF",X"F0",
		X"C7",X"F0",X"CE",X"F0",X"D7",X"F0",X"DE",X"F0",X"E7",X"F0",X"EC",X"F0",X"F5",X"F0",X"FA",X"F0",
		X"02",X"F1",X"08",X"F1",X"10",X"F1",X"18",X"F1",X"1E",X"F1",X"26",X"F1",X"2E",X"F1",X"34",X"F1",
		X"3C",X"F1",X"43",X"F1",X"4B",X"F1",X"51",X"F1",X"58",X"F1",X"60",X"F1",X"67",X"F1",X"6D",X"F1",
		X"77",X"F1",X"7C",X"F1",X"83",X"F1",X"8B",X"F1",X"91",X"F1",X"98",X"F1",X"9F",X"F1",X"A6",X"F1",
		X"AF",X"F1",X"B5",X"F1",X"BB",X"F1",X"C3",X"F1",X"CA",X"F1",X"D1",X"F1",X"D7",X"F1",X"DD",X"F1",
		X"E6",X"F1",X"ED",X"F1",X"F3",X"F1",X"F9",X"F1",X"02",X"F2",X"06",X"F2",X"0F",X"F2",X"14",X"F2",
		X"1D",X"F2",X"23",X"F2",X"2A",X"F2",X"2F",X"F2",X"37",X"F2",X"3D",X"F2",X"45",X"F2",X"4B",X"F2",
		X"51",X"F2",X"59",X"F2",X"5F",X"F2",X"67",X"F2",X"6C",X"F2",X"73",X"F2",X"7B",X"F2",X"7F",X"F2",
		X"86",X"F2",X"8C",X"F2",X"95",X"F2",X"9C",X"F2",X"A2",X"F2",X"A8",X"F2",X"B0",X"F2",X"B5",X"F2",
		X"BE",X"F2",X"C3",X"F2",X"CB",X"F2",X"CF",X"F2",X"D7",X"F2",X"DC",X"F2",X"E5",X"F2",X"E9",X"F2",
		X"F1",X"F2",X"F5",X"F2",X"FF",X"F2",X"FE",X"F2",X"38",X"F3",X"1A",X"F4",X"04",X"F5",X"EB",X"F5",
		X"CA",X"F6",X"A3",X"F7",X"78",X"F8",X"45",X"F9",X"0E",X"FA",X"D1",X"FA",X"8D",X"FB",X"42",X"FC",
		X"F8",X"FC",X"A3",X"FD",X"4B",X"FE",X"ED",X"FE",X"8B",X"FF",X"24",X"00",X"B8",X"00",X"49",X"01",
		X"D4",X"01",X"5B",X"02",X"E1",X"02",X"60",X"03",X"DD",X"03",X"54",X"04",X"CA",X"04",X"3A",X"05",
		X"A6",X"05",X"10",X"06",X"78",X"06",X"DB",X"06",X"3E",X"07",X"9A",X"07",X"F4",X"07",X"4D",X"08",
		X"A3",X"08",X"F4",X"08",X"45",X"09",X"93",X"09",X"DD",X"09",X"26",X"0A",X"6D",X"0A",X"B0",X"0A",
		X"F1",X"0A",X"34",X"0B",X"5A",X"0B",X"2D",X"0B",X"C6",X"0A",X"3A",X"0A",X"94",X"09",X"E1",X"08",
		X"24",X"08",X"64",X"07",X"A3",X"06",X"E5",X"05",X"27",X"05",X"6D",X"04",X"B8",X"03",X"07",X"03",
		X"59",X"02",X"B1",X"01",X"0C",X"01",X"6D",X"00",X"D3",X"FF",X"3E",X"FF",X"AC",X"FE",X"1E",X"FE",
		X"95",X"FD",X"0F",X"FD",X"8F",X"FC",X"10",X"FC",X"96",X"FB",X"20",X"FB",X"E9",X"FA",X"FE",X"FA",
		X"45",X"FB",X"AB",X"FB",X"28",X"FC",X"B2",X"FC",X"44",X"FD",X"D5",X"FD",X"6C",X"FE",X"00",X"FF",
		X"96",X"FF",X"23",X"00",X"B2",X"00",X"39",X"01",X"C4",X"01",X"43",X"02",X"C8",X"02",X"3E",X"03",
		X"BB",X"03",X"2C",X"04",X"A2",X"04",X"0A",X"05",X"7A",X"05",X"DD",X"05",X"45",X"06",X"A3",X"06",
		X"05",X"07",X"4D",X"07",X"49",X"07",X"02",X"07",X"95",X"06",X"0C",X"06",X"76",X"05",X"D0",X"04",
		X"2B",X"04",X"7F",X"03",X"D8",X"02",X"2E",X"02",X"8C",X"01",X"E9",X"00",X"4B",X"00",X"B1",X"FF",
		X"1C",X"FF",X"8B",X"FE",X"FC",X"FD",X"73",X"FD",X"ED",X"FC",X"6C",X"FC",X"EE",X"FB",X"74",X"FB",
		X"FD",X"FA",X"8B",X"FA",X"1A",X"FA",X"AF",X"F9",X"45",X"F9",X"E1",X"F8",X"7E",X"F8",X"20",X"F8",
		X"C0",X"F7",X"6A",X"F7",X"11",X"F7",X"BF",X"F6",X"6A",X"F6",X"1D",X"F6",X"CF",X"F5",X"86",X"F5",
		X"3D",X"F5",X"F9",X"F4",X"B7",X"F4",X"74",X"F4",X"35",X"F4",X"F9",X"F3",X"BE",X"F3",X"83",X"F3",
		X"4F",X"F3",X"18",X"F3",X"E7",X"F2",X"D6",X"F2",X"E6",X"F2",X"E4",X"F2",X"F4",X"F2",X"EF",X"F2",
		X"02",X"F3",X"FA",X"F2",X"10",X"F3",X"05",X"F3",X"1D",X"F3",X"11",X"F3",X"2D",X"F3",X"1D",X"F3",
		X"39",X"F3",X"2A",X"F3",X"48",X"F3",X"35",X"F3",X"56",X"F3",X"42",X"F3",X"64",X"F3",X"4D",X"F3",
		X"71",X"F3",X"5A",X"F3",X"7D",X"F3",X"67",X"F3",X"8A",X"F3",X"71",X"F3",X"96",X"F3",X"80",X"F3",
		X"A1",X"F3",X"8C",X"F3",X"AD",X"F3",X"99",X"F3",X"B8",X"F3",X"A9",X"F3",X"C1",X"F3",X"B6",X"F3",
		X"CC",X"F3",X"C5",X"F3",X"D6",X"F3",X"D6",X"F3",X"DD",X"F3",X"E4",X"F3",X"E7",X"F3",X"F7",X"F3",
		X"EB",X"F3",X"09",X"F4",X"F3",X"F3",X"19",X"F4",X"F7",X"F3",X"2E",X"F4",X"FC",X"F3",X"40",X"F4",
		X"FF",X"F3",X"57",X"F4",X"02",X"F4",X"6B",X"F4",X"04",X"F4",X"81",X"F4",X"04",X"F4",X"9A",X"F4",
		X"05",X"F4",X"B1",X"F4",X"03",X"F4",X"CA",X"F4",X"02",X"F4",X"E2",X"F4",X"00",X"F4",X"F9",X"F4",
		X"40",X"F4",X"5A",X"F6",X"06",X"F6",X"35",X"F8",X"B2",X"F7",X"FE",X"F9",X"47",X"F9",X"B2",X"FB",
		X"C1",X"FA",X"55",X"FD",X"22",X"FC",X"E3",X"FE",X"68",X"FD",X"65",X"00",X"90",X"FE",X"DA",X"01",
		X"96",X"FF",X"52",X"03",X"6B",X"00",X"ED",X"04",X"C7",X"00",X"7E",X"07",X"2F",X"F8",X"9C",X"FA",
		X"9C",X"15",X"24",X"0A",X"51",X"ED",X"7A",X"09",X"2F",X"02",X"BD",X"F0",X"52",X"0C",X"AB",X"16",
		X"A1",X"0D",X"48",X"FD",X"DC",X"09",X"6C",X"FD",X"23",X"0C",X"47",X"EF",X"B5",X"F9",X"49",X"11",
		X"6A",X"0F",X"C4",X"EF",X"37",X"F9",X"1C",X"EE",X"DF",X"09",X"24",X"00",X"18",X"06",X"96",X"17",
		X"8B",X"10",X"6A",X"14",X"04",X"13",X"A1",X"0D",X"12",X"F8",X"24",X"1A",X"D3",X"02",X"A9",X"F3",
		X"8E",X"F3",X"4B",X"F9",X"37",X"18",X"AD",X"03",X"58",X"01",X"F4",X"07",X"BB",X"ED",X"FB",X"F7",
		X"96",X"07",X"38",X"00",X"5B",X"09",X"F1",X"16",X"63",X"EB",X"59",X"03",X"91",X"0D",X"EE",X"1A",
		X"BC",X"FB",X"2A",X"09",X"34",X"0B",X"84",X"FC",X"3E",X"0C",X"2A",X"EC",X"CA",X"08",X"4E",X"02",
		X"57",X"EF",X"D4",X"F7",X"23",X"09",X"08",X"FD",X"55",X"EC",X"9C",X"01",X"08",X"05",X"95",X"01",
		X"F4",X"05",X"09",X"FF",X"B4",X"18",X"72",X"0E",X"C7",X"16",X"74",X"06",X"07",X"F0",X"7E",X"04",
		X"3A",X"16",X"AA",X"0F",X"1D",X"15",X"C4",X"F6",X"BF",X"11",X"A2",X"0C",X"83",X"FA",X"55",X"12",
		X"13",X"15",X"F2",X"02",X"FE",X"00",X"3F",X"07",X"A3",X"EA",X"45",X"10",X"DE",X"F7",X"8A",X"F2",
		X"CE",X"01",X"2C",X"19",X"38",X"F9",X"83",X"F4",X"9C",X"0A",X"3E",X"FC",X"0A",X"0D",X"25",X"17",
		X"F3",X"06",X"7C",X"F4",X"9C",X"F0",X"2E",X"04",X"4B",X"14",X"F8",X"11",X"84",X"FC",X"DD",X"EF",
		X"3E",X"F7",X"C5",X"EE",X"54",X"0A",X"94",X"FD",X"A0",X"07",X"28",X"FE",X"5A",X"08",X"7D",X"FB",
		X"E4",X"11",X"8A",X"0A",X"28",X"F8",X"A1",X"1B",X"D7",X"FC",X"67",X"F5",X"FC",X"EF",X"46",X"0D",
		X"84",X"10",X"9B",X"FA",X"89",X"0A",X"45",X"F6",X"A6",X"F0",X"2D",X"0D",X"0C",X"12",X"BD",X"12",
		X"62",X"10",X"46",X"14",X"3C",X"09",X"D9",X"EF",X"7B",X"00",X"D3",X"15",X"A9",X"0E",X"86",X"14",
		X"D6",X"0E",X"DC",X"13",X"91",X"F4",X"04",X"14",X"48",X"09",X"25",X"F5",X"6E",X"F0",X"EA",X"0F",
		X"DF",X"F1",X"98",X"FB",X"8E",X"07",X"82",X"FC",X"7D",X"11",X"21",X"15",X"40",X"FE",X"8E",X"04",
		X"4D",X"01",X"92",X"ED",X"C1",X"0F",X"38",X"0F",X"78",X"F4",X"26",X"F3",X"AD",X"F2",X"88",X"F4",
		X"CB",X"09",X"7A",X"FC",X"98",X"07",X"17",X"FD",X"27",X"08",X"7D",X"FA",X"EA",X"16",X"5B",X"0D",
		X"9F",X"15",X"B5",X"FA",X"DE",X"F1",X"FD",X"F3",X"D3",X"0E",X"2E",X"0F",X"BD",X"F0",X"EB",X"FA",
		X"12",X"15",X"75",X"04",X"48",X"EF",X"8C",X"F8",X"8D",X"12",X"AD",X"08",X"FF",X"F7",X"7C",X"1B",
		X"64",X"F9",X"53",X"08",X"BD",X"FC",X"46",X"07",X"4E",X"FC",X"C3",X"0A",X"DD",X"11",X"ED",X"ED",
		X"A3",X"FD",X"15",X"11",X"E4",X"11",X"FD",X"0F",X"12",X"12",X"60",X"10",X"CE",X"0B",X"77",X"EA",
		X"C7",X"06",X"92",X"FF",X"DF",X"01",X"44",X"16",X"85",X"F7",X"82",X"F2",X"D8",X"0E",X"FB",X"10",
		X"E8",X"10",X"57",X"11",X"BF",X"08",X"9D",X"EC",X"7D",X"F8",X"5F",X"EB",X"D5",X"00",X"56",X"02",
		X"4F",X"01",X"2D",X"02",X"06",X"01",X"92",X"03",X"1C",X"EC",X"D3",X"0C",X"A3",X"10",X"B4",X"F5",
		X"93",X"12",X"67",X"07",X"95",X"FC",X"0D",X"07",X"88",X"FA",X"FD",X"16",X"65",X"0C",X"0B",X"14",
		X"24",X"0D",X"13",X"15",X"24",X"00",X"7D",X"FE",X"D9",X"17",X"50",X"F7",X"98",X"F3",X"00",X"F0",
		X"EB",X"F5",X"4E",X"ED",X"E9",X"FD",X"F4",X"04",X"CC",X"FC",X"69",X"11",X"76",X"13",X"83",X"FB",
		X"45",X"06",X"0B",X"FC",X"74",X"09",X"EC",X"05",X"4E",X"FA",X"2C",X"1B",X"EB",X"F3",X"15",X"0C",
		X"2D",X"F7",X"96",X"0D",X"89",X"10",X"65",X"10",X"9B",X"10",X"80",X"08",X"50",X"EA",X"4E",X"07",
		X"CA",X"FD",X"A8",X"02",X"86",X"15",X"F0",X"F3",X"BD",X"F4",X"9A",X"0D",X"69",X"12",X"FC",X"FA",
		X"59",X"EF",X"D5",X"0C",X"85",X"F3",X"51",X"F6",X"AF",X"0F",X"35",X"12",X"6E",X"04",X"29",X"FA",
		X"35",X"18",X"15",X"FA",X"3E",X"F2",X"2B",X"F1",X"99",X"0A",X"72",X"F8",X"5E",X"0A",X"57",X"F2",
		X"7A",X"F2",X"B9",X"F1",X"66",X"F3",X"A8",X"0D",X"69",X"10",X"01",X"11",X"7F",X"08",X"00",X"EF",
		X"3D",X"F3",X"BE",X"FD",X"9B",X"18",X"66",X"F5",X"B6",X"0A",X"A2",X"F6",X"2E",X"F4",X"6A",X"0A",
		X"0E",X"F7",X"96",X"12",X"EC",X"F7",X"62",X"08",X"C1",X"F9",X"AB",X"09",X"07",X"F1",X"7B",X"FA",
		X"FE",X"0A",X"54",X"E8",X"C7",X"08",X"FE",X"FC",X"23",X"F1",X"57",X"F1",X"25",X"F4",X"E4",X"EE",
		X"CB",X"F9",X"E9",X"06",X"31",X"FB",X"D2",X"08",X"66",X"EE",X"AC",X"11",X"15",X"0A",X"6F",X"F3",
		X"91",X"EF",X"81",X"FE",X"4C",X"07",X"54",X"EB",X"05",X"F8",X"33",X"EC",X"1E",X"0E",X"47",X"F4",
		X"AE",X"F6",X"C7",X"08",X"AE",X"F5",X"5A",X"ED",X"C2",X"00",X"9A",X"04",X"97",X"EF",X"3C",X"F3",
		X"8A",X"F2",X"BE",X"F1",X"BC",X"F3",X"B5",X"F0",X"22",X"F5",X"6A",X"EE",X"58",X"0A",X"C7",X"F9",
		X"6E",X"F2",X"D3",X"0A",X"45",X"F9",X"F1",X"09",X"C1",X"F6",X"90",X"17",X"B8",X"FE",X"BC",X"00",
		X"B2",X"0F",X"5E",X"F3",X"CE",X"18",X"78",X"FE",X"81",X"01",X"13",X"04",X"C7",X"EB",X"A8",X"0A",
		X"7F",X"FA",X"73",X"EF",X"49",X"F6",X"24",X"0E",X"03",X"11",X"46",X"10",X"9E",X"08",X"F9",X"EA",
		X"74",X"06",X"DC",X"FF",X"43",X"EF",X"70",X"F3",X"F7",X"F9",X"99",X"18",X"FF",X"F9",X"16",X"06",
		X"8B",X"FD",X"A8",X"04",X"06",X"16",X"FB",X"08",X"46",X"FB",X"B0",X"07",X"A0",X"F8",X"38",X"14",
		X"22",X"0C",X"26",X"15",X"60",X"FA",X"89",X"05",X"C8",X"FD",X"20",X"EC",X"E5",X"01",X"F8",X"11",
		X"91",X"0E",X"20",X"11",X"01",X"0E",X"59",X"FA",X"FE",X"05",X"A7",X"FC",X"04",X"05",X"D1",X"FC",
		X"B5",X"05",X"4D",X"FA",X"FD",X"15",X"34",X"0B",X"FC",X"13",X"DB",X"F6",X"0E",X"F2",X"54",X"F1",
		X"85",X"F3",X"8F",X"EF",X"4A",X"08",X"69",X"FB",X"0C",X"06",X"38",X"FB",X"BA",X"0A",X"89",X"13",
		X"8F",X"0B",X"EB",X"14",X"C2",X"FF",X"1C",X"F2",X"A2",X"EF",X"0C",X"07",X"45",X"11",X"3A",X"F7",
		X"85",X"EF",X"C4",X"F4",X"77",X"EE",X"EE",X"08",X"FE",X"0F",X"14",X"F8",X"DA",X"0A",X"F4",X"0F",
		X"C9",X"EB",X"17",X"FF",X"72",X"0C",X"CD",X"15",X"1A",X"FA",X"EC",X"05",X"E7",X"FB",X"EC",X"05",
		X"4D",X"11",X"FB",X"F5",X"C7",X"0C",X"A5",X"12",X"12",X"F8",X"7F",X"08",X"45",X"0F",X"24",X"F7",
		X"79",X"09",X"E9",X"F2",X"37",X"EF",X"AC",X"FD",X"3F",X"10",X"B9",X"11",X"65",X"FB",X"48",X"04",
		X"2E",X"FD",X"3D",X"04",X"F3",X"FB",X"16",X"09",X"5D",X"14",X"07",X"05",X"A0",X"F1",X"32",X"F1",
		X"2C",X"F4",X"D3",X"0F",X"BB",X"08",X"06",X"F6",X"09",X"17",X"C4",X"FC",X"60",X"00",X"17",X"12",
		X"5E",X"0E",X"1C",X"FA",X"3F",X"EE",X"6F",X"F4",X"62",X"EF",X"35",X"F4",X"60",X"EF",X"85",X"F4",
		X"A8",X"EF",X"9E",X"11",X"FD",X"06",X"7D",X"FA",X"8F",X"0D",X"D9",X"13",X"7A",X"FD",X"FF",X"01",
		X"A2",X"FF",X"97",X"00",X"38",X"15",X"9A",X"F3",X"98",X"0B",X"C1",X"F4",X"20",X"12",X"53",X"06",
		X"25",X"EF",X"0D",X"FD",X"91",X"14",X"94",X"06",X"6A",X"F9",X"35",X"0F",X"AA",X"10",X"66",X"02",
		X"A8",X"ED",X"A5",X"F4",X"82",X"EE",X"50",X"0A",X"32",X"0E",X"CE",X"F6",X"71",X"0C",X"DE",X"10",
		X"4E",X"0C",X"55",X"13",X"AE",X"FE",X"86",X"FF",X"01",X"03",X"75",X"EA",X"74",X"F7",X"F1",X"EA",
		X"CF",X"03",X"B4",X"00",X"20",X"ED",X"0E",X"07",X"58",X"11",X"C6",X"0C",X"69",X"11",X"14",X"09",
		X"6C",X"F3",X"35",X"EE",X"29",X"FE",X"67",X"05",X"52",X"EC",X"83",X"F5",X"8E",X"ED",X"D1",X"FB",
		X"38",X"11",X"45",X"03",X"B7",X"EA",X"60",X"08",X"09",X"FB",X"96",X"EF",X"BA",X"0A",X"4C",X"11",
		X"70",X"09",X"F6",X"F2",X"29",X"EF",X"31",X"FC",X"3E",X"12",X"1C",X"01",X"C3",X"EA",X"F0",X"0A",
		X"D3",X"F5",X"D0",X"FD",X"92",X"03",X"1C",X"FB",X"49",X"17",X"D5",X"F5",X"C0",X"F2",X"AC",X"07",
		X"94",X"F9",X"E4",X"07",X"BA",X"F2",X"59",X"F0",X"22",X"FA",X"D5",X"15",X"B2",X"FA",X"5E",X"03",
		X"A3",X"FE",X"08",X"ED",X"DB",X"0B",X"87",X"10",X"BE",X"FF",X"AA",X"ED",X"67",X"F4",X"9B",X"EF",
		X"6A",X"0C",X"F3",X"0C",X"FF",X"F1",X"59",X"F2",X"A6",X"F0",X"AE",X"F3",X"1B",X"EE",X"6F",X"03",
		X"94",X"00",X"67",X"EC",X"24",X"0A",X"1E",X"10",X"3D",X"0C",X"35",X"F4",X"04",X"EF",X"29",X"08",
		X"AB",X"F9",X"A0",X"EF",X"13",X"F2",X"1E",X"F6",X"A0",X"0A",X"F7",X"EE",X"02",X"F3",X"0C",X"FB",
		X"3A",X"17",X"E6",X"F7",X"B1",X"05",X"D8",X"10",X"53",X"F7",X"4B",X"08",X"CB",X"F5",X"26",X"EE",
		X"ED",X"08",X"90",X"F9",X"20",X"07",X"8E",X"F8",X"A0",X"0D",X"A0",X"09",X"3B",X"F5",X"14",X"17",
		X"8A",X"FC",X"B8",X"FF",X"BA",X"13",X"B1",X"F8",X"A5",X"05",X"8B",X"12",X"01",X"0C",X"CF",X"10",
		X"7F",X"0D",X"20",X"0A",X"50",X"EC",X"66",X"0E",X"EF",X"EF",X"63",X"F8",X"24",X"0D",X"F1",X"0A",
		X"2C",X"E8",X"A0",X"06",X"EF",X"FB",X"9C",X"02",X"7E",X"10",X"A8",X"0E",X"4E",X"F6",X"4F",X"0A",
		X"2C",X"F1",X"05",X"F8",X"8B",X"0E",X"D9",X"0F",X"0D",X"0B",X"0A",X"F9",X"67",X"06",X"9B",X"F8",
		X"45",X"0F",X"BB",X"0E",X"43",X"0D",X"E7",X"10",X"4F",X"FC",X"53",X"EE",X"25",X"08",X"E1",X"F9",
		X"1A",X"05",X"E5",X"FA",X"65",X"05",X"B3",X"F8",X"B3",X"10",X"2A",X"0D",X"C6",X"0E",X"90",X"0E",
		X"4B",X"09",X"9A",X"ED",X"3E",X"F5",X"C8",X"EB",X"AA",X"05",X"D5",X"FB",X"4D",X"03",X"3F",X"FC",
		X"C2",X"04",X"51",X"13",X"23",X"0A",X"53",X"12",X"B4",X"04",X"CF",X"EF",X"CE",X"F2",X"59",X"EE",
		X"23",X"04",X"62",X"0A",X"A9",X"EE",X"63",X"F1",X"02",X"FD",X"15",X"12",X"23",X"0D",X"6A",X"FB",
		X"FE",X"02",X"96",X"FB",X"02",X"EB",X"30",X"F9",X"4E",X"0C",X"DC",X"09",X"41",X"EB",X"FE",X"F6",
		X"CD",X"EA",X"82",X"07",X"64",X"FB",X"1D",X"EE",X"B8",X"FB",X"8A",X"13",X"16",X"FD",X"8C",X"EE",
		X"B6",X"05",X"64",X"11",X"93",X"0A",X"7D",X"F8",X"35",X"07",X"61",X"F6",X"8F",X"12",X"15",X"01",
		X"34",X"FB",X"CE",X"12",X"34",X"0B",X"FB",X"0F",X"F5",X"0C",X"74",X"F6",X"EF",X"F9",X"61",X"16",
		X"6A",X"F7",X"E9",X"F1",X"07",X"05",X"B6",X"12",X"51",X"ED",X"F1",X"FA",X"20",X"03",X"39",X"FB",
		X"D9",X"0C",X"75",X"12",X"85",X"FA",X"37",X"03",X"39",X"FC",X"0B",X"03",X"7B",X"FB",X"EB",X"05",
		X"81",X"13",X"A5",X"F9",X"37",X"EF",X"0D",X"08",X"6E",X"0F",X"75",X"0D",X"D5",X"0A",X"62",X"EF",
		X"E5",X"F2",X"C9",X"EE",X"F0",X"FC",X"C0",X"13",X"C2",X"F8",X"D9",X"03",X"F7",X"FB",X"25",X"EC",
		X"5B",X"F5",X"86",X"EC",X"A2",X"05",X"BC",X"0E",X"EF",X"0D",X"64",X"0D",X"52",X"0E",X"27",X"0D",
		X"2E",X"0E",X"DB",X"0D",X"2B",X"06",X"32",X"E9",X"05",X"06",X"07",X"FB",X"BC",X"02",X"48",X"FC",
		X"41",X"EC",X"CE",X"0F",X"E3",X"06",X"EF",X"F7",X"C3",X"0D",X"07",X"0E",X"E5",X"F3",X"48",X"F3",
		X"DC",X"09",X"47",X"EF",X"DD",X"F2",X"31",X"EF",X"89",X"F3",X"4C",X"ED",X"27",X"05",X"6C",X"FC",
		X"25",X"ED",X"8A",X"0B",X"71",X"0D",X"3A",X"0E",X"18",X"0D",X"2C",X"0E",X"31",X"0D",X"E4",X"0C",
		X"38",X"F4",X"6D",X"0E",X"04",X"0B",X"0C",X"12",X"B3",X"FE",X"43",X"FE",X"FC",X"00",X"00",X"FC",
		X"F1",X"14",X"A0",X"07",X"AC",X"FB",X"56",X"02",X"92",X"F8",X"A1",X"E9",X"D7",X"FD",X"4C",X"0A",
		X"DE",X"11",X"BB",X"07",X"DB",X"14",X"04",X"FF",X"87",X"FF",X"31",X"FE",X"17",X"00",X"B3",X"FD",
		X"7B",X"00",X"9D",X"FD",X"90",X"EC",X"83",X"F2",X"BD",X"F2",X"7E",X"08",X"8C",X"F5",X"1B",X"0F",
		X"E9",X"0D",X"75",X"01",X"2B",X"F9",X"54",X"16",X"40",X"00",X"5E",X"FB",X"F6",X"0C",X"95",X"0F",
		X"E5",X"FD",X"CE",X"EC",X"7C",X"05",X"56",X"0F",X"D3",X"0B",X"CB",X"0C",X"5B",X"EF",X"5F",X"F3",
		X"C0",X"EC",X"E8",X"FC",X"20",X"0D",X"FE",X"0F",X"31",X"FA",X"73",X"F5",X"60",X"09",X"10",X"E9",
		X"78",X"02",X"B2",X"FF",X"9C",X"EB",X"BB",X"06",X"00",X"0E",X"46",X"F5",X"5E",X"EE",X"CC",X"F5",
		X"C3",X"0C",X"86",X"0D",X"D1",X"0C",X"21",X"0D",X"3A",X"0E",X"BC",X"FC",X"59",X"FD",X"07",X"17",
		X"09",X"FA",X"40",X"01",X"60",X"FE",X"72",X"EE",X"EB",X"F0",X"D3",X"F1",X"AD",X"05",X"2F",X"F9",
		X"1F",X"07",X"DC",X"13",X"43",X"FE",X"00",X"FF",X"A0",X"FE",X"E6",X"FE",X"D2",X"FE",X"2A",X"FE",
		X"7C",X"13",X"E5",X"07",X"87",X"12",X"D6",X"F9",X"C8",X"FF",X"09",X"12",X"AF",X"F3",X"6A",X"09",
		X"1A",X"0B",X"32",X"F1",X"7C",X"F0",X"26",X"F0",X"2F",X"F8",X"11",X"14",X"43",X"F9",X"7F",X"00",
		X"57",X"10",X"B9",X"F6",X"4B",X"EE",X"C4",X"F2",X"59",X"EE",X"7F",X"F3",X"21",X"ED",X"06",X"0A",
		X"62",X"0A",X"F3",X"F5",X"23",X"EB",X"96",X"FC",X"B1",X"00",X"16",X"FD",X"B0",X"00",X"91",X"FC",
		X"70",X"02",X"A4",X"E8",X"2B",X"0B",X"CB",X"F4",X"BB",X"08",X"AD",X"F1",X"6E",X"F1",X"9C",X"EF",
		X"84",X"07",X"DF",X"0D",X"39",X"F1",X"9C",X"F4",X"D0",X"0E",X"AE",X"05",X"46",X"EC",X"AD",X"FE",
		X"5F",X"0F",X"8F",X"0B",X"AD",X"0E",X"F7",X"F6",X"9A",X"EF",X"99",X"0B",X"B8",X"0C",X"64",X"0D",
		X"69",X"0C",X"54",X"0D",X"9E",X"0C",X"52",X"0B",X"82",X"EF",X"74",X"F6",X"19",X"10",X"28",X"01",
		X"33",X"F8",X"85",X"15",X"52",X"F5",X"6C",X"05",X"BE",X"F8",X"B0",X"ED",X"A7",X"F4",X"29",X"07",
		X"E5",X"F4",X"15",X"10",X"86",X"09",X"86",X"10",X"8C",X"06",X"70",X"F5",X"7E",X"EA",X"02",X"FF",
		X"DC",X"FE",X"11",X"FE",X"B6",X"FF",X"4C",X"FC",X"B6",X"13",X"4F",X"F3",X"49",X"08",X"CB",X"0E",
		X"53",X"07",X"64",X"F6",X"84",X"08",X"1B",X"EA",X"D9",X"FF",X"A1",X"0A",X"03",X"F4",X"8F",X"0F",
		X"8C",X"03",X"AF",X"EE",X"A6",X"F1",X"EE",X"EF",X"6B",X"F1",X"AB",X"EF",X"0C",X"06",X"AD",X"0F",
		X"3D",X"08",X"72",X"F6",X"9D",X"0B",X"93",X"0E",X"32",X"03",X"3B",X"ED",X"5C",X"F3",X"5E",X"ED",
		X"72",X"F9",X"E4",X"05",X"06",X"ED",X"A5",X"F3",X"4E",X"ED",X"44",X"03",X"D2",X"0E",X"AE",X"0B",
		X"EF",X"0C",X"CC",X"F1",X"DA",X"F1",X"1F",X"EE",X"93",X"FA",X"29",X"05",X"F1",X"EC",X"41",X"F2",
		X"2A",X"FE",X"E7",X"13",X"7D",X"00",X"B1",X"F1",X"1C",X"EF",X"3E",X"F3",X"97",X"ED",X"68",X"06",
		X"62",X"0D",X"EB",X"F5",X"86",X"ED",X"CB",X"F7",X"51",X"06",X"58",X"F0",X"AC",X"F0",X"46",X"F2",
		X"2F",X"EE",X"95",X"03",X"26",X"FD",X"34",X"EC",X"27",X"F5",X"69",X"EC",X"C2",X"02",X"C7",X"0D",
		X"11",X"0E",X"66",X"F6",X"71",X"F1",X"68",X"08",X"32",X"F6",X"9D",X"09",X"A6",X"EB",X"E8",X"FE",
		X"DE",X"02",X"B0",X"EC",X"AB",X"F4",X"65",X"ED",X"74",X"09",X"67",X"F4",X"7D",X"FC",X"88",X"11",
		X"F4",X"09",X"43",X"10",X"D3",X"F4",X"DA",X"F2",X"39",X"07",X"B1",X"F7",X"3F",X"07",X"B3",X"F4",
		X"19",X"15",X"B2",X"FA",X"E1",X"00",X"AE",X"FF",X"91",X"EB",X"72",X"09",X"19",X"0C",X"F1",X"F5",
		X"0E",X"0B",X"BC",X"0D",X"8C",X"0C",X"0F",X"0D",X"55",X"0D",X"FA",X"09",X"72",X"F5",X"13",X"0A",
		X"DC",X"EA",X"F3",X"FE",X"AF",X"0B",X"C9",X"10",X"68",X"F8",X"ED",X"03",X"4B",X"FA",X"CD",X"03",
		X"42",X"F9",X"82",X"06",X"7F",X"F0",X"32",X"05",X"AA",X"F9",X"87",X"05",X"29",X"10",X"19",X"0B",
		X"7B",X"09",X"9D",X"EC",X"D3",X"F4",X"B3",X"EC",X"13",X"01",X"1A",X"10",X"52",X"F8",X"BD",X"03",
		X"6E",X"F9",X"12",X"EE",X"2A",X"10",X"E4",X"08",X"A8",X"10",X"BF",X"08",X"1B",X"10",X"66",X"ED",
		X"94",X"F9",X"02",X"08",X"9F",X"13",X"5F",X"FB",X"26",X"01",X"C1",X"FC",X"87",X"00",X"83",X"FD",
		X"2B",X"EC",X"41",X"0B",X"5D",X"0A",X"F0",X"F3",X"27",X"10",X"D3",X"01",X"CD",X"F9",X"D3",X"0D",
		X"56",X"F2",X"24",X"EF",X"F8",X"F7",X"9E",X"0C",X"36",X"0F",X"E5",X"FD",X"DB",X"FC",X"C2",X"10",
		X"D4",X"0A",X"E5",X"F8",X"DD",X"04",X"C1",X"0E",X"EB",X"ED",X"8C",X"F4",X"12",X"EC",X"1C",X"FE",
		X"A8",X"02",X"42",X"EC",X"41",X"F7",X"9F",X"0C",X"EB",X"06",X"F8",X"E9",X"B4",X"02",X"11",X"FE",
		X"F5",X"EE",X"B4",X"F0",X"A4",X"06",X"97",X"F6",X"88",X"EF",X"EC",X"F0",X"DA",X"F5",X"73",X"0F",
		X"F6",X"03",X"CE",X"EA",X"2D",X"04",X"96",X"FB",X"EA",X"F5",X"4A",X"07",X"C2",X"F4",X"68",X"16",
		X"25",X"F7",X"C8",X"02",X"75",X"0E",X"12",X"0C",X"D1",X"0B",X"09",X"F5",X"86",X"09",X"38",X"ED",
		X"1A",X"FC",X"B7",X"03",X"AB",X"EE",X"CE",X"F0",X"61",X"00",X"A4",X"10",X"98",X"09",X"1E",X"10",
		X"01",X"FF",X"49",X"EE",X"EE",X"F2",X"5C",X"EF",X"E8",X"F2",X"FA",X"EF",X"C7",X"0B",X"26",X"ED",
		X"43",X"FC",X"F8",X"00",X"35",X"FD",X"80",X"00",X"7A",X"FD",X"6A",X"00",X"50",X"FD",X"EF",X"00",
		X"F5",X"E5",X"1A",X"07",X"77",X"F9",X"24",X"03",X"DB",X"FB",X"80",X"ED",X"A3",X"F3",X"C7",X"F0",
		X"19",X"10",X"6E",X"03",X"E9",X"F9",X"6B",X"06",X"C5",X"EA",X"60",X"02",X"C3",X"0D",X"04",X"0D",
		X"B4",X"F8",X"22",X"04",X"64",X"13",X"4B",X"F8",X"85",X"03",X"28",X"FB",X"C8",X"02",X"99",X"11",
		X"FF",X"06",X"92",X"F4",X"D9",X"ED",X"53",X"FA",X"1A",X"0E",X"F2",X"0B",X"1C",X"0D",X"EA",X"0B",
		X"BA",X"0D",X"68",X"F7",X"D1",X"EF",X"36",X"0A",X"D6",X"EF",X"EE",X"02",X"E7",X"0E",X"07",X"0B",
		X"D2",X"F5",X"87",X"F0",X"AF",X"0F",X"C1",X"03",X"DB",X"F7",X"89",X"10",X"0C",X"00",X"7A",X"EC",
		X"80",X"03",X"FE",X"0D",X"FC",X"0B",X"D1",X"0B",X"A3",X"F3",X"F2",X"EF",X"48",X"F2",X"84",X"EF",
		X"79",X"07",X"C7",X"F6",X"9A",X"09",X"8A",X"0A",X"96",X"ED",X"71",X"FA",X"DD",X"0D",X"FE",X"0B",
		X"4D",X"0C",X"79",X"0D",X"EF",X"F9",X"0D",X"EE",X"CB",X"09",X"1F",X"0D",X"A2",X"08",X"65",X"F4",
		X"17",X"10",X"9E",X"08",X"6A",X"F8",X"08",X"EB",X"E4",X"FA",X"22",X"02",X"DB",X"F9",X"E7",X"0C",
		X"22",X"0E",X"D7",X"FD",X"06",X"ED",X"6C",X"05",X"00",X"FA",X"51",X"ED",X"D1",X"0C",X"6E",X"EC",
		X"2D",X"FC",X"2A",X"01",X"0F",X"FB",X"EC",X"0B",X"00",X"F6",X"AE",X"09",X"32",X"10",X"AD",X"00",
		X"7D",X"FA",X"6A",X"0E",X"D1",X"0C",X"2D",X"FC",X"39",X"ED",X"4C",X"07",X"E8",X"F7",X"CD",X"04",
		X"AD",X"F7",X"E1",X"0A",X"79",X"0D",X"C0",X"0A",X"ED",X"0D",X"85",X"08",X"4C",X"F1",X"03",X"F6",
		X"9A",X"09",X"75",X"E7",X"1E",X"05",X"60",X"FA",X"C1",X"00",X"FB",X"0E",X"E6",X"F6",X"06",X"EE",
		X"28",X"F4",X"E7",X"EC",X"CF",X"F9",X"F6",X"09",X"8A",X"10",X"94",X"FD",X"77",X"F1",X"21",X"EE",
		X"CE",X"F9",X"6B",X"0A",X"F5",X"10",X"D0",X"FA",X"0F",X"01",X"95",X"FC",X"36",X"00",X"6A",X"10",
		X"AE",X"F3",X"25",X"08",X"2A",X"F2",X"C2",X"EF",X"02",X"F8",X"F0",X"0F",X"73",X"00",X"C3",X"EB",
		X"C4",X"04",X"FA",X"FA",X"A1",X"EE",X"24",X"F1",X"04",X"FC",X"F9",X"10",X"A5",X"08",X"BC",X"0F",
		X"5F",X"F4",X"63",X"F2",X"36",X"09",X"FD",X"0D",X"44",X"0A",X"55",X"0E",X"2F",X"09",X"B1",X"10",
		X"2D",X"FA",X"10",X"00",X"88",X"0E",X"B4",X"0B",X"D5",X"F3",X"AD",X"FC",X"E7",X"02",X"86",X"E8",
		X"C0",X"09",X"14",X"F5",X"C1",X"F1",X"1F",X"0A",X"59",X"09",X"BD",X"F2",X"F3",X"12",X"F4",X"FC",
		X"5F",X"FC",X"8D",X"0F",X"B2",X"FB",X"FD",X"EC",X"94",X"F4",X"69",X"ED",X"79",X"0F",X"80",X"F8",
		X"E8",X"02",X"CF",X"FA",X"0E",X"EE",X"39",X"F3",X"F5",X"09",X"E0",X"0B",X"BD",X"0D",X"D0",X"03",
		X"7D",X"EF",X"62",X"F0",X"E8",X"FD",X"09",X"11",X"6E",X"F7",X"BD",X"EF",X"59",X"08",X"87",X"0B",
		X"AF",X"F0",X"46",X"F2",X"5E",X"EF",X"36",X"07",X"7F",X"F6",X"3C",X"09",X"42",X"0C",X"B3",X"0D",
		X"BB",X"02",X"C0",X"F8",X"AD",X"06",X"26",X"E7",X"97",X"08",X"6D",X"F7",X"5F",X"F1",X"02",X"05",
		X"88",X"F9",X"5A",X"03",X"A2",X"F8",X"4B",X"0B",X"AC",X"0D",X"71",X"08",X"0F",X"F8",X"4F",X"04",
		X"13",X"F8",X"E8",X"06",X"1C",X"EB",X"E7",X"FF",X"6E",X"0C",X"8E",X"0D",X"47",X"F8",X"6C",X"03",
		X"74",X"0E",X"5D",X"F2",X"8B",X"0D",X"81",X"05",X"51",X"F0",X"6B",X"F1",X"77",X"F0",X"8A",X"F3",
		X"1A",X"0C",X"86",X"07",X"F3",X"EB",X"EC",X"FE",X"EC",X"00",X"57",X"EE",X"24",X"F1",X"A1",X"03",
		X"53",X"FA",X"F5",X"ED",X"77",X"0C",X"12",X"0B",X"1A",X"09",X"1B",X"EC",X"F8",X"FC",X"D1",X"0B",
		X"7D",X"F2",X"F8",X"F0",X"24",X"F1",X"97",X"F1",X"89",X"F0",X"AE",X"F2",X"71",X"EE",X"F4",X"03",
		X"C3",X"FB",X"94",X"ED",X"BB",X"0A",X"1F",X"0A",X"97",X"F1",X"73",X"F2",X"B9",X"EE",X"CF",X"FC",
		X"B7",X"03",X"3D",X"EC",X"65",X"F5",X"29",X"ED",X"75",X"FC",X"E4",X"04",X"DD",X"EA",X"AD",X"04",
		X"A7",X"FB",X"EE",X"00",X"EC",X"10",X"41",X"09",X"E8",X"0C",X"8C",X"F1",X"B3",X"12",X"75",X"FE",
		X"49",X"FE",X"48",X"00",X"AC",X"FB",X"56",X"11",X"AD",X"08",X"9F",X"0F",X"78",X"01",X"07",X"ED",
		X"44",X"02",X"98",X"FE",X"D1",X"EB",X"E6",X"09",X"FA",X"0A",X"EE",X"0D",X"9D",X"09",X"F3",X"0F",
		X"F3",X"00",X"16",X"FB",X"55",X"04",X"99",X"EB",X"FA",X"F4",X"2E",X"FE",X"C0",X"15",X"2B",X"F9",
		X"A7",X"02",X"41",X"FB",X"00",X"02",X"45",X"FB",X"6C",X"02",X"68",X"FA",X"ED",X"03",X"99",X"F7",
		X"4F",X"0C",X"87",X"0A",X"76",X"0F",X"0D",X"FD",X"50",X"FE",X"A0",X"00",X"BC",X"EA",X"51",X"09",
		X"65",X"0B",X"59",X"0C",X"7F",X"0C",X"4C",X"FC",X"CB",X"EC",X"8F",X"08",X"E8",X"F5",X"EC",X"08",
		X"C6",X"0D",X"83",X"05",X"0B",X"F5",X"49",X"13",X"34",X"FA",X"63",X"00",X"63",X"FE",X"10",X"ED",
		X"C7",X"F3",X"F1",X"04",X"8D",X"F6",X"A3",X"EE",X"9D",X"F2",X"EB",X"01",X"B0",X"10",X"F1",X"07",
		X"77",X"0F",X"A5",X"08",X"5B",X"0B",X"46",X"E8",X"1A",X"03",X"69",X"FB",X"B6",X"00",X"80",X"FD",
		X"4E",X"EE",X"31",X"F2",X"53",X"F2",X"D1",X"06",X"77",X"F6",X"79",X"0B",X"58",X"0C",X"AF",X"0A",
		X"5E",X"F7",X"E5",X"04",X"62",X"F7",X"5B",X"0B",X"55",X"0C",X"18",X"0B",X"87",X"0C",X"D3",X"0A",
		X"AB",X"0C",X"92",X"0A",X"A3",X"0C",X"28",X"F5",X"21",X"07",X"02",X"F2",X"73",X"F1",X"7A",X"F0",
		X"25",X"F2",X"CF",X"EF",X"A9",X"F4",X"67",X"0A",X"D1",X"0C",X"39",X"0A",X"47",X"0E",X"2F",X"FF",
		X"59",X"EE",X"18",X"F3",X"2E",X"EF",X"C7",X"06",X"E3",X"0B",X"3A",X"F3",X"E4",X"EF",X"78",X"F6",
		X"6C",X"0D",X"35",X"0A",X"90",X"F6",X"9A",X"08",X"50",X"0A",X"CD",X"EC",X"8C",X"FB",X"96",X"0B",
		X"B6",X"0D",X"3B",X"FD",X"4F",X"EE",X"1E",X"F3",X"DA",X"EF",X"56",X"08",X"DE",X"F2",X"67",X"F4",
		X"75",X"0C",X"41",X"0B",X"DE",X"0B",X"CA",X"0B",X"16",X"0B",X"10",X"0D",X"58",X"05",X"DA",X"EF",
		X"CC",X"F0",X"92",X"FB",X"38",X"11",X"D4",X"F8",X"B7",X"EF",X"9D",X"05",X"04",X"0E",X"84",X"09",
		X"14",X"0E",X"0B",X"05",X"69",X"F0",X"73",X"F1",X"11",X"F1",X"64",X"F1",X"FA",X"F0",X"E8",X"F1",
		X"C1",X"EF",X"AF",X"FA",X"43",X"10",X"62",X"FC",X"B0",X"ED",X"CA",X"05",X"92",X"F8",X"84",X"EF",
		X"77",X"0B",X"65",X"0B",X"46",X"08",X"82",X"EC",X"1E",X"FD",X"30",X"0C",X"06",X"0D",X"55",X"FC",
		X"8F",X"ED",X"D9",X"F4",X"7C",X"EC",X"F4",X"01",X"F3",X"FC",X"4C",X"FF",X"91",X"FE",X"C3",X"EA",
		X"F4",X"F7",X"FA",X"02",X"49",X"F7",X"31",X"EB",X"E6",X"FE",X"92",X"FF",X"A8",X"FC",X"DC",X"02",
		X"23",X"EA",X"59",X"08",X"2A",X"F7",X"F9",X"F0",X"6C",X"F0",X"4E",X"FF",X"6E",X"10",X"34",X"F7",
		X"E4",X"F0",X"5C",X"08",X"BC",X"0D",X"20",X"07",X"0C",X"F5",X"5A",X"11",X"F2",X"FD",X"48",X"FD",
		X"98",X"02",X"4A",X"EA",X"55",X"08",X"59",X"F7",X"1F",X"06",X"44",X"0E",X"AF",X"09",X"8A",X"0E",
		X"7B",X"F7",X"E4",X"F0",X"E6",X"F0",X"C5",X"F4",X"F1",X"09",X"BA",X"0E",X"B1",X"01",X"92",X"F9",
		X"D4",X"0E",X"58",X"0B",X"45",X"FD",X"7E",X"ED",X"4F",X"F4",X"5A",X"EF",X"A9",X"F4",X"41",X"0B",
		X"82",X"FC",X"95",X"ED",X"AD",X"F4",X"EA",X"EE",X"D7",X"F5",X"E5",X"0A",X"7E",X"07",X"BA",X"F3",
		X"29",X"15",X"55",X"F8",X"1C",X"03",X"68",X"FB",X"47",X"01",X"42",X"0F",X"23",X"F4",X"A4",X"F0",
		X"6F",X"F5",X"E2",X"0B",X"6B",X"0C",X"8A",X"F6",X"E2",X"F1",X"24",X"08",X"2E",X"F5",X"EB",X"0D",
		X"DB",X"09",X"BD",X"0D",X"93",X"09",X"D8",X"0E",X"88",X"FA",X"53",X"EF",X"40",X"06",X"C2",X"0D",
		X"08",X"0A",X"4F",X"0D",X"E3",X"09",X"98",X"0D",X"E3",X"08",X"EC",X"F8",X"77",X"03",X"6F",X"F6",
		X"88",X"EB",X"3D",X"FF",X"A3",X"FE",X"E3",X"FD",X"80",X"00",X"A9",X"ED",X"FD",X"F2",X"64",X"04",
		X"34",X"F9",X"34",X"06",X"3C",X"0F",X"D8",X"04",X"E0",X"F0",X"13",X"F2",X"C1",X"F1",X"37",X"0C",
		X"D4",X"05",X"9B",X"F7",X"9B",X"07",X"92",X"EA",X"88",X"02",X"8D",X"FD",X"6F",X"FD",X"60",X"12",
		X"5D",X"F2",X"9A",X"F5",X"A6",X"03",X"5F",X"FA",X"A4",X"03",X"43",X"F3",X"03",X"EE",X"56",X"FF",
		X"B0",X"0B",X"1F",X"0E",X"8E",X"03",X"09",X"F3",X"6E",X"ED",X"2D",X"02",X"72",X"FC",X"8E",X"00",
		X"22",X"FD",X"5D",X"ED",X"53",X"F4",X"31",X"F0",X"A9",X"F2",X"C2",X"F1",X"9D",X"F0",X"C7",X"FA",
		X"D7",X"0E",X"60",X"0A",X"07",X"0A",X"2D",X"ED",X"76",X"FD",X"4B",X"02",X"8C",X"F8",X"94",X"14",
		X"DB",X"F4",X"C7",X"06",X"17",X"F7",X"48",X"08",X"4B",X"09",X"EB",X"F6",X"0D",X"07",X"E7",X"EF",
		X"12",X"F2",X"E0",X"FA",X"90",X"12",X"55",X"F7",X"55",X"04",X"B2",X"06",X"40",X"ED",X"45",X"F5",
		X"D6",X"EE",X"1B",X"F5",X"44",X"EE",X"C7",X"09",X"DA",X"08",X"F6",X"F8",X"2C",X"04",X"D9",X"F8",
		X"B1",X"0B",X"EA",X"0D",X"CE",X"FF",X"C0",X"EF",X"32",X"F2",X"19",X"02",X"F8",X"10",X"47",X"FF",
		X"7D",X"F1",X"2C",X"F0",X"AB",X"03",X"C9",X"FB",X"8D",X"01",X"1B",X"FC",X"F6",X"03",X"A8",X"12",
		X"55",X"00",X"B1",X"FB",X"4D",X"0B",X"A7",X"0D",X"E4",X"08",X"01",X"10",X"20",X"F6",X"6A",X"06",
		X"8F",X"0B",X"10",X"0E",X"29",X"FC",X"69",X"F0",X"8E",X"F1",X"52",X"06",X"7E",X"F7",X"DD",X"08",
		X"E3",X"09",X"3F",X"EE",X"99",X"FB",X"37",X"05",X"2F",X"EB",X"F8",X"03",X"0E",X"FD",X"40",X"EE",
		X"46",X"07",X"F2",X"0C",X"60",X"09",X"A4",X"F2",X"0C",X"F2",X"5B",X"F1",X"1A",X"06",X"77",X"F8",
		X"D1",X"05",X"97",X"F3",X"93",X"F1",X"3A",X"F1",X"5C",X"FA",X"BE",X"10",X"A8",X"FC",X"B7",X"EE",
		X"9F",X"05",X"A1",X"F9",X"4B",X"EF",X"5F",X"F3",X"F7",X"F3",X"AF",X"0D",X"80",X"0A",X"56",X"F9",
		X"D5",X"03",X"41",X"F9",X"6E",X"09",X"34",X"09",X"4C",X"EC",X"AB",X"FE",X"57",X"0C",X"BC",X"0B",
		X"85",X"0C",X"0B",X"FA",X"3D",X"02",X"03",X"11",X"5A",X"05",X"DB",X"F8",X"80",X"0A",X"7D",X"07",
		X"96",X"EC",X"FF",X"0D",X"9B",X"04",X"C7",X"FA",X"74",X"03",X"4C",X"F3",X"45",X"EE",X"F0",X"00",
		X"AB",X"FF",X"BB",X"ED",X"29",X"05",X"F5",X"0D",X"5B",X"F3",X"77",X"F5",X"0F",X"06",X"FE",X"F6",
		X"8C",X"0D",X"85",X"0A",X"80",X"0C",X"D9",X"0A",X"74",X"0C",X"4C",X"0A",X"08",X"0E",X"50",X"00",
		X"BE",X"F9",X"97",X"12",X"88",X"F7",X"7F",X"F2",X"B2",X"F0",X"9B",X"08",X"02",X"F3",X"0D",X"F5",
		X"83",X"0D",X"74",X"03",X"40",X"F7",X"E1",X"11",X"56",X"04",X"BA",X"F5",X"3D",X"F2",X"E5",X"14",
		X"06",X"F9",X"E7",X"02",X"2C",X"FB",X"4D",X"01",X"ED",X"0C",X"2B",X"0C",X"9B",X"08",X"C3",X"F6",
		X"74",X"EC",X"0E",X"FD",X"FA",X"FF",X"30",X"FD",X"4A",X"01",X"01",X"F0",X"D3",X"F0",X"0A",X"F9",
		X"08",X"0B",X"E6",X"0E",X"E6",X"FB",X"1E",X"00",X"4A",X"FE",X"2E",X"EE",X"81",X"F3",X"CE",X"F2",
		X"D8",X"06",X"89",X"F7",X"42",X"06",X"76",X"F5",X"5A",X"12",X"BA",X"FB",X"EC",X"FD",X"07",X"10",
		X"3F",X"F8",X"7A",X"F0",X"60",X"F3",X"7E",X"EF",X"96",X"01",X"D5",X"FE",X"B1",X"EC",X"A7",X"F6",
		X"A9",X"03",X"27",X"12",X"46",X"01",X"2C",X"FD",X"64",X"00",X"FA",X"FC",X"56",X"01",X"7D",X"FA",
		X"FA",X"12",X"10",X"F5",X"0B",X"07",X"41",X"04",X"71",X"EB",X"D9",X"04",X"25",X"FB",X"35",X"01",
		X"0C",X"10",X"15",X"07",X"E8",X"F6",X"B0",X"ED",X"21",X"FB",X"81",X"04",X"DD",X"EE",X"6B",X"FD",
		X"80",X"0F",X"EE",X"07",X"BF",X"0F",X"17",X"F4",X"67",X"09",X"75",X"F0",X"C0",X"03",X"AB",X"FA",
		X"EA",X"02",X"AF",X"F9",X"B8",X"F0",X"1F",X"09",X"F5",X"F1",X"20",X"F2",X"EC",X"F2",X"E5",X"EF",
		X"75",X"FE",X"3B",X"0D",X"50",X"0C",X"5B",X"F9",X"91",X"03",X"BE",X"0D",X"DA",X"F3",X"2A",X"0C",
		X"45",X"0A",X"AD",X"0C",X"45",X"0A",X"9A",X"0C",X"1F",X"0A",X"D8",X"0C",X"65",X"09",X"6F",X"0E",
		X"3E",X"00",X"2E",X"F1",X"32",X"F0",X"20",X"03",X"A6",X"FB",X"2F",X"01",X"28",X"FC",X"6E",X"01",
		X"26",X"FB",X"DE",X"03",X"1A",X"F2",X"BA",X"04",X"DB",X"F9",X"62",X"03",X"40",X"F9",X"31",X"06",
		X"0D",X"EE",X"3E",X"FE",X"0F",X"02",X"05",X"EE",X"D1",X"F3",X"6F",X"01",X"01",X"10",X"F8",X"06",
		X"50",X"F8",X"4B",X"09",X"B8",X"07",X"69",X"F4",X"B9",X"11",X"0A",X"06",X"C5",X"0E",X"D5",X"EA",
		X"50",X"FF",X"3A",X"FE",X"7E",X"FE",X"38",X"00",X"5F",X"F0",X"EC",X"F0",X"FF",X"04",X"07",X"F9",
		X"A5",X"F0",X"A9",X"0A",X"5B",X"0B",X"E5",X"0A",X"CA",X"0C",X"7F",X"02",X"CD",X"EF",X"11",X"0D",
		X"05",X"05",X"51",X"F7",X"A9",X"0D",X"38",X"09",X"EA",X"0D",X"F5",X"FC",X"9D",X"EE",X"B7",X"04",
		X"EB",X"0C",X"EC",X"F4",X"EC",X"09",X"EE",X"07",X"1B",X"F1",X"8C",X"F2",X"99",X"F1",X"68",X"F2",
		X"5F",X"F1",X"A0",X"F5",X"77",X"0D",X"9D",X"08",X"6E",X"0F",X"D1",X"FB",X"65",X"FF",X"70",X"FF",
		X"31",X"EC",X"9F",X"09",X"19",X"09",X"51",X"F5",X"89",X"EF",X"26",X"F8",X"27",X"0D",X"FF",X"02",
		X"E4",X"EC",X"43",X"02",X"AE",X"FE",X"2D",X"EC",X"06",X"FE",X"4E",X"02",X"34",X"EF",X"B0",X"F3",
		X"5B",X"F1",X"72",X"F2",X"24",X"05",X"84",X"F8",X"28",X"EE",X"40",X"F9",X"33",X"05",X"84",X"F1",
		X"C1",X"F1",X"BD",X"FB",X"C3",X"11",X"76",X"F7",X"D5",X"04",X"FD",X"04",X"C8",X"F6",X"CE",X"13",
		X"9E",X"F7",X"D5",X"02",X"E2",X"0C",X"06",X"0B",X"8D",X"0A",X"55",X"F3",X"10",X"F5",X"43",X"0D",
		X"6B",X"09",X"6A",X"0D",X"A0",X"08",X"54",X"0F",X"7E",X"F8",X"2A",X"03",X"C4",X"FA",X"BC",X"ED",
		X"FD",X"FE",X"41",X"0F",X"E3",X"F8",X"67",X"02",X"84",X"0E",X"DA",X"08",X"7F",X"0D",X"3E",X"06",
		X"F1",X"F1",X"5C",X"F2",X"B5",X"F1",X"21",X"F3",X"F7",X"EF",X"F4",X"02",X"BD",X"FC",X"DC",X"ED",
		X"A6",X"0A",X"D2",X"09",X"FB",X"0C",X"40",X"09",X"86",X"0D",X"61",X"F5",X"28",X"F2",X"19",X"F3",
		X"BB",X"0D",X"8E",X"03",X"25",X"F3",X"04",X"EF",X"5D",X"00",X"AD",X"FF",X"E3",X"EE",X"92",X"F3",
		X"30",X"04",X"DD",X"F9",X"CA",X"05",X"A6",X"0E",X"40",X"08",X"48",X"0E",X"04",X"F5",X"FD",X"07",
		X"55",X"F2",X"97",X"F7",X"A9",X"05",X"D7",X"F5",X"60",X"12",X"6C",X"FA",X"88",X"00",X"DE",X"FE",
		X"22",X"ED",X"C5",X"08",X"B8",X"09",X"8E",X"F6",X"F5",X"09",X"54",X"0B",X"A2",X"0B",X"9D",X"F6",
		X"8F",X"F2",X"97",X"07",X"7E",X"F5",X"46",X"0D",X"4F",X"09",X"B1",X"0C",X"B4",X"09",X"24",X"0C",
		X"A7",X"0A",X"3F",X"FB",X"E7",X"ED",X"73",X"0A",X"A7",X"F0",X"E9",X"F8",X"61",X"03",X"9C",X"F8",
		X"16",X"0D",X"76",X"09",X"84",X"F2",X"C5",X"F6",X"FE",X"06",X"20",X"EE",X"8D",X"FC",X"8F",X"0E",
		X"A4",X"FC",X"DB",X"EF",X"7A",X"F3",X"C1",X"F1",X"90",X"06",X"CC",X"F7",X"72",X"05",X"35",X"F7",
		X"2A",X"08",X"29",X"EB",X"95",X"01",X"8F",X"09",X"E0",X"0E",X"2D",X"01",X"C9",X"FB",X"45",X"02",
		X"FE",X"F8",X"86",X"12",X"9B",X"F6",X"CE",X"03",X"08",X"0D",X"F9",X"08",X"E9",X"F4",X"43",X"F0",
		X"D9",X"F7",X"8D",X"0C",X"DD",X"09",X"3F",X"0C",X"4E",X"09",X"C5",X"0D",X"6D",X"02",X"A7",X"F9",
		X"44",X"05",X"87",X"EB",X"9C",X"02",X"83",X"0C",X"40",X"F9",X"0D",X"02",X"21",X"FB",X"B2",X"03",
		X"3D",X"11",X"CE",X"FF",X"56",X"FC",X"45",X"02",X"E4",X"EF",X"EB",X"F2",X"02",X"F2",X"FA",X"F1",
		X"D8",X"F2",X"BA",X"F0",X"13",X"FD",X"27",X"10",X"EC",X"F7",X"47",X"03",X"4B",X"FA",X"43",X"EE",
		X"26",X"F7",X"6F",X"08",X"91",X"0D",X"7D",X"03",X"F2",X"EE",X"14",X"FE",X"38",X"0D",X"90",X"0A",
		X"59",X"FB",X"66",X"EE",X"95",X"F5",X"79",X"EE",X"AE",X"01",X"35",X"0D",X"45",X"F9",X"9D",X"EF",
		X"C5",X"F4",X"87",X"EF",X"A3",X"F8",X"CC",X"05",X"DE",X"EF",X"44",X"FB",X"B9",X"0F",X"1A",X"FC",
		X"2D",X"F1",X"74",X"F2",X"FB",X"04",X"C6",X"0D",X"B3",X"08",X"7E",X"0E",X"CF",X"F8",X"C4",X"02",
		X"EE",X"0D",X"37",X"09",X"82",X"0C",X"8A",X"09",X"F4",X"0C",X"BC",X"03",X"A5",X"EE",X"58",X"FE",
		X"58",X"0D",X"74",X"09",X"25",X"0C",X"86",X"09",X"C0",X"F7",X"E0",X"ED",X"0E",X"03",X"D9",X"FC",
		X"4F",X"EE",X"79",X"08",X"52",X"09",X"4D",X"F6",X"15",X"0A",X"49",X"0B",X"35",X"0A",X"79",X"0C",
		X"F3",X"FF",X"AA",X"EE",X"FF",X"F4",X"63",X"EF",X"2B",X"07",X"E6",X"F6",X"96",X"06",X"D5",X"F2",
		X"11",X"F3",X"F5",X"F0",X"27",X"07",X"60",X"0B",X"08",X"0B",X"DE",X"0A",X"43",X"07",X"0B",X"ED",
		X"C7",X"FE",X"00",X"0A",X"15",X"0E",X"9E",X"F8",X"B7",X"02",X"56",X"0C",X"D0",X"F6",X"90",X"04",
		X"98",X"F8",X"52",X"05",X"E8",X"F0",X"80",X"05",X"C7",X"F8",X"64",X"04",X"6D",X"F4",X"3B",X"F4",
		X"F9",X"11",X"18",X"FB",X"33",X"00",X"60",X"FE",X"18",X"F0",X"9D",X"F2",X"3E",X"F3",X"4C",X"F0",
		X"6E",X"F7",X"7B",X"03",X"4F",X"FA",X"2F",X"03",X"A6",X"F8",X"1E",X"0F",X"89",X"06",X"E0",X"F2",
		X"A5",X"F6",X"04",X"0F",X"E7",X"FF",X"F6",X"F0",X"47",X"F2",X"5A",X"00",X"8C",X"0F",X"64",X"F4",
		X"75",X"F4",X"C4",X"07",X"EB",X"0A",X"B1",X"EC",X"04",X"FF",X"46",X"FF",X"DC",X"FC",X"32",X"0A",
		X"B9",X"F5",X"6A",X"08",X"B5",X"EC",X"A1",X"FF",X"92",X"01",X"D8",X"EC",X"B4",X"05",X"C0",X"F9",
		X"5E",X"03",X"36",X"0E",X"CC",X"08",X"78",X"0A",X"48",X"ED",X"2B",X"FE",X"A8",X"00",X"86",X"FA",
		X"15",X"10",X"85",X"03",X"30",X"F8",X"16",X"0D",X"11",X"09",X"BD",X"0C",X"80",X"08",X"13",X"0E",
		X"CF",X"F6",X"27",X"F3",X"F3",X"EF",X"27",X"F8",X"9D",X"02",X"5D",X"FB",X"7E",X"01",X"A1",X"FB",
		X"8E",X"02",X"22",X"EF",X"A4",X"F2",X"FD",X"03",X"00",X"05",X"FC",X"F6",X"6E",X"11",X"B2",X"05",
		X"12",X"10",X"40",X"F5",X"D8",X"06",X"BC",X"09",X"5C",X"F6",X"99",X"09",X"00",X"0C",X"62",X"04",
		X"32",X"EE",X"98",X"FE",X"68",X"0D",X"19",X"FC",X"3B",X"EE",X"A3",X"08",X"DE",X"01",X"1B",X"EE",
		X"F1",X"01",X"7A",X"FE",X"9E",X"EC",X"30",X"0A",X"6C",X"F2",X"44",X"F7",X"DB",X"06",X"30",X"10",
		X"F5",X"FD",X"9D",X"FE",X"FA",X"FE",X"F1",X"FC",X"43",X"0E",X"29",X"09",X"29",X"0B",X"9A",X"F6",
		X"35",X"EF",X"48",X"01",X"B7",X"0C",X"A2",X"F9",X"CF",X"EE",X"64",X"F6",X"61",X"ED",X"1F",X"FC",
		X"F2",X"FF",X"D1",X"FD",X"10",X"FF",X"7A",X"FE",X"92",X"FE",X"CB",X"FE",X"98",X"FE",X"4F",X"ED",
		X"E6",X"0A",X"CA",X"07",X"C2",X"F3",X"76",X"F2",X"01",X"F2",X"C1",X"06",X"2F",X"0A",X"60",X"F6",
		X"5A",X"07",X"2C",X"F0",X"39",X"FA",X"8D",X"0D",X"39",X"08",X"B0",X"0E",X"64",X"F8",X"82",X"03",
		X"A6",X"F9",X"56",X"F1",X"EB",X"07",X"9F",X"F5",X"42",X"0C",X"86",X"09",X"C6",X"0B",X"00",X"0A",
		X"20",X"0B",X"04",X"0B",X"15",X"06",X"7E",X"EF",X"29",X"F5",X"34",X"EF",X"D8",X"00",X"18",X"0D",
		X"9F",X"F9",X"C1",X"EF",X"F9",X"09",X"2C",X"07",X"7B",X"F7",X"F5",X"09",X"FF",X"0B",X"9F",X"F5",
		X"30",X"F4",X"AD",X"05",X"C6",X"F7",X"94",X"06",X"A6",X"EE",X"A7",X"FC",X"1D",X"0E",X"9E",X"FC",
		X"5C",X"F0",X"D6",X"F3",X"D8",X"F1",X"0A",X"F3",X"E6",X"F3",X"B8",X"0B",X"DD",X"05",X"E8",X"EF",
		X"C9",X"FB",X"97",X"0D",X"F8",X"06",X"77",X"F3",X"55",X"F2",X"01",X"F3",X"8B",X"F2",X"F2",X"F2",
		X"B4",X"F2",X"E2",X"F2",X"E4",X"F2",X"B3",X"F2",X"ED",X"F3",X"85",X"09",X"1F",X"09",X"33",X"EF",
		X"1D",X"FD",X"2C",X"02",X"EE",X"F9",X"E5",X"0E",X"85",X"EC",X"B8",X"FE",X"1C",X"00",X"C2",X"FC",
		X"58",X"03",X"7E",X"EC",X"69",X"06",X"DD",X"F9",X"99",X"03",X"76",X"0E",X"6D",X"08",X"31",X"0B",
		X"BE",X"EC",X"04",X"00",X"A1",X"FE",X"E6",X"FE",X"78",X"FF",X"80",X"FD",X"2F",X"10",X"38",X"07",
		X"A5",X"0E",X"8D",X"FE",X"56",X"EF",X"2E",X"04",X"A6",X"FB",X"D3",X"EF",X"CE",X"09",X"0C",X"0B",
		X"AB",X"07",X"1F",X"F5",X"B9",X"10",X"C4",X"FD",X"A9",X"FC",X"D6",X"0E",X"4F",X"FB",X"B6",X"EF",
		X"3E",X"FB",X"2C",X"0D",X"E3",X"08",X"C1",X"0D",X"50",X"F9",X"AE",X"02",X"1A",X"FB",X"89",X"EE",
		X"B6",X"F6",X"72",X"EE",X"53",X"FC",X"7F",X"02",X"18",X"F9",X"BB",X"10",X"8B",X"FA",X"FB",X"FF",
		X"ED",X"0E",X"46",X"F6",X"D9",X"F1",X"E5",X"FC",X"90",X"10",X"0B",X"F8",X"9E",X"F3",X"76",X"F1",
		X"9C",X"0A",X"6F",X"06",X"36",X"F9",X"46",X"05",X"E6",X"F1",X"ED",X"F2",X"FE",X"F3",X"92",X"F0",
		X"B2",X"03",X"42",X"FC",X"BC",X"EF",X"BC",X"09",X"30",X"0A",X"AA",X"0C",X"53",X"FB",X"6F",X"F0",
		X"F5",X"F4",X"1C",X"F2",X"71",X"0C",X"58",X"05",X"82",X"F4",X"45",X"F0",X"BC",X"FD",X"B6",X"0B",
		X"6F",X"0C",X"AF",X"FB",X"2E",X"F1",X"EF",X"F3",X"ED",X"F2",X"14",X"F3",X"A0",X"F3",X"90",X"F2",
		X"39",X"F4",X"4C",X"F2",X"21",X"0A",X"26",X"08",X"6E",X"F4",X"ED",X"F1",X"77",X"F5",X"A5",X"EF",
		X"7D",X"01",X"BA",X"FF",X"2C",X"F0",X"2C",X"F5",X"89",X"F2",X"BF",X"07",X"D9",X"F5",X"89",X"F2",
		X"44",X"F4",X"BD",X"F2",X"D2",X"F4",X"99",X"06",X"6C",X"F6",X"1A",X"F2",X"4D",X"F4",X"3D",X"F8",
		X"CD",X"11",X"5E",X"FC",X"D5",X"F4",X"76",X"F0",X"7B",X"07",X"39",X"F8",X"B5",X"F3",X"D8",X"F1",
		X"A2",X"F9",X"EA",X"04",X"3C",X"F9",X"F7",X"0D",X"96",X"F4",X"31",X"F6",X"66",X"09",X"D4",X"EE",
		X"E7",X"FF",X"49",X"00",X"84",X"FE",X"54",X"01",X"E3",X"FC",X"DC",X"12",X"AA",X"F3",X"7C",X"0A",
		X"7A",X"F2",X"81",X"F9",X"63",X"09",X"FE",X"0E",X"81",X"00",X"CE",X"F4",X"1D",X"09",X"52",X"0E",
		X"A4",X"03",X"C8",X"F4",X"24",X"F0",X"AB",X"02",X"BD",X"FD",X"23",X"01",X"16",X"FE",X"AA",X"01",
		X"22",X"10",X"F6",X"EF",X"B5",X"FB",X"64",X"03",X"51",X"FA",X"7C",X"0D",X"A3",X"0A",X"04",X"0A",
		X"CF",X"F1",X"E6",X"F9",X"CA",X"0D",X"62",X"02",X"68",X"EF",X"57",X"02",X"D6",X"0D",X"BA",X"F9",
		X"92",X"03",X"1B",X"FC",X"3B",X"03",X"AF",X"F8",X"39",X"EE",X"B7",X"FF",X"61",X"01",X"C7",X"F3",
		X"0E",X"F1",X"F6",X"04",X"69",X"06",X"C0",X"F2",X"54",X"F2",X"4B",X"00",X"B1",X"01",X"07",X"EE",
		X"78",X"08",X"6C",X"F8",X"D7",X"F2",X"16",X"F4",X"69",X"F6",X"72",X"0E",X"72",X"03",X"67",X"F2",
		X"00",X"F5",X"2C",X"F2",X"13",X"03",X"31",X"FF",X"F9",X"EC",X"05",X"03",X"DC",X"FE",X"9B",X"FE",
		X"A5",X"10",X"B9",X"F7",X"FA",X"05",X"24",X"FA",X"C5",X"05",X"48",X"F8",X"F9",X"0D",X"87",X"02",
		X"71",X"FB",X"6D",X"06",X"74",X"EB",X"F5",X"08",X"F4",X"F8",X"E6",X"F4",X"F6",X"F0",X"F2",X"01",
		X"92",X"00",X"4C",X"EF",X"D2",X"07",X"5B",X"F9",X"E7",X"F1",X"C0",X"F7",X"43",X"08",X"11",X"F1",
		X"CC",X"FD",X"A8",X"03",X"DC",X"F9",X"AA",X"13",X"35",X"F7",X"62",X"06",X"06",X"FA",X"DD",X"F2",
		X"27",X"0C",X"98",X"FE",X"FC",X"F0",X"80",X"F6",X"56",X"F2",X"42",X"0B",X"93",X"08",X"D1",X"F4",
		X"51",X"F7",X"64",X"11",X"FF",X"FD",X"EC",X"FF",X"0A",X"02",X"BE",X"EE",X"E1",X"07",X"E5",X"F9",
		X"FC",X"F1",X"61",X"F6",X"25",X"F1",X"15",X"06",X"59",X"FB",X"FD",X"04",X"85",X"0D",X"D3",X"F4",
		X"3D",X"0F",X"FD",X"02",X"30",X"FB",X"DA",X"0D",X"8F",X"0A",X"6B",X"0C",X"F6",X"0A",X"49",X"0C",
		X"B3",X"0A",X"F0",X"0C",X"E0",X"07",X"2D",X"F9",X"4A",X"07",X"C8",X"F1",X"0D",X"F6",X"B2",X"07",
		X"E3",X"0B",X"8E",X"F0",X"B5",X"FC",X"F9",X"04",X"C3",X"F0",X"25",X"FF",X"F8",X"0F",X"F3",X"F9",
		X"91",X"03",X"FD",X"0D",X"67",X"F6",X"57",X"0A",X"34",X"0B",X"09",X"0C",X"A8",X"0A",X"F6",X"0B",
		X"37",X"F6",X"2D",X"0C",X"3F",X"05",X"77",X"FA",X"0F",X"06",X"93",X"F0",X"EA",X"F5",X"0E",X"F3",
		X"D9",X"F3",X"76",X"04",X"18",X"FC",X"30",X"04",X"55",X"10",X"0F",X"04",X"34",X"FA",X"E1",X"0C",
		X"A5",X"03",X"13",X"F0",X"7D",X"F7",X"EA",X"EF",X"4B",X"FD",X"0F",X"04",X"45",X"F2",X"D4",X"F4",
		X"D6",X"F3",X"53",X"F4",X"F9",X"F3",X"1C",X"06",X"7E",X"0E",X"8A",X"06",X"6A",X"FA",X"A8",X"05",
		X"1B",X"F8",X"46",X"11",X"26",X"FD",X"1C",X"FF",X"36",X"0F",X"49",X"08",X"75",X"0F",X"DD",X"FE",
		X"F4",X"FD",X"38",X"0E",X"93",X"0A",X"97",X"FB",X"A8",X"02",X"D8",X"FC",X"15",X"03",X"B7",X"F8",
		X"4B",X"EF",X"20",X"FE",X"63",X"0A",X"68",X"0D",X"5A",X"08",X"9B",X"0F",X"17",X"01",X"73",X"FD",
		X"50",X"03",X"24",X"F1",X"40",X"F5",X"8E",X"F3",X"03",X"F4",X"E8",X"F4",X"7B",X"06",X"E8",X"F7",
		X"6A",X"F0",X"DB",X"FC",X"4C",X"03",X"A4",X"FA",X"28",X"0F",X"03",X"09",X"06",X"0D",X"EC",X"09",
		X"6A",X"0C",X"3D",X"0A",X"19",X"0C",X"6C",X"0A",X"CA",X"0B",X"C1",X"0A",X"A8",X"F9",X"86",X"05",
		X"E6",X"0E",X"D8",X"04",X"60",X"F5",X"FE",X"F1",X"6A",X"F6",X"3F",X"F0",X"C1",X"02",X"73",X"0B",
		X"34",X"0C",X"0C",X"09",X"A3",X"0E",X"73",X"FD",X"FE",X"F3",X"A1",X"F1",X"37",X"07",X"0A",X"F8",
		X"27",X"09",X"5C",X"07",X"11",X"FA",X"60",X"04",X"F0",X"F9",X"C6",X"0C",X"41",X"0C",X"07",X"FD",
		X"96",X"00",X"ED",X"FE",X"F6",X"EE",X"D9",X"0A",X"9A",X"F2",X"B2",X"01",X"E2",X"0D",X"F9",X"F8",
		X"05",X"F3",X"02",X"09",X"1F",X"0A",X"6C",X"F1",X"BA",X"FB",X"B2",X"04",X"BD",X"F1",X"1D",X"F4",
		X"E9",X"FE",X"2B",X"10",X"70",X"F7",X"E5",X"05",X"A8",X"F8",X"DC",X"F1",X"C7",X"F5",X"D3",X"F1",
		X"2D",X"06",X"30",X"0C",X"A9",X"09",X"12",X"F5",X"9B",X"F3",X"D2",X"F7",X"1E",X"10",X"4B",X"FE",
		X"24",X"FE",X"6C",X"0D",X"C0",X"0A",X"82",X"FB",X"53",X"F1",X"D2",X"09",X"94",X"0A",X"A8",X"0B",
		X"45",X"0A",X"C8",X"0B",X"2E",X"F8",X"F2",X"06",X"79",X"0D",X"49",X"05",X"3E",X"F8",X"7D",X"0E",
		X"13",X"01",X"A9",X"F0",X"40",X"01",X"63",X"0D",X"1A",X"09",X"93",X"0C",X"35",X"08",X"3E",X"F7",
		X"93",X"F0",X"83",X"FB",X"AA",X"04",X"FD",X"F1",X"C1",X"09",X"0B",X"09",X"32",X"F2",X"16",X"FA",
		X"F0",X"0B",X"A4",X"0A",X"58",X"0A",X"5F",X"0C",X"BA",X"FB",X"DA",X"F1",X"C8",X"F4",X"EA",X"07",
		X"32",X"09",X"18",X"F7",X"48",X"08",X"B7",X"EF",X"61",X"F7",X"2C",X"F0",X"8C",X"F9",X"E0",X"07",
		X"FB",X"0D",X"FB",X"06",X"2D",X"10",X"E5",X"FA",X"64",X"01",X"50",X"0B",X"31",X"0C",X"8F",X"F6",
		X"5F",X"09",X"9F",X"06",X"52",X"FA",X"98",X"03",X"30",X"FA",X"C3",X"0B",X"5C",X"0C",X"E4",X"FC",
		X"AC",X"F6",X"6F",X"07",X"BF",X"EF",X"4F",X"FD",X"33",X"0F",X"38",X"FA",X"9E",X"02",X"49",X"FC",
		X"E6",X"F0",X"16",X"F5",X"90",X"F3",X"C9",X"F2",X"83",X"F9",X"1E",X"0B",X"A4",X"0C",X"8B",X"FE",
		X"DC",X"FD",X"21",X"0E",X"D0",X"09",X"48",X"04",X"A3",X"F7",X"03",X"13",X"51",X"F7",X"E6",X"04",
		X"4A",X"FA",X"60",X"04",X"F5",X"0B",X"D4",X"F4",X"2F",X"0D",X"96",X"03",X"E5",X"F3",X"B6",X"F2",
		X"91",X"F5",X"9F",X"F0",X"B0",X"04",X"51",X"FB",X"B5",X"02",X"33",X"0F",X"C4",X"FD",X"2B",X"F2",
		X"CB",X"F4",X"FB",X"F2",X"BA",X"F4",X"B0",X"F3",X"93",X"0B",X"D0",X"05",X"AF",X"F4",X"B3",X"F1",
		X"A4",X"FD",X"D2",X"0B",X"EF",X"0B",X"77",X"FB",X"C3",X"01",X"4B",X"FD",X"D9",X"01",X"E5",X"11",
		X"A3",X"F7",X"1E",X"05",X"FA",X"F9",X"A5",X"04",X"0C",X"F9",X"F4",X"08",X"49",X"07",X"B9",X"F6",
		X"40",X"0F",X"F2",X"FF",X"80",X"F2",X"C2",X"F4",X"81",X"F2",X"3F",X"04",X"DB",X"0C",X"26",X"08",
		X"64",X"F8",X"EF",X"08",X"3C",X"0C",X"30",X"F9",X"89",X"04",X"62",X"0C",X"C1",X"F3",X"33",X"0F",
		X"14",X"00",X"18",X"FE",X"B3",X"00",X"82",X"FC",X"6D",X"0D",X"3D",X"0A",X"7B",X"FA",X"79",X"03",
		X"94",X"0C",X"60",X"F3",X"B3",X"F4",X"25",X"F3",X"2E",X"F4",X"C9",X"F3",X"5E",X"F4",X"78",X"0B",
		X"B8",X"04",X"1F",X"FA",X"5B",X"05",X"EA",X"F0",X"8F",X"F4",X"C3",X"FE",X"BC",X"0E",X"A5",X"07",
		X"B9",X"0C",X"AE",X"F5",X"05",X"0A",X"C7",X"09",X"6B",X"0B",X"99",X"09",X"5B",X"F9",X"62",X"F0",
		X"48",X"F9",X"E6",X"04",X"42",X"F4",X"F6",X"F2",X"5C",X"F5",X"4B",X"F1",X"B9",X"01",X"E4",X"0B",
		X"9F",X"0A",X"CD",X"F8",X"64",X"05",X"A9",X"F6",X"4A",X"F3",X"0A",X"F3",X"2F",X"FB",X"4B",X"05",
		X"53",X"F0",X"FB",X"0B",X"51",X"EE",X"37",X"FF",X"3A",X"00",X"E7",X"FC",X"FA",X"0B",X"9A",X"0B",
		X"D6",X"FB",X"27",X"F2",X"E6",X"F4",X"BF",X"07",X"CB",X"09",X"D0",X"F2",X"D4",X"F8",X"9D",X"0D",
		X"4E",X"01",X"15",X"F2",X"36",X"F5",X"AD",X"F2",X"6D",X"F9",X"3E",X"0D",X"27",X"08",X"43",X"0E",
		X"13",X"FB",X"48",X"01",X"8B",X"0D",X"7F",X"F7",X"53",X"F2",X"07",X"F8",X"48",X"05",X"1A",X"F9",
		X"4F",X"07",X"E7",X"ED",X"7D",X"02",X"9D",X"FF",X"4D",X"F0",X"01",X"FB",X"5D",X"0C",X"AC",X"02",
		X"A9",X"EE",X"06",X"05",X"85",X"FB",X"BC",X"02",X"BE",X"FB",X"77",X"F0",X"F8",X"F6",X"A7",X"F1",
		X"EC",X"F6",X"92",X"F0",X"7F",X"FF",X"94",X"02",X"3F",X"EF",X"CD",X"04",X"E7",X"0A",X"71",X"0C",
		X"AF",X"00",X"51",X"FB",X"99",X"11",X"21",X"F7",X"0A",X"06",X"27",X"F9",X"81",X"07",X"0C",X"09",
		X"55",X"F7",X"C1",X"08",X"5F",X"EE",X"14",X"01",X"04",X"01",X"C0",X"F0",X"04",X"03",X"32",X"0D",
		X"9C",X"08",X"F5",X"0C",X"D9",X"07",X"B9",X"0E",X"3F",X"F8",X"78",X"05",X"BB",X"F8",X"A7",X"F4",
		X"B5",X"08",X"3B",X"0D",X"B7",X"02",X"FB",X"FA",X"80",X"0B",X"64",X"0C",X"46",X"FC",X"2D",X"01",
		X"F9",X"FD",X"08",X"F0",X"75",X"F7",X"73",X"07",X"CF",X"0B",X"77",X"0A",X"96",X"FA",X"EE",X"F1",
		X"45",X"F5",X"CE",X"F3",X"6E",X"F3",X"8C",X"F9",X"AC",X"0B",X"AF",X"0B",X"57",X"FF",X"17",X"FD",
		X"8C",X"0F",X"F4",X"06",X"A7",X"0D",X"DC",X"06",X"5E",X"F8",X"50",X"F0",X"1B",X"05",X"D6",X"0A",
		X"9F",X"0A",X"89",X"F5",X"85",X"F6",X"F1",X"07",X"8A",X"F0",X"C3",X"FD",X"83",X"03",X"C7",X"EF",
		X"AC",X"01",X"77",X"0D",X"F5",X"F8",X"51",X"04",X"9F",X"FA",X"75",X"04",X"D4",X"F8",X"9A",X"0B",
		X"66",X"F9",X"5A",X"F3",X"39",X"08",X"50",X"0C",X"01",X"05",X"11",X"F9",X"F0",X"0B",X"19",X"0B",
		X"AE",X"FF",X"33",X"FC",X"21",X"11",X"C3",X"F5",X"48",X"07",X"4D",X"0A",X"C3",X"09",X"A4",X"F1",
		X"68",X"FB",X"84",X"04",X"89",X"F1",X"E5",X"F6",X"BD",X"06",X"62",X"F3",X"6B",X"F9",X"6E",X"0C",
		X"07",X"09",X"9F",X"0B",X"07",X"09",X"38",X"0C",X"7A",X"F9",X"8D",X"F2",X"DB",X"F5",X"48",X"08",
		X"EA",X"0B",X"28",X"05",X"8E",X"F2",X"DD",X"F4",X"9E",X"F4",X"33",X"0A",X"F2",X"09",X"80",X"0A",
		X"0B",X"0B",X"45",X"02",X"9C",X"F0",X"E8",X"F5",X"2C",X"FF",X"70",X"10",X"6F",X"F3",X"C3",X"0B",
		X"DF",X"03",X"BF",X"FC",X"DA",X"00",X"C5",X"FD",X"92",X"00",X"26",X"FD",X"D7",X"09",X"C9",X"F6",
		X"32",X"08",X"64",X"EE",X"95",X"00",X"60",X"01",X"F5",X"EE",X"E0",X"05",X"59",X"FA",X"0F",X"F3",
		X"EA",X"06",X"9C",X"F6",X"E7",X"F1",X"77",X"FA",X"4C",X"0A",X"5E",X"0C",X"8A",X"FE",X"8A",X"FD",
		X"6F",X"0E",X"03",X"08",X"E5",X"06",X"89",X"EC",X"2D",X"05",X"F9",X"FA",X"CA",X"02",X"BA",X"FB",
		X"65",X"03",X"1F",X"0C",X"C9",X"F4",X"FD",X"0C",X"6E",X"03",X"FB",X"F3",X"9B",X"F3",X"15",X"F5",
		X"38",X"F2",X"EB",X"02",X"F5",X"FD",X"35",X"EE",X"C0",X"01",X"86",X"FF",X"99",X"F2",X"D3",X"F3",
		X"D1",X"04",X"03",X"FA",X"1B",X"F3",X"97",X"0A",X"42",X"0A",X"AB",X"06",X"67",X"F0",X"F7",X"FD",
		X"0A",X"0D",X"14",X"FE",X"5C",X"F1",X"B9",X"F6",X"10",X"F1",X"97",X"FF",X"4E",X"02",X"91",X"EE",
		X"D4",X"06",X"B6",X"F9",X"0C",X"05",X"79",X"0C",X"BB",X"07",X"4C",X"F3",X"82",X"FA",X"E4",X"05",
		X"2E",X"F0",X"E6",X"F7",X"1A",X"F0",X"E0",X"05",X"83",X"FA",X"12",X"04",X"C7",X"F9",X"ED",X"F1",
		X"38",X"F6",X"1D",X"F3",X"8C",X"F5",X"3B",X"05",X"7F",X"0C",X"2E",X"F2",X"94",X"FA",X"DD",X"08",
		X"97",X"0D",X"17",X"00",X"39",X"F4",X"A1",X"F2",X"13",X"04",X"81",X"FC",X"B6",X"F1",X"3B",X"F6",
		X"92",X"F4",X"31",X"0D",X"FD",X"F9",X"A2",X"03",X"C8",X"0C",X"F7",X"F5",X"6D",X"0B",X"B3",X"05",
		X"07",X"F5",X"C2",X"F2",X"C2",X"FD",X"55",X"0C",X"A4",X"0A",X"8F",X"FD",X"FF",X"F0",X"3E",X"08",
		X"C3",X"09",X"79",X"F5",X"A9",X"F7",X"10",X"08",X"89",X"F0",X"FD",X"09",X"77",X"08",X"DA",X"0D",
		X"32",X"03",X"DB",X"FB",X"88",X"04",X"EF",X"F1",X"30",X"F6",X"B5",X"F2",X"D3",X"02",X"28",X"0D",
		X"2B",X"08",X"C6",X"F9",X"6C",X"F0",X"00",X"FC",X"F9",X"02",X"FF",X"FA",X"12",X"0C",X"3C",X"0A",
		X"37",X"0A",X"33",X"0B",X"60",X"09",X"F1",X"0B",X"54",X"08",X"B0",X"0D",X"02",X"FC",X"41",X"F4",
		X"2B",X"F3",X"C9",X"07",X"7F",X"08",X"91",X"F9",X"1F",X"05",X"A1",X"F5",X"E7",X"F1",X"7E",X"FE",
		X"64",X"09",X"58",X"F8",X"2E",X"09",X"F0",X"0C",X"F9",X"00",X"EB",X"FB",X"3C",X"0D",X"07",X"09",
		X"CE",X"0A",X"7C",X"0A",X"FB",X"F8",X"4E",X"05",X"75",X"F8",X"B9",X"0A",X"19",X"05",X"58",X"F3",
		X"6B",X"F4",X"46",X"F5",X"62",X"F2",X"E0",X"FA",X"CC",X"03",X"0A",X"FA",X"E9",X"0C",X"40",X"0A",
		X"35",X"FE",X"87",X"FE",X"12",X"10",X"8A",X"F4",X"9C",X"0A",X"9D",X"05",X"90",X"FA",X"72",X"04",
		X"89",X"F8",X"5F",X"0F",X"A9",X"FD",X"FF",X"F3",X"C7",X"F3",X"F7",X"F5",X"73",X"F1",X"31",X"00",
		X"43",X"00",X"E9",X"FC",X"3E",X"10",X"B7",X"F6",X"D0",X"F5",X"8C",X"06",X"20",X"0B",X"8E",X"F0",
		X"A4",X"FD",X"C7",X"01",X"21",X"FC",X"B2",X"04",X"66",X"ED",X"60",X"07",X"8E",X"F9",X"DE",X"F4",
		X"23",X"F2",X"73",X"01",X"BF",X"FF",X"4B",X"F1",X"7D",X"F6",X"4F",X"04",X"32",X"FA",X"E1",X"F0",
		X"D3",X"FA",X"F5",X"08",X"F6",X"0C",X"F5",X"00",X"49",X"F3",X"7B",X"F4",X"3F",X"01",X"92",X"0E",
		X"24",X"F6",X"11",X"0A",X"67",X"FE",X"B5",X"FE",X"67",X"0E",X"C2",X"07",X"F2",X"0B",X"90",X"F6",
		X"78",X"08",X"AD",X"F2",X"83",X"F7",X"65",X"F0",X"18",X"01",X"A3",X"FF",X"AF",X"FD",X"67",X"0F",
		X"45",X"F8",X"AA",X"F4",X"4B",X"F4",X"6C",X"F5",X"5C",X"F3",X"25",X"03",X"ED",X"0C",X"C6",X"F7",
		X"95",X"06",X"F5",X"F7",X"B5",X"0B",X"A4",X"04",X"A0",X"F3",X"27",X"F5",X"B8",X"F4",X"A9",X"F4",
		X"2A",X"F5",X"53",X"F4",X"A6",X"F5",X"AD",X"F3",X"F5",X"F7",X"12",X"09",X"85",X"0C",X"07",X"F9",
		X"C5",X"05",X"35",X"F8",X"41",X"F4",X"1A",X"F4",X"E7",X"FA",X"41",X"06",X"B2",X"F0",X"81",X"F8",
		X"F0",X"F0",X"FE",X"05",X"8C",X"FB",X"11",X"F3",X"2B",X"F7",X"3C",X"07",X"DE",X"F4",X"75",X"F9",
		X"C3",X"0C",X"31",X"F8",X"10",X"07",X"46",X"F6",X"56",X"F5",X"BF",X"F3",X"B1",X"FC",X"FF",X"05",
		X"1D",X"EE",X"C6",X"06",X"F8",X"FA",X"6E",X"04",X"5A",X"FB",X"3D",X"06",X"ED",X"0A",X"B0",X"F3",
		X"94",X"F6",X"F4",X"F3",X"D9",X"F6",X"89",X"06",X"66",X"F7",X"C7",X"F3",X"10",X"FA",X"CF",X"0E",
		X"16",X"FF",X"2E",X"FF",X"AC",X"02",X"49",X"EF",X"A1",X"08",X"6B",X"09",X"8C",X"F9",X"33",X"F2",
		X"C1",X"FA",X"AF",X"09",X"DC",X"0C",X"5B",X"02",X"7A",X"F2",X"AD",X"F9",X"94",X"06",X"5C",X"F4",
		X"35",X"F5",X"4C",X"FC",X"50",X"10",X"E7",X"FA",X"B0",X"02",X"2C",X"0D",X"68",X"09",X"27",X"0B",
		X"B7",X"F4",X"3E",X"F7",X"D8",X"F1",X"54",X"FF",X"9D",X"01",X"D1",X"FD",X"B5",X"03",X"06",X"EF",
		X"21",X"FE",X"D0",X"0A",X"60",X"04",X"38",X"EF",X"FE",X"05",X"C8",X"FC",X"91",X"F3",X"BE",X"06",
		X"95",X"FA",X"EF",X"05",X"BA",X"F6",X"83",X"F4",X"38",X"F6",X"90",X"F4",X"86",X"F6",X"B0",X"F3",
		X"25",X"03",X"E5",X"0D",X"5C",X"03",X"5D",X"F2",X"BA",X"00",X"4F",X"0D",X"22",X"09",X"BD",X"0C",
		X"C2",X"F7",X"C3",X"F6",X"F9",X"08",X"C6",X"0C",X"1B",X"05",X"ED",X"F3",X"44",X"FC",X"B9",X"10",
		X"10",X"FA",X"F4",X"04",X"1E",X"FB",X"D9",X"06",X"04",X"02",X"E4",X"FD",X"98",X"02",X"E6",X"FC",
		X"8D",X"12",X"E0",X"F2",X"70",X"FB",X"3A",X"02",X"6E",X"FE",X"D8",X"01",X"D5",X"FD",X"D4",X"03",
		X"83",X"F2",X"0B",X"F7",X"3A",X"F4",X"A7",X"F6",X"29",X"F4",X"94",X"0A",X"85",X"FF",X"79",X"FE",
		X"74",X"10",X"53",X"F7",X"D7",X"07",X"4C",X"0B",X"FF",X"08",X"A3",X"F4",X"F4",X"F5",X"D4",X"F9",
		X"8D",X"10",X"2D",X"FD",X"65",X"F6",X"E3",X"F2",X"1E",X"07",X"BB",X"F9",X"AB",X"F5",X"71",X"09",
		X"AE",X"0B",X"D0",X"09",X"11",X"0C",X"BE",X"08",X"A4",X"FA",X"F6",X"06",X"8E",X"0E",X"30",X"02",
		X"54",X"FC",X"1D",X"0C",X"73",X"0A",X"5F",X"0A",X"46",X"0B",X"B7",X"09",X"82",X"0B",X"B4",X"F6",
		X"D2",X"F5",X"42",X"F4",X"B4",X"F6",X"9F",X"F3",X"DC",X"F7",X"D8",X"05",X"18",X"0F",X"64",X"02",
		X"BD",X"FD",X"26",X"03",X"30",X"F5",X"DA",X"F2",X"19",X"04",X"E8",X"FC",X"20",X"03",X"0E",X"FC",
		X"03",X"F4",X"9B",X"08",X"14",X"F8",X"DD",X"08",X"01",X"F1",X"FB",X"09",X"9A",X"F6",X"1D",X"0C",
		X"91",X"07",X"62",X"0F",X"D1",X"FE",X"77",X"00",X"D3",X"FF",X"D1",X"FF",X"DC",X"00",X"5E",X"F0",
		X"8F",X"09",X"AA",X"09",X"C3",X"0B",X"5F",X"07",X"FB",X"F2",X"79",X"FD",X"91",X"04",X"66",X"F1",
		X"E6",X"F9",X"A4",X"09",X"D3",X"0A",X"4A",X"0B",X"D4",X"02",X"3E",X"F1",X"A0",X"02",X"11",X"0D",
		X"B3",X"F9",X"97",X"05",X"FE",X"0A",X"7A",X"F7",X"E3",X"08",X"48",X"F1",X"EA",X"FE",X"4E",X"03",
		X"5C",X"F2",X"FF",X"F8",X"DA",X"0A",X"D7",X"05",X"B0",X"F2",X"78",X"F7",X"54",X"F3",X"AA",X"F7",
		X"82",X"F2",X"38",X"07",X"8D",X"09",X"C8",X"FA",X"46",X"04",X"B3",X"FB",X"7C",X"05",X"89",X"F3",
		X"BB",X"FC",X"5A",X"0F",X"4D",X"FC",X"B8",X"F5",X"88",X"F3",X"37",X"FD",X"AC",X"0C",X"3A",X"01",
		X"2E",X"F0",X"8B",X"07",X"BD",X"F9",X"D5",X"06",X"A9",X"09",X"A9",X"F7",X"86",X"F2",X"AB",X"FD",
		X"A7",X"02",X"F4",X"FC",X"A2",X"04",X"B3",X"EF",X"84",X"05",X"C1",X"0B",X"51",X"04",X"27",X"F2",
		X"4F",X"F8",X"3C",X"F2",X"7A",X"05",X"DB",X"0A",X"0A",X"0B",X"4A",X"F6",X"DA",X"F8",X"2F",X"06",
		X"DD",X"F8",X"A5",X"0E",X"1F",X"00",X"A4",X"FC",X"A3",X"10",X"87",X"F8",X"4E",X"06",X"E9",X"F8",
		X"51",X"FD",X"D3",X"0C",X"AA",X"0A",X"7F",X"FC",X"82",X"02",X"06",X"0E",X"36",X"07",X"AF",X"F7",
		X"AE",X"F4",X"FB",X"F4",X"AF",X"FB",X"98",X"0C",X"98",X"0A",X"0F",X"FF",X"E7",X"FE",X"F6",X"0F",
		X"24",X"F6",X"4F",X"F6",X"02",X"FD",X"28",X"11",X"57",X"F7",X"0B",X"07",X"87",X"09",X"C3",X"0C",
		X"3B",X"05",X"9F",X"FB",X"F8",X"04",X"76",X"F4",X"4D",X"F5",X"51",X"F6",X"5A",X"F3",X"77",X"04",
		X"01",X"FD",X"D7",X"F2",X"B9",X"09",X"D2",X"09",X"50",X"0B",X"69",X"09",X"B8",X"0B",X"AB",X"F7",
		X"18",X"F7",X"61",X"06",X"71",X"F9",X"E2",X"07",X"2A",X"F0",X"A9",X"01",X"F7",X"00",X"F7",X"F2",
		X"D9",X"F6",X"89",X"F4",X"8C",X"F6",X"14",X"07",X"41",X"0C",X"C0",X"08",X"9E",X"0C",X"41",X"F9",
		X"A6",X"05",X"2E",X"FA",X"C6",X"06",X"66",X"F4",X"3B",X"FB",X"44",X"0B",X"29",X"0B",X"F8",X"00",
		X"B1",X"F1",X"3F",X"04",X"45",X"0C",X"98",X"F8",X"F0",X"07",X"9C",X"08",X"2C",X"F8",X"EB",X"0B",
		X"28",X"09",X"EC",X"0A",X"32",X"F6",X"F9",X"F7",X"1D",X"08",X"3C",X"F1",X"F1",X"FF",X"2A",X"01",
		X"09",X"FD",X"42",X"0E",X"D1",X"07",X"31",X"0C",X"4E",X"08",X"64",X"FA",X"7D",X"05",X"81",X"F6",
		X"28",X"F5",X"A0",X"F4",X"B1",X"FC",X"9F",X"0D",X"24",X"06",X"C2",X"F5",X"15",X"F9",X"C6",X"0E",
		X"CA",X"FE",X"D1",X"FD",X"CB",X"0E",X"4D",X"FA",X"42",X"F5",X"9C",X"F4",X"D1",X"F7",X"E6",X"05",
		X"57",X"F7",X"B2",X"F2",X"50",X"FE",X"4E",X"03",X"35",X"F3",X"D6",X"F5",X"44",X"F9",X"9B",X"07",
		X"C7",X"F0",X"6F",X"00",X"E5",X"0A",X"21",X"0B",X"2E",X"FD",X"92",X"F2",X"08",X"08",X"9E",X"F8",
		X"F6",X"07",X"EE",X"F3",X"71",X"F8",X"FD",X"F0",X"66",X"02",X"7A",X"FE",X"37",X"01",X"3C",X"FF",
		X"62",X"F3",X"16",X"F5",X"0C",X"FF",X"DA",X"02",X"DD",X"F1",X"6A",X"F7",X"3A",X"03",X"C0",X"0D",
		X"4A",X"07",X"B7",X"F7",X"43",X"F7",X"9E",X"0D",X"08",X"03",X"10",X"F3",X"1C",X"00",X"20",X"0C",
		X"8A",X"0A",X"40",X"FB",X"D0",X"F9",X"D6",X"0E",X"28",X"07",X"06",X"0D",X"49",X"08",X"E1",X"FD",
		X"CE",X"F0",X"71",X"0D",X"1F",X"03",X"75",X"FE",X"EF",X"00",X"37",X"FF",X"9A",X"00",X"2A",X"FF",
		X"71",X"01",X"59",X"F2",X"8D",X"F6",X"92",X"06",X"FD",X"02",X"F9",X"FA",X"9B",X"11",X"5D",X"F7",
		X"A4",X"06",X"9B",X"09",X"BF",X"F9",X"97",X"07",X"A7",X"0C",X"19",X"04",X"F9",X"F4",X"F2",X"F4",
		X"38",X"FE",X"2C",X"0F",X"7F",X"F9",X"D4",X"04",X"08",X"FB",X"CE",X"F3",X"5B",X"F6",X"96",X"F5",
		X"C1",X"F4",X"A5",X"05",X"DB",X"FA",X"B6",X"06",X"51",X"0B",X"E9",X"0A",X"66",X"04",X"C9",X"FA",
		X"C3",X"06",X"9C",X"EE",X"72",X"05",X"06",X"09",X"52",X"0C",X"CB",X"F7",X"EC",X"F6",X"1D",X"08",
		X"33",X"0C",X"D0",X"FB",X"B6",X"F3",X"85",X"07",X"52",X"F7",X"FD",X"F7",X"5C",X"07",X"CB",X"F3",
		X"E3",X"F6",X"F0",X"F4",X"7B",X"F5",X"FF",X"FF",X"AC",X"0E",X"AE",X"F8",X"88",X"F6",X"9E",X"05",
		X"D5",X"FA",X"1D",X"06",X"A8",X"F4",X"96",X"05",X"40",X"0B",X"07",X"F7",X"11",X"F5",X"10",X"F9",
		X"5C",X"0C",X"EB",X"03",X"82",X"F1",X"08",X"03",X"87",X"FE",X"01",X"01",X"36",X"FF",X"47",X"01",
		X"DD",X"0F",X"4B",X"05",X"BD",X"0F",X"8A",X"00",X"F1",X"FD",X"94",X"09",X"69",X"0C",X"17",X"05",
		X"2A",X"FB",X"2C",X"09",X"A8",X"0C",X"45",X"00",X"28",X"F5",X"FE",X"F3",X"86",X"04",X"4D",X"FC",
		X"A9",X"03",X"73",X"0D",X"13",X"06",X"07",X"F7",X"A4",X"F4",X"6C",X"F6",X"0A",X"F5",X"ED",X"F5",
		X"6D",X"F7",X"5B",X"0B",X"77",X"09",X"0C",X"06",X"54",X"EF",X"04",X"05",X"98",X"FC",X"33",X"02",
		X"14",X"0C",X"66",X"09",X"7B",X"F7",X"93",X"F7",X"B9",X"09",X"79",X"0B",X"82",X"03",X"10",X"F4",
		X"2A",X"F6",X"CA",X"F5",X"01",X"F5",X"33",X"F7",X"BE",X"F2",X"20",X"01",X"3C",X"00",X"81",X"FE",
		X"75",X"0E",X"63",X"07",X"1F",X"0C",X"FB",X"F5",X"FC",X"F6",X"A7",X"F3",X"23",X"FC",X"B3",X"05",
		X"E0",X"F1",X"6E",X"F9",X"0C",X"F1",X"81",X"07",X"3D",X"02",X"67",X"FE",X"70",X"01",X"D3",X"FE",
		X"20",X"01",X"15",X"FF",X"CD",X"00",X"2B",X"F0",X"DF",X"0B",X"46",X"F4",X"1C",X"10",X"30",X"FF",
		X"94",X"00",X"D9",X"FF",X"B6",X"FF",X"7D",X"01",X"16",X"F2",X"4B",X"F8",X"DD",X"F3",X"FD",X"F7",
		X"F5",X"F2",X"EE",X"03",X"83",X"FE",X"90",X"F2",X"BD",X"08",X"DF",X"F6",X"FB",X"F8",X"CD",X"06",
		X"0B",X"F5",X"EE",X"F5",X"77",X"FC",X"5C",X"0F",X"44",X"FC",X"25",X"F6",X"C8",X"F4",X"8B",X"07",
		X"1B",X"0A",X"24",X"0C",X"AF",X"FD",X"96",X"F4",X"55",X"F6",X"AD",X"06",X"A8",X"0B",X"38",X"08",
		X"5C",X"F4",X"8C",X"FC",X"57",X"05",X"E5",X"F2",X"4A",X"F8",X"86",X"F3",X"24",X"04",X"E6",X"0B",
		X"71",X"09",X"A4",X"0A",X"26",X"F5",X"4C",X"02",X"B2",X"0C",X"72",X"FA",X"BF",X"F4",X"F2",X"09",
		X"ED",X"08",X"FE",X"0C",X"9D",X"02",X"6E",X"FC",X"5B",X"0B",X"91",X"0B",X"6A",X"FD",X"90",X"01",
		X"14",X"FF",X"C8",X"F1",X"4A",X"0B",X"88",X"06",X"94",X"F7",X"AB",X"F4",X"2B",X"F7",X"C7",X"F4",
		X"07",X"F8",X"84",X"09",X"34",X"07",X"D3",X"F7",X"2F",X"10",X"80",X"FD",X"24",X"00",X"B5",X"0B",
		X"F2",X"09",X"09",X"0A",X"4A",X"0A",X"98",X"F8",X"42",X"09",X"C4",X"09",X"EF",X"0A",X"F3",X"08",
		X"21",X"FB",X"CB",X"F1",X"A5",X"FC",X"15",X"02",X"65",X"FE",X"55",X"01",X"E4",X"FE",X"F6",X"00",
		X"27",X"FF",X"CD",X"00",X"33",X"FF",X"5C",X"10",X"BE",X"03",X"C5",X"FD",X"70",X"02",X"38",X"FC",
		X"14",X"0A",X"25",X"0A",X"E7",X"F6",X"2F",X"F6",X"F0",X"F4",X"61",X"FA",X"E9",X"0D",X"DF",X"FE",
		X"5F",X"FF",X"0F",X"02",X"03",X"F1",X"76",X"F9",X"A9",X"02",X"77",X"0F",X"CF",X"02",X"15",X"FE",
		X"1E",X"02",X"86",X"FC",X"3B",X"0B",X"AD",X"08",X"71",X"F7",X"2D",X"0D",X"BA",X"01",X"83",X"FC",
		X"AD",X"0B",X"3C",X"09",X"E1",X"0A",X"46",X"FD",X"B0",X"F2",X"71",X"F8",X"D4",X"F3",X"03",X"0D",
		X"BC",X"02",X"D8",X"FC",X"78",X"08",X"8D",X"0D",X"02",X"FD",X"AF",X"00",X"C3",X"0B",X"F1",X"05",
		X"7C",X"F0",X"1B",X"03",X"AC",X"FD",X"8E",X"01",X"B1",X"FE",X"EC",X"F2",X"60",X"07",X"45",X"0A",
		X"46",X"F4",X"B2",X"FB",X"25",X"04",X"1A",X"F6",X"4E",X"F3",X"E1",X"01",X"B0",X"FF",X"00",X"F4",
		X"79",X"F5",X"9C",X"FC",X"A7",X"0B",X"4F",X"0A",X"B6",X"FE",X"62",X"F3",X"33",X"F7",X"B3",X"F5",
		X"D9",X"06",X"7F",X"F9",X"60",X"07",X"F3",X"F2",X"C8",X"FD",X"98",X"0A",X"F0",X"0A",X"0D",X"FF",
		X"43",X"F3",X"BA",X"F7",X"79",X"F4",X"4E",X"F7",X"BF",X"F4",X"35",X"F7",X"E4",X"F4",X"3C",X"F7",
		X"82",X"04",X"76",X"FC",X"03",X"04",X"F4",X"F8",X"91",X"F2",X"75",X"FF",X"F4",X"02",X"8A",X"F3",
		X"D5",X"F7",X"37",X"F4",X"BC",X"05",X"86",X"FB",X"D4",X"F3",X"2A",X"F8",X"D6",X"F3",X"C3",X"04",
		X"5E",X"0B",X"FF",X"F9",X"AC",X"05",X"43",X"FA",X"04",X"0A",X"B7",X"09",X"C8",X"0B",X"4D",X"01",
		X"55",X"FC",X"51",X"10",X"BE",X"F8",X"E5",X"05",X"C1",X"FA",X"A7",X"06",X"17",X"0B",X"55",X"0A",
		X"55",X"FD",X"35",X"F3",X"0C",X"F9",X"87",X"04",X"A0",X"FB",X"0B",X"08",X"41",X"0C",X"4B",X"07",
		X"4E",X"0E",X"33",X"FC",X"C6",X"02",X"A0",X"FD",X"7F",X"02",X"42",X"FD",X"AC",X"03",X"83",X"F9",
		X"93",X"F6",X"86",X"0D",X"C8",X"F8",X"E7",X"F5",X"7E",X"F7",X"28",X"07",X"5E",X"F8",X"E6",X"0C",
		X"6C",X"07",X"B5",X"0C",X"F0",X"06",X"11",X"0E",X"4E",X"F9",X"98",X"05",X"62",X"FA",X"0B",X"07",
		X"33",X"0A",X"F9",X"0A",X"CD",X"04",X"57",X"F5",X"65",X"05",X"EF",X"FB",X"3B",X"03",X"0A",X"FD",
		X"AA",X"02",X"34",X"FD",X"FA",X"02",X"D4",X"FB",X"E9",X"0E",X"51",X"06",X"C4",X"0C",X"E6",X"06",
		X"C9",X"FA",X"24",X"F2",X"6E",X"FC",X"4D",X"04",X"2D",X"F5",X"E1",X"F6",X"B5",X"06",X"33",X"F7",
		X"F9",X"F4",X"F3",X"FA",X"F7",X"0B",X"7F",X"08",X"D2",X"0A",X"95",X"09",X"44",X"FE",X"02",X"F2",
		X"5D",X"09",X"C8",X"07",X"00",X"0D",X"E7",X"02",X"29",X"FD",X"E5",X"02",X"7D",X"FB",X"74",X"0D",
		X"AF",X"05",X"A8",X"F5",X"03",X"FB",X"C4",X"06",X"63",X"EF",X"EF",X"04",X"AD",X"FC",X"D4",X"01",
		X"1E",X"0C",X"19",X"08",X"9B",X"F9",X"8D",X"08",X"C8",X"06",X"ED",X"F7",X"DA",X"0E",X"FB",X"FD",
		X"91",X"FF",X"0D",X"02",X"1B",X"F0",X"89",X"FF",X"EF",X"01",X"A9",X"F5",X"FE",X"F3",X"6A",X"03",
		X"5B",X"FD",X"0B",X"02",X"8E",X"FD",X"AD",X"02",X"9A",X"FA",X"0B",X"F2",X"52",X"FD",X"E2",X"08",
		X"E6",X"0B",X"8B",X"FF",X"4B",X"F4",X"85",X"F6",X"90",X"02",X"77",X"0E",X"97",X"FD",X"65",X"00",
		X"DC",X"00",X"A2",X"F1",X"09",X"07",X"EA",X"09",X"C0",X"08",X"88",X"F6",X"F8",X"F5",X"07",X"F6",
		X"E3",X"F5",X"44",X"F6",X"CE",X"F5",X"FC",X"F5",X"14",X"01",X"BD",X"0E",X"97",X"F4",X"5F",X"02",
		X"16",X"FE",X"C7",X"01",X"E6",X"FD",X"85",X"02",X"FD",X"FB",X"2F",X"F5",X"DC",X"07",X"8B",X"F8",
		X"5F",X"08",X"93",X"F0",X"C8",X"01",X"63",X"01",X"17",X"F2",X"83",X"05",X"FA",X"FB",X"ED",X"F4",
		X"9F",X"F5",X"E0",X"FF",X"48",X"0C",X"EF",X"08",X"41",X"FC",X"4F",X"F3",X"A2",X"F9",X"9F",X"05",
		X"01",X"F7",X"5A",X"F5",X"82",X"FB",X"B0",X"0E",X"7C",X"FC",X"2A",X"02",X"8B",X"FE",X"3C",X"01",
		X"08",X"0E",X"BC",X"05",X"5B",X"FB",X"D9",X"07",X"43",X"0B",X"89",X"08",X"F5",X"0A",X"A8",X"08",
		X"BC",X"0A",X"11",X"09",X"FF",X"06",X"B9",X"F0",X"93",X"02",X"CC",X"FE",X"9E",X"FF",X"7C",X"0C",
		X"60",X"08",X"DB",X"FA",X"FF",X"F3",X"77",X"F7",X"22",X"F5",X"89",X"F6",X"01",X"04",X"69",X"0C",
		X"71",X"07",X"00",X"0C",X"FC",X"06",X"74",X"0D",X"8B",X"FF",X"E0",X"FE",X"4A",X"02",X"5A",X"F2",
		X"8A",X"F8",X"FB",X"F3",X"2A",X"07",X"8A",X"F8",X"E3",X"F4",X"F9",X"F9",X"C3",X"06",X"F6",X"F2",
		X"F5",X"08",X"E4",X"08",X"C3",X"08",X"3C",X"F6",X"EC",X"0F",X"1D",X"FD",X"B9",X"01",X"88",X"FE",
		X"5C",X"00",X"71",X"0B",X"8F",X"09",X"28",X"08",X"68",X"FB",X"FE",X"02",X"44",X"FD",X"12",X"02",
		X"7F",X"FD",X"FD",X"02",X"3F",X"F4",X"B3",X"F5",X"62",X"FA",X"40",X"09",X"0C",X"0C",X"C0",X"FE",
		X"E0",X"FF",X"B5",X"00",X"CD",X"F2",X"B6",X"F7",X"84",X"F5",X"9F",X"F5",X"70",X"F9",X"11",X"05",
		X"BD",X"FA",X"41",X"06",X"8F",X"F1",X"0A",X"01",X"D1",X"0B",X"5B",X"04",X"DB",X"FA",X"B8",X"06",
		X"CF",X"EF",X"D1",X"04",X"DD",X"FC",X"1D",X"02",X"2A",X"FE",X"A0",X"F2",X"DD",X"0A",X"08",X"07",
		X"4A",X"0D",X"5B",X"01",X"96",X"FD",X"E1",X"03",X"EE",X"F1",X"BF",X"02",X"83",X"0A",X"19",X"0A",
		X"12",X"03",X"06",X"FA",X"C0",X"10",X"74",X"F8",X"87",X"05",X"B7",X"FA",X"8D",X"F5",X"C3",X"F6",
		X"9B",X"08",X"A6",X"F2",X"DD",X"FE",X"59",X"01",X"4A",X"FD",X"31",X"0B",X"13",X"0A",X"29",X"FD",
		X"34",X"F4",X"55",X"F7",X"CD",X"F4",X"63",X"FF",X"BC",X"0D",X"08",X"FA",X"CE",X"F6",X"70",X"F4",
		X"02",X"FA",X"88",X"03",X"0A",X"FD",X"9C",X"02",X"3A",X"FD",X"1F",X"03",X"5A",X"FB",X"E9",X"0F",
		X"D6",X"F8",X"17",X"05",X"3B",X"FB",X"12",X"F4",X"3C",X"F8",X"99",X"F3",X"73",X"05",X"90",X"FB",
		X"77",X"F5",X"2C",X"07",X"84",X"F7",X"2D",X"F5",X"3F",X"FB",X"71",X"0B",X"72",X"08",X"5B",X"0B",
		X"C5",X"FE",X"2A",X"F3",X"28",X"06",X"E2",X"09",X"79",X"09",X"71",X"F5",X"65",X"02",X"07",X"0B",
		X"3C",X"09",X"8C",X"F9",X"2D",X"F6",X"60",X"0A",X"7E",X"05",X"DA",X"F8",X"BE",X"0E",X"6C",X"FD",
		X"E2",X"00",X"41",X"00",X"84",X"F3",X"81",X"F7",X"FF",X"04",X"76",X"0B",X"6A",X"08",X"55",X"0A",
		X"10",X"09",X"B9",X"09",X"3E",X"09",X"0F",X"F7",X"08",X"F9",X"3B",X"06",X"13",X"F5",X"19",X"F6",
		X"F5",X"FC",X"98",X"0D",X"F8",X"FC",X"51",X"F4",X"3E",X"05",X"16",X"FB",X"0A",X"F5",X"8C",X"0A",
		X"D1",X"05",X"41",X"F5",X"2B",X"05",X"68",X"FB",X"D1",X"04",X"D1",X"F7",X"DF",X"F8",X"13",X"08",
		X"47",X"F0",X"0E",X"03",X"B7",X"FE",X"58",X"FF",X"92",X"0D",X"EB",X"F8",X"2F",X"06",X"15",X"09",
		X"A5",X"F8",X"C1",X"09",X"9A",X"09",X"D4",X"04",X"5C",X"F2",X"2E",X"FB",X"FE",X"02",X"F3",X"FC",
		X"1D",X"03",X"86",X"FB",X"D5",X"0B",X"02",X"09",X"B3",X"FF",X"AC",X"F2",X"05",X"F9",X"FE",X"F3",
		X"25",X"0A",X"0F",X"07",X"29",X"0D",X"00",X"01",X"4C",X"FE",X"4F",X"02",X"21",X"F6",X"26",X"07",
		X"03",X"F6",X"3C",X"F5",X"9A",X"FD",X"1B",X"04",X"0C",X"F2",X"8E",X"F9",X"10",X"F3",X"01",X"07",
		X"D9",X"08",X"D9",X"0A",X"8A",X"07",X"7E",X"0C",X"A8",X"01",X"A5",X"FD",X"AC",X"02",X"9B",X"FB",
		X"EF",X"0E",X"3F",X"02",X"03",X"F8",X"BF",X"F3",X"1C",X"FF",X"12",X"0C",X"1A",X"FD",X"4D",X"00",
		X"E1",X"0D",X"D4",X"F5",X"F4",X"F9",X"C8",X"03",X"64",X"FB",X"4D",X"09",X"74",X"05",X"B5",X"F0",
		X"53",X"03",X"75",X"07",X"66",X"0D",X"95",X"FF",X"EC",X"FF",X"9E",X"FF",X"03",X"00",X"9E",X"FF",
		X"A5",X"FF",X"5D",X"0D",X"21",X"F7",X"AD",X"F6",X"FD",X"F5",X"29",X"F6",X"F1",X"F6",X"98",X"F4",
		X"A6",X"FE",X"A2",X"0A",X"05",X"0A",X"C6",X"FC",X"75",X"01",X"F3",X"0D",X"5F",X"FE",X"2B",X"FE",
		X"08",X"0E",X"1C",X"F9",X"50",X"05",X"22",X"FA",X"87",X"07",X"AB",X"06",X"37",X"FA",X"CD",X"05",
		X"26",X"F4",X"A2",X"F6",X"29",X"FE",X"F0",X"0C",X"97",X"06",X"E7",X"0B",X"BF",X"F7",X"4C",X"F7",
		X"F5",X"F3",X"4E",X"03",X"33",X"FE",X"18",X"F3",X"7F",X"08",X"2A",X"08",X"63",X"0B",X"E6",X"03",
		X"B7",X"FA",X"84",X"0B",X"F9",X"01",X"E5",X"F1",X"7E",X"04",X"70",X"FC",X"B5",X"02",X"7E",X"FC",
		X"40",X"F3",X"B3",X"F8",X"AB",X"F3",X"AB",X"04",X"0E",X"0A",X"24",X"09",X"38",X"09",X"BE",X"09",
		X"47",X"06",X"E1",X"F3",X"22",X"FD",X"9F",X"0B",X"F1",X"FF",X"D6",X"F2",X"62",X"04",X"D5",X"09",
		X"07",X"09",X"0F",X"F8",X"0B",X"F6",X"10",X"F6",X"BD",X"F6",X"B4",X"F5",X"C7",X"06",X"F3",X"09",
		X"5B",X"07",X"EB",X"F4",X"5A",X"F8",X"FB",X"F2",X"55",X"01",X"A5",X"FF",X"CA",X"FE",X"E3",X"0C",
		X"04",X"07",X"8D",X"0A",X"05",X"F8",X"D0",X"08",X"4F",X"09",X"E3",X"05",X"71",X"F3",X"00",X"08",
		X"92",X"F7",X"0B",X"0B",X"02",X"03",X"F9",X"FB",X"3C",X"09",X"3A",X"0B",X"AE",X"FD",X"70",X"00",
		X"E8",X"FF",X"E1",X"F1",X"EE",X"08",X"83",X"06",X"8D",X"FA",X"AC",X"05",X"6D",X"F4",X"A6",X"FC",
		X"D4",X"0A",X"6B",X"07",X"FE",X"F5",X"A0",X"FA",X"84",X"05",X"C9",X"F3",X"3F",X"F7",X"6A",X"FD",
		X"99",X"0E",X"B5",X"F8",X"2F",X"05",X"85",X"09",X"CA",X"08",X"5F",X"F5",X"02",X"FB",X"FC",X"04",
		X"91",X"F4",X"49",X"F7",X"97",X"F5",X"F0",X"F6",X"BE",X"F5",X"20",X"F7",X"0B",X"F5",X"FA",X"FD",
		X"FE",X"0C",X"FF",X"FB",X"72",X"01",X"5D",X"0C",X"E6",X"F7",X"6E",X"07",X"68",X"F5",X"BF",X"FB",
		X"9C",X"03",X"81",X"FB",X"C8",X"05",X"01",X"F0",X"92",X"05",X"F1",X"03",X"45",X"FB",X"A8",X"0A",
		X"D7",X"08",X"EA",X"08",X"89",X"0A",X"9F",X"FB",X"DD",X"02",X"C1",X"FC",X"16",X"04",X"63",X"0C",
		X"3C",X"06",X"16",X"0C",X"AF",X"05",X"BD",X"0D",X"95",X"FB",X"71",X"02",X"AF",X"FD",X"ED",X"F4",
		X"75",X"F5",X"04",X"FF",X"93",X"02",X"19",X"F1",X"56",X"06",X"CE",X"FA",X"7A",X"F5",X"66",X"08",
		X"CD",X"06",X"7B",X"F8",X"74",X"0C",X"7D",X"00",X"BF",X"FC",X"FA",X"0B",X"0D",X"07",X"1C",X"0B",
		X"74",X"FA",X"B0",X"F4",X"D8",X"FD",X"E9",X"0C",X"FF",X"FB",X"B6",X"F5",X"3F",X"F6",X"A9",X"F6",
		X"BB",X"F5",X"88",X"F8",X"46",X"0A",X"B8",X"03",X"CC",X"F9",X"4D",X"0E",X"DE",X"FC",X"07",X"F7",
		X"58",X"F4",X"E4",X"05",X"15",X"FA",X"16",X"07",X"07",X"01",X"2D",X"F2",X"B3",X"05",X"71",X"FB",
		X"7B",X"03",X"19",X"FC",X"06",X"04",X"0D",X"F8",X"76",X"F4",X"14",X"FD",X"87",X"0B",X"EA",X"FF",
		X"2D",X"F3",X"1F",X"04",X"1A",X"0A",X"E4",X"F9",X"EF",X"F4",X"E7",X"F7",X"82",X"F4",X"3B",X"04",
		X"0B",X"0A",X"12",X"FA",X"C4",X"04",X"85",X"FA",X"8F",X"08",X"09",X"0A",X"B5",X"03",X"69",X"F2",
		X"75",X"02",X"79",X"FF",X"E4",X"F3",X"F7",X"F7",X"FA",X"F5",X"97",X"06",X"4F",X"F9",X"43",X"09",
		X"30",X"09",X"76",X"FB",X"64",X"F4",X"4E",X"F8",X"82",X"F4",X"89",X"FB",X"D8",X"05",X"57",X"F2",
		X"C8",X"01",X"6D",X"FF",X"B7",X"FF",X"DE",X"00",X"BE",X"F1",X"82",X"FA",X"DE",X"F2",X"28",X"FC",
		X"C9",X"03",X"C1",X"F7",X"74",X"F5",X"EC",X"F7",X"72",X"F6",X"01",X"0B",X"93",X"04",X"2F",X"F6",
		X"A5",X"FB",X"EB",X"0D",X"5F",X"FD",X"05",X"F7",X"3E",X"F5",X"CA",X"05",X"1A",X"09",X"70",X"FA",
		X"32",X"05",X"0D",X"FA",X"29",X"0B",X"23",X"03",X"B6",X"F4",X"38",X"F9",X"23",X"08",X"EE",X"09",
		X"DA",X"08",X"9E",X"09",X"10",X"09",X"31",X"09",X"EB",X"09",X"32",X"FD",X"3E",X"F4",X"10",X"07",
		X"5B",X"F9",X"99",X"08",X"AE",X"08",X"8F",X"0A",X"07",X"03",X"D4",X"F4",X"A8",X"F7",X"01",X"F6",
		X"BE",X"F6",X"6A",X"FA",X"97",X"0C",X"F5",X"05",X"74",X"0D",X"5F",X"FA",X"50",X"04",X"CD",X"FB",
		X"22",X"04",X"42",X"FB",X"71",X"05",X"96",X"F8",X"7C",X"0D",X"B9",X"FE",X"9E",X"00",X"33",X"FF",
		X"A7",X"00",X"84",X"06",X"AD",X"FA",X"D1",X"04",X"36",X"FA",X"60",X"0E",X"65",X"05",X"0E",X"0C",
		X"A8",X"06",X"98",X"0A",X"C6",X"F7",X"F7",X"07",X"E6",X"F3",X"ED",X"FC",X"1F",X"09",X"4A",X"09",
		X"3C",X"09",X"FC",X"FF",X"F3",X"F1",X"0A",X"FF",X"A6",X"02",X"2D",X"F4",X"CF",X"FF",X"D3",X"0C",
		X"D0",X"F9",X"AB",X"04",X"6D",X"FA",X"9A",X"F6",X"78",X"07",X"CF",X"F4",X"C3",X"FB",X"0C",X"0B",
		X"74",X"01",X"10",X"F4",X"B6",X"F8",X"12",X"F4",X"44",X"06",X"66",X"F9",X"14",X"FD",X"2B",X"0D",
		X"36",X"FC",X"E2",X"F5",X"FB",X"F6",X"35",X"05",X"0E",X"FA",X"2D",X"F4",X"1B",X"FC",X"C1",X"04",
		X"E5",X"F4",X"09",X"F8",X"15",X"F5",X"53",X"01",X"19",X"0C",X"ED",X"F9",X"3A",X"05",X"75",X"0A",
		X"37",X"08",X"4B",X"0A",X"96",X"FC",X"77",X"F4",X"F3",X"07",X"22",X"08",X"1A",X"0B",X"7E",X"03",
		X"AA",X"FB",X"9F",X"09",X"5D",X"0A",X"CE",X"FE",X"E8",X"FE",X"F3",X"0C",X"7B",X"F9",X"8B",X"F6",
		X"C9",X"06",X"2D",X"F6",X"DC",X"02",X"B8",X"FD",X"BC",X"01",X"CC",X"FD",X"74",X"02",X"B2",X"FA",
		X"FE",X"F2",X"3F",X"FE",X"A0",X"03",X"5E",X"F3",X"26",X"01",X"07",X"0A",X"66",X"09",X"36",X"FB",
		X"70",X"04",X"AA",X"09",X"F8",X"F7",X"3E",X"0A",X"AB",X"07",X"1E",X"0A",X"78",X"F8",X"5F",X"F7",
		X"7D",X"09",X"21",X"05",X"F5",X"F5",X"A5",X"F6",X"59",X"F7",X"BE",X"F4",X"08",X"03",X"E1",X"FD",
		X"6E",X"01",X"60",X"0C",X"68",X"F5",X"F1",X"FA",X"38",X"04",X"61",X"FA",X"3E",X"0B",X"42",X"F8",
		X"8C",X"07",X"CF",X"F4",X"48",X"FD",X"01",X"02",X"CC",X"FD",X"1D",X"02",X"CB",X"FC",X"E6",X"0C",
		X"FC",X"06",X"38",X"FD",X"1E",X"F4",X"37",X"08",X"93",X"F7",X"9F",X"0B",X"B4",X"02",X"E2",X"F6",
		X"DB",X"F5",X"09",X"F9",X"25",X"06",X"6D",X"F5",X"80",X"FC",X"46",X"05",X"CE",X"F1",X"DB",X"02",
		X"9A",X"08",X"A0",X"0A",X"EF",X"F9",X"CA",X"05",X"8A",X"08",X"8D",X"F7",X"A1",X"F5",X"A5",X"FB",
		X"D9",X"09",X"A1",X"09",X"84",X"00",X"79",X"F4",X"8F",X"F7",X"3A",X"FA",X"24",X"0C",X"85",X"06",
		X"40",X"0B",X"A0",X"06",X"A1",X"0B",X"18",X"F9",X"B6",X"F7",X"F5",X"05",X"1C",X"0B",X"5F",X"06",
		X"72",X"0C",X"A6",X"FF",X"3C",X"FE",X"B9",X"09",X"EB",X"09",X"86",X"03",X"E2",X"FB",X"89",X"04",
		X"7E",X"F3",X"04",X"F8",X"2A",X"FF",X"99",X"0D",X"A6",X"F7",X"60",X"07",X"0A",X"07",X"05",X"F8",
		X"C9",X"F7",X"29",X"0D",X"17",X"FF",X"89",X"FE",X"89",X"09",X"CF",X"09",X"92",X"FC",X"D9",X"F4",
		X"40",X"FC",X"5C",X"0D",X"9B",X"FB",X"6F",X"02",X"AD",X"FD",X"BB",X"F4",X"2C",X"F7",X"E3",X"F7",
		X"98",X"07",X"A5",X"0A",X"50",X"02",X"63",X"FC",X"95",X"04",X"52",X"F1",X"70",X"04",X"96",X"FD",
		X"00",X"F4",X"E5",X"07",X"2B",X"01",X"5A",X"F4",X"4D",X"F8",X"15",X"F5",X"63",X"05",X"00",X"FB",
		X"AF",X"05",X"83",X"0A",X"5D",X"07",X"4F",X"0A",X"EF",X"06",X"95",X"0B",X"A8",X"FD",X"70",X"FF",
		X"63",X"0C",X"2B",X"F9",X"49",X"05",X"93",X"F8",X"9A",X"FE",X"28",X"0C",X"1F",X"06",X"0D",X"0B",
		X"EC",X"05",X"79",X"FA",X"9A",X"F3",X"E5",X"F9",X"55",X"F2",X"DB",X"00",X"BB",X"FF",X"1F",X"FE",
		X"0E",X"0C",X"B5",X"FB",X"2D",X"F5",X"EE",X"F7",X"38",X"F5",X"BC",X"F9",X"E5",X"07",X"77",X"09",
		X"FC",X"07",X"41",X"FA",X"DC",X"F5",X"62",X"0A",X"62",X"06",X"D9",X"0B",X"7A",X"00",X"F6",X"F6",
		X"E9",X"F4",X"E7",X"01",X"6B",X"0A",X"21",X"FB",X"D4",X"F4",X"6B",X"F8",X"AE",X"F4",X"24",X"FB",
		X"AD",X"08",X"E8",X"FB",X"41",X"F4",X"B8",X"0A",X"2B",X"03",X"3D",X"FD",X"57",X"02",X"39",X"FC",
		X"68",X"0A",X"E2",X"08",X"DD",X"FE",X"C9",X"F3",X"75",X"05",X"AA",X"09",X"CD",X"06",X"DB",X"F9",
		X"3A",X"08",X"9C",X"09",X"20",X"03",X"E7",X"F4",X"47",X"09",X"23",X"05",X"B6",X"F9",X"32",X"0B",
		X"4C",X"01",X"F2",X"F5",X"BE",X"F5",X"F7",X"01",X"A2",X"FE",X"3C",X"00",X"2F",X"0D",X"D0",X"F3",
		X"C1",X"FC",X"D3",X"01",X"C9",X"FC",X"23",X"08",X"19",X"0A",X"76",X"06",X"BC",X"0B",X"C4",X"01",
		X"C5",X"FC",X"38",X"08",X"A7",X"0A",X"1B",X"FE",X"02",X"F6",X"28",X"F6",X"D1",X"F7",X"0C",X"03",
		X"75",X"FD",X"21",X"01",X"87",X"FE",X"78",X"00",X"E5",X"FE",X"7A",X"00",X"0E",X"FE",X"75",X"0A",
		X"F5",X"08",X"E4",X"02",X"17",X"FB",X"9A",X"0B",X"7B",X"06",X"83",X"0A",X"C4",X"FB",X"07",X"F5",
		X"20",X"06",X"1C",X"F9",X"A9",X"08",X"C6",X"04",X"63",X"F6",X"21",X"F6",X"D9",X"F7",X"29",X"F4",
		X"2D",X"03",X"14",X"FD",X"59",X"F9",X"84",X"0B",X"35",X"07",X"D8",X"01",X"41",X"F1",X"ED",X"06",
		X"81",X"F9",X"13",X"06",X"2A",X"08",X"28",X"0A",X"58",X"03",X"47",X"FB",X"44",X"09",X"54",X"09",
		X"B2",X"FF",X"AA",X"F4",X"8A",X"F7",X"53",X"F6",X"80",X"F6",X"7E",X"F7",X"B4",X"F4",X"32",X"03",
		X"26",X"FD",X"E8",X"01",X"9C",X"0B",X"66",X"05",X"97",X"F8",X"A4",X"F5",X"81",X"F7",X"34",X"F6",
		X"21",X"F7",X"A2",X"F6",X"C3",X"F6",X"27",X"F7",X"2E",X"F6",X"1F",X"F8",X"60",X"F4",X"81",X"02",
		X"50",X"FE",X"A3",X"00",X"DC",X"0B",X"C8",X"06",X"CE",X"08",X"CB",X"F7",X"EA",X"0A",X"02",X"06",
		X"1F",X"0C",X"4E",X"FE",X"F5",X"FE",X"D8",X"0A",X"41",X"07",X"9F",X"09",X"54",X"F9",X"D2",X"F6",
		X"22",X"09",X"E8",X"FD",X"44",X"F4",X"BD",X"05",X"F9",X"08",X"5E",X"08",X"E0",X"08",X"D9",X"05",
		X"EC",X"F3",X"AD",X"FE",X"F4",X"02",X"86",X"F2",X"4B",X"03",X"B2",X"08",X"11",X"09",X"93",X"F9",
		X"74",X"06",X"79",X"08",X"AA",X"09",X"37",X"FB",X"36",X"03",X"4F",X"FB",X"CF",X"F4",X"A0",X"F7",
		X"C7",X"F8",X"68",X"0B",X"98",X"01",X"3F",X"F4",X"1F",X"01",X"3E",X"00",X"4A",X"F3",X"5F",X"F9",
		X"6C",X"02",X"73",X"FD",X"0A",X"02",X"6E",X"FC",X"60",X"07",X"B4",X"09",X"D8",X"F8",X"5D",X"06",
		X"77",X"F6",X"10",X"F8",X"DA",X"F4",X"99",X"FD",X"A2",X"0A",X"94",X"FF",X"3B",X"F4",X"0D",X"F9",
		X"A9",X"F4",X"CC",X"07",X"23",X"06",X"E3",X"FA",X"14",X"07",X"8D",X"0A",X"F0",X"01",X"B5",X"F5",
		X"5F",X"F8",X"7A",X"08",X"01",X"08",X"30",X"09",X"B7",X"07",X"4F",X"09",X"95",X"07",X"42",X"09",
		X"DC",X"07",X"67",X"FC",X"31",X"F4",X"BD",X"08",X"09",X"F4",X"A6",X"FD",X"64",X"01",X"0B",X"FD",
		X"C5",X"08",X"D4",X"09",X"D0",X"03",X"27",X"FC",X"7A",X"03",X"35",X"F6",X"4C",X"F5",X"58",X"01",
		X"66",X"FF",X"6D",X"F4",X"D7",X"F7",X"43",X"05",X"FA",X"07",X"5F",X"F9",X"00",X"06",X"4E",X"F5",
		X"34",X"F7",X"A7",X"FC",X"D5",X"0B",X"22",X"06",X"16",X"08",X"45",X"F1",X"23",X"02",X"3C",X"FE",
		X"68",X"00",X"C6",X"FF",X"24",X"F4",X"66",X"F8",X"6A",X"04",X"85",X"0A",X"74",X"05",X"6B",X"F6",
		X"76",X"FB",X"B4",X"05",X"56",X"F1",X"C4",X"03",X"6E",X"FD",X"88",X"00",X"1C",X"0C",X"8B",X"00",
		X"4D",X"F6",X"45",X"F6",X"13",X"01",X"F0",X"0A",X"95",X"06",X"29",X"0A",X"85",X"06",X"CE",X"0A",
		X"F6",X"02",X"1F",X"FB",X"B0",X"0A",X"52",X"00",X"F5",X"FB",X"A5",X"0E",X"58",X"F7",X"93",X"07",
		X"1B",X"FF",X"FF",X"FF",X"01",X"FF",X"3E",X"00",X"A8",X"FE",X"B6",X"00",X"F9",X"FD",X"E1",X"01",
		X"A6",X"FA",X"98",X"F3",X"2E",X"FD",X"94",X"08",X"43",X"08",X"F8",X"08",X"DB",X"FE",X"92",X"F3",
		X"A1",X"05",X"A6",X"FA",X"F2",X"04",X"B7",X"0A",X"A9",X"FC",X"C1",X"F5",X"17",X"F7",X"86",X"F7",
		X"7D",X"05",X"C2",X"F7",X"93",X"F8",X"5C",X"0C",X"9F",X"FE",X"CD",X"FF",X"B8",X"FF",X"3B",X"FF",
		X"6A",X"00",X"80",X"F2",X"83",X"FA",X"8A",X"03",X"4D",X"0C",X"42",X"FB",X"19",X"F7",X"0F",X"F6",
		X"A1",X"F8",X"7F",X"04",X"77",X"FA",X"C5",X"08",X"55",X"04",X"76",X"F4",X"39",X"F9",X"F5",X"F3",
		X"8B",X"03",X"94",X"FD",X"F6",X"F4",X"3B",X"06",X"48",X"09",X"11",X"06",X"3C",X"F7",X"73",X"F6",
		X"88",X"04",X"5D",X"FB",X"82",X"05",X"9D",X"09",X"2E",X"08",X"50",X"04",X"12",X"F9",X"D2",X"0E",
		X"43",X"FA",X"72",X"03",X"C4",X"FC",X"0E",X"F6",X"03",X"F7",X"F0",X"07",X"2B",X"05",X"35",X"FB",
		X"B2",X"04",X"59",X"F5",X"94",X"F7",X"1F",X"F8",X"83",X"06",X"38",X"F5",X"59",X"FC",X"D2",X"09",
		X"21",X"07",X"65",X"0A",X"B8",X"FC",X"EB",X"00",X"6D",X"0B",X"BB",X"F7",X"0E",X"F8",X"39",X"F5",
		X"C0",X"FB",X"86",X"04",X"16",X"F5",X"36",X"F9",X"57",X"04",X"E4",X"FA",X"E1",X"07",X"AF",X"09",
		X"98",X"01",X"9A",X"FB",X"92",X"0D",X"D5",X"FA",X"0A",X"F8",X"39",X"F5",X"D1",X"07",X"6A",X"05",
		X"33",X"FC",X"B3",X"02",X"A7",X"FC",X"A4",X"03",X"25",X"F5",X"7E",X"F7",X"61",X"F9",X"61",X"06",
		X"DE",X"F3",X"C6",X"FE",X"05",X"09",X"FA",X"08",X"90",X"FE",X"6B",X"F4",X"4A",X"F9",X"3C",X"F5",
		X"BD",X"09",X"9B",X"03",X"F3",X"FC",X"AA",X"02",X"E8",X"FB",X"85",X"0A",X"41",X"07",X"64",X"09",
		X"F9",X"04",X"26",X"F5",X"38",X"F9",X"F3",X"F3",X"D7",X"02",X"67",X"FE",X"A9",X"F5",X"83",X"F7",
		X"70",X"05",X"B9",X"F8",X"44",X"F9",X"18",X"06",X"F0",X"F4",X"37",X"FD",X"46",X"0B",X"BB",X"FE",
		X"57",X"F6",X"B4",X"F6",X"FD",X"FB",X"FF",X"09",X"43",X"08",X"DC",X"00",X"0A",X"F3",X"E1",X"05",
		X"23",X"FB",X"32",X"04",X"18",X"FB",X"38",X"07",X"95",X"06",X"25",X"F4",X"B5",X"FE",X"8C",X"08",
		X"E0",X"09",X"4F",X"FD",X"F5",X"00",X"80",X"FF",X"A4",X"F1",X"33",X"03",X"AC",X"FE",X"9C",X"F6",
		X"83",X"F6",X"37",X"05",X"A1",X"08",X"6A",X"09",X"CA",X"04",X"7C",X"FB",X"E0",X"04",X"24",X"F5",
		X"73",X"F8",X"80",X"F6",X"B8",X"F7",X"2C",X"F7",X"21",X"F7",X"53",X"05",X"BE",X"F9",X"E7",X"F6",
		X"A3",X"F6",X"C3",X"03",X"D3",X"FC",X"D1",X"03",X"C1",X"09",X"EA",X"F5",X"92",X"F8",X"96",X"F9",
		X"4C",X"0D",X"45",X"FE",X"56",X"F8",X"0A",X"F5",X"E5",X"04",X"13",X"FC",X"3F",X"F6",X"EC",X"F7",
		X"3E",X"F7",X"A6",X"F7",X"22",X"F7",X"9B",X"04",X"C8",X"09",X"75",X"F7",X"78",X"F8",X"57",X"F6",
		X"EA",X"F8",X"ED",X"F5",X"A8",X"F9",X"7B",X"F4",X"65",X"04",X"5F",X"FD",X"95",X"F6",X"73",X"F7",
		X"8A",X"F9",X"24",X"05",X"04",X"FB",X"72",X"09",X"50",X"08",X"08",X"FB",X"37",X"05",X"2A",X"FA",
		X"AF",X"0A",X"1E",X"02",X"4A",X"FD",X"AE",X"04",X"27",X"F2",X"BB",X"05",X"3E",X"FC",X"82",X"03",
		X"EC",X"FC",X"8B",X"04",X"99",X"0B",X"CA",X"03",X"5F",X"F8",X"6E",X"F6",X"DD",X"F9",X"27",X"04",
		X"9D",X"FC",X"07",X"04",X"1F",X"FB",X"DD",X"0B",X"47",X"00",X"27",X"F6",X"C2",X"F8",X"54",X"F6",
		X"5E",X"05",X"48",X"09",X"F2",X"08",X"70",X"06",X"BC",X"F9",X"76",X"0B",X"A2",X"01",X"AE",X"F7",
		X"30",X"07",X"16",X"0A",X"00",X"04",X"30",X"FB",X"31",X"0B",X"94",X"06",X"05",X"0B",X"44",X"FD",
		X"95",X"F6",X"FA",X"F7",X"6F",X"F7",X"91",X"F7",X"16",X"F9",X"55",X"0A",X"07",X"03",X"82",X"FB",
		X"9C",X"0C",X"26",X"FE",X"01",X"F9",X"2D",X"0A",X"D1",X"03",X"0A",X"F5",X"EB",X"FF",X"EF",X"09",
		X"68",X"08",X"03",X"FE",X"B2",X"F4",X"72",X"08",X"BD",X"05",X"0A",X"FC",X"82",X"04",X"7C",X"F7",
		X"2D",X"F7",X"A0",X"F8",X"A9",X"F5",X"C8",X"02",X"A2",X"06",X"08",X"F5",X"42",X"FE",X"46",X"0B",
		X"D2",X"FE",X"65",X"F6",X"33",X"F8",X"91",X"F7",X"76",X"F7",X"53",X"F9",X"39",X"06",X"20",X"F7",
		X"A3",X"F8",X"53",X"F6",X"DD",X"FE",X"61",X"0B",X"76",X"FE",X"24",X"F5",X"C1",X"06",X"28",X"02",
		X"5E",X"FD",X"A6",X"04",X"06",X"F1",X"D5",X"08",X"BF",X"F8",X"81",X"08",X"FD",X"04",X"B6",X"FD",
		X"22",X"02",X"86",X"FE",X"36",X"02",X"30",X"FD",X"F2",X"0B",X"30",X"FE",X"7F",X"F5",X"54",X"FA",
		X"06",X"F4",X"37",X"03",X"2B",X"FE",X"38",X"02",X"40",X"FE",X"A5",X"02",X"E0",X"FC",X"85",X"F5",
		X"4F",X"F9",X"0B",X"F7",X"EE",X"F7",X"7B",X"FC",X"89",X"0C",X"8A",X"FE",X"47",X"F7",X"AD",X"F7",
		X"2D",X"04",X"53",X"FD",X"E5",X"F3",X"0D",X"04",X"9A",X"FE",X"A2",X"F6",X"38",X"F8",X"E8",X"F8",
		X"BA",X"05",X"AE",X"F9",X"FA",X"F5",X"51",X"FE",X"FF",X"03",X"CF",X"F5",X"50",X"F9",X"3B",X"F7",
		X"B4",X"F8",X"99",X"F7",X"F3",X"F8",X"14",X"06",X"51",X"F9",X"CD",X"F7",X"43",X"F8",X"40",X"F8",
		X"EF",X"F7",X"C1",X"F8",X"0B",X"F7",X"92",X"FC",X"C2",X"05",X"8B",X"F5",X"97",X"FA",X"54",X"F5",
		X"85",X"04",X"81",X"FE",X"7D",X"F6",X"87",X"06",X"CE",X"FB",X"CB",X"05",X"C0",X"F8",X"C5",X"F7",
		X"63",X"05",X"BD",X"FC",X"E1",X"04",X"87",X"FB",X"5F",X"0A",X"43",X"03",X"34",X"FD",X"CF",X"05",
		X"3B",X"F2",X"D2",X"06",X"7B",X"FC",X"5F",X"F8",X"BF",X"F7",X"53",X"09",X"84",X"05",X"C3",X"FC",
		X"61",X"05",X"AF",X"F6",X"BA",X"F9",X"BB",X"07",X"C9",X"07",X"75",X"F6",X"A2",X"FD",X"74",X"0A",
		X"EF",X"07",X"EB",X"0A",X"DC",X"FD",X"D5",X"01",X"2E",X"0C",X"A3",X"F8",X"C4",X"F9",X"FD",X"F5",
		X"DD",X"FD",X"B4",X"03",X"95",X"FC",X"C9",X"0B",X"F3",X"05",X"65",X"FB",X"0C",X"0A",X"57",X"04",
		X"27",X"F6",X"84",X"FF",X"82",X"0C",X"61",X"FC",X"BD",X"03",X"CE",X"FD",X"38",X"04",X"5A",X"0A",
		X"CF",X"F6",X"02",X"FA",X"93",X"F6",X"38",X"FA",X"C8",X"F5",X"DD",X"01",X"29",X"0A",X"49",X"06",
		X"08",X"F5",X"2B",X"01",X"83",X"01",X"65",X"FE",X"62",X"0D",X"2A",X"FB",X"A2",X"F8",X"8C",X"05",
		X"27",X"0B",X"7D",X"05",X"F7",X"F8",X"9A",X"FA",X"E3",X"0D",X"AC",X"FD",X"8E",X"02",X"2F",X"FF",
		X"D5",X"FA",X"55",X"06",X"95",X"F5",X"6D",X"F9",X"06",X"FF",X"92",X"0D",X"4E",X"FA",X"DA",X"05",
		X"9D",X"08",X"41",X"FB",X"21",X"06",X"E5",X"F7",X"FE",X"F8",X"73",X"F7",X"AF",X"F9",X"06",X"F6",
		X"13",X"04",X"AA",X"FE",X"03",X"F7",X"FD",X"F7",X"19",X"00",X"47",X"03",X"AA",X"F3",X"D5",X"06",
		X"3D",X"08",X"58",X"0A",X"6E",X"06",X"A6",X"FB",X"F9",X"08",X"B7",X"08",X"E1",X"09",X"66",X"02",
		X"42",X"F5",X"25",X"03",X"6D",X"0A",X"7B",X"07",X"5A",X"0B",X"40",X"FF",X"BC",X"00",X"73",X"01",
		X"AB",X"F4",X"FA",X"FA",X"25",X"04",X"F0",X"0B",X"02",X"06",X"43",X"0C",X"7E",X"01",X"E9",X"FD",
		X"EA",X"0A",X"B4",X"00",X"D3",X"F4",X"C9",X"05",X"76",X"FC",X"C9",X"04",X"DF",X"09",X"81",X"F6",
		X"F6",X"03",X"A8",X"FE",X"8A",X"F5",X"36",X"FB",X"E2",X"03",X"92",X"FD",X"AE",X"03",X"ED",X"FC",
		X"98",X"05",X"CC",X"F3",X"21",X"03",X"DB",X"08",X"6A",X"09",X"EA",X"07",X"05",X"0A",X"4E",X"06",
		X"C7",X"FB",X"DF",X"07",X"9B",X"09",X"90",X"07",X"10",X"FC",X"37",X"F5",X"61",X"FD",X"8C",X"03",
		X"75",X"F9",X"61",X"F5",X"51",X"02",X"AF",X"FF",X"75",X"00",X"20",X"0B",X"99",X"07",X"AD",X"FB",
		X"EE",X"F6",X"F8",X"F8",X"E4",X"F7",X"5D",X"F8",X"85",X"F8",X"A0",X"F7",X"98",X"FA",X"BB",X"05",
		X"81",X"F8",X"6B",X"F7",X"27",X"FE",X"B8",X"0A",X"B2",X"07",X"A2",X"09",X"1A",X"08",X"5D",X"09",
		X"32",X"08",X"45",X"09",X"24",X"08",X"52",X"09",X"ED",X"07",X"A4",X"09",X"C2",X"06",X"E9",X"FB",
		X"83",X"06",X"43",X"0B",X"57",X"01",X"B6",X"FE",X"0F",X"03",X"A3",X"F5",X"DB",X"F8",X"AC",X"02",
		X"DC",X"FE",X"2C",X"02",X"2B",X"0D",X"4E",X"02",X"ED",X"FE",X"E8",X"01",X"6B",X"FE",X"37",X"03",
		X"E0",X"F6",X"75",X"08",X"08",X"F5",X"8F",X"FB",X"BA",X"F3",X"C9",X"03",X"EA",X"FD",X"A7",X"02",
		X"1F",X"FE",X"EC",X"02",X"55",X"FD",X"3A",X"05",X"0F",X"0A",X"E5",X"07",X"83",X"08",X"C2",X"09",
		X"C8",X"00",X"13",X"FE",X"01",X"0C",X"F0",X"05",X"C4",X"0A",X"01",X"06",X"C6",X"0B",X"DF",X"FC",
		X"5E",X"02",X"A3",X"FE",X"87",X"01",X"18",X"FF",X"4F",X"01",X"16",X"FF",X"A2",X"01",X"02",X"FE",
		X"92",X"07",X"FE",X"0A",X"92",X"FD",X"C1",X"01",X"5B",X"FF",X"62",X"F5",X"BD",X"F9",X"AF",X"F6",
		X"72",X"F9",X"37",X"F6",X"AD",X"04",X"EF",X"FC",X"54",X"03",X"F3",X"FC",X"B7",X"05",X"01",X"0B",
		X"37",X"02",X"54",X"FC",X"31",X"0C",X"7C",X"FD",X"74",X"01",X"C2",X"FF",X"17",X"00",X"13",X"0E",
		X"8F",X"FC",X"A7",X"01",X"CB",X"08",X"05",X"09",X"2C",X"FB",X"62",X"F7",X"31",X"F8",X"23",X"F8",
		X"9B",X"F7",X"96",X"FB",X"EC",X"0B",X"A8",X"FE",X"6D",X"00",X"23",X"01",X"C1",X"F4",X"4F",X"FA",
		X"89",X"F6",X"DA",X"F8",X"ED",X"FE",X"D6",X"0C",X"24",X"FA",X"28",X"F9",X"0F",X"F7",X"68",X"09",
		X"5C",X"04",X"3B",X"FC",X"77",X"08",X"55",X"09",X"C3",X"01",X"19",X"F5",X"04",X"03",X"41",X"09",
		X"1D",X"08",X"70",X"FB",X"17",X"05",X"C9",X"F8",X"48",X"01",X"21",X"0B",X"1F",X"FA",X"5F",X"F8",
		X"BE",X"07",X"EC",X"05",X"7D",X"FA",X"35",X"0A",X"06",X"07",X"2D",X"09",X"24",X"08",X"EB",X"FF",
		X"75",X"F4",X"B7",X"06",X"82",X"FA",X"B5",X"06",X"73",X"08",X"4F",X"08",X"40",X"08",X"1F",X"FC",
		X"C8",X"F5",X"6B",X"FB",X"F4",X"03",X"B6",X"FB",X"F5",X"08",X"6A",X"08",X"68",X"02",X"DD",X"F3",
		X"C2",X"04",X"E0",X"FC",X"E8",X"02",X"7A",X"0A",X"8F",X"05",X"2C",X"FB",X"12",X"08",X"FD",X"07",
		X"8B",X"08",X"7F",X"07",X"41",X"09",X"EF",X"04",X"90",X"F8",X"5D",X"F6",X"8D",X"FE",X"B2",X"08",
		X"41",X"09",X"43",X"FD",X"DC",X"01",X"4D",X"FE",X"32",X"F5",X"5A",X"09",X"68",X"04",X"42",X"FB",
		X"98",X"09",X"71",X"02",X"5D",X"F6",X"8F",X"F8",X"5B",X"F9",X"96",X"09",X"B3",X"06",X"7B",X"09",
		X"6B",X"06",X"74",X"0A",X"70",X"FC",X"F6",X"01",X"1A",X"0A",X"23",X"F9",X"02",X"F8",X"99",X"F7",
		X"4A",X"F8",X"7D",X"F7",X"83",X"F8",X"25",X"F7",X"09",X"FA",X"45",X"07",X"E5",X"08",X"E0",X"06",
		X"4E",X"0A",X"EE",X"FE",X"BD",X"FF",X"74",X"01",X"5F",X"F3",X"76",X"07",X"74",X"F9",X"EE",X"06",
		X"30",X"F6",X"B3",X"FD",X"37",X"02",X"1A",X"FD",X"0A",X"09",X"19",X"09",X"74",X"FD",X"0E",X"FB",
		X"55",X"04",X"76",X"FB",X"A5",X"05",X"87",X"F1",X"18",X"06",X"FD",X"05",X"B3",X"0A",X"62",X"04",
		X"FE",X"FD",X"51",X"01",X"D6",X"FE",X"1E",X"01",X"83",X"FE",X"62",X"02",X"C7",X"F5",X"EF",X"F8",
		X"90",X"F7",X"FD",X"F7",X"72",X"F8",X"C3",X"F6",X"C5",X"00",X"D9",X"09",X"F6",X"06",X"E9",X"08",
		X"79",X"F9",X"45",X"F9",X"B7",X"05",X"64",X"F9",X"FF",X"0B",X"F7",X"FE",X"14",X"00",X"A8",X"00",
		X"49",X"FE",X"9A",X"0C",X"7E",X"F8",X"4F",X"FE",X"01",X"0A",X"79",X"FF",X"2D",X"F5",X"B1",X"04",
		X"2E",X"08",X"7A",X"08",X"32",X"06",X"0C",X"F9",X"80",X"F6",X"5D",X"FD",X"44",X"04",X"23",X"F4",
		X"FE",X"01",X"83",X"08",X"03",X"08",X"BD",X"07",X"50",X"08",X"55",X"07",X"20",X"09",X"CE",X"FD",
		X"34",X"F6",X"11",X"F9",X"7A",X"F7",X"0D",X"07",X"29",X"F6",X"9F",X"FD",X"62",X"02",X"B8",X"FC",
		X"91",X"09",X"3A",X"08",X"15",X"FE",X"E5",X"00",X"37",X"FF",X"F7",X"F3",X"78",X"FB",X"13",X"F4",
		X"29",X"05",X"3B",X"FC",X"A3",X"F7",X"D5",X"04",X"7E",X"FB",X"DD",X"06",X"67",X"06",X"4B",X"F4",
		X"C4",X"00",X"9D",X"00",X"D0",X"FD",X"49",X"0C",X"37",X"FA",X"7C",X"04",X"C3",X"FB",X"AE",X"04",
		X"B8",X"F8",X"8A",X"FA",X"13",X"09",X"5A",X"07",X"2B",X"08",X"07",X"08",X"4B",X"07",X"71",X"09",
		X"DD",X"01",X"28",X"FD",X"FD",X"03",X"27",X"F3",X"33",X"04",X"87",X"07",X"9F",X"08",X"70",X"06",
		X"66",X"FB",X"96",X"04",X"15",X"F8",X"0C",X"F8",X"EB",X"F7",X"51",X"05",X"44",X"FA",X"83",X"08",
		X"BC",X"03",X"29",X"F8",X"2F",X"F6",X"D4",X"00",X"01",X"00",X"04",X"FF",X"33",X"0B",X"A6",X"05",
		X"6C",X"09",X"A8",X"06",X"72",X"08",X"F8",X"07",X"A2",X"03",X"BB",X"FA",X"24",X"0B",X"30",X"F5",
		X"69",X"FD",X"32",X"02",X"54",X"FC",X"9F",X"09",X"07",X"01",X"82",X"F4",X"D2",X"03",X"7B",X"FD",
		X"19",X"F6",X"9D",X"06",X"5C",X"06",X"68",X"FA",X"21",X"06",X"78",X"F4",X"21",X"00",X"3F",X"01",
		X"B5",X"F6",X"9F",X"F7",X"E7",X"FB",X"A2",X"04",X"9C",X"F5",X"04",X"F9",X"46",X"FE",X"67",X"0C",
		X"7F",X"F9",X"40",X"05",X"A0",X"07",X"D7",X"07",X"19",X"F6",X"91",X"FD",X"21",X"02",X"40",X"FD",
		X"A6",X"03",X"39",X"F4",X"15",X"FB",X"84",X"F4",X"D6",X"FF",X"0D",X"01",X"64",X"FD",X"49",X"0B",
		X"D8",X"FC",X"C0",X"F6",X"9C",X"04",X"0F",X"FC",X"D9",X"03",X"47",X"FB",X"18",X"08",X"01",X"07",
		X"90",X"09",X"C9",X"FF",X"09",X"FE",X"98",X"0B",X"E5",X"FA",X"78",X"FB",X"57",X"0B",X"EA",X"FD",
		X"6C",X"00",X"77",X"00",X"62",X"F4",X"74",X"06",X"3C",X"07",X"57",X"08",X"5F",X"07",X"E5",X"05",
		X"B1",X"F4",X"FB",X"FF",X"88",X"01",X"2B",X"F6",X"6E",X"F8",X"BE",X"01",X"4A",X"FF",X"C7",X"F2",
		X"A1",X"03",X"8A",X"FD",X"3F",X"01",X"30",X"09",X"21",X"07",X"15",X"FB",X"9F",X"04",X"42",X"FA",
		X"30",X"09",X"8D",X"05",X"16",X"0B",X"7C",X"FD",X"58",X"01",X"A4",X"FE",X"AB",X"00",X"18",X"0A",
		X"5F",X"06",X"35",X"08",X"F1",X"07",X"5D",X"FE",X"80",X"F5",X"58",X"05",X"16",X"FB",X"5E",X"05",
		X"4B",X"09",X"3B",X"03",X"F6",X"FA",X"FA",X"0A",X"9C",X"FE",X"94",X"FE",X"ED",X"0A",X"3C",X"FB",
		X"AB",X"F7",X"36",X"04",X"C3",X"FB",X"41",X"04",X"C3",X"F7",X"97",X"02",X"8B",X"09",X"77",X"05",
		X"23",X"FB",X"CE",X"06",X"36",X"05",X"EA",X"F5",X"69",X"F9",X"9F",X"F6",X"08",X"F9",X"0C",X"F7",
		X"79",X"F8",X"D1",X"02",X"8D",X"FD",X"E6",X"01",X"67",X"FD",X"2A",X"03",X"01",X"F8",X"B5",X"03",
		X"8B",X"09",X"17",X"05",X"A3",X"F8",X"4A",X"FA",X"8A",X"09",X"8A",X"06",X"0A",X"03",X"D7",X"F2",
		X"67",X"05",X"7A",X"FB",X"B2",X"03",X"10",X"08",X"FC",X"F8",X"AD",X"F7",X"35",X"F8",X"CF",X"F7",
		X"57",X"F8",X"E0",X"04",X"7F",X"F9",X"3A",X"F9",X"A1",X"09",X"69",X"02",X"EB",X"F6",X"FA",X"F8",
		X"98",X"F6",X"0D",X"02",X"E6",X"08",X"13",X"07",X"B6",X"FA",X"FD",X"F7",X"43",X"08",X"86",X"06",
		X"68",X"09",X"15",X"01",X"BF",X"FC",X"18",X"0A",X"19",X"F4",X"99",X"FF",X"0C",X"00",X"95",X"FF",
		X"12",X"00",X"92",X"FF",X"28",X"00",X"42",X"FF",X"AF",X"0B",X"26",X"F7",X"33",X"FB",X"B9",X"03",
		X"11",X"F9",X"C3",X"F6",X"50",X"FD",X"65",X"0A",X"50",X"FE",X"90",X"F9",X"24",X"06",X"AC",X"F4",
		X"98",X"FF",X"FF",X"07",X"BE",X"07",X"56",X"07",X"D7",X"07",X"65",X"07",X"19",X"07",X"36",X"FA",
		X"F7",X"06",X"21",X"08",X"5F",X"03",X"45",X"FA",X"FA",X"0C",X"26",X"FB",X"F0",X"02",X"07",X"04",
		X"0C",X"F8",X"1F",X"F6",X"13",X"01",X"58",X"FF",X"6D",X"FF",X"5D",X"0A",X"B7",X"05",X"BF",X"08",
		X"C4",X"05",X"D3",X"F7",X"9A",X"FB",X"73",X"04",X"EC",X"F5",X"B5",X"F8",X"3C",X"FE",X"66",X"0B",
		X"E6",X"FA",X"C0",X"F7",X"58",X"FC",X"CE",X"0B",X"FD",X"FB",X"91",X"01",X"F2",X"08",X"38",X"FB",
		X"68",X"F6",X"BD",X"FA",X"26",X"04",X"7A",X"F8",X"67",X"F7",X"21",X"F9",X"18",X"F6",X"87",X"01",
		X"E8",X"FF",X"12",X"F5",X"6D",X"05",X"95",X"07",X"B2",X"07",X"51",X"07",X"B0",X"07",X"48",X"07",
		X"BC",X"07",X"99",X"06",X"54",X"FA",X"2B",X"07",X"06",X"07",X"77",X"08",X"03",X"02",X"A0",X"F5",
		X"36",X"00",X"0C",X"0A",X"31",X"FB",X"47",X"03",X"15",X"08",X"35",X"F9",X"B2",X"F6",X"6C",X"02",
		X"2C",X"FE",X"55",X"F5",X"AA",X"FA",X"71",X"03",X"51",X"FB",X"1C",X"08",X"C9",X"02",X"F2",X"FA",
		X"16",X"0C",X"28",X"FC",X"0D",X"01",X"4D",X"09",X"F3",X"FA",X"A1",X"03",X"AB",X"FA",X"E9",X"F7",
		X"0B",X"0A",X"52",X"FA",X"66",X"04",X"4F",X"07",X"DD",X"F8",X"15",X"F9",X"F5",X"09",X"94",X"00",
		X"F8",X"FD",X"94",X"02",X"E9",X"F4",X"33",X"FA",X"36",X"F6",X"DB",X"F9",X"14",X"F6",X"5B",X"FB",
		X"06",X"03",X"15",X"FC",X"62",X"07",X"C2",X"07",X"E8",X"F9",X"27",X"07",X"81",X"04",X"D5",X"FA",
		X"06",X"09",X"F9",X"05",X"6D",X"09",X"E5",X"FD",X"B8",X"FF",X"38",X"0A",X"36",X"05",X"31",X"09",
		X"A2",X"05",X"BA",X"07",X"64",X"F4",X"69",X"FF",X"FA",X"00",X"22",X"F8",X"7B",X"F6",X"4D",X"FC",
		X"AC",X"02",X"D0",X"FB",X"6B",X"09",X"B1",X"00",X"B0",X"F4",X"D0",X"03",X"E5",X"FC",X"11",X"F7",
		X"03",X"05",X"E6",X"08",X"E1",X"03",X"63",X"FB",X"D9",X"07",X"2A",X"07",X"40",X"07",X"57",X"07",
		X"6D",X"07",X"B8",X"04",X"5D",X"F5",X"94",X"FE",X"B9",X"08",X"61",X"FF",X"81",X"F5",X"12",X"FA",
		X"DB",X"F5",X"E9",X"FA",X"45",X"02",X"14",X"FD",X"BA",X"04",X"CC",X"0A",X"76",X"FE",X"05",X"00",
		X"E2",X"FF",X"93",X"F8",X"70",X"08",X"24",X"07",X"A5",X"02",X"9C",X"F4",X"B2",X"01",X"B6",X"07",
		X"8B",X"07",X"60",X"FB",X"D4",X"03",X"D9",X"07",X"70",X"F6",X"F5",X"FB",X"B2",X"07",X"0D",X"03",
		X"14",X"F4",X"90",X"02",X"63",X"FE",X"9F",X"F6",X"90",X"F8",X"FD",X"F7",X"70",X"F7",X"9F",X"FF",
		X"4F",X"0A",X"B5",X"FA",X"9A",X"03",X"66",X"08",X"77",X"06",X"3D",X"08",X"AB",X"03",X"1D",X"FA",
		X"6E",X"0B",X"1E",X"FD",X"D6",X"00",X"D9",X"FE",X"92",X"FF",X"F3",X"0A",X"D6",X"FF",X"C8",X"F6",
		X"AA",X"FF",X"1E",X"0A",X"A7",X"FA",X"70",X"03",X"E9",X"07",X"19",X"F8",X"B3",X"F8",X"04",X"F7",
		X"81",X"F9",X"8F",X"F5",X"EB",X"00",X"69",X"FF",X"C1",X"FE",X"AC",X"0A",X"D6",X"F9",X"60",X"04",
		X"07",X"09",X"F2",X"FD",X"67",X"FF",X"99",X"0A",X"1F",X"F9",X"2F",X"05",X"89",X"F9",X"61",X"08",
		X"52",X"02",X"2E",X"FC",X"DF",X"07",X"F3",X"07",X"B9",X"FE",X"A9",X"FE",X"C1",X"0A",X"57",X"F9",
		X"9F",X"F8",X"40",X"F7",X"C8",X"F8",X"71",X"F7",X"73",X"F8",X"06",X"03",X"93",X"FC",X"03",X"04",
		X"D4",X"07",X"18",X"F4",X"07",X"00",X"09",X"00",X"EB",X"FD",X"19",X"09",X"10",X"06",X"3E",X"08",
		X"29",X"FB",X"9B",X"03",X"BA",X"08",X"E1",X"05",X"43",X"08",X"F2",X"05",X"25",X"08",X"B2",X"F8",
		X"8D",X"F9",X"9A",X"06",X"0C",X"05",X"E4",X"F4",X"A0",X"FF",X"52",X"01",X"FC",X"F4",X"B2",X"02",
		X"FD",X"FD",X"86",X"F5",X"B3",X"06",X"F2",X"04",X"0F",X"FB",X"91",X"06",X"83",X"07",X"8D",X"06",
		X"C8",X"07",X"1A",X"05",X"F7",X"F9",X"B4",X"08",X"29",X"01",X"BB",X"FC",X"73",X"03",X"EE",X"F2",
		X"99",X"04",X"E6",X"FB",X"A1",X"F7",X"E7",X"03",X"60",X"FA",X"E6",X"F7",X"E4",X"09",X"71",X"00",
		X"42",X"FD",X"60",X"07",X"AB",X"F8",X"BA",X"F7",X"7F",X"F8",X"6C",X"F7",X"19",X"F9",X"3E",X"F6",
		X"57",X"01",X"79",X"FF",X"1F",X"F5",X"59",X"05",X"99",X"FA",X"8A",X"05",X"79",X"07",X"0B",X"07",
		X"08",X"07",X"3B",X"07",X"D3",X"06",X"61",X"07",X"92",X"06",X"AC",X"07",X"FE",X"05",X"DB",X"08",
		X"D7",X"FE",X"05",X"FE",X"6B",X"0A",X"6A",X"FA",X"22",X"03",X"D7",X"07",X"C3",X"F7",X"BE",X"FA",
		X"14",X"04",X"5F",X"F6",X"00",X"FD",X"9D",X"09",X"B6",X"FD",X"04",X"FF",X"58",X"0A",X"61",X"00",
		X"4B",X"FC",X"26",X"0A",X"E2",X"FC",X"D0",X"FF",X"93",X"09",X"BE",X"F9",X"2E",X"04",X"16",X"F9",
		X"BF",X"F9",X"11",X"05",X"05",X"F5",X"2D",X"FF",X"80",X"01",X"E3",X"F4",X"65",X"02",X"3F",X"FE",
		X"C4",X"F4",X"B1",X"FF",X"41",X"01",X"C9",X"F4",X"2A",X"03",X"37",X"FD",X"42",X"F6",X"6D",X"F9",
		X"E7",X"F6",X"7D",X"F9",X"42",X"F6",X"A8",X"FD",X"20",X"03",X"AC",X"F4",X"1C",X"02",X"9E",X"FE",
		X"5B",X"FF",X"98",X"0B",X"09",X"FE",X"18",X"FF",X"4E",X"08",X"7B",X"06",X"89",X"07",X"6E",X"FB",
		X"6F",X"03",X"E8",X"08",X"4A",X"05",X"D1",X"08",X"C2",X"04",X"25",X"0A",X"72",X"FD",X"44",X"00",
		X"74",X"FF",X"81",X"F5",X"35",X"04",X"84",X"07",X"E6",X"F7",X"31",X"00",X"38",X"08",X"99",X"06",
		X"BC",X"FB",X"A7",X"02",X"E1",X"FA",X"07",X"F6",X"73",X"FC",X"C8",X"03",X"BF",X"F4",X"0F",X"01",
		X"16",X"FF",X"B3",X"FE",X"15",X"0A",X"9B",X"04",X"1B",X"09",X"F1",X"03",X"77",X"FA",X"98",X"F5",
		X"6D",X"04",X"1B",X"FB",X"B7",X"03",X"99",X"F9",X"E9",X"F7",X"AD",X"F7",X"B8",X"FB",X"9A",X"09",
		X"D1",X"FE",X"FA",X"FD",X"79",X"0A",X"B9",X"FA",X"68",X"F8",X"A3",X"03",X"D6",X"08",X"03",X"05",
		X"4D",X"09",X"74",X"FA",X"DE",X"F8",X"3E",X"03",X"04",X"0A",X"5C",X"01",X"1F",X"FE",X"67",X"00",
		X"50",X"FE",X"A4",X"00",X"3E",X"FD",X"74",X"0A",X"02",X"FB",X"B7",X"F7",X"32",X"04",X"C7",X"F9",
		X"C2",X"F7",X"1B",X"F8",X"84",X"F8",X"A4",X"F7",X"FD",X"05",X"E6",X"04",X"39",X"FB",X"32",X"04",
		X"37",X"F6",X"B4",X"FD",X"59",X"09",X"26",X"FE",X"39",X"F7",X"92",X"F8",X"37",X"F8",X"F4",X"03",
		X"91",X"FA",X"C9",X"F6",X"D9",X"F9",X"10",X"F6",X"D1",X"FE",X"38",X"06",X"50",X"FB",X"D3",X"03",
		X"85",X"F8",X"66",X"F7",X"9C",X"FD",X"65",X"09",X"9E",X"FE",X"AD",X"F6",X"9D",X"F9",X"33",X"F7",
		X"A0",X"05",X"D9",X"F8",X"25",X"F9",X"24",X"F7",X"38",X"FA",X"93",X"F5",X"60",X"01",X"A8",X"FF",
		X"A1",X"F7",X"98",X"F7",X"D7",X"FD",X"03",X"03",X"0A",X"F6",X"1E",X"FA",X"ED",X"F6",X"67",X"03",
		X"46",X"08",X"DA",X"F9",X"76",X"F8",X"8E",X"F9",X"BC",X"09",X"98",X"00",X"B4",X"FE",X"83",X"01",
		X"4C",X"FD",X"F8",X"0A",X"32",X"04",X"79",X"0A",X"0E",X"FF",X"8F",X"FE",X"C2",X"09",X"17",X"FD",
		X"7A",X"F7",X"28",X"F9",X"A1",X"04",X"3B",X"08",X"92",X"06",X"8E",X"05",X"43",X"F5",X"18",X"00",
		X"79",X"01",X"ED",X"F5",X"05",X"02",X"7E",X"08",X"23",X"06",X"12",X"08",X"15",X"06",X"3C",X"08",
		X"B2",X"05",X"D2",X"08",X"E9",X"F9",X"54",X"F9",X"82",X"F6",X"F1",X"FC",X"E4",X"01",X"A5",X"FD",
		X"7E",X"02",X"48",X"F7",X"CC",X"F7",X"2A",X"02",X"0B",X"FE",X"AD",X"01",X"1A",X"09",X"AE",X"06",
		X"96",X"FF",X"9E",X"FE",X"0D",X"0B",X"DB",X"03",X"A0",X"09",X"D9",X"F5",X"F4",X"FD",X"FD",X"00",
		X"39",X"FE",X"1D",X"02",X"1F",X"F7",X"D9",X"F8",X"9A",X"F8",X"E4",X"F7",X"EE",X"03",X"B8",X"07",
		X"A4",X"F8",X"DF",X"FF",X"FC",X"09",X"F6",X"FA",X"A5",X"F8",X"7C",X"F8",X"49",X"06",X"91",X"F6",
		X"30",X"FE",X"7C",X"01",X"CE",X"FD",X"E7",X"02",X"E1",X"F4",X"F9",X"02",X"07",X"08",X"B5",X"FB",
		X"FB",X"F7",X"E5",X"05",X"AF",X"F7",X"9E",X"02",X"44",X"FE",X"0B",X"F6",X"A0",X"FA",X"73",X"F7",
		X"5D",X"0A",X"55",X"00",X"85",X"FF",X"3F",X"00",X"70",X"FF",X"85",X"00",X"A0",X"FE",X"E5",X"0A",
		X"9B",X"F9",X"65",X"F9",X"6D",X"F7",X"94",X"FB",X"7B",X"04",X"70",X"F7",X"99",X"F9",X"60",X"F8",
		X"88",X"06",X"AA",X"F6",X"33",X"FE",X"64",X"02",X"95",X"F8",X"3E",X"F7",X"D4",X"01",X"78",X"FF",
		X"B1",X"F6",X"E5",X"F9",X"63",X"F8",X"F9",X"06",X"73",X"05",X"27",X"F8",X"88",X"F9",X"CD",X"F7",
		X"BF",X"FA",X"B4",X"03",X"7B",X"FC",X"80",X"04",X"CC",X"F6",X"CD",X"FE",X"92",X"08",X"F6",X"06",
		X"AB",X"FF",X"75",X"F5",X"96",X"06",X"8E",X"F9",X"1D",X"FA",X"83",X"F6",X"61",X"FE",X"DA",X"01",
		X"AA",X"FD",X"BF",X"07",X"8E",X"FA",X"73",X"07",X"0B",X"05",X"8D",X"F5",X"55",X"01",X"99",X"FF",
		X"47",X"00",X"18",X"00",X"DA",X"FF",X"CF",X"0A",X"CB",X"F8",X"01",X"07",X"F6",X"F6",X"81",X"FD",
		X"82",X"06",X"86",X"08",X"B8",X"05",X"29",X"09",X"CC",X"04",X"B8",X"0A",X"27",X"FF",X"91",X"00",
		X"7B",X"FF",X"8C",X"00",X"68",X"FF",X"96",X"00",X"CE",X"09",X"BF",X"05",X"15",X"07",X"37",X"F8",
		X"3B",X"F9",X"C2",X"F8",X"00",X"F8",X"0F",X"FF",X"B4",X"08",X"F4",X"06",X"23",X"04",X"B0",X"FA",
		X"70",X"0B",X"8C",X"FD",X"38",X"00",X"55",X"09",X"2A",X"FC",X"0B",X"F8",X"87",X"05",X"C7",X"07",
		X"44",X"05",X"6E",X"F7",X"98",X"FD",X"09",X"04",X"A9",X"F4",X"23",X"03",X"BD",X"FE",X"03",X"F7",
		X"AF",X"04",X"9A",X"03",X"50",X"F4",X"4E",X"04",X"D2",X"FC",X"AD",X"02",X"03",X"08",X"DD",X"06",
		X"77",X"F8",X"66",X"FC",X"C4",X"02",X"49",X"FD",X"F0",X"02",X"FB",X"FB",X"BF",X"0B",X"C3",X"FB",
		X"79",X"F9",X"A8",X"F7",X"8B",X"06",X"CB",X"00",X"5C",X"F6",X"B3",X"02",X"6D",X"08",X"41",X"FB",
		X"3A",X"F8",X"09",X"F9",X"21",X"FA",X"3A",X"09",X"76",X"01",X"13",X"FD",X"7C",X"09",X"5F",X"05",
		X"26",X"09",X"06",X"FC",X"BD",X"F8",X"1D",X"04",X"CA",X"09",X"E9",X"FC",X"0D",X"02",X"21",X"FE",
		X"0D",X"02",X"07",X"09",X"9A",X"F7",X"D3",X"FB",X"7F",X"07",X"14",X"03",X"17",X"FB",X"22",X"0C",
		X"8B",X"FB",X"F6",X"02",X"AD",X"FD",X"8D",X"F7",X"62",X"F9",X"89",X"F8",X"1A",X"F9",X"5D",X"F8",
		X"D9",X"02",X"DC",X"08",X"DA",X"F8",X"73",X"FB",X"A0",X"03",X"DF",X"FB",X"3D",X"08",X"7B",X"06",
		X"8B",X"07",X"C1",X"06",X"59",X"07",X"CC",X"06",X"53",X"07",X"AB",X"06",X"9F",X"07",X"E5",X"04",
		X"95",X"F8",X"C7",X"F8",X"EC",X"03",X"DC",X"07",X"F4",X"F7",X"2C",X"FC",X"13",X"04",X"28",X"F7",
		X"FA",X"FD",X"D5",X"09",X"97",X"FD",X"71",X"00",X"7E",X"09",X"87",X"FA",X"36",X"F9",X"C8",X"05",
		X"79",X"07",X"9B",X"06",X"53",X"07",X"86",X"06",X"95",X"07",X"FD",X"04",X"C3",X"FA",X"75",X"08",
		X"22",X"02",X"AE",X"F7",X"43",X"F9",X"5F",X"F8",X"06",X"F9",X"90",X"F8",X"04",X"F9",X"B1",X"04",
		X"F5",X"07",X"12",X"06",X"1A",X"08",X"F0",X"02",X"CB",X"F6",X"6D",X"FF",X"56",X"07",X"36",X"F7",
		X"A9",X"FA",X"1D",X"F6",X"77",X"00",X"D5",X"00",X"51",X"F7",X"59",X"F9",X"C8",X"F8",X"9E",X"F8",
		X"99",X"05",X"A8",X"06",X"5B",X"08",X"63",X"02",X"6D",X"FD",X"AE",X"02",X"1E",X"FC",X"16",X"0B",
		X"BA",X"01",X"03",X"FD",X"69",X"07",X"73",X"06",X"1E",X"08",X"7E",X"FE",X"9E",X"FF",X"2A",X"0A",
		X"81",X"F9",X"52",X"FA",X"A3",X"03",X"A7",X"FB",X"65",X"07",X"5F",X"03",X"6B",X"F6",X"82",X"FF",
		X"01",X"09",X"58",X"FD",X"AA",X"00",X"46",X"0A",X"3A",X"FF",X"2F",X"FE",X"15",X"0A",X"CD",X"FB",
		X"A2",X"02",X"14",X"FD",X"4E",X"F7",X"9A",X"07",X"12",X"04",X"E0",X"F8",X"A5",X"F8",X"D9",X"F8",
		X"E2",X"F8",X"3D",X"F8",X"CB",X"00",X"95",X"09",X"D7",X"F9",X"3C",X"FE",X"49",X"08",X"98",X"06",
		X"0C",X"FF",X"E9",X"F5",X"FF",X"05",X"9E",X"F9",X"C6",X"F9",X"EE",X"F6",X"D7",X"FD",X"8E",X"02",
		X"85",X"F8",X"AD",X"F7",X"56",X"01",X"DB",X"FF",X"58",X"F6",X"BB",X"04",X"0A",X"08",X"64",X"00",
		X"FD",X"F6",X"3B",X"FA",X"AA",X"F7",X"C0",X"04",X"2F",X"FB",X"E7",X"F7",X"3B",X"FB",X"E2",X"07",
		X"2B",X"03",X"97",X"F6",X"18",X"00",X"0C",X"08",X"77",X"06",X"43",X"07",X"BB",X"06",X"0D",X"07",
		X"E0",X"06",X"C5",X"06",X"70",X"07",X"C3",X"FC",X"3F",X"02",X"A3",X"09",X"0E",X"03",X"12",X"FD",
		X"35",X"05",X"82",X"09",X"F1",X"FE",X"E5",X"FF",X"8B",X"00",X"FB",X"F6",X"50",X"F9",X"47",X"03",
		X"6E",X"FC",X"D2",X"04",X"01",X"06",X"E1",X"F7",X"60",X"F9",X"3F",X"03",X"AC",X"FC",X"5A",X"04",
		X"A6",X"08",X"E6",X"02",X"73",X"F8",X"9D",X"F8",X"13",X"FE",X"97",X"0A",X"43",X"FB",X"71",X"03",
		X"49",X"FC",X"4E",X"F8",X"6E",X"F8",X"4E",X"FB",X"59",X"06",X"EC",X"07",X"79",X"FA",X"27",X"06",
		X"33",X"04",X"08",X"FD",X"26",X"02",X"BA",X"FD",X"14",X"02",X"E6",X"FC",X"EF",X"09",X"AF",X"04",
		X"A3",X"08",X"CB",X"FA",X"AA",X"04",X"97",X"06",X"2E",X"F8",X"EA",X"F9",X"87",X"F7",X"93",X"FA",
		X"8E",X"F6",X"23",X"FD",X"60",X"01",X"D8",X"FE",X"9E",X"00",X"55",X"FF",X"47",X"00",X"7C",X"FF",
		X"87",X"00",X"2D",X"F6",X"8D",X"FA",X"13",X"04",X"F9",X"06",X"7C",X"F8",X"EA",X"F8",X"41",X"FC",
		X"95",X"08",X"F7",X"05",X"27",X"06",X"C5",X"F9",X"A4",X"09",X"5F",X"00",X"C6",X"FD",X"9E",X"08",
		X"84",X"05",X"44",X"08",X"33",X"FC",X"42",X"F8",X"77",X"F9",X"4F",X"06",X"B1",X"04",X"A5",X"FA",
		X"83",X"09",X"F2",X"FF",X"D3",X"FD",X"9B",X"09",X"8B",X"02",X"34",X"FC",X"37",X"08",X"8B",X"01",
		X"44",X"F6",X"9D",X"01",X"66",X"07",X"B9",X"06",X"37",X"FC",X"B0",X"02",X"FC",X"FC",X"C1",X"02",
		X"11",X"FC",X"55",X"07",X"EB",X"06",X"61",X"01",X"2E",X"F6",X"41",X"FB",X"E6",X"F5",X"FF",X"FF",
		X"6D",X"00",X"26",X"FE",X"E3",X"08",X"81",X"05",X"74",X"07",X"4B",X"06",X"35",X"06",X"DF",X"FA",
		X"CD",X"04",X"A0",X"F7",X"49",X"FA",X"C4",X"F6",X"8A",X"00",X"D6",X"00",X"CE",X"F5",X"38",X"04",
		X"8D",X"FC",X"2C",X"F7",X"7B",X"FF",X"46",X"09",X"5D",X"FC",X"03",X"02",X"70",X"08",X"10",X"05",
		X"5D",X"FA",X"A4",X"F9",X"A3",X"08",X"7C",X"04",X"C0",X"09",X"92",X"FD",X"0D",X"01",X"D1",X"FE",
		X"4C",X"00",X"47",X"09",X"7B",X"04",X"55",X"FB",X"66",X"F7",X"17",X"FA",X"D0",X"F7",X"F8",X"F9",
		X"C5",X"F7",X"0E",X"FB",X"F0",X"05",X"22",X"07",X"AF",X"06",X"D7",X"02",X"42",X"F5",X"D3",X"02",
		X"87",X"FE",X"4C",X"F7",X"FF",X"03",X"88",X"FC",X"10",X"03",X"E3",X"FA",X"1B",X"F7",X"32",X"04",
		X"3A",X"FC",X"DE",X"03",X"63",X"08",X"55",X"03",X"CA",X"FB",X"D1",X"07",X"51",X"06",X"F8",X"01",
		X"EF",X"F4",X"75",X"04",X"31",X"FC",X"42",X"03",X"F1",X"06",X"A8",X"FA",X"46",X"06",X"AC",X"06",
		X"A5",X"06",X"43",X"FC",X"73",X"02",X"3D",X"FD",X"46",X"02",X"CF",X"FC",X"BE",X"03",X"0F",X"F6",
		X"55",X"00",X"63",X"07",X"55",X"06",X"B1",X"06",X"A8",X"06",X"F6",X"05",X"39",X"FA",X"C2",X"F7",
		X"74",X"FC",X"CF",X"03",X"AA",X"F6",X"57",X"FB",X"32",X"03",X"3D",X"FA",X"DB",X"F7",X"34",X"FA",
		X"27",X"F7",X"12",X"00",X"8C",X"07",X"5B",X"06",X"AA",X"06",X"BA",X"06",X"4E",X"06",X"39",X"07",
		X"30",X"04",X"CA",X"FA",X"E9",X"08",X"6A",X"00",X"4C",X"F9",X"37",X"04",X"E7",X"FA",X"CF",X"07",
		X"6C",X"02",X"8B",X"F6",X"96",X"00",X"98",X"00",X"E1",X"F5",X"1E",X"04",X"66",X"06",X"C0",X"FB",
		X"76",X"03",X"FD",X"F9",X"5A",X"F8",X"64",X"F9",X"A0",X"F8",X"20",X"F9",X"DF",X"F9",X"7F",X"07",
		X"51",X"03",X"64",X"F7",X"7F",X"FE",X"1B",X"08",X"9E",X"05",X"6D",X"07",X"C7",X"05",X"3A",X"07",
		X"73",X"FA",X"EE",X"05",X"EE",X"05",X"07",X"08",X"3D",X"01",X"53",X"FD",X"38",X"03",X"87",X"F4",
		X"0F",X"04",X"03",X"03",X"0F",X"F8",X"39",X"FD",X"0E",X"0A",X"55",X"FC",X"8D",X"01",X"50",X"07",
		X"4B",X"06",X"FF",X"FA",X"96",X"04",X"14",X"F8",X"B7",X"FC",X"EC",X"05",X"5A",X"08",X"AA",X"FE",
		X"59",X"FF",X"AF",X"07",X"D2",X"06",X"CB",X"01",X"2B",X"FC",X"AB",X"09",X"B4",X"FD",X"92",X"F7",
		X"DD",X"02",X"20",X"07",X"6F",X"FA",X"14",X"F8",X"01",X"FA",X"FC",X"F6",X"BE",X"FE",X"15",X"01",
		X"4A",X"FD",X"D9",X"08",X"1A",X"05",X"42",X"07",X"0A",X"06",X"B7",X"FA",X"AB",X"FD",X"C9",X"09",
		X"F0",X"FB",X"F0",X"F8",X"9B",X"F8",X"27",X"05",X"85",X"05",X"8B",X"F8",X"6B",X"FB",X"74",X"08",
		X"27",X"00",X"3B",X"FD",X"BE",X"09",X"60",X"FC",X"D6",X"F8",X"9C",X"F8",X"65",X"F9",X"71",X"F8",
		X"87",X"F9",X"75",X"F8",X"72",X"F9",X"F2",X"02",X"FA",X"07",X"71",X"F7",X"38",X"FD",X"0E",X"02",
		X"93",X"FC",X"E8",X"07",X"84",X"05",X"DA",X"07",X"66",X"FD",X"AD",X"00",X"05",X"09",X"72",X"04",
		X"AC",X"07",X"43",X"F6",X"1D",X"04",X"FE",X"FB",X"2F",X"F9",X"4C",X"03",X"8D",X"FB",X"69",X"F6",
		X"7F",X"FE",X"42",X"01",X"0F",X"FD",X"C3",X"08",X"F0",X"FE",X"B9",X"F6",X"DE",X"03",X"3D",X"FC",
		X"10",X"F8",X"42",X"FA",X"9C",X"06",X"DD",X"03",X"F7",X"F7",X"08",X"04",X"E6",X"FB",X"BC",X"04",
		X"78",X"07",X"6B",X"05",X"12",X"08",X"4F",X"00",X"2C",X"FD",X"30",X"0A",X"56",X"FB",X"D4",X"02",
		X"C9",X"FC",X"85",X"02",X"47",X"FC",X"23",X"05",X"F3",X"06",X"1D",X"06",X"8D",X"06",X"D5",X"05",
		X"3B",X"F9",X"91",X"F9",X"A6",X"F7",X"C1",X"FD",X"88",X"06",X"90",X"07",X"15",X"FE",X"D0",X"FF",
		X"C3",X"08",X"AF",X"FA",X"11",X"04",X"9A",X"06",X"37",X"F7",X"C6",X"FD",X"75",X"01",X"FD",X"FC",
		X"2F",X"07",X"D4",X"F8",X"89",X"FA",X"78",X"08",X"1E",X"00",X"7C",X"FE",X"79",X"01",X"D6",X"F6",
		X"1A",X"FA",X"79",X"F8",X"49",X"F9",X"31",X"04",X"B3",X"F9",X"4D",X"FB",X"E3",X"03",X"10",X"F8",
		X"68",X"F9",X"47",X"F9",X"2A",X"F8",X"84",X"FC",X"BF",X"02",X"75",X"FC",X"27",X"04",X"94",X"F4",
		X"C7",X"03",X"2F",X"FD",X"A2",X"01",X"18",X"08",X"2E",X"FA",X"1D",X"06",X"CA",X"05",X"D3",X"07",
		X"99",X"01",X"5D",X"FC",X"B8",X"09",X"45",X"FD",X"65",X"00",X"42",X"08",X"21",X"05",X"7E",X"07",
		X"35",X"05",X"EB",X"07",X"43",X"FD",X"E8",X"F7",X"BF",X"03",X"68",X"FB",X"F3",X"F8",X"39",X"07",
		X"36",X"05",X"96",X"07",X"DF",X"04",X"62",X"08",X"1C",X"FE",X"97",X"F8",X"BE",X"F8",X"D0",X"F9",
		X"73",X"F7",X"71",X"00",X"75",X"00",X"10",X"F6",X"56",X"04",X"F4",X"FB",X"98",X"03",X"F5",X"07",
		X"1F",X"03",X"FE",X"FB",X"72",X"04",X"16",X"F5",X"36",X"02",X"1B",X"FE",X"B0",X"00",X"03",X"FF",
		X"A0",X"F6",X"F7",X"FA",X"29",X"F7",X"20",X"01",X"F3",X"07",X"0C",X"FC",X"DC",X"02",X"1B",X"07",
		X"DD",X"F9",X"3A",X"07",X"23",X"05",X"BC",X"07",X"A0",X"04",X"D3",X"08",X"14",X"FD",X"D1",X"00",
		X"5E",X"07",X"21",X"06",X"CC",X"05",X"BE",X"07",X"7B",X"FD",X"B1",X"00",X"B6",X"FE",X"84",X"F6",
		X"8C",X"06",X"E1",X"03",X"6E",X"FB",X"F9",X"06",X"4F",X"02",X"AD",X"F7",X"C9",X"F9",X"AB",X"F8",
		X"E9",X"F8",X"BF",X"01",X"FE",X"07",X"8B",X"04",X"D4",X"FB",X"09",X"05",X"BA",X"06",X"24",X"06",
		X"D9",X"FB",X"AA",X"03",X"19",X"06",X"48",X"F8",X"5E",X"F9",X"BB",X"FB",X"FD",X"08",X"24",X"FF",
		X"8B",X"F7",X"AD",X"01",X"A1",X"FE",X"65",X"F6",X"CF",X"FB",X"E6",X"01",X"33",X"FD",X"B5",X"02",
		X"A1",X"F8",X"6B",X"03",X"6B",X"FB",X"35",X"F9",X"BF",X"05",X"08",X"F6",X"C5",X"FF",X"72",X"00",
		X"78",X"FD",X"8B",X"09",X"EC",X"FB",X"26",X"02",X"53",X"FD",X"9B",X"F7",X"D9",X"06",X"F6",X"04",
		X"1C",X"08",X"72",X"01",X"42",X"F9",X"53",X"03",X"17",X"FC",X"05",X"05",X"5F",X"07",X"C3",X"04",
		X"9E",X"08",X"D7",X"FD",X"6A",X"00",X"05",X"FF",X"AB",X"FF",X"67",X"09",X"F8",X"02",X"9B",X"FD",
		X"37",X"01",X"8A",X"FD",X"35",X"02",X"57",X"F8",X"F5",X"F8",X"D8",X"FA",X"A5",X"03",X"B8",X"FA",
		X"E5",X"08",X"BE",X"FF",X"C1",X"F8",X"ED",X"F8",X"97",X"F9",X"6B",X"F8",X"A3",X"03",X"0B",X"FC",
		X"55",X"03",X"0B",X"FB",X"C5",X"07",X"10",X"01",X"1C",X"FD",X"B7",X"07",X"D9",X"05",X"47",X"04",
		X"87",X"FA",X"AF",X"08",X"D1",X"03",X"35",X"09",X"3A",X"FC",X"E7",X"01",X"64",X"FD",X"A0",X"01",
		X"B7",X"FC",X"FC",X"F6",X"35",X"FC",X"99",X"05",X"99",X"06",X"E6",X"05",X"3A",X"06",X"A3",X"06",
		X"82",X"FE",X"31",X"F7",X"99",X"FA",X"67",X"F7",X"89",X"FF",X"15",X"08",X"C2",X"FC",X"47",X"01",
		X"08",X"FE",X"76",X"01",X"86",X"09",X"2E",X"01",X"DA",X"FD",X"F8",X"01",X"3F",X"F8",X"A4",X"F9",
		X"3A",X"F8",X"40",X"01",X"2A",X"FF",X"BE",X"F5",X"18",X"00",X"0F",X"06",X"9C",X"06",X"F8",X"05",
		X"97",X"FD",X"0B",X"F7",X"DD",X"FA",X"52",X"F8",X"74",X"08",X"37",X"01",X"90",X"FA",X"AB",X"F6",
		X"4B",X"01",X"39",X"FF",X"5D",X"F8",X"F6",X"F8",X"7C",X"03",X"45",X"FB",X"CA",X"FD",X"B0",X"09",
		X"6A",X"FB",X"CF",X"02",X"CA",X"FC",X"99",X"02",X"06",X"FC",X"02",X"06",X"31",X"03",X"64",X"FB",
		X"AE",X"08",X"34",X"04",X"5C",X"08",X"10",X"FD",X"65",X"F8",X"2A",X"03",X"1F",X"FC",X"F7",X"F7",
		X"C1",X"F9",X"48",X"00",X"E8",X"08",X"94",X"03",X"F9",X"FD",X"BF",X"00",X"A4",X"FE",X"94",X"00",
		X"7F",X"FE",X"1D",X"01",X"1F",X"FD",X"64",X"09",X"8F",X"FC",X"F8",X"F8",X"40",X"F9",X"46",X"04",
		X"C0",X"06",X"E2",X"05",X"56",X"06",X"22",X"06",X"C2",X"05",X"CC",X"FB",X"D0",X"02",X"3B",X"FC",
		X"70",X"03",X"02",X"F8",X"8A",X"F9",X"CD",X"FD",X"4F",X"09",X"62",X"FC",X"F7",X"F8",X"AB",X"02",
		X"8E",X"FC",X"06",X"F8",X"3D",X"08",X"A8",X"01",X"3A",X"FA",X"FE",X"F7",X"65",X"06",X"7A",X"03",
		X"21",X"FB",X"99",X"F6",X"F4",X"FF",X"B8",X"FF",X"40",X"FF",X"B3",X"00",X"05",X"F7",X"A6",X"FA",
		X"87",X"F8",X"D5",X"04",X"C3",X"06",X"4B",X"04",X"DD",X"F8",X"B0",X"F9",X"FA",X"F8",X"4D",X"FA",
		X"77",X"04",X"88",X"F8",X"28",X"FD",X"59",X"03",X"16",X"F7",X"5A",X"FB",X"FA",X"F6",X"8B",X"03",
		X"E9",X"FC",X"B9",X"02",X"5E",X"07",X"07",X"06",X"89",X"04",X"AF",X"FA",X"07",X"09",X"93",X"FF",
		X"4F",X"FE",X"58",X"07",X"A1",X"F6",X"35",X"FF",X"81",X"00",X"DA",X"FE",X"EA",X"00",X"02",X"FE",
		X"3A",X"09",X"46",X"04",X"12",X"FE",X"FF",X"00",X"71",X"FE",X"56",X"01",X"4E",X"FD",X"09",X"06",
		X"7F",X"06",X"38",X"06",X"94",X"00",X"E8",X"F5",X"4E",X"FF",X"B2",X"00",X"C2",X"FD",X"86",X"07",
		X"07",X"06",X"A3",X"FE",X"58",X"F7",X"13",X"FB",X"79",X"02",X"FC",X"FB",X"AB",X"F8",X"F9",X"09",
		X"9F",X"FE",X"87",X"00",X"05",X"FF",X"54",X"00",X"63",X"FF",X"1E",X"F8",X"00",X"F9",X"02",X"FF",
		X"A8",X"01",X"09",X"F7",X"E1",X"FA",X"80",X"F8",X"20",X"FA",X"01",X"F9",X"87",X"FA",X"29",X"07",
		X"4E",X"02",X"14",X"FD",X"BA",X"03",X"B0",X"F5",X"EA",X"02",X"61",X"FE",X"44",X"00",X"0C",X"0A",
		X"04",X"FE",X"C0",X"00",X"80",X"FF",X"96",X"FF",X"27",X"09",X"30",X"FA",X"96",X"05",X"8D",X"04",
		X"8E",X"FB",X"DC",X"06",X"A4",X"05",X"CE",X"06",X"7A",X"05",X"52",X"07",X"12",X"FE",X"D6",X"F7",
		X"2B",X"04",X"07",X"FB",X"68",X"FE",X"AE",X"08",X"3E",X"04",X"F9",X"07",X"0E",X"04",X"9E",X"FD",
		X"8E",X"01",X"3C",X"FC",X"17",X"F6",X"8E",X"00",X"5B",X"FF",X"C4",X"FF",X"65",X"00",X"9D",X"F7",
		X"63",X"FA",X"EB",X"F8",X"32",X"FA",X"20",X"05",X"7A",X"06",X"06",X"06",X"5F",X"06",X"E5",X"FB",
		X"0A",X"F9",X"55",X"06",X"61",X"05",X"58",X"07",X"12",X"02",X"BE",X"F7",X"94",X"FF",X"65",X"07",
		X"B0",X"05",X"10",X"FE",X"4C",X"F7",X"46",X"FB",X"97",X"F7",X"9B",X"FC",X"79",X"05",X"2F",X"FE",
		X"E2",X"F6",X"92",X"07",X"33",X"02",X"7C",X"FE",X"C5",X"00",X"DB",X"FE",X"C3",X"00",X"83",X"FE",
		X"D7",X"01",X"BC",X"F5",X"E5",X"04",X"C6",X"FB",X"8D",X"03",X"AE",X"FB",X"30",X"06",X"8B",X"03",
		X"A1",X"F8",X"2A",X"FA",X"87",X"04",X"C2",X"05",X"65",X"F8",X"CA",X"FC",X"6F",X"07",X"34",X"01",
		X"E1",X"F7",X"CF",X"FA",X"17",X"F8",X"58",X"03",X"7A",X"06",X"AC",X"FB",X"A8",X"04",X"FB",X"06",
		X"4E",X"05",X"6F",X"07",X"1D",X"01",X"E2",X"F8",X"9B",X"06",X"9B",X"03",X"4F",X"F9",X"32",X"F9",
		X"A2",X"FD",X"16",X"09",X"25",X"FD",X"ED",X"00",X"AD",X"07",X"EC",X"04",X"A5",X"FC",X"D6",X"02",
		X"D5",X"FA",X"76",X"F8",X"C3",X"FA",X"B3",X"F7",X"52",X"00",X"4F",X"05",X"9E",X"F9",X"C7",X"F8",
		X"15",X"FE",X"F7",X"02",X"54",X"F6",X"18",X"02",X"D5",X"06",X"68",X"FD",X"16",X"F8",X"D3",X"05",
		X"9B",X"05",X"B6",X"05",X"C1",X"F6",X"06",X"00",X"2D",X"00",X"1C",X"FF",X"65",X"01",X"DA",X"F6",
		X"AF",X"FB",X"65",X"F7",X"D2",X"FF",X"8B",X"06",X"BE",X"06",X"39",X"FE",X"18",X"F8",X"D2",X"FA",
		X"78",X"F8",X"13",X"FB",X"A7",X"F7",X"97",X"FE",X"86",X"01",X"02",X"FE",X"EE",X"02",X"F5",X"F5",
		X"D2",X"03",X"CC",X"FD",X"DF",X"F7",X"57",X"FF",X"34",X"07",X"3C",X"06",X"CC",X"FE",X"A4",X"F7",
		X"16",X"05",X"2D",X"06",X"66",X"05",X"7C",X"FA",X"E3",X"08",X"0E",X"00",X"0A",X"FF",X"0A",X"02",
		X"B5",X"F6",X"1E",X"03",X"6E",X"FE",X"2C",X"F7",X"1F",X"00",X"4F",X"06",X"48",X"07",X"2A",X"FD",
		X"1E",X"02",X"A7",X"FD",X"5E",X"F8",X"3F",X"07",X"7C",X"03",X"69",X"F9",X"DC",X"FC",X"58",X"08",
		X"41",X"04",X"AE",X"08",X"44",X"FC",X"CA",X"02",X"33",X"FD",X"89",X"F8",X"5C",X"FA",X"5A",X"F9",
		X"FC",X"F9",X"A0",X"F9",X"FA",X"F9",X"E8",X"04",X"BD",X"05",X"B3",X"F8",X"71",X"FD",X"D4",X"03",
		X"A8",X"F6",X"C3",X"01",X"ED",X"FF",X"41",X"F8",X"B2",X"FA",X"54",X"F9",X"92",X"04",X"E1",X"FA",
		X"97",X"F9",X"FA",X"F9",X"CF",X"F9",X"23",X"FA",X"76",X"04",X"5A",X"FA",X"10",X"FC",X"45",X"04",
		X"E0",X"FA",X"04",X"0B",X"90",X"FC",X"B9",X"02",X"D3",X"FD",X"62",X"02",X"7C",X"FD",X"60",X"F9",
		X"E1",X"04",X"58",X"FB",X"AF",X"07",X"5E",X"FC",X"6B",X"03",X"08",X"07",X"40",X"F9",X"1C",X"FB",
		X"72",X"F8",X"DC",X"FB",X"16",X"F7",X"9C",X"02",X"6A",X"FE",X"AC",X"01",X"C8",X"FE",X"64",X"F8",
		X"B6",X"FA",X"CD",X"F9",X"9A",X"F9",X"B2",X"FC",X"30",X"07",X"DF",X"05",X"75",X"FB",X"7F",X"F9",
		X"9F",X"FB",X"70",X"08",X"BB",X"00",X"DF",X"FE",X"B7",X"02",X"64",X"F6",X"64",X"04",X"31",X"FD",
		X"ED",X"02",X"EF",X"FC",X"59",X"F9",X"45",X"08",X"50",X"02",X"9B",X"FA",X"ED",X"F8",X"4D",X"FC",
		X"CC",X"02",X"F3",X"FD",X"C2",X"02",X"DA",X"FC",X"E6",X"08",X"BA",X"FF",X"EF",X"F8",X"F6",X"FA",
		X"12",X"F9",X"A0",X"04",X"09",X"FC",X"18",X"06",X"02",X"04",X"C1",X"FC",X"93",X"04",X"F4",X"F6",
		X"42",X"01",X"9E",X"06",X"AD",X"06",X"FD",X"05",X"ED",X"06",X"B5",X"05",X"31",X"07",X"3F",X"05",
		X"FC",X"07",X"FE",X"FB",X"FD",X"03",X"78",X"FB",X"2A",X"FB",X"9A",X"05",X"DC",X"07",X"FA",X"00",
		X"EB",X"FE",X"08",X"02",X"3A",X"F8",X"3E",X"FA",X"3F",X"FD",X"4E",X"03",X"58",X"FC",X"B2",X"09",
		X"D2",X"03",X"6A",X"08",X"5B",X"04",X"2D",X"08",X"E2",X"03",X"86",X"FC",X"82",X"F7",X"E3",X"FE",
		X"4F",X"02",X"42",X"F9",X"40",X"FA",X"E3",X"F9",X"41",X"FA",X"65",X"F9",X"E5",X"FD",X"D2",X"07",
		X"5F",X"05",X"F6",X"06",X"08",X"06",X"15",X"FE",X"45",X"F8",X"71",X"06",X"1E",X"05",X"04",X"08",
		X"ED",X"01",X"69",X"FD",X"99",X"07",X"46",X"05",X"7C",X"07",X"24",X"FE",X"03",X"F9",X"64",X"FA",
		X"FB",X"F9",X"4B",X"F9",X"4D",X"01",X"44",X"00",X"FC",X"F6",X"5B",X"06",X"19",X"04",X"99",X"FD",
		X"D0",X"02",X"ED",X"FA",X"59",X"F8",X"1E",X"00",X"9C",X"01",X"F8",X"F7",X"8E",X"FB",X"97",X"F8",
		X"C1",X"04",X"D6",X"FB",X"1F",X"06",X"54",X"FF",X"E5",X"F8",X"82",X"FA",X"B8",X"03",X"48",X"07",
		X"FA",X"04",X"35",X"F9",X"1F",X"FE",X"6E",X"02",X"9B",X"FD",X"B3",X"03",X"C9",X"F5",X"7E",X"04",
		X"55",X"05",X"9C",X"07",X"5A",X"04",X"31",X"FD",X"A6",X"04",X"D3",X"07",X"3E",X"FC",X"17",X"FA",
		X"CF",X"04",X"C7",X"06",X"20",X"06",X"2B",X"04",X"D3",X"F7",X"89",X"FF",X"BF",X"07",X"E8",X"FE",
		X"D2",X"FF",X"5B",X"09",X"3D",X"FA",X"2C",X"06",X"BF",X"03",X"6E",X"FD",X"1F",X"03",X"C5",X"F9",
		X"B8",X"F9",X"58",X"FB",X"DB",X"03",X"C9",X"FA",X"E4",X"F8",X"B6",X"FE",X"02",X"03",X"06",X"F7",
		X"5A",X"02",X"71",X"06",X"71",X"06",X"C7",X"05",X"ED",X"06",X"4D",X"04",X"4E",X"FC",X"6A",X"06",
		X"0C",X"06",X"00",X"06",X"2E",X"FB",X"92",X"FA",X"64",X"07",X"86",X"02",X"B4",X"F9",X"E6",X"F9",
		X"7F",X"FA",X"0D",X"F9",X"26",X"02",X"28",X"07",X"B3",X"05",X"0A",X"06",X"4F",X"FA",X"7D",X"FA",
		X"F5",X"F8",X"86",X"FE",X"8A",X"02",X"7C",X"FC",X"B0",X"0A",X"17",X"00",X"11",X"00",X"67",X"00",
		X"24",X"FF",X"69",X"06",X"63",X"07",X"F9",X"FC",X"C7",X"02",X"31",X"FD",X"18",X"04",X"53",X"05",
		X"B9",X"FB",X"7B",X"06",X"A8",X"06",X"35",X"01",X"8A",X"FD",X"4D",X"09",X"B6",X"01",X"53",X"FD",
		X"48",X"07",X"3A",X"01",X"5A",X"F8",X"42",X"FB",X"A0",X"F8",X"85",X"03",X"A6",X"06",X"22",X"05",
		X"FD",X"FB",X"8A",X"04",X"64",X"F8",X"56",X"FE",X"00",X"07",X"46",X"01",X"DA",X"F6",X"17",X"04",
		X"03",X"02",X"FD",X"FD",X"EB",X"02",X"20",X"F7",X"E5",X"01",X"4D",X"07",X"A5",X"FC",X"F1",X"02",
		X"5B",X"FC",X"25",X"FA",X"98",X"05",X"6A",X"F7",X"E3",X"FF",X"32",X"01",X"A6",X"FD",X"87",X"09",
		X"5D",X"FC",X"FE",X"FA",X"E5",X"F7",X"37",X"01",X"7C",X"FF",X"7D",X"00",X"B9",X"FF",X"74",X"00",
		X"91",X"08",X"A7",X"F9",X"BC",X"FA",X"36",X"FB",X"7A",X"05",X"9B",X"F6",X"F6",X"00",X"48",X"05",
		X"CE",X"07",X"68",X"FD",X"01",X"FA",X"9C",X"F9",X"99",X"05",X"8D",X"00",X"09",X"F8",X"B5",X"02",
		X"EE",X"06",X"54",X"05",X"0C",X"FC",X"D4",X"F8",X"BE",X"FC",X"1B",X"06",X"2F",X"06",X"E8",X"05",
		X"3C",X"06",X"E0",X"05",X"23",X"06",X"0D",X"06",X"FA",X"FC",X"F4",X"02",X"32",X"08",X"0D",X"FE",
		X"49",X"F9",X"95",X"02",X"C0",X"07",X"98",X"03",X"95",X"FD",X"8A",X"02",X"FD",X"FA",X"23",X"F8",
		X"8A",X"00",X"4F",X"00",X"D5",X"FE",X"D2",X"08",X"04",X"FC",X"06",X"FA",X"59",X"04",X"8B",X"06",
		X"AB",X"05",X"1A",X"06",X"EF",X"05",X"95",X"FC",X"12",X"03",X"6B",X"FC",X"04",X"06",X"53",X"03",
		X"D1",X"F8",X"C9",X"FA",X"6E",X"F9",X"81",X"FA",X"B4",X"F9",X"37",X"FA",X"22",X"03",X"44",X"07",
		X"EA",X"04",X"F7",X"06",X"DE",X"04",X"1C",X"07",X"43",X"FB",X"AF",X"04",X"6A",X"F9",X"78",X"FD",
		X"36",X"02",X"7A",X"FD",X"6E",X"03",X"6E",X"F6",X"05",X"03",X"9E",X"FE",X"81",X"F8",X"80",X"04",
		X"59",X"05",X"F2",X"FB",X"72",X"05",X"92",X"06",X"8F",X"02",X"8C",X"F8",X"D9",X"FB",X"61",X"03",
		X"E9",X"FB",X"A0",X"07",X"CF",X"00",X"E2",X"FD",X"C2",X"07",X"C4",X"04",X"A8",X"06",X"5E",X"05",
		X"2E",X"FD",X"72",X"02",X"3D",X"FC",X"A9",X"F8",X"E6",X"FA",X"C0",X"FB",X"85",X"09",X"E6",X"FD",
		X"3A",X"FC",X"7A",X"04",X"1C",X"08",X"C5",X"FF",X"81",X"FF",X"31",X"01",X"3F",X"F8",X"F5",X"FA",
		X"7F",X"F9",X"64",X"FA",X"DF",X"F9",X"3A",X"FA",X"D3",X"F9",X"21",X"FC",X"39",X"08",X"D8",X"FF",
		X"A4",X"FE",X"2B",X"08",X"6C",X"02",X"AE",X"FC",X"73",X"07",X"6E",X"04",X"F0",X"07",X"7E",X"FD",
		X"50",X"01",X"02",X"07",X"7F",X"05",X"3A",X"05",X"F0",X"FB",X"36",X"04",X"B4",X"F8",X"E4",X"FD",
		X"55",X"07",X"59",X"00",X"FA",X"F7",X"7E",X"02",X"C8",X"FE",X"5A",X"F7",X"B5",X"00",X"E3",X"00",
		X"D6",X"F7",X"93",X"02",X"C1",X"06",X"D4",X"FB",X"35",X"FA",X"87",X"05",X"D2",X"05",X"D9",X"05",
		X"EB",X"05",X"86",X"05",X"B6",X"06",X"FB",X"FE",X"60",X"FF",X"25",X"09",X"64",X"F9",X"8D",X"00",
		X"6D",X"00",X"B0",X"F8",X"AD",X"FA",X"A9",X"F9",X"94",X"03",X"DB",X"06",X"B6",X"04",X"52",X"07",
		X"E5",X"01",X"8F",X"FA",X"4E",X"F8",X"4C",X"01",X"33",X"FF",X"63",X"00",X"9A",X"FF",X"34",X"00",
		X"D2",X"09",X"C1",X"FC",X"D9",X"01",X"C6",X"FE",X"84",X"F8",X"55",X"FB",X"DD",X"02",X"0F",X"FD",
		X"6B",X"03",X"39",X"F9",X"A5",X"FD",X"48",X"07",X"89",X"04",X"60",X"07",X"7E",X"FD",X"97",X"F9",
		X"36",X"FA",X"EF",X"03",X"09",X"FB",X"F6",X"F9",X"F7",X"F9",X"6B",X"FA",X"91",X"F9",X"79",X"FB",
		X"A6",X"03",X"65",X"FA",X"D6",X"FB",X"CE",X"08",X"A6",X"FE",X"9C",X"00",X"C1",X"FF",X"C5",X"FF",
		X"23",X"08",X"64",X"04",X"57",X"06",X"D4",X"FA",X"8C",X"06",X"D6",X"04",X"BC",X"06",X"D2",X"04",
		X"AF",X"06",X"EC",X"04",X"4D",X"05",X"1A",X"F7",X"7C",X"00",X"F9",X"FF",X"FE",X"FE",X"FD",X"06",
		X"A7",X"05",X"6D",X"FD",X"09",X"02",X"11",X"07",X"F8",X"F8",X"1B",X"FD",X"F2",X"02",X"53",X"F9",
		X"C0",X"FA",X"07",X"04",X"E0",X"06",X"DB",X"02",X"31",X"FC",X"AA",X"07",X"73",X"00",X"AC",X"F8",
		X"84",X"00",X"B1",X"07",X"0D",X"FC",X"E2",X"02",X"E9",X"FC",X"30",X"03",X"55",X"FA",X"FF",X"FB",
		X"9C",X"07",X"7A",X"00",X"16",X"FA",X"8D",X"04",X"3D",X"F9",X"36",X"FB",X"63",X"F8",X"BF",X"FF",
		X"E2",X"05",X"A9",X"06",X"5C",X"FD",X"BA",X"01",X"C1",X"06",X"7D",X"FB",X"EA",X"03",X"31",X"FA",
		X"1D",X"FA",X"29",X"FA",X"F0",X"F9",X"73",X"FA",X"9C",X"F9",X"F9",X"FA",X"B9",X"F8",X"DF",X"FE",
		X"BD",X"05",X"18",X"07",X"C3",X"FD",X"9A",X"01",X"54",X"FE",X"E6",X"01",X"D2",X"FC",X"49",X"FA",
		X"92",X"04",X"5B",X"FB",X"6B",X"05",X"89",X"F5",X"47",X"03",X"F4",X"FD",X"65",X"FC",X"9A",X"05",
		X"DF",X"06",X"79",X"00",X"9E",X"F9",X"A7",X"F9",X"1B",X"02",X"9E",X"FE",X"2E",X"F8",X"4F",X"FC",
		X"C2",X"03",X"A3",X"07",X"D0",X"01",X"C6",X"FA",X"A4",X"F8",X"04",X"01",X"F1",X"FF",X"29",X"FF",
		X"5B",X"09",X"3F",X"FF",X"96",X"FF",X"A8",X"01",X"2E",X"F7",X"DA",X"03",X"19",X"FD",X"D5",X"02",
		X"FE",X"06",X"17",X"04",X"1E",X"FA",X"87",X"FC",X"65",X"07",X"14",X"01",X"3C",X"F8",X"C7",X"01",
		X"52",X"FF",X"E3",X"FF",X"88",X"09",X"09",X"FE",X"71",X"00",X"1B",X"06",X"56",X"06",X"B5",X"FC",
		X"C8",X"02",X"F4",X"FC",X"55",X"04",X"78",X"06",X"57",X"03",X"FC",X"F7",X"77",X"00",X"4E",X"00",
		X"B9",X"FE",X"47",X"08",X"C5",X"03",X"66",X"07",X"8D",X"03",X"AD",X"FC",X"AA",X"F7",X"E5",X"03",
		X"96",X"FC",X"67",X"03",X"16",X"06",X"F9",X"04",X"9B",X"F8",X"BE",X"FE",X"43",X"01",X"F5",X"FD",
		X"D5",X"06",X"DF",X"05",X"FA",X"FD",X"50",X"01",X"5E",X"FE",X"23",X"02",X"7F",X"07",X"3B",X"04",
		X"A2",X"06",X"D2",X"04",X"DA",X"FC",X"50",X"F9",X"52",X"06",X"3F",X"03",X"30",X"F9",X"4F",X"FE",
		X"6C",X"02",X"F6",X"F7",X"3A",X"FB",X"EB",X"FF",X"44",X"08",X"58",X"03",X"C7",X"07",X"91",X"02",
		X"21",X"FC",X"02",X"F8",X"5E",X"04",X"68",X"04",X"60",X"FD",X"D5",X"01",X"9C",X"FD",X"D0",X"02",
		X"9A",X"F8",X"58",X"FF",X"E7",X"01",X"DE",X"F6",X"62",X"03",X"2B",X"05",X"A5",X"FD",X"4F",X"01",
		X"84",X"FE",X"3E",X"01",X"C9",X"FD",X"34",X"05",X"44",X"06",X"9E",X"04",X"A6",X"06",X"21",X"04",
		X"7D",X"07",X"28",X"00",X"07",X"FE",X"55",X"07",X"AF",X"FE",X"C4",X"F8",X"2B",X"FB",X"28",X"F9",
		X"45",X"05",X"AD",X"03",X"37",X"FC",X"F8",X"05",X"85",X"02",X"34",X"F8",X"7A",X"FC",X"47",X"02",
		X"8E",X"FB",X"3E",X"F8",X"6B",X"FF",X"50",X"01",X"CB",X"F8",X"F5",X"FA",X"66",X"F9",X"7F",X"02",
		X"CA",X"06",X"D2",X"03",X"08",X"FD",X"91",X"02",X"70",X"FC",X"AC",X"06",X"8E",X"04",X"B2",X"06",
		X"E7",X"02",X"1B",X"FD",X"A8",X"02",X"E9",X"FB",X"C2",X"08",X"B1",X"FD",X"2B",X"00",X"18",X"07",
		X"8D",X"FC",X"8D",X"F9",X"62",X"FA",X"D5",X"FA",X"F3",X"05",X"C7",X"04",X"58",X"06",X"52",X"04",
		X"50",X"07",X"AB",X"FD",X"E2",X"00",X"42",X"04",X"97",X"F7",X"97",X"FF",X"94",X"06",X"E6",X"FE",
		X"C2",X"F8",X"00",X"FB",X"39",X"02",X"39",X"07",X"C3",X"03",X"6F",X"07",X"3C",X"01",X"FF",X"FA",
		X"32",X"F8",X"17",X"01",X"5C",X"FF",X"69",X"F9",X"93",X"F9",X"7D",X"FE",X"F7",X"01",X"2A",X"F8",
		X"69",X"FB",X"5D",X"F9",X"BD",X"FA",X"CA",X"02",X"A0",X"06",X"EA",X"04",X"51",X"04",X"A4",X"FA",
		X"11",X"09",X"E8",X"FD",X"DA",X"00",X"07",X"FF",X"2B",X"00",X"B3",X"FF",X"42",X"F7",X"F5",X"06",
		X"B6",X"FD",X"23",X"01",X"AE",X"FE",X"B8",X"00",X"CC",X"FE",X"F8",X"00",X"55",X"FD",X"6C",X"F7",
		X"02",X"FF",X"05",X"04",X"E6",X"07",X"E5",X"FD",X"8C",X"00",X"E7",X"05",X"EF",X"05",X"CB",X"FB",
		X"8A",X"FA",X"D4",X"F8",X"EF",X"01",X"83",X"FE",X"20",X"F9",X"37",X"03",X"4F",X"FD",X"E0",X"01",
		X"EB",X"FD",X"BC",X"01",X"61",X"FD",X"40",X"06",X"FB",X"05",X"B4",X"FE",X"F1",X"FF",X"6B",X"07",
		X"29",X"04",X"55",X"06",X"C1",X"04",X"CC",X"05",X"61",X"05",X"56",X"FD",X"71",X"01",X"FA",X"FD",
		X"AB",X"01",X"D6",X"FB",X"40",X"F8",X"34",X"FF",X"7C",X"01",X"41",X"F8",X"BF",X"00",X"F9",X"06",
		X"61",X"FC",X"9C",X"02",X"DD",X"05",X"31",X"FA",X"8B",X"FA",X"E8",X"F9",X"74",X"FA",X"09",X"03",
		X"F6",X"05",X"73",X"F9",X"94",X"FB",X"3B",X"F8",X"B7",X"FF",X"8F",X"00",X"15",X"FE",X"08",X"08",
		X"16",X"FD",X"B7",X"F9",X"34",X"03",X"56",X"06",X"EA",X"03",X"85",X"FA",X"36",X"FA",X"38",X"FA",
		X"AF",X"FA",X"7D",X"03",X"37",X"FB",X"92",X"F9",X"09",X"FD",X"A0",X"06",X"57",X"04",X"20",X"07",
		X"BC",X"FD",X"14",X"01",X"E9",X"FE",X"3D",X"F8",X"B2",X"FB",X"16",X"FA",X"98",X"05",X"1F",X"F7",
		X"A6",X"00",X"F8",X"FF",X"AC",X"FB",X"4F",X"02",X"00",X"FE",X"A5",X"01",X"03",X"FE",X"73",X"02",
		X"19",X"F8",X"FB",X"FB",X"BC",X"F8",X"AA",X"03",X"91",X"FC",X"78",X"FA",X"27",X"04",X"6E",X"FB",
		X"6B",X"07",X"01",X"01",X"4C",X"FA",X"1D",X"FA",X"BC",X"FA",X"65",X"FB",X"E8",X"07",X"33",X"00",
		X"17",X"FB",X"A7",X"F8",X"7D",X"02",X"66",X"FE",X"BC",X"F9",X"9A",X"FA",X"C4",X"04",X"12",X"05",
		X"D8",X"06",X"91",X"01",X"DD",X"FD",X"07",X"06",X"4C",X"06",X"B4",X"FE",X"44",X"00",X"4E",X"07",
		X"5D",X"04",X"4D",X"06",X"CF",X"04",X"03",X"06",X"E8",X"04",X"03",X"06",X"01",X"FC",X"10",X"FA",
		X"46",X"FA",X"EA",X"FB",X"68",X"06",X"6F",X"04",X"E0",X"06",X"9C",X"FF",X"A1",X"F9",X"91",X"FA",
		X"89",X"FA",X"BA",X"F9",X"E3",X"FE",X"FE",X"06",X"49",X"04",X"C0",X"06",X"5F",X"FC",X"05",X"03",
		X"70",X"06",X"90",X"03",X"4C",X"FC",X"58",X"04",X"1F",X"F7",X"95",X"01",X"D2",X"FE",X"A5",X"00",
		X"6C",X"FF",X"13",X"F9",X"B7",X"FA",X"E3",X"04",X"60",X"FF",X"18",X"00",X"BF",X"FF",X"2D",X"00",
		X"56",X"FF",X"75",X"01",X"01",X"08",X"68",X"03",X"68",X"05",X"28",X"F6",X"70",X"02",X"23",X"FE",
		X"21",X"01",X"2E",X"FF",X"F8",X"F8",X"44",X"FB",X"BB",X"F9",X"3A",X"FB",X"33",X"F9",X"BF",X"02",
		X"CD",X"FD",X"45",X"02",X"00",X"07",X"88",X"03",X"3E",X"FA",X"67",X"FD",X"FC",X"02",X"DC",X"FB",
		X"E2",X"09",X"BA",X"FB",X"2A",X"03",X"10",X"FD",X"F9",X"02",X"8B",X"05",X"E2",X"FA",X"4D",X"FA",
		X"A8",X"FA",X"36",X"FA",X"0B",X"FB",X"90",X"03",X"15",X"FB",X"13",X"FC",X"91",X"04",X"3E",X"F7",
		X"88",X"01",X"C8",X"FF",X"27",X"FA",X"DF",X"F9",X"23",X"03",X"10",X"FD",X"F9",X"F9",X"61",X"FA",
		X"95",X"FC",X"C4",X"03",X"24",X"F9",X"63",X"04",X"80",X"FB",X"96",X"FA",X"38",X"FA",X"01",X"FD",
		X"54",X"07",X"80",X"00",X"BB",X"F9",X"33",X"FB",X"E3",X"F9",X"E5",X"02",X"D1",X"FD",X"EB",X"F8",
		X"08",X"FD",X"49",X"04",X"24",X"07",X"5B",X"01",X"7A",X"FA",X"C0",X"FA",X"8C",X"06",X"10",X"02",
		X"53",X"FE",X"24",X"02",X"41",X"FD",X"91",X"08",X"D3",X"FD",X"8C",X"FA",X"69",X"FA",X"95",X"03",
		X"3E",X"06",X"0C",X"05",X"0F",X"06",X"E5",X"04",X"8D",X"06",X"30",X"01",X"2C",X"F9",X"F4",X"FC",
		X"1D",X"03",X"4C",X"FC",X"A2",X"07",X"7E",X"03",X"0E",X"08",X"F4",X"FC",X"5E",X"02",X"0B",X"FE",
		X"8B",X"F9",X"BE",X"FB",X"C0",X"03",X"B1",X"FB",X"B0",X"07",X"28",X"00",X"01",X"FF",X"F2",X"05",
		X"24",X"06",X"76",X"02",X"97",X"FD",X"33",X"03",X"13",X"F8",X"04",X"01",X"12",X"06",X"4F",X"05",
		X"1E",X"FE",X"A4",X"F8",X"32",X"FD",X"A2",X"01",X"CC",X"FE",X"26",X"01",X"EF",X"FE",X"51",X"01",
		X"24",X"FE",X"AD",X"07",X"EF",X"03",X"ED",X"06",X"4E",X"01",X"8E",X"F9",X"88",X"FB",X"38",X"F9",
		X"E1",X"02",X"CF",X"FD",X"FE",X"F9",X"0B",X"04",X"75",X"FB",X"DB",X"F9",X"7D",X"FD",X"0C",X"06",
		X"5D",X"05",X"2E",X"05",X"5C",X"06",X"E5",X"FD",X"64",X"01",X"FE",X"06",X"5D",X"04",X"3C",X"06",
		X"B1",X"04",X"FD",X"05",X"D1",X"04",X"70",X"FD",X"9E",X"02",X"8E",X"07",X"6D",X"01",X"62",X"FE",
		X"29",X"02",X"93",X"F9",X"DE",X"FA",X"A5",X"FA",X"03",X"FA",X"98",X"02",X"01",X"06",X"3B",X"05",
		X"17",X"05",X"3C",X"06",X"6C",X"FD",X"EB",X"01",X"C0",X"FD",X"11",X"F9",X"9B",X"FB",X"C7",X"F9",
		X"3E",X"FB",X"14",X"FA",X"FF",X"FA",X"6E",X"FA",X"63",X"FA",X"2F",X"01",X"FD",X"06",X"2C",X"04",
		X"8A",X"06",X"1C",X"04",X"11",X"07",X"C7",X"FC",X"88",X"02",X"F9",X"05",X"5B",X"05",X"F5",X"03",
		X"03",X"FC",X"84",X"06",X"23",X"04",X"DE",X"06",X"5B",X"FF",X"F7",X"F9",X"9F",X"FA",X"C0",X"FA",
		X"4F",X"FA",X"B9",X"04",X"EE",X"03",X"71",X"FC",X"A1",X"05",X"37",X"05",X"78",X"FC",X"EE",X"F9",
		X"05",X"FB",X"10",X"FA",X"F6",X"FC",X"32",X"07",X"1B",X"00",X"44",X"FA",X"15",X"FA",X"B2",X"01",
		X"42",X"06",X"F6",X"04",X"FB",X"04",X"31",X"FB",X"11",X"FA",X"0F",X"FD",X"2D",X"06",X"94",X"04",
		X"F1",X"FB",X"16",X"FA",X"F3",X"FA",X"73",X"FA",X"B5",X"FA",X"D0",X"FA",X"0C",X"FA",X"B1",X"00",
		X"C2",X"06",X"6C",X"04",X"F8",X"05",X"96",X"FB",X"7C",X"05",X"43",X"03",X"AF",X"FA",X"18",X"FA",
		X"8C",X"FE",X"0A",X"07",X"05",X"03",X"6F",X"FB",X"91",X"F9",X"A5",X"FE",X"0D",X"06",X"2C",X"05",
		X"28",X"05",X"F6",X"05",X"06",X"FD",X"A6",X"02",X"72",X"FC",X"3A",X"FB",X"03",X"04",X"98",X"FB",
		X"A4",X"07",X"3C",X"03",X"8B",X"07",X"AB",X"01",X"8F",X"FE",X"CA",X"01",X"D5",X"FA",X"67",X"F9",
		X"F4",X"00",X"36",X"00",X"88",X"F8",X"A9",X"03",X"07",X"FD",X"65",X"03",X"81",X"05",X"F1",X"F8",
		X"CB",X"FE",X"EC",X"01",X"0C",X"FA",X"5D",X"FA",X"3F",X"00",X"17",X"07",X"05",X"02",X"8F",X"F9",
		X"30",X"FF",X"AA",X"06",X"49",X"04",X"67",X"06",X"C9",X"FC",X"3E",X"FA",X"53",X"FB",X"E2",X"04",
		X"70",X"05",X"85",X"03",X"50",X"F8",X"A9",X"00",X"8E",X"00",X"91",X"F9",X"14",X"FB",X"C6",X"FA",
		X"02",X"FA",X"45",X"FF",X"58",X"06",X"29",X"05",X"DB",X"FE",X"07",X"F9",X"70",X"04",X"47",X"FB",
		X"2E",X"FC",X"86",X"03",X"B9",X"FB",X"6A",X"08",X"6A",X"FE",X"F7",X"00",X"5B",X"FF",X"64",X"00",
		X"9C",X"06",X"57",X"05",X"B1",X"00",X"57",X"FE",X"93",X"07",X"F9",X"03",X"A5",X"FE",X"02",X"F9",
		X"00",X"05",X"19",X"FB",X"A2",X"06",X"C1",X"03",X"CE",X"06",X"86",X"03",X"68",X"07",X"CC",X"FD",
		X"F8",X"FA",X"BD",X"F9",X"0B",X"04",X"40",X"FB",X"AF",X"FF",X"14",X"07",X"42",X"FD",X"AB",X"01",
		X"05",X"07",X"F2",X"02",X"C0",X"FD",X"65",X"02",X"FE",X"FA",X"D0",X"F9",X"F7",X"FE",X"CE",X"06",
		X"02",X"FF",X"2F",X"F9",X"13",X"03",X"5A",X"05",X"82",X"FC",X"52",X"03",X"EA",X"FA",X"C9",X"FA",
		X"7E",X"FA",X"98",X"03",X"B9",X"05",X"32",X"04",X"AE",X"F9",X"50",X"FE",X"5E",X"02",X"68",X"F9",
		X"58",X"FB",X"89",X"FA",X"69",X"FA",X"92",X"02",X"CB",X"FD",X"76",X"02",X"10",X"FC",X"94",X"FB",
		X"50",X"06",X"77",X"04",X"86",X"FD",X"4D",X"02",X"5F",X"FD",X"8D",X"03",X"ED",X"F8",X"06",X"00",
		X"59",X"00",X"8C",X"FF",X"8C",X"00",X"42",X"FF",X"E1",X"07",X"7C",X"03",X"0D",X"06",X"50",X"FA",
		X"01",X"FB",X"D2",X"FC",X"E4",X"03",X"07",X"F8",X"B6",X"FD",X"D4",X"01",X"8E",X"FD",X"A7",X"05",
		X"26",X"02",X"41",X"F9",X"D4",X"FB",X"08",X"FA",X"39",X"FB",X"B8",X"01",X"DA",X"06",X"81",X"FA",
		X"FA",X"FB",X"1D",X"F9",X"F8",X"FE",X"7E",X"01",X"F9",X"FD",X"3D",X"06",X"1C",X"FB",X"77",X"05",
		X"56",X"F7",X"AF",X"01",X"E6",X"FE",X"1B",X"01",X"0E",X"FF",X"1F",X"01",X"E5",X"FE",X"A3",X"F9",
		X"42",X"04",X"28",X"FC",X"C1",X"05",X"F5",X"02",X"9C",X"F9",X"26",X"FC",X"31",X"F9",X"2C",X"FE",
		X"70",X"01",X"E6",X"FE",X"6B",X"01",X"38",X"FE",X"EF",X"06",X"66",X"04",X"05",X"06",X"82",X"FD",
		X"FC",X"F9",X"BF",X"04",X"4B",X"FA",X"67",X"FC",X"7C",X"F8",X"D0",X"00",X"98",X"FF",X"A1",X"00",
		X"90",X"FF",X"92",X"00",X"4C",X"06",X"CF",X"05",X"15",X"00",X"B9",X"FF",X"97",X"00",X"5B",X"FF",
		X"0C",X"08",X"43",X"03",X"62",X"06",X"68",X"FA",X"C1",X"07",X"3B",X"00",X"35",X"FF",X"B3",X"04",
		X"00",X"07",X"87",X"FD",X"29",X"02",X"8D",X"FD",X"0C",X"FE",X"72",X"02",X"E0",X"F8",X"95",X"FB",
		X"22",X"01",X"6A",X"FF",X"A1",X"00",X"55",X"FF",X"32",X"01",X"0D",X"FD",X"8E",X"F8",X"10",X"00",
		X"73",X"01",X"13",X"F9",X"A9",X"01",X"BB",X"FF",X"F4",X"F8",X"7B",X"FC",X"40",X"F9",X"CD",X"00",
		X"90",X"06",X"B0",X"FD",X"E8",X"01",X"0B",X"FE",X"20",X"FA",X"EF",X"04",X"FB",X"FA",X"31",X"08",
		X"86",X"FF",X"71",X"FF",X"E9",X"05",X"02",X"05",X"A3",X"05",X"C5",X"FD",X"CE",X"01",X"0E",X"FE",
		X"82",X"F8",X"86",X"02",X"0F",X"05",X"D0",X"05",X"3C",X"FC",X"7A",X"04",X"1E",X"04",X"CD",X"FA",
		X"FB",X"FA",X"00",X"FB",X"85",X"FA",X"60",X"FF",X"AA",X"07",X"CC",X"FC",X"A3",X"02",X"B4",X"FD",
		X"9F",X"02",X"F9",X"FC",X"74",X"05",X"29",X"FE",X"32",X"FA",X"55",X"FB",X"A5",X"04",X"E2",X"03",
		X"6A",X"FB",X"B4",X"F9",X"CA",X"FF",X"B6",X"00",X"6F",X"FF",X"E2",X"00",X"1B",X"FF",X"2A",X"08",
		X"09",X"03",X"12",X"07",X"8F",X"03",X"BB",X"06",X"B3",X"03",X"A3",X"06",X"2C",X"FB",X"40",X"FC",
		X"1C",X"04",X"E7",X"05",X"B8",X"04",X"18",X"03",X"D1",X"F7",X"45",X"02",X"29",X"FF",X"F1",X"F9",
		X"6C",X"02",X"38",X"06",X"4A",X"FB",X"00",X"06",X"FD",X"01",X"3C",X"FE",X"50",X"02",X"01",X"FA",
		X"FD",X"FA",X"58",X"FC",X"9D",X"03",X"0F",X"FA",X"3E",X"FB",X"08",X"FE",X"1C",X"08",X"1D",X"FD",
		X"E3",X"01",X"AC",X"05",X"01",X"05",X"19",X"FC",X"68",X"05",X"70",X"02",X"F1",X"FD",X"38",X"02",
		X"46",X"FD",X"EE",X"06",X"05",X"F9",X"87",X"FE",X"64",X"02",X"9A",X"F9",X"CE",X"FF",X"BA",X"01",
		X"00",X"F8",X"88",X"03",X"8F",X"04",X"12",X"06",X"E7",X"03",X"CD",X"06",X"8A",X"01",X"9E",X"FE",
		X"99",X"01",X"BD",X"FD",X"FC",X"06",X"C0",X"03",X"6B",X"06",X"D8",X"01",X"08",X"FA",X"C6",X"FE",
		X"5B",X"07",X"96",X"FD",X"36",X"01",X"4F",X"06",X"FE",X"FB",X"2F",X"FB",X"00",X"05",X"89",X"03",
		X"B8",X"F9",X"B3",X"FE",X"A8",X"02",X"B8",X"F7",X"0F",X"03",X"BE",X"FD",X"22",X"FD",X"F4",X"05",
		X"D6",X"04",X"CB",X"04",X"EC",X"05",X"85",X"FD",X"E8",X"01",X"C1",X"05",X"9F",X"FB",X"3B",X"FA",
		X"4C",X"FD",X"E0",X"02",X"13",X"FA",X"D3",X"FA",X"52",X"FF",X"9B",X"06",X"10",X"04",X"A9",X"05",
		X"D8",X"04",X"B5",X"01",X"23",X"F8",X"C3",X"02",X"4D",X"FE",X"05",X"FA",X"58",X"FB",X"02",X"FB",
		X"6D",X"05",X"E2",X"02",X"C9",X"FA",X"C3",X"FA",X"60",X"FB",X"F7",X"F9",X"0B",X"01",X"C3",X"05",
		X"F6",X"04",X"F0",X"FC",X"79",X"FA",X"C0",X"FA",X"86",X"00",X"D6",X"06",X"6B",X"FC",X"44",X"FB",
		X"22",X"03",X"FA",X"FC",X"AA",X"03",X"4B",X"F9",X"7F",X"FF",X"C9",X"01",X"EA",X"F8",X"7C",X"01",
		X"BC",X"05",X"B8",X"04",X"74",X"FD",X"A4",X"F9",X"5A",X"FC",X"33",X"F9",X"66",X"03",X"36",X"FD",
		X"E4",X"02",X"C5",X"FC",X"0F",X"05",X"E7",X"02",X"35",X"FB",X"DC",X"F9",X"4B",X"00",X"7B",X"00",
		X"E8",X"FE",X"CA",X"07",X"11",X"FC",X"26",X"03",X"38",X"FD",X"0C",X"03",X"67",X"FB",X"D2",X"FA",
		X"4D",X"FB",X"9C",X"FA",X"47",X"FC",X"40",X"03",X"58",X"FB",X"7B",X"FA",X"5A",X"FE",X"54",X"06",
		X"3C",X"04",X"29",X"06",X"2C",X"FE",X"34",X"FA",X"60",X"03",X"38",X"FD",X"3A",X"03",X"FF",X"FA",
		X"26",X"FD",X"3A",X"06",X"E2",X"FB",X"56",X"FB",X"76",X"FA",X"44",X"FD",X"70",X"05",X"0C",X"05",
		X"08",X"05",X"50",X"05",X"AE",X"04",X"D7",X"05",X"2D",X"FD",X"89",X"02",X"70",X"FD",X"F5",X"03",
		X"5C",X"05",X"53",X"05",X"2A",X"02",X"0D",X"FA",X"16",X"05",X"BE",X"03",X"5F",X"FA",X"1A",X"FE",
		X"F4",X"02",X"8D",X"F8",X"38",X"01",X"5E",X"05",X"F4",X"04",X"1E",X"05",X"DF",X"FC",X"66",X"FA",
		X"6C",X"FB",X"E2",X"FA",X"E4",X"FA",X"A9",X"FD",X"07",X"07",X"9B",X"FF",X"21",X"FA",X"31",X"FD",
		X"9C",X"05",X"B6",X"04",X"30",X"05",X"49",X"05",X"B5",X"FF",X"1F",X"F9",X"A6",X"03",X"E2",X"04",
		X"03",X"05",X"78",X"FA",X"A5",X"FD",X"C1",X"02",X"39",X"FA",X"83",X"FB",X"D9",X"FA",X"0F",X"FB",
		X"99",X"FC",X"47",X"06",X"C1",X"03",X"E3",X"06",X"5F",X"FE",X"F5",X"00",X"A7",X"FF",X"4F",X"F9",
		X"4B",X"FC",X"87",X"FA",X"00",X"06",X"63",X"02",X"A0",X"FB",X"05",X"FA",X"90",X"FF",X"A8",X"05",
		X"04",X"05",X"A0",X"04",X"1F",X"06",X"7F",X"00",X"12",X"FF",X"6F",X"01",X"F6",X"FD",X"E0",X"08",
		X"78",X"FA",X"72",X"05",X"5D",X"02",X"14",X"FF",X"84",X"00",X"C9",X"FF",X"19",X"00",X"14",X"00",
		X"E4",X"FF",X"31",X"00",X"FF",X"FF",X"73",X"F9",X"D8",X"FB",X"FB",X"FA",X"66",X"FA",X"AE",X"01",
		X"FA",X"FE",X"1A",X"01",X"88",X"06",X"E1",X"FA",X"C4",X"FB",X"6B",X"FA",X"6C",X"FD",X"DE",X"06",
		X"80",X"FF",X"01",X"00",X"84",X"00",X"30",X"FF",X"F2",X"07",X"FA",X"FA",X"24",X"05",X"DA",X"03",
		X"B2",X"06",X"D9",X"FC",X"B6",X"02",X"3F",X"05",X"47",X"05",X"7A",X"03",X"72",X"FB",X"40",X"FA",
		X"EE",X"FE",X"4D",X"02",X"89",X"F8",X"13",X"02",X"07",X"05",X"3B",X"05",X"8D",X"04",X"2A",X"05",
		X"47",X"FA",X"E7",X"01",X"EF",X"FE",X"CC",X"F9",X"1D",X"FC",X"99",X"03",X"C1",X"04",X"BE",X"F9",
		X"6D",X"FE",X"17",X"05",X"22",X"05",X"84",X"04",X"BD",X"05",X"32",X"FE",X"4A",X"FA",X"BF",X"FB",
		X"04",X"03",X"24",X"FC",X"A1",X"FA",X"81",X"FB",X"C2",X"FA",X"CC",X"FB",X"32",X"03",X"BD",X"FB",
		X"2E",X"FC",X"DD",X"06",X"40",X"00",X"B9",X"FE",X"58",X"06",X"04",X"04",X"EA",X"05",X"32",X"FD",
		X"DE",X"FA",X"F9",X"03",X"70",X"05",X"45",X"03",X"93",X"FA",X"95",X"FB",X"EF",X"FA",X"A0",X"04",
		X"86",X"04",X"C6",X"05",X"00",X"02",X"9E",X"FA",X"43",X"FB",X"30",X"FB",X"FD",X"FA",X"77",X"FB",
		X"BB",X"FA",X"8F",X"03",X"38",X"05",X"46",X"04",X"21",X"FA",X"8A",X"FE",X"4A",X"02",X"F4",X"F9",
		X"79",X"FC",X"5F",X"04",X"5A",X"05",X"D9",X"02",X"32",X"F9",X"6B",X"00",X"DA",X"04",X"F7",X"05",
		X"71",X"FD",X"49",X"02",X"76",X"FD",X"21",X"FB",X"DC",X"03",X"F9",X"FA",X"49",X"FB",X"61",X"FB",
		X"82",X"FA",X"EB",X"FF",X"31",X"06",X"F9",X"02",X"DD",X"F9",X"A2",X"FF",X"87",X"01",X"E2",X"F9",
		X"A3",X"FB",X"07",X"01",X"98",X"06",X"21",X"FC",X"9F",X"03",X"52",X"FC",X"F0",X"05",X"BF",X"01",
		X"76",X"FD",X"2E",X"07",X"CF",X"FE",X"2F",X"00",X"08",X"05",X"70",X"F8",X"E3",X"00",X"13",X"00",
		X"45",X"FF",X"87",X"06",X"F2",X"03",X"AC",X"05",X"4A",X"04",X"15",X"05",X"74",X"FA",X"D9",X"FD",
		X"9D",X"02",X"71",X"FA",X"51",X"FB",X"F1",X"FE",X"98",X"07",X"89",X"FC",X"2E",X"03",X"BD",X"01",
		X"7D",X"FA",X"CD",X"FA",X"68",X"01",X"45",X"FF",X"C8",X"00",X"B7",X"06",X"15",X"FB",X"DB",X"05",
		X"7B",X"03",X"B8",X"06",X"70",X"00",X"9C",X"FB",X"E1",X"F9",X"DC",X"01",X"24",X"FF",X"0D",X"FA",
		X"EA",X"FB",X"BD",X"FA",X"BE",X"FB",X"8C",X"FA",X"E7",X"01",X"F1",X"05",X"5D",X"FC",X"46",X"04",
		X"D5",X"03",X"46",X"FB",X"D9",X"FA",X"4F",X"FE",X"05",X"06",X"8A",X"04",X"78",X"00",X"BC",X"F8",
		X"33",X"04",X"C7",X"03",X"E9",X"06",X"ED",X"FD",X"AB",X"01",X"9D",X"FE",X"96",X"01",X"43",X"FE",
		X"F8",X"02",X"B7",X"04",X"8C",X"FB",X"40",X"07",X"1D",X"00",X"D0",X"FB",X"CA",X"F9",X"1D",X"02",
		X"AC",X"FE",X"38",X"01",X"3B",X"06",X"55",X"FB",X"AF",X"FB",X"E2",X"FA",X"7D",X"FB",X"05",X"02",
		X"78",X"06",X"BF",X"02",X"20",X"FE",X"21",X"02",X"57",X"FD",X"66",X"06",X"78",X"00",X"59",X"FA",
		X"DE",X"FB",X"C9",X"FA",X"C8",X"FB",X"CF",X"FA",X"E3",X"FB",X"8D",X"FA",X"5A",X"FD",X"06",X"05",
		X"FC",X"04",X"85",X"04",X"C3",X"FC",X"BE",X"04",X"43",X"03",X"AA",X"FA",X"72",X"FB",X"6C",X"FE",
		X"64",X"07",X"EB",X"FD",X"87",X"FB",X"B4",X"FA",X"E8",X"03",X"31",X"04",X"E7",X"FC",X"F6",X"04",
		X"18",X"03",X"D9",X"F9",X"E2",X"04",X"16",X"03",X"31",X"FE",X"C9",X"01",X"68",X"FE",X"0F",X"02",
		X"62",X"FD",X"F4",X"07",X"3B",X"FD",X"B7",X"01",X"B4",X"05",X"CB",X"FC",X"B1",X"03",X"47",X"04",
		X"EB",X"FB",X"EC",X"06",X"1F",X"00",X"FE",X"FE",X"AA",X"05",X"BF",X"04",X"4C",X"03",X"52",X"FA",
		X"27",X"FC",X"1E",X"FA",X"92",X"00",X"8C",X"05",X"BA",X"04",X"11",X"FE",X"88",X"01",X"BD",X"FE",
		X"6C",X"01",X"52",X"FE",X"F8",X"03",X"4F",X"06",X"B9",X"FF",X"47",X"FF",X"27",X"06",X"E9",X"03",
		X"BD",X"05",X"55",X"01",X"25",X"FA",X"2C",X"FC",X"1E",X"FA",X"44",X"02",X"27",X"05",X"48",X"FD",
		X"64",X"02",X"CC",X"FC",X"DD",X"F9",X"89",X"FE",X"AB",X"04",X"56",X"05",X"DE",X"03",X"45",X"06",
		X"41",X"FD",X"BC",X"FD",X"53",X"05",X"CC",X"04",X"41",X"04",X"D3",X"05",X"5A",X"FD",X"2D",X"02",
		X"B2",X"FD",X"24",X"03",X"80",X"04",X"21",X"FA",X"47",X"FE",X"D2",X"02",X"9B",X"F8",X"D2",X"01",
		X"55",X"FF",X"68",X"FA",X"CC",X"01",X"DA",X"06",X"C1",X"FE",X"86",X"00",X"0E",X"00",X"9E",X"F9",
		X"07",X"03",X"1F",X"05",X"69",X"FB",X"0D",X"FC",X"BE",X"F9",X"68",X"FF",X"B2",X"00",X"33",X"FF",
		X"45",X"01",X"C7",X"F9",X"C6",X"FB",X"CD",X"01",X"A8",X"05",X"AD",X"04",X"61",X"00",X"BB",X"F9",
		X"5B",X"FC",X"85",X"FA",X"88",X"03",X"5F",X"FC",X"BA",X"FA",X"3C",X"FD",X"1E",X"05",X"E8",X"04",
		X"81",X"01",X"1C",X"F9",X"22",X"02",X"21",X"FF",X"EC",X"F9",X"C2",X"03",X"8A",X"FC",X"E3",X"04",
		X"01",X"FF",X"7C",X"FA",X"B4",X"FB",X"8B",X"FB",X"40",X"03",X"DC",X"FC",X"0D",X"05",X"57",X"04",
		X"80",X"05",X"F6",X"00",X"B5",X"F9",X"50",X"01",X"B7",X"05",X"91",X"FD",X"C0",X"FA",X"52",X"04",
		X"6E",X"04",X"77",X"05",X"07",X"FE",X"9A",X"FA",X"20",X"FC",X"E6",X"02",X"FE",X"FC",X"04",X"05",
		X"30",X"04",X"BA",X"05",X"6B",X"00",X"B7",X"FA",X"35",X"FB",X"56",X"01",X"E2",X"05",X"F0",X"03",
		X"57",X"05",X"25",X"04",X"33",X"05",X"30",X"04",X"13",X"05",X"BC",X"FC",X"10",X"03",X"C7",X"FB",
		X"F8",X"FA",X"66",X"FD",X"4D",X"06",X"3E",X"00",X"16",X"FA",X"47",X"01",X"D4",X"FF",X"1D",X"F9",
		X"DF",X"04",X"E7",X"02",X"F5",X"FD",X"51",X"03",X"57",X"06",X"89",X"00",X"8E",X"FB",X"00",X"FB",
		X"2E",X"06",X"D3",X"00",X"59",X"FF",X"9D",X"00",X"35",X"FF",X"52",X"01",X"32",X"F9",X"5A",X"02",
		X"56",X"05",X"5A",X"FC",X"05",X"FC",X"13",X"03",X"96",X"FB",X"05",X"FB",X"E3",X"FB",X"7E",X"FA",
		X"3E",X"FD",X"F2",X"01",X"4C",X"FE",X"EA",X"01",X"86",X"FD",X"B7",X"06",X"5A",X"FF",X"32",X"FA",
		X"15",X"02",X"33",X"05",X"9F",X"04",X"F8",X"03",X"B7",X"FC",X"CC",X"04",X"70",X"04",X"DD",X"04",
		X"56",X"04",X"29",X"05",X"D5",X"02",X"29",X"FD",X"7C",X"03",X"B2",X"F8",X"3A",X"01",X"0A",X"00",
		X"11",X"FA",X"C8",X"01",X"B5",X"05",X"00",X"FC",X"3F",X"FC",X"0D",X"03",X"36",X"FB",X"37",X"FD",
		X"4D",X"06",X"38",X"00",X"73",X"FA",X"69",X"00",X"3A",X"06",X"0E",X"03",X"AD",X"06",X"B3",X"FE",
		X"82",X"00",X"1B",X"00",X"8F",X"F9",X"38",X"03",X"30",X"FD",X"85",X"FA",X"31",X"FC",X"2D",X"FA",
		X"B7",X"FE",X"1F",X"02",X"D4",X"F9",X"1A",X"00",X"4A",X"06",X"73",X"FD",X"1B",X"02",X"C3",X"02",
		X"BF",X"F8",X"F4",X"01",X"52",X"FF",X"56",X"FA",X"0B",X"FC",X"1C",X"FB",X"F4",X"03",X"CE",X"FA",
		X"26",X"FE",X"F3",X"01",X"96",X"FD",X"33",X"06",X"A7",X"03",X"66",X"05",X"05",X"04",X"18",X"05",
		X"2E",X"04",X"51",X"FC",X"47",X"FF",X"95",X"06",X"FE",X"02",X"1D",X"06",X"F2",X"02",X"7E",X"06",
		X"59",X"01",X"EA",X"FE",X"46",X"01",X"DF",X"FB",X"CC",X"F9",X"82",X"01",X"01",X"FF",X"83",X"00",
		X"F0",X"05",X"69",X"FC",X"6C",X"FB",X"F2",X"04",X"DC",X"FE",X"60",X"FA",X"A9",X"02",X"1D",X"05",
		X"43",X"FB",X"08",X"FD",X"04",X"04",X"9C",X"05",X"9E",X"00",X"38",X"FE",X"A4",X"06",X"48",X"FE",
		X"04",X"FB",X"63",X"FB",X"AF",X"02",X"EF",X"FC",X"CE",X"FA",X"78",X"FB",X"5E",X"01",X"31",X"FF",
		X"10",X"F9",X"51",X"FE",X"F4",X"00",X"2D",X"FF",X"EE",X"00",X"CD",X"FE",X"FC",X"01",X"1A",X"F9",
		X"2C",X"02",X"FF",X"FE",X"30",X"FA",X"57",X"FC",X"08",X"FB",X"65",X"05",X"44",X"02",X"CC",X"FB",
		X"EF",X"FA",X"1D",X"FC",X"25",X"FB",X"F8",X"05",X"1F",X"01",X"15",X"FF",X"1E",X"01",X"B5",X"FE",
		X"1A",X"02",X"6F",X"F8",X"C8",X"03",X"19",X"FD",X"10",X"03",X"B9",X"04",X"19",X"05",X"78",X"02",
		X"4E",X"FD",X"A1",X"05",X"B0",X"03",X"97",X"FC",X"0C",X"FB",X"83",X"FB",X"5B",X"FD",X"5E",X"06",
		X"11",X"00",X"89",X"FA",X"C6",X"00",X"1D",X"06",X"D6",X"FC",X"02",X"03",X"7C",X"04",X"2D",X"FC",
		X"CA",X"05",X"10",X"01",X"AC",X"FE",X"F3",X"01",X"63",X"FA",X"A1",X"05",X"BA",X"03",X"93",X"03",
		X"9A",X"F8",X"AC",X"01",X"80",X"FF",X"36",X"FB",X"00",X"FB",X"C9",X"02",X"48",X"FD",X"7B",X"FB",
		X"9F",X"04",X"4C",X"04",X"1A",X"05",X"C9",X"01",X"29",X"FA",X"AF",X"FC",X"FC",X"F9",X"E9",X"FE",
		X"45",X"01",X"8C",X"FE",X"4B",X"02",X"EB",X"F8",X"55",X"02",X"79",X"04",X"EB",X"04",X"F4",X"FC",
		X"0D",X"03",X"E1",X"FB",X"C2",X"FB",X"C7",X"FA",X"FF",X"FE",X"42",X"02",X"F4",X"F8",X"7E",X"02",
		X"BF",X"FE",X"CF",X"FA",X"E3",X"FB",X"80",X"FB",X"4B",X"FB",X"9F",X"00",X"4E",X"06",X"B5",X"FC",
		X"0A",X"03",X"03",X"FD",X"A5",X"04",X"BD",X"02",X"8E",X"FB",X"E3",X"FA",X"D6",X"FF",X"69",X"01",
		X"9E",X"F9",X"2E",X"FD",X"09",X"FA",X"C6",X"04",X"DE",X"FF",X"5D",X"FF",X"9C",X"06",X"7C",X"FD",
		X"80",X"FB",X"83",X"FB",X"E4",X"FB",X"46",X"FB",X"46",X"FC",X"8F",X"FA",X"9E",X"FF",X"AC",X"01",
		X"43",X"FA",X"8E",X"FC",X"16",X"FB",X"29",X"FC",X"8B",X"FB",X"DA",X"03",X"57",X"05",X"4D",X"FF",
		X"A5",X"FA",X"6D",X"FC",X"BC",X"02",X"41",X"05",X"DF",X"FA",X"F1",X"FC",X"10",X"FA",X"37",X"00",
		X"3C",X"01",X"BD",X"FA",X"54",X"FC",X"3B",X"FB",X"76",X"02",X"B4",X"05",X"7B",X"03",X"FF",X"FC",
		X"7B",X"FA",X"FC",X"02",X"F1",X"FD",X"69",X"FB",X"83",X"FB",X"7E",X"FD",X"AE",X"02",X"BB",X"FD",
		X"8F",X"03",X"D9",X"F8",X"68",X"02",X"79",X"FF",X"E7",X"FA",X"94",X"02",X"C0",X"05",X"5E",X"03",
		X"C8",X"FD",X"2C",X"04",X"46",X"05",X"21",X"04",X"45",X"05",X"4E",X"FB",X"22",X"FE",X"DF",X"01",
		X"B1",X"FE",X"03",X"02",X"DB",X"FD",X"52",X"07",X"34",X"FE",X"80",X"FB",X"37",X"02",X"C2",X"FE",
		X"1E",X"02",X"C3",X"06",X"59",X"01",X"BE",X"FE",X"81",X"04",X"60",X"05",X"2B",X"03",X"10",X"FD",
		X"12",X"FA",X"F4",X"FF",X"B4",X"00",X"8C",X"FF",X"69",X"01",X"10",X"FA",X"D1",X"FC",X"19",X"FB",
		X"6C",X"FC",X"B4",X"03",X"16",X"04",X"83",X"FC",X"69",X"06",X"D5",X"00",X"1D",X"FC",X"F4",X"02",
		X"AC",X"FD",X"48",X"03",X"A9",X"FA",X"FB",X"FC",X"2B",X"FA",X"BF",X"01",X"B9",X"FF",X"F7",X"FA",
		X"22",X"FC",X"F3",X"02",X"08",X"FD",X"52",X"FC",X"45",X"05",X"2F",X"04",X"76",X"05",X"35",X"01",
		X"5A",X"FA",X"0E",X"FE",X"E6",X"03",X"07",X"06",X"67",X"00",X"38",X"FF",X"CD",X"05",X"28",X"04",
		X"EB",X"04",X"94",X"04",X"A3",X"04",X"5C",X"04",X"8C",X"FB",X"9B",X"FC",X"53",X"FA",X"35",X"00",
		X"B3",X"00",X"31",X"FF",X"15",X"06",X"F1",X"03",X"E5",X"04",X"F0",X"04",X"F5",X"00",X"99",X"FA",
		X"77",X"FC",X"5C",X"FB",X"15",X"FC",X"C2",X"02",X"3E",X"FD",X"33",X"FB",X"2D",X"FC",X"B5",X"FB",
		X"86",X"FB",X"2E",X"FF",X"08",X"06",X"B6",X"03",X"78",X"05",X"E2",X"03",X"64",X"05",X"D6",X"03",
		X"7B",X"05",X"9D",X"03",X"E1",X"05",X"C1",X"FC",X"A6",X"03",X"23",X"04",X"BA",X"05",X"86",X"01",
		X"E2",X"FE",X"C8",X"01",X"45",X"FB",X"1D",X"FB",X"A0",X"01",X"19",X"FF",X"3F",X"01",X"A2",X"05",
		X"83",X"04",X"07",X"00",X"72",X"FF",X"E3",X"06",X"4C",X"FC",X"8D",X"FC",X"A6",X"02",X"52",X"FD",
		X"2C",X"05",X"86",X"01",X"68",X"FE",X"90",X"02",X"2F",X"F9",X"15",X"02",X"E9",X"04",X"1A",X"FE",
		X"CD",X"01",X"FE",X"FD",X"71",X"FA",X"E9",X"FC",X"94",X"FA",X"68",X"03",X"22",X"04",X"5C",X"FD",
		X"DE",X"03",X"10",X"05",X"7B",X"02",X"18",X"FA",X"A2",X"00",X"B4",X"00",X"92",X"FA",X"40",X"FC",
		X"BE",X"01",X"99",X"05",X"CF",X"FB",X"3E",X"FC",X"52",X"FB",X"48",X"FC",X"54",X"FB",X"8F",X"FC",
		X"57",X"03",X"80",X"05",X"62",X"02",X"BA",X"FB",X"80",X"FB",X"11",X"FF",X"96",X"06",X"11",X"FE",
		X"68",X"01",X"67",X"05",X"39",X"04",X"23",X"04",X"DB",X"FC",X"D6",X"04",X"2A",X"04",X"C3",X"04",
		X"40",X"FD",X"D1",X"02",X"24",X"FD",X"28",X"05",X"08",X"02",X"C3",X"FA",X"6C",X"FF",X"37",X"06",
		X"4B",X"FE",X"02",X"01",X"CA",X"05",X"93",X"FC",X"F3",X"03",X"87",X"03",X"AE",X"FB",X"DE",X"FB",
		X"B0",X"FB",X"25",X"FC",X"BC",X"03",X"F2",X"04",X"D0",X"02",X"FA",X"FA",X"9A",X"FC",X"9E",X"FA",
		X"D6",X"00",X"E3",X"04",X"BC",X"04",X"CF",X"FD",X"34",X"02",X"D2",X"FD",X"DE",X"03",X"2B",X"03",
		X"BD",X"FC",X"A0",X"06",X"CB",X"FF",X"C2",X"FB",X"62",X"FB",X"7F",X"FD",X"8E",X"05",X"DB",X"00",
		X"34",X"FE",X"0C",X"07",X"79",X"FD",X"D1",X"01",X"F9",X"04",X"16",X"04",X"FB",X"FC",X"67",X"04",
		X"CB",X"02",X"81",X"FB",X"89",X"FB",X"F5",X"FE",X"E6",X"05",X"36",X"03",X"DE",X"05",X"05",X"01",
		X"1A",X"FC",X"96",X"FA",X"60",X"01",X"70",X"FF",X"58",X"00",X"32",X"06",X"E0",X"FB",X"EB",X"FC",
		X"6F",X"03",X"89",X"05",X"38",X"01",X"7E",X"FE",X"74",X"02",X"60",X"F9",X"F0",X"FD",X"3E",X"F9",
		X"CC",X"00",X"9E",X"FF",X"8D",X"00",X"B4",X"FF",X"7B",X"00",X"E2",X"FF",X"2C",X"FA",X"1E",X"04",
		X"8C",X"03",X"25",X"FD",X"B8",X"03",X"9C",X"F9",X"D9",X"00",X"B4",X"FF",X"6E",X"00",X"DD",X"FF",
		X"37",X"00",X"EF",X"05",X"8F",X"03",X"E1",X"04",X"32",X"04",X"4D",X"04",X"D3",X"04",X"5C",X"FD",
		X"06",X"FC",X"86",X"02",X"0C",X"FE",X"0D",X"02",X"BD",X"FD",X"26",X"05",X"19",X"04",X"44",X"04",
		X"EB",X"04",X"68",X"FE",X"3C",X"FB",X"CC",X"FB",X"1B",X"FC",X"DC",X"FA",X"C5",X"01",X"09",X"FF",
		X"D1",X"FA",X"39",X"03",X"F0",X"FC",X"D3",X"FA",X"6C",X"FE",X"E4",X"01",X"BF",X"FD",X"05",X"06",
		X"21",X"03",X"C2",X"05",X"B5",X"FD",X"C3",X"01",X"64",X"05",X"20",X"03",X"E1",X"FC",X"AF",X"FA",
		X"84",X"02",X"24",X"FE",X"F8",X"01",X"7D",X"FD",X"CF",X"FA",X"C7",X"FC",X"91",X"FA",X"81",X"FF",
		X"6D",X"04",X"2A",X"05",X"9F",X"FE",X"07",X"01",X"49",X"FF",X"6A",X"FA",X"41",X"04",X"4B",X"FB",
		X"C3",X"FC",X"BA",X"FA",X"68",X"03",X"CF",X"03",X"29",X"FD",X"9A",X"FA",X"BA",X"FE",X"C0",X"01",
		X"C7",X"FD",X"74",X"06",X"0A",X"FF",X"BA",X"FB",X"79",X"FB",X"7F",X"02",X"E2",X"FD",X"1D",X"FB",
		X"59",X"FC",X"A5",X"FB",X"EC",X"FB",X"4B",X"02",X"11",X"FE",X"B0",X"FA",X"C6",X"FD",X"34",X"04",
		X"76",X"04",X"D3",X"04",X"B0",X"00",X"77",X"FE",X"49",X"07",X"7B",X"FC",X"31",X"03",X"27",X"FD",
		X"EA",X"03",X"2C",X"03",X"51",X"FC",X"0F",X"FB",X"16",X"FF",X"CD",X"04",X"7A",X"04",X"F1",X"03",
		X"5A",X"05",X"0B",X"01",X"CA",X"FE",X"2B",X"02",X"7D",X"F9",X"32",X"02",X"59",X"04",X"93",X"04",
		X"10",X"04",X"AA",X"04",X"E8",X"03",X"F7",X"04",X"02",X"02",X"32",X"FB",X"49",X"FC",X"6E",X"FB",
		X"69",X"FC",X"F7",X"FA",X"F0",X"FE",X"27",X"02",X"16",X"FA",X"DA",X"00",X"5B",X"05",X"1F",X"FE",
		X"87",X"01",X"71",X"05",X"80",X"FB",X"89",X"FD",X"C9",X"03",X"1D",X"05",X"65",X"01",X"BD",X"FA",
		X"1E",X"00",X"A5",X"05",X"F1",X"01",X"C4",X"FB",X"DC",X"FB",X"F0",X"FB",X"E8",X"FB",X"AF",X"FB",
		X"65",X"01",X"97",X"05",X"34",X"FC",X"0C",X"FD",X"A0",X"02",X"3C",X"FC",X"8C",X"FB",X"85",X"FC",
		X"DE",X"FA",X"EA",X"00",X"6B",X"00",X"4C",X"FA",X"60",X"FD",X"37",X"FA",X"39",X"01",X"E1",X"FF",
		X"DA",X"FF",X"53",X"06",X"C8",X"FC",X"4D",X"03",X"70",X"04",X"AD",X"04",X"A9",X"02",X"FB",X"FC",
		X"C5",X"06",X"CD",X"FE",X"EC",X"00",X"A6",X"FF",X"65",X"00",X"BF",X"05",X"93",X"03",X"9E",X"04",
		X"A6",X"04",X"F1",X"FE",X"CE",X"00",X"7D",X"FF",X"FE",X"F9",X"EB",X"FD",X"FD",X"02",X"39",X"05",
		X"BC",X"03",X"B0",X"02",X"4B",X"F9",X"11",X"02",X"4C",X"FF",X"26",X"FB",X"22",X"02",X"81",X"05",
		X"42",X"00",X"BF",X"FA",X"5E",X"01",X"07",X"05",X"CC",X"03",X"E0",X"FD",X"53",X"02",X"AD",X"FC",
		X"AA",X"FB",X"CA",X"FB",X"63",X"FE",X"E4",X"05",X"A7",X"FF",X"BA",X"FA",X"48",X"02",X"77",X"FE",
		X"C2",X"01",X"1B",X"FE",X"AD",X"03",X"7D",X"FF",X"3B",X"00",X"2F",X"06",X"EB",X"02",X"D3",X"04",
		X"B8",X"FB",X"46",X"06",X"6F",X"00",X"CF",X"FC",X"56",X"FA",X"84",X"01",X"AD",X"FF",X"C6",X"FA",
		X"A4",X"02",X"F3",X"FD",X"EF",X"FA",X"6D",X"FD",X"49",X"04",X"AF",X"FE",X"1E",X"01",X"D6",X"05",
		X"D0",X"FA",X"71",X"FE",X"F4",X"02",X"18",X"06",X"A7",X"FF",X"BD",X"FF",X"90",X"04",X"C0",X"04",
		X"61",X"FE",X"73",X"FB",X"DF",X"02",X"96",X"04",X"12",X"FB",X"8B",X"FE",X"E0",X"01",X"D8",X"FB",
		X"53",X"02",X"64",X"FE",X"A8",X"01",X"51",X"FE",X"E8",X"03",X"55",X"05",X"9E",X"FF",X"BC",X"FF",
		X"30",X"05",X"02",X"04",X"2C",X"FE",X"ED",X"01",X"6C",X"05",X"7A",X"02",X"67",X"FC",X"42",X"FB",
		X"B1",X"FE",X"ED",X"04",X"9E",X"FB",X"78",X"FD",X"3B",X"04",X"A5",X"02",X"C7",X"F9",X"41",X"01",
		X"D5",X"FF",X"7C",X"FB",X"AC",X"FB",X"7C",X"02",X"DA",X"FD",X"A0",X"02",X"22",X"FC",X"8D",X"FD",
		X"53",X"04",X"C7",X"04",X"86",X"00",X"1A",X"FC",X"28",X"03",X"D2",X"FC",X"A5",X"05",X"D5",X"02",
		X"F3",X"05",X"58",X"FE",X"2B",X"01",X"2F",X"FF",X"E0",X"00",X"ED",X"FE",X"80",X"FA",X"08",X"06",
		X"A8",X"00",X"52",X"FF",X"6A",X"01",X"16",X"FB",X"A3",X"FF",X"2A",X"06",X"BA",X"00",X"E9",X"FE",
		X"FF",X"03",X"1F",X"05",X"3E",X"FF",X"B7",X"FB",X"86",X"FB",X"A2",X"02",X"3D",X"04",X"84",X"04",
		X"D3",X"02",X"F7",X"FB",X"42",X"FD",X"61",X"06",X"C1",X"FE",X"B6",X"00",X"D5",X"FF",X"1E",X"FB",
		X"E9",X"FB",X"95",X"FE",X"98",X"05",X"92",X"FF",X"9D",X"FA",X"7E",X"02",X"02",X"FE",X"C2",X"FB",
		X"F7",X"02",X"34",X"FD",X"66",X"04",X"E7",X"03",X"58",X"04",X"F2",X"03",X"4E",X"04",X"E3",X"03",
		X"79",X"04",X"0A",X"FE",X"DE",X"FA",X"B2",X"FF",X"72",X"05",X"97",X"FE",X"65",X"FB",X"27",X"FC",
		X"0E",X"FC",X"83",X"03",X"53",X"04",X"D6",X"03",X"A7",X"04",X"4B",X"01",X"F0",X"FA",X"AF",X"FC",
		X"FD",X"FA",X"FA",X"01",X"B5",X"FE",X"2A",X"01",X"5E",X"06",X"D9",X"FD",X"92",X"01",X"AB",X"FE",
		X"50",X"01",X"A6",X"FE",X"8E",X"01",X"1E",X"FE",X"A9",X"02",X"8B",X"FA",X"FD",X"FF",X"9D",X"00",
		X"C5",X"FE",X"29",X"06",X"A3",X"FD",X"BB",X"FB",X"CB",X"02",X"01",X"04",X"19",X"FC",X"BA",X"FB",
		X"7D",X"01",X"FF",X"04",X"7C",X"FC",X"8A",X"FC",X"0C",X"04",X"C9",X"03",X"C7",X"04",X"FD",X"00",
		X"6C",X"FB",X"C3",X"FB",X"99",X"00",X"18",X"05",X"7F",X"03",X"2D",X"04",X"16",X"FD",X"DB",X"02",
		X"CC",X"FB",X"04",X"FC",X"FF",X"01",X"FE",X"FD",X"4E",X"FB",X"56",X"05",X"50",X"01",X"AD",X"FC",
		X"8E",X"FA",X"D5",X"00",X"CA",X"FF",X"BE",X"FF",X"9A",X"05",X"05",X"03",X"EA",X"04",X"32",X"03",
		X"12",X"05",X"AA",X"01",X"D9",X"FD",X"DA",X"04",X"26",X"03",X"16",X"FD",X"F4",X"FA",X"3E",X"FE",
		X"C6",X"03",X"F8",X"04",X"93",X"FF",X"CE",X"FF",X"A1",X"00",X"04",X"FA",X"69",X"FD",X"0B",X"01",
		X"29",X"FF",X"D0",X"00",X"FA",X"FE",X"88",X"01",X"B3",X"FB",X"3E",X"FC",X"26",X"03",X"95",X"FB",
		X"E5",X"FD",X"69",X"04",X"B7",X"03",X"AC",X"04",X"89",X"FF",X"68",X"FF",X"42",X"06",X"39",X"FC",
		X"85",X"03",X"7B",X"03",X"29",X"04",X"FC",X"F9",X"29",X"00",X"DC",X"FF",X"09",X"00",X"09",X"00",
		X"C5",X"FC",X"52",X"02",X"CE",X"FD",X"6F",X"02",X"48",X"FA",X"C2",X"FC",X"C2",X"FF",X"E7",X"05",
		X"72",X"02",X"73",X"05",X"6E",X"02",X"D8",X"05",X"7D",X"00",X"6E",X"FF",X"85",X"00",X"1D",X"FF",
		X"4B",X"01",X"04",X"FA",X"88",X"FD",X"18",X"FA",X"8F",X"00",X"F6",X"FF",X"66",X"FF",X"38",X"05",
		X"6A",X"03",X"65",X"FE",X"64",X"01",X"C8",X"FD",X"9C",X"FB",X"7A",X"05",X"59",X"02",X"FB",X"05",
		X"CC",X"FE",X"2C",X"00",X"3E",X"04",X"60",X"04",X"76",X"01",X"5B",X"FB",X"2C",X"FC",X"D5",X"FB",
		X"0F",X"FC",X"C4",X"FB",X"0A",X"02",X"FB",X"FD",X"42",X"FB",X"4B",X"05",X"E6",X"00",X"EE",X"FE",
		X"7D",X"01",X"38",X"FB",X"01",X"FC",X"34",X"00",X"84",X"05",X"0E",X"FD",X"3D",X"FC",X"3E",X"FB",
		X"81",X"00",X"A0",X"04",X"D0",X"03",X"07",X"FE",X"3B",X"FB",X"73",X"FC",X"6A",X"FC",X"19",X"05",
		X"37",X"01",X"CE",X"FB",X"03",X"FC",X"1D",X"FC",X"EF",X"FB",X"2A",X"FC",X"F3",X"FB",X"50",X"FC",
		X"30",X"03",X"39",X"04",X"1F",X"04",X"BF",X"FE",X"F4",X"FA",X"DA",X"03",X"C8",X"02",X"EB",X"FD",
		X"46",X"02",X"1B",X"FD",X"42",X"06",X"BA",X"FE",X"B5",X"00",X"A4",X"FF",X"21",X"00",X"9F",X"05",
		X"9A",X"02",X"2D",X"FE",X"C7",X"02",X"AA",X"04",X"87",X"03",X"57",X"FE",X"BE",X"01",X"A0",X"04",
		X"AE",X"FB",X"25",X"06",X"B0",X"FF",X"9E",X"FF",X"95",X"03",X"29",X"05",X"F3",X"FD",X"8D",X"01",
		X"77",X"FE",X"7C",X"01",X"40",X"FE",X"15",X"02",X"33",X"FC",X"11",X"FC",X"E7",X"FB",X"0C",X"03",
		X"F2",X"03",X"44",X"04",X"3A",X"02",X"89",X"FB",X"5C",X"FC",X"8A",X"FB",X"CD",X"FF",X"A7",X"05",
		X"4C",X"FD",X"35",X"02",X"78",X"FD",X"5E",X"FC",X"B1",X"02",X"2A",X"FD",X"B6",X"04",X"60",X"03",
		X"09",X"04",X"AD",X"FC",X"4B",X"04",X"29",X"03",X"02",X"05",X"61",X"00",X"F2",X"FB",X"51",X"FB",
		X"56",X"01",X"2E",X"FF",X"E9",X"FA",X"EC",X"FC",X"BA",X"02",X"71",X"04",X"8C",X"03",X"05",X"04",
		X"19",X"04",X"F3",X"00",X"B4",X"FA",X"12",X"FD",X"D0",X"FA",X"21",X"FF",X"CA",X"01",X"1B",X"FA",
		X"94",X"01",X"07",X"FF",X"A7",X"00",X"65",X"FF",X"86",X"00",X"5D",X"FF",X"BC",X"00",X"E6",X"FE",
		X"C0",X"01",X"13",X"FB",X"CB",X"FF",X"21",X"01",X"F6",X"FA",X"76",X"06",X"68",X"FF",X"C8",X"FF",
		X"93",X"03",X"F4",X"04",X"57",X"FE",X"11",X"FC",X"A4",X"FB",X"24",X"03",X"1C",X"FC",X"C4",X"FD",
		X"DE",X"01",X"B5",X"FD",X"1D",X"05",X"6D",X"00",X"D8",X"FA",X"F6",X"00",X"E7",X"04",X"19",X"01",
		X"F3",X"FD",X"A7",X"05",X"5B",X"02",X"89",X"05",X"2F",X"FD",X"98",X"FC",X"C8",X"01",X"05",X"05",
		X"13",X"FA",X"F3",X"FF",X"C1",X"FF",X"45",X"00",X"93",X"FF",X"63",X"00",X"AB",X"FF",X"A5",X"FB",
		X"5A",X"FB",X"03",X"00",X"25",X"00",X"C2",X"FF",X"6A",X"00",X"8C",X"FA",X"01",X"FD",X"40",X"02",
		X"EA",X"03",X"D0",X"FC",X"6C",X"03",X"3E",X"FA",X"F3",X"FF",X"A1",X"03",X"B7",X"04",X"DD",X"FE",
		X"B8",X"FB",X"09",X"FC",X"FC",X"02",X"EA",X"00",X"C0",X"FA",X"1A",X"FD",X"4A",X"FB",X"0A",X"FD",
		X"84",X"01",X"C7",X"FE",X"6C",X"01",X"35",X"FD",X"B8",X"FA",X"22",X"00",X"C6",X"00",X"5C",X"FB",
		X"87",X"FC",X"06",X"FC",X"45",X"FC",X"2D",X"FC",X"3A",X"FC",X"31",X"FC",X"51",X"FC",X"04",X"FC",
		X"3C",X"02",X"44",X"FE",X"2A",X"02",X"B2",X"FC",X"5E",X"FD",X"D0",X"04",X"9D",X"03",X"97",X"01",
		X"06",X"FA",X"38",X"02",X"98",X"03",X"A5",X"04",X"BC",X"FC",X"12",X"FD",X"24",X"03",X"D7",X"04",
		X"FA",X"FD",X"16",X"FC",X"BB",X"02",X"A0",X"04",X"2F",X"03",X"07",X"05",X"DF",X"00",X"7D",X"FE",
		X"49",X"05",X"A7",X"FF",X"16",X"FB",X"F3",X"01",X"47",X"04",X"C9",X"03",X"E5",X"03",X"F7",X"03",
		X"B6",X"03",X"32",X"04",X"A9",X"FD",X"CD",X"FB",X"58",X"FC",X"30",X"FC",X"F3",X"FB",X"1E",X"FE",
		X"2C",X"05",X"3C",X"00",X"0E",X"FB",X"6B",X"01",X"8C",X"FF",X"B0",X"FA",X"FF",X"03",X"75",X"02",
		X"6C",X"FE",X"AE",X"01",X"03",X"FE",X"B6",X"04",X"00",X"03",X"D0",X"FD",X"86",X"02",X"DC",X"FB",
		X"B4",X"FC",X"75",X"FB",X"C3",X"FF",X"F9",X"04",X"1F",X"FF",X"26",X"FB",X"BD",X"02",X"B0",X"FD",
		X"12",X"03",X"57",X"03",X"98",X"FB",X"41",X"FE",X"FF",X"04",X"58",X"00",X"A1",X"FB",X"62",X"FC",
		X"6D",X"FD",X"04",X"05",X"C2",X"02",X"72",X"05",X"6E",X"FE",X"30",X"01",X"16",X"FF",X"07",X"01",
		X"E9",X"FE",X"04",X"02",X"50",X"04",X"89",X"FA",X"7E",X"FF",X"49",X"03",X"12",X"05",X"1E",X"FF",
		X"4B",X"FD",X"AA",X"02",X"58",X"FB",X"E6",X"FC",X"A4",X"FB",X"F3",X"FC",X"42",X"FB",X"5A",X"02",
		X"28",X"FE",X"54",X"02",X"D4",X"03",X"DF",X"FC",X"C8",X"04",X"7C",X"01",X"BD",X"FB",X"C4",X"FC",
		X"6E",X"FB",X"57",X"01",X"8F",X"FF",X"03",X"FB",X"48",X"FD",X"38",X"FB",X"B3",X"00",X"DB",X"04",
		X"36",X"FE",X"79",X"01",X"20",X"05",X"51",X"02",X"19",X"FE",X"95",X"03",X"18",X"04",X"E2",X"03",
		X"5D",X"01",X"32",X"FA",X"25",X"02",X"40",X"03",X"47",X"05",X"7F",X"FF",X"56",X"00",X"DE",X"FF",
		X"3A",X"00",X"DF",X"FF",X"50",X"00",X"79",X"FF",X"EC",X"F9",X"76",X"FF",X"8F",X"00",X"69",X"FF",
		X"35",X"01",X"DE",X"FB",X"F3",X"FB",X"02",X"01",X"E4",X"FF",X"8F",X"FA",X"42",X"04",X"DA",X"FF",
		X"19",X"FC",X"F2",X"FB",X"C8",X"01",X"5B",X"04",X"37",X"FD",X"62",X"FC",X"8F",X"04",X"B4",X"01",
		X"AC",X"FC",X"4C",X"FB",X"91",X"00",X"62",X"00",X"88",X"FB",X"72",X"FC",X"07",X"02",X"24",X"04",
		X"20",X"FD",X"7B",X"FB",X"D2",X"01",X"D6",X"FE",X"64",X"01",X"B5",X"FE",X"FE",X"01",X"BA",X"FC",
		X"DA",X"FD",X"BD",X"02",X"ED",X"FA",X"89",X"FD",X"1E",X"FB",X"90",X"01",X"35",X"04",X"D5",X"03",
		X"BA",X"FD",X"BE",X"FB",X"94",X"FD",X"05",X"04",X"DD",X"FE",X"5F",X"FB",X"87",X"03",X"AB",X"FC",
		X"26",X"05",X"AE",X"00",X"C8",X"FF",X"6F",X"00",X"EB",X"FF",X"57",X"00",X"F6",X"FF",X"6F",X"00",
		X"8E",X"FA",X"CC",X"03",X"79",X"FC",X"CA",X"FC",X"0E",X"FC",X"C1",X"FC",X"2C",X"FC",X"D4",X"FC",
		X"9F",X"03",X"BE",X"02",X"BF",X"FD",X"26",X"03",X"37",X"FA",X"23",X"01",X"7E",X"03",X"F1",X"04",
		X"E3",X"FD",X"23",X"02",X"32",X"04",X"19",X"04",X"AD",X"02",X"9C",X"FD",X"CF",X"04",X"34",X"01",
		X"89",X"FB",X"3B",X"FD",X"52",X"FB",X"29",X"FF",X"57",X"01",X"84",X"FE",X"0B",X"05",X"3E",X"03",
		X"49",X"04",X"B4",X"03",X"86",X"FE",X"58",X"FB",X"EE",X"FD",X"E6",X"01",X"42",X"FE",X"A8",X"02",
		X"BB",X"FA",X"97",X"00",X"40",X"03",X"E3",X"FC",X"99",X"FB",X"77",X"FF",X"3B",X"01",X"90",X"FE",
		X"A6",X"05",X"8D",X"02",X"26",X"05",X"3C",X"FD",X"AE",X"02",X"9D",X"FD",X"13",X"03",X"69",X"FB",
		X"33",X"FF",X"9F",X"03",X"C3",X"04",X"87",X"FF",X"59",X"FC",X"B9",X"FB",X"78",X"FF",X"1D",X"01",
		X"BA",X"FE",X"62",X"05",X"E5",X"02",X"8A",X"04",X"59",X"03",X"F3",X"03",X"27",X"FD",X"02",X"04",
		X"71",X"02",X"7A",X"FB",X"60",X"FF",X"27",X"04",X"30",X"04",X"34",X"FF",X"58",X"00",X"7C",X"05",
		X"6E",X"00",X"8A",X"FB",X"C2",X"00",X"5D",X"00",X"8F",X"FA",X"74",X"03",X"CD",X"FC",X"80",X"FD",
		X"18",X"02",X"F0",X"FD",X"36",X"04",X"D6",X"03",X"24",X"01",X"E6",X"FA",X"CE",X"FD",X"C4",X"FA",
		X"DB",X"03",X"DE",X"FF",X"17",X"00",X"91",X"00",X"4E",X"FB",X"09",X"FD",X"24",X"FC",X"FA",X"02",
		X"99",X"03",X"CB",X"FC",X"63",X"05",X"21",X"00",X"F1",X"FF",X"7A",X"00",X"62",X"FF",X"06",X"05",
		X"28",X"03",X"22",X"04",X"9E",X"03",X"C5",X"03",X"E7",X"03",X"72",X"03",X"49",X"04",X"7C",X"FD",
		X"BF",X"FC",X"5F",X"02",X"17",X"FD",X"95",X"FB",X"EB",X"FE",X"EF",X"03",X"F2",X"03",X"4B",X"03",
		X"8F",X"04",X"30",X"FE",X"50",X"FC",X"19",X"FC",X"08",X"FD",X"4F",X"FB",X"06",X"02",X"9D",X"FE",
		X"2F",X"FC",X"27",X"02",X"95",X"FE",X"58",X"01",X"FF",X"FE",X"25",X"01",X"04",X"FF",X"56",X"01",
		X"5C",X"FE",X"54",X"06",X"F1",X"FC",X"8E",X"02",X"DC",X"FD",X"62",X"02",X"E7",X"FC",X"1F",X"FC",
		X"85",X"01",X"A3",X"04",X"0F",X"03",X"00",X"04",X"41",X"FB",X"4C",X"FF",X"05",X"01",X"AB",X"FE",
		X"A6",X"04",X"43",X"03",X"FF",X"03",X"87",X"03",X"CE",X"03",X"B8",X"FD",X"BA",X"02",X"82",X"03",
		X"4A",X"FB",X"0F",X"FF",X"76",X"03",X"3D",X"FE",X"7F",X"01",X"8A",X"FE",X"E1",X"02",X"03",X"05",
		X"B0",X"FF",X"F8",X"FF",X"90",X"00",X"46",X"FB",X"FE",X"FC",X"13",X"FC",X"CB",X"FC",X"BD",X"02",
		X"36",X"FC",X"57",X"FE",X"03",X"02",X"D4",X"FB",X"7F",X"FC",X"5A",X"FD",X"34",X"02",X"09",X"FE",
		X"53",X"02",X"36",X"FD",X"97",X"06",X"8A",X"FD",X"FA",X"01",X"67",X"FE",X"C2",X"01",X"F9",X"FD",
		X"7A",X"FC",X"B9",X"03",X"E4",X"03",X"E7",X"01",X"B8",X"FB",X"CA",X"FC",X"E5",X"FC",X"1A",X"03",
		X"5C",X"FB",X"26",X"FF",X"FF",X"03",X"8C",X"03",X"0C",X"04",X"72",X"FF",X"44",X"FB",X"D2",X"02",
		X"59",X"03",X"B1",X"FD",X"4A",X"03",X"C4",X"03",X"DB",X"03",X"8C",X"01",X"F4",X"FA",X"B0",X"00",
		X"56",X"04",X"DB",X"01",X"7C",X"FD",X"D4",X"05",X"A2",X"FE",X"CA",X"00",X"CC",X"FF",X"60",X"FB",
		X"1F",X"FD",X"E1",X"FB",X"70",X"FD",X"25",X"03",X"33",X"04",X"AA",X"01",X"B3",X"FB",X"22",X"FD",
		X"8A",X"FB",X"3F",X"01",X"E2",X"03",X"1F",X"04",X"98",X"00",X"BE",X"FE",X"46",X"05",X"65",X"02",
		X"DD",X"04",X"19",X"FD",X"C0",X"02",X"B4",X"FC",X"E3",X"FC",X"92",X"FB",X"36",X"FF",X"9A",X"01",
		X"2A",X"FB",X"76",X"00",X"A7",X"04",X"6F",X"FE",X"F1",X"FB",X"ED",X"02",X"14",X"01",X"89",X"FA",
		X"62",X"02",X"63",X"FE",X"56",X"FC",X"26",X"FC",X"B9",X"FD",X"D1",X"01",X"6A",X"FE",X"18",X"02",
		X"B0",X"FB",X"BD",X"FC",X"82",X"FF",X"86",X"05",X"84",X"FD",X"26",X"02",X"13",X"FE",X"DF",X"02",
		X"8B",X"00",X"B9",X"FA",X"DA",X"02",X"C9",X"FD",X"B7",X"02",X"3B",X"03",X"B8",X"FC",X"26",X"FC",
		X"89",X"FE",X"62",X"04",X"2C",X"03",X"46",X"04",X"5E",X"FF",X"72",X"FB",X"97",X"02",X"EB",X"FD",
		X"70",X"02",X"81",X"FC",X"FF",X"00",X"5E",X"04",X"3B",X"03",X"AD",X"FD",X"80",X"FC",X"4B",X"04",
		X"A3",X"01",X"DA",X"FD",X"63",X"05",X"26",X"FF",X"5A",X"00",X"5A",X"00",X"F1",X"FA",X"E0",X"02",
		X"87",X"03",X"BF",X"03",X"A3",X"03",X"92",X"02",X"A6",X"FB",X"B3",X"02",X"67",X"03",X"F2",X"FC",
		X"6A",X"FC",X"7B",X"FC",X"BB",X"FC",X"EC",X"FB",X"0F",X"00",X"01",X"01",X"A3",X"FA",X"8F",X"02",
		X"5A",X"03",X"53",X"FE",X"07",X"02",X"F4",X"04",X"1D",X"01",X"9F",X"FE",X"F4",X"03",X"81",X"03",
		X"BB",X"03",X"9B",X"02",X"16",X"FD",X"85",X"05",X"4C",X"FF",X"43",X"00",X"5A",X"00",X"8A",X"FB",
		X"FF",X"FC",X"43",X"FC",X"CC",X"FC",X"3B",X"03",X"A5",X"02",X"71",X"FD",X"BA",X"04",X"BC",X"00",
		X"05",X"FC",X"DD",X"FC",X"30",X"FC",X"0B",X"FD",X"AB",X"FB",X"E0",X"FF",X"18",X"01",X"52",X"FB",
		X"6E",X"FD",X"CE",X"FB",X"78",X"02",X"F8",X"03",X"CC",X"02",X"E0",X"FD",X"72",X"02",X"29",X"FD",
		X"E9",X"05",X"BD",X"FE",X"BF",X"00",X"90",X"02",X"F7",X"FD",X"A6",X"02",X"8F",X"FA",X"42",X"01",
		X"A6",X"FF",X"FE",X"FF",X"09",X"05",X"77",X"02",X"BB",X"FE",X"DD",X"FA",X"3D",X"FF",X"AF",X"00",
		X"7D",X"FF",X"D6",X"00",X"EA",X"FE",X"BC",X"04",X"E8",X"02",X"37",X"04",X"8F",X"01",X"48",X"FB",
		X"99",X"00",X"84",X"00",X"08",X"FB",X"68",X"02",X"5B",X"FE",X"A0",X"01",X"70",X"FE",X"B2",X"02",
		X"44",X"04",X"CD",X"02",X"A9",X"04",X"E1",X"FF",X"78",X"FC",X"0B",X"FC",X"A8",X"01",X"BC",X"03",
		X"01",X"04",X"36",X"00",X"FA",X"FB",X"85",X"FC",X"79",X"01",X"E4",X"FE",X"A9",X"FB",X"25",X"04",
		X"D0",X"01",X"2A",X"FE",X"F5",X"03",X"35",X"03",X"1F",X"04",X"E7",X"FF",X"AD",X"FB",X"35",X"FD",
		X"F3",X"FB",X"2A",X"03",X"A8",X"00",X"1A",X"FB",X"EA",X"01",X"CF",X"FE",X"33",X"01",X"B2",X"04",
		X"92",X"02",X"9A",X"04",X"57",X"01",X"D8",X"FC",X"E0",X"FB",X"C8",X"FF",X"79",X"04",X"3C",X"FF",
		X"98",X"FB",X"6C",X"02",X"A6",X"03",X"7B",X"03",X"BD",X"03",X"66",X"FF",X"6D",X"FB",X"8E",X"FD",
		X"80",X"FB",X"50",X"FE",X"7A",X"01",X"6D",X"FD",X"4D",X"FB",X"51",X"00",X"7B",X"00",X"31",X"FC",
		X"45",X"FC",X"BB",X"01",X"AC",X"FE",X"CD",X"01",X"D2",X"03",X"D8",X"FC",X"B4",X"04",X"A5",X"FD",
		X"3B",X"02",X"9F",X"03",X"EC",X"03",X"F3",X"01",X"5D",X"FE",X"E6",X"01",X"AC",X"FD",X"BD",X"05",
		X"90",X"FE",X"E1",X"FC",X"12",X"FC",X"42",X"FD",X"CA",X"FB",X"0E",X"FE",X"90",X"01",X"68",X"FE",
		X"84",X"03",X"CB",X"03",X"D9",X"02",X"9B",X"FD",X"96",X"FB",X"29",X"FF",X"1B",X"01",X"CD",X"FE",
		X"F7",X"01",X"45",X"FA",X"96",X"02",X"3B",X"FE",X"B4",X"01",X"7A",X"FE",X"33",X"02",X"77",X"04",
		X"7C",X"01",X"30",X"FE",X"61",X"04",X"DC",X"02",X"20",X"04",X"C8",X"02",X"7C",X"04",X"AC",X"00",
		X"9E",X"FE",X"EE",X"04",X"FC",X"FE",X"23",X"00",X"CA",X"04",X"4A",X"02",X"18",X"FF",X"9B",X"00",
		X"95",X"FF",X"5E",X"00",X"B1",X"FF",X"65",X"00",X"65",X"FF",X"4A",X"03",X"79",X"FD",X"AC",X"03",
		X"B2",X"03",X"F1",X"00",X"CC",X"FB",X"FA",X"FC",X"60",X"FC",X"AF",X"FC",X"B4",X"FC",X"F3",X"01",
		X"6B",X"FE",X"A2",X"01",X"21",X"FE",X"CA",X"03",X"4C",X"03",X"7A",X"03",X"8C",X"03",X"88",X"02",
		X"DC",X"FB",X"DF",X"FE",X"E5",X"03",X"69",X"03",X"49",X"00",X"ED",X"FA",X"90",X"02",X"E1",X"FD",
		X"58",X"02",X"42",X"03",X"4B",X"FC",X"28",X"FE",X"79",X"02",X"A6",X"FA",X"20",X"01",X"7E",X"FF",
		X"0F",X"00",X"67",X"04",X"08",X"03",X"AF",X"01",X"91",X"FA",X"D6",X"01",X"CD",X"FE",X"E2",X"00",
		X"42",X"04",X"EE",X"02",X"53",X"03",X"15",X"FC",X"38",X"FE",X"DD",X"03",X"3F",X"01",X"15",X"FB",
		X"20",X"01",X"B4",X"FF",X"A4",X"FB",X"3E",X"FD",X"0B",X"FC",X"3B",X"FD",X"C6",X"FB",X"52",X"01",
		X"BD",X"03",X"68",X"03",X"FF",X"02",X"CF",X"FD",X"66",X"02",X"EF",X"FB",X"04",X"FF",X"BB",X"01",
		X"37",X"FB",X"D8",X"FD",X"36",X"FB",X"82",X"02",X"DE",X"FD",X"E4",X"FC",X"B6",X"FB",X"51",X"01",
		X"30",X"FF",X"BB",X"00",X"5B",X"04",X"16",X"FD",X"77",X"FC",X"CF",X"FD",X"6B",X"02",X"CB",X"FB",
		X"6D",X"FD",X"CB",X"FB",X"7D",X"00",X"4E",X"04",X"91",X"FE",X"2C",X"FC",X"01",X"FD",X"D5",X"FC",
		X"AD",X"03",X"FF",X"02",X"15",X"04",X"85",X"FD",X"33",X"FD",X"FB",X"01",X"4A",X"FE",X"34",X"02",
		X"DA",X"FB",X"3A",X"FF",X"9C",X"04",X"6F",X"FF",X"59",X"FC",X"AC",X"FC",X"DB",X"01",X"FF",X"03",
		X"1F",X"03",X"AE",X"03",X"3C",X"03",X"9D",X"03",X"1D",X"03",X"2D",X"FE",X"C4",X"01",X"22",X"FE",
		X"65",X"03",X"A8",X"03",X"3A",X"01",X"57",X"FB",X"BA",X"00",X"1A",X"04",X"87",X"FE",X"16",X"01",
		X"72",X"04",X"FC",X"FB",X"8F",X"FE",X"8B",X"01",X"C3",X"FC",X"95",X"01",X"54",X"04",X"9A",X"FB",
		X"40",X"FF",X"81",X"00",X"B2",X"FF",X"5C",X"00",X"AE",X"FF",X"AC",X"00",X"9A",X"FB",X"1D",X"FD",
		X"9D",X"01",X"BE",X"03",X"7A",X"FD",X"8D",X"02",X"54",X"FC",X"09",X"FD",X"75",X"FC",X"1B",X"FD",
		X"39",X"03",X"42",X"02",X"E7",X"FD",X"C5",X"02",X"79",X"FA",X"93",X"01",X"34",X"FF",X"75",X"00",
		X"37",X"04",X"FB",X"02",X"A4",X"03",X"38",X"03",X"80",X"03",X"3C",X"03",X"A5",X"03",X"57",X"01",
		X"5A",X"FB",X"97",X"FE",X"0A",X"01",X"18",X"FF",X"08",X"01",X"B2",X"FE",X"29",X"04",X"5C",X"03",
		X"2F",X"FF",X"7F",X"00",X"95",X"FF",X"F2",X"FA",X"C3",X"FE",X"F1",X"00",X"FD",X"FE",X"88",X"01",
		X"24",X"FC",X"0D",X"FD",X"68",X"FC",X"22",X"FD",X"11",X"FC",X"16",X"FF",X"93",X"03",X"D9",X"03",
		X"66",X"FF",X"16",X"00",X"92",X"04",X"90",X"02",X"EA",X"03",X"0C",X"03",X"B7",X"02",X"35",X"FD",
		X"B9",X"04",X"F8",X"01",X"0A",X"05",X"57",X"FE",X"2A",X"01",X"25",X"FF",X"11",X"FC",X"EC",X"FC",
		X"BF",X"FC",X"53",X"FC",X"EC",X"00",X"FD",X"03",X"F8",X"02",X"87",X"03",X"4A",X"03",X"92",X"02",
		X"3E",X"FC",X"2D",X"FD",X"0D",X"FC",X"A5",X"FF",X"6F",X"04",X"E5",X"FE",X"63",X"FC",X"91",X"FC",
		X"08",X"FF",X"53",X"04",X"A2",X"02",X"DC",X"03",X"E2",X"02",X"B2",X"FE",X"8A",X"FB",X"31",X"FE",
		X"79",X"02",X"23",X"03",X"8C",X"FA",X"21",X"01",X"41",X"FF",X"9A",X"00",X"AD",X"FF",X"2A",X"FC",
		X"AE",X"FC",X"E4",X"02",X"17",X"00",X"56",X"FF",X"FC",X"04",X"9A",X"FD",X"E7",X"01",X"08",X"FE",
		X"27",X"FC",X"24",X"FD",X"47",X"FD",X"28",X"05",X"3D",X"FF",X"75",X"00",X"CE",X"FF",X"FA",X"FF",
		X"5F",X"04",X"B9",X"02",X"A8",X"03",X"D2",X"02",X"6D",X"FC",X"48",X"01",X"15",X"FF",X"FE",X"00",
		X"25",X"04",X"A0",X"FC",X"70",X"04",X"AA",X"00",X"FB",X"FE",X"46",X"03",X"FB",X"03",X"1C",X"FF",
		X"70",X"00",X"CE",X"FF",X"59",X"FB",X"C2",X"FD",X"D2",X"FB",X"A9",X"FD",X"AD",X"FB",X"41",X"02",
		X"FC",X"02",X"5A",X"FE",X"EE",X"01",X"A1",X"04",X"7B",X"00",X"7B",X"FF",X"A2",X"00",X"2D",X"FF",
		X"4C",X"01",X"9A",X"FA",X"C9",X"02",X"CC",X"FD",X"1D",X"02",X"71",X"FD",X"7A",X"FC",X"DF",X"FD",
		X"07",X"04",X"8E",X"02",X"10",X"04",X"49",X"02",X"9C",X"04",X"5A",X"00",X"9D",X"FF",X"7E",X"00",
		X"22",X"FF",X"28",X"04",X"D8",X"02",X"5B",X"03",X"49",X"03",X"F8",X"02",X"B2",X"03",X"E9",X"01",
		X"0B",X"FD",X"32",X"FC",X"75",X"FD",X"A7",X"FB",X"B5",X"FE",X"9C",X"00",X"99",X"FF",X"2D",X"00",
		X"EC",X"FF",X"E4",X"FF",X"36",X"00",X"95",X"FF",X"90",X"00",X"22",X"FF",X"3D",X"01",X"AB",X"FD",
		X"87",X"FD",X"ED",X"01",X"35",X"FE",X"CB",X"01",X"D7",X"FD",X"4F",X"05",X"91",X"01",X"B9",X"04",
		X"9F",X"01",X"24",X"05",X"62",X"FE",X"0D",X"01",X"F6",X"FE",X"D4",X"00",X"EC",X"FE",X"F8",X"FB",
		X"66",X"03",X"AB",X"02",X"E3",X"03",X"16",X"01",X"57",X"FC",X"E6",X"FC",X"A5",X"FC",X"B5",X"FC",
		X"C5",X"FD",X"90",X"04",X"A0",X"FF",X"BB",X"FF",X"BD",X"00",X"06",X"FB",X"63",X"02",X"01",X"FE",
		X"A8",X"FC",X"10",X"03",X"4C",X"02",X"96",X"FC",X"B3",X"FC",X"99",X"FE",X"C5",X"04",X"C7",X"FE",
		X"60",X"00",X"F5",X"03",X"E3",X"02",X"8A",X"01",X"C1",X"FA",X"E2",X"01",X"87",X"FE",X"3F",X"01",
		X"A6",X"FE",X"7F",X"01",X"8E",X"FD",X"62",X"FD",X"9E",X"02",X"53",X"FB",X"0F",X"00",X"DD",X"00",
		X"5D",X"FB",X"68",X"01",X"2D",X"03",X"BF",X"03",X"48",X"00",X"DC",X"FE",X"E6",X"04",X"04",X"FE",
		X"39",X"01",X"C1",X"03",X"C4",X"02",X"8A",X"03",X"AF",X"02",X"E3",X"03",X"BE",X"00",X"65",X"FE",
		X"76",X"04",X"49",X"FF",X"1C",X"FC",X"1A",X"01",X"D5",X"03",X"45",X"FD",X"FE",X"02",X"97",X"FF",
		X"19",X"FC",X"00",X"FD",X"5E",X"01",X"8C",X"FE",X"D2",X"01",X"F5",X"03",X"4D",X"02",X"32",X"04",
		X"F3",X"FF",X"F7",X"FE",X"62",X"04",X"AC",X"FE",X"6B",X"FC",X"D1",X"FC",X"F7",X"FC",X"FF",X"01",
		X"2B",X"FD",X"58",X"FC",X"6C",X"01",X"A2",X"FE",X"0B",X"FC",X"AC",X"03",X"59",X"01",X"8E",X"FE",
		X"A4",X"01",X"D2",X"FB",X"8E",X"FD",X"C8",X"FB",X"61",X"01",X"12",X"FF",X"11",X"FC",X"5E",X"02",
		X"AA",X"FD",X"29",X"03",X"F2",X"01",X"3C",X"FC",X"29",X"02",X"08",X"03",X"7A",X"FD",X"56",X"03",
		X"98",X"02",X"16",X"04",X"D1",X"FF",X"AB",X"FF",X"58",X"00",X"25",X"FF",X"EB",X"04",X"A2",X"01",
		X"8A",X"04",X"28",X"01",X"0F",X"FF",X"D6",X"00",X"45",X"FD",X"19",X"FC",X"28",X"03",X"BD",X"01",
		X"69",X"FE",X"7C",X"02",X"02",X"04",X"1F",X"00",X"AC",X"FC",X"7F",X"FC",X"44",X"FD",X"09",X"FC",
		X"5B",X"02",X"6E",X"02",X"82",X"FE",X"F1",X"00",X"EB",X"FE",X"E5",X"00",X"88",X"FE",X"C8",X"03",
		X"F0",X"02",X"22",X"02",X"85",X"FD",X"0E",X"04",X"1E",X"02",X"4D",X"04",X"9A",X"FE",X"8C",X"00",
		X"60",X"FF",X"B4",X"FB",X"C5",X"02",X"B8",X"02",X"94",X"03",X"8B",X"01",X"75",X"FC",X"07",X"FD",
		X"4B",X"FC",X"E4",X"FF",X"D2",X"03",X"81",X"02",X"8F",X"03",X"74",X"02",X"ED",X"03",X"F9",X"FE",
		X"DD",X"FF",X"36",X"04",X"49",X"FD",X"47",X"FD",X"5D",X"01",X"45",X"FE",X"90",X"01",X"30",X"FC",
		X"BC",X"FE",X"35",X"04",X"FD",X"FE",X"CC",X"FF",X"37",X"04",X"A1",X"00",X"68",X"FC",X"F8",X"FC",
		X"98",X"FC",X"F8",X"FC",X"90",X"FC",X"21",X"FD",X"5B",X"01",X"87",X"FE",X"4A",X"01",X"38",X"FD",
		X"2B",X"FC",X"34",X"FF",X"83",X"03",X"C0",X"02",X"7F",X"03",X"84",X"FE",X"C5",X"FD",X"66",X"04",
		X"C3",X"01",X"94",X"04",X"AD",X"FD",X"97",X"01",X"0F",X"FE",X"BC",X"01",X"14",X"FD",X"DC",X"FD",
		X"C2",X"01",X"1F",X"FC",X"E5",X"FE",X"1C",X"04",X"55",X"FF",X"3A",X"FC",X"F8",X"00",X"4F",X"FF",
		X"03",X"FB",X"21",X"01",X"46",X"FF",X"B4",X"FC",X"74",X"FC",X"2C",X"02",X"7F",X"02",X"5A",X"FE",
		X"1D",X"01",X"AF",X"FE",X"30",X"01",X"17",X"FE",X"9F",X"04",X"F5",X"FE",X"C2",X"FC",X"99",X"FC",
		X"9C",X"01",X"35",X"FE",X"49",X"FC",X"41",X"FD",X"92",X"FC",X"16",X"FD",X"4D",X"01",X"DF",X"FE",
		X"04",X"01",X"A8",X"FE",X"94",X"02",X"BD",X"03",X"99",X"00",X"13",X"FC",X"24",X"00",X"10",X"04",
		X"4B",X"FE",X"9B",X"FC",X"39",X"FD",X"52",X"02",X"B3",X"03",X"B4",X"FE",X"BB",X"00",X"31",X"FF",
		X"BB",X"FB",X"21",X"04",X"B7",X"00",X"65",X"FF",X"77",X"00",X"56",X"FF",X"B5",X"00",X"BC",X"FE",
		X"0A",X"05",X"59",X"FD",X"12",X"02",X"B3",X"02",X"0B",X"FE",X"6B",X"02",X"7A",X"03",X"8A",X"02",
		X"A4",X"03",X"F4",X"01",X"A7",X"FE",X"E5",X"00",X"CF",X"FE",X"35",X"01",X"74",X"FC",X"B5",X"FC",
		X"F5",X"FF",X"CA",X"03",X"8A",X"02",X"50",X"03",X"8A",X"FD",X"AF",X"FC",X"12",X"FD",X"7F",X"FC",
		X"97",X"FE",X"57",X"03",X"BE",X"FD",X"E6",X"01",X"9E",X"FD",X"D9",X"03",X"84",X"00",X"9D",X"FE",
		X"39",X"04",X"4B",X"FF",X"33",X"FC",X"4E",X"01",X"72",X"03",X"9B",X"02",X"3E",X"FD",X"B0",X"FD",
		X"F0",X"01",X"67",X"FD",X"C4",X"04",X"3D",X"FF",X"1D",X"FD",X"FC",X"FC",X"8E",X"04",X"84",X"FF",
		X"24",X"00",X"A5",X"FF",X"1F",X"00",X"9A",X"FF",X"38",X"00",X"5F",X"FF",X"D9",X"FB",X"66",X"03",
		X"61",X"02",X"91",X"03",X"7B",X"02",X"65",X"03",X"CC",X"02",X"85",X"00",X"21",X"FB",X"AE",X"FF",
		X"50",X"00",X"CE",X"FE",X"EF",X"03",X"6B",X"FF",X"3C",X"FC",X"4E",X"FD",X"E9",X"00",X"0F",X"FF",
		X"05",X"01",X"B8",X"04",X"FB",X"FF",X"BE",X"FF",X"07",X"00",X"50",X"FF",X"57",X"03",X"14",X"03",
		X"78",X"02",X"EB",X"03",X"A9",X"FF",X"6C",X"FF",X"4E",X"03",X"28",X"03",X"6A",X"FE",X"A5",X"FC",
		X"BE",X"FC",X"4D",X"FD",X"14",X"FC",X"0D",X"FF",X"99",X"00",X"C7",X"FE",X"51",X"03",X"44",X"03",
		X"F4",X"FE",X"3A",X"00",X"0B",X"04",X"5C",X"00",X"E5",X"FB",X"87",X"00",X"19",X"03",X"23",X"03",
		X"E1",X"FD",X"F9",X"FC",X"4C",X"02",X"AC",X"02",X"A2",X"FB",X"B9",X"FF",X"46",X"00",X"F9",X"FC",
		X"1B",X"FC",X"4A",X"01",X"A5",X"FE",X"EE",X"FC",X"21",X"FC",X"9D",X"00",X"51",X"FF",X"5D",X"00",
		X"59",X"FF",X"1A",X"FC",X"77",X"FD",X"A8",X"02",X"C7",X"01",X"5C",X"FE",X"63",X"01",X"09",X"FE",
		X"55",X"04",X"DC",X"01",X"1A",X"04",X"DD",X"FD",X"70",X"01",X"41",X"FE",X"1A",X"02",X"4D",X"00",
		X"55",X"FB",X"47",X"02",X"A9",X"FD",X"79",X"FD",X"76",X"01",X"B6",X"FD",X"F2",X"FB",X"A3",X"FF",
		X"71",X"00",X"D8",X"FE",X"45",X"04",X"B5",X"FE",X"A1",X"FC",X"24",X"FD",X"09",X"FD",X"1C",X"02",
		X"89",X"FD",X"B6",X"03",X"F7",X"FD",X"31",X"FD",X"63",X"FC",X"61",X"FE",X"06",X"01",X"FF",X"FE",
		X"EF",X"00",X"D0",X"FE",X"93",X"01",X"F6",X"FA",X"25",X"02",X"57",X"FE",X"7B",X"01",X"29",X"03",
		X"55",X"FD",X"C3",X"FC",X"32",X"FE",X"64",X"03",X"97",X"02",X"3E",X"FE",X"CC",X"01",X"F8",X"FC",
		X"52",X"FE",X"4C",X"03",X"25",X"03",X"32",X"00",X"01",X"FF",X"C1",X"04",X"98",X"FD",X"72",X"FD",
		X"9D",X"FC",X"2C",X"03",X"50",X"02",X"E3",X"03",X"AC",X"00",X"15",X"FD",X"DC",X"FC",X"59",X"03",
		X"44",X"01",X"9E",X"FE",X"DC",X"02",X"94",X"03",X"A3",X"FF",X"97",X"FF",X"E9",X"03",X"4C",X"02",
		X"71",X"03",X"42",X"02",X"D4",X"FD",X"56",X"FC",X"7F",X"FE",X"F7",X"02",X"ED",X"02",X"EB",X"02",
		X"76",X"02",X"B2",X"FC",X"71",X"FD",X"49",X"FC",X"85",X"FF",X"33",X"03",X"E6",X"02",X"C2",X"02",
		X"33",X"03",X"0D",X"FE",X"A6",X"01",X"75",X"03",X"B1",X"01",X"F6",X"FD",X"3B",X"02",X"F7",X"FA",
		X"3A",X"01",X"DF",X"FE",X"75",X"FE",X"A9",X"00",X"42",X"FF",X"4B",X"00",X"7C",X"FF",X"2C",X"00",
		X"6D",X"FF",X"27",X"04",X"0F",X"02",X"67",X"FE",X"F4",X"01",X"4A",X"02",X"B4",X"FD",X"2F",X"02",
		X"52",X"FB",X"59",X"00",X"D1",X"02",X"FD",X"02",X"E4",X"02",X"70",X"01",X"A2",X"FB",X"70",X"00",
		X"04",X"00",X"C5",X"FB",X"C9",X"01",X"1C",X"FE",X"13",X"FD",X"CA",X"01",X"47",X"FD",X"BF",X"FC",
		X"69",X"FD",X"4D",X"FC",X"EE",X"FF",X"07",X"03",X"3F",X"03",X"90",X"FE",X"E2",X"FC",X"A0",X"FC",
		X"DA",X"FF",X"42",X"03",X"00",X"03",X"A1",X"FE",X"9E",X"FC",X"52",X"FD",X"A3",X"02",X"F5",X"01",
		X"FD",X"FC",X"DD",X"FC",X"7A",X"FD",X"2E",X"FC",X"E5",X"00",X"74",X"FF",X"A4",X"FC",X"F6",X"FC",
		X"A0",X"02",X"C4",X"FF",X"E4",X"FF",X"44",X"00",X"A5",X"FB",X"9E",X"02",X"64",X"02",X"A8",X"FD",
		X"BB",X"FC",X"2A",X"FE",X"00",X"04",X"C4",X"FF",X"DF",X"FF",X"3A",X"00",X"75",X"FF",X"56",X"04",
		X"E0",X"01",X"B9",X"03",X"30",X"02",X"76",X"03",X"7B",X"02",X"45",X"FF",X"EF",X"FB",X"0F",X"03",
		X"23",X"02",X"BF",X"03",X"CA",X"01",X"4E",X"04",X"40",X"FF",X"25",X"00",X"E5",X"FF",X"8C",X"FC",
		X"05",X"FD",X"74",X"01",X"55",X"FE",X"08",X"02",X"7A",X"02",X"76",X"FC",X"52",X"01",X"41",X"03",
		X"3F",X"FD",X"DA",X"FD",X"A0",X"01",X"04",X"FD",X"D4",X"FC",X"00",X"FF",X"D7",X"03",X"78",X"FF",
		X"52",X"FC",X"52",X"01",X"1C",X"03",X"03",X"FE",X"A2",X"01",X"6F",X"FD",X"E3",X"FC",X"44",X"FD",
		X"F1",X"FC",X"68",X"02",X"55",X"02",X"18",X"FD",X"1B",X"FD",X"23",X"FD",X"06",X"FD",X"48",X"FD",
		X"BE",X"FC",X"B4",X"00",X"A4",X"03",X"07",X"FE",X"A4",X"01",X"3E",X"FE",X"AF",X"02",X"02",X"02",
		X"30",X"FC",X"8F",X"FF",X"2A",X"03",X"E2",X"02",X"23",X"02",X"71",X"FC",X"14",X"FF",X"48",X"03",
		X"9E",X"02",X"14",X"03",X"9B",X"02",X"2E",X"03",X"27",X"FE",X"8A",X"01",X"B1",X"FD",X"A6",X"FD",
		X"4C",X"02",X"C7",X"FB",X"F4",X"FF",X"9B",X"02",X"86",X"03",X"17",X"01",X"E3",X"FE",X"2D",X"01",
		X"AE",X"FC",X"EB",X"FC",X"51",X"00",X"19",X"00",X"C6",X"FB",X"6B",X"02",X"B8",X"FD",X"BE",X"02",
		X"C6",X"01",X"06",X"FE",X"A8",X"03",X"7D",X"00",X"A1",X"FC",X"79",X"FD",X"AD",X"FC",X"BA",X"FE",
		X"CE",X"01",X"87",X"FB",X"14",X"01",X"68",X"FF",X"2D",X"00",X"CF",X"03",X"DB",X"FD",X"27",X"FD",
		X"DE",X"02",X"9D",X"01",X"8B",X"FE",X"84",X"01",X"FC",X"FD",X"B4",X"04",X"B0",X"FE",X"87",X"FD",
		X"58",X"FC",X"9D",X"FF",X"06",X"01",X"05",X"FC",X"C2",X"00",X"38",X"03",X"B7",X"02",X"A3",X"FE",
		X"13",X"01",X"E9",X"FE",X"44",X"01",X"80",X"FD",X"A3",X"FC",X"5A",X"FF",X"A2",X"03",X"C7",X"FF",
		X"38",X"FC",X"9C",X"01",X"EF",X"02",X"FB",X"02",X"85",X"02",X"7B",X"03",X"A6",X"FE",X"F0",X"00",
		X"08",X"FF",X"06",X"01",X"26",X"FE",X"57",X"FD",X"C6",X"02",X"38",X"FB",X"F7",X"00",X"6C",X"FF",
		X"24",X"00",X"26",X"03",X"0A",X"03",X"2B",X"FE",X"CB",X"01",X"51",X"FD",X"7E",X"00",X"D5",X"FF",
		X"34",X"FC",X"CC",X"FD",X"EA",X"FC",X"10",X"03",X"C2",X"01",X"F8",X"FC",X"90",X"FE",X"0E",X"04",
		X"66",X"FF",X"DF",X"FF",X"9E",X"03",X"67",X"02",X"ED",X"FE",X"33",X"FC",X"6C",X"FE",X"E9",X"01",
		X"C5",X"03",X"F5",X"FD",X"9F",X"FD",X"28",X"01",X"24",X"FF",X"BB",X"00",X"3C",X"FF",X"FE",X"00",
		X"0F",X"FD",X"B4",X"FC",X"B7",X"00",X"D3",X"FF",X"58",X"FC",X"C7",X"FD",X"B9",X"FC",X"20",X"FE",
		X"CB",X"01",X"2A",X"FD",X"47",X"FD",X"8D",X"01",X"7C",X"FE",X"72",X"FC",X"9F",X"FE",X"DB",X"02",
		X"AC",X"01",X"D3",X"FB",X"BB",X"00",X"AA",X"02",X"7A",X"03",X"64",X"FE",X"5D",X"FD",X"71",X"01",
		X"FB",X"FE",X"12",X"01",X"D1",X"FE",X"CF",X"02",X"01",X"03",X"B2",X"FD",X"26",X"03",X"3B",X"01",
		X"FB",X"FE",X"5B",X"01",X"B6",X"FC",X"47",X"FD",X"F7",X"FF",X"04",X"04",X"24",X"FE",X"94",X"01",
		X"56",X"FE",X"2C",X"FD",X"5B",X"03",X"6E",X"01",X"D6",X"FC",X"37",X"FF",X"58",X"03",X"3D",X"FD",
		X"F0",X"03",X"5B",X"00",X"8D",X"FF",X"ED",X"00",X"9B",X"FC",X"90",X"FD",X"21",X"FD",X"57",X"FD",
		X"46",X"FD",X"70",X"FD",X"B3",X"02",X"1F",X"02",X"E4",X"FC",X"CC",X"FE",X"D1",X"03",X"EC",X"FF",
		X"86",X"FD",X"7D",X"02",X"1C",X"FC",X"19",X"00",X"5F",X"00",X"85",X"FF",X"11",X"01",X"78",X"FB",
		X"9D",X"02",X"D7",X"FD",X"EC",X"FD",X"7E",X"01",X"A8",X"FE",X"AB",X"02",X"1C",X"03",X"81",X"02",
		X"48",X"03",X"3D",X"02",X"C0",X"03",X"84",X"00",X"80",X"FF",X"C4",X"00",X"FB",X"FE",X"1F",X"04",
		X"D8",X"01",X"B4",X"03",X"A3",X"FD",X"DD",X"FD",X"A9",X"01",X"A0",X"FD",X"DC",X"FD",X"33",X"04",
		X"9D",X"FF",X"DB",X"FF",X"1C",X"03",X"04",X"03",X"D8",X"FE",X"F6",X"FC",X"52",X"FD",X"79",X"FD",
		X"C6",X"FC",X"41",X"01",X"35",X"FF",X"C2",X"FC",X"2C",X"02",X"19",X"FE",X"C9",X"02",X"C5",X"02",
		X"C7",X"02",X"0A",X"03",X"86",X"00",X"2A",X"FC",X"3C",X"01",X"F6",X"02",X"C8",X"02",X"05",X"FE",
		X"2C",X"FD",X"1F",X"FD",X"B9",X"00",X"88",X"03",X"1F",X"02",X"CE",X"FE",X"48",X"01",X"F9",X"FD",
		X"9E",X"FC",X"2C",X"FF",X"6D",X"03",X"16",X"00",X"2D",X"FF",X"9D",X"04",X"7E",X"FD",X"48",X"02",
		X"AC",X"FD",X"41",X"03",X"D1",X"FE",X"0A",X"01",X"15",X"FF",X"E6",X"FC",X"44",X"FD",X"1D",X"FE",
		X"A5",X"01",X"3D",X"FE",X"A0",X"03",X"8D",X"00",X"7B",X"FC",X"84",X"00",X"68",X"03",X"D4",X"FE",
		X"CD",X"FC",X"81",X"02",X"36",X"02",X"98",X"FD",X"20",X"FD",X"8B",X"FD",X"58",X"01",X"BF",X"03",
		X"41",X"01",X"2B",X"FF",X"F6",X"00",X"DB",X"FE",X"3A",X"03",X"CE",X"02",X"1A",X"00",X"36",X"FC",
		X"DD",X"01",X"90",X"FE",X"FF",X"FC",X"6B",X"FD",X"EC",X"FD",X"29",X"03",X"6C",X"02",X"1B",X"03",
		X"3F",X"02",X"AB",X"FD",X"FD",X"FD",X"66",X"02",X"B7",X"FB",X"CA",X"00",X"CD",X"FF",X"D0",X"FF",
		X"D0",X"03",X"67",X"FE",X"34",X"01",X"1A",X"FF",X"EB",X"00",X"2B",X"FF",X"0D",X"01",X"AC",X"FE",
		X"6C",X"03",X"0C",X"02",X"F7",X"FD",X"C3",X"FC",X"04",X"FF",X"96",X"01",X"2A",X"FC",X"69",X"00",
		X"0B",X"03",X"9B",X"02",X"EE",X"02",X"5C",X"FE",X"52",X"FD",X"12",X"02",X"F2",X"FD",X"50",X"03",
		X"23",X"02",X"71",X"03",X"9A",X"01",X"0D",X"FF",X"EC",X"00",X"F4",X"FE",X"9C",X"02",X"6A",X"03",
		X"71",X"FF",X"4D",X"00",X"DC",X"FF",X"16",X"00",X"01",X"04",X"A8",X"01",X"BD",X"03",X"0A",X"01",
		X"FF",X"FD",X"54",X"FC",X"20",X"00",X"7C",X"00",X"97",X"FC",X"67",X"FE",X"26",X"03",X"F6",X"00",
		X"9D",X"FC",X"E4",X"FF",X"B9",X"03",X"98",X"FE",X"F8",X"00",X"2A",X"03",X"C2",X"FD",X"25",X"FD",
		X"27",X"FE",X"DF",X"02",X"C1",X"02",X"07",X"01",X"53",X"FC",X"3A",X"FE",X"43",X"FC",X"AF",X"FF",
		X"97",X"00",X"04",X"FF",X"BD",X"03",X"71",X"FF",X"A4",X"FC",X"8F",X"01",X"E8",X"02",X"63",X"02",
		X"0B",X"FE",X"51",X"02",X"26",X"FC",X"2D",X"00",X"02",X"00",X"FC",X"FF",X"1F",X"00",X"C6",X"FF",
		X"B9",X"03",X"38",X"02",X"4D",X"01",X"C5",X"FB",X"69",X"01",X"54",X"FF",X"B4",X"FC",X"F2",X"01",
		X"0A",X"FE",X"45",X"FD",X"42",X"FD",X"B2",X"FD",X"AC",X"FC",X"14",X"00",X"57",X"00",X"67",X"FF",
		X"DD",X"03",X"E9",X"01",X"42",X"03",X"BB",X"FD",X"42",X"FD",X"0D",X"00",X"D4",X"03",X"22",X"FE",
		X"79",X"FD",X"62",X"FD",X"D2",X"02",X"BC",X"01",X"28",X"FD",X"B8",X"FE",X"D8",X"03",X"7B",X"FF",
		X"D7",X"FF",X"C3",X"03",X"53",X"FE",X"5C",X"01",X"9F",X"FE",X"C3",X"FC",X"F8",X"FD",X"B4",X"FC",
		X"CF",X"01",X"7F",X"FE",X"F4",X"01",X"5B",X"02",X"E4",X"FD",X"8D",X"03",X"7E",X"00",X"E5",X"FE",
		X"FE",X"03",X"ED",X"FE",X"82",X"00",X"46",X"03",X"5E",X"02",X"9D",X"02",X"0E",X"FE",X"1D",X"02",
		X"B0",X"FC",X"C9",X"01",X"86",X"FE",X"BF",X"01",X"1B",X"03",X"B0",X"01",X"1D",X"FD",X"B7",X"FD",
		X"D9",X"FC",X"03",X"00",X"2A",X"03",X"68",X"02",X"C8",X"02",X"9E",X"02",X"5C",X"02",X"4C",X"FE",
		X"AB",X"01",X"08",X"FE",X"85",X"03",X"B6",X"FD",X"37",X"02",X"03",X"FD",X"FD",X"FE",X"E1",X"00",
		X"EA",X"FE",X"EE",X"02",X"F5",X"02",X"61",X"FF",X"47",X"00",X"D3",X"FF",X"43",X"FC",X"C5",X"02",
		X"17",X"02",X"4A",X"03",X"17",X"01",X"58",X"FD",X"63",X"FD",X"24",X"02",X"4F",X"02",X"E6",X"FC",
		X"0B",X"FF",X"48",X"01",X"B3",X"FC",X"A6",X"FD",X"AB",X"FF",X"05",X"04",X"D7",X"FD",X"E9",X"01",
		X"3F",X"02",X"1D",X"FE",X"9B",X"FC",X"57",X"FF",X"B8",X"00",X"22",X"FF",X"42",X"01",X"05",X"FC",
		X"93",X"FE",X"17",X"FC",X"48",X"00",X"24",X"00",X"74",X"FF",X"9D",X"03",X"04",X"FF",X"E5",X"FC",
		X"E4",X"01",X"BF",X"02",X"39",X"02",X"BC",X"FD",X"C6",X"03",X"E9",X"FF",X"F3",X"FF",X"33",X"00",
		X"93",X"FF",X"73",X"03",X"39",X"02",X"AD",X"02",X"F0",X"02",X"DB",X"FF",X"86",X"FF",X"C7",X"03",
		X"3D",X"FE",X"55",X"FD",X"0F",X"02",X"12",X"02",X"3E",X"FE",X"D7",X"01",X"7D",X"FC",X"8D",X"FF",
		X"4C",X"03",X"6E",X"FF",X"D7",X"FF",X"DE",X"03",X"19",X"00",X"07",X"FF",X"BD",X"03",X"CF",X"FE",
		X"A1",X"00",X"68",X"FF",X"95",X"FC",X"F6",X"FD",X"F9",X"FC",X"D0",X"FD",X"F7",X"FC",X"EE",X"FE",
		X"7A",X"03",X"A3",X"FF",X"BB",X"FF",X"66",X"03",X"2E",X"02",X"D3",X"FE",X"5B",X"FE",X"76",X"04",
		X"1F",X"FE",X"60",X"01",X"A9",X"FE",X"67",X"01",X"7B",X"02",X"38",X"FE",X"B1",X"01",X"25",X"FD",
		X"9A",X"FD",X"5A",X"FD",X"4F",X"FD",X"E7",X"FF",X"B7",X"03",X"2C",X"FE",X"88",X"01",X"A9",X"02",
		X"D9",X"02",X"A7",X"FF",X"D0",X"FC",X"D7",X"FD",X"26",X"FD",X"57",X"02",X"F8",X"01",X"9A",X"FD",
		X"2A",X"FD",X"F4",X"FE",X"31",X"03",X"10",X"02",X"34",X"03",X"0C",X"FF",X"28",X"FD",X"83",X"FD",
		X"AE",X"FD",X"CF",X"01",X"92",X"FD",X"81",X"FD",X"60",X"FD",X"8E",X"01",X"6A",X"FE",X"FC",X"FC",
		X"F3",X"FD",X"DA",X"FC",X"65",X"FF",X"C0",X"02",X"D7",X"02",X"E3",X"FF",X"A7",X"FC",X"77",X"01",
		X"C9",X"02",X"13",X"FE",X"46",X"FD",X"28",X"FE",X"0D",X"03",X"8C",X"FE",X"60",X"FD",X"59",X"FD",
		X"4D",X"FE",X"93",X"01",X"4F",X"FE",X"67",X"03",X"E5",X"01",X"73",X"03",X"4B",X"FF",X"67",X"FD",
		X"4D",X"FD",X"C7",X"01",X"61",X"02",X"7A",X"FE",X"84",X"01",X"60",X"FE",X"29",X"03",X"14",X"02",
		X"69",X"FE",X"FF",X"FC",X"FD",X"FD",X"F0",X"FC",X"47",X"FF",X"35",X"03",X"25",X"00",X"DF",X"FC",
		X"FF",X"FD",X"25",X"FD",X"E0",X"FD",X"79",X"FD",X"31",X"02",X"C1",X"FD",X"C4",X"03",X"10",X"00",
		X"AD",X"FF",X"68",X"02",X"63",X"FE",X"63",X"02",X"F6",X"02",X"FC",X"00",X"D0",X"FC",X"15",X"00",
		X"28",X"03",X"4B",X"02",X"79",X"FF",X"71",X"FC",X"DA",X"FE",X"AB",X"00",X"95",X"FF",X"94",X"00",
		X"52",X"FF",X"8F",X"02",X"0A",X"03",X"62",X"01",X"EF",X"FE",X"28",X"02",X"76",X"03",X"9C",X"FF",
		X"40",X"00",X"F6",X"FF",X"F1",X"FF",X"A5",X"03",X"E3",X"FD",X"AE",X"FD",X"4C",X"FD",X"56",X"FE",
		X"DA",X"02",X"36",X"02",X"20",X"03",X"11",X"00",X"1D",X"FD",X"C2",X"FD",X"4E",X"FD",X"EA",X"FE",
		X"B5",X"03",X"52",X"FF",X"2E",X"00",X"27",X"03",X"43",X"02",X"9C",X"02",X"5F",X"FE",X"A4",X"01",
		X"B9",X"FD",X"52",X"FD",X"DE",X"FE",X"74",X"03",X"EB",X"FF",X"2D",X"FD",X"C4",X"FD",X"61",X"FD",
		X"CB",X"FD",X"25",X"FD",X"0A",X"00",X"2D",X"03",X"20",X"02",X"FC",X"02",X"2F",X"FE",X"C1",X"FD",
		X"40",X"02",X"AE",X"02",X"69",X"02",X"AE",X"02",X"60",X"02",X"B4",X"02",X"51",X"02",X"C5",X"02",
		X"2C",X"02",X"0F",X"03",X"48",X"00",X"18",X"FD",X"C8",X"FD",X"3D",X"FD",X"41",X"01",X"1A",X"FF",
		X"10",X"01",X"A4",X"03",X"9B",X"00",X"72",X"FF",X"D2",X"00",X"7B",X"FD",X"02",X"FD",X"D0",X"00",
		X"83",X"FF",X"78",X"00",X"87",X"FF",X"A1",X"FC",X"41",X"03",X"1D",X"FF",X"81",X"FD",X"69",X"FD",
		X"97",X"01",X"A6",X"FE",X"81",X"01",X"3F",X"FE",X"4B",X"03",X"55",X"00",X"43",X"FF",X"10",X"03",
		X"68",X"02",X"B5",X"FF",X"A8",X"FC",X"F1",X"01",X"66",X"FE",X"B2",X"01",X"A4",X"FD",X"A7",X"FD",
		X"75",X"FD",X"B8",X"FD",X"67",X"FD",X"21",X"FE",X"B9",X"02",X"41",X"01",X"5A",X"FE",X"FF",X"03",
		X"0C",X"FF",X"93",X"00",X"DE",X"FF",X"C2",X"FC",X"E8",X"01",X"A2",X"02",X"10",X"02",X"A5",X"FD",
		X"7D",X"FD",X"23",X"01",X"0C",X"03",X"16",X"02",X"DB",X"02",X"32",X"02",X"02",X"02",X"19",X"FC",
		X"D7",X"00",X"80",X"FF",X"76",X"00",X"9F",X"FF",X"79",X"00",X"7E",X"FF",X"F0",X"00",X"11",X"03",
		X"8E",X"FC",X"90",X"FF",X"E5",X"00",X"49",X"FD",X"F5",X"FD",X"36",X"02",X"B9",X"02",X"3E",X"01",
		X"50",X"FE",X"FE",X"03",X"FD",X"FE",X"70",X"00",X"B7",X"02",X"8D",X"02",X"81",X"FE",X"A1",X"01",
		X"C7",X"02",X"C9",X"01",X"F9",X"FC",X"7A",X"FF",X"09",X"01",X"B6",X"FC",X"AA",X"FE",X"8B",X"01",
		X"0B",X"FD",X"7D",X"FF",X"27",X"01",X"5A",X"FC",X"F3",X"00",X"8B",X"02",X"85",X"02",X"5D",X"02",
		X"5A",X"02",X"FB",X"FD",X"F1",X"02",X"C4",X"00",X"19",X"FF",X"46",X"01",X"72",X"FC",X"F9",X"FE",
		X"20",X"01",X"B1",X"FD",X"68",X"FD",X"E3",X"FD",X"17",X"FD",X"87",X"00",X"DB",X"02",X"45",X"02",
		X"78",X"02",X"36",X"FE",X"34",X"FD",X"AE",X"FE",X"84",X"01",X"26",X"FD",X"C4",X"FD",X"48",X"FF",
		X"D4",X"03",X"88",X"FE",X"09",X"FE",X"BD",X"FC",X"78",X"00",X"EE",X"FF",X"DC",X"FF",X"3B",X"03",
		X"0A",X"02",X"95",X"02",X"63",X"FE",X"86",X"01",X"60",X"FE",X"E4",X"02",X"FF",X"00",X"CE",X"FC",
		X"31",X"00",X"A4",X"02",X"A6",X"02",X"D0",X"FE",X"A4",X"FE",X"83",X"03",X"BA",X"FF",X"FF",X"FC",
		X"19",X"01",X"44",X"FF",X"CF",X"00",X"19",X"03",X"03",X"FD",X"F4",X"FE",X"19",X"02",X"DA",X"02",
		X"DF",X"01",X"40",X"03",X"15",X"FF",X"81",X"00",X"C8",X"FF",X"56",X"FC",X"7B",X"00",X"2D",X"00",
		X"19",X"FD",X"C3",X"FD",X"EF",X"00",X"46",X"FF",X"98",X"FC",X"0F",X"FF",X"D8",X"00",X"FB",X"FE",
		X"8D",X"02",X"7C",X"02",X"46",X"02",X"9F",X"02",X"1E",X"02",X"CD",X"02",X"53",X"FE",X"BD",X"01",
		X"6D",X"02",X"A8",X"02",X"34",X"FF",X"22",X"FD",X"AD",X"01",X"6C",X"02",X"6F",X"FD",X"B4",X"FE",
		X"6B",X"01",X"FA",X"FC",X"76",X"FF",X"51",X"03",X"18",X"FF",X"79",X"00",X"B4",X"FF",X"A2",X"FC",
		X"96",X"FE",X"54",X"01",X"61",X"03",X"71",X"FE",X"33",X"01",X"90",X"02",X"63",X"02",X"45",X"02",
		X"80",X"02",X"49",X"02",X"6B",X"01",X"30",X"FC",X"02",X"01",X"33",X"FF",X"8C",X"00",X"6A",X"FF",
		X"FD",X"FC",X"1B",X"FE",X"E1",X"01",X"7A",X"02",X"61",X"02",X"3C",X"02",X"7B",X"02",X"C4",X"FD",
		X"F4",X"FD",X"E6",X"FC",X"8C",X"FF",X"56",X"00",X"87",X"FF",X"73",X"00",X"31",X"FF",X"B7",X"03",
		X"1A",X"FE",X"68",X"01",X"76",X"02",X"7A",X"FD",X"B2",X"FE",X"12",X"01",X"95",X"FE",X"E9",X"02",
		X"A6",X"FD",X"2F",X"FE",X"5C",X"02",X"22",X"02",X"D2",X"02",X"38",X"00",X"6A",X"FD",X"59",X"FD",
		X"D8",X"00",X"3F",X"FF",X"A3",X"00",X"F4",X"FE",X"EE",X"FC",X"2B",X"FE",X"36",X"FD",X"09",X"FE",
		X"4A",X"FD",X"36",X"FE",X"FE",X"01",X"7B",X"02",X"7B",X"02",X"DF",X"00",X"88",X"FE",X"F9",X"03",
		X"7A",X"FE",X"EC",X"00",X"65",X"02",X"8F",X"02",X"C2",X"01",X"A8",X"FE",X"CE",X"01",X"CD",X"02",
		X"BB",X"01",X"2F",X"03",X"8A",X"FF",X"D4",X"FD",X"E8",X"FC",X"A7",X"FF",X"23",X"00",X"C2",X"FF",
		X"0B",X"00",X"DE",X"FF",X"F0",X"FF",X"FC",X"FF",X"B9",X"FF",X"5F",X"FC",X"20",X"FF",X"BE",X"00",
		X"C1",X"FE",X"E3",X"02",X"22",X"00",X"69",X"FF",X"D6",X"00",X"2C",X"FC",X"B6",X"FF",X"F3",X"01",
		X"B1",X"02",X"1C",X"02",X"3B",X"00",X"5F",X"FC",X"E4",X"01",X"D9",X"01",X"FA",X"02",X"2B",X"01",
		X"67",X"FE",X"B1",X"FC",X"ED",X"FF",X"4C",X"00",X"98",X"FD",X"36",X"FD",X"FA",X"00",X"1E",X"FF",
		X"71",X"FE",X"89",X"03",X"43",X"FF",X"F5",X"FF",X"29",X"03",X"6D",X"FE",X"BD",X"FD",X"86",X"01",
		X"DE",X"02",X"13",X"01",X"B1",X"FE",X"90",X"02",X"28",X"02",X"61",X"02",X"35",X"02",X"72",X"02",
		X"1C",X"FF",X"00",X"FD",X"3E",X"02",X"DE",X"FF",X"49",X"FD",X"CA",X"FD",X"A7",X"FD",X"A4",X"FD",
		X"E5",X"01",X"C4",X"01",X"4A",X"FE",X"A3",X"02",X"F6",X"00",X"B6",X"FC",X"84",X"00",X"A6",X"FF",
		X"10",X"00",X"D9",X"FF",X"0A",X"00",X"84",X"03",X"79",X"FC",X"7E",X"01",X"A3",X"FE",X"1D",X"01",
		X"B1",X"FE",X"7C",X"01",X"81",X"02",X"B7",X"01",X"DF",X"FC",X"CD",X"FF",X"49",X"00",X"29",X"FF",
		X"48",X"03",X"F3",X"FE",X"56",X"FD",X"62",X"01",X"45",X"02",X"ED",X"FD",X"77",X"FD",X"8E",X"00",
		X"DD",X"02",X"31",X"FE",X"B3",X"01",X"56",X"02",X"4E",X"02",X"21",X"02",X"92",X"02",X"7C",X"00",
		X"EB",X"FC",X"3B",X"00",X"D7",X"02",X"A0",X"FE",X"CA",X"00",X"00",X"FF",X"C3",X"00",X"BD",X"FE",
		X"07",X"02",X"5C",X"02",X"07",X"02",X"79",X"FE",X"3E",X"01",X"AA",X"FD",X"DD",X"FD",X"3F",X"FD",
		X"8F",X"FF",X"6B",X"02",X"79",X"02",X"24",X"FF",X"4C",X"00",X"E4",X"02",X"E2",X"FD",X"13",X"02",
		X"84",X"01",X"77",X"FD",X"E8",X"FD",X"60",X"FD",X"54",X"FE",X"00",X"01",X"3C",X"FE",X"E3",X"FC",
		X"F4",X"FF",X"EF",X"FF",X"D9",X"FF",X"EE",X"FF",X"E5",X"FF",X"E6",X"FF",X"AB",X"FC",X"98",X"FE",
		X"74",X"01",X"21",X"02",X"01",X"FD",X"61",X"FE",X"F7",X"FC",X"21",X"00",X"1C",X"02",X"33",X"FD",
		X"48",X"FF",X"F4",X"00",X"3F",X"FD",X"D2",X"FD",X"EE",X"FF",X"32",X"03",X"72",X"FE",X"D6",X"FD",
		X"4D",X"01",X"B6",X"FE",X"80",X"01",X"3A",X"FD",X"61",X"FF",X"53",X"02",X"A2",X"02",X"93",X"FF",
		X"1E",X"FE",X"AB",X"02",X"0E",X"02",X"44",X"02",X"8B",X"02",X"7E",X"FF",X"F6",X"FF",X"2B",X"03",
		X"07",X"FE",X"C8",X"01",X"3E",X"02",X"40",X"02",X"51",X"02",X"22",X"01",X"BB",X"FC",X"5A",X"00",
		X"0D",X"00",X"EB",X"FC",X"1F",X"FF",X"71",X"02",X"AA",X"00",X"9E",X"FC",X"0A",X"01",X"2B",X"FF",
		X"7D",X"00",X"E8",X"02",X"73",X"01",X"D2",X"FE",X"01",X"01",X"81",X"FE",X"B5",X"02",X"B2",X"01",
		X"E9",X"02",X"57",X"FF",X"A5",X"FD",X"81",X"FD",X"58",X"01",X"28",X"02",X"AB",X"02",X"32",X"FF",
		X"48",X"00",X"8B",X"FF",X"FB",X"FC",X"16",X"02",X"F7",X"01",X"67",X"02",X"1D",X"02",X"39",X"01",
		X"A2",X"FC",X"46",X"00",X"13",X"02",X"7B",X"02",X"C2",X"01",X"B7",X"02",X"70",X"FD",X"5B",X"00",
		X"7A",X"FF",X"F7",X"FF",X"CE",X"02",X"B8",X"01",X"9B",X"FE",X"1C",X"01",X"9B",X"FD",X"DA",X"FE",
		X"02",X"01",X"F8",X"FC",X"BB",X"FF",X"E4",X"02",X"CA",X"FE",X"99",X"00",X"FE",X"FE",X"75",X"FD",
		X"C3",X"01",X"87",X"02",X"EB",X"FE",X"87",X"00",X"F8",X"FE",X"7B",X"FD",X"95",X"01",X"9B",X"FD",
		X"CE",X"FD",X"DF",X"FD",X"48",X"FD",X"31",X"00",X"C2",X"FF",X"E6",X"FF",X"E0",X"FF",X"C1",X"FC",
		X"9F",X"FE",X"3C",X"01",X"AC",X"02",X"EA",X"01",X"3B",X"FF",X"12",X"FD",X"72",X"FE",X"93",X"01",
		X"E3",X"01",X"1B",X"FD",X"62",X"FE",X"15",X"FD",X"0E",X"00",X"9C",X"02",X"5A",X"FF",X"3F",X"FD",
		X"36",X"FE",X"5B",X"FD",X"97",X"FE",X"34",X"01",X"C6",X"FD",X"D3",X"FD",X"E4",X"FD",X"81",X"01",
		X"FF",X"FD",X"EC",X"FD",X"7E",X"FD",X"55",X"FF",X"7E",X"02",X"4C",X"02",X"ED",X"FF",X"08",X"FD",
		X"5E",X"01",X"4D",X"02",X"3D",X"02",X"CC",X"01",X"2E",X"FE",X"F4",X"02",X"30",X"00",X"6E",X"FF",
		X"25",X"02",X"66",X"FE",X"04",X"02",X"97",X"02",X"67",X"00",X"25",X"FF",X"B7",X"02",X"20",X"02",
		X"61",X"FF",X"42",X"00",X"84",X"FF",X"FB",X"FC",X"BC",X"02",X"EB",X"00",X"0E",X"FE",X"69",X"FE",
		X"71",X"03",X"3A",X"FF",X"98",X"FE",X"87",X"01",X"15",X"03",X"C9",X"FF",X"F3",X"FF",X"E9",X"FF",
		X"D7",X"FF",X"1E",X"00",X"CB",X"FC",X"DB",X"01",X"C6",X"01",X"31",X"FE",X"A7",X"FD",X"E5",X"FD",
		X"DC",X"FD",X"96",X"FD",X"C1",X"FF",X"A5",X"02",X"0E",X"02",X"41",X"01",X"3E",X"FE",X"A9",X"03",
		X"D3",X"FE",X"A6",X"00",X"77",X"FF",X"71",X"FD",X"F0",X"FD",X"11",X"FE",X"75",X"01",X"E4",X"FD",
		X"D8",X"FD",X"E7",X"FD",X"A8",X"FD",X"A7",X"FF",X"20",X"03",X"D5",X"FE",X"C7",X"00",X"88",X"02",
		X"26",X"02",X"60",X"00",X"D4",X"FC",X"38",X"01",X"19",X"02",X"6B",X"02",X"9B",X"01",X"BD",X"FE",
		X"C1",X"01",X"83",X"02",X"AF",X"01",X"E7",X"02",X"6F",X"FF",X"19",X"00",X"F6",X"FF",X"05",X"FD",
		X"75",X"FE",X"2D",X"FD",X"34",X"00",X"68",X"02",X"08",X"02",X"37",X"02",X"1A",X"02",X"FD",X"01",
		X"E6",X"FD",X"FA",X"FD",X"9F",X"FD",X"32",X"FE",X"3E",X"FD",X"52",X"00",X"0A",X"00",X"46",X"FD",
		X"2A",X"FE",X"C0",X"FD",X"BF",X"FD",X"D8",X"FF",X"D0",X"02",X"B6",X"01",X"85",X"02",X"D0",X"01",
		X"79",X"02",X"CE",X"01",X"81",X"02",X"AC",X"01",X"CF",X"02",X"E4",X"FF",X"75",X"FF",X"BA",X"02",
		X"B5",X"01",X"7D",X"02",X"73",X"FE",X"C7",X"FD",X"D0",X"FD",X"F6",X"FD",X"A2",X"FD",X"FA",X"00",
		X"6C",X"02",X"EB",X"01",X"51",X"02",X"6B",X"01",X"59",X"FD",X"6C",X"FF",X"D5",X"00",X"D8",X"FC",
		X"9E",X"00",X"22",X"02",X"42",X"02",X"95",X"FE",X"CF",X"FD",X"DE",X"01",X"9F",X"01",X"64",X"FD",
		X"2A",X"01",X"15",X"02",X"67",X"FE",X"67",X"FD",X"FD",X"FE",X"E2",X"00",X"C8",X"FD",X"85",X"FD",
		X"2E",X"00",X"E3",X"FF",X"DD",X"FF",X"0E",X"00",X"B4",X"FC",X"FE",X"FE",X"F3",X"00",X"00",X"03",
		X"40",X"01",X"00",X"03",X"BE",X"FD",X"5C",X"02",X"CE",X"00",X"70",X"FF",X"4A",X"00",X"77",X"FF",
		X"96",X"00",X"59",X"FD",X"31",X"FE",X"93",X"FD",X"F6",X"00",X"2D",X"FF",X"D2",X"00",X"F3",X"02",
		X"D4",X"00",X"46",X"FE",X"75",X"FD",X"60",X"FE",X"85",X"FD",X"B8",X"02",X"7E",X"00",X"86",X"FF",
		X"75",X"00",X"1F",X"FF",X"EA",X"02",X"76",X"FF",X"80",X"FD",X"3A",X"FE",X"8E",X"FD",X"84",X"FE",
		X"15",X"01",X"52",X"FE",X"88",X"FD",X"69",X"FE",X"31",X"FD",X"73",X"00",X"7C",X"01",X"F5",X"FE",
		X"0A",X"01",X"E3",X"FE",X"87",X"01",X"44",X"FC",X"AF",X"01",X"BA",X"FE",X"44",X"01",X"B6",X"FE",
		X"CC",X"01",X"68",X"01",X"15",X"FF",X"D4",X"00",X"37",X"FF",X"07",X"01",X"37",X"FD",X"57",X"FE",
		X"C5",X"FD",X"FC",X"FD",X"28",X"FE",X"6C",X"FD",X"9A",X"00",X"B8",X"FF",X"5F",X"00",X"B5",X"FF",
		X"89",X"00",X"37",X"FF",X"4B",X"FD",X"7C",X"FE",X"9A",X"FD",X"4B",X"FE",X"C8",X"FD",X"22",X"FE",
		X"F7",X"FD",X"F2",X"FD",X"41",X"FE",X"73",X"FD",X"59",X"00",X"0D",X"00",X"1B",X"00",X"1C",X"00",
		X"24",X"00",X"1E",X"03",X"F6",X"FD",X"16",X"02",X"EB",X"FD",X"7E",X"03",X"A2",X"FF",X"54",X"00",
		X"0B",X"00",X"DB",X"FF",X"FE",X"02",X"D8",X"FE",X"D7",X"FD",X"38",X"FE",X"AB",X"FD",X"8B",X"00",
		X"8C",X"02",X"FC",X"01",X"FF",X"FE",X"65",X"01",X"31",X"02",X"88",X"FD",X"99",X"FE",X"50",X"FD",
		X"1E",X"00",X"2B",X"02",X"7D",X"02",X"64",X"FF",X"B4",X"FD",X"64",X"01",X"60",X"02",X"BE",X"FD",
		X"AB",X"00",X"61",X"02",X"22",X"02",X"CF",X"FE",X"8C",X"01",X"4F",X"02",X"2C",X"02",X"4E",X"01",
		X"75",X"FD",X"8F",X"FE",X"4B",X"FD",X"F7",X"00",X"86",X"FF",X"84",X"00",X"C4",X"02",X"12",X"FE",
		X"7E",X"FE",X"3F",X"02",X"59",X"FF",X"92",X"00",X"F0",X"02",X"38",X"01",X"1E",X"FF",X"C4",X"01",
		X"62",X"02",X"FC",X"01",X"FC",X"00",X"C7",X"FC",X"47",X"01",X"51",X"FF",X"E1",X"FD",X"F8",X"FD",
		X"37",X"FE",X"BC",X"FD",X"E3",X"FE",X"19",X"02",X"3E",X"02",X"D6",X"01",X"ED",X"FE",X"41",X"01",
		X"2B",X"FE",X"01",X"FE",X"F6",X"FD",X"6D",X"FF",X"17",X"03",X"4B",X"FF",X"0C",X"FE",X"DF",X"FD",
		X"88",X"01",X"FF",X"01",X"8D",X"FE",X"58",X"02",X"FE",X"00",X"E0",X"FE",X"E1",X"02",X"78",X"01",
		X"D3",X"02",X"B1",X"00",X"5A",X"FF",X"2A",X"01",X"19",X"FD",X"AF",X"00",X"E2",X"FF",X"FD",X"FF",
		X"14",X"03",X"49",X"01",X"F1",X"02",X"D1",X"00",X"7D",X"FF",X"CB",X"00",X"23",X"FE",X"BD",X"FD",
		X"AD",X"FE",X"82",X"01",X"BD",X"02",X"8E",X"00",X"4C",X"FE",X"63",X"FD",X"B5",X"00",X"B4",X"FF",
		X"42",X"00",X"BA",X"02",X"A2",X"01",X"CC",X"FE",X"9D",X"FD",X"DE",X"FE",X"5C",X"02",X"BF",X"00",
		X"DD",X"FE",X"6D",X"03",X"D4",X"FE",X"53",X"FF",X"A4",X"00",X"78",X"FF",X"DC",X"00",X"6E",X"FD",
		X"39",X"FE",X"89",X"00",X"D4",X"FF",X"2A",X"FD",X"D5",X"FE",X"40",X"FD",X"84",X"FF",X"B7",X"00",
		X"21",X"FF",X"C5",X"02",X"09",X"00",X"A7",X"FD",X"6E",X"FE",X"9F",X"FD",X"BC",X"FF",X"04",X"01",
		X"EB",X"FC",X"51",X"01",X"36",X"FF",X"E8",X"00",X"2A",X"FF",X"E5",X"FD",X"31",X"02",X"F4",X"01",
		X"32",X"02",X"07",X"02",X"18",X"02",X"20",X"02",X"F1",X"01",X"60",X"02",X"F3",X"FE",X"FC",X"FE",
		X"0E",X"03",X"70",X"FF",X"28",X"00",X"B1",X"02",X"95",X"01",X"85",X"02",X"62",X"01",X"B2",X"FE",
		X"87",X"FD",X"B7",X"FE",X"38",X"FD",X"53",X"00",X"BB",X"01",X"D6",X"02",X"AE",X"FE",X"59",X"01",
		X"A0",X"FE",X"10",X"02",X"85",X"FF",X"8F",X"00",X"81",X"FF",X"BE",X"00",X"10",X"FF",X"27",X"FE",
		X"4E",X"01",X"12",X"FF",X"F1",X"00",X"3B",X"FF",X"ED",X"00",X"00",X"FF",X"3B",X"03",X"21",X"01",
		X"D1",X"02",X"4C",X"01",X"A7",X"02",X"44",X"FD",X"48",X"01",X"0D",X"FF",X"FC",X"00",X"2C",X"02",
		X"1C",X"02",X"BA",X"01",X"92",X"02",X"69",X"00",X"8F",X"FF",X"B2",X"00",X"9F",X"FD",X"03",X"FE",
		X"B5",X"00",X"88",X"FF",X"91",X"00",X"60",X"FF",X"3A",X"01",X"66",X"02",X"D5",X"01",X"3F",X"FF",
		X"B7",X"00",X"0A",X"FF",X"87",X"FD",X"79",X"FE",X"C9",X"FD",X"46",X"FE",X"0B",X"FE",X"DB",X"FD",
		X"82",X"00",X"D6",X"FF",X"34",X"00",X"E7",X"FF",X"47",X"00",X"A7",X"FF",X"2B",X"01",X"B7",X"02",
		X"5B",X"01",X"89",X"02",X"04",X"FE",X"83",X"02",X"33",X"01",X"11",X"03",X"98",X"FF",X"54",X"00",
		X"CE",X"FF",X"33",X"00",X"FD",X"FF",X"5E",X"FD",X"92",X"FE",X"A9",X"FD",X"CA",X"FE",X"B4",X"01",
		X"58",X"02",X"B0",X"00",X"E3",X"FD",X"98",X"01",X"1E",X"FE",X"3C",X"FE",X"E5",X"FD",X"69",X"FE",
		X"94",X"FD",X"71",X"00",X"1D",X"00",X"7A",X"FD",X"8C",X"FE",X"D5",X"FD",X"E2",X"01",X"D7",X"01",
		X"4D",X"02",X"0C",X"01",X"B5",X"FD",X"A7",X"FF",X"7C",X"02",X"B0",X"01",X"CB",X"01",X"1B",X"FD",
		X"57",X"00",X"FD",X"FF",X"F8",X"FF",X"66",X"00",X"2E",X"FD",X"86",X"01",X"D6",X"01",X"DF",X"FE",
		X"91",X"01",X"39",X"02",X"BF",X"01",X"52",X"02",X"79",X"00",X"7B",X"FD",X"6A",X"00",X"6B",X"02",
		X"EF",X"00",X"91",X"FD",X"E3",X"FF",X"50",X"02",X"C8",X"01",X"17",X"02",X"DE",X"01",X"F6",X"01",
		X"77",X"FE",X"01",X"FE",X"30",X"FE",X"04",X"FE",X"46",X"FE",X"CF",X"FD",X"F4",X"FF",X"8D",X"02",
		X"6E",X"FF",X"86",X"FD",X"D4",X"FF",X"C3",X"00",X"45",X"FD",X"B6",X"00",X"48",X"02",X"0D",X"FF",
		X"D5",X"FD",X"7E",X"FE",X"D4",X"01",X"72",X"01",X"D7",X"FD",X"5B",X"FE",X"FC",X"FD",X"45",X"FE",
		X"1A",X"FE",X"15",X"FE",X"DB",X"00",X"7F",X"FF",X"4A",X"FD",X"95",X"00",X"02",X"02",X"34",X"02",
		X"01",X"FF",X"FF",X"FD",X"2A",X"FE",X"9F",X"FE",X"8C",X"01",X"A8",X"FD",X"C2",X"FE",X"5C",X"FD",
		X"CD",X"00",X"9C",X"FF",X"83",X"00",X"AF",X"FF",X"BA",X"FD",X"37",X"FE",X"1B",X"00",X"77",X"00",
		X"40",X"FD",X"ED",X"FE",X"A5",X"FD",X"4B",X"02",X"24",X"01",X"A8",X"FE",X"A0",X"FD",X"E4",X"FF",
		X"D3",X"00",X"54",X"FD",X"F7",X"00",X"9E",X"FF",X"7B",X"00",X"CE",X"FF",X"94",X"00",X"37",X"03",
		X"BF",X"FE",X"30",X"01",X"1E",X"FF",X"2C",X"FE",X"FD",X"FD",X"0E",X"FF",X"F9",X"00",X"44",X"FF",
		X"35",X"01",X"8E",X"FD",X"B7",X"FE",X"D6",X"FD",X"A4",X"FE",X"D2",X"FD",X"B2",X"01",X"A9",X"01",
		X"0F",X"FF",X"4C",X"01",X"10",X"FE",X"1C",X"01",X"4D",X"02",X"47",X"FE",X"87",X"FE",X"CC",X"FD",
		X"A1",X"FF",X"F7",X"00",X"C6",X"FD",X"9C",X"FE",X"E1",X"FD",X"DB",X"00",X"57",X"02",X"C2",X"01",
		X"07",X"FF",X"A7",X"01",X"BD",X"01",X"C6",X"FD",X"BF",X"FE",X"D8",X"FD",X"56",X"02",X"F5",X"00",
		X"8F",X"FF",X"C3",X"00",X"4C",X"FF",X"9B",X"02",X"2E",X"00",X"80",X"FD",X"52",X"01",X"2E",X"FF",
		X"2F",X"01",X"2A",X"02",X"29",X"02",X"25",X"01",X"30",X"FF",X"4B",X"01",X"8E",X"FD",X"FF",X"FE",
		X"88",X"01",X"54",X"02",X"AF",X"01",X"54",X"02",X"96",X"01",X"9C",X"02",X"4E",X"FF",X"A9",X"00",
		X"B3",X"FF",X"9D",X"FD",X"ED",X"FE",X"65",X"01",X"80",X"02",X"CF",X"00",X"39",X"FE",X"31",X"FE",
		X"67",X"FE",X"09",X"FE",X"10",X"FF",X"2B",X"02",X"D5",X"01",X"3B",X"02",X"36",X"00",X"95",X"FD",
		X"0B",X"01",X"1F",X"02",X"E7",X"01",X"13",X"02",X"7C",X"01",X"C1",X"FE",X"5E",X"02",X"8A",X"01",
		X"84",X"02",X"EB",X"FF",X"14",X"FE",X"44",X"FE",X"56",X"FE",X"23",X"FE",X"7B",X"FE",X"E5",X"FD",
		X"94",X"00",X"3F",X"02",X"D7",X"01",X"00",X"02",X"FC",X"01",X"98",X"01",X"23",X"FE",X"7B",X"FE",
		X"E1",X"FD",X"FC",X"FF",X"B5",X"00",X"68",X"FD",X"0B",X"FF",X"5E",X"FD",X"6A",X"00",X"13",X"00",
		X"ED",X"FF",X"60",X"02",X"E7",X"01",X"44",X"FF",X"DE",X"00",X"41",X"FF",X"91",X"01",X"85",X"01",
		X"98",X"FE",X"D2",X"02",X"1C",X"01",X"F7",X"02",X"EA",X"FE",X"18",X"01",X"17",X"FF",X"6C",X"01",
		X"47",X"00",X"D1",X"FF",X"8E",X"00",X"4F",X"FD",X"04",X"FF",X"99",X"FD",X"31",X"FF",X"C0",X"00",
		X"62",X"FF",X"B3",X"01",X"63",X"02",X"3C",X"00",X"22",X"FE",X"1F",X"FE",X"B9",X"00",X"CC",X"FF",
		X"86",X"FD",X"62",X"02",X"78",X"FF",X"82",X"00",X"E4",X"FF",X"B4",X"FD",X"A6",X"01",X"F4",X"01",
		X"DC",X"01",X"2E",X"02",X"CC",X"00",X"26",X"FF",X"7B",X"02",X"AE",X"01",X"4F",X"00",X"4F",X"FD",
		X"A2",X"01",X"CB",X"FE",X"93",X"01",X"9D",X"01",X"2F",X"FE",X"A1",X"00",X"76",X"02",X"69",X"FE",
		X"CE",X"FE",X"0B",X"01",X"15",X"FF",X"FD",X"01",X"FD",X"01",X"A7",X"00",X"6C",X"FD",X"F9",X"00",
		X"89",X"FF",X"84",X"00",X"7D",X"02",X"73",X"01",X"53",X"02",X"10",X"01",X"3F",X"FE",X"E9",X"00",
		X"37",X"02",X"6C",X"FE",X"30",X"02",X"E2",X"00",X"7B",X"FE",X"D1",X"FD",X"23",X"00",X"78",X"00",
		X"86",X"FD",X"F6",X"00",X"0F",X"02",X"FE",X"FE",X"31",X"01",X"57",X"02",X"EC",X"00",X"12",X"FF",
		X"33",X"02",X"8C",X"01",X"D0",X"FE",X"E7",X"FD",X"28",X"FF",X"E1",X"01",X"0D",X"02",X"74",X"00",
		X"C0",X"FD",X"B6",X"FE",X"D0",X"FD",X"44",X"01",X"D3",X"01",X"15",X"02",X"44",X"01",X"8C",X"FE",
		X"E6",X"FD",X"97",X"FF",X"0C",X"02",X"A0",X"01",X"87",X"FE",X"84",X"02",X"2C",X"00",X"E9",X"FF",
		X"47",X"00",X"B1",X"FF",X"5A",X"02",X"BB",X"01",X"47",X"FF",X"C7",X"00",X"3A",X"FF",X"70",X"01",
		X"85",X"01",X"D0",X"FD",X"73",X"FF",X"6F",X"02",X"CD",X"FF",X"9F",X"FE",X"5D",X"01",X"D4",X"FD",
		X"7B",X"FF",X"8E",X"02",X"7D",X"FF",X"5A",X"00",X"F3",X"FF",X"9F",X"FD",X"9E",X"01",X"97",X"01",
		X"73",X"FE",X"4F",X"FE",X"31",X"FE",X"86",X"FE",X"DA",X"FD",X"5A",X"00",X"36",X"00",X"A0",X"FD",
		X"7D",X"FF",X"19",X"02",X"8E",X"01",X"59",X"02",X"52",X"FF",X"99",X"00",X"95",X"FF",X"EC",X"FD",
		X"84",X"01",X"BD",X"FE",X"8E",X"01",X"98",X"FD",X"E8",X"FF",X"B6",X"01",X"4B",X"02",X"6E",X"FF",
		X"79",X"00",X"C5",X"FF",X"B0",X"FD",X"C4",X"FE",X"F4",X"FD",X"A7",X"FE",X"08",X"FE",X"A0",X"FE",
		X"CC",X"00",X"82",X"FF",X"BD",X"00",X"DB",X"FE",X"B8",X"FD",X"F6",X"FF",X"AE",X"00",X"9D",X"FD",
		X"C5",X"00",X"C5",X"FF",X"46",X"00",X"FC",X"FF",X"16",X"FD",X"34",X"01",X"50",X"FF",X"B2",X"00",
		X"0C",X"02",X"02",X"FF",X"ED",X"FD",X"22",X"FF",X"7A",X"01",X"60",X"02",X"5A",X"00",X"6F",X"FE",
		X"EE",X"FD",X"BA",X"00",X"C9",X"FF",X"F6",X"FD",X"9F",X"FE",X"4F",X"01",X"15",X"02",X"AB",X"01",
		X"12",X"02",X"21",X"FF",X"02",X"01",X"15",X"02",X"F8",X"FD",X"5F",X"FF",X"97",X"01",X"5A",X"02",
		X"F6",X"FF",X"DD",X"FF",X"48",X"02",X"9B",X"01",X"EF",X"01",X"BC",X"01",X"B9",X"FE",X"57",X"FE",
		X"28",X"FE",X"DA",X"00",X"85",X"FF",X"A4",X"00",X"4D",X"FF",X"A6",X"FD",X"92",X"FF",X"DB",X"00",
		X"14",X"FE",X"A3",X"FF",X"A5",X"02",X"41",X"FF",X"91",X"00",X"20",X"02",X"B2",X"01",X"B8",X"01",
		X"6A",X"FE",X"CF",X"FE",X"35",X"02",X"ED",X"FE",X"25",X"01",X"C2",X"FE",X"59",X"FE",X"2B",X"FE",
		X"5E",X"FF",X"EB",X"01",X"11",X"02",X"DC",X"FF",X"18",X"00",X"40",X"00",X"80",X"FD",X"11",X"FF",
		X"E4",X"FD",X"6E",X"02",X"80",X"00",X"B0",X"FF",X"B2",X"00",X"43",X"FE",X"94",X"01",X"A1",X"01",
		X"DE",X"FD",X"C6",X"FF",X"9C",X"00",X"40",X"FF",X"D2",X"02",X"18",X"FF",X"C6",X"00",X"86",X"FF",
		X"A2",X"00",X"7E",X"FF",X"1D",X"01",X"49",X"02",X"50",X"01",X"63",X"02",X"17",X"00",X"7C",X"FE",
		X"CD",X"01",X"29",X"01",X"B6",X"FE",X"D2",X"02",X"84",X"FF",X"37",X"00",X"E3",X"01",X"F3",X"01",
		X"18",X"FF",X"46",X"FE",X"57",X"FE",X"70",X"FE",X"A7",X"FE",X"81",X"02",X"0E",X"00",X"C9",X"FF",
		X"EA",X"01",X"F5",X"01",X"DD",X"00",X"1F",X"FF",X"3D",X"02",X"58",X"00",X"AF",X"FD",X"C2",X"00",
		X"BB",X"01",X"FE",X"01",X"9F",X"FE",X"D1",X"FE",X"EB",X"00",X"D5",X"FE",X"AD",X"FD",X"3E",X"00",
		X"F8",X"FF",X"30",X"00",X"EF",X"FF",X"3E",X"00",X"78",X"01",X"9A",X"FD",X"05",X"00",X"55",X"02",
		X"4E",X"FF",X"A6",X"00",X"7C",X"FF",X"C5",X"00",X"F8",X"FE",X"9B",X"FE",X"5A",X"01",X"22",X"FE",
		X"62",X"FE",X"9D",X"FF",X"32",X"02",X"A2",X"01",X"D0",X"FF",X"D7",X"FD",X"D2",X"FE",X"F5",X"FD",
		X"34",X"00",X"4D",X"02",X"28",X"FF",X"CB",X"00",X"63",X"FF",X"E6",X"00",X"B4",X"FE",X"DF",X"FE",
		X"6C",X"01",X"91",X"FD",X"3A",X"00",X"BF",X"01",X"F7",X"01",X"98",X"FF",X"F0",X"FD",X"8F",X"01",
		X"5A",X"00",X"0E",X"FE",X"80",X"FE",X"7B",X"00",X"49",X"02",X"43",X"01",X"1E",X"FF",X"E1",X"FD",
		X"64",X"FF",X"9B",X"01",X"F5",X"01",X"7F",X"01",X"09",X"02",X"60",X"01",X"3F",X"02",X"DA",X"FE",
		X"3E",X"01",X"9D",X"01",X"28",X"02",X"4E",X"FF",X"A4",X"00",X"80",X"FF",X"C4",X"00",X"00",X"02",
		X"07",X"FE",X"5C",X"FF",X"FE",X"00",X"E2",X"FD",X"E8",X"FF",X"22",X"02",X"CF",X"FF",X"DD",X"FD",
		X"2F",X"01",X"16",X"FF",X"30",X"FE",X"CC",X"FE",X"C6",X"01",X"97",X"01",X"E6",X"01",X"5E",X"01",
		X"3E",X"FF",X"CE",X"00",X"32",X"FF",X"BC",X"01",X"D7",X"01",X"7B",X"00",X"AE",X"FD",X"CD",X"00",
		X"99",X"FF",X"64",X"00",X"B5",X"FF",X"8D",X"FD",X"89",X"FF",X"80",X"00",X"77",X"FF",X"A7",X"01",
		X"3C",X"FF",X"EC",X"00",X"61",X"02",X"71",X"00",X"87",X"FF",X"9C",X"01",X"11",X"02",X"D7",X"FF",
		X"4A",X"FE",X"49",X"FE",X"F1",X"00",X"C2",X"01",X"F2",X"FE",X"24",X"01",X"5A",X"FE",X"1D",X"FF",
		X"19",X"02",X"3A",X"01",X"4A",X"FF",X"D5",X"00",X"AD",X"FE",X"11",X"FE",X"A4",X"FF",X"0D",X"02",
		X"21",X"00",X"BA",X"FD",X"18",X"01",X"3A",X"FF",X"ED",X"00",X"C2",X"01",X"A3",X"FE",X"14",X"02",
		X"8A",X"00",X"48",X"FF",X"23",X"02",X"52",X"01",X"10",X"02",X"C7",X"00",X"7E",X"FE",X"23",X"FE",
		X"E4",X"FF",X"E8",X"01",X"B6",X"01",X"7D",X"FF",X"64",X"00",X"C2",X"FF",X"4F",X"00",X"B1",X"FF",
		X"E7",X"00",X"8C",X"02",X"BA",X"FF",X"35",X"00",X"F3",X"FF",X"F0",X"FF",X"29",X"02",X"C8",X"00",
		X"C4",X"FD",X"5B",X"00",X"F1",X"FF",X"EC",X"FF",X"46",X"02",X"F8",X"FE",X"3E",X"FE",X"A7",X"FE",
		X"04",X"FE",X"80",X"FF",X"7D",X"00",X"9E",X"FF",X"78",X"00",X"8E",X"FF",X"B3",X"00",X"52",X"FD",
		X"FF",X"FF",X"63",X"01",X"F6",X"01",X"53",X"01",X"F6",X"01",X"4D",X"01",X"FD",X"01",X"3B",X"01",
		X"25",X"02",X"AA",X"00",X"8A",X"FF",X"77",X"00",X"7D",X"FF",X"C3",X"00",X"AA",X"FD",X"7E",X"00",
		X"F5",X"01",X"0D",X"FF",X"37",X"FF",X"53",X"02",X"BA",X"FF",X"10",X"FE",X"BB",X"00",X"80",X"FF",
		X"0C",X"FE",X"7B",X"01",X"4F",X"FE",X"9B",X"FE",X"CB",X"FE",X"8F",X"02",X"8E",X"FF",X"21",X"00",
		X"B6",X"01",X"D2",X"01",X"16",X"FF",X"EB",X"00",X"C0",X"01",X"B4",X"01",X"C9",X"FF",X"EF",X"FD",
		X"0B",X"01",X"2C",X"FF",X"D1",X"00",X"D8",X"FE",X"15",X"FE",X"65",X"FF",X"C5",X"01",X"88",X"01",
		X"A8",X"01",X"89",X"01",X"BC",X"01",X"43",X"FF",X"20",X"FE",X"C5",X"FE",X"49",X"01",X"B5",X"01",
		X"94",X"01",X"45",X"FF",X"A1",X"00",X"17",X"02",X"22",X"01",X"15",X"02",X"72",X"00",X"6E",X"FE",
		X"50",X"FE",X"91",X"FE",X"48",X"FE",X"9A",X"FE",X"44",X"FE",X"AA",X"FE",X"05",X"01",X"F5",X"01",
		X"E4",X"00",X"5C",X"FE",X"C2",X"00",X"49",X"FF",X"F8",X"FD",X"19",X"FF",X"89",X"01",X"F2",X"00",
		X"04",X"FE",X"A8",X"FE",X"94",X"FF",X"83",X"02",X"EF",X"FE",X"A2",X"FE",X"A5",X"00",X"60",X"FF",
		X"BE",X"FD",X"8F",X"FF",X"2F",X"01",X"13",X"02",X"61",X"FE",X"2A",X"FF",X"8D",X"00",X"89",X"FF",
		X"A9",X"00",X"64",X"FE",X"4C",X"FE",X"FB",X"FF",X"29",X"02",X"30",X"FF",X"A1",X"00",X"7F",X"FF",
		X"BE",X"00",X"29",X"02",X"B7",X"00",X"7D",X"FE",X"36",X"FF",X"18",X"02",X"5B",X"FE",X"27",X"02",
		X"4C",X"00",X"B7",X"FF",X"89",X"00",X"3B",X"FE",X"8A",X"FE",X"7D",X"FE",X"70",X"FE",X"8E",X"FE",
		X"E6",X"00",X"03",X"02",X"E6",X"00",X"D6",X"FE",X"FA",X"FD",X"FA",X"FF",X"45",X"00",X"A1",X"FF",
		X"CA",X"01",X"5F",X"FE",X"A9",X"02",X"8C",X"FF",X"54",X"00",X"DB",X"FF",X"10",X"00",X"F8",X"01",
		X"6B",X"01",X"27",X"FF",X"16",X"01",X"B6",X"01",X"8F",X"01",X"6F",X"01",X"EB",X"01",X"FD",X"FF",
		X"CF",X"FF",X"6B",X"00",X"9B",X"FD",X"CD",X"FF",X"71",X"01",X"BC",X"01",X"52",X"01",X"E5",X"01",
		X"3C",X"FF",X"81",X"00",X"7A",X"FF",X"D2",X"FD",X"73",X"FF",X"65",X"00",X"96",X"FF",X"78",X"00",
		X"4C",X"FF",X"3C",X"02",X"93",X"FF",X"20",X"FE",X"83",X"FF",X"D4",X"00",X"B2",X"FD",X"90",X"00",
		X"DE",X"FF",X"11",X"FE",X"CC",X"FE",X"44",X"FE",X"A7",X"01",X"E1",X"00",X"4E",X"FF",X"E5",X"00",
		X"29",X"FE",X"C2",X"FE",X"31",X"FE",X"4F",X"00",X"F1",X"01",X"39",X"FF",X"29",X"FE",X"E8",X"FF",
		X"DE",X"01",X"78",X"01",X"B4",X"FF",X"FB",X"FD",X"F2",X"FE",X"3F",X"FE",X"09",X"02",X"81",X"00",
		X"ED",X"FE",X"D7",X"FD",X"79",X"00",X"C5",X"FF",X"43",X"00",X"EA",X"FF",X"18",X"FE",X"C4",X"FE",
		X"41",X"01",X"3A",X"00",X"FE",X"FD",X"EF",X"FE",X"36",X"FE",X"5B",X"01",X"80",X"01",X"70",X"01",
		X"0F",X"FE",X"C8",X"FF",X"7B",X"00",X"54",X"FF",X"69",X"02",X"3D",X"FF",X"8F",X"00",X"AE",X"FF",
		X"13",X"FE",X"8E",X"01",X"29",X"FE",X"D5",X"00",X"70",X"FF",X"A3",X"00",X"6A",X"FF",X"05",X"01",
		X"7F",X"01",X"3B",X"FE",X"DA",X"FE",X"45",X"FE",X"E4",X"FE",X"15",X"FE",X"AC",X"00",X"C6",X"FF",
		X"29",X"FE",X"30",X"01",X"F3",X"FE",X"63",X"FE",X"1C",X"FF",X"B9",X"01",X"6C",X"01",X"BB",X"01",
		X"2C",X"01",X"16",X"FF",X"9B",X"01",X"75",X"01",X"C1",X"01",X"5D",X"00",X"03",X"FE",X"81",X"00",
		X"CF",X"01",X"4B",X"FF",X"41",X"FE",X"06",X"FF",X"DA",X"00",X"31",X"FF",X"A5",X"01",X"7F",X"01",
		X"8C",X"01",X"9A",X"01",X"26",X"01",X"83",X"FE",X"85",X"FE",X"6C",X"FF",X"11",X"02",X"11",X"01",
		X"1B",X"02",X"12",X"FF",X"D8",X"00",X"87",X"01",X"14",X"FF",X"3F",X"01",X"61",X"01",X"D7",X"FD",
		X"2D",X"00",X"23",X"00",X"D0",X"FE",X"E8",X"00",X"D0",X"FE",X"0F",X"FE",X"2F",X"00",X"FE",X"FF",
		X"1D",X"00",X"F7",X"FF",X"2C",X"00",X"E0",X"FF",X"FC",X"FD",X"17",X"FF",X"50",X"01",X"0F",X"01",
		X"12",X"FF",X"3C",X"01",X"94",X"FD",X"AC",X"00",X"F2",X"00",X"2B",X"FF",X"D3",X"01",X"78",X"00",
		X"3B",X"FE",X"DE",X"FE",X"3C",X"FE",X"CD",X"00",X"88",X"FF",X"40",X"FE",X"9B",X"01",X"35",X"01",
		X"09",X"02",X"3B",X"00",X"DB",X"FF",X"49",X"00",X"C7",X"FF",X"6B",X"00",X"4A",X"FE",X"95",X"02",
		X"9F",X"FF",X"2F",X"00",X"3F",X"00",X"04",X"FE",X"E5",X"00",X"73",X"FF",X"56",X"FE",X"82",X"01",
		X"20",X"01",X"83",X"FE",X"41",X"FF",X"F3",X"01",X"40",X"00",X"1E",X"FE",X"8D",X"00",X"D7",X"FF",
		X"1B",X"00",X"6F",X"02",X"8B",X"FF",X"2D",X"00",X"B1",X"01",X"79",X"01",X"78",X"01",X"7B",X"01",
		X"E7",X"FE",X"93",X"01",X"D5",X"00",X"9E",X"FE",X"5A",X"FE",X"F6",X"FF",X"7E",X"00",X"D6",X"FD",
		X"EC",X"00",X"6E",X"01",X"A5",X"01",X"44",X"01",X"D8",X"01",X"8F",X"FF",X"76",X"FE",X"9F",X"FE",
		X"F2",X"00",X"2B",X"FF",X"12",X"01",X"53",X"FE",X"8F",X"FF",X"6E",X"01",X"D6",X"01",X"B3",X"FF",
		X"34",X"00",X"FF",X"FF",X"10",X"FE",X"05",X"FF",X"DB",X"00",X"ED",X"01",X"96",X"FF",X"4D",X"FE",
		X"F6",X"00",X"7A",X"01",X"E1",X"FE",X"6E",X"FE",X"E2",X"FE",X"25",X"FE",X"13",X"00",X"27",X"00",
		X"DF",X"FF",X"61",X"00",X"DC",X"FD",X"2E",X"01",X"5D",X"01",X"02",X"FF",X"7B",X"FE",X"B5",X"FE",
		X"9C",X"FE",X"9D",X"FE",X"B9",X"FE",X"7F",X"FE",X"E6",X"FE",X"33",X"FE",X"E5",X"FF",X"4C",X"00",
		X"D0",X"FF",X"7B",X"00",X"23",X"FE",X"E2",X"FE",X"91",X"00",X"D4",X"01",X"BC",X"FE",X"A7",X"FE",
		X"13",X"FF",X"B3",X"01",X"5E",X"01",X"35",X"FF",X"63",X"FE",X"2E",X"FF",X"26",X"01",X"0E",X"FE",
		X"3B",X"00",X"10",X"00",X"14",X"00",X"1C",X"00",X"10",X"00",X"17",X"00",X"F8",X"FD",X"B9",X"01",
		X"2B",X"FE",X"C7",X"FF",X"6D",X"00",X"96",X"FF",X"9F",X"01",X"FD",X"FE",X"8A",X"01",X"F7",X"00",
		X"74",X"FE",X"E4",X"FE",X"67",X"FE",X"28",X"00",X"EC",X"01",X"7B",X"FF",X"7A",X"FE",X"22",X"01",
		X"94",X"01",X"7F",X"01",X"25",X"01",X"3B",X"FE",X"ED",X"FF",X"94",X"00",X"36",X"FE",X"13",X"FF",
		X"3C",X"FE",X"DD",X"FF",X"82",X"00",X"68",X"FF",X"5A",X"02",X"41",X"FF",X"9B",X"00",X"B3",X"01",
		X"1A",X"FF",X"AE",X"FE",X"99",X"01",X"3B",X"01",X"E9",X"01",X"34",X"00",X"B4",X"FF",X"CC",X"01",
		X"65",X"01",X"10",X"01",X"5A",X"FE",X"FD",X"FE",X"51",X"FE",X"4A",X"00",X"A9",X"01",X"73",X"01",
		X"78",X"FF",X"59",X"FE",X"03",X"FF",X"4F",X"FE",X"9A",X"FF",X"A0",X"00",X"5F",X"FF",X"F4",X"01",
		X"1A",X"01",X"EC",X"01",X"56",X"FF",X"4D",X"FF",X"ED",X"01",X"30",X"00",X"41",X"FE",X"8A",X"00",
		X"9C",X"01",X"74",X"01",X"16",X"FF",X"DC",X"FE",X"02",X"01",X"21",X"FF",X"AA",X"01",X"76",X"01",
		X"64",X"00",X"69",X"FF",X"70",X"02",X"F4",X"FE",X"1B",X"FF",X"0F",X"FE",X"88",X"00",X"D6",X"FF",
		X"25",X"00",X"E1",X"01",X"38",X"FF",X"C7",X"00",X"EB",X"01",X"A2",X"00",X"A7",X"FF",X"7B",X"00",
		X"A7",X"FF",X"96",X"00",X"5A",X"FF",X"73",X"02",X"E7",X"FE",X"02",X"01",X"48",X"01",X"D5",X"01",
		X"A9",X"FF",X"2D",X"00",X"D9",X"01",X"2B",X"FF",X"9F",X"FE",X"5B",X"01",X"12",X"01",X"A2",X"FE",
		X"3D",X"FF",X"10",X"02",X"C1",X"FF",X"27",X"00",X"27",X"00",X"3D",X"FE",X"FA",X"FE",X"B2",X"00",
		X"D1",X"01",X"10",X"01",X"DB",X"01",X"33",X"FF",X"C5",X"00",X"42",X"FF",X"B1",X"FE",X"43",X"01",
		X"47",X"FE",X"C8",X"FF",X"99",X"00",X"5E",X"FE",X"F4",X"FE",X"70",X"FE",X"9E",X"00",X"A1",X"01",
		X"48",X"01",X"89",X"01",X"43",X"01",X"A7",X"01",X"61",X"FF",X"97",X"00",X"A5",X"01",X"DA",X"FE",
		X"55",X"01",X"17",X"FE",X"18",X"00",X"0D",X"00",X"0F",X"00",X"0C",X"00",X"16",X"00",X"FF",X"FF",
		X"29",X"00",X"E2",X"FF",X"5C",X"00",X"5C",X"FF",X"4A",X"FE",X"07",X"FF",X"70",X"00",X"FA",X"01",
		X"BC",X"00",X"38",X"FF",X"33",X"FE",X"DA",X"FF",X"98",X"00",X"38",X"FE",X"61",X"00",X"16",X"00",
		X"42",X"FE",X"0C",X"FF",X"AB",X"00",X"B6",X"01",X"56",X"FE",X"9F",X"FF",X"A5",X"00",X"9F",X"FE",
		X"CA",X"FE",X"AE",X"FE",X"11",X"FF",X"9A",X"01",X"B7",X"00",X"4F",X"FE",X"15",X"00",X"81",X"01",
		X"8E",X"01",X"7B",X"FF",X"8D",X"00",X"92",X"FF",X"D2",X"00",X"A5",X"01",X"58",X"01",X"CA",X"00",
		X"24",X"FF",X"17",X"02",X"A4",X"00",X"4B",X"FF",X"25",X"FE",X"03",X"00",X"47",X"00",X"9A",X"FF",
		X"FB",X"01",X"8E",X"FF",X"A1",X"FE",X"C6",X"FE",X"BD",X"FE",X"DA",X"FE",X"7C",X"01",X"C1",X"00",
		X"48",X"FF",X"B9",X"01",X"23",X"01",X"AC",X"01",X"D8",X"FF",X"53",X"FE",X"C2",X"FF",X"A9",X"00",
		X"4B",X"FE",X"20",X"FF",X"55",X"FE",X"DE",X"00",X"6F",X"FF",X"A4",X"FE",X"3D",X"01",X"6C",X"01",
		X"53",X"01",X"88",X"01",X"90",X"00",X"52",X"FE",X"25",X"00",X"C3",X"01",X"7F",X"FF",X"A7",X"FE",
		X"AC",X"FE",X"DA",X"FF",X"B9",X"01",X"3D",X"01",X"D3",X"FF",X"45",X"FE",X"2F",X"FF",X"58",X"FE",
		X"70",X"FF",X"26",X"01",X"27",X"01",X"E4",X"FD",X"A8",X"00",X"A9",X"FF",X"6B",X"00",X"CA",X"FF",
		X"99",X"FE",X"A4",X"FE",X"13",X"00",X"5A",X"00",X"44",X"FE",X"26",X"FF",X"83",X"FE",X"24",X"01",
		X"0E",X"FF",X"89",X"01",X"A9",X"00",X"6C",X"FF",X"94",X"01",X"64",X"01",X"40",X"00",X"40",X"FE",
		X"C2",X"00",X"7B",X"01",X"3D",X"FF",X"AB",X"FE",X"C5",X"FE",X"3C",X"00",X"CF",X"01",X"01",X"01",
		X"AA",X"FF",X"66",X"00",X"CB",X"FF",X"63",X"00",X"B4",X"FF",X"AA",X"00",X"58",X"FE",X"2A",X"00",
		X"C4",X"01",X"7B",X"FF",X"AD",X"FE",X"E4",X"FE",X"00",X"01",X"D6",X"FE",X"47",X"00",X"CC",X"01",
		X"25",X"FF",X"D3",X"FE",X"B1",X"FE",X"32",X"FF",X"6D",X"01",X"DD",X"00",X"31",X"FE",X"6B",X"00",
		X"EF",X"FF",X"2B",X"00",X"1B",X"00",X"45",X"FE",X"35",X"FF",X"7C",X"FE",X"50",X"FF",X"54",X"01",
		X"C1",X"FF",X"6D",X"FE",X"2A",X"FF",X"7D",X"FE",X"78",X"FF",X"D8",X"00",X"8E",X"FE",X"E0",X"FF",
		X"A8",X"00",X"3D",X"FE",X"58",X"FF",X"51",X"FE",X"36",X"01",X"0A",X"FF",X"34",X"FF",X"B9",X"00",
		X"8E",X"FF",X"CF",X"00",X"9D",X"FE",X"15",X"FF",X"10",X"01",X"A4",X"01",X"B1",X"00",X"60",X"FF",
		X"C4",X"01",X"0E",X"01",X"C0",X"01",X"B5",X"FF",X"A8",X"FE",X"C1",X"00",X"96",X"01",X"D4",X"FE",
		X"42",X"FF",X"45",X"01",X"7B",X"01",X"37",X"01",X"95",X"01",X"E7",X"00",X"79",X"FF",X"CD",X"00",
		X"BD",X"FE",X"CC",X"FE",X"C7",X"FF",X"F4",X"01",X"79",X"FF",X"77",X"00",X"A1",X"01",X"2E",X"01",
		X"84",X"01",X"F8",X"00",X"D4",X"FE",X"E8",X"FE",X"B0",X"FE",X"D6",X"FF",X"BA",X"01",X"CF",X"00",
		X"E4",X"FE",X"D4",X"FE",X"DA",X"FE",X"E6",X"FE",X"B6",X"FE",X"57",X"00",X"A6",X"01",X"26",X"01",
		X"81",X"01",X"32",X"01",X"7B",X"01",X"2F",X"01",X"90",X"01",X"7E",X"00",X"76",X"FE",X"2E",X"00",
		X"8E",X"01",X"41",X"01",X"DE",X"00",X"3A",X"FE",X"60",X"00",X"25",X"00",X"72",X"FE",X"A9",X"00",
		X"89",X"01",X"25",X"FF",X"2E",X"01",X"FF",X"00",X"E6",X"FE",X"A4",X"FE",X"DD",X"FF",X"7B",X"00",
		X"77",X"FF",X"38",X"02",X"03",X"FF",X"C5",X"FF",X"47",X"01",X"7B",X"01",X"0F",X"01",X"B5",X"01",
		X"44",X"FF",X"CA",X"00",X"41",X"FF",X"FE",X"FE",X"E5",X"00",X"34",X"FF",X"A5",X"01",X"66",X"00",
		X"85",X"FE",X"1C",X"00",X"B3",X"01",X"7A",X"FF",X"71",X"00",X"C8",X"01",X"01",X"00",X"B5",X"FE",
		X"EC",X"FE",X"C5",X"FE",X"B5",X"00",X"95",X"FF",X"8B",X"00",X"94",X"FF",X"BF",X"00",X"AD",X"FE",
		X"A5",X"FF",X"BB",X"01",X"F6",X"FF",X"86",X"FE",X"A8",X"00",X"B0",X"FF",X"6D",X"00",X"9D",X"FF",
		X"46",X"FE",X"BB",X"00",X"37",X"01",X"78",X"01",X"04",X"01",X"46",X"FF",X"C2",X"FE",X"EB",X"01",
		X"00",X"00",X"1D",X"00",X"14",X"00",X"08",X"00",X"3A",X"00",X"66",X"FE",X"29",X"FF",X"B3",X"FE",
		X"37",X"01",X"3C",X"01",X"5C",X"01",X"39",X"01",X"57",X"01",X"3B",X"01",X"35",X"01",X"B3",X"FE",
		X"8A",X"FF",X"AD",X"00",X"3C",X"FF",X"16",X"02",X"68",X"FF",X"86",X"00",X"B2",X"FF",X"6B",X"00",
		X"B9",X"FF",X"71",X"00",X"A0",X"FF",X"B0",X"00",X"C8",X"FE",X"C0",X"00",X"62",X"FF",X"C9",X"FE",
		X"76",X"01",X"06",X"01",X"89",X"01",X"ED",X"00",X"C1",X"01",X"91",X"FF",X"67",X"00",X"C3",X"FF",
		X"5D",X"00",X"AC",X"FF",X"73",X"FE",X"31",X"FF",X"99",X"FE",X"22",X"FF",X"9D",X"FE",X"3A",X"FF",
		X"D0",X"00",X"9F",X"01",X"D9",X"00",X"D7",X"01",X"D7",X"FF",X"30",X"00",X"FE",X"FF",X"1C",X"00",
		X"14",X"00",X"5D",X"FE",X"1F",X"01",X"25",X"FF",X"0A",X"01",X"98",X"FE",X"A9",X"FF",X"4F",X"01",
		X"31",X"01",X"1D",X"FF",X"6B",X"01",X"8B",X"00",X"7A",X"FF",X"76",X"01",X"38",X"01",X"37",X"00",
		X"4E",X"FE",X"E4",X"00",X"67",X"FF",X"C4",X"00",X"3E",X"01",X"0B",X"FF",X"8F",X"01",X"5F",X"00",
		X"80",X"FF",X"B0",X"01",X"E2",X"FF",X"F2",X"FE",X"9A",X"01",X"59",X"00",X"E6",X"FE",X"A5",X"FE",
		X"4A",X"00",X"15",X"00",X"68",X"FE",X"F1",X"00",X"37",X"01",X"47",X"01",X"29",X"01",X"54",X"01",
		X"B2",X"00",X"72",X"FE",X"25",X"00",X"42",X"00",X"79",X"FE",X"31",X"FF",X"8E",X"FE",X"DC",X"FF",
		X"7A",X"01",X"0D",X"00",X"6D",X"FE",X"CD",X"00",X"77",X"FF",X"CB",X"FE",X"22",X"01",X"FE",X"00",
		X"BE",X"FE",X"1E",X"FF",X"8A",X"FE",X"2E",X"00",X"30",X"00",X"A4",X"FE",X"F0",X"FE",X"AC",X"00",
		X"AB",X"00",X"76",X"FE",X"26",X"FF",X"F5",X"FF",X"E6",X"01",X"F0",X"FE",X"2A",X"01",X"F7",X"00",
		X"A3",X"01",X"51",X"00",X"D2",X"FF",X"5F",X"00",X"94",X"FF",X"C3",X"01",X"A3",X"FF",X"CF",X"FE",
		X"F2",X"FE",X"BF",X"00",X"6F",X"01",X"01",X"01",X"7A",X"01",X"75",X"FF",X"D7",X"FE",X"E4",X"FE",
		X"00",X"FF",X"BC",X"FE",X"8D",X"FF",X"A7",X"00",X"48",X"FF",X"F7",X"01",X"79",X"FF",X"73",X"00",
		X"D1",X"FF",X"AE",X"FE",X"0D",X"FF",X"0E",X"01",X"22",X"00",X"8E",X"FE",X"30",X"FF",X"BC",X"FE",
		X"00",X"01",X"02",X"FF",X"4A",X"FF",X"EB",X"00",X"84",X"FE",X"0B",X"00",X"62",X"00",X"9B",X"FE",
		X"2B",X"FF",X"BC",X"FE",X"BF",X"00",X"50",X"01",X"0D",X"FF",X"08",X"FF",X"BF",X"FE",X"B5",X"00",
		X"91",X"FF",X"C3",X"FE",X"28",X"FF",X"55",X"01",X"8F",X"00",X"A2",X"FF",X"98",X"00",X"6C",X"FF",
		X"F3",X"01",X"7A",X"FF",X"FA",X"FE",X"80",X"00",X"9C",X"01",X"BA",X"00",X"91",X"FF",X"FD",X"00",
		X"6F",X"01",X"F5",X"00",X"86",X"01",X"A5",X"00",X"B5",X"FF",X"67",X"00",X"BF",X"FF",X"74",X"00",
		X"88",X"FF",X"D0",X"01",X"92",X"FF",X"DC",X"FE",X"9E",X"00",X"A5",X"FF",X"9D",X"00",X"A4",X"01",
		X"68",X"00",X"9E",X"FF",X"3E",X"01",X"65",X"FF",X"B1",X"00",X"2B",X"FF",X"CA",X"FE",X"29",X"FF",
		X"A3",X"FE",X"2B",X"00",X"47",X"00",X"73",X"FE",X"CD",X"00",X"8B",X"FF",X"D6",X"FE",X"1D",X"01",
		X"25",X"01",X"4C",X"01",X"AD",X"00",X"9A",X"FE",X"08",X"00",X"4C",X"01",X"3B",X"01",X"BA",X"00",
		X"DA",X"FE",X"EB",X"FE",X"DD",X"FF",X"7D",X"01",X"0F",X"01",X"DE",X"FF",X"8D",X"FE",X"51",X"FF",
		X"9B",X"FE",X"96",X"FF",X"9D",X"00",X"ED",X"FE",X"89",X"FF",X"BD",X"01",X"C2",X"FF",X"0E",X"FF",
		X"B4",X"FE",X"E3",X"FF",X"68",X"00",X"8C",X"FF",X"E0",X"01",X"59",X"FF",X"9E",X"00",X"98",X"FF",
		X"A6",X"00",X"5E",X"01",X"1F",X"01",X"DD",X"00",X"C4",X"FE",X"11",X"FF",X"A0",X"FF",X"D4",X"01",
		X"6B",X"FF",X"9A",X"FF",X"A3",X"00",X"BD",X"FE",X"22",X"FF",X"E0",X"FE",X"1E",X"FF",X"D3",X"FE",
		X"C6",X"00",X"3A",X"01",X"3C",X"01",X"D4",X"00",X"50",X"FF",X"7C",X"01",X"54",X"00",X"CC",X"FE",
		X"2A",X"FF",X"C1",X"FE",X"9D",X"00",X"B5",X"FF",X"BA",X"FE",X"39",X"FF",X"BD",X"FE",X"6E",X"00",
		X"5A",X"01",X"11",X"01",X"3F",X"01",X"1B",X"01",X"0A",X"01",X"B2",X"FE",X"CA",X"FF",X"1B",X"01",
		X"6B",X"01",X"DC",X"FF",X"12",X"00",X"85",X"01",X"E4",X"00",X"74",X"01",X"13",X"00",X"CF",X"FE",
		X"1C",X"FF",X"E9",X"FE",X"19",X"FF",X"BD",X"00",X"47",X"01",X"B2",X"FE",X"C7",X"FF",X"78",X"00",
		X"02",X"FF",X"C7",X"FE",X"56",X"00",X"FC",X"FF",X"13",X"00",X"A3",X"01",X"17",X"FF",X"05",X"01",
		X"D5",X"FE",X"7B",X"00",X"36",X"01",X"32",X"01",X"31",X"FF",X"44",X"FF",X"AB",X"00",X"84",X"FF",
		X"BE",X"00",X"B5",X"FE",X"32",X"FF",X"EE",X"FE",X"FC",X"FE",X"73",X"00",X"D6",X"FF",X"50",X"00",
		X"D5",X"FF",X"75",X"00",X"3C",X"FF",X"3E",X"00",X"A0",X"01",X"E9",X"FE",X"59",X"FF",X"9D",X"FE",
		X"DC",X"FF",X"73",X"00",X"FF",X"FE",X"FD",X"FE",X"1D",X"FF",X"F6",X"FE",X"17",X"FF",X"81",X"00",
		X"D4",X"FF",X"56",X"00",X"DA",X"FF",X"74",X"00",X"39",X"FF",X"DA",X"FE",X"04",X"01",X"28",X"FF",
		X"76",X"01",X"51",X"00",X"E5",X"FF",X"5D",X"00",X"AF",X"FF",X"A5",X"01",X"AF",X"FF",X"F2",X"FE",
		X"1D",X"FF",X"0C",X"FF",X"0C",X"01",X"F0",X"00",X"EF",X"FE",X"96",X"FF",X"62",X"01",X"DF",X"00",
		X"8E",X"FF",X"B3",X"00",X"03",X"FF",X"87",X"FF",X"92",X"01",X"01",X"00",X"06",X"FF",X"F2",X"FE",
		X"87",X"00",X"49",X"01",X"1B",X"01",X"FD",X"00",X"5E",X"FF",X"EC",X"00",X"A8",X"FE",X"00",X"00",
		X"1A",X"01",X"53",X"01",X"97",X"00",X"AD",X"FF",X"8C",X"00",X"80",X"FF",X"A6",X"01",X"D9",X"FF",
		X"DA",X"FE",X"90",X"00",X"C0",X"FF",X"C0",X"FE",X"65",X"FF",X"FE",X"00",X"DA",X"00",X"33",X"FF",
		X"CC",X"01",X"BA",X"FF",X"37",X"00",X"26",X"01",X"51",X"01",X"52",X"00",X"B2",X"FF",X"5D",X"01",
		X"11",X"01",X"05",X"00",X"A4",X"FE",X"EC",X"00",X"F1",X"00",X"86",X"FF",X"A6",X"00",X"23",X"FF",
		X"FB",X"FE",X"2D",X"FF",X"E1",X"FE",X"1E",X"00",X"6F",X"01",X"9B",X"FF",X"5F",X"FF",X"B2",X"01",
		X"B9",X"FF",X"45",X"00",X"0B",X"00",X"C5",X"FE",X"3E",X"FF",X"F5",X"FE",X"2A",X"FF",X"06",X"FF",
		X"1D",X"FF",X"17",X"FF",X"03",X"FF",X"D7",X"FF",X"96",X"01",X"9E",X"FF",X"5E",X"00",X"53",X"01",
		X"0D",X"01",X"6B",X"00",X"87",X"FE",X"AF",X"00",X"FF",X"00",X"4F",X"01",X"1E",X"FF",X"6F",X"FF",
		X"C4",X"00",X"8F",X"01",X"0F",X"00",X"1E",X"00",X"0E",X"00",X"27",X"00",X"01",X"00",X"37",X"00",
		X"EC",X"FF",X"CC",X"FE",X"0E",X"01",X"31",X"01",X"C8",X"FF",X"4C",X"00",X"E8",X"FF",X"4C",X"00",
		X"D4",X"FF",X"7B",X"00",X"40",X"FF",X"FB",X"FE",X"29",X"FF",X"16",X"FF",X"FD",X"FE",X"58",X"00",
		X"08",X"00",X"B2",X"FE",X"09",X"01",X"00",X"01",X"30",X"01",X"11",X"01",X"CF",X"FF",X"D0",X"FE",
		X"F2",X"00",X"4F",X"FF",X"F8",X"00",X"B5",X"FE",X"07",X"00",X"48",X"00",X"B9",X"FF",X"94",X"01",
		X"9F",X"FF",X"54",X"00",X"60",X"01",X"37",X"FF",X"49",X"FF",X"F3",X"00",X"2E",X"01",X"FB",X"00",
		X"31",X"01",X"3E",X"FF",X"48",X"FF",X"08",X"01",X"D6",X"00",X"AA",X"FE",X"2F",X"00",X"22",X"00",
		X"E5",X"FF",X"70",X"01",X"D5",X"00",X"42",X"01",X"47",X"FF",X"1D",X"FF",X"12",X"FF",X"25",X"FF",
		X"13",X"FF",X"24",X"FF",X"23",X"FF",X"07",X"01",X"D4",X"00",X"FA",X"FE",X"A3",X"FF",X"6C",X"01",
		X"05",X"00",X"E1",X"FF",X"95",X"01",X"60",X"FF",X"AA",X"00",X"81",X"FF",X"DF",X"00",X"D2",X"00",
		X"75",X"FF",X"CF",X"00",X"B8",X"FE",X"73",X"FF",X"C3",X"FE",X"B8",X"FF",X"C7",X"00",X"80",X"01",
		X"EA",X"FF",X"31",X"00",X"05",X"00",X"25",X"00",X"14",X"00",X"B4",X"FE",X"77",X"FF",X"A8",X"00",
		X"58",X"01",X"8D",X"00",X"0B",X"FF",X"B0",X"FF",X"69",X"01",X"9A",X"00",X"9F",X"FF",X"F0",X"00",
		X"3F",X"01",X"46",X"00",X"FB",X"FE",X"1E",X"FF",X"2D",X"00",X"70",X"01",X"4D",X"FF",X"E0",X"00",
		X"D2",X"00",X"89",X"FF",X"AA",X"00",X"05",X"FF",X"2A",X"FF",X"23",X"FF",X"09",X"FF",X"37",X"00",
		X"5F",X"01",X"5F",X"00",X"04",X"FF",X"35",X"FF",X"11",X"FF",X"3C",X"FF",X"01",X"FF",X"BA",X"00",
		X"01",X"01",X"7F",X"FF",X"A9",X"00",X"6E",X"FF",X"5A",X"01",X"34",X"00",X"B2",X"FF",X"95",X"01",
		X"84",X"FF",X"87",X"00",X"92",X"00",X"7A",X"FF",X"A2",X"01",X"9E",X"FF",X"49",X"00",X"40",X"01",
		X"81",X"FF",X"9D",X"00",X"49",X"01",X"93",X"00",X"89",X"FF",X"32",X"01",X"64",X"00",X"DA",X"FE",
		X"67",X"FF",X"D0",X"FE",X"AB",X"00",X"E7",X"00",X"5A",X"01",X"D2",X"FF",X"42",X"00",X"EC",X"FF",
		X"40",X"00",X"E1",X"FF",X"58",X"00",X"9F",X"FF",X"D4",X"FE",X"A9",X"FF",X"22",X"01",X"63",X"00",
		X"ED",X"FE",X"43",X"FF",X"1A",X"FF",X"1C",X"FF",X"96",X"00",X"9B",X"FF",X"D0",X"00",X"19",X"00",
		X"F0",X"FF",X"80",X"01",X"A9",X"00",X"3F",X"01",X"25",X"FF",X"13",X"01",X"9C",X"FE",X"36",X"00",
		X"07",X"00",X"16",X"00",X"31",X"00",X"E9",X"FE",X"46",X"FF",X"1D",X"FF",X"29",X"FF",X"49",X"FF",
		X"F1",X"00",X"0B",X"01",X"F8",X"00",X"0E",X"01",X"5A",X"FF",X"42",X"FF",X"0C",X"01",X"B0",X"00",
		X"E3",X"FE",X"F1",X"FF",X"15",X"01",X"13",X"01",X"F0",X"FF",X"E1",X"FE",X"B5",X"00",X"FE",X"00",
		X"6A",X"FF",X"F8",X"00",X"B7",X"00",X"FB",X"FE",X"B5",X"00",X"78",X"FF",X"10",X"FF",X"31",X"FF",
		X"71",X"FF",X"47",X"01",X"B9",X"00",X"62",X"01",X"B4",X"FF",X"54",X"00",X"EC",X"FF",X"EA",X"FE",
		X"DA",X"00",X"EB",X"00",X"21",X"FF",X"8C",X"FF",X"0C",X"01",X"FE",X"00",X"E2",X"00",X"5C",X"FF",
		X"05",X"FF",X"60",X"FF",X"D8",X"FE",X"2A",X"00",X"15",X"00",X"0B",X"00",X"33",X"00",X"CD",X"FE",
		X"6C",X"FF",X"89",X"00",X"1C",X"01",X"2E",X"FF",X"5E",X"01",X"2B",X"00",X"D6",X"FF",X"02",X"01",
		X"64",X"FF",X"08",X"01",X"9F",X"00",X"02",X"FF",X"5B",X"FF",X"EE",X"FE",X"50",X"00",X"14",X"00",
		X"D3",X"FE",X"C9",X"00",X"EE",X"00",X"14",X"01",X"D5",X"00",X"36",X"01",X"47",X"00",X"C8",X"FF",
		X"8B",X"00",X"AA",X"FE",X"E3",X"FF",X"44",X"00",X"DD",X"FF",X"5C",X"00",X"A9",X"FF",X"7B",X"01",
		X"9F",X"FF",X"27",X"FF",X"7F",X"00",X"AE",X"FF",X"03",X"FF",X"3D",X"01",X"A0",X"00",X"6F",X"01",
		X"E1",X"FF",X"33",X"00",X"FC",X"FF",X"23",X"00",X"D6",X"00",X"ED",X"FE",X"4B",X"FF",X"C6",X"FF",
		X"78",X"01",X"82",X"FF",X"7C",X"00",X"BE",X"FF",X"62",X"00",X"C6",X"FF",X"6A",X"00",X"A5",X"FF",
		X"FF",X"00",X"F4",X"00",X"F0",X"00",X"F9",X"00",X"EA",X"00",X"F7",X"00",X"F5",X"00",X"72",X"00",
		X"B4",X"FE",X"82",X"00",X"C5",X"FF",X"47",X"00",X"26",X"01",X"57",X"FF",X"27",X"FF",X"40",X"FF",
		X"10",X"FF",X"B5",X"FF",X"0F",X"01",X"E8",X"00",X"EC",X"00",X"0B",X"01",X"B8",X"FF",X"49",X"00",
		X"55",X"01",X"E1",X"FF",X"F9",X"FF",X"51",X"01",X"75",X"FF",X"8B",X"00",X"93",X"FF",X"B6",X"00",
		X"D5",X"00",X"F7",X"FE",X"D1",X"FF",X"84",X"00",X"BD",X"FE",X"66",X"00",X"F4",X"FF",X"F9",X"FE",
		X"90",X"00",X"AB",X"FF",X"D5",X"FE",X"6B",X"00",X"E4",X"FF",X"0C",X"FF",X"48",X"FF",X"9B",X"00",
		X"66",X"FF",X"23",X"FF",X"76",X"FF",X"4B",X"01",X"F9",X"FF",X"17",X"00",X"15",X"00",X"08",X"00",
		X"24",X"00",X"C5",X"FE",X"F4",X"00",X"CB",X"00",X"E6",X"00",X"FC",X"FE",X"75",X"FF",X"FB",X"FE",
		X"F5",X"00",X"94",X"00",X"AA",X"FF",X"C5",X"00",X"28",X"01",X"29",X"00",X"33",X"FF",X"14",X"FF",
		X"4E",X"00",X"09",X"01",X"E1",X"00",X"EA",X"00",X"EF",X"00",X"DF",X"00",X"F5",X"00",X"DD",X"00",
		X"A9",X"FF",X"08",X"FF",X"F2",X"00",X"DA",X"FE",X"03",X"00",X"12",X"00",X"11",X"00",X"06",X"00",
		X"1C",X"00",X"FC",X"FF",X"29",X"00",X"EE",X"FF",X"3E",X"00",X"D1",X"FF",X"6D",X"00",X"43",X"FF",
		X"92",X"FF",X"1E",X"01",X"C6",X"00",X"DA",X"00",X"4E",X"FF",X"3A",X"01",X"24",X"00",X"CF",X"FF",
		X"0B",X"01",X"E3",X"00",X"F7",X"FF",X"EE",X"FE",X"74",X"FF",X"59",X"00",X"B9",X"FF",X"C3",X"FE",
		X"02",X"00",X"19",X"00",X"01",X"00",X"2C",X"00",X"50",X"FF",X"9D",X"00",X"42",X"FF",X"0E",X"FF",
		X"01",X"00",X"44",X"00",X"01",X"FF",X"56",X"FF",X"34",X"FF",X"38",X"FF",X"51",X"FF",X"16",X"FF",
		X"AB",X"FF",X"65",X"00",X"C4",X"FF",X"69",X"00",X"A2",X"FF",X"5C",X"01",X"52",X"00",X"B7",X"FF",
		X"F3",X"00",X"D4",X"00",X"09",X"01",X"EC",X"FF",X"09",X"00",X"3C",X"01",X"9D",X"00",X"19",X"01",
		X"10",X"FF",X"BD",X"FF",X"55",X"00",X"B7",X"FF",X"F3",X"00",X"E6",X"00",X"CD",X"00",X"08",X"01",
		X"64",X"00",X"49",X"FF",X"09",X"FF",X"30",X"00",X"09",X"00",X"FD",X"FF",X"38",X"01",X"A0",X"00",
		X"08",X"01",X"21",X"FF",X"A2",X"FF",X"82",X"00",X"1E",X"FF",X"C3",X"FF",X"33",X"01",X"DE",X"FF",
		X"37",X"FF",X"29",X"FF",X"94",X"00",X"68",X"00",X"E6",X"FE",X"3E",X"00",X"0B",X"01",X"A8",X"FF",
		X"5B",X"00",X"C8",X"FF",X"60",X"00",X"79",X"FF",X"54",X"FF",X"4A",X"01",X"00",X"00",X"62",X"FF",
		X"F8",X"FE",X"7C",X"00",X"C0",X"FF",X"39",X"FF",X"20",X"FF",X"1D",X"00",X"31",X"00",X"E8",X"FE",
		X"9A",X"00",X"A9",X"FF",X"1D",X"FF",X"6B",X"FF",X"13",X"FF",X"C8",X"FF",X"6F",X"00",X"29",X"FF",
		X"42",X"FF",X"03",X"00",X"31",X"01",X"A3",X"FF",X"3C",X"FF",X"99",X"00",X"FE",X"00",X"BD",X"00",
		X"08",X"01",X"9D",X"FF",X"75",X"00",X"FE",X"00",X"C8",X"00",X"E8",X"00",X"D4",X"00",X"DA",X"00",
		X"EB",X"00",X"36",X"00",X"F6",X"FE",X"54",X"00",X"FB",X"00",X"94",X"FF",X"86",X"00",X"DA",X"00",
		X"65",X"FF",X"F9",X"00",X"BB",X"00",X"BD",X"FF",X"14",X"FF",X"E0",X"00",X"FC",X"FE",X"E2",X"FF",
		X"9D",X"00",X"36",X"01",X"C1",X"FF",X"48",X"00",X"DA",X"FF",X"42",X"00",X"D3",X"FF",X"5B",X"00",
		X"15",X"01",X"7F",X"00",X"55",X"FF",X"3B",X"FF",X"76",X"00",X"BE",X"FF",X"53",X"00",X"CB",X"FF",
		X"57",X"00",X"AC",X"FF",X"FE",X"00",X"BD",X"00",X"DF",X"00",X"C8",X"00",X"DE",X"00",X"A6",X"FF",
		X"19",X"FF",X"86",X"FF",X"A2",X"00",X"09",X"01",X"3B",X"00",X"B9",X"FF",X"09",X"01",X"88",X"00",
		X"8D",X"FF",X"E8",X"00",X"63",X"00",X"01",X"FF",X"20",X"00",X"2A",X"00",X"F8",X"FE",X"85",X"FF",
		X"11",X"FF",X"CA",X"00",X"A9",X"00",X"09",X"01",X"54",X"00",X"67",X"FF",X"0B",X"FF",X"1C",X"00",
		X"A5",X"00",X"99",X"FF",X"88",X"00",X"20",X"FF",X"6A",X"FF",X"1B",X"FF",X"36",X"00",X"14",X"00",
		X"EE",X"FE",X"BB",X"00",X"9D",X"00",X"B7",X"FF",X"5A",X"00",X"B1",X"FF",X"D1",X"00",X"D4",X"00",
		X"BE",X"00",X"DE",X"00",X"B5",X"00",X"E7",X"00",X"A4",X"00",X"07",X"01",X"EC",X"FF",X"F5",X"FF",
		X"15",X"01",X"99",X"FF",X"3E",X"FF",X"46",X"FF",X"68",X"FF",X"C3",X"00",X"CC",X"00",X"C2",X"00",
		X"DF",X"00",X"29",X"00",X"15",X"FF",X"6E",X"FF",X"2B",X"FF",X"6C",X"FF",X"1E",X"FF",X"04",X"00",
		X"00",X"01",X"CD",X"FF",X"28",X"FF",X"66",X"FF",X"6C",X"00",X"AC",X"FF",X"9D",X"00",X"F0",X"00",
		X"5A",X"00",X"1B",X"FF",X"FE",X"FF",X"EA",X"00",X"C1",X"00",X"DF",X"FF",X"0E",X"FF",X"87",X"FF",
		X"08",X"FF",X"52",X"00",X"F4",X"FF",X"12",X"FF",X"98",X"00",X"7F",X"FF",X"66",X"FF",X"BD",X"00",
		X"E0",X"00",X"49",X"00",X"B7",X"FF",X"84",X"00",X"BF",X"FE",X"A1",X"00",X"96",X"FF",X"7B",X"00",
		X"87",X"FF",X"DD",X"FF",X"19",X"01",X"B5",X"FF",X"43",X"FF",X"56",X"FF",X"84",X"00",X"8F",X"FF",
		X"CB",X"00",X"73",X"00",X"47",X"FF",X"3D",X"FF",X"01",X"00",X"44",X"00",X"E9",X"FE",X"98",X"00",
		X"A2",X"FF",X"4D",X"FF",X"A1",X"00",X"40",X"FF",X"55",X"00",X"D9",X"FF",X"41",X"00",X"0A",X"01",
		X"7C",X"00",X"70",X"FF",X"7C",X"FF",X"10",X"01",X"1B",X"00",X"43",X"FF",X"61",X"FF",X"3B",X"FF",
		X"62",X"00",X"CF",X"FF",X"4B",X"00",X"C6",X"FF",X"8D",X"00",X"E7",X"00",X"AD",X"00",X"C1",X"FF",
		X"5B",X"00",X"0C",X"01",X"51",X"00",X"B9",X"FF",X"CA",X"00",X"BD",X"00",X"CF",X"00",X"14",X"00",
		X"06",X"FF",X"84",X"00",X"AE",X"FF",X"6D",X"00",X"EC",X"00",X"78",X"00",X"61",X"FF",X"4A",X"FF",
		X"64",X"FF",X"49",X"FF",X"61",X"FF",X"70",X"FF",X"F8",X"00",X"7F",X"00",X"1E",X"01",X"C0",X"FF",
		X"46",X"00",X"D3",X"FF",X"48",X"00",X"C6",X"FF",X"66",X"00",X"7A",X"FF",X"93",X"FF",X"65",X"00",
		X"B9",X"FF",X"69",X"00",X"27",X"FF",X"5F",X"FF",X"9C",X"FF",X"6A",X"00",X"B6",X"FF",X"66",X"00",
		X"A1",X"FF",X"2C",X"01",X"6D",X"00",X"04",X"01",X"7C",X"00",X"03",X"01",X"5A",X"00",X"D4",X"FF",
		X"46",X"00",X"B7",X"FF",X"E9",X"00",X"23",X"00",X"26",X"FF",X"84",X"FF",X"26",X"FF",X"DE",X"FF",
		X"C5",X"00",X"C3",X"00",X"AB",X"00",X"D9",X"00",X"B7",X"FF",X"43",X"FF",X"70",X"FF",X"89",X"00",
		X"56",X"FF",X"A4",X"FF",X"CA",X"00",X"C0",X"00",X"3C",X"00",X"09",X"FF",X"5E",X"00",X"7E",X"00",
		X"2B",X"FF",X"E5",X"FF",X"F3",X"00",X"EA",X"FF",X"42",X"FF",X"62",X"FF",X"5C",X"00",X"BE",X"FF",
		X"19",X"FF",X"CE",X"FF",X"42",X"00",X"CD",X"FF",X"62",X"00",X"21",X"FF",X"8D",X"FF",X"2C",X"FF",
		X"67",X"00",X"C4",X"00",X"C5",X"00",X"2D",X"00",X"0D",X"FF",X"72",X"00",X"C3",X"FF",X"50",X"00",
		X"BC",X"FF",X"33",X"FF",X"84",X"FF",X"41",X"FF",X"80",X"FF",X"41",X"FF",X"88",X"FF",X"2D",X"FF",
		X"54",X"00",X"B9",X"00",X"D9",X"00",X"26",X"00",X"55",X"FF",X"50",X"FF",X"4A",X"00",X"E8",X"FF",
		X"31",X"FF",X"7F",X"FF",X"6F",X"FF",X"A3",X"00",X"3A",X"FF",X"95",X"FF",X"2B",X"FF",X"1A",X"00",
		X"C7",X"00",X"BB",X"00",X"B9",X"00",X"CA",X"FF",X"47",X"00",X"18",X"01",X"AE",X"FF",X"5B",X"00",
		X"CC",X"FF",X"5B",X"00",X"D2",X"00",X"B8",X"00",X"7F",X"00",X"98",X"FF",X"E6",X"00",X"38",X"00",
		X"26",X"FF",X"45",X"00",X"F3",X"FF",X"1A",X"00",X"F9",X"00",X"84",X"00",X"E1",X"00",X"89",X"00",
		X"E8",X"00",X"A1",X"FF",X"6B",X"FF",X"51",X"FF",X"9A",X"FF",X"94",X"00",X"DF",X"00",X"3A",X"00",
		X"6A",X"FF",X"41",X"FF",X"3A",X"00",X"F5",X"FF",X"18",X"00",X"F9",X"00",X"75",X"00",X"C3",X"FF",
		X"81",X"00",X"D6",X"00",X"92",X"00",X"CF",X"00",X"70",X"FF",X"7C",X"FF",X"42",X"FF",X"CF",X"FF",
		X"67",X"00",X"27",X"FF",X"21",X"00",X"2B",X"00",X"19",X"FF",X"7A",X"00",X"AD",X"00",X"BC",X"00",
		X"A6",X"00",X"9E",X"00",X"39",X"FF",X"DE",X"FF",X"B0",X"00",X"C4",X"00",X"78",X"00",X"AA",X"FF",
		X"AE",X"00",X"BC",X"00",X"42",X"00",X"23",X"FF",X"3F",X"00",X"02",X"00",X"2D",X"FF",X"8B",X"00",
		X"9F",X"00",X"8E",X"FF",X"53",X"FF",X"83",X"FF",X"45",X"FF",X"EB",X"FF",X"B2",X"00",X"8D",X"FF",
		X"B5",X"00",X"9B",X"00",X"CB",X"00",X"30",X"00",X"3E",X"FF",X"19",X"00",X"E8",X"00",X"A2",X"FF",
		X"64",X"00",X"AF",X"FF",X"91",X"00",X"7F",X"00",X"A2",X"FF",X"BD",X"00",X"B6",X"00",X"18",X"00",
		X"DF",X"FF",X"CD",X"00",X"0D",X"FF",X"0F",X"00",X"34",X"00",X"38",X"FF",X"30",X"00",X"0A",X"00",
		X"2E",X"FF",X"9C",X"FF",X"4B",X"00",X"B1",X"FF",X"5F",X"FF",X"F0",X"00",X"25",X"00",X"6D",X"FF",
		X"D2",X"FF",X"00",X"01",X"59",X"00",X"0A",X"01",X"E8",X"FF",X"22",X"00",X"FE",X"FF",X"03",X"00",
		X"D4",X"00",X"C6",X"FF",X"42",X"FF",X"A9",X"FF",X"40",X"00",X"DF",X"FF",X"3D",X"00",X"8E",X"FF",
		X"2C",X"FF",X"3D",X"00",X"E5",X"FF",X"31",X"00",X"E0",X"FF",X"A7",X"FF",X"D7",X"00",X"9B",X"00",
		X"16",X"00",X"2F",X"FF",X"6A",X"00",X"B0",X"00",X"90",X"FF",X"84",X"FF",X"9E",X"00",X"BA",X"00",
		X"42",X"00",X"B3",X"FF",X"F8",X"00",X"D1",X"FF",X"17",X"00",X"DD",X"00",X"96",X"FF",X"81",X"FF",
		X"46",X"FF",X"41",X"00",X"E8",X"FF",X"29",X"00",X"EB",X"FF",X"2E",X"FF",X"C0",X"FF",X"58",X"00",
		X"73",X"FF",X"B7",X"FF",X"D7",X"00",X"7C",X"00",X"C9",X"00",X"7F",X"00",X"C9",X"00",X"78",X"00",
		X"CD",X"00",X"43",X"FF",X"55",X"00",X"CF",X"FF",X"3E",X"00",X"B4",X"00",X"9C",X"FF",X"4F",X"FF",
		X"C8",X"FF",X"45",X"00",X"C6",X"FF",X"B3",X"00",X"B4",X"00",X"ED",X"FF",X"15",X"00",X"0B",X"00",
		X"2C",X"FF",X"A5",X"00",X"86",X"00",X"BC",X"00",X"84",X"00",X"BB",X"00",X"80",X"00",X"C2",X"00",
		X"5A",X"00",X"C4",X"FF",X"52",X"00",X"66",X"FF",X"76",X"FF",X"75",X"FF",X"6E",X"FF",X"7D",X"FF",
		X"64",X"FF",X"62",X"00",X"AF",X"00",X"93",X"00",X"AD",X"00",X"62",X"00",X"60",X"FF",X"84",X"FF",
		X"74",X"FF",X"84",X"00",X"60",X"FF",X"9A",X"FF",X"3E",X"FF",X"16",X"00",X"1B",X"00",X"63",X"FF",
		X"6B",X"FF",X"51",X"00",X"CC",X"FF",X"56",X"00",X"B7",X"00",X"9A",X"00",X"64",X"00",X"A3",X"FF",
		X"D0",X"00",X"7A",X"FF",X"B1",X"00",X"4F",X"00",X"BE",X"FF",X"AD",X"00",X"90",X"00",X"AD",X"00",
		X"07",X"00",X"3F",X"FF",X"65",X"00",X"BF",X"FF",X"6A",X"FF",X"95",X"00",X"8E",X"00",X"B1",X"00",
		X"43",X"00",X"66",X"FF",X"79",X"FF",X"9B",X"FF",X"69",X"00",X"9E",X"FF",X"CC",X"00",X"6C",X"00",
		X"CE",X"00",X"DF",X"FF",X"6B",X"FF",X"33",X"00",X"CB",X"00",X"78",X"FF",X"B4",X"00",X"38",X"00",
		X"E9",X"FF",X"1E",X"00",X"EE",X"FF",X"29",X"00",X"62",X"FF",X"6D",X"FF",X"D6",X"FF",X"39",X"00",
		X"D6",X"FF",X"47",X"00",X"3B",X"FF",X"9D",X"FF",X"1D",X"00",X"D3",X"00",X"67",X"00",X"B3",X"00",
		X"3F",X"FF",X"F7",X"FF",X"1C",X"00",X"ED",X"FF",X"38",X"00",X"4B",X"FF",X"9B",X"FF",X"64",X"FF",
		X"93",X"FF",X"66",X"FF",X"98",X"FF",X"5A",X"FF",X"42",X"00",X"A2",X"00",X"9B",X"00",X"7D",X"00",
		X"BD",X"FF",X"52",X"00",X"BC",X"FF",X"70",X"00",X"2F",X"FF",X"37",X"00",X"F5",X"FF",X"11",X"00",
		X"13",X"00",X"28",X"FF",X"2A",X"00",X"16",X"00",X"5B",X"FF",X"34",X"00",X"BA",X"00",X"A4",X"FF",
		X"89",X"FF",X"85",X"00",X"7B",X"00",X"67",X"FF",X"9B",X"FF",X"5C",X"FF",X"09",X"00",X"B5",X"00",
		X"F0",X"FF",X"57",X"FF",X"6F",X"00",X"90",X"00",X"9E",X"00",X"85",X"00",X"A4",X"00",X"7E",X"00",
		X"A9",X"00",X"86",X"FF",X"AE",X"FF",X"71",X"00",X"C2",X"00",X"11",X"00",X"FB",X"FF",X"1E",X"00",
		X"E7",X"FF",X"C6",X"00",X"76",X"00",X"DB",X"FF",X"33",X"00",X"C7",X"FF",X"58",X"FF",X"9F",X"FF",
		X"1F",X"00",X"CD",X"00",X"73",X"FF",X"B9",X"00",X"2F",X"00",X"E6",X"FF",X"6F",X"00",X"CD",X"00",
		X"D5",X"FF",X"30",X"00",X"E4",X"FF",X"31",X"00",X"DB",X"FF",X"71",X"FF",X"72",X"00",X"90",X"FF",
		X"75",X"FF",X"4F",X"00",X"C8",X"FF",X"7B",X"FF",X"79",X"00",X"75",X"FF",X"C4",X"FF",X"A1",X"00",
		X"7C",X"00",X"A9",X"00",X"F9",X"FF",X"63",X"FF",X"44",X"00",X"A6",X"00",X"98",X"FF",X"8F",X"FF",
		X"72",X"FF",X"C4",X"FF",X"95",X"00",X"C6",X"FF",X"40",X"00",X"C3",X"FF",X"4A",X"FF",X"FC",X"FF",
		X"1A",X"00",X"F5",X"FF",X"2F",X"00",X"64",X"FF",X"93",X"FF",X"2F",X"00",X"B1",X"00",X"96",X"FF",
		X"93",X"FF",X"77",X"FF",X"C4",X"FF",X"9A",X"00",X"81",X"00",X"AF",X"FF",X"7C",X"FF",X"8F",X"FF",
		X"B1",X"FF",X"C0",X"00",X"11",X"00",X"86",X"FF",X"86",X"FF",X"92",X"FF",X"83",X"FF",X"96",X"FF",
		X"82",X"FF",X"94",X"FF",X"9A",X"FF",X"B5",X"00",X"2C",X"00",X"92",X"FF",X"7A",X"FF",X"C2",X"FF",
		X"49",X"00",X"CD",X"FF",X"62",X"00",X"49",X"FF",X"39",X"00",X"FA",X"FF",X"16",X"00",X"10",X"00",
		X"4E",X"FF",X"9C",X"00",X"6C",X"FF",X"EB",X"FF",X"26",X"00",X"F9",X"FF",X"28",X"00",X"E5",X"FF",
		X"B4",X"00",X"76",X"00",X"9D",X"00",X"49",X"00",X"58",X"FF",X"34",X"00",X"F8",X"FF",X"1D",X"00",
		X"FF",X"FF",X"21",X"00",X"BA",X"00",X"72",X"FF",X"BB",X"FF",X"61",X"FF",X"FD",X"FF",X"7E",X"00",
		X"A1",X"00",X"6C",X"00",X"AD",X"00",X"5C",X"00",X"CA",X"00",X"E6",X"FF",X"2A",X"00",X"F2",X"FF",
		X"29",X"00",X"EB",X"FF",X"39",X"00",X"96",X"00",X"AE",X"FF",X"63",X"00",X"8F",X"FF",X"83",X"FF",
		X"FC",X"FF",X"2D",X"00",X"DC",X"FF",X"CD",X"00",X"50",X"00",X"B8",X"00",X"52",X"00",X"C5",X"00",
		X"C3",X"FF",X"40",X"00",X"DF",X"FF",X"84",X"FF",X"65",X"00",X"9C",X"00",X"4F",X"00",X"A2",X"FF",
		X"71",X"FF",X"0D",X"00",X"19",X"00",X"EF",X"FF",X"B6",X"00",X"67",X"00",X"EB",X"FF",X"28",X"00",
		X"CC",X"00",X"C1",X"FF",X"40",X"00",X"E1",X"FF",X"7F",X"FF",X"A5",X"FF",X"77",X"00",X"65",X"00",
		X"7F",X"FF",X"D3",X"FF",X"B0",X"00",X"F8",X"FF",X"01",X"00",X"A4",X"00",X"70",X"00",X"DE",X"FF",
		X"38",X"00",X"A3",X"00",X"60",X"FF",X"5F",X"00",X"C6",X"FF",X"4D",X"00",X"C2",X"FF",X"71",X"00",
		X"61",X"00",X"87",X"FF",X"CE",X"FF",X"B5",X"00",X"EC",X"FF",X"0E",X"00",X"93",X"00",X"80",X"00",
		X"C8",X"FF",X"52",X"00",X"78",X"00",X"AE",X"FF",X"8B",X"00",X"73",X"00",X"80",X"00",X"B9",X"FF",
		X"65",X"00",X"90",X"00",X"3B",X"00",X"C2",X"FF",X"AC",X"00",X"00",X"00",X"7E",X"FF",X"25",X"00",
		X"9F",X"00",X"B6",X"FF",X"4E",X"00",X"B2",X"FF",X"85",X"FF",X"C7",X"FF",X"8C",X"00",X"6D",X"00",
		X"89",X"00",X"6B",X"00",X"90",X"00",X"3D",X"00",X"88",X"FF",X"D8",X"FF",X"AE",X"00",X"D4",X"FF",
		X"1F",X"00",X"ED",X"FF",X"7B",X"FF",X"53",X"00",X"BC",X"FF",X"5F",X"00",X"91",X"00",X"28",X"00",
		X"CA",X"FF",X"8D",X"00",X"89",X"FF",X"C6",X"FF",X"45",X"00",X"72",X"FF",X"FF",X"FF",X"1E",X"00",
		X"78",X"FF",X"AE",X"FF",X"8A",X"FF",X"A3",X"FF",X"9B",X"FF",X"6C",X"00",X"83",X"00",X"45",X"00",
		X"C0",X"FF",X"A1",X"00",X"5A",X"00",X"85",X"00",X"6C",X"FF",X"FC",X"FF",X"14",X"00",X"F0",X"FF",
		X"31",X"00",X"61",X"FF",X"49",X"00",X"DD",X"FF",X"2F",X"00",X"9A",X"00",X"4A",X"00",X"B4",X"FF",
		X"86",X"FF",X"B1",X"FF",X"82",X"FF",X"BA",X"FF",X"75",X"FF",X"ED",X"FF",X"22",X"00",X"EE",X"FF",
		X"32",X"00",X"81",X"FF",X"AC",X"FF",X"9A",X"FF",X"9C",X"FF",X"4B",X"00",X"7A",X"00",X"A9",X"FF",
		X"98",X"FF",X"C6",X"FF",X"92",X"00",X"24",X"00",X"80",X"FF",X"16",X"00",X"94",X"00",X"D7",X"FF",
		X"94",X"FF",X"9F",X"FF",X"F2",X"FF",X"AC",X"00",X"C7",X"FF",X"3C",X"00",X"7E",X"00",X"79",X"00",
		X"5D",X"00",X"AA",X"FF",X"93",X"FF",X"DD",X"FF",X"8A",X"00",X"63",X"00",X"8D",X"00",X"E6",X"FF",
		X"1A",X"00",X"A4",X"00",X"09",X"00",X"9D",X"FF",X"9E",X"FF",X"A9",X"FF",X"96",X"FF",X"52",X"00",
		X"71",X"00",X"AE",X"FF",X"9F",X"FF",X"A7",X"FF",X"97",X"FF",X"E7",X"FF",X"A0",X"00",X"E9",X"FF",
		X"13",X"00",X"91",X"00",X"5C",X"00",X"7F",X"00",X"99",X"FF",X"1B",X"00",X"89",X"00",X"D5",X"FF",
		X"93",X"FF",X"B9",X"FF",X"5C",X"00",X"68",X"00",X"7A",X"FF",X"06",X"00",X"19",X"00",X"EF",X"FF",
		X"90",X"00",X"67",X"00",X"EF",X"FF",X"1F",X"00",X"97",X"00",X"8F",X"FF",X"C7",X"FF",X"7C",X"FF",
		X"5C",X"00",X"5A",X"00",X"92",X"00",X"2F",X"00",X"F8",X"FF",X"17",X"00",X"01",X"00",X"11",X"00",
		X"01",X"00",X"1A",X"00",X"85",X"FF",X"B1",X"FF",X"37",X"00",X"7C",X"00",X"A8",X"FF",X"C0",X"FF",
		X"7C",X"00",X"D5",X"FF",X"A2",X"FF",X"4E",X"00",X"BF",X"FF",X"92",X"FF",X"E0",X"FF",X"70",X"00",
		X"77",X"00",X"19",X"00",X"82",X"FF",X"38",X"00",X"F1",X"FF",X"8C",X"FF",X"C2",X"FF",X"92",X"FF",
		X"C4",X"FF",X"88",X"FF",X"F7",X"FF",X"63",X"00",X"D2",X"FF",X"86",X"FF",X"F1",X"FF",X"24",X"00",
		X"F1",X"FF",X"34",X"00",X"8C",X"FF",X"C0",X"FF",X"95",X"FF",X"41",X"00",X"E3",X"FF",X"96",X"FF",
		X"BC",X"FF",X"B2",X"FF",X"90",X"00",X"22",X"00",X"AE",X"FF",X"A7",X"FF",X"B6",X"FF",X"B9",X"FF",
		X"94",X"00",X"17",X"00",X"B9",X"FF",X"92",X"FF",X"32",X"00",X"FC",X"FF",X"9C",X"FF",X"B6",X"FF",
		X"B4",X"FF",X"5E",X"00",X"77",X"00",X"44",X"00",X"9E",X"FF",X"F3",X"FF",X"8A",X"00",X"3D",X"00",
		X"E6",X"FF",X"38",X"00",X"D7",X"FF",X"8C",X"00",X"4E",X"00",X"8D",X"00",X"DB",X"FF",X"30",X"00",
		X"78",X"00",X"C1",X"FF",X"B9",X"FF",X"71",X"00",X"5D",X"00",X"7A",X"00",X"53",X"00",X"8B",X"00",
		X"E7",X"FF",X"25",X"00",X"4B",X"00",X"A1",X"FF",X"AF",X"FF",X"01",X"00",X"82",X"00",X"58",X"00",
		X"74",X"00",X"D4",X"FF",X"39",X"00",X"D6",X"FF",X"8E",X"FF",X"FB",X"FF",X"1F",X"00",X"F9",X"FF",
		X"25",X"00",X"E8",X"FF",X"A1",X"00",X"C2",X"FF",X"EC",X"FF",X"7D",X"00",X"10",X"00",X"94",X"FF",
		X"31",X"00",X"74",X"00",X"D2",X"FF",X"A8",X"FF",X"CA",X"FF",X"4E",X"00",X"9D",X"FF",X"F7",X"FF",
		X"35",X"00",X"8C",X"FF",X"2B",X"00",X"09",X"00",X"91",X"FF",X"58",X"00",X"BF",X"FF",X"04",X"00",
		X"7A",X"00",X"56",X"00",X"70",X"00",X"D4",X"FF",X"3E",X"00",X"D8",X"FF",X"5E",X"00",X"63",X"00",
		X"6B",X"00",X"27",X"00",X"95",X"FF",X"1D",X"00",X"77",X"00",X"E4",X"FF",X"AA",X"FF",X"4A",X"00",
		X"CC",X"FF",X"A5",X"FF",X"2F",X"00",X"F7",X"FF",X"98",X"FF",X"D7",X"FF",X"35",X"00",X"DD",X"FF",
		X"6B",X"00",X"2D",X"00",X"D6",X"FF",X"9B",X"00",X"D9",X"FF",X"2D",X"00",X"F3",X"FF",X"A7",X"FF",
		X"4C",X"00",X"C8",X"FF",X"B1",X"FF",X"BE",X"FF",X"B0",X"FF",X"49",X"00",X"5C",X"00",X"D2",X"FF",
		X"5E",X"00",X"69",X"00",X"2D",X"00",X"D7",X"FF",X"98",X"00",X"D8",X"FF",X"31",X"00",X"F0",X"FF",
		X"AF",X"FF",X"40",X"00",X"E3",X"FF",X"35",X"00",X"DE",X"FF",X"69",X"00",X"D9",X"FF",X"AB",X"FF",
		X"D7",X"FF",X"3F",X"00",X"B2",X"FF",X"E7",X"FF",X"79",X"00",X"45",X"00",X"7F",X"00",X"DA",X"FF",
		X"36",X"00",X"E5",X"FF",X"39",X"00",X"CD",X"FF",X"BC",X"FF",X"B0",X"FF",X"ED",X"FF",X"62",X"00",
		X"DB",X"FF",X"38",X"00",X"CE",X"FF",X"A1",X"FF",X"0B",X"00",X"13",X"00",X"05",X"00",X"17",X"00",
		X"FD",X"FF",X"86",X"00",X"3F",X"00",X"6F",X"00",X"BB",X"FF",X"78",X"00",X"1F",X"00",X"F1",X"FF",
		X"5F",X"00",X"5D",X"00",X"56",X"00",X"4F",X"00",X"9C",X"FF",X"0F",X"00",X"14",X"00",X"FA",X"FF",
		X"6D",X"00",X"57",X"00",X"EF",X"FF",X"27",X"00",X"6C",X"00",X"B7",X"FF",X"C9",X"FF",X"B5",X"FF",
		X"C3",X"FF",X"E7",X"FF",X"83",X"00",X"F1",X"FF",X"BE",X"FF",X"D3",X"FF",X"81",X"00",X"FB",X"FF",
		X"0B",X"00",X"5F",X"00",X"62",X"00",X"E0",X"FF",X"32",X"00",X"60",X"00",X"5B",X"00",X"3B",X"00",
		X"DE",X"FF",X"43",X"00",X"97",X"FF",X"1F",X"00",X"0D",X"00",X"A6",X"FF",X"F4",X"FF",X"33",X"00",
		X"A0",X"FF",X"17",X"00",X"5D",X"00",X"58",X"00",X"53",X"00",X"5C",X"00",X"CA",X"FF",X"D6",X"FF",
		X"34",X"00",X"E4",X"FF",X"35",X"00",X"D4",X"FF",X"8A",X"00",X"E4",X"FF",X"D4",X"FF",X"A4",X"FF",
		X"0F",X"00",X"0F",X"00",X"FF",X"FF",X"66",X"00",X"51",X"00",X"EE",X"FF",X"B6",X"FF",X"42",X"00",
		X"D7",X"FF",X"57",X"00",X"37",X"00",X"AC",X"FF",X"05",X"00",X"57",X"00",X"5D",X"00",X"F3",X"FF",
		X"18",X"00",X"69",X"00",X"CB",X"FF",X"BF",X"FF",X"0D",X"00",X"6A",X"00",X"40",X"00",X"5E",X"00",
		X"CA",X"FF",X"C7",X"FF",X"D0",X"FF",X"62",X"00",X"43",X"00",X"60",X"00",X"40",X"00",X"68",X"00",
		X"ED",X"FF",X"BE",X"FF",X"2E",X"00",X"60",X"00",X"B8",X"FF",X"1C",X"00",X"5A",X"00",X"ED",X"FF",
		X"1C",X"00",X"FF",X"FF",X"14",X"00",X"02",X"00",X"12",X"00",X"03",X"00",X"17",X"00",X"F5",X"FF",
		X"6C",X"00",X"F0",X"FF",X"B7",X"FF",X"3C",X"00",X"49",X"00",X"E0",X"FF",X"32",X"00",X"C7",X"FF",
		X"C2",X"FF",X"36",X"00",X"55",X"00",X"4C",X"00",X"41",X"00",X"B1",X"FF",X"00",X"00",X"20",X"00",
		X"B5",X"FF",X"D0",X"FF",X"C2",X"FF",X"C9",X"FF",X"2B",X"00",X"ED",X"FF",X"2B",X"00",X"D7",X"FF",
		X"C1",X"FF",X"CB",X"FF",X"2C",X"00",X"ED",X"FF",X"2E",X"00",X"CF",X"FF",X"CA",X"FF",X"BE",X"FF",
		X"05",X"00",X"1F",X"00",X"B3",X"FF",X"D3",X"FF",X"1C",X"00",X"62",X"00",X"3A",X"00",X"D7",X"FF",
		X"D9",X"FF",X"3B",X"00",X"D5",X"FF",X"6F",X"00",X"26",X"00",X"FC",X"FF",X"1B",X"00",X"F7",X"FF",
		X"2A",X"00",X"B2",X"FF",X"15",X"00",X"14",X"00",X"AE",X"FF",X"36",X"00",X"4A",X"00",X"48",X"00",
		X"DA",X"FF",X"4F",X"00",X"2C",X"00",X"C4",X"FF",X"D0",X"FF",X"C9",X"FF",X"DB",X"FF",X"4C",X"00",
		X"33",X"00",X"B6",X"FF",X"0A",X"00",X"4D",X"00",X"4D",X"00",X"43",X"00",X"54",X"00",X"DC",X"FF",
		X"39",X"00",X"CB",X"FF",X"EF",X"FF",X"1F",X"00",X"FA",X"FF",X"1C",X"00",X"FA",X"FF",X"23",X"00",
		X"AC",X"FF",X"FD",X"FF",X"4B",X"00",X"19",X"00",X"ED",X"FF",X"72",X"00",X"DB",X"FF",X"2F",X"00",
		X"44",X"00",X"4E",X"00",X"3C",X"00",X"5A",X"00",X"18",X"00",X"FD",X"FF",X"1B",X"00",X"F3",X"FF",
		X"5E",X"00",X"39",X"00",X"38",X"00",X"B6",X"FF",X"E6",X"FF",X"B7",X"FF",X"21",X"00",X"43",X"00",
		X"4C",X"00",X"3C",X"00",X"4C",X"00",X"C5",X"FF",X"F3",X"FF",X"1E",X"00",X"F1",X"FF",X"4D",X"00",
		X"47",X"00",X"0A",X"00",X"BB",X"FF",X"2B",X"00",X"46",X"00",X"43",X"00",X"42",X"00",X"4C",X"00",
		X"FA",X"FF",X"C4",X"FF",X"DC",X"FF",X"2C",X"00",X"52",X"00",X"23",X"00",X"ED",X"FF",X"2D",X"00",
		X"B4",X"FF",X"19",X"00",X"0B",X"00",X"C2",X"FF",X"24",X"00",X"50",X"00",X"CF",X"FF",X"14",X"00",
		X"05",X"00",X"0A",X"00",X"54",X"00",X"34",X"00",X"EB",X"FF",X"33",X"00",X"30",X"00",X"E1",X"FF",
		X"32",X"00",X"B0",X"FF",X"18",X"00",X"09",X"00",X"C2",X"FF",X"2C",X"00",X"EC",X"FF",X"D0",X"FF",
		X"CC",X"FF",X"19",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"18",X"00",X"ED",X"FF",X"C7",X"FF",
		X"DD",X"FF",X"E8",X"FF",X"5B",X"00",X"02",X"00",X"D0",X"FF",X"15",X"00",X"4E",X"00",X"33",X"00",
		X"F1",X"FF",X"2B",X"00",X"3E",X"00",X"C2",X"FF",X"31",X"00",X"39",X"00",X"46",X"00",X"27",X"00",
		X"EF",X"FF",X"2B",X"00",X"C4",X"FF",X"09",X"00",X"19",X"00",X"BF",X"FF",X"22",X"00",X"3E",X"00",
		X"3C",X"00",X"3A",X"00",X"41",X"00",X"2C",X"00",X"D4",X"FF",X"DA",X"FF",X"D4",X"FF",X"DF",X"FF",
		X"36",X"00",X"30",X"00",X"C9",X"FF",X"FE",X"FF",X"3E",X"00",X"3E",X"00",X"37",X"00",X"45",X"00",
		X"EE",X"FF",X"D7",X"FF",X"D5",X"FF",X"E9",X"FF",X"25",X"00",X"DD",X"FF",X"D0",X"FF",X"01",X"00",
		X"3A",X"00",X"DF",X"FF",X"D0",X"FF",X"FA",X"FF",X"1C",X"00",X"F2",X"FF",X"4F",X"00",X"29",X"00",
		X"4A",X"00",X"E8",X"FF",X"2A",X"00",X"36",X"00",X"ED",X"FF",X"24",X"00",X"ED",X"FF",X"2E",X"00",
		X"BF",X"FF",X"16",X"00",X"29",X"00",X"E4",X"FF",X"CD",X"FF",X"09",X"00",X"11",X"00",X"FC",X"FF",
		X"4C",X"00",X"F5",X"FF",X"D6",X"FF",X"27",X"00",X"37",X"00",X"DF",X"FF",X"E9",X"FF",X"3E",X"00",
		X"30",X"00",X"45",X"00",X"04",X"00",X"05",X"00",X"47",X"00",X"17",X"00",X"EF",X"FF",X"4B",X"00",
		X"FC",X"FF",X"0B",X"00",X"06",X"00",X"CF",X"FF",X"E7",X"FF",X"DC",X"FF",X"35",X"00",X"32",X"00",
		X"39",X"00",X"30",X"00",X"3B",X"00",X"0F",X"00",X"CD",X"FF",X"15",X"00",X"FC",X"FF",X"D7",X"FF",
		X"E1",X"FF",X"FF",X"FF",X"49",X"00",X"F2",X"FF",X"E0",X"FF",X"DC",X"FF",X"E4",X"FF",X"E2",X"FF",
		X"3C",X"00",X"28",X"00",X"45",X"00",X"02",X"00",X"0D",X"00",X"08",X"00",X"07",X"00",X"44",X"00",
		X"ED",X"FF",X"DC",X"FF",X"09",X"00",X"3D",X"00",X"30",X"00",X"FC",X"FF",X"D6",X"FF",X"2D",X"00",
		X"E0",X"FF",X"F1",X"FF",X"34",X"00",X"2F",X"00",X"39",X"00",X"0B",X"00",X"DA",X"FF",X"E4",X"FF",
		X"14",X"00",X"3C",X"00",X"2A",X"00",X"37",X"00",X"2C",X"00",X"34",X"00",X"2E",X"00",X"F3",X"FF",
		X"0A",X"00",X"39",X"00",X"D3",X"FF",X"FC",X"FF",X"00",X"00",X"FD",X"FF",X"03",X"00",X"E2",X"FF",
		X"DB",X"FF",X"14",X"00",X"F3",X"FF",X"14",X"00",X"34",X"00",X"2F",X"00",X"01",X"00",X"DB",X"FF",
		X"E8",X"FF",X"E4",X"FF",X"1A",X"00",X"F2",X"FF",X"18",X"00",X"E8",X"FF",X"3D",X"00",X"FF",X"FF",
		X"00",X"00",X"32",X"00",X"30",X"00",X"F1",X"FF",X"08",X"00",X"F5",X"FF",X"11",X"00",X"3B",X"00",
		X"EE",X"FF",X"0A",X"00",X"34",X"00",X"24",X"00",X"E7",X"FF",X"E7",X"FF",X"E4",X"FF",X"F1",X"FF",
		X"2C",X"00",X"2B",X"00",X"2F",X"00",X"FC",X"FF",X"DE",X"FF",X"09",X"00",X"F0",X"FF",X"E2",X"FF",
		X"F1",X"FF",X"10",X"00",X"E2",X"FF",X"12",X"00",X"ED",X"FF",X"EE",X"FF",X"13",X"00",X"E2",X"FF",
		X"FA",X"FF",X"30",X"00",X"06",X"00",X"E0",X"FF",X"F1",X"FF",X"E4",X"FF",X"21",X"00",X"EB",X"FF",
		X"F5",X"FF",X"1D",X"00",X"E5",X"FF",X"ED",X"FF",X"E8",X"FF",X"EB",X"FF",X"EB",X"FF",X"EA",X"FF",
		X"FB",X"FF",X"38",X"00",X"05",X"00",X"EA",X"FF",X"E8",X"FF",X"1B",X"00",X"FC",X"FF",X"E5",X"FF",
		X"F4",X"FF",X"2B",X"00",X"1D",X"00",X"E8",X"FF",X"ED",X"FF",X"03",X"00",X"36",X"00",X"16",X"00",
		X"FE",X"FF",X"2C",X"00",X"28",X"00",X"2B",X"00",X"09",X"00",X"E1",X"FF",X"1D",X"00",X"27",X"00",
		X"29",X"00",X"26",X"00",X"2A",X"00",X"24",X"00",X"2B",X"00",X"11",X"00",X"E3",X"FF",X"11",X"00",
		X"0C",X"00",X"DE",X"FF",X"0A",X"00",X"22",X"00",X"32",X"00",X"FF",X"FF",X"13",X"00",X"02",X"00",
		X"E7",X"FF",X"F6",X"FF",X"1B",X"00",X"F8",X"FF",X"2D",X"00",X"11",X"00",X"01",X"00",X"2F",X"00",
		X"20",X"00",X"28",X"00",X"24",X"00",X"18",X"00",X"E1",X"FF",X"0F",X"00",X"03",X"00",X"09",X"00",
		X"07",X"00",X"E5",X"FF",X"FB",X"FF",X"E5",X"FF",X"03",X"00",X"10",X"00",X"03",X"00",X"24",X"00",
		X"2B",X"00",X"03",X"00",X"0E",X"00",X"28",X"00",X"24",X"00",X"0F",X"00",X"EA",X"FF",X"F2",X"FF",
		X"0E",X"00",X"2B",X"00",X"F6",X"FF",X"F3",X"FF",X"F0",X"FF",X"FA",X"FF",X"25",X"00",X"20",X"00",
		X"27",X"00",X"0C",X"00",X"EE",X"FF",X"F6",X"FF",X"F1",X"FF",X"18",X"00",X"FE",X"FF",X"EC",X"FF",
		X"12",X"00",X"25",X"00",X"21",X"00",X"FB",X"FF",X"F3",X"FF",X"1D",X"00",X"F2",X"FF",X"00",X"00",
		X"23",X"00",X"22",X"00",X"0F",X"00",X"E8",X"FF",X"19",X"00",X"FE",X"FF",X"15",X"00",X"01",X"00",
		X"17",X"00",X"F5",X"FF",X"10",X"00",X"26",X"00",X"FB",X"FF",X"F2",X"FF",X"FA",X"FF",X"18",X"00",
		X"FA",X"FF",X"29",X"00",X"06",X"00",X"0A",X"00",X"23",X"00",X"1F",X"00",X"03",X"00",X"F0",X"FF",
		X"FE",X"FF",X"15",X"00",X"FE",X"FF",X"20",X"00",X"01",X"00",X"F3",X"FF",X"1C",X"00",X"1C",X"00",
		X"1F",X"00",X"1C",X"00",X"21",X"00",X"0C",X"00",X"F5",X"FF",X"F7",X"FF",X"0F",X"00",X"23",X"00",
		X"FC",X"FF",X"17",X"00",X"FA",X"FF",X"FF",X"FF",X"17",X"00",X"F4",X"FF",X"FB",X"FF",X"18",X"00",
		X"1A",X"00",X"FB",X"FF",X"22",X"00",X"15",X"00",X"23",X"00",X"06",X"00",X"F9",X"FF",X"F5",X"FF",
		X"14",X"00",X"02",X"00",X"F9",X"FF",X"FB",X"FF",X"1E",X"00",X"0F",X"00",X"02",X"00",X"1F",X"00",
		X"1B",X"00",X"15",X"00",X"FF",X"FF",X"16",X"00",X"F1",X"FF",X"0D",X"00",X"0A",X"00",X"07",X"00",
		X"22",X"00",X"FE",X"FF",X"15",X"00",X"FE",X"FF",X"FC",X"FF",X"FB",X"FF",X"FC",X"FF",X"00",X"00",
		X"22",X"00",X"05",X"00",X"0F",X"00",X"13",X"00",X"04",X"00",X"12",X"00",X"F8",X"FF",X"FB",X"FF",
		X"0A",X"00",X"1B",X"00",X"15",X"00",X"04",X"00",X"FC",X"FF",X"19",X"00",X"15",X"00",X"1B",X"00",
		X"15",X"00",X"1C",X"00",X"06",X"00",X"0A",X"00",X"09",X"00",X"FD",X"FF",X"1C",X"00",X"0B",X"00",
		X"FB",X"FF",X"0D",X"00",X"08",X"00",X"0C",X"00",X"09",X"00",X"0A",X"00",X"0A",X"00",X"0D",X"00",
		X"09",X"00",X"0D",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"FC",X"FF",X"10",X"00",X"10",X"00",
		X"FA",X"FF",X"0F",X"00",X"0A",X"00",X"FE",X"FF",X"02",X"00",X"0F",X"00",X"19",X"00",X"12",X"00",
		X"05",X"00",X"15",X"00",X"14",X"00",X"17",X"00",X"08",X"00",X"0B",X"00",X"0B",X"00",X"0A",X"00",
		X"1A",X"00",X"0F",X"00",X"19",X"00",X"04",X"00",X"08",X"00",X"06",X"00",X"FF",X"FF",X"03",X"00",
		X"00",X"00",X"05",X"00",X"13",X"00",X"14",X"00",X"0C",X"00",X"05",X"00",X"18",X"00",X"06",X"00",
		X"02",X"00",X"0E",X"00",X"08",X"00",X"0F",X"00",X"16",X"00",X"04",X"00",X"0C",X"00",X"05",X"00",
		X"0C",X"00",X"13",X"00",X"0E",X"00",X"00",X"00",X"11",X"00",X"0C",X"00",X"01",X"00",X"02",X"00",
		X"06",X"00",X"08",X"00",X"00",X"00",X"0D",X"00",X"11",X"00",X"10",X"00",X"10",X"00",X"08",X"00",
		X"02",X"00",X"05",X"00",X"02",X"00",X"0D",X"00",X"10",X"00",X"0C",X"00",X"01",X"00",X"07",X"00",
		X"08",X"00",X"09",X"00",X"07",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"07",X"00",X"05",X"00",
		X"0D",X"00",X"05",X"00",X"09",X"00",X"0F",X"00",X"0C",X"00",X"07",X"00",X"07",X"00",X"09",X"00",
		X"06",X"00",X"0E",X"00",X"07",X"00",X"04",X"00",X"06",X"00",X"08",X"00",X"0B",X"00",X"09",X"00",
		X"0C",X"00",X"09",X"00",X"0F",X"00",X"08",X"00",X"0B",X"00",X"0B",X"00",X"05",X"00",X"08",X"00",
		X"09",X"00",X"08",X"00",X"07",X"00",X"07",X"00",X"08",X"00",X"08",X"00",X"0B",X"00",X"09",X"00",
		X"0B",X"00",X"0A",X"00",X"0B",X"00",X"0C",X"00",X"0A",X"00",X"0A",X"00",X"09",X"00",X"0A",X"00",
		X"0B",X"00",X"0B",X"00",X"09",X"00",X"09",X"00",X"09",X"00",X"0B",X"00",X"0B",X"00",X"09",X"00",
		X"0A",X"00",X"0A",X"00",X"0A",X"00",X"09",X"00",X"0B",X"00",X"09",X"00",X"0A",X"00",X"0A",X"00",
		X"0C",X"00",X"0B",X"00",X"0B",X"00",X"0B",X"00",X"0B",X"00",X"0B",X"00",X"0A",X"00",X"0A",X"00",
		X"0B",X"00",X"0C",X"00",X"0B",X"00",X"0D",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0D",X"00",
		X"0C",X"00",X"0C",X"00",X"0B",X"00",X"0E",X"00",X"0C",X"00",X"0D",X"00",X"0D",X"00",X"0E",X"00",
		X"0C",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",
		X"0F",X"00",X"0E",X"00",X"0E",X"00",X"0D",X"00",X"0E",X"00",X"0E",X"00",X"0F",X"00",X"0D",X"00",
		X"0E",X"00",X"0E",X"00",X"0F",X"00",X"0E",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",
		X"0E",X"00",X"0E",X"00",X"0F",X"00",X"10",X"00",X"0F",X"00",X"0F",X"00",X"0E",X"00",X"10",X"00",
		X"10",X"00",X"10",X"00",X"11",X"00",X"0F",X"00",X"10",X"00",X"0F",X"00",X"10",X"00",X"12",X"00",
		X"10",X"00",X"0F",X"00",X"10",X"00",X"10",X"00",X"11",X"00",X"12",X"00",X"11",X"00",X"11",X"00",
		X"11",X"00",X"10",X"00",X"13",X"00",X"10",X"00",X"10",X"00",X"10",X"00",X"11",X"00",X"12",X"00",
		X"12",X"00",X"12",X"00",X"13",X"00",X"11",X"00",X"12",X"00",X"12",X"00",X"11",X"00",X"12",X"00",
		X"13",X"00",X"11",X"00",X"12",X"00",X"13",X"00",X"11",X"00",X"13",X"00",X"13",X"00",X"15",X"00",
		X"14",X"00",X"13",X"00",X"13",X"00",X"13",X"00",X"12",X"00",X"14",X"00",X"14",X"00",X"12",X"00",
		X"13",X"00",X"12",X"00",X"15",X"00",X"14",X"00",X"14",X"00",X"14",X"00",X"14",X"00",X"15",X"00",
		X"14",X"00",X"13",X"00",X"14",X"00",X"14",X"00",X"14",X"00",X"14",X"00",X"14",X"00",X"14",X"00",
		X"15",X"00",X"16",X"00",X"16",X"00",X"15",X"00",X"13",X"00",X"15",X"00",X"15",X"00",X"15",X"00",
		X"15",X"00",X"15",X"00",X"15",X"00",X"14",X"00",X"16",X"00",X"17",X"00",X"15",X"00",X"17",X"00",
		X"16",X"00",X"16",X"00",X"16",X"00",X"16",X"00",X"15",X"00",X"14",X"00",X"16",X"00",X"16",X"00",
		X"16",X"00",X"18",X"00",X"16",X"00",X"16",X"00",X"15",X"00",X"17",X"00",X"17",X"00",X"17",X"00",
		X"18",X"00",X"18",X"00",X"16",X"00",X"17",X"00",X"17",X"00",X"17",X"00",X"17",X"00",X"18",X"00",
		X"16",X"00",X"17",X"00",X"17",X"00",X"18",X"00",X"18",X"00",X"17",X"00",X"19",X"00",X"17",X"00",
		X"17",X"00",X"18",X"00",X"16",X"00",X"17",X"00",X"19",X"00",X"19",X"00",X"19",X"00",X"18",X"00",
		X"1A",X"00",X"18",X"00",X"17",X"00",X"18",X"00",X"19",X"00",X"19",X"00",X"19",X"00",X"19",X"00",
		X"18",X"00",X"19",X"00",X"18",X"00",X"17",X"00",X"19",X"00",X"19",X"00",X"18",X"00",X"19",X"00",
		X"19",X"00",X"18",X"00",X"19",X"00",X"19",X"00",X"1A",X"00",X"1A",X"00",X"1A",X"00",X"1A",X"00",
		X"1A",X"00",X"1A",X"00",X"1A",X"00",X"19",X"00",X"1A",X"00",X"1A",X"00",X"1B",X"00",X"1A",X"00",
		X"1B",X"00",X"1B",X"00",X"1A",X"00",X"1A",X"00",X"1A",X"00",X"1A",X"00",X"1B",X"00",X"1B",X"00",
		X"1C",X"00",X"1A",X"00",X"1C",X"00",X"1C",X"00",X"1B",X"00",X"1B",X"00",X"1B",X"00",X"1B",X"00",
		X"1B",X"00",X"1B",X"00",X"1B",X"00",X"1A",X"00",X"1B",X"00",X"1B",X"00",X"1B",X"00",X"1C",X"00",
		X"1C",X"00",X"1C",X"00",X"1D",X"00",X"1B",X"00",X"1B",X"00",X"1C",X"00",X"1C",X"00",X"1B",X"00",
		X"1B",X"00",X"1C",X"00",X"1C",X"00",X"1E",X"00",X"1C",X"00",X"1C",X"00",X"1C",X"00",X"1B",X"00",
		X"1C",X"00",X"1D",X"00",X"1D",X"00",X"1E",X"00",X"1E",X"00",X"1E",X"00",X"1E",X"00",X"1D",X"00",
		X"1D",X"00",X"1B",X"00",X"1D",X"00",X"1D",X"00",X"1D",X"00",X"1D",X"00",X"1C",X"00",X"1D",X"00",
		X"1D",X"00",X"1D",X"00",X"1E",X"00",X"1D",X"00",X"1D",X"00",X"1E",X"00",X"1D",X"00",X"1E",X"00",
		X"1E",X"00",X"1D",X"00",X"1D",X"00",X"1F",X"00",X"1E",X"00",X"1F",X"00",X"1E",X"00",X"1E",X"00",
		X"1F",X"00",X"1E",X"00",X"1E",X"00",X"1E",X"00",X"1E",X"00",X"1E",X"00",X"1D",X"00",X"1D",X"00",
		X"1E",X"00",X"20",X"00",X"1F",X"00",X"1E",X"00",X"1E",X"00",X"1E",X"00",X"1F",X"00",X"1F",X"00",
		X"1F",X"00",X"1E",X"00",X"1E",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",
		X"1F",X"00",X"1F",X"00",X"20",X"00",X"1F",X"00",X"20",X"00",X"1F",X"00",X"1F",X"00",X"21",X"00",
		X"20",X"00",X"20",X"00",X"21",X"00",X"1F",X"00",X"1F",X"00",X"21",X"00",X"20",X"00",X"1F",X"00",
		X"20",X"00",X"20",X"00",X"20",X"00",X"1F",X"00",X"22",X"00",X"20",X"00",X"21",X"00",X"20",X"00",
		X"20",X"00",X"21",X"00",X"21",X"00",X"1F",X"00",X"20",X"00",X"20",X"00",X"21",X"00",X"21",X"00",
		X"22",X"00",X"21",X"00",X"22",X"00",X"21",X"00",X"22",X"00",X"21",X"00",X"22",X"00",X"21",X"00",
		X"21",X"00",X"21",X"00",X"20",X"00",X"20",X"00",X"21",X"00",X"22",X"00",X"21",X"00",X"22",X"00",
		X"21",X"00",X"21",X"00",X"21",X"00",X"21",X"00",X"21",X"00",X"22",X"00",X"21",X"00",X"21",X"00",
		X"20",X"00",X"20",X"00",X"21",X"00",X"24",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FE",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FE",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"1C",X"00",X"7B",X"00",
		X"2E",X"01",X"43",X"02",X"AF",X"03",X"76",X"05",X"87",X"07",X"DF",X"09",X"6F",X"0C",X"32",X"0F",
		X"17",X"12",X"21",X"15",X"3A",X"18",X"72",X"1B",X"03",X"1E",X"5E",X"1F",X"FA",X"1F",X"04",X"20",
		X"B8",X"1F",X"2B",X"1F",X"7B",X"1E",X"B0",X"1D",X"D6",X"1C",X"F2",X"1B",X"0E",X"1B",X"28",X"1A",
		X"45",X"19",X"66",X"18",X"8B",X"17",X"B6",X"16",X"E5",X"15",X"19",X"15",X"53",X"14",X"95",X"13",
		X"DA",X"12",X"27",X"12",X"76",X"11",X"CD",X"10",X"28",X"10",X"8A",X"0F",X"EA",X"0E",X"76",X"0E",
		X"4D",X"0F",X"4E",X"11",X"05",X"14",X"34",X"17",X"A9",X"1A",X"44",X"1E",X"EC",X"21",X"98",X"25",
		X"38",X"29",X"C9",X"2C",X"44",X"30",X"A9",X"33",X"F5",X"36",X"26",X"3A",X"3A",X"3D",X"39",X"40",
		X"1B",X"43",X"E4",X"45",X"93",X"48",X"2A",X"4B",X"A8",X"4D",X"12",X"50",X"61",X"52",X"9D",X"54",
		X"C1",X"56",X"D4",X"58",X"D0",X"5A",X"BA",X"5C",X"90",X"5E",X"55",X"60",X"07",X"62",X"A9",X"63",
		X"38",X"65",X"B8",X"66",X"29",X"68",X"8A",X"69",X"DB",X"6A",X"21",X"6C",X"57",X"6D",X"80",X"6E",
		X"9A",X"6F",X"A9",X"70",X"AD",X"71",X"A4",X"72",X"8F",X"73",X"70",X"74",X"45",X"75",X"10",X"76",
		X"D1",X"76",X"87",X"77",X"35",X"78",X"DB",X"78",X"76",X"79",X"08",X"7A",X"93",X"7A",X"15",X"7B",
		X"8F",X"7B",X"02",X"7C",X"6D",X"7C",X"D4",X"7C",X"2F",X"7D",X"86",X"7D",X"D5",X"7D",X"20",X"7E",
		X"64",X"7E",X"A1",X"7E",X"DA",X"7E",X"0C",X"7F",X"3A",X"7F",X"62",X"7F",X"84",X"7F",X"A4",X"7F",
		X"BC",X"7F",X"D4",X"7F",X"E2",X"7F",X"F0",X"7F",X"F8",X"7F",X"FE",X"7F",X"FD",X"7F",X"FE",X"7F",
		X"F1",X"7F",X"F4",X"7F",X"7A",X"7F",X"90",X"7D",X"AD",X"7A",X"27",X"77",X"41",X"73",X"1F",X"6F",
		X"E2",X"6A",X"9A",X"66",X"59",X"62",X"24",X"5E",X"01",X"5A",X"F8",X"55",X"06",X"52",X"30",X"4E",
		X"76",X"4A",X"D4",X"46",X"51",X"43",X"E8",X"3F",X"99",X"3C",X"64",X"39",X"4B",X"36",X"46",X"33",
		X"5C",X"30",X"88",X"2D",X"CB",X"2A",X"24",X"28",X"92",X"25",X"17",X"23",X"AE",X"20",X"58",X"1E",
		X"18",X"1C",X"E7",X"19",X"C8",X"17",X"BD",X"15",X"C1",X"13",X"D5",X"11",X"FA",X"0F",X"2C",X"0E",
		X"6E",X"0C",X"C0",X"0A",X"1D",X"09",X"8A",X"07",X"04",X"06",X"8D",X"04",X"1C",X"03",X"BE",X"01",
		X"66",X"00",X"1F",X"FF",X"DD",X"FD",X"A8",X"FC",X"7C",X"FB",X"5D",X"FA",X"43",X"F9",X"3B",X"F8",
		X"2B",X"F7",X"7D",X"F6",X"36",X"F7",X"01",X"F9",X"7B",X"FB",X"66",X"FE",X"90",X"01",X"E2",X"04",
		X"41",X"08",X"A2",X"0B",X"FB",X"0E",X"46",X"12",X"7C",X"15",X"9E",X"18",X"A9",X"1B",X"9E",X"1E",
		X"79",X"21",X"3D",X"24",X"E9",X"26",X"7F",X"29",X"FD",X"2B",X"66",X"2E",X"B6",X"30",X"F3",X"32",
		X"1C",X"35",X"30",X"37",X"32",X"39",X"21",X"3B",X"FC",X"3C",X"C6",X"3E",X"80",X"40",X"28",X"42",
		X"BF",X"43",X"49",X"45",X"C1",X"46",X"2E",X"48",X"8A",X"49",X"D8",X"4A",X"19",X"4C",X"4E",X"4D",
		X"75",X"4E",X"91",X"4F",X"9F",X"50",X"A4",X"51",X"9C",X"52",X"8D",X"53",X"70",X"54",X"49",X"55",
		X"19",X"56",X"E0",X"56",X"9D",X"57",X"52",X"58",X"FE",X"58",X"A2",X"59",X"3A",X"5A",X"D3",X"5A",
		X"30",X"5B",X"36",X"5A",X"14",X"58",X"40",X"55",X"F3",X"51",X"62",X"4E",X"A9",X"4A",X"E1",X"46",
		X"17",X"43",X"57",X"3F",X"A4",X"3B",X"05",X"38",X"7B",X"34",X"09",X"31",X"B1",X"2D",X"70",X"2A",
		X"47",X"27",X"39",X"24",X"41",X"21",X"62",X"1E",X"99",X"1B",X"E9",X"18",X"4C",X"16",X"C6",X"13",
		X"55",X"11",X"F6",X"0E",X"AB",X"0C",X"76",X"0A",X"4F",X"08",X"3D",X"06",X"3D",X"04",X"4D",X"02",
		X"6D",X"00",X"9D",X"FE",X"DC",X"FC",X"2A",X"FB",X"85",X"F9",X"F0",X"F7",X"69",X"F6",X"ED",X"F4",
		X"7F",X"F3",X"1F",X"F2",X"C8",X"F0",X"7E",X"EF",X"3F",X"EE",X"0B",X"ED",X"E3",X"EB",X"C5",X"EA",
		X"B0",X"E9",X"A4",X"E8",X"A3",X"E7",X"A9",X"E6",X"BA",X"E5",X"D3",X"E4",X"F5",X"E3",X"1E",X"E3",
		X"50",X"E2",X"87",X"E1",X"C6",X"E0",X"0F",X"E0",X"5D",X"DF",X"B1",X"DE",X"0D",X"DE",X"6E",X"DD",
		X"D6",X"DC",X"44",X"DC",X"B6",X"DB",X"2F",X"DB",X"AD",X"DA",X"2F",X"DA",X"B9",X"D9",X"45",X"D9",
		X"D9",X"D8",X"6E",X"D8",X"0A",X"D8",X"A9",X"D7",X"4D",X"D7",X"F3",X"D6",X"9F",X"D6",X"50",X"D6",
		X"02",X"D6",X"BA",X"D5",X"74",X"D5",X"31",X"D5",X"F1",X"D4",X"B5",X"D4",X"7D",X"D4",X"47",X"D4",
		X"14",X"D4",X"E3",X"D3",X"B7",X"D3",X"8D",X"D3",X"63",X"D3",X"3D",X"D3",X"1B",X"D3",X"F7",X"D2",
		X"D8",X"D2",X"BA",X"D2",X"A0",X"D2",X"88",X"D2",X"71",X"D2",X"5C",X"D2",X"48",X"D2",X"37",X"D2",
		X"2A",X"D2",X"1A",X"D2",X"0E",X"D2",X"03",X"D2",X"F9",X"D1",X"F0",X"D1",X"EB",X"D1",X"E6",X"D1",
		X"E3",X"D1",X"DF",X"D1",X"DE",X"D1",X"DD",X"D1",X"DE",X"D1",X"E1",X"D1",X"E5",X"D1",X"E9",X"D1",
		X"EE",X"D1",X"F4",X"D1",X"FC",X"D1",X"04",X"D2",X"0D",X"D2",X"16",X"D2",X"22",X"D2",X"2D",X"D2",
		X"3A",X"D2",X"47",X"D2",X"56",X"D2",X"61",X"D2",X"73",X"D2",X"81",X"D2",X"94",X"D2",X"A2",X"D2",
		X"B7",X"D2",X"BE",X"D2",X"2D",X"D3",X"03",X"D5",X"D8",X"D7",X"54",X"DB",X"32",X"DF",X"4A",X"E3",
		X"7D",X"E7",X"B9",X"EB",X"ED",X"EF",X"13",X"F4",X"23",X"F8",X"1C",X"FC",X"F7",X"FF",X"B8",X"03",
		X"5B",X"07",X"DF",X"0A",X"47",X"0E",X"95",X"11",X"C5",X"14",X"DB",X"17",X"D4",X"1A",X"B6",X"1D",
		X"7C",X"20",X"2C",X"23",X"BF",X"25",X"43",X"28",X"A6",X"2A",X"FC",X"2C",X"4A",X"2E",X"2C",X"2E",
		X"31",X"2D",X"96",X"2B",X"A2",X"29",X"6A",X"27",X"12",X"25",X"A9",X"22",X"3B",X"20",X"CD",X"1D",
		X"69",X"1B",X"0D",X"19",X"C1",X"16",X"82",X"14",X"56",X"12",X"37",X"10",X"29",X"0E",X"2B",X"0C",
		X"3D",X"0A",X"5F",X"08",X"91",X"06",X"D0",X"04",X"1E",X"03",X"7A",X"01",X"E6",X"FF",X"5D",X"FE",
		X"E2",X"FC",X"74",X"FB",X"11",X"FA",X"B9",X"F8",X"6F",X"F7",X"2D",X"F6",X"FA",X"F4",X"CF",X"F3",
		X"B0",X"F2",X"98",X"F1",X"8B",X"F0",X"86",X"EF",X"8D",X"EE",X"9A",X"ED",X"B0",X"EC",X"CF",X"EB",
		X"F6",X"EA",X"24",X"EA",X"5A",X"E9",X"97",X"E8",X"DB",X"E7",X"26",X"E7",X"77",X"E6",X"CE",X"E5",
		X"2D",X"E5",X"90",X"E4",X"FA",X"E3",X"69",X"E3",X"E0",X"E2",X"5A",X"E2",X"D9",X"E1",X"5E",X"E1",
		X"E7",X"E0",X"76",X"E0",X"07",X"E0",X"9E",X"DF",X"3B",X"DF",X"D9",X"DE",X"7E",X"DE",X"25",X"DE",
		X"CF",X"DD",X"7E",X"DD",X"32",X"DD",X"E7",X"DC",X"A0",X"DC",X"5C",X"DC",X"1C",X"DC",X"DE",X"DB",
		X"A6",X"DB",X"6C",X"DB",X"38",X"DB",X"03",X"DB",X"D8",X"DA",X"A8",X"DA",X"82",X"DA",X"4E",X"DA",
		X"C4",X"DA",X"A7",X"DC",X"6E",X"DF",X"D0",X"E2",X"89",X"E6",X"79",X"EA",X"7F",X"EE",X"8C",X"F2",
		X"91",X"F6",X"89",X"FA",X"68",X"FE",X"33",X"02",X"E2",X"05",X"76",X"09",X"EF",X"0C",X"4A",X"10",
		X"8A",X"13",X"AF",X"16",X"BA",X"19",X"A9",X"1C",X"7F",X"1F",X"3C",X"22",X"E1",X"24",X"6D",X"27",
		X"E4",X"29",X"42",X"2C",X"8C",X"2E",X"C1",X"30",X"E2",X"32",X"EF",X"34",X"E9",X"36",X"CF",X"38",
		X"A6",X"3A",X"6B",X"3C",X"1E",X"3E",X"C0",X"3F",X"53",X"41",X"D5",X"42",X"4C",X"44",X"B1",X"45",
		X"09",X"47",X"52",X"48",X"90",X"49",X"C1",X"4A",X"E6",X"4B",X"FB",X"4C",X"09",X"4E",X"09",X"4F",
		X"02",X"50",X"EA",X"50",X"CE",X"51",X"A2",X"52",X"75",X"53",X"31",X"54",X"FA",X"54",X"38",X"55",
		X"03",X"54",X"D2",X"51",X"FB",X"4E",X"BE",X"4B",X"43",X"48",X"A7",X"44",X"FE",X"40",X"57",X"3D",
		X"B8",X"39",X"28",X"36",X"AD",X"32",X"46",X"2F",X"F6",X"2B",X"BF",X"28",X"A0",X"25",X"98",X"22",
		X"A7",X"1F",X"CF",X"1C",X"0D",X"1A",X"62",X"17",X"CC",X"14",X"4C",X"12",X"E0",X"0F",X"89",X"0D",
		X"44",X"0B",X"12",X"09",X"F2",X"06",X"E4",X"04",X"EA",X"02",X"FE",X"00",X"23",X"FF",X"57",X"FD",
		X"9C",X"FB",X"ED",X"F9",X"51",X"F8",X"BD",X"F6",X"39",X"F5",X"C1",X"F3",X"59",X"F2",X"FB",X"F0",
		X"A9",X"EF",X"62",X"EE",X"28",X"ED",X"F8",X"EB",X"D2",X"EA",X"B6",X"E9",X"A7",X"E8",X"9C",X"E7",
		X"9F",X"E6",X"A9",X"E5",X"BE",X"E4",X"D8",X"E3",X"FE",X"E2",X"23",X"E2",X"A7",X"E1",X"98",X"E2",
		X"96",X"E4",X"3F",X"E7",X"55",X"EA",X"AE",X"ED",X"29",X"F1",X"B1",X"F4",X"3B",X"F8",X"BB",X"FB",
		X"2A",X"FF",X"87",X"02",X"CC",X"05",X"FD",X"08",X"13",X"0C",X"12",X"0F",X"F6",X"11",X"C4",X"14",
		X"7A",X"17",X"18",X"1A",X"9D",X"1C",X"11",X"1F",X"68",X"21",X"B2",X"23",X"DE",X"25",X"02",X"28",
		X"06",X"2A",X"04",X"2C",X"0B",X"2D",X"A2",X"2C",X"5B",X"2B",X"75",X"29",X"36",X"27",X"B5",X"24",
		X"18",X"22",X"66",X"1F",X"B6",X"1C",X"06",X"1A",X"62",X"17",X"CB",X"14",X"43",X"12",X"CC",X"0F",
		X"67",X"0D",X"14",X"0B",X"D1",X"08",X"A2",X"06",X"85",X"04",X"79",X"02",X"7C",X"00",X"94",X"FE",
		X"B8",X"FC",X"EE",X"FA",X"30",X"F9",X"84",X"F7",X"E0",X"F5",X"84",X"F4",X"88",X"F4",X"B3",X"F5",
		X"9B",X"F7",X"F8",X"F9",X"A4",X"FC",X"7A",X"FF",X"63",X"02",X"53",X"05",X"42",X"08",X"24",X"0B",
		X"FA",X"0D",X"BB",X"10",X"6B",X"13",X"05",X"16",X"8E",X"18",X"FE",X"1A",X"5D",X"1D",X"A5",X"1F",
		X"DB",X"21",X"FB",X"23",X"0B",X"26",X"04",X"28",X"F1",X"29",X"C5",X"2B",X"92",X"2D",X"3F",X"2F",
		X"F1",X"30",X"D7",X"31",X"43",X"31",X"CA",X"2F",X"AA",X"2D",X"2E",X"2B",X"6D",X"28",X"90",X"25",
		X"9F",X"22",X"B1",X"1F",X"C3",X"1C",X"E4",X"19",X"11",X"17",X"52",X"14",X"A2",X"11",X"07",X"0F",
		X"7F",X"0C",X"0C",X"0A",X"AC",X"07",X"60",X"05",X"25",X"03",X"FD",X"00",X"E9",X"FE",X"E7",X"FC",
		X"F0",X"FA",X"0F",X"F9",X"3C",X"F7",X"77",X"F5",X"DF",X"F3",X"92",X"F3",X"84",X"F4",X"36",X"F6",
		X"6E",X"F8",X"F3",X"FA",X"AC",X"FD",X"79",X"00",X"50",X"03",X"25",X"06",X"F4",X"08",X"B2",X"0B",
		X"63",X"0E",X"00",X"11",X"89",X"13",X"FF",X"15",X"62",X"18",X"B0",X"1A",X"E7",X"1C",X"0F",X"1F",
		X"22",X"21",X"25",X"23",X"11",X"25",X"F2",X"26",X"B9",X"28",X"79",X"2A",X"1E",X"2C",X"C7",X"2D",
		X"CC",X"2E",X"54",X"2E",X"E9",X"2C",X"D0",X"2A",X"51",X"28",X"8F",X"25",X"AB",X"22",X"B5",X"1F",
		X"BB",X"1C",X"C5",X"19",X"DB",X"16",X"FF",X"13",X"35",X"11",X"7D",X"0E",X"DA",X"0B",X"49",X"09",
		X"CD",X"06",X"65",X"04",X"11",X"02",X"D0",X"FF",X"A1",X"FD",X"84",X"FB",X"7A",X"F9",X"80",X"F7",
		X"9A",X"F5",X"C0",X"F3",X"FA",X"F1",X"4A",X"F0",X"C9",X"EF",X"99",X"F0",X"33",X"F2",X"5D",X"F4",
		X"D7",X"F6",X"88",X"F9",X"51",X"FC",X"28",X"FF",X"FB",X"01",X"C9",X"04",X"89",X"07",X"3A",X"0A",
		X"D8",X"0C",X"63",X"0F",X"DB",X"11",X"3F",X"14",X"8E",X"16",X"CB",X"18",X"F3",X"1A",X"08",X"1D",
		X"0B",X"1F",X"FC",X"20",X"DD",X"22",X"AA",X"24",X"6A",X"26",X"13",X"28",X"BC",X"29",X"E9",X"2A",
		X"9E",X"2A",X"4C",X"29",X"45",X"27",X"D2",X"24",X"17",X"22",X"36",X"1F",X"44",X"1C",X"4A",X"19",
		X"54",X"16",X"6B",X"13",X"8E",X"10",X"C3",X"0D",X"0B",X"0B",X"67",X"08",X"D4",X"05",X"57",X"03",
		X"EE",X"00",X"9A",X"FE",X"57",X"FC",X"29",X"FA",X"0B",X"F8",X"01",X"F6",X"05",X"F4",X"20",X"F2",
		X"45",X"F0",X"81",X"EE",X"C5",X"EC",X"13",X"EC",X"C5",X"EC",X"4D",X"EE",X"6B",X"F0",X"DE",X"F2",
		X"8E",X"F5",X"55",X"F8",X"2E",X"FB",X"06",X"FE",X"D6",X"00",X"99",X"03",X"4E",X"06",X"F2",X"08",
		X"80",X"0B",X"FC",X"0D",X"66",X"10",X"BB",X"12",X"FC",X"14",X"28",X"17",X"43",X"19",X"4B",X"1B",
		X"40",X"1D",X"23",X"1F",X"F8",X"20",X"BA",X"22",X"6D",X"24",X"0E",X"26",X"A2",X"27",X"26",X"29",
		X"9D",X"2A",X"06",X"2C",X"5F",X"2D",X"AD",X"2E",X"F0",X"2F",X"25",X"31",X"4E",X"32",X"6C",X"33",
		X"7E",X"34",X"85",X"35",X"82",X"36",X"75",X"37",X"5E",X"38",X"3E",X"39",X"14",X"3A",X"E1",X"3A",
		X"A6",X"3B",X"62",X"3C",X"17",X"3D",X"C2",X"3D",X"67",X"3E",X"03",X"3F",X"99",X"3F",X"27",X"40",
		X"B1",X"40",X"32",X"41",X"AD",X"41",X"21",X"42",X"91",X"42",X"F9",X"42",X"5E",X"43",X"BC",X"43",
		X"13",X"44",X"68",X"44",X"B7",X"44",X"00",X"45",X"45",X"45",X"87",X"45",X"C4",X"45",X"FA",X"45",
		X"30",X"46",X"5F",X"46",X"8E",X"46",X"B5",X"46",X"DC",X"46",X"FD",X"46",X"1D",X"47",X"37",X"47",
		X"52",X"47",X"62",X"47",X"7A",X"47",X"82",X"47",X"9C",X"47",X"00",X"47",X"FA",X"44",X"14",X"42",
		X"90",X"3E",X"B9",X"3A",X"AB",X"36",X"87",X"32",X"5A",X"2E",X"38",X"2A",X"23",X"26",X"23",X"22",
		X"3B",X"1E",X"6C",X"1A",X"B7",X"16",X"22",X"13",X"A6",X"0F",X"47",X"0C",X"01",X"09",X"D7",X"05",
		X"C6",X"02",X"D1",X"FF",X"F6",X"FC",X"30",X"FA",X"83",X"F7",X"EC",X"F4",X"6C",X"F2",X"FF",X"EF",
		X"BD",X"ED",X"C3",X"EC",X"14",X"ED",X"2E",X"EE",X"D4",X"EF",X"D1",X"F1",X"03",X"F4",X"50",X"F6",
		X"B0",X"F8",X"0E",X"FB",X"6B",X"FD",X"BD",X"FF",X"04",X"02",X"3B",X"04",X"62",X"06",X"7A",X"08",
		X"83",X"0A",X"78",X"0C",X"60",X"0E",X"35",X"10",X"F9",X"11",X"B0",X"13",X"57",X"15",X"F0",X"16",
		X"79",X"18",X"F6",X"19",X"63",X"1B",X"C5",X"1C",X"1B",X"1E",X"5F",X"1F",X"9D",X"20",X"CD",X"21",
		X"F0",X"22",X"0B",X"24",X"19",X"25",X"1E",X"26",X"1A",X"27",X"0B",X"28",X"F3",X"28",X"D0",X"29",
		X"A6",X"2A",X"72",X"2B",X"39",X"2C",X"F4",X"2C",X"A9",X"2D",X"58",X"2E",X"FD",X"2E",X"9B",X"2F",
		X"33",X"30",X"C5",X"30",X"50",X"31",X"D4",X"31",X"52",X"32",X"CB",X"32",X"3F",X"33",X"AB",X"33",
		X"13",X"34",X"76",X"34",X"D4",X"34",X"2E",X"35",X"82",X"35",X"D2",X"35",X"1E",X"36",X"64",X"36",
		X"A8",X"36",X"E6",X"36",X"21",X"37",X"58",X"37",X"8D",X"37",X"BC",X"37",X"E9",X"37",X"12",X"38",
		X"38",X"38",X"5A",X"38",X"7A",X"38",X"97",X"38",X"B2",X"38",X"C9",X"38",X"E0",X"38",X"EF",X"38",
		X"02",X"39",X"09",X"39",X"20",X"39",X"D2",X"38",X"1C",X"37",X"62",X"34",X"01",X"31",X"39",X"2D",
		X"36",X"29",X"16",X"25",X"EB",X"20",X"C7",X"1C",X"B0",X"18",X"AB",X"14",X"BF",X"10",X"EB",X"0C",
		X"34",X"09",X"9A",X"05",X"1A",X"02",X"B9",X"FE",X"71",X"FB",X"45",X"F8",X"33",X"F5",X"3C",X"F2",
		X"5A",X"EF",X"97",X"EC",X"E7",X"E9",X"52",X"E7",X"CD",X"E4",X"68",X"E2",X"0D",X"E0",X"B3",X"DE",
		X"CB",X"DE",X"BB",X"DF",X"4F",X"E1",X"3D",X"E3",X"6B",X"E5",X"BB",X"E7",X"20",X"EA",X"86",X"EC",
		X"EA",X"EE",X"47",X"F1",X"99",X"F3",X"DB",X"F5",X"10",X"F8",X"32",X"FA",X"47",X"FC",X"49",X"FE",
		X"3B",X"00",X"1C",X"02",X"EE",X"03",X"AF",X"05",X"64",X"07",X"08",X"09",X"9E",X"0A",X"26",X"0C",
		X"9F",X"0D",X"0C",X"0F",X"6E",X"10",X"C1",X"11",X"08",X"13",X"44",X"14",X"74",X"15",X"9B",X"16",
		X"B4",X"17",X"C5",X"18",X"CC",X"19",X"C7",X"1A",X"BB",X"1B",X"A5",X"1C",X"85",X"1D",X"5E",X"1E",
		X"2F",X"1F",X"F8",X"1F",X"B6",X"20",X"71",X"21",X"1F",X"22",X"CD",X"22",X"6E",X"23",X"0C",X"24",
		X"9F",X"24",X"32",X"25",X"B8",X"25",X"41",X"26",X"B7",X"26",X"3C",X"27",X"F4",X"26",X"40",X"25",
		X"B2",X"22",X"8B",X"1F",X"0D",X"1C",X"59",X"18",X"8F",X"14",X"BA",X"10",X"EE",X"0C",X"2C",X"09",
		X"82",X"05",X"E9",X"01",X"6C",X"FE",X"06",X"FB",X"BC",X"F7",X"8A",X"F4",X"73",X"F1",X"74",X"EE",
		X"90",X"EB",X"C4",X"E8",X"0F",X"E6",X"72",X"E3",X"EC",X"E0",X"7C",X"DE",X"21",X"DC",X"DC",X"D9",
		X"A8",X"D7",X"AA",X"D5",X"FE",X"D4",X"92",X"D5",X"E9",X"D6",X"C9",X"D8",X"FA",X"DA",X"60",X"DD",
		X"DE",X"DF",X"6D",X"E2",X"F8",X"E4",X"7F",X"E7",X"FD",X"E9",X"6F",X"EC",X"CD",X"EE",X"1F",X"F1",
		X"5D",X"F3",X"8B",X"F5",X"A7",X"F7",X"B2",X"F9",X"AA",X"FB",X"96",X"FD",X"6D",X"FF",X"36",X"01",
		X"EF",X"02",X"9A",X"04",X"36",X"06",X"C4",X"07",X"43",X"09",X"B8",X"0A",X"1D",X"0C",X"77",X"0D",
		X"C3",X"0E",X"06",X"10",X"3B",X"11",X"68",X"12",X"87",X"13",X"9D",X"14",X"A8",X"15",X"A9",X"16",
		X"A3",X"17",X"90",X"18",X"77",X"19",X"57",X"1A",X"2A",X"1B",X"F8",X"1B",X"BB",X"1C",X"79",X"1D",
		X"2F",X"1E",X"DE",X"1E",X"85",X"1F",X"26",X"20",X"C0",X"20",X"54",X"21",X"E3",X"21",X"6C",X"22",
		X"EC",X"22",X"6A",X"23",X"E0",X"23",X"53",X"24",X"BF",X"24",X"27",X"25",X"89",X"25",X"EB",X"25",
		X"42",X"26",X"9A",X"26",X"EA",X"26",X"36",X"27",X"80",X"27",X"C5",X"27",X"07",X"28",X"45",X"28",
		X"80",X"28",X"B7",X"28",X"EA",X"28",X"1D",X"29",X"49",X"29",X"75",X"29",X"9C",X"29",X"C3",X"29",
		X"E3",X"29",X"06",X"2A",X"1D",X"2A",X"44",X"2A",X"F5",X"29",X"38",X"28",X"83",X"25",X"28",X"22",
		X"6A",X"1E",X"74",X"1A",X"61",X"16",X"45",X"12",X"30",X"0E",X"27",X"0A",X"36",X"06",X"58",X"02",
		X"97",X"FE",X"F0",X"FA",X"64",X"F7",X"F4",X"F3",X"A1",X"F0",X"6A",X"ED",X"4D",X"EA",X"4A",X"E7",
		X"61",X"E4",X"92",X"E1",X"DA",X"DE",X"39",X"DC",X"B3",X"D9",X"40",X"D7",X"E4",X"D4",X"9C",X"D2",
		X"69",X"D0",X"4A",X"CE",X"3E",X"CC",X"45",X"CA",X"5D",X"C8",X"89",X"C6",X"C3",X"C4",X"10",X"C3",
		X"6B",X"C1",X"D7",X"BF",X"51",X"BE",X"D9",X"BC",X"70",X"BB",X"16",X"BA",X"C8",X"B8",X"86",X"B7",
		X"51",X"B6",X"28",X"B5",X"0A",X"B4",X"FA",X"B2",X"F3",X"B1",X"F7",X"B0",X"08",X"B0",X"20",X"AF",
		X"41",X"AE",X"6E",X"AD",X"A1",X"AC",X"E0",X"AB",X"26",X"AB",X"75",X"AA",X"CA",X"A9",X"28",X"A9",
		X"8F",X"A8",X"FD",X"A7",X"70",X"A7",X"EC",X"A6",X"6E",X"A6",X"F6",X"A5",X"84",X"A5",X"1B",X"A5",
		X"B3",X"A4",X"54",X"A4",X"FA",X"A3",X"A6",X"A3",X"56",X"A3",X"0C",X"A3",X"C5",X"A2",X"85",X"A2",
		X"47",X"A2",X"10",X"A2",X"D9",X"A1",X"AE",X"A1",X"7C",X"A1",X"5C",X"A1",X"2D",X"A1",X"DE",X"A1",
		X"F4",X"A3",X"DC",X"A6",X"58",X"AA",X"23",X"AE",X"25",X"B2",X"38",X"B6",X"55",X"BA",X"65",X"BE",
		X"69",X"C2",X"57",X"C6",X"30",X"CA",X"EB",X"CD",X"8F",X"D1",X"16",X"D5",X"85",X"D8",X"D5",X"DB",
		X"0D",X"DF",X"29",X"E2",X"2C",X"E5",X"16",X"E8",X"E9",X"EA",X"A3",X"ED",X"47",X"F0",X"D5",X"F2",
		X"4D",X"F5",X"AF",X"F7",X"FE",X"F9",X"38",X"FC",X"60",X"FE",X"73",X"00",X"77",X"02",X"69",X"04",
		X"49",X"06",X"19",X"08",X"D8",X"09",X"89",X"0B",X"2A",X"0D",X"BF",X"0E",X"44",X"10",X"BC",X"11",
		X"24",X"13",X"83",X"14",X"D2",X"15",X"19",X"17",X"51",X"18",X"80",X"19",X"A0",X"1A",X"BB",X"1B",
		X"C5",X"1C",X"CC",X"1D",X"C3",X"1E",X"B9",X"1F",X"99",X"20",X"83",X"21",X"B5",X"21",X"76",X"20",
		X"4E",X"1E",X"87",X"1B",X"64",X"18",X"07",X"15",X"8F",X"11",X"0B",X"0E",X"8A",X"0A",X"13",X"07",
		X"AB",X"03",X"58",X"00",X"1B",X"FD",X"F5",X"F9",X"E6",X"F6",X"F0",X"F3",X"11",X"F1",X"4C",X"EE",
		X"9B",X"EB",X"06",X"E9",X"81",X"E6",X"18",X"E4",X"BC",X"E1",X"7D",X"DF",X"4B",X"DD",X"36",X"DB",
		X"1F",X"D9",X"AA",X"D7",X"B4",X"D7",X"BA",X"D8",X"6E",X"DA",X"8C",X"DC",X"F2",X"DE",X"7C",X"E1",
		X"1C",X"E4",X"C0",X"E6",X"65",X"E9",X"FF",X"EB",X"8D",X"EE",X"0B",X"F1",X"7A",X"F3",X"D6",X"F5",
		X"20",X"F8",X"58",X"FA",X"81",X"FC",X"94",X"FE",X"97",X"00",X"89",X"02",X"6C",X"04",X"3C",X"06",
		X"FE",X"07",X"B0",X"09",X"55",X"0B",X"E7",X"0C",X"66",X"0E",X"BE",X"0E",X"C2",X"0D",X"FD",X"0B",
		X"A8",X"09",X"02",X"07",X"25",X"04",X"33",X"01",X"34",X"FE",X"39",X"FB",X"42",X"F8",X"5F",X"F5",
		X"88",X"F2",X"C4",X"EF",X"16",X"ED",X"7B",X"EA",X"F5",X"E7",X"86",X"E5",X"29",X"E3",X"E1",X"E0",
		X"AC",X"DE",X"8A",X"DC",X"7D",X"DA",X"80",X"D8",X"97",X"D6",X"BC",X"D4",X"F7",X"D2",X"35",X"D1",
		X"E9",X"CF",X"13",X"D0",X"4D",X"D1",X"38",X"D3",X"94",X"D5",X"37",X"D8",X"00",X"DB",X"E0",X"DD",
		X"C2",X"E0",X"A1",X"E3",X"7A",X"E6",X"45",X"E9",X"FA",X"EB",X"A2",X"EE",X"34",X"F1",X"B4",X"F3",
		X"1F",X"F6",X"76",X"F8",X"BC",X"FA",X"EE",X"FC",X"0D",X"FF",X"1B",X"01",X"15",X"03",X"00",X"05",
		X"DC",X"06",X"A4",X"08",X"5E",X"0A",X"08",X"0C",X"A4",X"0D",X"33",X"0F",X"B2",X"10",X"25",X"12",
		X"8B",X"13",X"E2",X"14",X"2F",X"16",X"70",X"17",X"A4",X"18",X"CE",X"19",X"ED",X"1A",X"00",X"1C",
		X"0A",X"1D",X"0B",X"1E",X"01",X"1F",X"EE",X"1F",X"D3",X"20",X"AE",X"21",X"81",X"22",X"4C",X"23",
		X"0E",X"24",X"C9",X"24",X"7D",X"25",X"28",X"26",X"CE",X"26",X"6C",X"27",X"03",X"28",X"95",X"28",
		X"1F",X"29",X"A5",X"29",X"25",X"2A",X"9D",X"2A",X"11",X"2B",X"80",X"2B",X"EB",X"2B",X"4E",X"2C",
		X"AE",X"2C",X"09",X"2D",X"60",X"2D",X"B2",X"2D",X"00",X"2E",X"4A",X"2E",X"90",X"2E",X"D2",X"2E",
		X"10",X"2F",X"4A",X"2F",X"82",X"2F",X"B6",X"2F",X"E5",X"2F",X"12",X"30",X"3D",X"30",X"65",X"30",
		X"88",X"30",X"A9",X"30",X"C8",X"30",X"E4",X"30",X"FE",X"30",X"16",X"31",X"29",X"31",X"3C",X"31",
		X"4B",X"31",X"59",X"31",X"65",X"31",X"6F",X"31",X"77",X"31",X"7D",X"31",X"82",X"31",X"83",X"31",
		X"84",X"31",X"84",X"31",X"7F",X"31",X"7D",X"31",X"78",X"31",X"70",X"31",X"66",X"31",X"5E",X"31",
		X"53",X"31",X"46",X"31",X"38",X"31",X"29",X"31",X"19",X"31",X"0C",X"31",X"D7",X"30",X"5C",X"2F",
		X"B3",X"2C",X"5D",X"29",X"91",X"25",X"82",X"21",X"4F",X"1D",X"15",X"19",X"D8",X"14",X"AC",X"10",
		X"91",X"0C",X"8F",X"08",X"A6",X"04",X"DB",X"00",X"2A",X"FD",X"99",X"F9",X"23",X"F6",X"CB",X"F2",
		X"8A",X"EF",X"6A",X"EC",X"62",X"E9",X"73",X"E6",X"9E",X"E3",X"E3",X"E0",X"3E",X"DE",X"B2",X"DB",
		X"3A",X"D9",X"DB",X"D6",X"91",X"D4",X"59",X"D2",X"37",X"D0",X"28",X"CE",X"2A",X"CC",X"40",X"CA",
		X"65",X"C8",X"9F",X"C6",X"E7",X"C4",X"41",X"C3",X"A8",X"C1",X"20",X"C0",X"A6",X"BE",X"3A",X"BD",
		X"DC",X"BB",X"8C",X"BA",X"49",X"B9",X"12",X"B8",X"E7",X"B6",X"C8",X"B5",X"B5",X"B4",X"AB",X"B3",
		X"AD",X"B2",X"B9",X"B1",X"D1",X"B0",X"F0",X"AF",X"1A",X"AF",X"5C",X"AE",X"D1",X"AE",X"8C",X"B0",
		X"06",X"B3",X"09",X"B6",X"57",X"B9",X"D2",X"BC",X"60",X"C0",X"F7",X"C3",X"85",X"C7",X"08",X"CB",
		X"78",X"CE",X"D6",X"D1",X"1C",X"D5",X"4C",X"D8",X"64",X"DB",X"64",X"DE",X"4A",X"E1",X"1C",X"E4",
		X"D5",X"E6",X"79",X"E9",X"07",X"EC",X"7D",X"EE",X"E2",X"F0",X"31",X"F3",X"6D",X"F5",X"97",X"F7",
		X"AE",X"F9",X"B1",X"FB",X"A4",X"FD",X"86",X"FF",X"57",X"01",X"1B",X"03",X"CE",X"04",X"73",X"06",
		X"08",X"08",X"8F",X"09",X"0A",X"0B",X"77",X"0C",X"D6",X"0D",X"2C",X"0F",X"74",X"10",X"AE",X"11",
		X"E1",X"12",X"08",X"14",X"23",X"15",X"32",X"16",X"3B",X"17",X"39",X"18",X"2C",X"19",X"18",X"1A",
		X"F9",X"1A",X"D5",X"1B",X"A5",X"1C",X"6F",X"1D",X"30",X"1E",X"EB",X"1E",X"9E",X"1F",X"49",X"20",
		X"EE",X"20",X"8D",X"21",X"24",X"22",X"B4",X"22",X"41",X"23",X"C7",X"23",X"47",X"24",X"C2",X"24",
		X"39",X"25",X"A7",X"25",X"11",X"26",X"78",X"26",X"D9",X"26",X"36",X"27",X"8E",X"27",X"E2",X"27",
		X"32",X"28",X"7D",X"28",X"C5",X"28",X"0A",X"29",X"4A",X"29",X"87",X"29",X"C0",X"29",X"F6",X"29",
		X"29",X"2A",X"5A",X"2A",X"87",X"2A",X"AF",X"2A",X"D7",X"2A",X"FB",X"2A",X"1E",X"2B",X"3D",X"2B",
		X"5A",X"2B",X"74",X"2B",X"8B",X"2B",X"A0",X"2B",X"B5",X"2B",X"C6",X"2B",X"D6",X"2B",X"E1",X"2B",
		X"EE",X"2B",X"F6",X"2B",X"00",X"2C",X"05",X"2C",X"09",X"2C",X"0C",X"2C",X"0C",X"2C",X"0C",X"2C",
		X"0A",X"2C",X"06",X"2C",X"02",X"2C",X"FA",X"2B",X"F5",X"2B",X"ED",X"2B",X"E3",X"2B",X"D6",X"2B",
		X"CB",X"2B",X"BD",X"2B",X"B0",X"2B",X"A0",X"2B",X"91",X"2B",X"7F",X"2B",X"6D",X"2B",X"5B",X"2B",
		X"47",X"2B",X"32",X"2B",X"1D",X"2B",X"07",X"2B",X"F2",X"2A",X"D8",X"2A",X"C1",X"2A",X"A8",X"2A",
		X"8E",X"2A",X"76",X"2A",X"5A",X"2A",X"3F",X"2A",X"24",X"2A",X"05",X"2A",X"EE",X"29",X"A2",X"29",
		X"05",X"28",X"48",X"25",X"DD",X"21",X"02",X"1E",X"E8",X"19",X"AD",X"15",X"68",X"11",X"27",X"0D",
		X"F5",X"08",X"D6",X"04",X"D1",X"00",X"E4",X"FC",X"14",X"F9",X"64",X"F5",X"CC",X"F1",X"55",X"EE",
		X"F9",X"EA",X"B9",X"E7",X"95",X"E4",X"8F",X"E1",X"9E",X"DE",X"CB",X"DB",X"0D",X"D9",X"6B",X"D6",
		X"DB",X"D3",X"6A",X"D1",X"FF",X"CE",X"61",X"CD",X"41",X"CD",X"0C",X"CE",X"85",X"CF",X"64",X"D1",
		X"88",X"D3",X"D0",X"D5",X"32",X"D8",X"97",X"DA",X"FB",X"DC",X"58",X"DF",X"AE",X"E1",X"F2",X"E3",
		X"2B",X"E6",X"54",X"E8",X"6E",X"EA",X"73",X"EC",X"6D",X"EE",X"55",X"F0",X"2E",X"F2",X"F7",X"F3",
		X"B3",X"F5",X"5E",X"F7",X"FB",X"F8",X"8A",X"FA",X"0E",X"FC",X"82",X"FD",X"EB",X"FE",X"48",X"00",
		X"99",X"01",X"DE",X"02",X"18",X"04",X"47",X"05",X"6A",X"06",X"86",X"07",X"95",X"08",X"9E",X"09",
		X"99",X"0A",X"90",X"0B",X"7B",X"0C",X"60",X"0D",X"3A",X"0E",X"0E",X"0F",X"D9",X"0F",X"9E",X"10",
		X"57",X"11",X"10",X"12",X"BD",X"12",X"66",X"13",X"07",X"14",X"A5",X"14",X"36",X"15",X"CD",X"15",
		X"4F",X"16",X"E1",X"16",X"DE",X"16",X"6A",X"15",X"06",X"13",X"FE",X"0F",X"98",X"0C",X"F6",X"08",
		X"3B",X"05",X"73",X"01",X"B2",X"FD",X"FB",X"F9",X"57",X"F6",X"C8",X"F2",X"52",X"EF",X"F5",X"EB",
		X"B1",X"E8",X"88",X"E5",X"7A",X"E2",X"85",X"DF",X"A7",X"DC",X"E6",X"D9",X"38",X"D7",X"A6",X"D4",
		X"25",X"D2",X"C1",X"CF",X"6C",X"CD",X"36",X"CB",X"02",X"C9",X"51",X"C7",X"1A",X"C7",X"F2",X"C7",
		X"81",X"C9",X"80",X"CB",X"C9",X"CD",X"3E",X"D0",X"C6",X"D2",X"5A",X"D5",X"EC",X"D7",X"78",X"DA",
		X"F8",X"DC",X"6A",X"DF",X"CD",X"E1",X"1F",X"E4",X"60",X"E6",X"90",X"E8",X"B0",X"EA",X"BE",X"EC",
		X"B9",X"EE",X"A6",X"F0",X"83",X"F2",X"50",X"F4",X"0D",X"F6",X"BB",X"F7",X"5D",X"F9",X"EF",X"FA",
		X"75",X"FC",X"ED",X"FD",X"58",X"FF",X"B7",X"00",X"0B",X"02",X"50",X"03",X"8E",X"04",X"BF",X"05",
		X"E4",X"06",X"02",X"08",X"13",X"09",X"1D",X"0A",X"1E",X"0B",X"14",X"0C",X"00",X"0D",X"E6",X"0D",
		X"C3",X"0E",X"97",X"0F",X"63",X"10",X"2A",X"11",X"E8",X"11",X"9E",X"12",X"4F",X"13",X"F8",X"13",
		X"9A",X"14",X"39",X"15",X"CE",X"15",X"5F",X"16",X"EB",X"16",X"6F",X"17",X"EF",X"17",X"6B",X"18",
		X"E1",X"18",X"51",X"19",X"BD",X"19",X"26",X"1A",X"8A",X"1A",X"E9",X"1A",X"42",X"1B",X"9B",X"1B",
		X"EC",X"1B",X"3B",X"1C",X"86",X"1C",X"CD",X"1C",X"13",X"1D",X"54",X"1D",X"93",X"1D",X"CD",X"1D",
		X"04",X"1E",X"39",X"1E",X"6B",X"1E",X"9A",X"1E",X"C6",X"1E",X"EF",X"1E",X"17",X"1F",X"3E",X"1F",
		X"5F",X"1F",X"7D",X"1F",X"9B",X"1F",X"B8",X"1F",X"D1",X"1F",X"E8",X"1F",X"FF",X"1F",X"13",X"20",
		X"24",X"20",X"35",X"20",X"43",X"20",X"4F",X"20",X"5C",X"20",X"66",X"20",X"6E",X"20",X"74",X"20",
		X"7A",X"20",X"7E",X"20",X"80",X"20",X"82",X"20",X"84",X"20",X"83",X"20",X"80",X"20",X"7C",X"20",
		X"79",X"20",X"73",X"20",X"71",X"20",X"42",X"20",X"C9",X"1E",X"2A",X"1C",X"DA",X"18",X"15",X"15",
		X"12",X"11",X"EC",X"0C",X"BA",X"08",X"8B",X"04",X"6B",X"00",X"5D",X"FC",X"68",X"F8",X"8B",X"F4",
		X"CB",X"F0",X"29",X"ED",X"A2",X"E9",X"38",X"E6",X"EA",X"E2",X"BB",X"DF",X"A4",X"DC",X"AB",X"D9",
		X"C7",X"D6",X"03",X"D4",X"50",X"D1",X"BA",X"CE",X"36",X"CC",X"D4",X"C9",X"73",X"C7",X"D2",X"C5",
		X"B2",X"C5",X"84",X"C6",X"04",X"C8",X"E9",X"C9",X"18",X"CC",X"6B",X"CE",X"D6",X"D0",X"46",X"D3",
		X"B8",X"D5",X"20",X"D8",X"80",X"DA",X"D0",X"DC",X"13",X"DF",X"46",X"E1",X"69",X"E3",X"7D",X"E5",
		X"80",X"E7",X"71",X"E9",X"55",X"EB",X"28",X"ED",X"ED",X"EE",X"A1",X"F0",X"4A",X"F2",X"E2",X"F3",
		X"6F",X"F5",X"EE",X"F6",X"4F",X"F8",X"72",X"F8",X"51",X"F7",X"6E",X"F5",X"02",X"F3",X"49",X"F0",
		X"5D",X"ED",X"5D",X"EA",X"53",X"E7",X"4D",X"E4",X"51",X"E1",X"64",X"DE",X"89",X"DB",X"C2",X"D8",
		X"10",X"D6",X"74",X"D3",X"E9",X"D0",X"79",X"CE",X"1D",X"CC",X"D5",X"C9",X"A1",X"C7",X"82",X"C5",
		X"74",X"C3",X"7D",X"C1",X"95",X"BF",X"C0",X"BD",X"FB",X"BB",X"48",X"BA",X"A3",X"B8",X"11",X"B7",
		X"8D",X"B5",X"17",X"B4",X"AF",X"B2",X"57",X"B1",X"0B",X"B0",X"CD",X"AE",X"9A",X"AD",X"77",X"AC",
		X"5B",X"AB",X"4E",X"AA",X"4A",X"A9",X"52",X"A8",X"65",X"A7",X"80",X"A6",X"A8",X"A5",X"D8",X"A4",
		X"11",X"A4",X"52",X"A3",X"A0",X"A2",X"F1",X"A1",X"4E",X"A1",X"AF",X"A0",X"1C",X"A0",X"8B",X"9F",
		X"0A",X"9F",X"8D",X"9E",X"26",X"9F",X"12",X"A1",X"C5",X"A3",X"03",X"A7",X"8D",X"AA",X"4A",X"AE",
		X"17",X"B2",X"ED",X"B5",X"BA",X"B9",X"7A",X"BD",X"28",X"C1",X"BF",X"C4",X"3F",X"C8",X"A8",X"CB",
		X"F5",X"CE",X"2A",X"D2",X"46",X"D5",X"49",X"D8",X"34",X"DB",X"07",X"DE",X"C4",X"E0",X"6A",X"E3",
		X"FB",X"E5",X"74",X"E8",X"DD",X"EA",X"29",X"ED",X"71",X"EF",X"4C",X"F1",X"AE",X"F1",X"FC",X"F0",
		X"90",X"EF",X"B0",X"ED",X"83",X"EB",X"2D",X"E9",X"BD",X"E6",X"47",X"E4",X"CE",X"E1",X"61",X"DF",
		X"FD",X"DC",X"A9",X"DA",X"62",X"D8",X"2E",X"D6",X"0C",X"D4",X"FB",X"D1",X"FA",X"CF",X"0D",X"CE",
		X"2F",X"CC",X"67",X"CA",X"A8",X"C8",X"FE",X"C6",X"61",X"C5",X"D5",X"C3",X"54",X"C2",X"EA",X"C0",
		X"82",X"BF",X"0D",X"BF",X"05",X"C0",X"D2",X"C1",X"3B",X"C4",X"FA",X"C6",X"F6",X"C9",X"0A",X"CD",
		X"2D",X"D0",X"4E",X"D3",X"69",X"D6",X"76",X"D9",X"74",X"DC",X"5C",X"DF",X"33",X"E2",X"F2",X"E4",
		X"9E",X"E7",X"36",X"EA",X"B6",X"EC",X"24",X"EF",X"7D",X"F1",X"C4",X"F3",X"F7",X"F5",X"17",X"F8",
		X"25",X"FA",X"24",X"FC",X"0E",X"FE",X"EE",X"FF",X"86",X"01",X"B9",X"01",X"C1",X"00",X"13",X"FF",
		X"E6",X"FC",X"6D",X"FA",X"C5",X"F7",X"0A",X"F5",X"44",X"F2",X"82",X"EF",X"C6",X"EC",X"1C",X"EA",
		X"7F",X"E7",X"F5",X"E4",X"7A",X"E2",X"17",X"E0",X"C6",X"DD",X"88",X"DB",X"5F",X"D9",X"46",X"D7",
		X"41",X"D5",X"4D",X"D3",X"6D",X"D1",X"9C",X"CF",X"DC",X"CD",X"2D",X"CC",X"8D",X"CA",X"FD",X"C8",
		X"7A",X"C7",X"06",X"C6",X"A0",X"C4",X"48",X"C3",X"FC",X"C1",X"BD",X"C0",X"89",X"BF",X"64",X"BE",
		X"47",X"BD",X"38",X"BC",X"31",X"BB",X"38",X"BA",X"47",X"B9",X"61",X"B8",X"83",X"B7",X"B0",X"B6",
		X"E5",X"B5",X"22",X"B5",X"6A",X"B4",X"B8",X"B3",X"0D",X"B3",X"6C",X"B2",X"D1",X"B1",X"3D",X"B1",
		X"B1",X"B0",X"2B",X"B0",X"AC",X"AF",X"34",X"AF",X"C1",X"AE",X"54",X"AE",X"ED",X"AD",X"8C",X"AD",
		X"30",X"AD",X"DA",X"AC",X"87",X"AC",X"3C",X"AC",X"F5",X"AB",X"B0",X"AB",X"71",X"AB",X"36",X"AB",
		X"01",X"AB",X"CF",X"AA",X"A0",X"AA",X"75",X"AA",X"50",X"AA",X"2C",X"AA",X"0C",X"AA",X"F1",X"A9",
		X"D7",X"A9",X"C0",X"A9",X"AE",X"A9",X"9F",X"A9",X"91",X"A9",X"86",X"A9",X"7E",X"A9",X"79",X"A9",
		X"77",X"A9",X"76",X"A9",X"77",X"A9",X"7B",X"A9",X"83",X"A9",X"8B",X"A9",X"95",X"A9",X"A2",X"A9",
		X"B1",X"A9",X"C1",X"A9",X"D3",X"A9",X"E8",X"A9",X"FC",X"A9",X"13",X"AA",X"2B",X"AA",X"46",X"AA",
		X"60",X"AA",X"7E",X"AA",X"9C",X"AA",X"BB",X"AA",X"DB",X"AA",X"FD",X"AA",X"1F",X"AB",X"46",X"AB",
		X"68",X"AB",X"90",X"AB",X"C1",X"AB",X"12",X"AD",X"A8",X"AF",X"FA",X"B2",X"CE",X"B6",X"E8",X"BA",
		X"2B",X"BF",X"7B",X"C3",X"CD",X"C7",X"11",X"CC",X"44",X"D0",X"5E",X"D4",X"61",X"D8",X"45",X"DC",
		X"0E",X"E0",X"BA",X"E3",X"49",X"E7",X"BA",X"EA",X"12",X"EE",X"4D",X"F1",X"6D",X"F4",X"74",X"F7",
		X"5F",X"FA",X"33",X"FD",X"EE",X"FF",X"92",X"02",X"21",X"05",X"97",X"07",X"FB",X"09",X"47",X"0C",
		X"82",X"0E",X"A7",X"10",X"BC",X"12",X"BB",X"14",X"A9",X"16",X"88",X"18",X"54",X"1A",X"11",X"1C",
		X"BE",X"1D",X"5C",X"1F",X"EC",X"20",X"6B",X"22",X"DF",X"23",X"44",X"25",X"9F",X"26",X"E8",X"27",
		X"29",X"29",X"5C",X"2A",X"85",X"2B",X"A0",X"2C",X"B3",X"2D",X"B8",X"2E",X"B9",X"2F",X"A8",X"30",
		X"9B",X"31",X"33",X"32",X"63",X"31",X"7E",X"2F",X"EA",X"2C",X"E4",X"29",X"9C",X"26",X"2C",X"23",
		X"AF",X"1F",X"2F",X"1C",X"B8",X"18",X"4E",X"15",X"F7",X"11",X"B5",X"0E",X"88",X"0B",X"75",X"08",
		X"79",X"05",X"94",X"02",X"C6",X"FF",X"10",X"FD",X"6F",X"FA",X"E6",X"F7",X"72",X"F5",X"12",X"F3",
		X"C9",X"F0",X"91",X"EE",X"6E",X"EC",X"5C",X"EA",X"5D",X"E8",X"71",X"E6",X"94",X"E4",X"C8",X"E2",
		X"0C",X"E1",X"60",X"DF",X"C4",X"DD",X"35",X"DC",X"B7",X"DA",X"42",X"D9",X"DF",X"D7",X"86",X"D6",
		X"3A",X"D5",X"FB",X"D3",X"C9",X"D2",X"A0",X"D1",X"83",X"D0",X"70",X"CF",X"6A",X"CE",X"6B",X"CD",
		X"78",X"CC",X"8D",X"CB",X"AC",X"CA",X"D2",X"C9",X"04",X"C9",X"3D",X"C8",X"7E",X"C7",X"C6",X"C6",
		X"18",X"C6",X"6F",X"C5",X"CE",X"C4",X"33",X"C4",X"A1",X"C3",X"13",X"C3",X"8D",X"C2",X"0E",X"C2",
		X"94",X"C1",X"1D",X"C1",X"B1",X"C0",X"45",X"C0",X"E1",X"BF",X"81",X"BF",X"27",X"BF",X"D0",X"BE",
		X"82",X"BE",X"33",X"BE",X"EE",X"BD",X"A7",X"BD",X"69",X"BD",X"2B",X"BD",X"F4",X"BC",X"BD",X"BC",
		X"92",X"BC",X"5E",X"BC",X"3C",X"BC",X"07",X"BC",X"89",X"BC",X"76",X"BE",X"45",X"C1",X"B0",X"C4",
		X"6F",X"C8",X"67",X"CC",X"74",X"D0",X"89",X"D4",X"96",X"D8",X"95",X"DC",X"80",X"E0",X"53",X"E4",
		X"0A",X"E8",X"AB",X"EB",X"2D",X"EF",X"95",X"F2",X"E1",X"F5",X"10",X"F9",X"28",X"FC",X"24",X"FF",
		X"08",X"02",X"D4",X"04",X"86",X"07",X"22",X"0A",X"A6",X"0C",X"17",X"0F",X"72",X"11",X"A2",X"13",
		X"89",X"14",X"27",X"14",X"FF",X"12",X"47",X"11",X"3C",X"0F",X"F9",X"0C",X"9C",X"0A",X"2F",X"08",
		X"C0",X"05",X"54",X"03",X"F5",X"00",X"A0",X"FE",X"5A",X"FC",X"24",X"FA",X"FF",X"F7",X"EA",X"F5",
		X"E7",X"F3",X"F2",X"F1",X"0F",X"F0",X"3C",X"EE",X"7A",X"EC",X"C4",X"EA",X"21",X"E9",X"8B",X"E7",
		X"03",X"E6",X"89",X"E4",X"1B",X"E3",X"BA",X"E1",X"67",X"E0",X"1F",X"DF",X"E4",X"DD",X"B1",X"DC",
		X"8E",X"DB",X"73",X"DA",X"63",X"D9",X"5D",X"D8",X"61",X"D7",X"6E",X"D6",X"85",X"D5",X"A4",X"D4",
		X"CD",X"D3",X"FE",X"D2",X"35",X"D2",X"75",X"D1",X"BF",X"D0",X"0D",X"D0",X"65",X"CF",X"C3",X"CE",
		X"27",X"CE",X"92",X"CD",X"03",X"CD",X"7C",X"CC",X"F8",X"CB",X"7E",X"CB",X"0C",X"CB",X"B3",X"CB",
		X"AB",X"CD",X"64",X"D0",X"A8",X"D3",X"34",X"D7",X"F1",X"DA",X"BF",X"DE",X"93",X"E2",X"5E",X"E6",
		X"1B",X"EA",X"C1",X"ED",X"55",X"F1",X"CD",X"F4",X"2C",X"F8",X"70",X"FB",X"9C",X"FE",X"AD",X"01",
		X"A7",X"04",X"85",X"07",X"4D",X"0A",X"FB",X"0C",X"93",X"0F",X"14",X"12",X"81",X"14",X"D6",X"16",
		X"19",X"19",X"46",X"1B",X"60",X"1D",X"68",X"1F",X"5E",X"21",X"41",X"23",X"13",X"25",X"D6",X"26",
		X"88",X"28",X"2A",X"2A",X"BD",X"2B",X"40",X"2D",X"B6",X"2E",X"1E",X"30",X"7A",X"31",X"C6",X"32",
		X"08",X"34",X"3D",X"35",X"66",X"36",X"83",X"37",X"96",X"38",X"9E",X"39",X"9C",X"3A",X"8D",X"3B",
		X"76",X"3C",X"55",X"3D",X"2C",X"3E",X"FA",X"3E",X"BE",X"3F",X"7B",X"40",X"30",X"41",X"DB",X"41",
		X"80",X"42",X"1F",X"43",X"B2",X"43",X"43",X"44",X"CB",X"44",X"4C",X"45",X"C8",X"45",X"3F",X"46",
		X"AC",X"46",X"17",X"47",X"7B",X"47",X"DA",X"47",X"32",X"48",X"88",X"48",X"D7",X"48",X"22",X"49",
		X"69",X"49",X"A9",X"49",X"E6",X"49",X"1F",X"4A",X"54",X"4A",X"86",X"4A",X"B3",X"4A",X"DD",X"4A",
		X"02",X"4B",X"26",X"4B",X"44",X"4B",X"61",X"4B",X"79",X"4B",X"90",X"4B",X"A3",X"4B",X"B1",X"4B",
		X"BF",X"4B",X"C9",X"4B",X"D4",X"4B",X"D8",X"4B",X"DC",X"4B",X"DC",X"4B",X"DC",X"4B",X"D8",X"4B",
		X"D3",X"4B",X"CC",X"4B",X"C1",X"4B",X"B5",X"4B",X"A8",X"4B",X"98",X"4B",X"8A",X"4B",X"74",X"4B",
		X"63",X"4B",X"4A",X"4B",X"37",X"4B",X"19",X"4B",X"0B",X"4B",X"34",X"4A",X"F5",X"47",X"E1",X"44",
		X"36",X"41",X"39",X"3D",X"09",X"39",X"C6",X"34",X"7D",X"30",X"40",X"2C",X"10",X"28",X"FB",X"23",
		X"F7",X"1F",X"17",X"1C",X"4C",X"18",X"A0",X"14",X"10",X"11",X"A0",X"0D",X"48",X"0A",X"0C",X"07",
		X"EB",X"03",X"E7",X"00",X"FA",X"FD",X"26",X"FB",X"6A",X"F8",X"C7",X"F5",X"39",X"F3",X"C0",X"F0",
		X"5E",X"EE",X"10",X"EC",X"D6",X"E9",X"B0",X"E7",X"9E",X"E5",X"9D",X"E3",X"AF",X"E1",X"CF",X"DF",
		X"03",X"DE",X"46",X"DC",X"9A",X"DA",X"FD",X"D8",X"6D",X"D7",X"ED",X"D5",X"7B",X"D4",X"15",X"D3",
		X"BE",X"D1",X"71",X"D0",X"33",X"CF",X"00",X"CE",X"D8",X"CC",X"BC",X"CB",X"AB",X"CA",X"A4",X"C9",
		X"A7",X"C8",X"B3",X"C7",X"CB",X"C6",X"E9",X"C5",X"12",X"C5",X"46",X"C4",X"80",X"C3",X"C2",X"C2",
		X"0C",X"C2",X"5F",X"C1",X"B7",X"C0",X"19",X"C0",X"80",X"BF",X"EF",X"BE",X"64",X"BE",X"DF",X"BD",
		X"62",X"BD",X"E8",X"BC",X"77",X"BC",X"09",X"BC",X"A4",X"BB",X"40",X"BB",X"E4",X"BA",X"8C",X"BA",
		X"37",X"BA",X"EA",X"B9",X"9F",X"B9",X"5A",X"B9",X"19",X"B9",X"DA",X"B8",X"A2",X"B8",X"6B",X"B8",
		X"3A",X"B8",X"0C",X"B8",X"E3",X"B7",X"BA",X"B7",X"96",X"B7",X"77",X"B7",X"57",X"B7",X"3C",X"B7",
		X"25",X"B7",X"0F",X"B7",X"FE",X"B6",X"ED",X"B6",X"DF",X"B6",X"D4",X"B6",X"CB",X"B6",X"C6",X"B6",
		X"C1",X"B6",X"BF",X"B6",X"BF",X"B6",X"C1",X"B6",X"C6",X"B6",X"CC",X"B6",X"D2",X"B6",X"DD",X"B6",
		X"E6",X"B6",X"F5",X"B6",X"02",X"B7",X"12",X"B7",X"24",X"B7",X"36",X"B7",X"4A",X"B7",X"5F",X"B7",
		X"76",X"B7",X"8D",X"B7",X"A9",X"B7",X"C1",X"B7",X"DD",X"B7",X"FA",X"B7",X"17",X"B8",X"35",X"B8",
		X"54",X"B8",X"74",X"B8",X"95",X"B8",X"B8",X"B8",X"DB",X"B8",X"FF",X"B8",X"22",X"B9",X"48",X"B9",
		X"6E",X"B9",X"95",X"B9",X"BB",X"B9",X"E3",X"B9",X"0C",X"BA",X"35",X"BA",X"5F",X"BA",X"8A",X"BA",
		X"B2",X"BA",X"DE",X"BA",X"0A",X"BB",X"36",X"BB",X"61",X"BB",X"90",X"BB",X"BB",X"BB",X"EA",X"BB",
		X"18",X"BC",X"48",X"BC",X"75",X"BC",X"A5",X"BC",X"D4",X"BC",X"04",X"BD",X"32",X"BD",X"63",X"BD",
		X"92",X"BD",X"C3",X"BD",X"F5",X"BD",X"25",X"BE",X"57",X"BE",X"88",X"BE",X"BA",X"BE",X"EC",X"BE",
		X"1D",X"BF",X"50",X"BF",X"81",X"BF",X"B4",X"BF",X"E8",X"BF",X"19",X"C0",X"4C",X"C0",X"7F",X"C0",
		X"B1",X"C0",X"E4",X"C0",X"16",X"C1",X"4B",X"C1",X"7C",X"C1",X"AF",X"C1",X"E3",X"C1",X"18",X"C2",
		X"4A",X"C2",X"7E",X"C2",X"AF",X"C2",X"E4",X"C2",X"18",X"C3",X"4B",X"C3",X"7C",X"C3",X"B1",X"C3",
		X"E3",X"C3",X"18",X"C4",X"49",X"C4",X"7F",X"C4",X"AC",X"C4",X"10",X"C5",X"C4",X"C6",X"96",X"C9",
		X"16",X"CD",X"05",X"D1",X"32",X"D5",X"80",X"D9",X"D7",X"DD",X"2A",X"E2",X"70",X"E6",X"A0",X"EA",
		X"B6",X"EE",X"B4",X"F2",X"94",X"F6",X"56",X"FA",X"FA",X"FD",X"82",X"01",X"EC",X"04",X"3A",X"08",
		X"6B",X"0B",X"84",X"0E",X"7F",X"11",X"63",X"14",X"2B",X"17",X"DD",X"19",X"77",X"1C",X"FA",X"1E",
		X"66",X"21",X"BC",X"23",X"FD",X"25",X"2A",X"28",X"45",X"2A",X"4C",X"2C",X"40",X"2E",X"21",X"30",
		X"F2",X"31",X"B1",X"33",X"60",X"35",X"FF",X"36",X"91",X"38",X"13",X"3A",X"84",X"3B",X"E9",X"3C",
		X"3E",X"3E",X"8B",X"3F",X"C6",X"40",X"F7",X"41",X"1D",X"43",X"35",X"44",X"42",X"45",X"46",X"46",
		X"3E",X"47",X"2C",X"48",X"0F",X"49",X"EB",X"49",X"BB",X"4A",X"83",X"4B",X"40",X"4C",X"F8",X"4C",
		X"A5",X"4D",X"4C",X"4E",X"EA",X"4E",X"82",X"4F",X"11",X"50",X"9A",X"50",X"1B",X"51",X"98",X"51",
		X"0D",X"52",X"7B",X"52",X"E1",X"52",X"45",X"53",X"A0",X"53",X"FB",X"53",X"4C",X"54",X"9B",X"54",
		X"E1",X"54",X"27",X"55",X"62",X"55",X"9F",X"55",X"D1",X"55",X"07",X"56",X"2D",X"56",X"65",X"56",
		X"08",X"56",X"3B",X"54",X"7F",X"51",X"20",X"4E",X"68",X"4A",X"73",X"46",X"66",X"42",X"4E",X"3E",
		X"3D",X"3A",X"38",X"36",X"46",X"32",X"6D",X"2E",X"AD",X"2A",X"05",X"27",X"7A",X"23",X"08",X"20",
		X"B3",X"1C",X"77",X"19",X"57",X"16",X"50",X"13",X"62",X"10",X"8C",X"0D",X"CF",X"0A",X"25",X"08",
		X"96",X"05",X"18",X"03",X"B5",X"00",X"6B",X"FE",X"4F",X"FD",X"8B",X"FD",X"98",X"FE",X"39",X"00",
		X"30",X"02",X"63",X"04",X"B3",X"06",X"13",X"09",X"75",X"0B",X"D5",X"0D",X"2A",X"10",X"73",X"12",
		X"AE",X"14",X"D7",X"16",X"F2",X"18",X"FC",X"1A",X"F2",X"1C",X"DB",X"1E",X"B3",X"20",X"79",X"22",
		X"31",X"24",X"D7",X"25",X"70",X"27",X"F8",X"28",X"75",X"2A",X"DE",X"2B",X"49",X"2D",X"3E",X"2E",
		X"BF",X"2D",X"37",X"2C",X"FB",X"29",X"55",X"27",X"68",X"24",X"58",X"21",X"35",X"1E",X"0E",X"1B",
		X"ED",X"17",X"D8",X"14",X"D2",X"11",X"E2",X"0E",X"02",X"0C",X"39",X"09",X"83",X"06",X"E5",X"03",
		X"59",X"01",X"E7",X"FE",X"85",X"FC",X"38",X"FA",X"FE",X"F7",X"D9",X"F5",X"C4",X"F3",X"C5",X"F1",
		X"D1",X"EF",X"F7",X"ED",X"23",X"EC",X"55",X"EB",X"F0",X"EB",X"5F",X"ED",X"69",X"EF",X"CA",X"F1",
		X"69",X"F4",X"1F",X"F7",X"E9",X"F9",X"B0",X"FC",X"72",X"FF",X"29",X"02",X"D3",X"04",X"67",X"07",
		X"EB",X"09",X"5D",X"0C",X"BC",X"0E",X"05",X"11",X"3F",X"13",X"63",X"15",X"75",X"17",X"74",X"19",
		X"62",X"1B",X"3E",X"1D",X"0D",X"1F",X"C9",X"20",X"75",X"22",X"11",X"24",X"A0",X"25",X"20",X"27",
		X"92",X"28",X"F8",X"29",X"4C",X"2B",X"9A",X"2C",X"D7",X"2D",X"0A",X"2F",X"31",X"30",X"4B",X"31",
		X"5C",X"32",X"62",X"33",X"5E",X"34",X"50",X"35",X"36",X"36",X"17",X"37",X"EC",X"37",X"B9",X"38",
		X"7D",X"39",X"3A",X"3A",X"ED",X"3A",X"9D",X"3B",X"3F",X"3C",X"E1",X"3C",X"73",X"3D",X"07",X"3E",
		X"8A",X"3E",X"19",X"3F",X"D2",X"3E",X"20",X"3D",X"96",X"3A",X"74",X"37",X"FB",X"33",X"4B",X"30",
		X"86",X"2C",X"B7",X"28",X"EF",X"24",X"33",X"21",X"8C",X"1D",X"F5",X"19",X"7A",X"16",X"17",X"13",
		X"CD",X"0F",X"9C",X"0C",X"85",X"09",X"87",X"06",X"A2",X"03",X"D5",X"00",X"21",X"FE",X"83",X"FB",
		X"F9",X"F8",X"87",X"F6",X"2B",X"F4",X"E1",X"F1",X"A7",X"EF",X"A8",X"ED",X"04",X"ED",X"98",X"ED",
		X"EE",X"EE",X"CD",X"F0",X"F7",X"F2",X"59",X"F5",X"D1",X"F7",X"57",X"FA",X"DB",X"FC",X"5D",X"FF",
		X"D1",X"01",X"39",X"04",X"90",X"06",X"D9",X"08",X"0F",X"0B",X"35",X"0D",X"46",X"0F",X"48",X"11",
		X"38",X"13",X"18",X"15",X"E6",X"16",X"A8",X"18",X"55",X"1A",X"F8",X"1B",X"87",X"1D",X"0D",X"1F",
		X"81",X"20",X"EB",X"21",X"45",X"23",X"94",X"24",X"D7",X"25",X"0D",X"27",X"38",X"28",X"57",X"29",
		X"6C",X"2A",X"77",X"2B",X"75",X"2C",X"6D",X"2D",X"58",X"2E",X"3D",X"2F",X"17",X"30",X"E9",X"30",
		X"B1",X"31",X"72",X"32",X"2D",X"33",X"DD",X"33",X"88",X"34",X"2A",X"35",X"C6",X"35",X"5A",X"36",
		X"E9",X"36",X"71",X"37",X"F3",X"37",X"6E",X"38",X"D5",X"38",X"0B",X"38",X"FE",X"35",X"37",X"33",
		X"E9",X"2F",X"55",X"2C",X"94",X"28",X"C2",X"24",X"EC",X"20",X"22",X"1D",X"64",X"19",X"BC",X"15",
		X"28",X"12",X"B0",X"0E",X"4D",X"0B",X"09",X"08",X"DA",X"04",X"C8",X"01",X"CE",X"FE",X"EE",X"FB",
		X"26",X"F9",X"73",X"F6",X"D9",X"F3",X"56",X"F1",X"E7",X"EE",X"8E",X"EC",X"49",X"EA",X"1A",X"E8",
		X"FA",X"E5",X"F1",X"E3",X"F7",X"E1",X"11",X"E0",X"3A",X"DE",X"75",X"DC",X"C0",X"DA",X"19",X"D9",
		X"83",X"D7",X"FA",X"D5",X"80",X"D4",X"14",X"D3",X"B5",X"D1",X"62",X"D0",X"1D",X"CF",X"E3",X"CD",
		X"B6",X"CC",X"93",X"CB",X"7D",X"CA",X"6F",X"C9",X"6E",X"C8",X"74",X"C7",X"88",X"C6",X"A1",X"C5",
		X"C9",X"C4",X"F3",X"C3",X"2E",X"C3",X"6C",X"C2",X"BE",X"C2",X"65",X"C4",X"D4",X"C6",X"D3",X"C9",
		X"20",X"CD",X"A2",X"D0",X"36",X"D4",X"D2",X"D7",X"68",X"DB",X"F2",X"DE",X"6A",X"E2",X"CE",X"E5",
		X"1B",X"E9",X"50",X"EC",X"6C",X"EF",X"71",X"F2",X"5D",X"F5",X"32",X"F8",X"EF",X"FA",X"95",X"FD",
		X"25",X"00",X"9C",X"02",X"03",X"05",X"52",X"07",X"91",X"09",X"B6",X"0B",X"D6",X"0D",X"8C",X"0F",
		X"CF",X"0F",X"F9",X"0E",X"6A",X"0D",X"65",X"0B",X"15",X"09",X"99",X"06",X"06",X"04",X"6B",X"01",
		X"D2",X"FE",X"40",X"FC",X"BA",X"F9",X"42",X"F7",X"DC",X"F4",X"87",X"F2",X"42",X"F0",X"10",X"EE",
		X"F2",X"EB",X"E4",X"E9",X"EA",X"E7",X"FD",X"E5",X"25",X"E4",X"5A",X"E2",X"A0",X"E0",X"F6",X"DE",
		X"5B",X"DD",X"CE",X"DB",X"50",X"DA",X"DD",X"D8",X"7B",X"D7",X"24",X"D6",X"DB",X"D4",X"9B",X"D3",
		X"6B",X"D2",X"44",X"D1",X"29",X"D0",X"17",X"CF",X"11",X"CE",X"13",X"CD",X"22",X"CC",X"38",X"CB",
		X"59",X"CA",X"80",X"C9",X"B3",X"C8",X"EC",X"C7",X"30",X"C7",X"78",X"C6",X"CC",X"C5",X"22",X"C5",
		X"85",X"C4",X"E9",X"C3",X"5B",X"C3",X"C9",X"C2",X"4D",X"C2",X"C0",X"C1",X"FC",X"C1",X"A5",X"C3",
		X"2B",X"C6",X"4D",X"C9",X"C4",X"CC",X"72",X"D0",X"3A",X"D4",X"0B",X"D8",X"D5",X"DB",X"94",X"DF",
		X"3F",X"E3",X"D6",X"E6",X"53",X"EA",X"B9",X"ED",X"03",X"F1",X"35",X"F4",X"4C",X"F7",X"4C",X"FA",
		X"32",X"FD",X"FF",X"FF",X"B5",X"02",X"52",X"05",X"DB",X"07",X"4F",X"0A",X"AC",X"0C",X"F6",X"0E",
		X"2C",X"11",X"32",X"13",X"E6",X"13",X"5A",X"13",X"08",X"12",X"2E",X"10",X"02",X"0E",X"A2",X"0B",
		X"27",X"09",X"9F",X"06",X"17",X"04",X"94",X"01",X"1D",X"FF",X"B3",X"FC",X"58",X"FA",X"0C",X"F8",
		X"D3",X"F5",X"AC",X"F3",X"94",X"F1",X"90",X"EF",X"9B",X"ED",X"B9",X"EB",X"E4",X"E9",X"24",X"E8",
		X"6E",X"E6",X"CE",X"E4",X"33",X"E3",X"B2",X"E1",X"2B",X"E0",X"48",X"DF",X"E1",X"DF",X"6A",X"E1",
		X"A1",X"E3",X"3A",X"E6",X"14",X"E9",X"0F",X"EC",X"1B",X"EF",X"2A",X"F2",X"31",X"F5",X"2C",X"F8",
		X"19",X"FB",X"F2",X"FD",X"B7",X"00",X"68",X"03",X"03",X"06",X"89",X"08",X"FC",X"0A",X"57",X"0D",
		X"A1",X"0F",X"D7",X"11",X"F9",X"13",X"06",X"16",X"08",X"18",X"F1",X"19",X"CD",X"1B",X"96",X"1D",
		X"46",X"1F",X"C5",X"1F",X"F3",X"1E",X"58",X"1D",X"2C",X"1B",X"AE",X"18",X"F9",X"15",X"2C",X"13",
		X"52",X"10",X"79",X"0D",X"A5",X"0A",X"E1",X"07",X"2A",X"05",X"87",X"02",X"F5",X"FF",X"77",X"FD",
		X"0D",X"FB",X"B5",X"F8",X"70",X"F6",X"3E",X"F4",X"20",X"F2",X"13",X"F0",X"19",X"EE",X"2D",X"EC",
		X"56",X"EA",X"8B",X"E8",X"D8",X"E6",X"23",X"E5",X"EB",X"E3",X"2C",X"E4",X"75",X"E5",X"6F",X"E7",
		X"D7",X"E9",X"85",X"EC",X"57",X"EF",X"40",X"F2",X"29",X"F5",X"11",X"F8",X"EE",X"FA",X"BC",X"FD",
		X"77",X"00",X"21",X"03",X"B8",X"05",X"39",X"08",X"A6",X"0A",X"00",X"0D",X"48",X"0F",X"7A",X"11",
		X"9A",X"13",X"A7",X"15",X"A2",X"17",X"8C",X"19",X"65",X"1B",X"2C",X"1D",X"E6",X"1E",X"8E",X"20",
		X"26",X"22",X"B2",X"23",X"2E",X"25",X"9C",X"26",X"FE",X"27",X"52",X"29",X"9A",X"2A",X"D7",X"2B",
		X"06",X"2D",X"29",X"2E",X"44",X"2F",X"51",X"30",X"58",X"31",X"50",X"32",X"42",X"33",X"28",X"34",
		X"04",X"35",X"D9",X"35",X"A5",X"36",X"68",X"37",X"23",X"38",X"D6",X"38",X"83",X"39",X"27",X"3A",
		X"C4",X"3A",X"5B",X"3B",X"EA",X"3B",X"73",X"3C",X"F4",X"3C",X"72",X"3D",X"E7",X"3D",X"59",X"3E",
		X"C2",X"3E",X"2B",X"3F",X"8A",X"3F",X"E6",X"3F",X"3C",X"40",X"8E",X"40",X"DB",X"40",X"24",X"41",
		X"68",X"41",X"A8",X"41",X"E4",X"41",X"1C",X"42",X"51",X"42",X"82",X"42",X"AE",X"42",X"D9",X"42",
		X"FF",X"42",X"23",X"43",X"42",X"43",X"5E",X"43",X"79",X"43",X"8F",X"43",X"A4",X"43",X"B5",X"43",
		X"C5",X"43",X"D0",X"43",X"DA",X"43",X"E3",X"43",X"E9",X"43",X"ED",X"43",X"EE",X"43",X"EE",X"43",
		X"EA",X"43",X"E5",X"43",X"DF",X"43",X"D8",X"43",X"CC",X"43",X"C3",X"43",X"B5",X"43",X"A6",X"43",
		X"95",X"43",X"85",X"43",X"70",X"43",X"5B",X"43",X"46",X"43",X"2F",X"43",X"16",X"43",X"FD",X"42",
		X"E2",X"42",X"C9",X"42",X"86",X"42",X"F6",X"40",X"3F",X"3E",X"DA",X"3A",X"FF",X"36",X"E7",X"32",
		X"AA",X"2E",X"64",X"2A",X"1E",X"26",X"E7",X"21",X"C1",X"1D",X"B7",X"19",X"C4",X"15",X"ED",X"11",
		X"34",X"0E",X"99",X"0A",X"19",X"07",X"B6",X"03",X"6D",X"00",X"42",X"FD",X"2F",X"FA",X"38",X"F7",
		X"5A",X"F4",X"95",X"F1",X"E6",X"EE",X"51",X"EC",X"CF",X"E9",X"66",X"E7",X"10",X"E5",X"D1",X"E2",
		X"A4",X"E0",X"8B",X"DE",X"85",X"DC",X"91",X"DA",X"AE",X"D8",X"DD",X"D6",X"1B",X"D5",X"6B",X"D3",
		X"C8",X"D1",X"37",X"D0",X"B4",X"CE",X"3F",X"CD",X"D7",X"CB",X"7D",X"CA",X"30",X"C9",X"EE",X"C7",
		X"BA",X"C6",X"91",X"C5",X"75",X"C4",X"62",X"C3",X"5C",X"C2",X"5E",X"C1",X"6A",X"C0",X"81",X"BF",
		X"A1",X"BE",X"DD",X"BD",X"52",X"BE",X"09",X"C0",X"7F",X"C2",X"79",X"C5",X"BE",X"C8",X"31",X"CC",
		X"B6",X"CF",X"46",X"D3",X"C9",X"D6",X"43",X"DA",X"A9",X"DD",X"FE",X"E0",X"38",X"E4",X"5E",X"E7",
		X"6B",X"EA",X"60",X"ED",X"40",X"F0",X"07",X"F3",X"B5",X"F5",X"50",X"F8",X"D3",X"FA",X"43",X"FD",
		X"9D",X"FF",X"E2",X"01",X"14",X"04",X"33",X"06",X"40",X"08",X"3C",X"0A",X"26",X"0C",X"FF",X"0D",
		X"C8",X"0F",X"80",X"11",X"2A",X"13",X"C6",X"14",X"52",X"16",X"D1",X"17",X"42",X"19",X"A6",X"1A",
		X"FE",X"1B",X"48",X"1D",X"87",X"1E",X"BB",X"1F",X"E3",X"20",X"FF",X"21",X"13",X"23",X"1B",X"24",
		X"19",X"25",X"0E",X"26",X"FB",X"26",X"DB",X"27",X"B9",X"28",X"87",X"29",X"52",X"2A",X"0E",X"2B",
		X"C6",X"2B",X"66",X"2B",X"B1",X"29",X"36",X"27",X"30",X"24",X"DC",X"20",X"56",X"1D",X"BD",X"19",
		X"1C",X"16",X"83",X"12",X"F4",X"0E",X"7B",X"0B",X"16",X"08",X"C8",X"04",X"92",X"01",X"75",X"FE",
		X"71",X"FB",X"83",X"F8",X"B0",X"F5",X"F5",X"F2",X"50",X"F0",X"C0",X"ED",X"49",X"EB",X"E4",X"E8",
		X"99",X"E6",X"5C",X"E4",X"3A",X"E2",X"1C",X"E0",X"6E",X"DE",X"38",X"DE",X"15",X"DF",X"AB",X"E0",
		X"B6",X"E2",X"0B",X"E5",X"8B",X"E7",X"25",X"EA",X"C1",X"EC",X"61",X"EF",X"F8",X"F1",X"83",X"F4",
		X"FE",X"F6",X"6A",X"F9",X"C5",X"FB",X"0E",X"FE",X"43",X"00",X"68",X"02",X"7B",X"04",X"7D",X"06",
		X"6D",X"08",X"4E",X"0A",X"1D",X"0C",X"E0",X"0D",X"8C",X"0F",X"31",X"11",X"C0",X"12",X"4C",X"14",
		X"E2",X"14",X"0B",X"14",X"60",X"12",X"19",X"10",X"7D",X"0D",X"A2",X"0A",X"B0",X"07",X"AD",X"04",
		X"AF",X"01",X"B4",X"FE",X"CA",X"FB",X"ED",X"F8",X"25",X"F6",X"6F",X"F3",X"D1",X"F0",X"44",X"EE",
		X"CF",X"EB",X"6B",X"E9",X"1E",X"E7",X"E4",X"E4",X"BD",X"E2",X"A8",X"E0",X"A8",X"DE",X"B8",X"DC",
		X"DB",X"DA",X"0D",X"D9",X"50",X"D7",X"A4",X"D5",X"06",X"D4",X"79",X"D2",X"F7",X"D0",X"84",X"CF",
		X"21",X"CE",X"C9",X"CC",X"7E",X"CB",X"40",X"CA",X"0E",X"C9",X"E7",X"C7",X"CC",X"C6",X"BC",X"C5",
		X"B8",X"C4",X"BC",X"C3",X"CA",X"C2",X"E2",X"C1",X"04",X"C1",X"30",X"C0",X"62",X"BF",X"A0",X"BE",
		X"E3",X"BD",X"31",X"BD",X"85",X"BC",X"E1",X"BB",X"45",X"BB",X"AE",X"BA",X"1F",X"BA",X"97",X"B9",
		X"16",X"B9",X"9B",X"B8",X"25",X"B8",X"B6",X"B7",X"4C",X"B7",X"E8",X"B6",X"88",X"B6",X"2E",X"B6",
		X"D9",X"B5",X"8A",X"B5",X"3D",X"B5",X"F8",X"B4",X"B4",X"B4",X"76",X"B4",X"3C",X"B4",X"06",X"B4",
		X"D5",X"B3",X"A5",X"B3",X"7B",X"B3",X"53",X"B3",X"2F",X"B3",X"10",X"B3",X"F0",X"B2",X"D8",X"B2",
		X"C1",X"B2",X"AB",X"B2",X"9A",X"B2",X"8B",X"B2",X"7F",X"B2",X"74",X"B2",X"6E",X"B2",X"69",X"B2",
		X"66",X"B2",X"66",X"B2",X"67",X"B2",X"6A",X"B2",X"71",X"B2",X"78",X"B2",X"82",X"B2",X"8E",X"B2",
		X"9B",X"B2",X"AA",X"B2",X"BA",X"B2",X"CB",X"B2",X"E0",X"B2",X"F5",X"B2",X"0C",X"B3",X"22",X"B3",
		X"3E",X"B3",X"56",X"B3",X"71",X"B3",X"8E",X"B3",X"AE",X"B3",X"CC",X"B3",X"ED",X"B3",X"0D",X"B4",
		X"30",X"B4",X"53",X"B4",X"78",X"B4",X"9B",X"B4",X"C1",X"B4",X"E8",X"B4",X"0F",X"B5",X"39",X"B5",
		X"61",X"B5",X"89",X"B5",X"B4",X"B5",X"DF",X"B5",X"0A",X"B6",X"36",X"B6",X"64",X"B6",X"93",X"B6",
		X"C0",X"B6",X"ED",X"B6",X"1D",X"B7",X"4C",X"B7",X"7C",X"B7",X"AB",X"B7",X"DB",X"B7",X"0E",X"B8",
		X"40",X"B8",X"6F",X"B8",X"A3",X"B8",X"D6",X"B8",X"08",X"B9",X"3B",X"B9",X"6D",X"B9",X"A2",X"B9",
		X"D5",X"B9",X"0A",X"BA",X"3D",X"BA",X"71",X"BA",X"A7",X"BA",X"DB",X"BA",X"11",X"BB",X"46",X"BB",
		X"7A",X"BB",X"B1",X"BB",X"E6",X"BB",X"1B",X"BC",X"51",X"BC",X"89",X"BC",X"BD",X"BC",X"F4",X"BC",
		X"29",X"BD",X"61",X"BD",X"94",X"BD",X"D0",X"BD",X"05",X"BE",X"3F",X"BF",X"C9",X"C1",X"19",X"C5",
		X"EE",X"C8",X"0D",X"CD",X"57",X"D1",X"B2",X"D5",X"0D",X"DA",X"5A",X"DE",X"95",X"E2",X"BA",X"E6",
		X"C4",X"EA",X"B1",X"EE",X"82",X"F2",X"35",X"F6",X"CB",X"F9",X"43",X"FD",X"9F",X"00",X"DE",X"03",
		X"03",X"07",X"0D",X"0A",X"FB",X"0C",X"D2",X"0F",X"8F",X"12",X"37",X"15",X"C3",X"17",X"44",X"1A",
		X"5E",X"1C",X"03",X"1D",X"87",X"1C",X"50",X"1B",X"9F",X"19",X"9D",X"17",X"6F",X"15",X"24",X"13",
		X"D0",X"10",X"78",X"0E",X"27",X"0C",X"DF",X"09",X"A2",X"07",X"73",X"05",X"56",X"03",X"45",X"01",
		X"48",X"FF",X"58",X"FD",X"79",X"FB",X"AA",X"F9",X"EA",X"F7",X"39",X"F6",X"94",X"F4",X"00",X"F3",
		X"79",X"F1",X"00",X"F0",X"93",X"EE",X"34",X"ED",X"DE",X"EB",X"98",X"EA",X"5B",X"E9",X"2A",X"E8",
		X"04",X"E7",X"E8",X"E5",X"D8",X"E4",X"D2",X"E3",X"D1",X"E2",X"DE",X"E1",X"F1",X"E0",X"10",X"E0",
		X"36",X"DF",X"63",X"DE",X"98",X"DD",X"D7",X"DC",X"1B",X"DC",X"69",X"DB",X"BB",X"DA",X"16",X"DA",
		X"75",X"D9",X"DE",X"D8",X"4B",X"D8",X"BF",X"D7",X"39",X"D7",X"B8",X"D6",X"3B",X"D6",X"C7",X"D5",
		X"54",X"D5",X"E7",X"D4",X"82",X"D4",X"1F",X"D4",X"C1",X"D3",X"69",X"D3",X"12",X"D3",X"C0",X"D2",
		X"74",X"D2",X"2A",X"D2",X"E5",X"D1",X"A3",X"D1",X"66",X"D1",X"2B",X"D1",X"F3",X"D0",X"BF",X"D0",
		X"8D",X"D0",X"5E",X"D0",X"33",X"D0",X"0B",X"D0",X"E5",X"CF",X"C2",X"CF",X"A1",X"CF",X"84",X"CF",
		X"68",X"CF",X"4F",X"CF",X"38",X"CF",X"23",X"CF",X"0F",X"CF",X"FF",X"CE",X"F0",X"CE",X"E3",X"CE",
		X"D9",X"CE",X"CF",X"CE",X"C8",X"CE",X"C1",X"CE",X"BE",X"CE",X"BA",X"CE",X"B9",X"CE",X"B9",X"CE",
		X"BD",X"CE",X"BF",X"CE",X"C4",X"CE",X"C8",X"CE",X"D0",X"CE",X"D7",X"CE",X"E2",X"CE",X"ED",X"CE",
		X"F7",X"CE",X"04",X"CF",X"11",X"CF",X"1F",X"CF",X"2F",X"CF",X"3F",X"CF",X"51",X"CF",X"63",X"CF",
		X"76",X"CF",X"8A",X"CF",X"9E",X"CF",X"B2",X"CF",X"CA",X"CF",X"DF",X"CF",X"F7",X"CF",X"0E",X"D0",
		X"28",X"D0",X"40",X"D0",X"5B",X"D0",X"74",X"D0",X"90",X"D0",X"AA",X"D0",X"C6",X"D0",X"E1",X"D0",
		X"FF",X"D0",X"1C",X"D1",X"3A",X"D1",X"55",X"D1",X"76",X"D1",X"91",X"D1",X"B4",X"D1",X"CE",X"D1",
		X"F4",X"D1",X"08",X"D2",X"A5",X"D2",X"AD",X"D4",X"A5",X"D7",X"3E",X"DB",X"2F",X"DF",X"57",X"E3",
		X"98",X"E7",X"DF",X"EB",X"1F",X"F0",X"4E",X"F4",X"67",X"F8",X"67",X"FC",X"4B",X"00",X"13",X"04",
		X"BD",X"07",X"4B",X"0B",X"BA",X"0E",X"0E",X"12",X"45",X"15",X"61",X"18",X"62",X"1B",X"4B",X"1E",
		X"16",X"21",X"CE",X"23",X"68",X"26",X"EF",X"28",X"5D",X"2B",X"B0",X"2D",X"DA",X"2E",X"A5",X"2E",
		X"9D",X"2D",X"00",X"2C",X"0A",X"2A",X"D6",X"27",X"86",X"25",X"20",X"23",X"BA",X"20",X"56",X"1E",
		X"FA",X"1B",X"A8",X"19",X"66",X"17",X"2F",X"15",X"0D",X"13",X"F6",X"10",X"F3",X"0E",X"FE",X"0C",
		X"18",X"0B",X"43",X"09",X"7D",X"07",X"C5",X"05",X"1D",X"04",X"81",X"02",X"F4",X"00",X"74",X"FF",
		X"01",X"FE",X"9A",X"FC",X"41",X"FB",X"F0",X"F9",X"AE",X"F8",X"74",X"F7",X"47",X"F6",X"24",X"F5",
		X"0B",X"F4",X"FC",X"F2",X"F5",X"F1",X"F8",X"F0",X"05",X"F0",X"19",X"EF",X"36",X"EE",X"5C",X"ED",
		X"89",X"EC",X"BF",X"EB",X"F9",X"EA",X"3E",X"EA",X"86",X"E9",X"DA",X"E8",X"31",X"E8",X"8F",X"E7",
		X"F1",X"E6",X"5E",X"E6",X"CB",X"E5",X"46",X"E5",X"BB",X"E4",X"25",X"E5",X"F1",X"E6",X"88",X"E9",
		X"B1",X"EC",X"28",X"F0",X"D4",X"F3",X"92",X"F7",X"58",X"FB",X"13",X"FF",X"C3",X"02",X"5F",X"06",
		X"E5",X"09",X"51",X"0D",X"A5",X"10",X"DF",X"13",X"FE",X"16",X"04",X"1A",X"F0",X"1C",X"C2",X"1F",
		X"7C",X"22",X"1F",X"25",X"AA",X"27",X"20",X"2A",X"7C",X"2C",X"C7",X"2E",X"F9",X"30",X"21",X"33",
		X"F3",X"34",X"5C",X"35",X"9C",X"34",X"1F",X"33",X"24",X"31",X"DC",X"2E",X"62",X"2C",X"D3",X"29",
		X"37",X"27",X"9A",X"24",X"03",X"22",X"7B",X"1F",X"FD",X"1C",X"92",X"1A",X"34",X"18",X"E8",X"15",
		X"AE",X"13",X"86",X"11",X"6E",X"0F",X"67",X"0D",X"70",X"0B",X"8C",X"09",X"B7",X"07",X"F1",X"05",
		X"39",X"04",X"8F",X"02",X"F4",X"00",X"68",X"FF",X"E8",X"FD",X"76",X"FC",X"0E",X"FB",X"B6",X"F9",
		X"66",X"F8",X"23",X"F7",X"EB",X"F5",X"BE",X"F4",X"9B",X"F3",X"82",X"F2",X"72",X"F1",X"6F",X"F0",
		X"71",X"EF",X"7F",X"EE",X"93",X"ED",X"B2",X"EC",X"D7",X"EB",X"06",X"EB",X"3C",X"EA",X"79",X"E9",
		X"BD",X"E8",X"09",X"E8",X"5A",X"E7",X"B3",X"E6",X"11",X"E6",X"77",X"E5",X"E0",X"E4",X"70",X"E4",
		X"49",X"E5",X"53",X"E7",X"14",X"EA",X"51",X"ED",X"D2",X"F0",X"7B",X"F4",X"34",X"F8",X"F0",X"FB",
		X"A0",X"FF",X"40",X"03",X"CD",X"06",X"45",X"0A",X"A1",X"0D",X"E6",X"10",X"0F",X"14",X"20",X"17",
		X"16",X"1A",X"F5",X"1C",X"B8",X"1F",X"65",X"22",X"FB",X"24",X"79",X"27",X"E2",X"29",X"35",X"2C",
		X"73",X"2E",X"9C",X"30",X"B1",X"32",X"B5",X"34",X"A2",X"36",X"82",X"38",X"4F",X"3A",X"09",X"3C",
		X"B4",X"3D",X"52",X"3F",X"DC",X"40",X"58",X"42",X"C6",X"43",X"26",X"45",X"79",X"46",X"BF",X"47",
		X"F7",X"48",X"23",X"4A",X"41",X"4B",X"58",X"4C",X"5F",X"4D",X"60",X"4E",X"50",X"4F",X"3D",X"50",
		X"19",X"51",X"F0",X"51",X"BB",X"52",X"80",X"53",X"35",X"54",X"F3",X"54",X"2A",X"55",X"F1",X"53",
		X"BB",X"51",X"DE",X"4E",X"9A",X"4B",X"18",X"48",X"74",X"44",X"C5",X"40",X"18",X"3D",X"74",X"39",
		X"E1",X"35",X"5E",X"32",X"F4",X"2E",X"A1",X"2B",X"65",X"28",X"42",X"25",X"36",X"22",X"43",X"1F",
		X"68",X"1C",X"A3",X"19",X"F6",X"16",X"5E",X"14",X"DD",X"11",X"6D",X"0F",X"17",X"0D",X"CF",X"0A",
		X"A1",X"08",X"82",X"06",X"7D",X"05",X"DD",X"05",X"0B",X"07",X"D4",X"08",X"F0",X"0A",X"49",X"0D",
		X"C0",X"0F",X"46",X"12",X"CA",X"14",X"4E",X"17",X"C5",X"19",X"30",X"1C",X"8A",X"1E",X"D5",X"20",
		X"0B",X"23",X"30",X"25",X"43",X"27",X"45",X"29",X"35",X"2B",X"13",X"2D",X"E2",X"2E",X"9F",X"30",
		X"4C",X"32",X"E9",X"33",X"78",X"35",X"F7",X"36",X"69",X"38",X"CD",X"39",X"23",X"3B",X"6B",X"3C",
		X"A6",X"3D",X"D8",X"3E",X"FB",X"3F",X"14",X"41",X"20",X"42",X"23",X"43",X"1A",X"44",X"09",X"45",
		X"ED",X"45",X"C7",X"46",X"9A",X"47",X"60",X"48",X"20",X"49",X"D8",X"49",X"86",X"4A",X"2D",X"4B",
		X"CC",X"4B",X"64",X"4C",X"F5",X"4C",X"7E",X"4D",X"00",X"4E",X"7D",X"4E",X"F3",X"4E",X"62",X"4F",
		X"CE",X"4F",X"30",X"50",X"90",X"50",X"E8",X"50",X"3B",X"51",X"8A",X"51",X"D3",X"51",X"19",X"52",
		X"59",X"52",X"95",X"52",X"CC",X"52",X"00",X"53",X"2F",X"53",X"5A",X"53",X"81",X"53",X"A5",X"53",
		X"C6",X"53",X"E3",X"53",X"FB",X"53",X"12",X"54",X"27",X"54",X"36",X"54",X"41",X"54",X"4D",X"54",
		X"54",X"54",X"5B",X"54",X"5A",X"54",X"60",X"54",X"2C",X"54",X"A6",X"52",X"00",X"50",X"A9",X"4C",
		X"E1",X"48",X"DA",X"44",X"AF",X"40",X"79",X"3C",X"45",X"38",X"1E",X"34",X"0A",X"30",X"0E",X"2C",
		X"2A",X"28",X"60",X"24",X"B4",X"20",X"22",X"1D",X"AE",X"19",X"53",X"16",X"17",X"13",X"F4",X"0F",
		X"EA",X"0C",X"F8",X"09",X"24",X"07",X"60",X"04",X"BB",X"01",X"24",X"FF",X"AF",X"FC",X"3D",X"FA",
		X"97",X"F8",X"72",X"F8",X"36",X"F9",X"A7",X"FA",X"7A",X"FC",X"93",X"FE",X"D0",X"00",X"22",X"03",
		X"7B",X"05",X"D4",X"07",X"22",X"0A",X"69",X"0C",X"9F",X"0E",X"C7",X"10",X"E0",X"12",X"E7",X"14",
		X"DD",X"16",X"C5",X"18",X"9B",X"1A",X"61",X"1C",X"17",X"1E",X"BF",X"1F",X"57",X"21",X"E2",X"22",
		X"5D",X"24",X"CB",X"25",X"2E",X"27",X"68",X"28",X"5C",X"28",X"12",X"27",X"0A",X"25",X"7B",X"22",
		X"9F",X"1F",X"93",X"1C",X"75",X"19",X"4B",X"16",X"29",X"13",X"0D",X"10",X"04",X"0D",X"0A",X"0A",
		X"25",X"07",X"55",X"04",X"9A",X"01",X"F4",X"FE",X"65",X"FC",X"E9",X"F9",X"84",X"F7",X"30",X"F5",
		X"F4",X"F2",X"C7",X"F0",X"B1",X"EE",X"A9",X"EC",X"B5",X"EA",X"D2",X"E8",X"00",X"E7",X"3E",X"E5",
		X"8B",X"E3",X"E7",X"E1",X"53",X"E0",X"CC",X"DE",X"55",X"DD",X"EB",X"DB",X"8C",X"DA",X"3B",X"D9",
		X"F6",X"D7",X"BE",X"D6",X"91",X"D5",X"6F",X"D4",X"57",X"D3",X"4B",X"D2",X"48",X"D1",X"4F",X"D0",
		X"61",X"CF",X"7B",X"CE",X"9F",X"CD",X"C9",X"CC",X"FF",X"CB",X"3B",X"CB",X"80",X"CA",X"CC",X"C9",
		X"1F",X"C9",X"7C",X"C8",X"DE",X"C7",X"46",X"C7",X"B5",X"C6",X"2B",X"C6",X"A8",X"C5",X"28",X"C5",
		X"B1",X"C4",X"3E",X"C4",X"D1",X"C3",X"69",X"C3",X"08",X"C3",X"AA",X"C2",X"51",X"C2",X"FD",X"C1",
		X"AC",X"C1",X"61",X"C1",X"1B",X"C1",X"D9",X"C0",X"99",X"C0",X"5D",X"C0",X"26",X"C0",X"F2",X"BF",
		X"C2",X"BF",X"95",X"BF",X"6B",X"BF",X"45",X"BF",X"21",X"BF",X"02",X"BF",X"E3",X"BE",X"C9",X"BE",
		X"B2",X"BE",X"9C",X"BE",X"89",X"BE",X"78",X"BE",X"6B",X"BE",X"5F",X"BE",X"56",X"BE",X"4D",X"BE",
		X"49",X"BE",X"45",X"BE",X"44",X"BE",X"44",X"BE",X"46",X"BE",X"4B",X"BE",X"50",X"BE",X"58",X"BE",
		X"60",X"BE",X"6C",X"BE",X"76",X"BE",X"86",X"BE",X"93",X"BE",X"A6",X"BE",X"B5",X"BE",X"C9",X"BE",
		X"DB",X"BE",X"F1",X"BE",X"06",X"BF",X"1F",X"BF",X"36",X"BF",X"4F",X"BF",X"6A",X"BF",X"86",X"BF",
		X"A0",X"BF",X"BE",X"BF",X"DC",X"BF",X"FA",X"BF",X"1A",X"C0",X"3B",X"C0",X"5B",X"C0",X"7C",X"C0",
		X"9E",X"C0",X"C2",X"C0",X"E4",X"C0",X"0A",X"C1",X"2E",X"C1",X"53",X"C1",X"78",X"C1",X"A0",X"C1",
		X"C5",X"C1",X"ED",X"C1",X"14",X"C2",X"40",X"C2",X"5F",X"C2",X"C8",X"C2",X"8A",X"C4",X"5F",X"C7",
		X"E0",X"CA",X"CC",X"CE",X"F4",X"D2",X"39",X"D7",X"8B",X"DB",X"D5",X"DF",X"14",X"E4",X"3A",X"E8",
		X"4B",X"EC",X"3F",X"F0",X"18",X"F4",X"D3",X"F7",X"6F",X"FB",X"F1",X"FE",X"55",X"02",X"9C",X"05",
		X"CA",X"08",X"DA",X"0B",X"D1",X"0E",X"AD",X"11",X"73",X"14",X"1D",X"17",X"B7",X"19",X"2D",X"1C",
		X"A1",X"1E",X"30",X"20",X"43",X"20",X"75",X"1F",X"FA",X"1D",X"20",X"1C",X"02",X"1A",X"C3",X"17",
		X"6C",X"15",X"0E",X"13",X"B2",X"10",X"5F",X"0E",X"15",X"0C",X"D9",X"09",X"AA",X"07",X"8C",X"05",
		X"7F",X"03",X"81",X"01",X"93",X"FF",X"B5",X"FD",X"E7",X"FB",X"27",X"FA",X"76",X"F8",X"D5",X"F6",
		X"41",X"F5",X"BB",X"F3",X"42",X"F2",X"D4",X"F0",X"98",X"EF",X"B1",X"EF",X"FC",X"F0",X"02",X"F3",
		X"8B",X"F5",X"5A",X"F8",X"5A",X"FB",X"6D",X"FE",X"87",X"01",X"9B",X"04",X"A8",X"07",X"A1",X"0A",
		X"8A",X"0D",X"5D",X"10",X"1F",X"13",X"C9",X"15",X"5E",X"18",X"DB",X"1A",X"45",X"1D",X"99",X"1F",
		X"DB",X"21",X"07",X"24",X"20",X"26",X"26",X"28",X"1A",X"2A",X"FC",X"2B",X"CD",X"2D",X"8D",X"2F",
		X"3E",X"31",X"DD",X"32",X"6F",X"34",X"EF",X"35",X"65",X"37",X"C9",X"38",X"23",X"3A",X"6B",X"3B",
		X"AC",X"3C",X"DC",X"3D",X"04",X"3F",X"1D",X"40",X"2D",X"41",X"31",X"42",X"2D",X"43",X"1A",X"44",
		X"02",X"45",X"DE",X"45",X"B0",X"46",X"7A",X"47",X"3A",X"48",X"F2",X"48",X"A3",X"49",X"4D",X"4A",
		X"EC",X"4A",X"86",X"4B",X"19",X"4C",X"93",X"4C",X"DD",X"4B",X"E2",X"49",X"29",X"47",X"EF",X"43",
		X"69",X"40",X"B7",X"3C",X"F3",X"38",X"29",X"35",X"6B",X"31",X"B7",X"2D",X"19",X"2A",X"8F",X"26",
		X"1F",X"23",X"C7",X"1F",X"86",X"1C",X"60",X"19",X"52",X"16",X"5E",X"13",X"81",X"10",X"BC",X"0D",
		X"0E",X"0B",X"76",X"08",X"F3",X"05",X"88",X"03",X"2E",X"01",X"ED",X"FE",X"BD",X"FC",X"A7",X"FB",
		X"FE",X"FB",X"24",X"FD",X"E3",X"FE",X"FA",X"00",X"4C",X"03",X"BC",X"05",X"3E",X"08",X"BD",X"0A",
		X"3E",X"0D",X"AF",X"0F",X"17",X"12",X"6D",X"14",X"B5",X"16",X"E9",X"18",X"0D",X"1B",X"1D",X"1D",
		X"1F",X"1F",X"0D",X"21",X"EB",X"22",X"B9",X"24",X"75",X"26",X"22",X"28",X"BF",X"29",X"4E",X"2B",
		X"CF",X"2C",X"41",X"2E",X"A5",X"2F",X"FC",X"30",X"48",X"32",X"85",X"33",X"B7",X"34",X"DD",X"35",
		X"F9",X"36",X"08",X"38",X"0E",X"39",X"08",X"3A",X"F8",X"3A",X"E0",X"3B",X"BD",X"3C",X"92",X"3D",
		X"5E",X"3E",X"21",X"3F",X"DB",X"3F",X"8E",X"40",X"3A",X"41",X"DE",X"41",X"79",X"42",X"0C",X"43",
		X"9C",X"43",X"21",X"44",X"A3",X"44",X"1E",X"45",X"93",X"45",X"01",X"46",X"69",X"46",X"CD",X"46",
		X"2B",X"47",X"86",X"47",X"D9",X"47",X"27",X"48",X"72",X"48",X"B7",X"48",X"F8",X"48",X"37",X"49",
		X"70",X"49",X"A4",X"49",X"D5",X"49",X"03",X"4A",X"2B",X"4A",X"52",X"4A",X"74",X"4A",X"93",X"4A",
		X"B1",X"4A",X"C9",X"4A",X"DF",X"4A",X"F3",X"4A",X"03",X"4B",X"11",X"4B",X"1D",X"4B",X"26",X"4B",
		X"2B",X"4B",X"2D",X"4B",X"30",X"4B",X"2F",X"4B",X"2C",X"4B",X"26",X"4B",X"21",X"4B",X"17",X"4B",
		X"0C",X"4B",X"FF",X"4A",X"F1",X"4A",X"E2",X"4A",X"CF",X"4A",X"BB",X"4A",X"A8",X"4A",X"92",X"4A",
		X"78",X"4A",X"5F",X"4A",X"46",X"4A",X"28",X"4A",X"0E",X"4A",X"ED",X"49",X"D0",X"49",X"AE",X"49",
		X"8F",X"49",X"69",X"49",X"4B",X"49",X"1F",X"49",X"05",X"49",X"28",X"48",X"DD",X"45",X"B9",X"42",
		X"FD",X"3E",X"F0",X"3A",X"AC",X"36",X"58",X"32",X"FB",X"2D",X"AB",X"29",X"68",X"25",X"40",X"21",
		X"2E",X"1D",X"3A",X"19",X"60",X"15",X"A7",X"11",X"06",X"0E",X"86",X"0A",X"22",X"07",X"DA",X"03",
		X"AD",X"00",X"9C",X"FD",X"A3",X"FA",X"C3",X"F7",X"FE",X"F4",X"4F",X"F2",X"B7",X"EF",X"36",X"ED",
		X"CB",X"EA",X"75",X"E8",X"32",X"E6",X"05",X"E4",X"EB",X"E1",X"E4",X"DF",X"EE",X"DD",X"09",X"DC",
		X"38",X"DA",X"75",X"D8",X"C4",X"D6",X"1F",X"D5",X"8C",X"D3",X"06",X"D2",X"91",X"D0",X"27",X"CF",
		X"CD",X"CD",X"7C",X"CC",X"3B",X"CB",X"04",X"CA",X"DA",X"C8",X"B9",X"C7",X"A8",X"C6",X"9C",X"C5",
		X"A1",X"C4",X"A8",X"C3",X"C3",X"C2",X"D5",X"C1",X"8A",X"C1",X"B7",X"C2",X"D6",X"C4",X"9C",X"C7",
		X"C2",X"CA",X"29",X"CE",X"AC",X"D1",X"3C",X"D5",X"CA",X"D8",X"4F",X"DC",X"C5",X"DF",X"28",X"E3",
		X"72",X"E6",X"A9",X"E9",X"C7",X"EC",X"CB",X"EF",X"B9",X"F2",X"8F",X"F5",X"4E",X"F8",X"F6",X"FA",
		X"88",X"FD",X"03",X"00",X"6A",X"02",X"BB",X"04",X"FA",X"06",X"25",X"09",X"3C",X"0B",X"36",X"0D",
		X"FD",X"0D",X"6A",X"0D",X"0C",X"0C",X"1B",X"0A",X"D6",X"07",X"57",X"05",X"C0",X"02",X"16",X"00",
		X"71",X"FD",X"CC",X"FA",X"38",X"F8",X"AF",X"F5",X"37",X"F3",X"CE",X"F0",X"7A",X"EE",X"36",X"EC",
		X"09",X"EA",X"E9",X"E7",X"DF",X"E5",X"E5",X"E3",X"FD",X"E1",X"24",X"E0",X"5F",X"DE",X"A9",X"DC",
		X"00",X"DB",X"68",X"D9",X"DF",X"D7",X"64",X"D6",X"F4",X"D4",X"94",X"D3",X"42",X"D2",X"F9",X"D0",
		X"BF",X"CF",X"8F",X"CE",X"6B",X"CD",X"53",X"CC",X"45",X"CB",X"40",X"CA",X"48",X"C9",X"59",X"C8",
		X"73",X"C7",X"96",X"C6",X"C1",X"C5",X"F7",X"C4",X"34",X"C4",X"7A",X"C3",X"C6",X"C2",X"1B",X"C2",
		X"75",X"C1",X"DB",X"C0",X"43",X"C0",X"B7",X"BF",X"2B",X"BF",X"AD",X"BE",X"2F",X"BE",X"B7",X"BE",
		X"9C",X"C0",X"4D",X"C3",X"90",X"C6",X"20",X"CA",X"E3",X"CD",X"B9",X"D1",X"97",X"D5",X"6A",X"D9",
		X"33",X"DD",X"E7",X"E0",X"86",X"E4",X"0B",X"E8",X"76",X"EB",X"C9",X"EE",X"00",X"F2",X"1F",X"F5",
		X"24",X"F8",X"0E",X"FB",X"E3",X"FD",X"9C",X"00",X"41",X"03",X"CE",X"05",X"46",X"08",X"A9",X"0A",
		X"F7",X"0C",X"30",X"0F",X"56",X"11",X"6A",X"13",X"6B",X"15",X"5B",X"17",X"39",X"19",X"06",X"1B",
		X"C2",X"1C",X"70",X"1E",X"0E",X"20",X"9D",X"21",X"1E",X"23",X"93",X"24",X"F8",X"25",X"53",X"27",
		X"9D",X"28",X"DC",X"29",X"10",X"2B",X"3A",X"2C",X"55",X"2D",X"6A",X"2E",X"70",X"2F",X"6E",X"30",
		X"60",X"31",X"4D",X"32",X"2A",X"33",X"07",X"34",X"D0",X"34",X"A0",X"35",X"92",X"35",X"14",X"34",
		X"BB",X"31",X"C9",X"2E",X"80",X"2B",X"FD",X"27",X"65",X"24",X"C1",X"20",X"23",X"1D",X"90",X"19",
		X"0E",X"16",X"A0",X"12",X"49",X"0F",X"0A",X"0C",X"E4",X"08",X"D6",X"05",X"E0",X"02",X"02",X"00",
		X"3E",X"FD",X"90",X"FA",X"F8",X"F7",X"76",X"F5",X"0B",X"F3",X"B4",X"F0",X"71",X"EE",X"41",X"EC",
		X"25",X"EA",X"1C",X"E8",X"24",X"E6",X"3E",X"E4",X"68",X"E2",X"A5",X"E0",X"ED",X"DE",X"4A",X"DD",
		X"B3",X"DB",X"2B",X"DA",X"B2",X"D8",X"46",X"D7",X"E6",X"D5",X"95",X"D4",X"4F",X"D3",X"16",X"D2",
		X"E7",X"D0",X"C7",X"CF",X"AC",X"CE",X"A2",X"CD",X"9E",X"CC",X"A8",X"CB",X"B7",X"CA",X"D4",X"C9",
		X"F5",X"C8",X"24",X"C8",X"55",X"C7",X"9A",X"C6",X"D1",X"C5",X"BF",X"C5",X"25",X"C7",X"72",X"C9",
		X"61",X"CC",X"AD",X"CF",X"36",X"D3",X"D6",X"D6",X"85",X"DA",X"2C",X"DE",X"CC",X"E1",X"5A",X"E5",
		X"D4",X"E8",X"35",X"EC",X"81",X"EF",X"B2",X"F2",X"CC",X"F5",X"CA",X"F8",X"B3",X"FB",X"82",X"FE",
		X"39",X"01",X"DB",X"03",X"66",X"06",X"DA",X"08",X"3C",X"0B",X"86",X"0D",X"BC",X"0F",X"E0",X"11",
		X"F3",X"13",X"F0",X"15",X"DD",X"17",X"BB",X"19",X"85",X"1B",X"41",X"1D",X"EC",X"1E",X"89",X"20",
		X"17",X"22",X"96",X"23",X"07",X"25",X"6C",X"26",X"C2",X"27",X"0C",X"29",X"4B",X"2A",X"7F",X"2B",
		X"A6",X"2C",X"C2",X"2D",X"D3",X"2E",X"D9",X"2F",X"D5",X"30",X"C8",X"31",X"AF",X"32",X"91",X"33",
		X"67",X"34",X"36",X"35",X"FA",X"35",X"B7",X"36",X"6D",X"37",X"1D",X"38",X"C3",X"38",X"63",X"39",
		X"F9",X"39",X"8C",X"3A",X"15",X"3B",X"9C",X"3B",X"1A",X"3C",X"93",X"3C",X"05",X"3D",X"72",X"3D",
		X"D9",X"3D",X"3D",X"3E",X"99",X"3E",X"F3",X"3E",X"44",X"3F",X"97",X"3F",X"DC",X"3F",X"28",X"40",
		X"65",X"40",X"A8",X"40",X"DD",X"40",X"18",X"41",X"44",X"41",X"7D",X"41",X"97",X"41",X"EF",X"41",
		X"A1",X"42",X"B4",X"42",X"DA",X"42",X"F2",X"42",X"0F",X"43",X"23",X"43",X"38",X"43",X"46",X"43",
		X"58",X"43",X"60",X"43",X"6D",X"43",X"72",X"43",X"77",X"43",X"7A",X"43",X"7C",X"43",X"7A",X"43",
		X"78",X"43",X"72",X"43",X"6C",X"43",X"61",X"43",X"59",X"43",X"4B",X"43",X"3F",X"43",X"2E",X"43",
		X"22",X"43",X"0B",X"43",X"FD",X"42",X"F9",X"41",X"8F",X"3F",X"5C",X"3C",X"96",X"38",X"84",X"34",
		X"42",X"30",X"F1",X"2B",X"9A",X"27",X"50",X"23",X"14",X"1F",X"F1",X"1A",X"E9",X"16",X"FC",X"12",
		X"2A",X"0F",X"78",X"0B",X"E1",X"07",X"68",X"04",X"0C",X"01",X"CD",X"FD",X"A8",X"FA",X"9B",X"F7",
		X"AC",X"F4",X"D4",X"F1",X"15",X"EF",X"6D",X"EC",X"DF",X"E9",X"5E",X"E7",X"34",X"E5",X"80",X"E4",
		X"FC",X"E4",X"3A",X"E6",X"FA",X"E7",X"0B",X"EA",X"4B",X"EC",X"A9",X"EE",X"11",X"F1",X"7D",X"F3",
		X"E1",X"F5",X"3C",X"F8",X"8B",X"FA",X"CE",X"FC",X"FD",X"FE",X"1A",X"01",X"2B",X"03",X"2A",X"05",
		X"18",X"07",X"F6",X"08",X"C4",X"0A",X"83",X"0C",X"32",X"0E",X"D4",X"0F",X"66",X"11",X"EA",X"12",
		X"61",X"14",X"CB",X"15",X"29",X"17",X"78",X"18",X"BF",X"19",X"F6",X"1A",X"24",X"1C",X"47",X"1D",
		X"5E",X"1E",X"6C",X"1F",X"70",X"20",X"6A",X"21",X"5A",X"22",X"42",X"23",X"20",X"24",X"F8",X"24",
		X"C5",X"25",X"8C",X"26",X"49",X"27",X"00",X"28",X"AF",X"28",X"58",X"29",X"F9",X"29",X"93",X"2A",
		X"27",X"2B",X"B5",X"2B",X"3E",X"2C",X"BE",X"2C",X"3A",X"2D",X"B2",X"2D",X"23",X"2E",X"8E",X"2E",
		X"F6",X"2E",X"58",X"2F",X"B7",X"2F",X"0F",X"30",X"65",X"30",X"B4",X"30",X"FF",X"30",X"47",X"31",
		X"8D",X"31",X"CB",X"31",X"0A",X"32",X"42",X"32",X"79",X"32",X"AA",X"32",X"DB",X"32",X"06",X"33",
		X"30",X"33",X"55",X"33",X"7B",X"33",X"97",X"33",X"B9",X"33",X"D2",X"33",X"EE",X"33",X"FF",X"33",
		X"1F",X"34",X"9C",X"33",X"A3",X"31",X"C1",X"2E",X"3C",X"2B",X"5D",X"27",X"44",X"23",X"15",X"1F",
		X"DE",X"1A",X"B0",X"16",X"8F",X"12",X"85",X"0E",X"92",X"0A",X"BD",X"06",X"01",X"03",X"64",X"FF",
		X"E2",X"FB",X"7C",X"F8",X"33",X"F5",X"03",X"F2",X"F1",X"EE",X"F7",X"EB",X"18",X"E9",X"53",X"E6",
		X"A4",X"E3",X"0E",X"E1",X"8D",X"DE",X"24",X"DC",X"DD",X"D9",X"D9",X"D8",X"2E",X"D9",X"51",X"DA",
		X"0C",X"DC",X"1D",X"DE",X"6A",X"E0",X"D1",X"E2",X"4C",X"E5",X"C9",X"E7",X"43",X"EA",X"B3",X"EC",
		X"17",X"EF",X"6A",X"F1",X"AF",X"F3",X"E2",X"F5",X"07",X"F8",X"1A",X"FA",X"1C",X"FC",X"0D",X"FE",
		X"EF",X"FF",X"BE",X"01",X"81",X"03",X"33",X"05",X"D8",X"06",X"6D",X"08",X"F4",X"09",X"6E",X"0B",
		X"DC",X"0C",X"3C",X"0E",X"91",X"0F",X"DB",X"10",X"19",X"12",X"49",X"13",X"71",X"14",X"8C",X"15",
		X"A0",X"16",X"A7",X"17",X"A6",X"18",X"9B",X"19",X"87",X"1A",X"6A",X"1B",X"48",X"1C",X"19",X"1D",
		X"E4",X"1D",X"A5",X"1E",X"62",X"1F",X"17",X"20",X"C3",X"20",X"6C",X"21",X"09",X"22",X"A5",X"22",
		X"35",X"23",X"C6",X"23",X"4A",X"24",X"CA",X"24",X"3F",X"24",X"53",X"22",X"9D",X"1F",X"57",X"1C",
		X"C4",X"18",X"FC",X"14",X"23",X"11",X"44",X"0D",X"6F",X"09",X"A6",X"05",X"F3",X"01",X"55",X"FE",
		X"D3",X"FA",X"68",X"F7",X"1A",X"F4",X"E5",X"F0",X"CA",X"ED",X"C9",X"EA",X"E4",X"E7",X"15",X"E5",
		X"5F",X"E2",X"C0",X"DF",X"38",X"DD",X"C7",X"DA",X"6E",X"D8",X"26",X"D6",X"F5",X"D3",X"D8",X"D1",
		X"CD",X"CF",X"D5",X"CD",X"EF",X"CB",X"1B",X"CA",X"57",X"C8",X"A5",X"C6",X"01",X"C5",X"6E",X"C3",
		X"EA",X"C1",X"74",X"C0",X"0C",X"BF",X"B3",X"BD",X"66",X"BC",X"28",X"BB",X"F5",X"B9",X"CD",X"B8",
		X"B1",X"B7",X"A2",X"B6",X"9C",X"B5",X"A3",X"B4",X"B3",X"B3",X"CD",X"B2",X"F0",X"B1",X"1E",X"B1",
		X"53",X"B0",X"93",X"AF",X"DB",X"AE",X"2A",X"AE",X"83",X"AD",X"E3",X"AC",X"4A",X"AC",X"B9",X"AB",
		X"31",X"AB",X"AC",X"AA",X"30",X"AA",X"B8",X"A9",X"4A",X"A9",X"DF",X"A8",X"7D",X"A8",X"1F",X"A8",
		X"C6",X"A7",X"71",X"A7",X"23",X"A7",X"DC",X"A6",X"97",X"A6",X"58",X"A6",X"1D",X"A6",X"E5",X"A5",
		X"B4",X"A5",X"84",X"A5",X"5D",X"A5",X"33",X"A5",X"12",X"A5",X"F0",X"A4",X"00",X"A5",X"6C",X"A6",
		X"01",X"A9",X"4A",X"AC",X"0A",X"B0",X"0D",X"B4",X"33",X"B8",X"68",X"BC",X"99",X"C0",X"C1",X"C4",
		X"D5",X"C8",X"D4",X"CC",X"B8",X"D0",X"81",X"D4",X"30",X"D8",X"C3",X"DB",X"37",X"DF",X"93",X"E2",
		X"D4",X"E5",X"F9",X"E8",X"03",X"EC",X"F8",X"EE",X"CE",X"F1",X"92",X"F4",X"38",X"F7",X"D3",X"F9",
		X"49",X"FC",X"BE",X"FE",X"68",X"00",X"8C",X"00",X"BD",X"FF",X"3F",X"FE",X"5B",X"FC",X"2F",X"FA",
		X"DF",X"F7",X"78",X"F5",X"0D",X"F3",X"A1",X"F0",X"40",X"EE",X"E7",X"EB",X"9F",X"E9",X"66",X"E7",
		X"3E",X"E5",X"24",X"E3",X"21",X"E1",X"2A",X"DF",X"45",X"DD",X"71",X"DB",X"AE",X"D9",X"FA",X"D7",
		X"57",X"D6",X"BF",X"D4",X"3A",X"D3",X"C0",X"D1",X"56",X"D0",X"0E",X"CF",X"0F",X"CF",X"5C",X"D0",
		X"69",X"D2",X"03",X"D5",X"EA",X"D7",X"01",X"DB",X"31",X"DE",X"68",X"E1",X"9B",X"E4",X"C5",X"E7",
		X"DE",X"EA",X"E6",X"ED",X"DC",X"F0",X"BB",X"F3",X"83",X"F6",X"38",X"F9",X"D4",X"FB",X"5C",X"FE",
		X"D0",X"00",X"2D",X"03",X"79",X"05",X"AE",X"07",X"D5",X"09",X"E4",X"0B",X"E7",X"0D",X"CE",X"0F",
		X"B7",X"11",X"05",X"13",X"CD",X"12",X"94",X"11",X"AA",X"0F",X"56",X"0D",X"BA",X"0A",X"FA",X"07",
		X"27",X"05",X"4E",X"02",X"78",X"FF",X"B1",X"FC",X"F4",X"F9",X"49",X"F7",X"AF",X"F4",X"2B",X"F2",
		X"B8",X"EF",X"5A",X"ED",X"10",X"EB",X"DA",X"E8",X"B4",X"E6",X"A4",X"E4",X"A5",X"E2",X"B7",X"E0",
		X"D9",X"DE",X"0F",X"DD",X"54",X"DB",X"A6",X"D9",X"0A",X"D8",X"7D",X"D6",X"FE",X"D4",X"8D",X"D3",
		X"28",X"D2",X"D2",X"D0",X"87",X"CF",X"4A",X"CE",X"17",X"CD",X"F2",X"CB",X"D8",X"CA",X"C5",X"C9",
		X"C2",X"C8",X"C5",X"C7",X"D5",X"C6",X"EC",X"C5",X"0E",X"C5",X"37",X"C4",X"6E",X"C3",X"A7",X"C2",
		X"EE",X"C1",X"36",X"C1",X"8E",X"C0",X"E4",X"BF",X"4E",X"BF",X"AE",X"BE",X"2A",X"BE",X"8C",X"BD",
		X"75",X"BD",X"3A",X"BE",X"63",X"C0",X"82",X"C3",X"F1",X"C6",X"B6",X"CA",X"8B",X"CE",X"7A",X"D2",
		X"5C",X"D6",X"3D",X"DA",X"04",X"DE",X"BD",X"E1",X"59",X"E5",X"DE",X"E8",X"47",X"EC",X"9B",X"EF",
		X"CE",X"F2",X"EC",X"F5",X"EE",X"F8",X"D7",X"FB",X"A8",X"FE",X"60",X"01",X"02",X"04",X"8E",X"06",
		X"07",X"09",X"62",X"0B",X"B7",X"0D",X"AE",X"0F",X"2A",X"10",X"7A",X"0F",X"0A",X"0E",X"19",X"0C",
		X"D9",X"09",X"68",X"07",X"E0",X"04",X"4C",X"02",X"B9",X"FF",X"2D",X"FD",X"AA",X"FA",X"37",X"F8",
		X"D4",X"F5",X"81",X"F3",X"40",X"F1",X"12",X"EF",X"F5",X"EC",X"EA",X"EA",X"F1",X"E8",X"08",X"E7",
		X"31",X"E5",X"6A",X"E3",X"B3",X"E1",X"0A",X"E0",X"71",X"DE",X"E6",X"DC",X"6A",X"DB",X"FA",X"D9",
		X"9A",X"D8",X"44",X"D7",X"FC",X"D5",X"C0",X"D4",X"8F",X"D3",X"6A",X"D2",X"52",X"D1",X"41",X"D0",
		X"3E",X"CF",X"40",X"CE",X"51",X"CD",X"69",X"CC",X"8A",X"CB",X"B4",X"CA",X"E8",X"C9",X"23",X"C9",
		X"66",X"C8",X"B2",X"C7",X"05",X"C7",X"5F",X"C6",X"C0",X"C5",X"29",X"C5",X"98",X"C4",X"0D",X"C4",
		X"89",X"C3",X"09",X"C3",X"91",X"C2",X"1F",X"C2",X"B2",X"C1",X"4B",X"C1",X"E9",X"C0",X"8C",X"C0",
		X"33",X"C0",X"DF",X"BF",X"91",X"BF",X"46",X"BF",X"FE",X"BE",X"BE",X"BE",X"7D",X"BE",X"44",X"BE",
		X"0E",X"BE",X"DB",X"BD",X"AB",X"BD",X"80",X"BD",X"57",X"BD",X"33",X"BD",X"10",X"BD",X"F1",X"BC",
		X"D4",X"BC",X"BB",X"BC",X"A6",X"BC",X"91",X"BC",X"80",X"BC",X"71",X"BC",X"63",X"BC",X"5A",X"BC",
		X"52",X"BC",X"4D",X"BC",X"49",X"BC",X"46",X"BC",X"47",X"BC",X"4A",X"BC",X"4D",X"BC",X"53",X"BC",
		X"5B",X"BC",X"64",X"BC",X"6F",X"BC",X"7C",X"BC",X"89",X"BC",X"9A",X"BC",X"A8",X"BC",X"BC",X"BC",
		X"D0",X"BC",X"E2",X"BC",X"FB",X"BC",X"10",X"BD",X"28",X"BD",X"42",X"BD",X"5C",X"BD",X"76",X"BD",
		X"92",X"BD",X"C1",X"BD",X"26",X"BF",X"D0",X"C1",X"39",X"C5",X"24",X"C9",X"55",X"CD",X"AF",X"D1",
		X"14",X"D6",X"7C",X"DA",X"D3",X"DE",X"1A",X"E3",X"47",X"E7",X"5B",X"EB",X"50",X"EF",X"2A",X"F3",
		X"E4",X"F6",X"84",X"FA",X"02",X"FE",X"65",X"01",X"A9",X"04",X"D5",X"07",X"E3",X"0A",X"DA",X"0D",
		X"B7",X"10",X"7B",X"13",X"25",X"16",X"BB",X"18",X"35",X"1B",X"9F",X"1D",X"F0",X"1F",X"2E",X"22",
		X"57",X"24",X"6D",X"26",X"6E",X"28",X"61",X"2A",X"40",X"2C",X"0E",X"2E",X"CB",X"2F",X"78",X"31",
		X"16",X"33",X"A4",X"34",X"22",X"36",X"94",X"37",X"F8",X"38",X"4D",X"3A",X"96",X"3B",X"D2",X"3C",
		X"03",X"3E",X"27",X"3F",X"3F",X"40",X"4C",X"41",X"4F",X"42",X"46",X"43",X"37",X"44",X"17",X"45",
		X"F0",X"45",X"AE",X"45",X"09",X"44",X"95",X"41",X"8D",X"3E",X"36",X"3B",X"A8",X"37",X"05",X"34",
		X"5A",X"30",X"B4",X"2C",X"19",X"29",X"93",X"25",X"1E",X"22",X"C1",X"1E",X"7B",X"1B",X"51",X"18",
		X"3C",X"15",X"42",X"12",X"5D",X"0F",X"92",X"0C",X"DC",X"09",X"40",X"07",X"B5",X"04",X"43",X"02",
		X"E7",X"FF",X"9D",X"FD",X"66",X"FB",X"42",X"F9",X"32",X"F7",X"34",X"F5",X"46",X"F3",X"69",X"F1",
		X"9B",X"EF",X"DE",X"ED",X"31",X"EC",X"93",X"EA",X"05",X"E9",X"80",X"E7",X"0D",X"E6",X"A5",X"E4",
		X"4B",X"E3",X"FE",X"E1",X"BC",X"E0",X"85",X"DF",X"59",X"DE",X"3A",X"DD",X"23",X"DC",X"18",X"DB",
		X"18",X"DA",X"1F",X"D9",X"33",X"D8",X"4B",X"D7",X"70",X"D6",X"9A",X"D5",X"D3",X"D4",X"09",X"D4",
		X"30",X"D4",X"C8",X"D5",X"38",X"D8",X"45",X"DB",X"A7",X"DE",X"3F",X"E2",X"EE",X"E5",X"A7",X"E9",
		X"59",X"ED",X"03",X"F1",X"95",X"F4",X"16",X"F8",X"7B",X"FB",X"CB",X"FE",X"00",X"02",X"1D",X"05",
		X"20",X"08",X"09",X"0B",X"DA",X"0D",X"94",X"10",X"35",X"13",X"C2",X"15",X"37",X"18",X"95",X"1A",
		X"E3",X"1C",X"17",X"1F",X"3F",X"21",X"1B",X"23",X"88",X"23",X"BE",X"22",X"31",X"21",X"20",X"1F",
		X"BF",X"1C",X"2B",X"1A",X"80",X"17",X"C8",X"14",X"13",X"12",X"63",X"0F",X"C0",X"0C",X"2A",X"0A",
		X"A7",X"07",X"33",X"05",X"D4",X"02",X"86",X"00",X"4B",X"FE",X"21",X"FC",X"0C",X"FA",X"06",X"F8",
		X"12",X"F6",X"2F",X"F4",X"5D",X"F2",X"9A",X"F0",X"E6",X"EE",X"40",X"ED",X"AC",X"EB",X"23",X"EA",
		X"A7",X"E8",X"3C",X"E7",X"DB",X"E5",X"87",X"E4",X"3F",X"E3",X"04",X"E2",X"D5",X"E0",X"B0",X"DF",
		X"94",X"DE",X"85",X"DD",X"7E",X"DC",X"82",X"DB",X"90",X"DA",X"A6",X"D9",X"C4",X"D8",X"EC",X"D7",
		X"1D",X"D7",X"53",X"D6",X"94",X"D5",X"DB",X"D4",X"2B",X"D4",X"82",X"D3",X"E0",X"D2",X"43",X"D2",
		X"AE",X"D1",X"1E",X"D1",X"96",X"D0",X"14",X"D0",X"95",X"CF",X"1D",X"CF",X"AB",X"CE",X"3D",X"CE",
		X"D5",X"CD",X"72",X"CD",X"14",X"CD",X"BA",X"CC",X"65",X"CC",X"13",X"CC",X"C9",X"CB",X"7D",X"CB",
		X"3B",X"CB",X"F8",X"CA",X"BB",X"CA",X"80",X"CA",X"4B",X"CA",X"17",X"CA",X"E8",X"C9",X"BB",X"C9",
		X"94",X"C9",X"6B",X"C9",X"4A",X"C9",X"24",X"C9",X"0D",X"C9",X"E3",X"C8",X"53",X"C9",X"3E",X"CB",
		X"1A",X"CE",X"9C",X"D1",X"7C",X"D5",X"96",X"D9",X"CB",X"DD",X"06",X"E2",X"3A",X"E6",X"61",X"EA",
		X"71",X"EE",X"6A",X"F2",X"48",X"F6",X"08",X"FA",X"AD",X"FD",X"35",X"01",X"A1",X"04",X"EF",X"07",
		X"24",X"0B",X"3B",X"0E",X"3A",X"11",X"1E",X"14",X"E8",X"16",X"9B",X"19",X"35",X"1C",X"B9",X"1E",
		X"29",X"21",X"81",X"23",X"C3",X"25",X"F2",X"27",X"0D",X"2A",X"15",X"2C",X"0C",X"2E",X"EF",X"2F",
		X"C1",X"31",X"82",X"33",X"33",X"35",X"D4",X"36",X"65",X"38",X"E7",X"39",X"5B",X"3B",X"C3",X"3C",
		X"1B",X"3E",X"65",X"3F",X"A5",X"40",X"D7",X"41",X"FC",X"42",X"18",X"44",X"26",X"45",X"2B",X"46",
		X"24",X"47",X"14",X"48",X"F8",X"48",X"D4",X"49",X"A6",X"4A",X"6F",X"4B",X"30",X"4C",X"E8",X"4C",
		X"97",X"4D",X"40",X"4E",X"DD",X"4E",X"78",X"4F",X"06",X"50",X"92",X"50",X"13",X"51",X"91",X"51",
		X"04",X"52",X"78",X"52",X"DF",X"52",X"46",X"53",X"A0",X"53",X"FC",X"53",X"4C",X"54",X"9E",X"54",
		X"E4",X"54",X"2E",X"55",X"68",X"55",X"AA",X"55",X"DA",X"55",X"16",X"56",X"38",X"56",X"72",X"56",
		X"81",X"56",X"E6",X"56",X"BB",X"57",X"C7",X"57",X"EB",X"57",X"F9",X"57",X"10",X"58",X"1B",X"58",
		X"2C",X"58",X"31",X"58",X"3A",X"58",X"3D",X"58",X"40",X"58",X"3F",X"58",X"3A",X"58",X"35",X"58",
		X"2B",X"58",X"24",X"58",X"16",X"58",X"08",X"58",X"F5",X"57",X"E4",X"57",X"CE",X"57",X"BA",X"57",
		X"9E",X"57",X"88",X"57",X"69",X"57",X"55",X"57",X"F4",X"56",X"29",X"55",X"3F",X"52",X"A4",X"4E",
		X"96",X"4A",X"4C",X"46",X"DD",X"41",X"66",X"3D",X"F3",X"38",X"8E",X"34",X"3D",X"30",X"07",X"2C",
		X"E9",X"27",X"EB",X"23",X"07",X"20",X"45",X"1C",X"9D",X"18",X"17",X"15",X"A9",X"11",X"5A",X"0E",
		X"24",X"0B",X"0B",X"08",X"0A",X"05",X"24",X"02",X"55",X"FF",X"A1",X"FC",X"01",X"FA",X"7B",X"F7",
		X"07",X"F5",X"AB",X"F2",X"61",X"F0",X"2E",X"EE",X"0A",X"EC",X"FD",X"E9",X"FF",X"E7",X"14",X"E6",
		X"39",X"E4",X"71",X"E2",X"B8",X"E0",X"0F",X"DF",X"73",X"DD",X"E7",X"DB",X"68",X"DA",X"FA",X"D8",
		X"96",X"D7",X"40",X"D6",X"F7",X"D4",X"BA",X"D3",X"89",X"D2",X"63",X"D1",X"48",X"D0",X"38",X"CF",
		X"33",X"CE",X"37",X"CD",X"45",X"CC",X"5D",X"CB",X"7F",X"CA",X"A7",X"C9",X"DC",X"C8",X"15",X"C8",
		X"59",X"C7",X"A3",X"C6",X"F7",X"C5",X"52",X"C5",X"B0",X"C4",X"19",X"C4",X"88",X"C3",X"FE",X"C2",
		X"7A",X"C2",X"FB",X"C1",X"82",X"C1",X"11",X"C1",X"A4",X"C0",X"3B",X"C0",X"DA",X"BF",X"7D",X"BF",
		X"25",X"BF",X"D2",X"BE",X"82",X"BE",X"38",X"BE",X"F2",X"BD",X"B0",X"BD",X"71",X"BD",X"37",X"BD",
		X"00",X"BD",X"CE",X"BC",X"9F",X"BC",X"74",X"BC",X"4C",X"BC",X"26",X"BC",X"05",X"BC",X"E7",X"BB",
		X"CA",X"BB",X"B2",X"BB",X"9B",X"BB",X"87",X"BB",X"77",X"BB",X"68",X"BB",X"5C",X"BB",X"53",X"BB",
		X"4C",X"BB",X"46",X"BB",X"42",X"BB",X"42",X"BB",X"42",X"BB",X"45",X"BB",X"4A",X"BB",X"52",X"BB",
		X"58",X"BB",X"63",X"BB",X"6C",X"BB",X"7B",X"BB",X"8A",X"BB",X"99",X"BB",X"AA",X"BB",X"BE",X"BB",
		X"D1",X"BB",X"E7",X"BB",X"FD",X"BB",X"14",X"BC",X"2C",X"BC",X"47",X"BC",X"62",X"BC",X"7D",X"BC",
		X"9B",X"BC",X"B8",X"BC",X"D8",X"BC",X"F7",X"BC",X"19",X"BD",X"39",X"BD",X"5C",X"BD",X"7F",X"BD",
		X"A2",X"BD",X"C7",X"BD",X"EB",X"BD",X"11",X"BE",X"37",X"BE",X"5E",X"BE",X"85",X"BE",X"AE",X"BE",
		X"D7",X"BE",X"FE",X"BE",X"29",X"BF",X"51",X"BF",X"7E",X"BF",X"A8",X"BF",X"D4",X"BF",X"00",X"C0",
		X"2B",X"C0",X"58",X"C0",X"85",X"C0",X"B2",X"C0",X"DF",X"C0",X"0E",X"C1",X"3C",X"C1",X"6A",X"C1",
		X"98",X"C1",X"C8",X"C1",X"F6",X"C1",X"26",X"C2",X"55",X"C2",X"86",X"C2",X"B5",X"C2",X"E4",X"C2",
		X"14",X"C3",X"44",X"C3",X"75",X"C3",X"A5",X"C3",X"D7",X"C3",X"08",X"C4",X"39",X"C4",X"6A",X"C4",
		X"9B",X"C4",X"CD",X"C4",X"FF",X"C4",X"2E",X"C5",X"60",X"C5",X"92",X"C5",X"C3",X"C5",X"F4",X"C5",
		X"26",X"C6",X"5A",X"C6",X"8A",X"C6",X"BC",X"C6",X"ED",X"C6",X"22",X"C7",X"50",X"C7",X"84",X"C7",
		X"B4",X"C7",X"E8",X"C7",X"15",X"C8",X"4D",X"C8",X"78",X"C8",X"98",X"C9",X"22",X"CC",X"7D",X"CF",
		X"6D",X"D3",X"A8",X"D7",X"17",X"DC",X"94",X"E0",X"17",X"E5",X"89",X"E9",X"EE",X"ED",X"35",X"F2",
		X"64",X"F6",X"74",X"FA",X"68",X"FE",X"3C",X"02",X"F2",X"05",X"87",X"09",X"01",X"0D",X"5D",X"10",
		X"9C",X"13",X"BF",X"16",X"C8",X"19",X"B4",X"1C",X"8A",X"1F",X"43",X"22",X"E8",X"24",X"73",X"27",
		X"E8",X"29",X"48",X"2C",X"90",X"2E",X"C6",X"30",X"E6",X"32",X"F2",X"34",X"ED",X"36",X"D4",X"38",
		X"AA",X"3A",X"70",X"3C",X"23",X"3E",X"C6",X"3F",X"5A",X"41",X"DE",X"42",X"54",X"44",X"BD",X"45",
		X"15",X"47",X"64",X"48",X"A1",X"49",X"D5",X"4A",X"F9",X"4B",X"17",X"4D",X"23",X"4E",X"29",X"4F",
		X"1D",X"50",X"12",X"51",X"ED",X"51",X"D5",X"52",X"E8",X"52",X"7B",X"51",X"25",X"4F",X"2C",X"4C",
		X"D5",X"48",X"42",X"45",X"93",X"41",X"DA",X"3D",X"22",X"3A",X"76",X"36",X"DB",X"32",X"53",X"2F",
		X"E2",X"2B",X"89",X"28",X"48",X"25",X"21",X"22",X"10",X"1F",X"18",X"1C",X"39",X"19",X"73",X"16",
		X"C2",X"13",X"27",X"11",X"A0",X"0E",X"33",X"0C",X"D6",X"09",X"8F",X"07",X"56",X"05",X"53",X"03",
		X"B0",X"02",X"58",X"03",X"C9",X"04",X"C9",X"06",X"1A",X"09",X"A1",X"0B",X"42",X"0E",X"F0",X"10",
		X"9D",X"13",X"43",X"16",X"DE",X"18",X"6A",X"1B",X"E4",X"1D",X"4E",X"20",X"A2",X"22",X"E7",X"24",
		X"15",X"27",X"32",X"29",X"3A",X"2B",X"32",X"2D",X"19",X"2F",X"EE",X"30",X"B1",X"32",X"64",X"34",
		X"08",X"36",X"9D",X"37",X"21",X"39",X"99",X"3A",X"00",X"3C",X"5C",X"3D",X"A9",X"3E",X"EA",X"3F",
		X"1D",X"41",X"46",X"42",X"64",X"43",X"75",X"44",X"7A",X"45",X"75",X"46",X"66",X"47",X"4E",X"48",
		X"2B",X"49",X"00",X"4A",X"CA",X"4A",X"8C",X"4B",X"45",X"4C",X"F6",X"4C",X"A1",X"4D",X"41",X"4E",
		X"D9",X"4E",X"6C",X"4F",X"F8",X"4F",X"7C",X"50",X"FB",X"50",X"71",X"51",X"D7",X"51",X"08",X"51",
		X"E6",X"4E",X"FA",X"4B",X"83",X"48",X"C2",X"44",X"CF",X"40",X"CB",X"3C",X"C4",X"38",X"C5",X"34",
		X"D4",X"30",X"F8",X"2C",X"35",X"29",X"89",X"25",X"F9",X"21",X"82",X"1E",X"26",X"1B",X"E8",X"17",
		X"C2",X"14",X"B4",X"11",X"C0",X"0E",X"E5",X"0B",X"25",X"09",X"76",X"06",X"E4",X"03",X"60",X"01",
		X"FE",X"FE",X"9B",X"FC",X"C3",X"FA",X"78",X"FA",X"43",X"FB",X"C9",X"FC",X"C3",X"FE",X"0B",X"01",
		X"7E",X"03",X"0A",X"06",X"9D",X"08",X"2F",X"0B",X"B8",X"0D",X"39",X"10",X"A6",X"12",X"07",X"15",
		X"54",X"17",X"90",X"19",X"B7",X"1B",X"D0",X"1D",X"D5",X"1F",X"C9",X"21",X"AB",X"23",X"7F",X"25",
		X"3E",X"27",X"F1",X"28",X"90",X"2A",X"26",X"2C",X"A4",X"2D",X"1E",X"2F",X"7E",X"2F",X"6F",X"2E",
		X"89",X"2C",X"05",X"2A",X"2B",X"27",X"16",X"24",X"E7",X"20",X"A9",X"1D",X"6F",X"1A",X"3C",X"17",
		X"1A",X"14",X"06",X"11",X"08",X"0E",X"1F",X"0B",X"4C",X"08",X"8F",X"05",X"E7",X"02",X"56",X"00",
		X"D9",X"FD",X"71",X"FB",X"1B",X"F9",X"DE",X"F6",X"B0",X"F4",X"98",X"F2",X"8D",X"F0",X"9E",X"EE",
		X"AC",X"EC",X"25",X"EB",X"07",X"EB",X"F7",X"EB",X"D7",X"ED",X"2F",X"F0",X"D8",X"F2",X"AA",X"F5",
		X"95",X"F8",X"88",X"FB",X"78",X"FE",X"5D",X"01",X"35",X"04",X"FD",X"06",X"AF",X"09",X"50",X"0C",
		X"DC",X"0E",X"55",X"11",X"B5",X"13",X"06",X"16",X"40",X"18",X"69",X"1A",X"7C",X"1C",X"7F",X"1E",
		X"6F",X"20",X"50",X"22",X"1F",X"24",X"DB",X"25",X"88",X"27",X"27",X"29",X"B8",X"2A",X"3A",X"2C",
		X"AA",X"2D",X"11",X"2F",X"68",X"30",X"B5",X"31",X"F1",X"32",X"25",X"34",X"4B",X"35",X"66",X"36",
		X"78",X"37",X"7D",X"38",X"78",X"39",X"6A",X"3A",X"52",X"3B",X"30",X"3C",X"03",X"3D",X"D1",X"3D",
		X"95",X"3E",X"50",X"3F",X"02",X"40",X"AE",X"40",X"54",X"41",X"EF",X"41",X"85",X"42",X"14",X"43",
		X"9B",X"43",X"1D",X"44",X"98",X"44",X"0C",X"45",X"7D",X"45",X"E6",X"45",X"4A",X"46",X"AA",X"46",
		X"03",X"47",X"57",X"47",X"A8",X"47",X"F1",X"47",X"38",X"48",X"7B",X"48",X"B8",X"48",X"F1",X"48",
		X"27",X"49",X"58",X"49",X"87",X"49",X"B3",X"49",X"D8",X"49",X"FB",X"49",X"1A",X"4A",X"37",X"4A",
		X"50",X"4A",X"68",X"4A",X"7D",X"4A",X"76",X"4A",X"27",X"49",X"90",X"46",X"38",X"43",X"5D",X"3F",
		X"3C",X"3B",X"EE",X"36",X"94",X"32",X"3A",X"2E",X"EC",X"29",X"AF",X"25",X"8D",X"21",X"84",X"1D",
		X"95",X"19",X"C5",X"15",X"11",X"12",X"7A",X"0E",X"00",X"0B",X"A4",X"07",X"62",X"04",X"3C",X"01",
		X"32",X"FE",X"42",X"FB",X"67",X"F8",X"A9",X"F5",X"FB",X"F2",X"72",X"F0",X"E8",X"ED",X"09",X"EC",
		X"BD",X"EB",X"7E",X"EC",X"F7",X"ED",X"E5",X"EF",X"21",X"F2",X"84",X"F4",X"00",X"F7",X"83",X"F9",
		X"06",X"FC",X"82",X"FE",X"F4",X"00",X"55",X"03",X"A8",X"05",X"EB",X"07",X"1D",X"0A",X"3B",X"0C",
		X"4B",X"0E",X"46",X"10",X"33",X"12",X"0C",X"14",X"D9",X"15",X"92",X"17",X"40",X"19",X"DB",X"1A",
		X"6A",X"1C",X"E9",X"1D",X"54",X"1F",X"8E",X"1F",X"60",X"1E",X"62",X"1C",X"CB",X"19",X"E0",X"16",
		X"BC",X"13",X"82",X"10",X"39",X"0D",X"F8",X"09",X"BC",X"06",X"93",X"03",X"7A",X"00",X"78",X"FD",
		X"8A",X"FA",X"B3",X"F7",X"F1",X"F4",X"47",X"F2",X"B1",X"EF",X"33",X"ED",X"CA",X"EA",X"75",X"E8",
		X"35",X"E6",X"09",X"E4",X"EF",X"E1",X"EA",X"DF",X"F3",X"DD",X"13",X"DC",X"40",X"DA",X"7F",X"D8",
		X"CE",X"D6",X"2A",X"D5",X"99",X"D3",X"14",X"D2",X"9D",X"D0",X"36",X"CF",X"DB",X"CD",X"8D",X"CC",
		X"4C",X"CB",X"17",X"CA",X"EE",X"C8",X"CE",X"C7",X"BB",X"C6",X"B4",X"C5",X"B5",X"C4",X"C1",X"C3",
		X"D8",X"C2",X"F8",X"C1",X"1F",X"C1",X"52",X"C0",X"8B",X"BF",X"D0",X"BE",X"19",X"BE",X"6C",X"BD",
		X"C5",X"BC",X"28",X"BC",X"90",X"BB",X"FF",X"BA",X"76",X"BA",X"F2",X"B9",X"77",X"B9",X"FF",X"B8",
		X"8D",X"B8",X"22",X"B8",X"BC",X"B7",X"5D",X"B7",X"01",X"B7",X"AC",X"B6",X"5B",X"B6",X"10",X"B6",
		X"C6",X"B5",X"83",X"B5",X"44",X"B5",X"0B",X"B5",X"D2",X"B4",X"A0",X"B4",X"70",X"B4",X"44",X"B4",
		X"1D",X"B4",X"F9",X"B3",X"D7",X"B3",X"BB",X"B3",X"9A",X"B3",X"BF",X"B3",X"53",X"B5",X"0E",X"B8",
		X"7C",X"BB",X"62",X"BF",X"87",X"C3",X"D1",X"C7",X"27",X"CC",X"7A",X"D0",X"C1",X"D4",X"F3",X"D8",
		X"0C",X"DD",X"0D",X"E1",X"EF",X"E4",X"B6",X"E8",X"5F",X"EC",X"EC",X"EF",X"5C",X"F3",X"AE",X"F6",
		X"E6",X"F9",X"05",X"FD",X"07",X"00",X"F0",X"02",X"C0",X"05",X"78",X"08",X"1A",X"0B",X"A3",X"0D",
		X"17",X"10",X"77",X"12",X"C0",X"14",X"F6",X"16",X"17",X"19",X"29",X"1B",X"24",X"1D",X"0E",X"1F",
		X"E8",X"20",X"B2",X"22",X"6A",X"24",X"14",X"26",X"AE",X"27",X"3B",X"29",X"B5",X"2A",X"25",X"2C",
		X"84",X"2D",X"DA",X"2E",X"21",X"30",X"5C",X"31",X"8B",X"32",X"AE",X"33",X"C8",X"34",X"D7",X"35",
		X"D8",X"36",X"D1",X"37",X"C0",X"38",X"A8",X"39",X"62",X"3A",X"BC",X"39",X"D7",X"37",X"2C",X"35",
		X"00",X"32",X"87",X"2E",X"E2",X"2A",X"2A",X"27",X"6E",X"23",X"B8",X"1F",X"12",X"1C",X"7F",X"18",
		X"03",X"15",X"9D",X"11",X"51",X"0E",X"1D",X"0B",X"03",X"08",X"02",X"05",X"19",X"02",X"47",X"FF",
		X"90",X"FC",X"EC",X"F9",X"63",X"F7",X"EB",X"F4",X"8F",X"F2",X"3C",X"F0",X"0D",X"EE",X"D9",X"EB",
		X"64",X"EA",X"7E",X"EA",X"99",X"EB",X"68",X"ED",X"A3",X"EF",X"26",X"F2",X"CE",X"F4",X"8F",X"F7",
		X"51",X"FA",X"12",X"FD",X"C7",X"FF",X"72",X"02",X"0A",X"05",X"91",X"07",X"05",X"0A",X"69",X"0C",
		X"B6",X"0E",X"F3",X"10",X"1A",X"13",X"31",X"15",X"33",X"17",X"27",X"19",X"08",X"1B",X"DA",X"1C",
		X"97",X"1E",X"4A",X"20",X"E9",X"21",X"6E",X"23",X"AC",X"23",X"8F",X"22",X"9F",X"20",X"1F",X"1E",
		X"49",X"1B",X"3F",X"18",X"1B",X"15",X"ED",X"11",X"C2",X"0E",X"9E",X"0B",X"8A",X"08",X"87",X"05",
		X"9A",X"02",X"C0",X"FF",X"FD",X"FC",X"4F",X"FA",X"B7",X"F7",X"35",X"F5",X"C4",X"F2",X"6C",X"F0",
		X"26",X"EE",X"F7",X"EB",X"D6",X"E9",X"CF",X"E7",X"D1",X"E5",X"EE",X"E3",X"0A",X"E2",X"B5",X"E0",
		X"EE",X"E0",X"36",X"E2",X"3C",X"E4",X"AF",X"E6",X"70",X"E9",X"53",X"EC",X"51",X"EF",X"50",X"F2",
		X"4D",X"F5",X"3C",X"F8",X"20",X"FB",X"F1",X"FD",X"AF",X"00",X"57",X"03",X"ED",X"05",X"6D",X"08",
		X"DA",X"0A",X"30",X"0D",X"77",X"0F",X"A6",X"11",X"C5",X"13",X"CE",X"15",X"C8",X"17",X"AD",X"19",
		X"88",X"1B",X"49",X"1D",X"FF",X"1E",X"94",X"1F",X"B5",X"1E",X"FF",X"1C",X"A9",X"1A",X"FC",X"17",
		X"10",X"15",X"0D",X"12",X"F9",X"0E",X"E7",X"0B",X"DA",X"08",X"DF",X"05",X"EE",X"02",X"16",X"00",
		X"50",X"FD",X"A1",X"FA",X"05",X"F8",X"7E",X"F5",X"0D",X"F3",X"B0",X"F0",X"65",X"EE",X"2F",X"EC",
		X"0E",X"EA",X"FF",X"E7",X"01",X"E6",X"15",X"E4",X"3A",X"E2",X"70",X"E0",X"B5",X"DE",X"0B",X"DD",
		X"71",X"DB",X"E3",X"D9",X"66",X"D8",X"F5",X"D6",X"92",X"D5",X"3C",X"D4",X"F3",X"D2",X"B6",X"D1",
		X"84",X"D0",X"5E",X"CF",X"45",X"CE",X"32",X"CD",X"31",X"CC",X"32",X"CB",X"43",X"CA",X"58",X"C9",
		X"7C",X"C8",X"A5",X"C7",X"D9",X"C6",X"12",X"C6",X"5A",X"C5",X"A2",X"C4",X"FA",X"C3",X"4D",X"C3",
		X"B8",X"C2",X"15",X"C2",X"97",X"C1",X"DC",X"C0",X"D4",X"BF",X"60",X"BF",X"E1",X"BE",X"72",X"BE",
		X"03",X"BE",X"9D",X"BD",X"3A",X"BD",X"DE",X"BC",X"85",X"BC",X"31",X"BC",X"E2",X"BB",X"99",X"BB",
		X"52",X"BB",X"11",X"BB",X"D4",X"BA",X"9A",X"BA",X"65",X"BA",X"32",X"BA",X"04",X"BA",X"DA",X"B9",
		X"B2",X"B9",X"8F",X"B9",X"6E",X"B9",X"4F",X"B9",X"36",X"B9",X"1C",X"B9",X"08",X"B9",X"F6",X"B8",
		X"E5",X"B8",X"D7",X"B8",X"CD",X"B8",X"C5",X"B8",X"C0",X"B8",X"BA",X"B8",X"B8",X"B8",X"B9",X"B8",
		X"BB",X"B8",X"BE",X"B8",X"C4",X"B8",X"CE",X"B8",X"D5",X"B8",X"E1",X"B8",X"EF",X"B8",X"FE",X"B8",
		X"0C",X"B9",X"1F",X"B9",X"30",X"B9",X"47",X"B9",X"5A",X"B9",X"74",X"B9",X"87",X"B9",X"A8",X"B9",
		X"B4",X"B9",X"83",X"BA",X"D2",X"BC",X"0D",X"C0",X"E9",X"C3",X"1E",X"C8",X"8A",X"CC",X"0C",X"D1",
		X"96",X"D5",X"14",X"DA",X"81",X"DE",X"D9",X"E2",X"15",X"E7",X"34",X"EB",X"34",X"EF",X"19",X"F3",
		X"DB",X"F6",X"82",X"FA",X"0A",X"FE",X"73",X"01",X"C1",X"04",X"F3",X"07",X"08",X"0B",X"06",X"0E",
		X"E5",X"10",X"B2",X"13",X"5C",X"16",X"03",X"19",X"F8",X"1A",X"53",X"1B",X"A0",X"1A",X"32",X"19",
		X"52",X"17",X"22",X"15",X"CB",X"12",X"59",X"10",X"DE",X"0D",X"63",X"0B",X"F1",X"08",X"87",X"06",
		X"2B",X"04",X"DE",X"01",X"A5",X"FF",X"79",X"FD",X"5E",X"FB",X"56",X"F9",X"5F",X"F7",X"76",X"F5",
		X"9F",X"F3",X"D6",X"F1",X"21",X"F0",X"76",X"EE",X"DB",X"EC",X"4F",X"EB",X"D3",X"E9",X"6A",X"E8",
		X"3E",X"E8",X"76",X"E9",X"83",X"EB",X"26",X"EE",X"1D",X"F1",X"4B",X"F4",X"91",X"F7",X"E4",X"FA",
		X"2F",X"FE",X"73",X"01",X"A4",X"04",X"C5",X"07",X"D2",X"0A",X"C5",X"0D",X"A4",X"10",X"6A",X"13",
		X"1B",X"16",X"B5",X"18",X"38",X"1B",X"A6",X"1D",X"FF",X"1F",X"41",X"22",X"71",X"24",X"8B",X"26",
		X"98",X"28",X"89",X"2A",X"7A",X"2C",X"E6",X"2D",X"C3",X"2D",X"86",X"2C",X"89",X"2A",X"17",X"28",
		X"57",X"25",X"6D",X"22",X"6E",X"1F",X"69",X"1C",X"68",X"19",X"70",X"16",X"86",X"13",X"AD",X"10",
		X"E8",X"0D",X"38",X"0B",X"99",X"08",X"12",X"06",X"9D",X"03",X"3E",X"01",X"F0",X"FE",X"B9",X"FC",
		X"90",X"FA",X"7E",X"F8",X"7A",X"F6",X"8C",X"F4",X"AA",X"F2",X"DE",X"F0",X"1A",X"EF",X"6F",X"EE",
		X"3E",X"EF",X"ED",X"F0",X"3E",X"F3",X"EA",X"F5",X"D4",X"F8",X"D9",X"FB",X"EE",X"FE",X"01",X"02",
		X"0F",X"05",X"0E",X"08",X"FC",X"0A",X"D6",X"0D",X"9C",X"10",X"4C",X"13",X"E8",X"15",X"6F",X"18",
		X"DF",X"1A",X"3B",X"1D",X"83",X"1F",X"B7",X"21",X"D7",X"23",X"E4",X"25",X"DD",X"27",X"C7",X"29",
		X"9B",X"2B",X"69",X"2D",X"DB",X"2E",X"CC",X"2E",X"8C",X"2D",X"87",X"2B",X"04",X"29",X"32",X"26",
		X"32",X"23",X"1B",X"20",X"FF",X"1C",X"E4",X"19",X"D3",X"16",X"D2",X"13",X"E3",X"10",X"07",X"0E",
		X"3E",X"0B",X"8D",X"08",X"EE",X"05",X"64",X"03",X"F2",X"00",X"93",X"FE",X"46",X"FC",X"0E",X"FA",
		X"EB",X"F7",X"D6",X"F5",X"D6",X"F3",X"E4",X"F1",X"0C",X"F0",X"33",X"EE",X"46",X"ED",X"E5",X"ED",
		X"6F",X"EF",X"A8",X"F1",X"3E",X"F4",X"1A",X"F7",X"12",X"FA",X"1D",X"FD",X"26",X"00",X"2C",X"03",
		X"24",X"06",X"0C",X"09",X"E1",X"0B",X"A3",X"0E",X"4F",X"11",X"E7",X"13",X"6A",X"16",X"D7",X"18",
		X"2D",X"1B",X"73",X"1D",X"A2",X"1F",X"C1",X"21",X"C9",X"23",X"C1",X"25",X"A7",X"27",X"7C",X"29",
		X"41",X"2B",X"F3",X"2C",X"98",X"2E",X"2D",X"30",X"B2",X"31",X"2A",X"33",X"94",X"34",X"EF",X"35",
		X"3E",X"37",X"80",X"38",X"B6",X"39",X"DF",X"3A",X"FE",X"3B",X"10",X"3D",X"19",X"3E",X"16",X"3F",
		X"0A",X"40",X"F0",X"40",X"D2",X"41",X"A7",X"42",X"77",X"43",X"38",X"44",X"F9",X"44",X"A9",X"45",
		X"59",X"46",X"F8",X"46",X"9C",X"47",X"29",X"48",X"C6",X"48",X"A8",X"48",X"05",X"47",X"6A",X"44",
		X"26",X"41",X"83",X"3D",X"A0",X"39",X"A3",X"35",X"9B",X"31",X"95",X"2D",X"9D",X"29",X"BA",X"25",
		X"EB",X"21",X"37",X"1E",X"9B",X"1A",X"1B",X"17",X"B6",X"13",X"6A",X"10",X"3B",X"0D",X"24",X"0A",
		X"28",X"07",X"46",X"04",X"79",X"01",X"C8",X"FE",X"2B",X"FC",X"A5",X"F9",X"35",X"F7",X"DA",X"F4",
		X"92",X"F2",X"5F",X"F0",X"40",X"EE",X"32",X"EC",X"37",X"EA",X"4E",X"E8",X"74",X"E6",X"AC",X"E4",
		X"F4",X"E2",X"4B",X"E1",X"B2",X"DF",X"26",X"DE",X"AA",X"DC",X"39",X"DB",X"D7",X"D9",X"82",X"D8",
		X"3A",X"D7",X"FD",X"D5",X"CC",X"D4",X"A6",X"D3",X"8A",X"D2",X"7B",X"D1",X"76",X"D0",X"7B",X"CF",
		X"8A",X"CE",X"9F",X"CD",X"C1",X"CC",X"EA",X"CB",X"1C",X"CB",X"58",X"CA",X"9B",X"C9",X"E5",X"C8",
		X"37",X"C8",X"91",X"C7",X"F2",X"C6",X"59",X"C6",X"C8",X"C5",X"3C",X"C5",X"B8",X"C4",X"39",X"C4",
		X"C0",X"C3",X"4C",X"C3",X"E0",X"C2",X"77",X"C2",X"14",X"C2",X"B6",X"C1",X"5B",X"C1",X"08",X"C1",
		X"B8",X"C0",X"6D",X"C0",X"26",X"C0",X"E3",X"BF",X"A5",X"BF",X"6A",X"BF",X"32",X"BF",X"FF",X"BE",
		X"D0",X"BE",X"A4",X"BE",X"79",X"BE",X"54",X"BE",X"30",X"BE",X"10",X"BE",X"F3",X"BD",X"DA",X"BD",
		X"C3",X"BD",X"AE",X"BD",X"9C",X"BD",X"8B",X"BD",X"7E",X"BD",X"74",X"BD",X"6A",X"BD",X"66",X"BD",
		X"60",X"BD",X"5F",X"BD",X"5C",X"BD",X"60",X"BD",X"61",X"BD",X"69",X"BD",X"6D",X"BD",X"79",X"BD",
		X"7F",X"BD",X"90",X"BD",X"93",X"BD",X"F6",X"BD",X"D5",X"BF",X"C9",X"C2",X"71",X"C6",X"87",X"CA",
		X"DC",X"CE",X"4F",X"D3",X"CD",X"D7",X"46",X"DC",X"AF",X"E0",X"04",X"E5",X"3D",X"E9",X"5D",X"ED",
		X"5D",X"F1",X"40",X"F5",X"03",X"F9",X"AA",X"FC",X"32",X"00",X"9C",X"03",X"EA",X"06",X"1C",X"0A",
		X"32",X"0D",X"2E",X"10",X"11",X"13",X"D8",X"15",X"8C",X"18",X"23",X"1B",X"A6",X"1D",X"14",X"20",
		X"6C",X"22",X"AB",X"24",X"D9",X"26",X"F3",X"28",X"F9",X"2A",X"EE",X"2C",X"D1",X"2E",X"A2",X"30",
		X"62",X"32",X"10",X"34",X"B4",X"35",X"42",X"37",X"C6",X"38",X"35",X"3A",X"9F",X"3B",X"F3",X"3C",
		X"41",X"3E",X"7C",X"3F",X"B0",X"40",X"D2",X"41",X"F0",X"42",X"F9",X"43",X"03",X"45",X"F6",X"45",
		X"EA",X"46",X"C9",X"47",X"AE",X"48",X"6E",X"49",X"6E",X"4A",X"CE",X"4B",X"77",X"4C",X"32",X"4D",
		X"D5",X"4D",X"79",X"4E",X"10",X"4F",X"A5",X"4F",X"2F",X"50",X"B4",X"50",X"31",X"51",X"A9",X"51",
		X"1A",X"52",X"85",X"52",X"E9",X"52",X"49",X"53",X"A2",X"53",X"F7",X"53",X"46",X"54",X"91",X"54",
		X"D6",X"54",X"17",X"55",X"54",X"55",X"8B",X"55",X"BF",X"55",X"ED",X"55",X"1A",X"56",X"41",X"56",
		X"65",X"56",X"84",X"56",X"A0",X"56",X"B9",X"56",X"CF",X"56",X"E3",X"56",X"F4",X"56",X"FF",X"56",
		X"08",X"57",X"0F",X"57",X"15",X"57",X"15",X"57",X"16",X"57",X"12",X"57",X"0E",X"57",X"05",X"57",
		X"FB",X"56",X"EE",X"56",X"E1",X"56",X"D0",X"56",X"BE",X"56",X"AA",X"56",X"94",X"56",X"7C",X"56",
		X"65",X"56",X"48",X"56",X"2C",X"56",X"0F",X"56",X"EF",X"55",X"CE",X"55",X"AC",X"55",X"89",X"55",
		X"65",X"55",X"3F",X"55",X"19",X"55",X"F0",X"54",X"C7",X"54",X"9C",X"54",X"72",X"54",X"45",X"54",
		X"15",X"54",X"E9",X"53",X"BA",X"53",X"8A",X"53",X"5B",X"53",X"28",X"53",X"F7",X"52",X"C3",X"52",
		X"90",X"52",X"5C",X"52",X"27",X"52",X"F3",X"51",X"BC",X"51",X"86",X"51",X"4F",X"51",X"17",X"51",
		X"DF",X"50",X"A8",X"50",X"6D",X"50",X"35",X"50",X"FA",X"4F",X"C2",X"4F",X"86",X"4F",X"4C",X"4F",
		X"10",X"4F",X"D5",X"4E",X"98",X"4E",X"5D",X"4E",X"20",X"4E",X"E5",X"4D",X"A8",X"4D",X"6C",X"4D",
		X"2D",X"4D",X"F0",X"4C",X"B1",X"4C",X"76",X"4C",X"35",X"4C",X"FB",X"4B",X"B6",X"4B",X"86",X"4B",
		X"DA",X"4A",X"A8",X"48",X"6D",X"45",X"83",X"41",X"33",X"3D",X"A5",X"38",X"FC",X"33",X"4B",X"2F",
		X"A1",X"2A",X"0B",X"26",X"88",X"21",X"21",X"1D",X"DA",X"18",X"B0",X"14",X"A7",X"10",X"BB",X"0C",
		X"F0",X"08",X"43",X"05",X"B5",X"01",X"46",X"FE",X"F3",X"FA",X"B9",X"F7",X"A1",X"F4",X"9E",X"F1",
		X"B9",X"EE",X"E7",X"EB",X"36",X"E9",X"96",X"E6",X"1F",X"E5",X"2B",X"E5",X"1D",X"E6",X"BA",X"E7",
		X"B6",X"E9",X"F8",X"EB",X"5A",X"EE",X"D3",X"F0",X"4F",X"F3",X"CA",X"F5",X"3B",X"F8",X"A3",X"FA",
		X"FB",X"FC",X"42",X"FF",X"7A",X"01",X"9F",X"03",X"B5",X"05",X"BA",X"07",X"AE",X"09",X"91",X"0B",
		X"64",X"0D",X"27",X"0F",X"DA",X"10",X"7D",X"12",X"16",X"14",X"99",X"15",X"1D",X"17",X"40",X"18",
		X"DC",X"17",X"4E",X"16",X"FB",X"13",X"30",X"11",X"17",X"0E",X"D3",X"0A",X"79",X"07",X"1F",X"04",
		X"C9",X"00",X"7F",X"FD",X"47",X"FA",X"22",X"F7",X"13",X"F4",X"1D",X"F1",X"3C",X"EE",X"74",X"EB",
		X"C1",X"E8",X"27",X"E6",X"A0",X"E3",X"32",X"E1",X"D6",X"DE",X"93",X"DC",X"5F",X"DA",X"45",X"D8",
		X"36",X"D6",X"44",X"D4",X"55",X"D2",X"5E",X"D1",X"F5",X"D1",X"77",X"D3",X"A8",X"D5",X"3B",X"D8",
		X"12",X"DB",X"07",X"DE",X"11",X"E1",X"1B",X"E4",X"21",X"E7",X"17",X"EA",X"02",X"ED",X"D8",X"EF",
		X"9B",X"F2",X"4A",X"F5",X"E6",X"F7",X"6C",X"FA",X"DF",X"FC",X"3B",X"FF",X"85",X"01",X"BC",X"03",
		X"DE",X"05",X"EF",X"07",X"F1",X"09",X"DF",X"0B",X"B9",X"0D",X"8C",X"0F",X"1C",X"11",X"39",X"11",
		X"0E",X"10",X"1A",X"0E",X"9F",X"0B",X"D0",X"08",X"D1",X"05",X"BC",X"02",X"9D",X"FF",X"83",X"FC",
		X"6F",X"F9",X"6E",X"F6",X"7B",X"F3",X"9F",X"F0",X"D7",X"ED",X"24",X"EB",X"87",X"E8",X"01",X"E6",
		X"8E",X"E3",X"31",X"E1",X"E8",X"DE",X"B7",X"DC",X"94",X"DA",X"88",X"D8",X"8D",X"D6",X"A4",X"D4",
		X"CC",X"D2",X"06",X"D1",X"4E",X"CF",X"A9",X"CD",X"10",X"CC",X"8A",X"CA",X"0F",X"C9",X"A5",X"C7",
		X"45",X"C6",X"F7",X"C4",X"B1",X"C3",X"7A",X"C2",X"4E",X"C1",X"30",X"C0",X"1C",X"BF",X"12",X"BE",
		X"12",X"BD",X"20",X"BC",X"36",X"BB",X"54",X"BA",X"7C",X"B9",X"AF",X"B8",X"E8",X"B7",X"2A",X"B7",
		X"77",X"B6",X"CB",X"B5",X"25",X"B5",X"88",X"B4",X"F1",X"B3",X"78",X"B3",X"4D",X"B4",X"78",X"B6",
		X"6C",X"B9",X"ED",X"BC",X"B7",X"C0",X"B4",X"C4",X"BF",X"C8",X"D1",X"CC",X"D9",X"D0",X"D1",X"D4",
		X"B3",X"D8",X"81",X"DC",X"31",X"E0",X"C7",X"E3",X"43",X"E7",X"A5",X"EA",X"E9",X"ED",X"16",X"F1",
		X"25",X"F4",X"1E",X"F7",X"FC",X"F9",X"C3",X"FC",X"71",X"FF",X"09",X"02",X"8A",X"04",X"F7",X"06",
		X"4D",X"09",X"8F",X"0B",X"BF",X"0D",X"DC",X"0F",X"E4",X"11",X"DF",X"13",X"C3",X"15",X"9B",X"17",
		X"5E",X"19",X"15",X"1B",X"BA",X"1C",X"53",X"1E",X"D9",X"1F",X"54",X"21",X"C0",X"22",X"1F",X"24",
		X"72",X"25",X"B7",X"26",X"F4",X"27",X"22",X"29",X"46",X"2A",X"5F",X"2B",X"6C",X"2C",X"6F",X"2D",
		X"6A",X"2E",X"57",X"2F",X"41",X"30",X"1A",X"31",X"EB",X"31",X"8C",X"31",X"C3",X"2F",X"26",X"2D",
		X"F2",X"29",X"6C",X"26",X"AF",X"22",X"DF",X"1E",X"05",X"1B",X"35",X"17",X"70",X"13",X"BF",X"0F",
		X"23",X"0C",X"A2",X"08",X"38",X"05",X"E9",X"01",X"B6",X"FE",X"9B",X"FB",X"9A",X"F8",X"B2",X"F5",
		X"E4",X"F2",X"2C",X"F0",X"8D",X"ED",X"01",X"EB",X"91",X"E8",X"30",X"E6",X"ED",X"E3",X"AC",X"E1",
		X"E7",X"DF",X"B3",X"DF",X"A9",X"E0",X"60",X"E2",X"94",X"E4",X"19",X"E7",X"CB",X"E9",X"96",X"EC",
		X"68",X"EF",X"3A",X"F2",X"04",X"F5",X"C0",X"F7",X"6C",X"FA",X"06",X"FD",X"8E",X"FF",X"01",X"02",
		X"64",X"04",X"B0",X"06",X"EC",X"08",X"13",X"0B",X"29",X"0D",X"2E",X"0F",X"1F",X"11",X"00",X"13",
		X"D2",X"14",X"92",X"16",X"42",X"18",X"E3",X"19",X"76",X"1B",X"FC",X"1C",X"72",X"1E",X"DC",X"1F",
		X"3A",X"21",X"87",X"22",X"CC",X"23",X"04",X"25",X"31",X"26",X"51",X"27",X"67",X"28",X"73",X"29",
		X"74",X"2A",X"6C",X"2B",X"5B",X"2C",X"3F",X"2D",X"1C",X"2E",X"F0",X"2E",X"B8",X"2F",X"7D",X"30",
		X"37",X"31",X"EA",X"31",X"95",X"32",X"3A",X"33",X"D7",X"33",X"6E",X"34",X"FF",X"34",X"88",X"35",
		X"0C",X"36",X"89",X"36",X"01",X"37",X"74",X"37",X"E0",X"37",X"48",X"38",X"AA",X"38",X"09",X"39",
		X"60",X"39",X"B6",X"39",X"03",X"3A",X"50",X"3A",X"94",X"3A",X"D9",X"3A",X"17",X"3B",X"54",X"3B",
		X"88",X"3B",X"BE",X"3B",X"ED",X"3B",X"1D",X"3C",X"42",X"3C",X"6C",X"3C",X"8B",X"3C",X"B1",X"3C",
		X"C9",X"3C",X"E9",X"3C",X"FA",X"3C",X"1A",X"3D",X"1C",X"3D",X"5A",X"3D",X"EA",X"3D",X"EC",X"3D",
		X"FB",X"3D",X"FF",X"3D",X"07",X"3E",X"07",X"3E",X"0B",X"3E",X"09",X"3E",X"08",X"3E",X"03",X"3E",
		X"FE",X"3D",X"F7",X"3D",X"EE",X"3D",X"E3",X"3D",X"D7",X"3D",X"CB",X"3D",X"BD",X"3D",X"AB",X"3D",
		X"9A",X"3D",X"88",X"3D",X"73",X"3D",X"5F",X"3D",X"48",X"3D",X"34",X"3D",X"FB",X"3C",X"67",X"3B",
		X"8A",X"38",X"EE",X"34",X"CD",X"30",X"68",X"2C",X"D8",X"27",X"40",X"23",X"A5",X"1E",X"1B",X"1A",
		X"A5",X"15",X"4B",X"11",X"0A",X"0D",X"E9",X"08",X"E6",X"04",X"04",X"01",X"42",X"FD",X"9B",X"F9",
		X"13",X"F6",X"AC",X"F2",X"61",X"EF",X"2F",X"EC",X"1B",X"E9",X"21",X"E6",X"44",X"E3",X"79",X"E0",
		X"D2",X"DD",X"2E",X"DB",X"46",X"D9",X"02",X"D9",X"C9",X"D9",X"52",X"DB",X"4C",X"DD",X"95",X"DF",
		X"08",X"E2",X"97",X"E4",X"29",X"E7",X"C0",X"E9",X"4C",X"EC",X"CE",X"EE",X"42",X"F1",X"A7",X"F3",
		X"F9",X"F5",X"3B",X"F8",X"6C",X"FA",X"8B",X"FC",X"96",X"FE",X"93",X"00",X"7F",X"02",X"5A",X"04",
		X"24",X"06",X"E1",X"07",X"8E",X"09",X"2C",X"0B",X"BB",X"0C",X"3F",X"0E",X"B3",X"0F",X"1B",X"11",
		X"75",X"12",X"C4",X"13",X"08",X"15",X"3F",X"16",X"6C",X"17",X"8E",X"18",X"A7",X"19",X"B2",X"1A",
		X"B6",X"1B",X"AF",X"1C",X"A0",X"1D",X"87",X"1E",X"66",X"1F",X"3D",X"20",X"0C",X"21",X"D1",X"21",
		X"8F",X"22",X"48",X"23",X"F7",X"23",X"A2",X"24",X"43",X"25",X"DE",X"25",X"73",X"26",X"03",X"27",
		X"8C",X"27",X"10",X"28",X"8D",X"28",X"06",X"29",X"78",X"29",X"E7",X"29",X"4E",X"2A",X"B5",X"2A",
		X"12",X"2B",X"6E",X"2B",X"C2",X"2B",X"17",X"2C",X"64",X"2C",X"AE",X"2C",X"F6",X"2C",X"39",X"2D",
		X"76",X"2D",X"B4",X"2D",X"EA",X"2D",X"20",X"2E",X"50",X"2E",X"80",X"2E",X"AB",X"2E",X"D6",X"2E",
		X"F9",X"2E",X"1F",X"2F",X"3A",X"2F",X"63",X"2F",X"2D",X"2F",X"78",X"2D",X"9F",X"2A",X"10",X"27",
		X"0D",X"23",X"C8",X"1E",X"62",X"1A",X"F3",X"15",X"86",X"11",X"28",X"0D",X"E1",X"08",X"B0",X"04",
		X"9E",X"00",X"A9",X"FC",X"D2",X"F8",X"18",X"F5",X"7D",X"F1",X"01",X"EE",X"9F",X"EA",X"5D",X"E7",
		X"36",X"E4",X"2B",X"E1",X"39",X"DE",X"61",X"DB",X"A2",X"D8",X"FD",X"D5",X"6F",X"D3",X"F7",X"D0",
		X"97",X"CE",X"4C",X"CC",X"14",X"CA",X"F2",X"C7",X"E4",X"C5",X"E7",X"C3",X"FF",X"C1",X"28",X"C0",
		X"61",X"BE",X"AD",X"BC",X"08",X"BB",X"73",X"B9",X"EE",X"B7",X"76",X"B6",X"0F",X"B5",X"B6",X"B3",
		X"68",X"B2",X"29",X"B1",X"F6",X"AF",X"D1",X"AE",X"B6",X"AD",X"A8",X"AC",X"A4",X"AB",X"AC",X"AA",
		X"BF",X"A9",X"DB",X"A8",X"01",X"A8",X"31",X"A7",X"6A",X"A6",X"AD",X"A5",X"F8",X"A4",X"4C",X"A4",
		X"A7",X"A3",X"0C",X"A3",X"76",X"A2",X"EA",X"A1",X"63",X"A1",X"E6",X"A0",X"6D",X"A0",X"FC",X"9F",
		X"8F",X"9F",X"2D",X"9F",X"CD",X"9E",X"74",X"9E",X"1F",X"9E",X"D3",X"9D",X"89",X"9D",X"49",X"9D",
		X"06",X"9D",X"CF",X"9C",X"97",X"9C",X"6A",X"9C",X"39",X"9C",X"19",X"9C",X"E5",X"9B",X"7D",X"9C",
		X"A0",X"9E",X"B4",X"A1",X"70",X"A5",X"8A",X"A9",X"DF",X"AD",X"4A",X"B2",X"C0",X"B6",X"2C",X"BB",
		X"8A",X"BF",X"D1",X"C3",X"02",X"C8",X"14",X"CC",X"0C",X"D0",X"E5",X"D3",X"A0",X"D7",X"40",X"DB",
		X"C2",X"DE",X"27",X"E2",X"71",X"E5",X"9F",X"E8",X"B4",X"EB",X"AC",X"EE",X"8F",X"F1",X"58",X"F4",
		X"0B",X"F7",X"A6",X"F9",X"14",X"FC",X"18",X"FD",X"BB",X"FC",X"86",X"FB",X"B7",X"F9",X"91",X"F7",
		X"2F",X"F5",X"B0",X"F2",X"21",X"F0",X"8F",X"ED",X"03",X"EB",X"80",X"E8",X"0C",X"E6",X"A8",X"E3",
		X"54",X"E1",X"13",X"DF",X"E5",X"DC",X"C6",X"DA",X"BC",X"D8",X"C3",X"D6",X"DE",X"D4",X"06",X"D3",
		X"42",X"D1",X"8A",X"CF",X"E8",X"CD",X"4C",X"CC",X"CD",X"CA",X"45",X"C9",X"65",X"C8",X"1E",X"C9",
		X"E1",X"CA",X"5F",X"CD",X"4A",X"D0",X"7F",X"D3",X"D5",X"D6",X"3F",X"DA",X"AA",X"DD",X"0F",X"E1",
		X"66",X"E4",X"AD",X"E7",X"DC",X"EA",X"F8",X"ED",X"FC",X"F0",X"E9",X"F3",X"BF",X"F6",X"80",X"F9",
		X"28",X"FC",X"BB",X"FE",X"38",X"01",X"9F",X"03",X"F1",X"05",X"32",X"08",X"5D",X"0A",X"79",X"0C",
		X"7D",X"0E",X"6C",X"10",X"19",X"11",X"52",X"10",X"B0",X"0E",X"6E",X"0C",X"D5",X"09",X"FD",X"06",
		X"0A",X"04",X"07",X"01",X"09",X"FE",X"0D",X"FB",X"22",X"F8",X"42",X"F5",X"7A",X"F2",X"C4",X"EF",
		X"23",X"ED",X"95",X"EA",X"21",X"E8",X"BC",X"E5",X"6F",X"E3",X"34",X"E1",X"0F",X"DF",X"FA",X"DC",
		X"F9",X"DA",X"0A",X"D9",X"2D",X"D7",X"60",X"D5",X"A4",X"D3",X"F7",X"D1",X"5C",X"D0",X"CE",X"CE",
		X"4F",X"CD",X"DE",X"CB",X"7C",X"CA",X"26",X"C9",X"DD",X"C7",X"A0",X"C6",X"70",X"C5",X"4C",X"C4",
		X"33",X"C3",X"25",X"C2",X"22",X"C1",X"29",X"C0",X"3A",X"BF",X"54",X"BE",X"79",X"BD",X"A8",X"BC",
		X"DD",X"BB",X"1D",X"BB",X"64",X"BA",X"B2",X"B9",X"0A",X"B9",X"6B",X"B8",X"D0",X"B7",X"3E",X"B7",
		X"B2",X"B6",X"2C",X"B6",X"AD",X"B5",X"35",X"B5",X"C3",X"B4",X"57",X"B4",X"F1",X"B3",X"90",X"B3",
		X"35",X"B3",X"DD",X"B2",X"8C",X"B2",X"40",X"B2",X"F8",X"B1",X"B5",X"B1",X"76",X"B1",X"3A",X"B1",
		X"06",X"B1",X"D2",X"B0",X"A4",X"B0",X"79",X"B0",X"51",X"B0",X"2E",X"B0",X"0F",X"B0",X"F2",X"AF",
		X"D9",X"AF",X"C2",X"AF",X"AD",X"AF",X"9D",X"AF",X"8E",X"AF",X"84",X"AF",X"7C",X"AF",X"75",X"AF",
		X"71",X"AF",X"71",X"AF",X"72",X"AF",X"75",X"AF",X"7C",X"AF",X"83",X"AF",X"8C",X"AF",X"98",X"AF",
		X"A7",X"AF",X"B5",X"AF",X"C6",X"AF",X"DA",X"AF",X"EF",X"AF",X"02",X"B0",X"1B",X"B0",X"33",X"B0",
		X"51",X"B0",X"69",X"B0",X"88",X"B0",X"A3",X"B0",X"C7",X"B0",X"E3",X"B0",X"0D",X"B1",X"22",X"B1",
		X"18",X"B2",X"8E",X"B4",X"EF",X"B7",X"EE",X"BB",X"44",X"C0",X"D3",X"C4",X"75",X"C9",X"1A",X"CE",
		X"B9",X"D2",X"43",X"D7",X"B5",X"DB",X"0C",X"E0",X"46",X"E4",X"5F",X"E8",X"5E",X"EC",X"38",X"F0",
		X"F7",X"F3",X"94",X"F7",X"16",X"FB",X"79",X"FE",X"C0",X"01",X"EA",X"04",X"FC",X"07",X"F0",X"0A",
		X"CF",X"0D",X"91",X"10",X"41",X"13",X"AF",X"15",X"AC",X"16",X"47",X"16",X"24",X"15",X"84",X"13",
		X"5A",X"11",X"FB",X"0E",X"7D",X"0C",X"EE",X"09",X"5D",X"07",X"D1",X"04",X"50",X"02",X"DC",X"FF",
		X"78",X"FD",X"22",X"FB",X"E1",X"F8",X"AD",X"F6",X"8E",X"F4",X"7F",X"F2",X"82",X"F0",X"97",X"EE",
		X"BB",X"EC",X"EF",X"EA",X"36",X"E9",X"86",X"E7",X"EB",X"E5",X"5B",X"E4",X"DC",X"E2",X"69",X"E1",
		X"03",X"E0",X"AB",X"DE",X"5F",X"DD",X"1E",X"DC",X"EB",X"DA",X"C0",X"D9",X"A4",X"D8",X"8F",X"D7",
		X"87",X"D6",X"87",X"D5",X"93",X"D4",X"A7",X"D3",X"C4",X"D2",X"EA",X"D1",X"18",X"D1",X"50",X"D0",
		X"90",X"CF",X"D6",X"CE",X"26",X"CE",X"7B",X"CD",X"D8",X"CC",X"3D",X"CC",X"A7",X"CB",X"19",X"CB",
		X"90",X"CA",X"0F",X"CA",X"A2",X"C9",X"7E",X"CA",X"BD",X"CC",X"CA",X"CF",X"69",X"D3",X"55",X"D7",
		X"73",X"DB",X"A1",X"DF",X"D3",X"E3",X"FC",X"E7",X"13",X"EC",X"16",X"F0",X"FE",X"F3",X"CB",X"F7",
		X"7C",X"FB",X"12",X"FF",X"88",X"02",X"E4",X"05",X"24",X"09",X"4A",X"0C",X"53",X"0F",X"45",X"12",
		X"19",X"15",X"D9",X"17",X"7D",X"1A",X"10",X"1D",X"82",X"1F",X"F2",X"21",X"C8",X"23",X"FD",X"23",
		X"12",X"23",X"61",X"21",X"37",X"1F",X"BC",X"1C",X"18",X"1A",X"56",X"17",X"8F",X"14",X"C8",X"11",
		X"0A",X"0F",X"57",X"0C",X"B6",X"09",X"25",X"07",X"A6",X"04",X"39",X"02",X"E1",X"FF",X"9C",X"FD",
		X"68",X"FB",X"47",X"F9",X"38",X"F7",X"3A",X"F5",X"4F",X"F3",X"73",X"F1",X"AA",X"EF",X"EA",X"ED",
		X"42",X"EC",X"A7",X"EA",X"35",X"EA",X"44",X"EB",X"35",X"ED",X"C6",X"EF",X"B2",X"F2",X"DC",X"F5",
		X"1E",X"F9",X"72",X"FC",X"BF",X"FF",X"06",X"03",X"3E",X"06",X"63",X"09",X"71",X"0C",X"6A",X"0F",
		X"4E",X"12",X"18",X"15",X"CE",X"17",X"6B",X"1A",X"F3",X"1C",X"63",X"1F",X"C1",X"21",X"06",X"24",
		X"3C",X"26",X"58",X"28",X"67",X"2A",X"5B",X"2C",X"4A",X"2E",X"2E",X"2F",X"7E",X"2E",X"E4",X"2C",
		X"9D",X"2A",X"F2",X"27",X"04",X"25",X"F7",X"21",X"D9",X"1E",X"BB",X"1B",X"A1",X"18",X"95",X"15",
		X"97",X"12",X"AD",X"0F",X"D7",X"0C",X"15",X"0A",X"69",X"07",X"D2",X"04",X"50",X"02",X"E4",X"FF",
		X"8B",X"FD",X"47",X"FB",X"15",X"F9",X"F6",X"F6",X"E9",X"F4",X"EE",X"F2",X"07",X"F1",X"28",X"EF",
		X"95",X"ED",X"88",X"ED",X"BF",X"EE",X"C3",X"F0",X"4C",X"F3",X"2B",X"F6",X"36",X"F9",X"59",X"FC",
		X"87",X"FF",X"AE",X"02",X"CC",X"05",X"DD",X"08",X"DB",X"0B",X"C3",X"0E",X"96",X"11",X"53",X"14",
		X"FA",X"16",X"8B",X"19",X"06",X"1C",X"6D",X"1E",X"BC",X"20",X"FA",X"22",X"21",X"25",X"3B",X"27",
		X"38",X"29",X"2E",X"2B",X"05",X"2D",X"E1",X"2E",X"DD",X"2F",X"3C",X"2F",X"A1",X"2D",X"50",X"2B",
		X"98",X"28",X"9C",X"25",X"7B",X"22",X"48",X"1F",X"13",X"1C",X"E3",X"18",X"C2",X"15",X"AF",X"12",
		X"B2",X"0F",X"C6",X"0C",X"F4",X"09",X"33",X"07",X"8B",X"04",X"F8",X"01",X"78",X"FF",X"0F",X"FD",
		X"B9",X"FA",X"78",X"F8",X"4B",X"F6",X"2F",X"F4",X"26",X"F2",X"2E",X"F0",X"45",X"EE",X"90",X"EC",
		X"40",X"EC",X"4F",X"ED",X"32",X"EF",X"A5",X"F1",X"71",X"F4",X"72",X"F7",X"89",X"FA",X"AE",X"FD",
		X"CF",X"00",X"EA",X"03",X"F1",X"06",X"EB",X"09",X"CF",X"0C",X"9E",X"0F",X"59",X"12",X"FE",X"14",
		X"8A",X"17",X"03",X"1A",X"66",X"1C",X"B6",X"1E",X"EF",X"20",X"17",X"23",X"29",X"25",X"2B",X"27",
		X"18",X"29",X"F8",X"2A",X"C2",X"2C",X"7E",X"2E",X"29",X"30",X"C6",X"31",X"52",X"33",X"D2",X"34",
		X"40",X"36",X"A4",X"37",X"F6",X"38",X"3F",X"3A",X"78",X"3B",X"A9",X"3C",X"CD",X"3D",X"E3",X"3E",
		X"F2",X"3F",X"F3",X"40",X"EA",X"41",X"DA",X"42",X"BD",X"43",X"96",X"44",X"68",X"45",X"2F",X"46",
		X"EF",X"46",X"A7",X"47",X"55",X"48",X"FB",X"48",X"9B",X"49",X"34",X"4A",X"C4",X"4A",X"4E",X"4B",
		X"D2",X"4B",X"50",X"4C",X"C6",X"4C",X"36",X"4D",X"A0",X"4D",X"05",X"4E",X"64",X"4E",X"BF",X"4E",
		X"12",X"4F",X"63",X"4F",X"AE",X"4F",X"F4",X"4F",X"34",X"50",X"72",X"50",X"AB",X"50",X"DF",X"50",
		X"0F",X"51",X"3C",X"51",X"64",X"51",X"8A",X"51",X"AB",X"51",X"CB",X"51",X"E5",X"51",X"FC",X"51",
		X"12",X"52",X"23",X"52",X"32",X"52",X"3E",X"52",X"46",X"52",X"4E",X"52",X"50",X"52",X"52",X"52",
		X"51",X"52",X"4E",X"52",X"49",X"52",X"41",X"52",X"38",X"52",X"2B",X"52",X"1E",X"52",X"0E",X"52",
		X"FD",X"51",X"EA",X"51",X"D5",X"51",X"BF",X"51",X"A7",X"51",X"8D",X"51",X"72",X"51",X"56",X"51",
		X"38",X"51",X"1A",X"51",X"F9",X"50",X"D7",X"50",X"B3",X"50",X"91",X"50",X"6B",X"50",X"44",X"50",
		X"1E",X"50",X"F6",X"4F",X"CF",X"4F",X"A4",X"4F",X"7A",X"4F",X"4E",X"4F",X"21",X"4F",X"F3",X"4E",
		X"C5",X"4E",X"95",X"4E",X"66",X"4E",X"35",X"4E",X"07",X"4E",X"D5",X"4D",X"A1",X"4D",X"70",X"4D",
		X"3D",X"4D",X"08",X"4D",X"D5",X"4C",X"A0",X"4C",X"6D",X"4C",X"35",X"4C",X"01",X"4C",X"C7",X"4B",
		X"99",X"4B",X"1C",X"4B",X"1F",X"49",X"FA",X"45",X"1A",X"42",X"C7",X"3D",X"30",X"39",X"79",X"34",
		X"B7",X"2F",X"FB",X"2A",X"4F",X"26",X"BA",X"21",X"40",X"1D",X"E3",X"18",X"A5",X"14",X"87",X"10",
		X"88",X"0C",X"AC",X"08",X"ED",X"04",X"4D",X"01",X"CD",X"FD",X"6A",X"FA",X"23",X"F7",X"F8",X"F3",
		X"EA",X"F0",X"F3",X"ED",X"18",X"EB",X"56",X"E8",X"AA",X"E5",X"16",X"E3",X"9C",X"E0",X"34",X"DE",
		X"E3",X"DB",X"A7",X"D9",X"7F",X"D7",X"69",X"D5",X"69",X"D3",X"77",X"D1",X"9C",X"CF",X"CD",X"CD",
		X"12",X"CC",X"67",X"CA",X"CB",X"C8",X"3F",X"C7",X"C1",X"C5",X"50",X"C4",X"F0",X"C2",X"9B",X"C1",
		X"54",X"C0",X"19",X"BF",X"EB",X"BD",X"C9",X"BC",X"B1",X"BB",X"A5",X"BA",X"A5",X"B9",X"AD",X"B8",
		X"C3",X"B7",X"DF",X"B6",X"07",X"B6",X"37",X"B5",X"72",X"B4",X"B2",X"B3",X"FF",X"B2",X"4F",X"B2",
		X"AB",X"B1",X"0A",X"B1",X"78",X"B0",X"E5",X"AF",X"60",X"AF",X"DC",X"AE",X"64",X"AE",X"EB",X"AD",
		X"82",X"AD",X"14",X"AD",X"B8",X"AC",X"56",X"AC",X"04",X"AC",X"AB",X"AB",X"64",X"AB",X"13",X"AB",
		X"DA",X"AA",X"8F",X"AA",X"63",X"AA",X"17",X"AA",X"98",X"AA",X"96",X"AC",X"AC",X"AF",X"23",X"B3",
		X"99",X"B6",X"04",X"BB",X"6B",X"BF",X"EE",X"C3",X"5D",X"C8",X"C6",X"CC",X"14",X"D1",X"4C",X"D5",
		X"64",X"D9",X"62",X"DD",X"40",X"E1",X"04",X"E5",X"A5",X"E8",X"2C",X"EC",X"94",X"EF",X"E1",X"F2",
		X"13",X"F6",X"2C",X"F9",X"27",X"FC",X"0D",X"FF",X"D5",X"01",X"89",X"04",X"25",X"07",X"98",X"09",
		X"A6",X"0A",X"46",X"0A",X"06",X"09",X"26",X"07",X"EC",X"04",X"70",X"02",X"DA",X"FF",X"30",X"FD",
		X"87",X"FA",X"DF",X"F7",X"43",X"F5",X"B5",X"F2",X"37",X"F0",X"CA",X"ED",X"73",X"EB",X"2A",X"E9",
		X"F5",X"E6",X"D5",X"E4",X"C5",X"E2",X"C8",X"E0",X"DB",X"DE",X"01",X"DD",X"35",X"DB",X"7E",X"D9",
		X"D0",X"D7",X"3C",X"D6",X"A2",X"D4",X"A1",X"D3",X"44",X"D4",X"FE",X"D5",X"76",X"D8",X"62",X"DB",
		X"99",X"DE",X"F5",X"E1",X"67",X"E5",X"D7",X"E8",X"46",X"EC",X"A3",X"EF",X"F0",X"F2",X"27",X"F6",
		X"4A",X"F9",X"53",X"FC",X"46",X"FF",X"20",X"02",X"E6",X"04",X"92",X"07",X"2B",X"0A",X"AA",X"0C",
		X"16",X"0F",X"69",X"11",X"AF",X"13",X"DA",X"15",X"F9",X"17",X"FD",X"19",X"F2",X"1B",X"AC",X"1C",
		X"E3",X"1B",X"37",X"1A",X"E5",X"17",X"37",X"15",X"48",X"12",X"3E",X"0F",X"23",X"0C",X"08",X"09",
		X"F4",X"05",X"EF",X"02",X"FC",X"FF",X"1A",X"FD",X"4B",X"FA",X"92",X"F7",X"EF",X"F4",X"62",X"F2",
		X"E7",X"EF",X"85",X"ED",X"36",X"EB",X"F9",X"E8",X"D4",X"E6",X"BC",X"E4",X"BC",X"E2",X"C9",X"E0",
		X"EE",X"DE",X"15",X"DD",X"AE",X"DB",X"E2",X"DB",X"46",X"DD",X"72",X"DF",X"1B",X"E2",X"15",X"E5",
		X"3B",X"E8",X"76",X"EB",X"B8",X"EE",X"F5",X"F1",X"27",X"F5",X"4B",X"F8",X"59",X"FB",X"52",X"FE",
		X"36",X"01",X"05",X"04",X"BE",X"06",X"5F",X"09",X"EB",X"0B",X"61",X"0E",X"C3",X"10",X"10",X"13",
		X"48",X"15",X"6D",X"17",X"7F",X"19",X"80",X"1B",X"70",X"1D",X"4B",X"1F",X"18",X"21",X"D3",X"22",
		X"80",X"24",X"1C",X"26",X"AB",X"27",X"2A",X"29",X"9B",X"2A",X"FE",X"2B",X"56",X"2D",X"A1",X"2E",
		X"DF",X"2F",X"10",X"31",X"35",X"32",X"50",X"33",X"61",X"34",X"67",X"35",X"62",X"36",X"54",X"37",
		X"3C",X"38",X"1A",X"39",X"F0",X"39",X"BB",X"3A",X"81",X"3B",X"3C",X"3C",X"F0",X"3C",X"9C",X"3D",
		X"40",X"3E",X"DD",X"3E",X"74",X"3F",X"03",X"40",X"8C",X"40",X"0E",X"41",X"8C",X"41",X"01",X"42",
		X"72",X"42",X"DC",X"42",X"41",X"43",X"A2",X"43",X"FC",X"43",X"51",X"44",X"A3",X"44",X"F0",X"44",
		X"38",X"45",X"7B",X"45",X"BA",X"45",X"F6",X"45",X"2B",X"46",X"5F",X"46",X"8F",X"46",X"BB",X"46",
		X"E3",X"46",X"0A",X"47",X"2B",X"47",X"49",X"47",X"65",X"47",X"7E",X"47",X"92",X"47",X"A6",X"47",
		X"B5",X"47",X"C3",X"47",X"CF",X"47",X"D7",X"47",X"DE",X"47",X"E3",X"47",X"E3",X"47",X"E3",X"47",
		X"E1",X"47",X"DD",X"47",X"D6",X"47",X"D0",X"47",X"C6",X"47",X"B9",X"47",X"AC",X"47",X"9D",X"47",
		X"8D",X"47",X"7A",X"47",X"67",X"47",X"50",X"47",X"3B",X"47",X"24",X"47",X"0A",X"47",X"F1",X"46",
		X"D6",X"46",X"B9",X"46",X"9B",X"46",X"7D",X"46",X"5D",X"46",X"3C",X"46",X"1B",X"46",X"F8",X"45",
		X"D3",X"45",X"B0",X"45",X"8C",X"45",X"65",X"45",X"3F",X"45",X"18",X"45",X"EF",X"44",X"C7",X"44",
		X"9D",X"44",X"74",X"44",X"48",X"44",X"1D",X"44",X"F1",X"43",X"C5",X"43",X"99",X"43",X"6C",X"43",
		X"3D",X"43",X"0F",X"43",X"E1",X"42",X"B2",X"42",X"83",X"42",X"54",X"42",X"22",X"42",X"F2",X"41",
		X"C0",X"41",X"8F",X"41",X"5E",X"41",X"2C",X"41",X"FA",X"40",X"C8",X"40",X"95",X"40",X"63",X"40",
		X"2F",X"40",X"FE",X"3F",X"CA",X"3F",X"96",X"3F",X"63",X"3F",X"2F",X"3F",X"FB",X"3E",X"C7",X"3E",
		X"93",X"3E",X"60",X"3E",X"2A",X"3E",X"F5",X"3D",X"C1",X"3D",X"8C",X"3D",X"58",X"3D",X"21",X"3D",
		X"ED",X"3C",X"B9",X"3C",X"83",X"3C",X"4E",X"3C",X"19",X"3C",X"E5",X"3B",X"B0",X"3B",X"79",X"3B",
		X"44",X"3B",X"0E",X"3B",X"DA",X"3A",X"A5",X"3A",X"70",X"3A",X"3B",X"3A",X"05",X"3A",X"D1",X"39",
		X"9C",X"39",X"68",X"39",X"31",X"39",X"FC",X"38",X"C9",X"38",X"92",X"38",X"5E",X"38",X"29",X"38",
		X"F6",X"37",X"C0",X"37",X"8B",X"37",X"58",X"37",X"23",X"37",X"EF",X"36",X"BB",X"36",X"86",X"36",
		X"52",X"36",X"1F",X"36",X"EA",X"35",X"B6",X"35",X"82",X"35",X"4F",X"35",X"1B",X"35",X"E9",X"34",
		X"B4",X"34",X"81",X"34",X"4F",X"34",X"1B",X"34",X"E8",X"33",X"B5",X"33",X"82",X"33",X"50",X"33",
		X"1C",X"33",X"EB",X"32",X"B9",X"32",X"86",X"32",X"53",X"32",X"22",X"32",X"F0",X"31",X"BE",X"31",
		X"8D",X"31",X"5C",X"31",X"2A",X"31",X"F9",X"30",X"C8",X"30",X"97",X"30",X"66",X"30",X"35",X"30",
		X"05",X"30",X"D3",X"2F",X"A3",X"2F",X"74",X"2F",X"43",X"2F",X"13",X"2F",X"E4",X"2E",X"B3",X"2E",
		X"84",X"2E",X"54",X"2E",X"25",X"2E",X"F7",X"2D",X"C8",X"2D",X"98",X"2D",X"6B",X"2D",X"3B",X"2D",
		X"0D",X"2D",X"DD",X"2C",X"B1",X"2C",X"81",X"2C",X"54",X"2C",X"26",X"2C",X"F9",X"2B",X"C9",X"2B",
		X"9C",X"2B",X"70",X"2B",X"42",X"2B",X"15",X"2B",X"E9",X"2A",X"BB",X"2A",X"8F",X"2A",X"62",X"2A",
		X"36",X"2A",X"0B",X"2A",X"DE",X"29",X"B0",X"29",X"85",X"29",X"5A",X"29",X"2E",X"29",X"03",X"29",
		X"D9",X"28",X"AC",X"28",X"82",X"28",X"55",X"28",X"30",X"28",X"D8",X"27",X"0D",X"26",X"03",X"23",
		X"3A",X"1F",X"F1",X"1A",X"66",X"16",X"B3",X"11",X"F6",X"0C",X"3D",X"08",X"94",X"03",X"01",X"FF",
		X"89",X"FA",X"30",X"F6",X"F6",X"F1",X"DB",X"ED",X"E3",X"E9",X"0A",X"E6",X"53",X"E2",X"BB",X"DE",
		X"40",X"DB",X"E5",X"D7",X"A7",X"D4",X"86",X"D1",X"7F",X"CE",X"94",X"CB",X"C3",X"C8",X"0C",X"C6",
		X"6E",X"C3",X"E7",X"C0",X"76",X"BE",X"1D",X"BC",X"D8",X"B9",X"AC",X"B7",X"90",X"B5",X"8C",X"B3",
		X"98",X"B1",X"BB",X"AF",X"EA",X"AD",X"30",X"AC",X"82",X"AA",X"EC",X"A8",X"5D",X"A7",X"E4",X"A5",
		X"75",X"A4",X"1A",X"A3",X"C7",X"A1",X"89",X"A0",X"50",X"9F",X"2D",X"9E",X"0D",X"9D",X"03",X"9C",
		X"F9",X"9A",X"07",X"9A",X"13",X"99",X"39",X"98",X"57",X"97",X"94",X"96",X"C1",X"95",X"20",X"95",
		X"1F",X"94",X"8F",X"92",X"03",X"92",X"5C",X"91",X"D5",X"90",X"43",X"90",X"C6",X"8F",X"47",X"8F",
		X"D7",X"8E",X"68",X"8E",X"05",X"8E",X"A1",X"8D",X"4A",X"8D",X"F4",X"8C",X"AA",X"8C",X"60",X"8C",
		X"21",X"8C",X"E0",X"8B",X"AC",X"8B",X"75",X"8B",X"4B",X"8B",X"1E",X"8B",X"00",X"8B",X"D2",X"8A",
		X"3E",X"8B",X"46",X"8D",X"59",X"90",X"23",X"94",X"58",X"98",X"CF",X"9C",X"62",X"A1",X"01",X"A6",
		X"99",X"AA",X"24",X"AF",X"95",X"B3",X"F2",X"B7",X"30",X"BC",X"52",X"C0",X"54",X"C4",X"3C",X"C8",
		X"00",X"CC",X"AB",X"CF",X"35",X"D3",X"A5",X"D6",X"F7",X"D9",X"32",X"DD",X"4D",X"E0",X"54",X"E3",
		X"3C",X"E6",X"12",X"E9",X"CA",X"EB",X"6A",X"EE",X"C1",X"EF",X"91",X"EF",X"7A",X"EE",X"B7",X"EC",
		X"95",X"EA",X"30",X"E8",X"AA",X"E5",X"10",X"E3",X"75",X"E0",X"DB",X"DD",X"4F",X"DB",X"CE",X"D8",
		X"5D",X"D6",X"FD",X"D3",X"B3",X"D1",X"78",X"CF",X"53",X"CD",X"3F",X"CB",X"3C",X"C9",X"4E",X"C7",
		X"6F",X"C5",X"A5",X"C3",X"E8",X"C1",X"3E",X"C0",X"A2",X"BE",X"17",X"BD",X"9B",X"BB",X"2B",X"BA",
		X"CC",X"B8",X"79",X"B7",X"34",X"B6",X"FB",X"B4",X"CF",X"B3",X"AF",X"B2",X"9A",X"B1",X"92",X"B0",
		X"94",X"AF",X"A2",X"AE",X"B8",X"AD",X"DA",X"AC",X"05",X"AC",X"39",X"AB",X"76",X"AA",X"BD",X"A9",
		X"0B",X"A9",X"63",X"A8",X"C1",X"A7",X"29",X"A7",X"96",X"A6",X"0C",X"A6",X"86",X"A5",X"0F",X"A5",
		X"95",X"A4",X"2D",X"A4",X"BB",X"A3",X"5A",X"A4",X"84",X"A6",X"91",X"A9",X"44",X"AD",X"4C",X"B1",
		X"8F",X"B5",X"EB",X"B9",X"4A",X"BE",X"A4",X"C2",X"ED",X"C6",X"23",X"CB",X"3C",X"CF",X"3C",X"D3",
		X"20",X"D7",X"E6",X"DA",X"8F",X"DE",X"1A",X"E2",X"8A",X"E5",X"DF",X"E8",X"16",X"EC",X"34",X"EF",
		X"38",X"F2",X"24",X"F5",X"F5",X"F7",X"B1",X"FA",X"51",X"FD",X"E5",X"FF",X"1D",X"02",X"C3",X"02",
		X"1B",X"02",X"A2",X"00",X"9B",X"FE",X"3C",X"FC",X"A8",X"F9",X"F7",X"F6",X"3E",X"F4",X"80",X"F1",
		X"CC",X"EE",X"22",X"EC",X"88",X"E9",X"FF",X"E6",X"8A",X"E4",X"28",X"E2",X"D6",X"DF",X"99",X"DD",
		X"72",X"DB",X"5B",X"D9",X"58",X"D7",X"66",X"D5",X"87",X"D3",X"B3",X"D1",X"F9",X"CF",X"46",X"CE",
		X"AF",X"CC",X"12",X"CB",X"61",X"CA",X"4D",X"CB",X"35",X"CD",X"D4",X"CF",X"D7",X"D2",X"22",X"D6",
		X"89",X"D9",X"06",X"DD",X"7E",X"E0",X"F3",X"E3",X"55",X"E7",X"A7",X"EA",X"E4",X"ED",X"09",X"F1",
		X"18",X"F4",X"0F",X"F7",X"F0",X"F9",X"B9",X"FC",X"6A",X"FF",X"02",X"02",X"88",X"04",X"F6",X"06",
		X"53",X"09",X"96",X"0B",X"CF",X"0D",X"E8",X"0F",X"01",X"12",X"57",X"13",X"02",X"13",X"A3",X"11",
		X"84",X"0F",X"F4",X"0C",X"1A",X"0A",X"1B",X"07",X"06",X"04",X"ED",X"00",X"DA",X"FD",X"D3",X"FA",
		X"DA",X"F7",X"F5",X"F4",X"23",X"F2",X"66",X"EF",X"BE",X"EC",X"2D",X"EA",X"AF",X"E7",X"49",X"E5",
		X"F6",X"E2",X"B8",X"E0",X"8E",X"DE",X"76",X"DC",X"73",X"DA",X"80",X"D8",X"A0",X"D6",X"D0",X"D4",
		X"11",X"D3",X"62",X"D1",X"C4",X"CF",X"32",X"CE",X"B1",X"CC",X"3F",X"CB",X"DB",X"C9",X"82",X"C8",
		X"38",X"C7",X"F9",X"C5",X"C8",X"C4",X"A0",X"C3",X"87",X"C2",X"77",X"C1",X"75",X"C0",X"79",X"BF",
		X"8B",X"BE",X"A2",X"BD",X"C8",X"BC",X"F3",X"BB",X"2B",X"BB",X"65",X"BA",X"AE",X"B9",X"FA",X"B8",
		X"56",X"B8",X"B1",X"B7",X"1D",X"B7",X"7B",X"B6",X"69",X"B6",X"F2",X"B7",X"96",X"BA",X"F2",X"BD",
		X"BD",X"C1",X"CF",X"C5",X"01",X"CA",X"3F",X"CE",X"7A",X"D2",X"AA",X"D6",X"C7",X"DA",X"CD",X"DE",
		X"B6",X"E2",X"87",X"E6",X"3A",X"EA",X"D1",X"ED",X"4B",X"F1",X"A8",X"F4",X"EA",X"F7",X"13",X"FB",
		X"1F",X"FE",X"12",X"01",X"EB",X"03",X"AF",X"06",X"56",X"09",X"EF",X"0B",X"66",X"0E",X"CF",X"10",
		X"FA",X"11",X"9B",X"11",X"50",X"10",X"59",X"0E",X"03",X"0C",X"67",X"09",X"AD",X"06",X"DE",X"03",
		X"0E",X"01",X"42",X"FE",X"81",X"FB",X"CE",X"F8",X"2E",X"F6",X"9D",X"F3",X"21",X"F1",X"B9",X"EE",
		X"64",X"EC",X"22",X"EA",X"F2",X"E7",X"D8",X"E5",X"CE",X"E3",X"D9",X"E1",X"F1",X"DF",X"20",X"DE",
		X"58",X"DC",X"A8",X"DA",X"FA",X"D8",X"B8",X"D7",X"11",X"D8",X"9F",X"D9",X"F6",X"DB",X"CE",X"DE",
		X"F3",X"E1",X"45",X"E5",X"AD",X"E8",X"1A",X"EC",X"84",X"EF",X"DF",X"F2",X"2A",X"F6",X"60",X"F9",
		X"82",X"FC",X"8A",X"FF",X"7D",X"02",X"57",X"05",X"1C",X"08",X"C7",X"0A",X"5F",X"0D",X"DF",X"0F",
		X"4B",X"12",X"9D",X"14",X"E0",X"16",X"0A",X"19",X"29",X"1B",X"2A",X"1D",X"29",X"1F",X"1C",X"20",
		X"75",X"1F",X"DB",X"1D",X"8E",X"1B",X"DE",X"18",X"E6",X"15",X"D1",X"12",X"A7",X"0F",X"7F",X"0C",
		X"5A",X"09",X"45",X"06",X"3F",X"03",X"4E",X"00",X"6F",X"FD",X"A7",X"FA",X"F5",X"F7",X"59",X"F5",
		X"CF",X"F2",X"5E",X"F0",X"FF",X"ED",X"B7",X"EB",X"84",X"E9",X"61",X"E7",X"51",X"E5",X"57",X"E3",
		X"6A",X"E1",X"91",X"DF",X"C7",X"DD",X"0E",X"DC",X"67",X"DA",X"CA",X"D8",X"40",X"D7",X"C4",X"D5",
		X"55",X"D4",X"F3",X"D2",X"A0",X"D1",X"57",X"D0",X"1B",X"CF",X"EC",X"CD",X"CA",X"CC",X"B0",X"CB",
		X"A3",X"CA",X"9F",X"C9",X"A7",X"C8",X"B6",X"C7",X"D1",X"C6",X"F4",X"C5",X"23",X"C5",X"56",X"C4",
		X"96",X"C3",X"D9",X"C2",X"2A",X"C2",X"7A",X"C1",X"E0",X"C0",X"35",X"C0",X"5F",X"C0",X"25",X"C2",
		X"E3",X"C4",X"51",X"C8",X"21",X"CC",X"32",X"D0",X"5E",X"D4",X"94",X"D8",X"C3",X"DC",X"E9",X"E0",
		X"F6",X"E4",X"EF",X"E8",X"CC",X"EC",X"8D",X"F0",X"32",X"F4",X"BA",X"F7",X"26",X"FB",X"76",X"FE",
		X"AA",X"01",X"C4",X"04",X"C5",X"07",X"A9",X"0A",X"78",X"0D",X"2D",X"10",X"CA",X"12",X"51",X"15",
		X"C3",X"17",X"1C",X"1A",X"64",X"1C",X"95",X"1E",X"B4",X"20",X"BF",X"22",X"BA",X"24",X"A0",X"26",
		X"77",X"28",X"3D",X"2A",X"F0",X"2B",X"96",X"2D",X"2C",X"2F",X"B3",X"30",X"2C",X"32",X"97",X"33",
		X"F4",X"34",X"44",X"36",X"88",X"37",X"BE",X"38",X"E8",X"39",X"0A",X"3B",X"1D",X"3C",X"26",X"3D",
		X"26",X"3E",X"1A",X"3F",X"05",X"40",X"E4",X"40",X"C6",X"41",X"09",X"42",X"A4",X"40",X"3B",X"3E",
		X"04",X"3B",X"98",X"37",X"2B",X"34",X"1A",X"30",X"0D",X"2C",X"F8",X"27",X"F6",X"23",X"01",X"20",
		X"24",X"1C",X"5F",X"18",X"B5",X"14",X"26",X"11",X"B4",X"0D",X"5C",X"0A",X"1F",X"07",X"FF",X"03",
		X"F6",X"00",X"09",X"FE",X"33",X"FB",X"77",X"F8",X"D0",X"F5",X"42",X"F3",X"C7",X"F0",X"66",X"EE",
		X"1F",X"EC",X"27",X"EB",X"B7",X"EB",X"2F",X"ED",X"4A",X"EF",X"C8",X"F1",X"85",X"F4",X"61",X"F7",
		X"4D",X"FA",X"3C",X"FD",X"23",X"00",X"FE",X"02",X"CE",X"05",X"89",X"08",X"31",X"0B",X"C6",X"0D",
		X"45",X"10",X"B0",X"12",X"07",X"15",X"4B",X"17",X"79",X"19",X"97",X"1B",X"A1",X"1D",X"99",X"1F",
		X"7F",X"21",X"57",X"23",X"16",X"25",X"D8",X"26",X"15",X"28",X"AD",X"27",X"19",X"26",X"BE",X"23",
		X"E4",X"20",X"BD",X"1D",X"6B",X"1A",X"03",X"17",X"98",X"13",X"2E",X"10",X"D6",X"0C",X"8C",X"09",
		X"57",X"06",X"38",X"03",X"32",X"00",X"42",X"FD",X"69",X"FA",X"A7",X"F7",X"FD",X"F4",X"67",X"F2",
		X"E9",X"EF",X"81",X"ED",X"2D",X"EB",X"ED",X"E8",X"BF",X"E6",X"A7",X"E4",X"A1",X"E2",X"AE",X"E0",
		X"CA",X"DE",X"F9",X"DC",X"39",X"DB",X"88",X"D9",X"E7",X"D7",X"57",X"D6",X"D1",X"D4",X"5A",X"D3",
		X"F4",X"D1",X"9B",X"D0",X"4C",X"CF",X"0B",X"CE",X"D5",X"CC",X"AD",X"CB",X"8D",X"CA",X"7B",X"C9",
		X"73",X"C8",X"76",X"C7",X"82",X"C6",X"98",X"C5",X"B9",X"C4",X"E2",X"C3",X"14",X"C3",X"4D",X"C2",
		X"8F",X"C1",X"DB",X"C0",X"2E",X"C0",X"88",X"BF",X"EA",X"BE",X"52",X"BE",X"C1",X"BD",X"38",X"BD",
		X"B5",X"BC",X"39",X"BC",X"C1",X"BB",X"50",X"BB",X"E5",X"BA",X"7F",X"BA",X"1F",X"BA",X"C4",X"B9",
		X"6F",X"B9",X"1D",X"B9",X"D0",X"B8",X"89",X"B8",X"45",X"B8",X"07",X"B8",X"CB",X"B7",X"95",X"B7",
		X"60",X"B7",X"33",X"B7",X"07",X"B7",X"DF",X"B6",X"BA",X"B6",X"98",X"B6",X"7B",X"B6",X"60",X"B6",
		X"49",X"B6",X"34",X"B6",X"21",X"B6",X"11",X"B6",X"05",X"B6",X"FB",X"B5",X"F3",X"B5",X"ED",X"B5",
		X"E8",X"B5",X"E8",X"B5",X"E9",X"B5",X"ED",X"B5",X"F2",X"B5",X"F9",X"B5",X"03",X"B6",X"0F",X"B6",
		X"1B",X"B6",X"28",X"B6",X"39",X"B6",X"4C",X"B6",X"5E",X"B6",X"73",X"B6",X"89",X"B6",X"A0",X"B6",
		X"B9",X"B6",X"D4",X"B6",X"EF",X"B6",X"0D",X"B7",X"2A",X"B7",X"4A",X"B7",X"69",X"B7",X"89",X"B7",
		X"AC",X"B7",X"CE",X"B7",X"F4",X"B7",X"19",X"B8",X"3E",X"B8",X"65",X"B8",X"8C",X"B8",X"B4",X"B8",
		X"DB",X"B8",X"05",X"B9",X"31",X"B9",X"5B",X"B9",X"86",X"B9",X"B4",X"B9",X"DF",X"B9",X"0D",X"BA",
		X"3A",X"BA",X"68",X"BA",X"98",X"BA",X"C6",X"BA",X"F6",X"BA",X"26",X"BB",X"57",X"BB",X"86",X"BB",
		X"B8",X"BB",X"EA",X"BB",X"1C",X"BC",X"4E",X"BC",X"82",X"BC",X"B5",X"BC",X"E8",X"BC",X"1B",X"BD",
		X"4E",X"BD",X"84",X"BD",X"B7",X"BD",X"EB",X"BD",X"20",X"BE",X"55",X"BE",X"88",X"BE",X"BF",X"BE",
		X"F3",X"BE",X"2B",X"BF",X"5F",X"BF",X"97",X"BF",X"CA",X"BF",X"05",X"C0",X"35",X"C0",X"71",X"C0",
		X"99",X"C0",X"54",X"C1",X"A7",X"C3",X"09",X"C7",X"21",X"CB",X"A4",X"CF",X"64",X"D4",X"3E",X"D9",
		X"21",X"DE",X"FA",X"E2",X"C1",X"E7",X"70",X"EC",X"04",X"F1",X"76",X"F5",X"C8",X"F9",X"FB",X"FD",
		X"0A",X"02",X"F9",X"05",X"C8",X"09",X"79",X"0D",X"07",X"11",X"7A",X"14",X"CE",X"17",X"06",X"1B",
		X"20",X"1E",X"20",X"21",X"05",X"24",X"D2",X"26",X"85",X"29",X"21",X"2C",X"A3",X"2E",X"11",X"31",
		X"67",X"33",X"A9",X"35",X"D5",X"37",X"F0",X"39",X"F4",X"3B",X"E8",X"3D",X"C8",X"3F",X"98",X"41",
		X"53",X"43",X"01",X"45",X"9D",X"46",X"2A",X"48",X"A9",X"49",X"1A",X"4B",X"78",X"4C",X"CD",X"4D",
		X"11",X"4F",X"4D",X"50",X"77",X"51",X"98",X"52",X"AA",X"53",X"B6",X"54",X"AE",X"55",X"AD",X"56",
		X"39",X"57",X"2A",X"56",X"EC",X"53",X"E8",X"50",X"68",X"4D",X"9E",X"49",X"AB",X"45",X"A8",X"41",
		X"A2",X"3D",X"A6",X"39",X"BB",X"35",X"E4",X"31",X"25",X"2E",X"80",X"2A",X"F5",X"26",X"84",X"23",
		X"2E",X"20",X"F1",X"1C",X"D1",X"19",X"C8",X"16",X"DA",X"13",X"02",X"11",X"45",X"0E",X"99",X"0B",
		X"0C",X"09",X"8A",X"06",X"2B",X"04",X"D1",X"01",X"8D",X"00",X"E9",X"00",X"39",X"02",X"40",X"04",
		X"A9",X"06",X"5C",X"09",X"31",X"0C",X"19",X"0F",X"02",X"12",X"E6",X"14",X"C0",X"17",X"8B",X"1A",
		X"42",X"1D",X"E8",X"1F",X"77",X"22",X"F5",X"24",X"5C",X"27",X"AE",X"29",X"EE",X"2B",X"19",X"2E",
		X"30",X"30",X"34",X"32",X"26",X"34",X"05",X"36",X"D5",X"37",X"90",X"39",X"45",X"3B",X"A9",X"3C",
		X"7E",X"3C",X"06",X"3B",X"BD",X"38",X"E9",X"35",X"C2",X"32",X"68",X"2F",X"FA",X"2B",X"81",X"28",
		X"0D",X"25",X"A4",X"21",X"4D",X"1E",X"08",X"1B",X"DB",X"17",X"C2",X"14",X"C2",X"11",X"D8",X"0E",
		X"07",X"0C",X"4A",X"09",X"A8",X"06",X"17",X"04",X"9E",X"01",X"3C",X"FF",X"EB",X"FC",X"B0",X"FA",
		X"87",X"F8",X"70",X"F6",X"6D",X"F4",X"7B",X"F2",X"99",X"F0",X"C8",X"EE",X"09",X"ED",X"57",X"EB",
		X"B5",X"E9",X"20",X"E8",X"9C",X"E6",X"25",X"E5",X"BA",X"E3",X"5C",X"E2",X"0C",X"E1",X"C8",X"DF",
		X"90",X"DE",X"62",X"DD",X"3F",X"DC",X"28",X"DB",X"1B",X"DA",X"17",X"D9",X"1F",X"D8",X"30",X"D7",
		X"48",X"D6",X"6B",X"D5",X"96",X"D4",X"CB",X"D3",X"06",X"D3",X"4A",X"D2",X"95",X"D1",X"E7",X"D0",
		X"40",X"D0",X"A2",X"CF",X"09",X"CF",X"78",X"CE",X"EB",X"CD",X"66",X"CD",X"E7",X"CC",X"6C",X"CC",
		X"F9",X"CB",X"8A",X"CB",X"20",X"CB",X"BC",X"CA",X"5D",X"CA",X"01",X"CA",X"AB",X"C9",X"59",X"C9",
		X"0C",X"C9",X"C3",X"C8",X"7E",X"C8",X"3D",X"C8",X"00",X"C8",X"C7",X"C7",X"90",X"C7",X"5E",X"C7",
		X"2E",X"C7",X"02",X"C7",X"D9",X"C6",X"B3",X"C6",X"91",X"C6",X"71",X"C6",X"54",X"C6",X"3A",X"C6",
		X"20",X"C6",X"0D",X"C6",X"F8",X"C5",X"E9",X"C5",X"D9",X"C5",X"CE",X"C5",X"C3",X"C5",X"BD",X"C5",
		X"B6",X"C5",X"B3",X"C5",X"AF",X"C5",X"B1",X"C5",X"AF",X"C5",X"B5",X"C5",X"B8",X"C5",X"BF",X"C5",
		X"C8",X"C5",X"D1",X"C5",X"DA",X"C5",X"E8",X"C5",X"F3",X"C5",X"11",X"C6",X"68",X"C7",X"3B",X"CA",
		X"D4",X"CD",X"13",X"D2",X"75",X"D6",X"DB",X"DA",X"AE",X"DF",X"76",X"E4",X"38",X"E9",X"E1",X"ED",
		X"73",X"F2",X"E6",X"F6",X"39",X"FB",X"6B",X"FF",X"7B",X"03",X"6E",X"07",X"3E",X"0B",X"F1",X"0E",
		X"82",X"12",X"F7",X"15",X"4C",X"19",X"87",X"1C",X"A3",X"1F",X"A6",X"22",X"8A",X"25",X"59",X"28",
		X"0E",X"2B",X"AA",X"2D",X"2E",X"30",X"9C",X"32",X"F6",X"34",X"39",X"37",X"66",X"39",X"80",X"3B",
		X"87",X"3D",X"7A",X"3F",X"5B",X"41",X"2B",X"43",X"E8",X"44",X"95",X"46",X"33",X"48",X"C0",X"49",
		X"3F",X"4B",X"AE",X"4C",X"10",X"4E",X"62",X"4F",X"A9",X"50",X"DE",X"51",X"0E",X"53",X"2B",X"54",
		X"41",X"55",X"48",X"56",X"47",X"57",X"35",X"58",X"21",X"59",X"E5",X"58",X"1A",X"57",X"65",X"54",
		X"08",X"51",X"52",X"4D",X"5C",X"49",X"50",X"45",X"39",X"41",X"29",X"3D",X"22",X"39",X"31",X"35",
		X"57",X"31",X"94",X"2D",X"EC",X"29",X"63",X"26",X"F1",X"22",X"9B",X"1F",X"5F",X"1C",X"3F",X"19",
		X"37",X"16",X"48",X"13",X"72",X"10",X"B4",X"0D",X"0D",X"0B",X"78",X"08",X"02",X"06",X"92",X"03",
		X"8A",X"01",X"25",X"01",X"07",X"02",X"BC",X"03",X"FE",X"05",X"93",X"08",X"5D",X"0B",X"42",X"0E",
		X"30",X"11",X"1E",X"14",X"03",X"17",X"D9",X"19",X"A1",X"1C",X"52",X"1F",X"F2",X"21",X"7B",X"24",
		X"F2",X"26",X"53",X"29",X"9F",X"2B",X"D6",X"2D",X"FC",X"2F",X"0C",X"32",X"0C",X"34",X"F7",X"35",
		X"D1",X"37",X"99",X"39",X"53",X"3B",X"FA",X"3C",X"93",X"3E",X"1B",X"40",X"95",X"41",X"00",X"43",
		X"5F",X"44",X"AE",X"45",X"F3",X"46",X"27",X"48",X"52",X"49",X"6F",X"4A",X"84",X"4B",X"8A",X"4C",
		X"87",X"4D",X"78",X"4E",X"60",X"4F",X"3E",X"50",X"12",X"51",X"DC",X"51",X"A0",X"52",X"58",X"53",
		X"08",X"54",X"B0",X"54",X"52",X"55",X"E9",X"55",X"7C",X"56",X"03",X"57",X"8B",X"57",X"DB",X"57",
		X"B0",X"56",X"2C",X"54",X"DE",X"50",X"04",X"4D",X"DF",X"48",X"8A",X"44",X"27",X"40",X"BE",X"3B",
		X"66",X"37",X"1C",X"33",X"EA",X"2E",X"D0",X"2A",X"D7",X"26",X"F6",X"22",X"34",X"1F",X"8F",X"1B",
		X"0B",X"18",X"9E",X"14",X"4F",X"11",X"1C",X"0E",X"04",X"0B",X"06",X"08",X"1F",X"05",X"52",X"02",
		X"9E",X"FF",X"00",X"FD",X"79",X"FA",X"07",X"F8",X"AB",X"F5",X"62",X"F3",X"2D",X"F1",X"0B",X"EF",
		X"FE",X"EC",X"FF",X"EA",X"17",X"E9",X"3C",X"E7",X"74",X"E5",X"BA",X"E3",X"11",X"E2",X"77",X"E0",
		X"EB",X"DE",X"6E",X"DD",X"FE",X"DB",X"9A",X"DA",X"45",X"D9",X"FB",X"D7",X"BE",X"D6",X"8E",X"D5",
		X"66",X"D4",X"4B",X"D3",X"3C",X"D2",X"38",X"D1",X"3C",X"D0",X"48",X"CF",X"75",X"CE",X"01",X"CF",
		X"FE",X"D0",X"D1",X"D3",X"3D",X"D7",X"FC",X"DA",X"F1",X"DE",X"F9",X"E2",X"07",X"E7",X"0C",X"EB",
		X"04",X"EF",X"E5",X"F2",X"B1",X"F6",X"5F",X"FA",X"F5",X"FD",X"6E",X"01",X"CC",X"04",X"10",X"08",
		X"37",X"0B",X"45",X"0E",X"36",X"11",X"11",X"14",X"D0",X"16",X"7B",X"19",X"0B",X"1C",X"89",X"1E",
		X"EC",X"20",X"37",X"23",X"33",X"24",X"A1",X"23",X"26",X"22",X"02",X"20",X"79",X"1D",X"B0",X"1A",
		X"C9",X"17",X"CC",X"14",X"D1",X"11",X"D9",X"0E",X"EF",X"0B",X"11",X"09",X"48",X"06",X"91",X"03",
		X"EF",X"00",X"63",X"FE",X"EA",X"FB",X"85",X"F9",X"32",X"F7",X"F6",X"F4",X"CA",X"F2",X"B3",X"F0",
		X"AC",X"EE",X"BA",X"EC",X"D4",X"EA",X"07",X"E9",X"38",X"E7",X"E9",X"E5",X"41",X"E6",X"CD",X"E7",
		X"23",X"EA",X"F7",X"EC",X"1F",X"F0",X"6F",X"F3",X"D7",X"F6",X"42",X"FA",X"A8",X"FD",X"01",X"01",
		X"4A",X"04",X"7E",X"07",X"9D",X"0A",X"A2",X"0D",X"90",X"10",X"68",X"13",X"29",X"16",X"D1",X"18",
		X"65",X"1B",X"DE",X"1D",X"47",X"20",X"95",X"22",X"D3",X"24",X"F8",X"26",X"11",X"29",X"0E",X"2B",
		X"04",X"2D",X"DA",X"2D",X"12",X"2D",X"57",X"2B",X"E9",X"28",X"19",X"26",X"02",X"23",X"CD",X"1F",
		X"86",X"1C",X"3F",X"19",X"FD",X"15",X"CA",X"12",X"AA",X"0F",X"9C",X"0C",X"A1",X"09",X"BF",X"06",
		X"F3",X"03",X"3B",X"01",X"9D",X"FE",X"12",X"FC",X"9C",X"F9",X"3C",X"F7",X"F0",X"F4",X"B8",X"F2",
		X"94",X"F0",X"81",X"EE",X"83",X"EC",X"8B",X"EA",X"EF",X"E8",X"E9",X"E8",X"31",X"EA",X"4B",X"EC",
		X"F1",X"EE",X"E9",X"F1",X"17",X"F5",X"5B",X"F8",X"A5",X"FB",X"EF",X"FE",X"2C",X"02",X"5A",X"05",
		X"74",X"08",X"79",X"0B",X"6A",X"0E",X"42",X"11",X"03",X"14",X"AD",X"16",X"43",X"19",X"C1",X"1B",
		X"2A",X"1E",X"7D",X"20",X"BC",X"22",X"E7",X"24",X"00",X"27",X"04",X"29",X"F8",X"2A",X"D6",X"2C",
		X"A8",X"2E",X"65",X"30",X"14",X"32",X"B2",X"33",X"42",X"35",X"C2",X"36",X"35",X"38",X"99",X"39",
		X"F0",X"3A",X"39",X"3C",X"77",X"3D",X"A6",X"3E",X"CD",X"3F",X"E6",X"40",X"F4",X"41",X"F7",X"42",
		X"F0",X"43",X"DF",X"44",X"C4",X"45",X"9E",X"46",X"72",X"47",X"39",X"48",X"FB",X"48",X"B0",X"49",
		X"61",X"4A",X"08",X"4B",X"AA",X"4B",X"40",X"4C",X"D4",X"4C",X"5E",X"4D",X"E1",X"4D",X"5D",X"4E",
		X"D4",X"4E",X"42",X"4F",X"B0",X"4F",X"13",X"50",X"72",X"50",X"CA",X"50",X"20",X"51",X"6E",X"51",
		X"BB",X"51",X"FE",X"51",X"40",X"52",X"7C",X"52",X"B6",X"52",X"E6",X"52",X"19",X"53",X"43",X"53",
		X"6D",X"53",X"8F",X"53",X"B4",X"53",X"CC",X"53",X"ED",X"53",X"FA",X"53",X"1D",X"54",X"8B",X"53",
		X"57",X"51",X"1B",X"4E",X"2C",X"4A",X"D5",X"45",X"3F",X"41",X"90",X"3C",X"D5",X"37",X"24",X"33",
		X"81",X"2E",X"F9",X"29",X"87",X"25",X"37",X"21",X"04",X"1D",X"F1",X"18",X"FD",X"14",X"28",X"11",
		X"73",X"0D",X"DD",X"09",X"64",X"06",X"09",X"03",X"C9",X"FF",X"A8",X"FC",X"9D",X"F9",X"AF",X"F6",
		X"D8",X"F3",X"1B",X"F1",X"82",X"EE",X"50",X"ED",X"9E",X"ED",X"D7",X"EE",X"B7",X"F0",X"F7",X"F2",
		X"79",X"F5",X"1E",X"F8",X"D4",X"FA",X"8C",X"FD",X"3F",X"00",X"EA",X"02",X"86",X"05",X"12",X"08",
		X"8C",X"0A",X"F4",X"0C",X"48",X"0F",X"8C",X"11",X"B8",X"13",X"D7",X"15",X"DF",X"17",X"D9",X"19",
		X"BF",X"1B",X"97",X"1D",X"5A",X"1F",X"14",X"21",X"B4",X"22",X"59",X"24",X"69",X"25",X"D4",X"24",
		X"12",X"23",X"8F",X"20",X"89",X"1D",X"4D",X"1A",X"07",X"17",X"6F",X"13",X"DC",X"0F",X"4A",X"0C",
		X"CC",X"08",X"5B",X"05",X"03",X"02",X"C1",X"FE",X"98",X"FB",X"85",X"F8",X"8F",X"F5",X"AD",X"F2",
		X"E5",X"EF",X"34",X"ED",X"9C",X"EA",X"17",X"E8",X"AC",X"E5",X"53",X"E3",X"12",X"E1",X"DF",X"DE",
		X"C8",X"DC",X"BE",X"DA",X"EE",X"D9",X"B8",X"DA",X"71",X"DC",X"D8",X"DE",X"A0",X"E1",X"B2",X"E4",
		X"DD",X"E7",X"1D",X"EB",X"5A",X"EE",X"93",X"F1",X"BA",X"F4",X"D4",X"F7",X"D9",X"FA",X"C9",X"FD",
		X"A2",X"00",X"65",X"03",X"11",X"06",X"A8",X"08",X"29",X"0B",X"97",X"0D",X"EC",X"0F",X"32",X"12",
		X"61",X"14",X"7D",X"16",X"87",X"18",X"80",X"1A",X"65",X"1C",X"3A",X"1E",X"FF",X"1F",X"B5",X"21",
		X"59",X"23",X"F1",X"24",X"76",X"26",X"F0",X"27",X"5B",X"29",X"BA",X"2A",X"0A",X"2C",X"4F",X"2D",
		X"87",X"2E",X"B6",X"2F",X"D6",X"30",X"ED",X"31",X"F8",X"32",X"F8",X"33",X"F1",X"34",X"DD",X"35",
		X"C1",X"36",X"9C",X"37",X"6D",X"38",X"36",X"39",X"F8",X"39",X"B0",X"3A",X"63",X"3B",X"0A",X"3C",
		X"AC",X"3C",X"48",X"3D",X"DC",X"3D",X"69",X"3E",X"F0",X"3E",X"70",X"3F",X"EA",X"3F",X"5E",X"40",
		X"CD",X"40",X"34",X"41",X"9A",X"41",X"F7",X"41",X"51",X"42",X"A4",X"42",X"F4",X"42",X"3F",X"43",
		X"86",X"43",X"C8",X"43",X"07",X"44",X"41",X"44",X"78",X"44",X"AA",X"44",X"D8",X"44",X"05",X"45",
		X"2B",X"45",X"50",X"45",X"71",X"45",X"8F",X"45",X"AA",X"45",X"C3",X"45",X"D7",X"45",X"EB",X"45",
		X"FA",X"45",X"07",X"46",X"12",X"46",X"1D",X"46",X"21",X"46",X"26",X"46",X"26",X"46",X"28",X"46",
		X"23",X"46",X"20",X"46",X"18",X"46",X"13",X"46",X"06",X"46",X"FE",X"45",X"F0",X"45",X"E1",X"45",
		X"CF",X"45",X"BF",X"45",X"AA",X"45",X"98",X"45",X"7E",X"45",X"6D",X"45",X"4C",X"45",X"41",X"45",
		X"6A",X"44",X"EF",X"41",X"78",X"3E",X"4E",X"3A",X"C2",X"35",X"FB",X"30",X"1D",X"2C",X"37",X"27",
		X"5D",X"22",X"92",X"1D",X"E4",X"18",X"51",X"14",X"DD",X"0F",X"88",X"0B",X"58",X"07",X"46",X"03",
		X"59",X"FF",X"88",X"FB",X"D9",X"F7",X"46",X"F4",X"D6",X"F0",X"80",X"ED",X"48",X"EA",X"2B",X"E7",
		X"2C",X"E4",X"43",X"E1",X"76",X"DE",X"C3",X"DB",X"27",X"D9",X"A0",X"D6",X"31",X"D4",X"D9",X"D1",
		X"95",X"CF",X"65",X"CD",X"4B",X"CB",X"44",X"C9",X"50",X"C7",X"6C",X"C5",X"9D",X"C3",X"DD",X"C1",
		X"2D",X"C0",X"8E",X"BE",X"FE",X"BC",X"7E",X"BB",X"0D",X"BA",X"A8",X"B8",X"54",X"B7",X"0B",X"B6",
		X"D0",X"B4",X"A0",X"B3",X"7D",X"B2",X"69",X"B1",X"5C",X"B0",X"5C",X"AF",X"67",X"AE",X"7C",X"AD",
		X"9A",X"AC",X"C3",X"AB",X"F6",X"AA",X"30",X"AA",X"74",X"A9",X"C2",X"A8",X"17",X"A8",X"73",X"A7",
		X"DA",X"A6",X"49",X"A6",X"BB",X"A5",X"37",X"A5",X"BA",X"A4",X"41",X"A4",X"D1",X"A3",X"67",X"A3",
		X"03",X"A3",X"A4",X"A2",X"4A",X"A2",X"F9",X"A1",X"AB",X"A1",X"63",X"A1",X"1F",X"A1",X"E1",X"A0",
		X"A6",X"A0",X"73",X"A0",X"49",X"A0",X"5C",X"A1",X"F3",X"A3",X"66",X"A7",X"77",X"AB",X"DB",X"AF",
		X"75",X"B4",X"1E",X"B9",X"CE",X"BD",X"71",X"C2",X"06",X"C7",X"7D",X"CB",X"DD",X"CF",X"1C",X"D4",
		X"3E",X"D8",X"40",X"DC",X"25",X"E0",X"E8",X"E3",X"8E",X"E7",X"16",X"EB",X"81",X"EE",X"D2",X"F1",
		X"04",X"F5",X"1E",X"F8",X"19",X"FB",X"03",X"FE",X"C8",X"00",X"80",X"03",X"09",X"05",X"EE",X"04",
		X"DC",X"03",X"11",X"02",X"DE",X"FF",X"62",X"FD",X"C2",X"FA",X"0B",X"F8",X"53",X"F5",X"9A",X"F2",
		X"EF",X"EF",X"4D",X"ED",X"C0",X"EA",X"40",X"E8",X"D6",X"E5",X"7E",X"E3",X"3B",X"E1",X"07",X"DF",
		X"EB",X"DC",X"DF",X"DA",X"E5",X"D8",X"FD",X"D6",X"28",X"D5",X"61",X"D3",X"AC",X"D1",X"06",X"D0",
		X"6E",X"CE",X"E7",X"CC",X"6E",X"CB",X"03",X"CA",X"A5",X"C8",X"55",X"C7",X"12",X"C6",X"DA",X"C4",
		X"AF",X"C3",X"91",X"C2",X"7B",X"C1",X"75",X"C0",X"74",X"BF",X"80",X"BE",X"95",X"BD",X"B6",X"BC",
		X"DE",X"BB",X"12",X"BB",X"48",X"BA",X"8F",X"B9",X"D7",X"B8",X"2E",X"B8",X"86",X"B7",X"EE",X"B6",
		X"54",X"B6",X"C8",X"B5",X"3A",X"B5",X"C2",X"B4",X"39",X"B4",X"A3",X"B4",X"AE",X"B6",X"B1",X"B9",
		X"64",X"BD",X"78",X"C1",X"CA",X"C5",X"36",X"CA",X"AB",X"CE",X"18",X"D3",X"78",X"D7",X"BD",X"DB",
		X"EE",X"DF",X"02",X"E4",X"F8",X"E7",X"CF",X"EB",X"89",X"EF",X"27",X"F3",X"A6",X"F6",X"08",X"FA",
		X"4E",X"FD",X"78",X"00",X"87",X"03",X"7D",X"06",X"5A",X"09",X"1D",X"0C",X"C7",X"0E",X"60",X"11",
		X"B6",X"13",X"80",X"14",X"DE",X"13",X"5F",X"12",X"44",X"10",X"CD",X"0D",X"1B",X"0B",X"4A",X"08",
		X"6B",X"05",X"8C",X"02",X"B4",X"FF",X"E7",X"FC",X"2A",X"FA",X"7E",X"F7",X"E5",X"F4",X"5F",X"F2",
		X"EE",X"EF",X"91",X"ED",X"46",X"EB",X"10",X"E9",X"EE",X"E6",X"DA",X"E4",X"DE",X"E2",X"F1",X"E0",
		X"19",X"DF",X"4A",X"DD",X"96",X"DB",X"DD",X"D9",X"ED",X"D8",X"B0",X"D9",X"85",X"DB",X"1C",X"DE",
		X"1F",X"E1",X"72",X"E4",X"E6",X"E7",X"6E",X"EB",X"F5",X"EE",X"76",X"F2",X"E9",X"F5",X"4A",X"F9",
		X"93",X"FC",X"C9",X"FF",X"E4",X"02",X"E8",X"05",X"D2",X"08",X"A6",X"0B",X"62",X"0E",X"07",X"11",
		X"94",X"13",X"0D",X"16",X"6E",X"18",X"BE",X"1A",X"F4",X"1C",X"1D",X"1F",X"2D",X"21",X"1C",X"23",
		X"A2",X"23",X"AB",X"22",X"CE",X"20",X"4E",X"1E",X"73",X"1B",X"59",X"18",X"24",X"15",X"E0",X"11",
		X"A0",X"0E",X"65",X"0B",X"39",X"08",X"20",X"05",X"1C",X"02",X"2C",X"FF",X"53",X"FC",X"8F",X"F9",
		X"E1",X"F6",X"4C",X"F4",X"CA",X"F1",X"60",X"EF",X"08",X"ED",X"C6",X"EA",X"96",X"E8",X"7D",X"E6",
		X"72",X"E4",X"81",X"E2",X"8D",X"E0",X"37",X"DF",X"96",X"DF",X"1A",X"E1",X"6B",X"E3",X"33",X"E6",
		X"4F",X"E9",X"92",X"EC",X"EC",X"EF",X"48",X"F3",X"A3",X"F6",X"EE",X"F9",X"2A",X"FD",X"50",X"00",
		X"63",X"03",X"5C",X"06",X"43",X"09",X"0D",X"0C",X"C4",X"0E",X"63",X"11",X"ED",X"13",X"5E",X"16",
		X"BE",X"18",X"06",X"1B",X"3B",X"1D",X"5B",X"1F",X"6C",X"21",X"65",X"23",X"53",X"25",X"28",X"27",
		X"F4",X"28",X"A5",X"2A",X"55",X"2C",X"E1",X"2D",X"8D",X"2F",X"71",X"31",X"D7",X"32",X"40",X"34",
		X"91",X"35",X"DD",X"36",X"17",X"38",X"49",X"39",X"6A",X"3A",X"85",X"3B",X"92",X"3C",X"95",X"3D",
		X"8E",X"3E",X"7C",X"3F",X"61",X"40",X"3D",X"41",X"0F",X"42",X"D8",X"42",X"9A",X"43",X"52",X"44",
		X"02",X"45",X"AB",X"45",X"4C",X"46",X"E6",X"46",X"78",X"47",X"02",X"48",X"89",X"48",X"06",X"49",
		X"7F",X"49",X"EF",X"49",X"5D",X"4A",X"C3",X"4A",X"24",X"4B",X"7E",X"4B",X"D8",X"4B",X"27",X"4C",
		X"74",X"4C",X"BC",X"4C",X"FF",X"4C",X"3D",X"4D",X"78",X"4D",X"AD",X"4D",X"E0",X"4D",X"0F",X"4E",
		X"39",X"4E",X"5F",X"4E",X"85",X"4E",X"A3",X"4E",X"C1",X"4E",X"D9",X"4E",X"F0",X"4E",X"04",X"4F",
		X"15",X"4F",X"21",X"4F",X"2E",X"4F",X"36",X"4F",X"3D",X"4F",X"3F",X"4F",X"41",X"4F",X"3E",X"4F",
		X"3C",X"4F",X"35",X"4F",X"2F",X"4F",X"24",X"4F",X"19",X"4F",X"0B",X"4F",X"FC",X"4E",X"EB",X"4E",
		X"D7",X"4E",X"C2",X"4E",X"AD",X"4E",X"94",X"4E",X"7D",X"4E",X"61",X"4E",X"48",X"4E",X"27",X"4E",
		X"11",X"4E",X"B9",X"4D",X"DA",X"4B",X"AE",X"48",X"B7",X"44",X"3D",X"40",X"7A",X"3B",X"8F",X"36",
		X"99",X"31",X"A7",X"2C",X"C3",X"27",X"F7",X"22",X"47",X"1E",X"B5",X"19",X"46",X"15",X"F4",X"10",
		X"C6",X"0C",X"B9",X"08",X"CD",X"04",X"01",X"01",X"55",X"FD",X"CA",X"F9",X"57",X"F6",X"07",X"F3",
		X"D0",X"EF",X"BA",X"EC",X"B6",X"E9",X"DB",X"E6",X"01",X"E4",X"15",X"E2",X"E7",X"E1",X"CA",X"E2",
		X"76",X"E4",X"95",X"E6",X"09",X"E9",X"A3",X"EB",X"5B",X"EE",X"16",X"F1",X"D4",X"F3",X"86",X"F6",
		X"2F",X"F9",X"C7",X"FB",X"4F",X"FE",X"C2",X"00",X"25",X"03",X"75",X"05",X"B1",X"07",X"D9",X"09",
		X"F3",X"0B",X"F9",X"0D",X"ED",X"0F",X"CF",X"11",X"A2",X"13",X"64",X"15",X"18",X"17",X"BC",X"18",
		X"50",X"1A",X"D7",X"1B",X"50",X"1D",X"BC",X"1E",X"1B",X"20",X"6C",X"21",X"B2",X"22",X"EB",X"23",
		X"18",X"25",X"3B",X"26",X"53",X"27",X"61",X"28",X"64",X"29",X"5E",X"2A",X"4D",X"2B",X"35",X"2C",
		X"11",X"2D",X"E8",X"2D",X"B1",X"2E",X"78",X"2F",X"33",X"30",X"EA",X"30",X"93",X"31",X"3C",X"32",
		X"D6",X"32",X"75",X"33",X"FE",X"33",X"98",X"34",X"84",X"34",X"C7",X"32",X"F1",X"2F",X"5E",X"2C",
		X"5E",X"28",X"17",X"24",X"B1",X"1F",X"40",X"1B",X"D4",X"16",X"76",X"12",X"2D",X"0E",X"FC",X"09",
		X"E7",X"05",X"F0",X"01",X"1A",X"FE",X"5F",X"FA",X"C3",X"F6",X"45",X"F3",X"E4",X"EF",X"A1",X"EC",
		X"77",X"E9",X"6A",X"E6",X"78",X"E3",X"9F",X"E0",X"DD",X"DD",X"38",X"DB",X"A8",X"D8",X"2E",X"D6",
		X"CC",X"D3",X"7F",X"D1",X"46",X"CF",X"23",X"CD",X"11",X"CB",X"14",X"C9",X"28",X"C7",X"51",X"C5",
		X"89",X"C3",X"D2",X"C1",X"2A",X"C0",X"94",X"BE",X"0D",X"BD",X"96",X"BB",X"2A",X"BA",X"CF",X"B8",
		X"7E",X"B7",X"3F",X"B6",X"09",X"B5",X"E2",X"B3",X"C4",X"B2",X"B5",X"B1",X"AC",X"B0",X"B6",X"AF",
		X"C0",X"AE",X"E2",X"AD",X"F8",X"AC",X"91",X"AC",X"D6",X"AD",X"4B",X"B0",X"86",X"B3",X"3D",X"B7",
		X"3F",X"BB",X"66",X"BF",X"A1",X"C3",X"D9",X"C7",X"08",X"CC",X"23",X"D0",X"29",X"D4",X"17",X"D8",
		X"E6",X"DB",X"9C",X"DF",X"35",X"E3",X"B3",X"E6",X"14",X"EA",X"5B",X"ED",X"85",X"F0",X"95",X"F3",
		X"8C",X"F6",X"6B",X"F9",X"30",X"FC",X"DF",X"FE",X"75",X"01",X"F7",X"03",X"63",X"06",X"B9",X"08",
		X"FB",X"0A",X"2B",X"0D",X"47",X"0F",X"51",X"11",X"48",X"13",X"2E",X"15",X"03",X"17",X"CA",X"18",
		X"7D",X"1A",X"23",X"1C",X"B9",X"1D",X"44",X"1F",X"BC",X"20",X"2A",X"22",X"86",X"23",X"DB",X"24",
		X"21",X"26",X"5E",X"27",X"8A",X"28",X"B0",X"29",X"C5",X"2A",X"D7",X"2B",X"D5",X"2C",X"D6",X"2D",
		X"BC",X"2E",X"B0",X"2F",X"A3",X"2F",X"F1",X"2D",X"43",X"2B",X"E2",X"27",X"21",X"24",X"1E",X"20",
		X"00",X"1C",X"D5",X"17",X"B1",X"13",X"99",X"0F",X"95",X"0B",X"AA",X"07",X"D9",X"03",X"22",X"00",
		X"8A",X"FC",X"0E",X"F9",X"AE",X"F5",X"68",X"F2",X"3F",X"EF",X"31",X"EC",X"3D",X"E9",X"64",X"E6",
		X"A1",X"E3",X"F9",X"E0",X"65",X"DE",X"EC",X"DB",X"82",X"D9",X"61",X"D7",X"D3",X"D6",X"AC",X"D7",
		X"66",X"D9",X"B9",X"DB",X"65",X"DE",X"4E",X"E1",X"53",X"E4",X"63",X"E7",X"76",X"EA",X"7F",X"ED",
		X"7C",X"F0",X"68",X"F3",X"42",X"F6",X"08",X"F9",X"B7",X"FB",X"53",X"FE",X"DB",X"00",X"4B",X"03",
		X"AA",X"05",X"F3",X"07",X"2A",X"0A",X"4B",X"0C",X"5F",X"0E",X"5A",X"10",X"4D",X"12",X"22",X"14",
		X"FB",X"15",X"02",X"17",X"4E",X"16",X"8E",X"14",X"09",X"12",X"15",X"0F",X"D5",X"0B",X"71",X"08",
		X"F8",X"04",X"80",X"01",X"0F",X"FE",X"AD",X"FA",X"5C",X"F7",X"20",X"F4",X"FB",X"F0",X"EF",X"ED",
		X"FA",X"EA",X"1D",X"E8",X"58",X"E5",X"AA",X"E2",X"15",X"E0",X"95",X"DD",X"29",X"DB",X"D6",X"D8",
		X"98",X"D6",X"6C",X"D4",X"55",X"D2",X"50",X"D0",X"5D",X"CE",X"7E",X"CC",X"AF",X"CA",X"F1",X"C8",
		X"44",X"C7",X"A5",X"C5",X"18",X"C4",X"99",X"C2",X"2A",X"C1",X"C4",X"BF",X"70",X"BE",X"27",X"BD",
		X"EE",X"BB",X"BD",X"BA",X"9C",X"B9",X"82",X"B8",X"78",X"B7",X"77",X"B6",X"82",X"B5",X"93",X"B4",
		X"B3",X"B3",X"D9",X"B2",X"0D",X"B2",X"43",X"B1",X"8A",X"B0",X"D0",X"AF",X"2B",X"AF",X"77",X"AE",
		X"63",X"AE",X"FD",X"AF",X"B5",X"B2",X"2F",X"B6",X"19",X"BA",X"4F",X"BE",X"A3",X"C2",X"06",X"C7",
		X"65",X"CB",X"BA",X"CF",X"F9",X"D3",X"22",X"D8",X"2F",X"DC",X"1E",X"E0",X"F1",X"E3",X"A7",X"E7",
		X"40",X"EB",X"BB",X"EE",X"1B",X"F2",X"5F",X"F5",X"87",X"F8",X"94",X"FB",X"88",X"FE",X"63",X"01",
		X"24",X"04",X"CF",X"06",X"63",X"09",X"E1",X"0B",X"49",X"0E",X"9E",X"10",X"D9",X"12",X"06",X"15",
		X"1D",X"17",X"24",X"19",X"16",X"1B",X"F9",X"1C",X"C9",X"1E",X"8B",X"20",X"39",X"22",X"DD",X"23",
		X"6E",X"25",X"F3",X"26",X"67",X"28",X"D0",X"29",X"2A",X"2B",X"7B",X"2C",X"B9",X"2D",X"F1",X"2E",
		X"19",X"30",X"3B",X"31",X"4B",X"32",X"58",X"33",X"54",X"34",X"4B",X"35",X"32",X"36",X"19",X"37",
		X"EC",X"37",X"C0",X"38",X"82",X"39",X"4A",X"3A",X"F0",X"3A",X"CD",X"3B",X"F5",X"3C",X"89",X"3D",
		X"2B",X"3E",X"BA",X"3E",X"4B",X"3F",X"CE",X"3F",X"51",X"40",X"C9",X"40",X"40",X"41",X"AC",X"41",
		X"16",X"42",X"79",X"42",X"D7",X"42",X"2F",X"43",X"86",X"43",X"D2",X"43",X"20",X"44",X"61",X"44",
		X"A9",X"44",X"E0",X"44",X"23",X"45",X"50",X"44",X"E0",X"41",X"81",X"3E",X"75",X"3A",X"0F",X"36",
		X"6E",X"31",X"B9",X"2C",X"F9",X"27",X"46",X"23",X"A4",X"1E",X"1D",X"1A",X"AF",X"15",X"62",X"11",
		X"31",X"0D",X"24",X"09",X"32",X"05",X"65",X"01",X"B4",X"FD",X"24",X"FA",X"B2",X"F6",X"5C",X"F3",
		X"23",X"F0",X"06",X"ED",X"05",X"EA",X"1B",X"E7",X"4D",X"E4",X"97",X"E1",X"F9",X"DE",X"71",X"DC",
		X"01",X"DA",X"A4",X"D7",X"62",X"D5",X"30",X"D3",X"13",X"D1",X"09",X"CF",X"14",X"CD",X"2D",X"CB",
		X"5B",X"C9",X"99",X"C7",X"E8",X"C5",X"45",X"C4",X"B5",X"C2",X"30",X"C1",X"BD",X"BF",X"57",X"BE",
		X"00",X"BD",X"B2",X"BB",X"77",X"BA",X"44",X"B9",X"20",X"B8",X"02",X"B7",X"F8",X"B5",X"EF",X"B4",
		X"01",X"B4",X"05",X"B3",X"F2",X"B2",X"91",X"B4",X"36",X"B7",X"95",X"BA",X"5B",X"BE",X"66",X"C2",
		X"8F",X"C6",X"C6",X"CA",X"F7",X"CE",X"1E",X"D3",X"30",X"D7",X"2D",X"DB",X"0D",X"DF",X"D4",X"E2",
		X"7D",X"E6",X"0C",X"EA",X"7C",X"ED",X"D3",X"F0",X"0D",X"F4",X"2E",X"F7",X"33",X"FA",X"20",X"FD",
		X"F3",X"FF",X"B0",X"02",X"52",X"05",X"DF",X"07",X"5B",X"0A",X"9D",X"0C",X"53",X"0D",X"95",X"0C",
		X"EF",X"0A",X"AC",X"08",X"08",X"06",X"29",X"03",X"2C",X"00",X"20",X"FD",X"16",X"FA",X"11",X"F7",
		X"1A",X"F4",X"35",X"F1",X"62",X"EE",X"A3",X"EB",X"F8",X"E8",X"66",X"E6",X"E6",X"E3",X"7D",X"E1",
		X"26",X"DF",X"E7",X"DC",X"B9",X"DA",X"A0",X"D8",X"96",X"D6",X"A7",X"D4",X"C0",X"D2",X"F6",X"D0",
		X"26",X"CF",X"17",X"CE",X"C2",X"CE",X"8C",X"D0",X"20",X"D3",X"27",X"D6",X"7F",X"D9",X"FB",X"DC",
		X"8C",X"E0",X"1E",X"E4",X"AE",X"E7",X"2B",X"EB",X"99",X"EE",X"EF",X"F1",X"31",X"F5",X"59",X"F8",
		X"68",X"FB",X"61",X"FE",X"40",X"01",X"08",X"04",X"B9",X"06",X"52",X"09",X"D7",X"0B",X"43",X"0E",
		X"9D",X"10",X"E2",X"12",X"14",X"15",X"2F",X"17",X"2E",X"19",X"CB",X"19",X"DA",X"18",X"FC",X"16",
		X"76",X"14",X"90",X"11",X"6A",X"0E",X"28",X"0B",X"D5",X"07",X"85",X"04",X"3E",X"01",X"04",X"FE",
		X"DD",X"FA",X"CA",X"F7",X"CD",X"F4",X"E6",X"F1",X"18",X"EF",X"60",X"EC",X"BF",X"E9",X"33",X"E7",
		X"C0",X"E4",X"60",X"E2",X"17",X"E0",X"DD",X"DD",X"BD",X"DB",X"AB",X"D9",X"B5",X"D7",X"BC",X"D5",
		X"55",X"D4",X"AA",X"D4",X"33",X"D6",X"8D",X"D8",X"67",X"DB",X"93",X"DE",X"EA",X"E1",X"5C",X"E5",
		X"CF",X"E8",X"40",X"EC",X"A4",X"EF",X"F7",X"F2",X"34",X"F6",X"5E",X"F9",X"70",X"FC",X"6B",X"FF",
		X"4B",X"02",X"16",X"05",X"C8",X"07",X"69",X"0A",X"EE",X"0C",X"60",X"0F",X"BB",X"11",X"04",X"14",
		X"35",X"16",X"58",X"18",X"60",X"1A",X"60",X"1C",X"27",X"1D",X"4B",X"1C",X"76",X"1A",X"EF",X"17",
		X"06",X"15",X"D4",X"11",X"89",X"0E",X"27",X"0B",X"CA",X"07",X"70",X"04",X"29",X"01",X"F1",X"FD",
		X"D4",X"FA",X"C6",X"F7",X"D3",X"F4",X"F4",X"F1",X"30",X"EF",X"7F",X"EC",X"E8",X"E9",X"65",X"E7",
		X"FB",X"E4",X"A4",X"E2",X"63",X"E0",X"34",X"DE",X"19",X"DC",X"11",X"DA",X"1B",X"D8",X"38",X"D6",
		X"67",X"D4",X"A3",X"D2",X"F3",X"D0",X"50",X"CF",X"BF",X"CD",X"3B",X"CC",X"C7",X"CA",X"5E",X"C9",
		X"07",X"C8",X"B9",X"C6",X"7B",X"C5",X"46",X"C4",X"1F",X"C3",X"02",X"C2",X"F2",X"C0",X"EC",X"BF",
		X"F1",X"BE",X"FE",X"BD",X"18",X"BD",X"3B",X"BC",X"68",X"BB",X"9A",X"BA",X"D8",X"B9",X"1D",X"B9",
		X"6D",X"B8",X"BD",X"B7",X"4E",X"B7",X"6D",X"B8",X"E7",X"BA",X"35",X"BE",X"0F",X"C2",X"38",X"C6",
		X"8F",X"CA",X"FA",X"CE",X"63",X"D3",X"C3",X"D7",X"11",X"DC",X"47",X"E0",X"63",X"E4",X"61",X"E8",
		X"44",X"EC",X"07",X"F0",X"AD",X"F3",X"37",X"F7",X"A2",X"FA",X"F4",X"FD",X"27",X"01",X"3E",X"04",
		X"3E",X"07",X"22",X"0A",X"EE",X"0C",X"A0",X"0F",X"3D",X"12",X"C3",X"14",X"34",X"17",X"8C",X"19",
		X"D2",X"1B",X"04",X"1E",X"21",X"20",X"2A",X"22",X"24",X"24",X"09",X"26",X"DF",X"27",X"A3",X"29",
		X"58",X"2B",X"FB",X"2C",X"91",X"2E",X"17",X"30",X"8E",X"31",X"F7",X"32",X"54",X"34",X"A3",X"35",
		X"E7",X"36",X"1D",X"38",X"48",X"39",X"66",X"3A",X"7A",X"3B",X"83",X"3C",X"81",X"3D",X"76",X"3E",
		X"60",X"3F",X"40",X"40",X"17",X"41",X"E5",X"41",X"AB",X"42",X"69",X"43",X"1D",X"44",X"C9",X"44",
		X"6E",X"45",X"0E",X"46",X"A4",X"46",X"34",X"47",X"BD",X"47",X"3E",X"48",X"BA",X"48",X"2E",X"49",
		X"9F",X"49",X"09",X"4A",X"6D",X"4A",X"CC",X"4A",X"25",X"4B",X"79",X"4B",X"C9",X"4B",X"13",X"4C",
		X"59",X"4C",X"9B",X"4C",X"D7",X"4C",X"11",X"4D",X"46",X"4D",X"77",X"4D",X"A4",X"4D",X"CD",X"4D",
		X"F2",X"4D",X"17",X"4E",X"33",X"4E",X"4F",X"4E",X"69",X"4E",X"7D",X"4E",X"90",X"4E",X"A0",X"4E",
		X"AC",X"4E",X"B7",X"4E",X"BF",X"4E",X"C3",X"4E",X"C7",X"4E",X"C7",X"4E",X"C6",X"4E",X"C1",X"4E",
		X"BB",X"4E",X"B2",X"4E",X"A9",X"4E",X"9E",X"4E",X"8F",X"4E",X"7F",X"4E",X"6E",X"4E",X"5A",X"4E",
		X"45",X"4E",X"30",X"4E",X"19",X"4E",X"FF",X"4D",X"E4",X"4D",X"CB",X"4D",X"AB",X"4D",X"8D",X"4D",
		X"6D",X"4D",X"4C",X"4D",X"2A",X"4D",X"06",X"4D",X"E3",X"4C",X"BD",X"4C",X"98",X"4C",X"71",X"4C",
		X"4A",X"4C",X"20",X"4C",X"F8",X"4B",X"CC",X"4B",X"A1",X"4B",X"75",X"4B",X"48",X"4B",X"1B",X"4B",
		X"EC",X"4A",X"BE",X"4A",X"8F",X"4A",X"60",X"4A",X"30",X"4A",X"FE",X"49",X"CE",X"49",X"9D",X"49",
		X"68",X"49",X"36",X"49",X"03",X"49",X"CF",X"48",X"9C",X"48",X"67",X"48",X"32",X"48",X"FC",X"47",
		X"C7",X"47",X"91",X"47",X"5B",X"47",X"24",X"47",X"F0",X"46",X"B8",X"46",X"82",X"46",X"4A",X"46",
		X"12",X"46",X"DB",X"45",X"A1",X"45",X"6A",X"45",X"32",X"45",X"FB",X"44",X"C1",X"44",X"89",X"44",
		X"51",X"44",X"17",X"44",X"DE",X"43",X"A5",X"43",X"6D",X"43",X"33",X"43",X"FA",X"42",X"C1",X"42",
		X"87",X"42",X"4E",X"42",X"14",X"42",X"DA",X"41",X"A0",X"41",X"67",X"41",X"2D",X"41",X"F3",X"40",
		X"BA",X"40",X"80",X"40",X"47",X"40",X"0D",X"40",X"D4",X"3F",X"9A",X"3F",X"61",X"3F",X"28",X"3F",
		X"EF",X"3E",X"B5",X"3E",X"7B",X"3E",X"41",X"3E",X"09",X"3E",X"CF",X"3D",X"97",X"3D",X"5D",X"3D",
		X"24",X"3D",X"EC",X"3C",X"B3",X"3C",X"79",X"3C",X"42",X"3C",X"09",X"3C",X"D0",X"3B",X"99",X"3B",
		X"60",X"3B",X"28",X"3B",X"EE",X"3A",X"B7",X"3A",X"7F",X"3A",X"48",X"3A",X"0F",X"3A",X"DA",X"39",
		X"A0",X"39",X"6A",X"39",X"33",X"39",X"FD",X"38",X"C2",X"38",X"90",X"38",X"51",X"38",X"98",X"37",
		X"2C",X"35",X"5C",X"31",X"FE",X"2C",X"2D",X"28",X"2E",X"23",X"10",X"1E",X"F5",X"18",X"E0",X"13",
		X"E4",X"0E",X"FF",X"09",X"3D",X"05",X"9B",X"00",X"1C",X"FC",X"BD",X"F7",X"85",X"F3",X"6B",X"EF",
		X"78",X"EB",X"A3",X"E7",X"F0",X"E3",X"5C",X"E0",X"E9",X"DC",X"92",X"D9",X"5C",X"D6",X"3F",X"D3",
		X"3F",X"D0",X"56",X"CD",X"8E",X"CA",X"D9",X"C7",X"3F",X"C5",X"BD",X"C2",X"53",X"C0",X"FC",X"BD",
		X"BE",X"BB",X"93",X"B9",X"7F",X"B7",X"7B",X"B5",X"8D",X"B3",X"AE",X"B1",X"E6",X"AF",X"2B",X"AE",
		X"85",X"AC",X"EB",X"AA",X"65",X"A9",X"EB",X"A7",X"83",X"A6",X"25",X"A5",X"DA",X"A3",X"97",X"A2",
		X"69",X"A1",X"40",X"A0",X"2B",X"9F",X"17",X"9E",X"20",X"9D",X"18",X"9C",X"D8",X"9B",X"51",X"9D",
		X"E3",X"9F",X"39",X"A3",X"FE",X"A6",X"0F",X"AB",X"3F",X"AF",X"81",X"B3",X"BD",X"B7",X"F1",X"BB",
		X"13",X"C0",X"1E",X"C4",X"0D",X"C8",X"E4",X"CB",X"9E",X"CF",X"3C",X"D3",X"BE",X"D6",X"25",X"DA",
		X"71",X"DD",X"A1",X"E0",X"B7",X"E3",X"B5",X"E6",X"98",X"E9",X"66",X"EC",X"18",X"EF",X"B8",X"F1",
		X"40",X"F4",X"A6",X"F6",X"98",X"F7",X"FD",X"F6",X"73",X"F5",X"3F",X"F3",X"A7",X"F0",X"CD",X"ED",
		X"D6",X"EA",X"CD",X"E7",X"C5",X"E4",X"C1",X"E1",X"CD",X"DE",X"E9",X"DB",X"18",X"D9",X"5B",X"D6",
		X"B4",X"D3",X"23",X"D1",X"A7",X"CE",X"41",X"CC",X"F0",X"C9",X"B3",X"C7",X"8A",X"C5",X"78",X"C3",
		X"75",X"C1",X"87",X"BF",X"A8",X"BD",X"E4",X"BB",X"1D",X"BA",X"F0",X"B8",X"82",X"B9",X"45",X"BB",
		X"DB",X"BD",X"EE",X"C0",X"54",X"C4",X"E5",X"C7",X"8D",X"CB",X"37",X"CF",X"DB",X"D2",X"73",X"D6",
		X"F9",X"D9",X"69",X"DD",X"C2",X"E0",X"03",X"E4",X"2B",X"E7",X"3D",X"EA",X"35",X"ED",X"13",X"F0",
		X"DC",X"F2",X"8D",X"F5",X"28",X"F8",X"AC",X"FA",X"1C",X"FD",X"77",X"FF",X"BC",X"01",X"EF",X"03",
		X"10",X"06",X"1E",X"08",X"1A",X"0A",X"04",X"0C",X"DD",X"0D",X"A9",X"0F",X"61",X"11",X"0D",X"13",
		X"A7",X"14",X"35",X"16",X"B4",X"17",X"26",X"19",X"8A",X"1A",X"E4",X"1B",X"2F",X"1D",X"70",X"1E",
		X"A4",X"1F",X"CD",X"20",X"EA",X"21",X"FF",X"22",X"05",X"24",X"07",X"25",X"FB",X"25",X"EA",X"26",
		X"C9",X"27",X"A8",X"28",X"75",X"29",X"49",X"2A",X"B5",X"2A",X"79",X"29",X"FB",X"26",X"AC",X"23",
		X"DB",X"1F",X"BD",X"1B",X"73",X"17",X"1D",X"13",X"C3",X"0E",X"78",X"0A",X"3D",X"06",X"1F",X"02",
		X"16",X"FE",X"2D",X"FA",X"60",X"F6",X"B5",X"F2",X"23",X"EF",X"B2",X"EB",X"5B",X"E8",X"21",X"E5",
		X"03",X"E2",X"FF",X"DE",X"19",X"DC",X"48",X"D9",X"94",X"D6",X"F6",X"D3",X"6F",X"D1",X"01",X"CF",
		X"A8",X"CC",X"64",X"CA",X"35",X"C8",X"1B",X"C6",X"12",X"C4",X"1E",X"C2",X"3B",X"C0",X"6D",X"BE",
		X"AC",X"BC",X"FE",X"BA",X"5F",X"B9",X"D2",X"B7",X"52",X"B6",X"E3",X"B4",X"80",X"B3",X"2E",X"B2",
		X"E5",X"B0",X"AD",X"AF",X"7E",X"AE",X"5F",X"AD",X"4A",X"AC",X"42",X"AB",X"43",X"AA",X"51",X"A9",
		X"67",X"A8",X"8B",X"A7",X"AF",X"A6",X"19",X"A6",X"15",X"A7",X"72",X"A9",X"A5",X"AC",X"68",X"B0",
		X"7D",X"B4",X"C1",X"B8",X"19",X"BD",X"75",X"C1",X"C5",X"C5",X"07",X"CA",X"2F",X"CE",X"41",X"D2",
		X"35",X"D6",X"0D",X"DA",X"C8",X"DD",X"67",X"E1",X"EA",X"E4",X"4F",X"E8",X"98",X"EB",X"C7",X"EE",
		X"DB",X"F1",X"D7",X"F4",X"B7",X"F7",X"7F",X"FA",X"32",X"FD",X"CC",X"FF",X"4F",X"02",X"BF",X"04",
		X"18",X"07",X"5F",X"09",X"90",X"0B",X"AE",X"0D",X"BB",X"0F",X"B6",X"11",X"9D",X"13",X"75",X"15",
		X"3D",X"17",X"F5",X"18",X"9D",X"1A",X"36",X"1C",X"C0",X"1D",X"3E",X"1F",X"AD",X"20",X"0F",X"22",
		X"64",X"23",X"AD",X"24",X"E9",X"25",X"19",X"27",X"41",X"28",X"5A",X"29",X"69",X"2A",X"6F",X"2B",
		X"6B",X"2C",X"5D",X"2D",X"46",X"2E",X"27",X"2F",X"FC",X"2F",X"CA",X"30",X"91",X"31",X"4F",X"32",
		X"05",X"33",X"B2",X"33",X"59",X"34",X"FA",X"34",X"93",X"35",X"25",X"36",X"B2",X"36",X"37",X"37",
		X"B7",X"37",X"2F",X"38",X"A5",X"38",X"15",X"39",X"7E",X"39",X"E1",X"39",X"3F",X"3A",X"9A",X"3A",
		X"EF",X"3A",X"41",X"3B",X"8C",X"3B",X"D7",X"3B",X"18",X"3C",X"4F",X"3C",X"36",X"3B",X"91",X"38",
		X"0E",X"35",X"EA",X"30",X"74",X"2C",X"C7",X"27",X"09",X"23",X"44",X"1E",X"90",X"19",X"EA",X"14",
		X"64",X"10",X"F6",X"0B",X"AA",X"07",X"7B",X"03",X"70",X"FF",X"81",X"FB",X"B7",X"F7",X"09",X"F4",
		X"7C",X"F0",X"0A",X"ED",X"B8",X"E9",X"83",X"E6",X"69",X"E3",X"6A",X"E0",X"85",X"DD",X"BB",X"DA",
		X"0A",X"D8",X"6E",X"D5",X"ED",X"D2",X"7F",X"D0",X"2A",X"CE",X"E9",X"CB",X"BD",X"C9",X"A5",X"C7",
		X"9F",X"C5",X"AF",X"C3",X"CF",X"C1",X"01",X"C0",X"45",X"BE",X"99",X"BC",X"FC",X"BA",X"70",X"B9",
		X"F2",X"B7",X"85",X"B6",X"23",X"B5",X"D1",X"B3",X"8B",X"B2",X"55",X"B1",X"28",X"B0",X"0A",X"AF",
		X"F4",X"AD",X"F0",X"AC",X"EE",X"AB",X"01",X"AB",X"14",X"AA",X"55",X"AA",X"38",X"AC",X"0D",X"AF",
		X"92",X"B2",X"76",X"B6",X"99",X"BA",X"D8",X"BE",X"20",X"C3",X"61",X"C7",X"96",X"CB",X"B5",X"CF",
		X"BE",X"D3",X"AB",X"D7",X"7E",X"DB",X"32",X"DF",X"C9",X"E2",X"47",X"E6",X"A9",X"E9",X"EC",X"EC",
		X"17",X"F0",X"26",X"F3",X"1D",X"F6",X"FB",X"F8",X"C0",X"FB",X"6D",X"FE",X"02",X"01",X"85",X"03",
		X"EF",X"05",X"45",X"08",X"86",X"0A",X"B6",X"0C",X"D0",X"0E",X"DC",X"10",X"CE",X"12",X"C3",X"14",
		X"C8",X"16",X"8D",X"18",X"49",X"1A",X"F1",X"1B",X"8E",X"1D",X"19",X"1F",X"98",X"20",X"06",X"22",
		X"6B",X"23",X"C0",X"24",X"0A",X"26",X"47",X"27",X"7A",X"28",X"9F",X"29",X"BD",X"2A",X"CC",X"2B",
		X"D3",X"2C",X"CD",X"2D",X"C0",X"2E",X"AB",X"2F",X"8A",X"30",X"61",X"31",X"2F",X"32",X"F6",X"32",
		X"B2",X"33",X"69",X"34",X"19",X"35",X"BF",X"35",X"60",X"36",X"F9",X"36",X"8C",X"37",X"16",X"38",
		X"9F",X"38",X"1D",X"39",X"96",X"39",X"09",X"3A",X"79",X"3A",X"E1",X"3A",X"47",X"3B",X"A4",X"3B",
		X"FE",X"3B",X"52",X"3C",X"A4",X"3C",X"EF",X"3C",X"38",X"3D",X"7A",X"3D",X"BE",X"3D",X"CF",X"3D",
		X"56",X"3C",X"77",X"39",X"C2",X"35",X"7C",X"31",X"E8",X"2C",X"26",X"28",X"55",X"23",X"87",X"1E",
		X"C3",X"19",X"17",X"15",X"85",X"10",X"0F",X"0C",X"B9",X"07",X"85",X"03",X"70",X"FF",X"7D",X"FB",
		X"AA",X"F7",X"F8",X"F3",X"63",X"F0",X"EF",X"EC",X"94",X"E9",X"5D",X"E6",X"3B",X"E3",X"3C",X"E0",
		X"4B",X"DD",X"86",X"DA",X"BF",X"D7",X"D6",X"D5",X"B8",X"D5",X"BD",X"D6",X"94",X"D8",X"E5",X"DA",
		X"8D",X"DD",X"5F",X"E0",X"4F",X"E3",X"43",X"E6",X"37",X"E9",X"20",X"EC",X"FE",X"EE",X"CC",X"F1",
		X"87",X"F4",X"2F",X"F7",X"C1",X"F9",X"40",X"FC",X"AA",X"FE",X"01",X"01",X"46",X"03",X"74",X"05",
		X"93",X"07",X"9F",X"09",X"99",X"0B",X"80",X"0D",X"5B",X"0F",X"22",X"11",X"C8",X"12",X"FA",X"12",
		X"A1",X"11",X"5D",X"0F",X"76",X"0C",X"2F",X"09",X"AE",X"05",X"11",X"02",X"6B",X"FE",X"C7",X"FA",
		X"2E",X"F7",X"A6",X"F3",X"35",X"F0",X"DB",X"EC",X"9A",X"E9",X"72",X"E6",X"61",X"E3",X"6B",X"E0",
		X"90",X"DD",X"C9",X"DA",X"21",X"D8",X"8A",X"D5",X"0E",X"D3",X"A4",X"D0",X"56",X"CE",X"16",X"CC",
		X"F6",X"C9",X"D2",X"C7",X"57",X"C6",X"A2",X"C6",X"21",X"C8",X"73",X"CA",X"47",X"CD",X"6E",X"D0",
		X"C2",X"D3",X"2E",X"D7",X"A0",X"DA",X"0F",X"DE",X"6F",X"E1",X"C1",X"E4",X"FD",X"E7",X"25",X"EB",
		X"37",X"EE",X"31",X"F1",X"14",X"F4",X"E0",X"F6",X"94",X"F9",X"34",X"FC",X"BB",X"FE",X"2F",X"01",
		X"8C",X"03",X"D7",X"05",X"0C",X"08",X"31",X"0A",X"3F",X"0C",X"3D",X"0E",X"EE",X"0E",X"F8",X"0D",
		X"0F",X"0C",X"72",X"09",X"74",X"06",X"2E",X"03",X"CC",X"FF",X"58",X"FC",X"E8",X"F8",X"7F",X"F5",
		X"26",X"F2",X"DF",X"EE",X"B0",X"EB",X"95",X"E8",X"96",X"E5",X"AC",X"E2",X"DC",X"DF",X"21",X"DD",
		X"80",X"DA",X"F5",X"D7",X"82",X"D5",X"20",X"D3",X"D8",X"D0",X"A4",X"CE",X"83",X"CC",X"76",X"CA",
		X"7C",X"C8",X"95",X"C6",X"BF",X"C4",X"FA",X"C2",X"47",X"C1",X"A3",X"BF",X"10",X"BE",X"8A",X"BC",
		X"14",X"BB",X"AE",X"B9",X"56",X"B8",X"09",X"B7",X"CC",X"B5",X"99",X"B4",X"72",X"B3",X"59",X"B2",
		X"4A",X"B1",X"47",X"B0",X"4D",X"AF",X"60",X"AE",X"7E",X"AD",X"A4",X"AC",X"D3",X"AB",X"0F",X"AB",
		X"4E",X"AA",X"9C",X"A9",X"EB",X"A8",X"4E",X"A8",X"A8",X"A7",X"18",X"A8",X"33",X"AA",X"4A",X"AD",
		X"15",X"B1",X"40",X"B5",X"AD",X"B9",X"30",X"BE",X"C1",X"C2",X"47",X"C7",X"C1",X"CB",X"22",X"D0",
		X"6A",X"D4",X"94",X"D8",X"A4",X"DC",X"95",X"E0",X"66",X"E4",X"19",X"E8",X"B0",X"EB",X"26",X"EF",
		X"82",X"F2",X"C3",X"F5",X"E8",X"F8",X"F0",X"FB",X"E1",X"FE",X"B7",X"01",X"76",X"04",X"1F",X"07",
		X"AE",X"09",X"29",X"0C",X"8D",X"0E",X"DE",X"10",X"19",X"13",X"42",X"15",X"57",X"17",X"5A",X"19",
		X"4A",X"1B",X"2A",X"1D",X"F8",X"1E",X"B7",X"20",X"66",X"22",X"05",X"24",X"94",X"25",X"17",X"27",
		X"8B",X"28",X"F2",X"29",X"4A",X"2B",X"98",X"2C",X"D5",X"2D",X"0D",X"2F",X"32",X"30",X"53",X"31",
		X"61",X"32",X"6F",X"33",X"62",X"34",X"66",X"35",X"81",X"35",X"E3",X"33",X"37",X"31",X"CD",X"2D",
		X"F9",X"29",X"DD",X"25",X"A4",X"21",X"5C",X"1D",X"1A",X"19",X"E3",X"14",X"C4",X"10",X"B9",X"0C",
		X"CD",X"08",X"F9",X"04",X"45",X"01",X"AB",X"FD",X"32",X"FA",X"D2",X"F6",X"8F",X"F3",X"6A",X"F0",
		X"5F",X"ED",X"6B",X"EA",X"95",X"E7",X"D6",X"E4",X"2F",X"E2",X"9E",X"DF",X"27",X"DD",X"C3",X"DA",
		X"75",X"D8",X"3D",X"D6",X"19",X"D4",X"07",X"D2",X"08",X"D0",X"1D",X"CE",X"43",X"CC",X"7B",X"CA",
		X"C2",X"C8",X"1A",X"C7",X"83",X"C5",X"F9",X"C3",X"80",X"C2",X"15",X"C1",X"B7",X"BF",X"66",X"BE",
		X"23",X"BD",X"ED",X"BB",X"C2",X"BA",X"A4",X"B9",X"91",X"B8",X"8A",X"B7",X"8E",X"B6",X"9A",X"B5",
		X"B2",X"B4",X"D3",X"B3",X"FF",X"B2",X"32",X"B2",X"70",X"B1",X"B6",X"B0",X"06",X"B0",X"5B",X"AF",
		X"BA",X"AE",X"21",X"AE",X"8F",X"AD",X"03",X"AD",X"80",X"AC",X"01",X"AC",X"8D",X"AB",X"1A",X"AB",
		X"B2",X"AA",X"4C",X"AA",X"F0",X"A9",X"94",X"A9",X"41",X"A9",X"F2",X"A8",X"AB",X"A8",X"64",X"A8",
		X"27",X"A8",X"E9",X"A7",X"B5",X"A7",X"7E",X"A7",X"59",X"A7",X"20",X"A7",X"71",X"A7",X"77",X"A9",
		X"AB",X"AC",X"A6",X"B0",X"18",X"B5",X"D1",X"B9",X"AD",X"BE",X"94",X"C3",X"75",X"C8",X"49",X"CD",
		X"02",X"D2",X"A3",X"D6",X"24",X"DB",X"85",X"DF",X"C6",X"E3",X"E8",X"E7",X"E5",X"EB",X"C7",X"EF",
		X"85",X"F3",X"27",X"F7",X"A8",X"FA",X"0E",X"FE",X"53",X"01",X"80",X"04",X"8F",X"07",X"89",X"0A",
		X"62",X"0D",X"29",X"10",X"AB",X"11",X"7C",X"11",X"4C",X"10",X"60",X"0E",X"0A",X"0C",X"68",X"09",
		X"A0",X"06",X"C3",X"03",X"E4",X"00",X"07",X"FE",X"34",X"FB",X"6F",X"F8",X"BB",X"F5",X"1A",X"F3",
		X"8B",X"F0",X"13",X"EE",X"AE",X"EB",X"5B",X"E9",X"1F",X"E7",X"F3",X"E4",X"DC",X"E2",X"D8",X"E0",
		X"E5",X"DE",X"05",X"DD",X"32",X"DB",X"76",X"D9",X"BD",X"D7",X"6B",X"D6",X"CE",X"D6",X"81",X"D8",
		X"10",X"DB",X"28",X"DE",X"94",X"E1",X"32",X"E5",X"E8",X"E8",X"A3",X"EC",X"59",X"F0",X"00",X"F4",
		X"94",X"F7",X"13",X"FB",X"7A",X"FE",X"C8",X"01",X"FD",X"04",X"18",X"08",X"1B",X"0B",X"01",X"0E",
		X"D4",X"10",X"89",X"13",X"2C",X"16",X"B2",X"18",X"2B",X"1B",X"84",X"1D",X"D2",X"1F",X"FF",X"21",
		X"2D",X"24",X"48",X"25",X"A8",X"24",X"FC",X"22",X"91",X"20",X"B6",X"1D",X"91",X"1A",X"43",X"17",
		X"F3",X"13",X"B7",X"10",X"4F",X"0D",X"FF",X"09",X"BB",X"06",X"8F",X"03",X"75",X"00",X"77",X"FD",
		X"8B",X"FA",X"BB",X"F7",X"00",X"F5",X"5C",X"F2",X"CD",X"EF",X"56",X"ED",X"F4",X"EA",X"A7",X"E8",
		X"6D",X"E6",X"48",X"E4",X"34",X"E2",X"36",X"E0",X"46",X"DE",X"6A",X"DC",X"9F",X"DA",X"E5",X"D8",
		X"39",X"D7",X"9D",X"D5",X"0F",X"D4",X"93",X"D2",X"23",X"D1",X"BF",X"CF",X"6B",X"CE",X"21",X"CD",
		X"E5",X"CB",X"B5",X"CA",X"91",X"C9",X"76",X"C8",X"6B",X"C7",X"65",X"C6",X"6E",X"C5",X"7D",X"C4",
		X"9A",X"C3",X"BB",X"C2",X"EB",X"C1",X"1F",X"C1",X"61",X"C0",X"A2",X"BF",X"FA",X"BE",X"3F",X"BE",
		X"60",X"BE",X"3A",X"C0",X"2C",X"C3",X"DC",X"C6",X"F9",X"CA",X"5F",X"CF",X"E1",X"D3",X"6F",X"D8",
		X"F7",X"DC",X"73",X"E1",X"D8",X"E5",X"24",X"EA",X"53",X"EE",X"62",X"F2",X"56",X"F6",X"29",X"FA",
		X"DD",X"FD",X"74",X"01",X"EC",X"04",X"46",X"08",X"87",X"0B",X"A9",X"0E",X"B2",X"11",X"9F",X"14",
		X"75",X"17",X"31",X"1A",X"D4",X"1C",X"60",X"1F",X"D7",X"21",X"37",X"24",X"82",X"26",X"B8",X"28",
		X"DB",X"2A",X"EA",X"2C",X"E5",X"2E",X"D0",X"30",X"A8",X"32",X"6F",X"34",X"26",X"36",X"CB",X"37",
		X"63",X"39",X"EB",X"3A",X"64",X"3C",X"CE",X"3D",X"2C",X"3F",X"7B",X"40",X"BF",X"41",X"F5",X"42",
		X"20",X"44",X"3C",X"45",X"4F",X"46",X"56",X"47",X"53",X"48",X"47",X"49",X"30",X"4A",X"0D",X"4B",
		X"E2",X"4B",X"AF",X"4C",X"71",X"4D",X"2B",X"4E",X"DD",X"4E",X"87",X"4F",X"28",X"50",X"C4",X"50",
		X"57",X"51",X"E1",X"51",X"66",X"52",X"E6",X"52",X"5D",X"53",X"D0",X"53",X"39",X"54",X"A0",X"54",
		X"FF",X"54",X"58",X"55",X"AD",X"55",X"FD",X"55",X"48",X"56",X"8C",X"56",X"CE",X"56",X"0A",X"57",
		X"43",X"57",X"76",X"57",X"A5",X"57",X"D1",X"57",X"F7",X"57",X"1D",X"58",X"3C",X"58",X"59",X"58",
		X"71",X"58",X"88",X"58",X"9B",X"58",X"AB",X"58",X"B6",X"58",X"C1",X"58",X"C6",X"58",X"CC",X"58",
		X"CB",X"58",X"CD",X"58",X"C8",X"58",X"C3",X"58",X"B9",X"58",X"AF",X"58",X"A2",X"58",X"95",X"58",
		X"82",X"58",X"73",X"58",X"5C",X"58",X"49",X"58",X"2B",X"58",X"1E",X"58",X"A0",X"57",X"6F",X"55",
		X"04",X"52",X"CF",X"4D",X"1D",X"49",X"24",X"44",X"08",X"3F",X"E1",X"39",X"C0",X"34",X"B2",X"2F",
		X"B8",X"2A",X"E0",X"25",X"26",X"21",X"8E",X"1C",X"19",X"18",X"C4",X"13",X"95",X"0F",X"87",X"0B",
		X"99",X"07",X"CE",X"03",X"21",X"00",X"93",X"FC",X"24",X"F9",X"D3",X"F5",X"9D",X"F2",X"84",X"EF",
		X"84",X"EC",X"A1",X"E9",X"D5",X"E6",X"22",X"E4",X"87",X"E1",X"05",X"DF",X"96",X"DC",X"3F",X"DA",
		X"FC",X"D7",X"CD",X"D5",X"B2",X"D3",X"AC",X"D1",X"B7",X"CF",X"D4",X"CD",X"01",X"CC",X"42",X"CA",
		X"92",X"C8",X"F4",X"C6",X"63",X"C5",X"E2",X"C3",X"70",X"C2",X"0B",X"C1",X"B4",X"BF",X"69",X"BE",
		X"2B",X"BD",X"FC",X"BB",X"D8",X"BA",X"BF",X"B9",X"B1",X"B8",X"AF",X"B7",X"B7",X"B6",X"C9",X"B5",
		X"E5",X"B4",X"0C",X"B4",X"3C",X"B3",X"76",X"B2",X"B7",X"B1",X"01",X"B1",X"53",X"B0",X"AE",X"AF",
		X"10",X"AF",X"79",X"AE",X"EA",X"AD",X"64",X"AD",X"E1",X"AC",X"68",X"AC",X"F4",X"AB",X"87",X"AB",
		X"1E",X"AB",X"BF",X"AA",X"5F",X"AA",X"0C",X"AA",X"B8",X"A9",X"70",X"A9",X"22",X"A9",X"E9",X"A8",
		X"9D",X"A8",X"3E",X"A9",X"96",X"AB",X"F6",X"AE",X"11",X"B3",X"91",X"B7",X"53",X"BC",X"2D",X"C1",
		X"13",X"C6",X"EE",X"CA",X"B9",X"CF",X"6A",X"D4",X"01",X"D9",X"77",X"DD",X"D1",X"E1",X"06",X"E6",
		X"1E",X"EA",X"11",X"EE",X"E7",X"F1",X"9D",X"F5",X"33",X"F9",X"AD",X"FC",X"08",X"00",X"47",X"03",
		X"6C",X"06",X"74",X"09",X"62",X"0C",X"37",X"0F",X"F3",X"11",X"98",X"14",X"26",X"17",X"9C",X"19",
		X"01",X"1C",X"4B",X"1E",X"84",X"20",X"A7",X"22",X"B9",X"24",X"B8",X"26",X"A2",X"28",X"7D",X"2A",
		X"47",X"2C",X"01",X"2E",X"AA",X"2F",X"43",X"31",X"CE",X"32",X"4A",X"34",X"B8",X"35",X"18",X"37",
		X"6D",X"38",X"B2",X"39",X"EA",X"3A",X"18",X"3C",X"3B",X"3D",X"50",X"3E",X"5D",X"3F",X"5F",X"40",
		X"53",X"41",X"41",X"42",X"23",X"43",X"FD",X"43",X"CC",X"44",X"93",X"45",X"51",X"46",X"08",X"47",
		X"B6",X"47",X"5E",X"48",X"FC",X"48",X"94",X"49",X"24",X"4A",X"AE",X"4A",X"31",X"4B",X"AD",X"4B",
		X"22",X"4C",X"92",X"4C",X"FD",X"4C",X"61",X"4D",X"C1",X"4D",X"1A",X"4E",X"6E",X"4E",X"BD",X"4E",
		X"09",X"4F",X"4F",X"4F",X"90",X"4F",X"CC",X"4F",X"05",X"50",X"3B",X"50",X"6B",X"50",X"96",X"50",
		X"BF",X"50",X"E4",X"50",X"06",X"51",X"25",X"51",X"40",X"51",X"58",X"51",X"6B",X"51",X"7E",X"51",
		X"8C",X"51",X"97",X"51",X"A3",X"51",X"A8",X"51",X"AE",X"51",X"AF",X"51",X"AE",X"51",X"AB",X"51",
		X"A6",X"51",X"9E",X"51",X"96",X"51",X"89",X"51",X"7C",X"51",X"6F",X"51",X"5C",X"51",X"49",X"51",
		X"36",X"51",X"1E",X"51",X"07",X"51",X"EE",X"50",X"D3",X"50",X"B8",X"50",X"9B",X"50",X"7C",X"50",
		X"5B",X"50",X"3B",X"50",X"19",X"50",X"F4",X"4F",X"D1",X"4F",X"AB",X"4F",X"84",X"4F",X"5C",X"4F",
		X"34",X"4F",X"0A",X"4F",X"E0",X"4E",X"B4",X"4E",X"88",X"4E",X"5D",X"4E",X"2E",X"4E",X"00",X"4E",
		X"D1",X"4D",X"A1",X"4D",X"73",X"4D",X"41",X"4D",X"0F",X"4D",X"DD",X"4C",X"AB",X"4C",X"79",X"4C",
		X"44",X"4C",X"11",X"4C",X"DB",X"4B",X"A7",X"4B",X"70",X"4B",X"3B",X"4B",X"05",X"4B",X"CF",X"4A",
		X"96",X"4A",X"61",X"4A",X"2A",X"4A",X"F2",X"49",X"B7",X"49",X"82",X"49",X"47",X"49",X"11",X"49",
		X"D5",X"48",X"9F",X"48",X"61",X"48",X"2D",X"48",X"ED",X"47",X"BE",X"47",X"85",X"46",X"A0",X"43",
		X"C3",X"3F",X"36",X"3B",X"4D",X"36",X"2A",X"31",X"F1",X"2B",X"B4",X"26",X"86",X"21",X"6C",X"1C",
		X"70",X"17",X"90",X"12",X"D6",X"0D",X"3B",X"09",X"C5",X"04",X"73",X"00",X"46",X"FC",X"38",X"F8",
		X"4D",X"F4",X"83",X"F0",X"DB",X"EC",X"51",X"E9",X"E5",X"E5",X"98",X"E2",X"67",X"DF",X"53",X"DC",
		X"56",X"D9",X"AB",X"D6",X"B0",X"D5",X"28",X"D6",X"8E",X"D7",X"8F",X"D9",X"FA",X"DB",X"9B",X"DE",
		X"67",X"E1",X"2B",X"E4",X"CF",X"E6",X"B0",X"E9",X"7C",X"EC",X"41",X"EF",X"EF",X"F1",X"8D",X"F4",
		X"18",X"F7",X"90",X"F9",X"F6",X"FB",X"44",X"FE",X"82",X"00",X"AC",X"02",X"C6",X"04",X"C9",X"06",
		X"C1",X"08",X"A2",X"0A",X"7A",X"0C",X"36",X"0E",X"F9",X"0F",X"D3",X"10",X"E5",X"0F",X"DD",X"0D",
		X"0B",X"0B",X"C7",X"07",X"36",X"04",X"82",X"00",X"BC",X"FC",X"F6",X"F8",X"37",X"F5",X"8B",X"F1",
		X"F0",X"ED",X"72",X"EA",X"08",X"E7",X"BB",X"E3",X"88",X"E0",X"6E",X"DD",X"70",X"DA",X"8B",X"D7",
		X"BF",X"D4",X"0C",X"D2",X"71",X"CF",X"EE",X"CC",X"80",X"CA",X"28",X"C8",X"E8",X"C5",X"BB",X"C3",
		X"A4",X"C1",X"9C",X"BF",X"AB",X"BD",X"CC",X"BB",X"FE",X"B9",X"41",X"B8",X"96",X"B6",X"F9",X"B4",
		X"6F",X"B3",X"F2",X"B1",X"86",X"B0",X"24",X"AF",X"D5",X"AD",X"8D",X"AC",X"59",X"AB",X"2E",X"AA",
		X"11",X"A9",X"FE",X"A7",X"FA",X"A6",X"FD",X"A5",X"10",X"A5",X"28",X"A4",X"50",X"A3",X"79",X"A2",
		X"B7",X"A1",X"F1",X"A0",X"44",X"A0",X"85",X"9F",X"7B",X"9F",X"34",X"A1",X"16",X"A4",X"C2",X"A7",
		X"E4",X"AB",X"50",X"B0",X"E2",X"B4",X"7E",X"B9",X"19",X"BE",X"A8",X"C2",X"1F",X"C7",X"82",X"CB",
		X"C4",X"CF",X"EB",X"D3",X"F0",X"D7",X"DC",X"DB",X"A6",X"DF",X"52",X"E3",X"DF",X"E6",X"52",X"EA",
		X"A6",X"ED",X"E0",X"F0",X"FE",X"F3",X"04",X"F7",X"ED",X"F9",X"C1",X"FC",X"77",X"FF",X"13",X"02",
		X"46",X"03",X"D2",X"02",X"61",X"01",X"3A",X"FF",X"AA",X"FC",X"D2",X"F9",X"D9",X"F6",X"CC",X"F3",
		X"BE",X"F0",X"B4",X"ED",X"B8",X"EA",X"CB",X"E7",X"F1",X"E4",X"2C",X"E2",X"7D",X"DF",X"E2",X"DC",
		X"5C",X"DA",X"EE",X"D7",X"94",X"D5",X"51",X"D3",X"1E",X"D1",X"01",X"CF",X"F6",X"CC",X"02",X"CB",
		X"18",X"C9",X"4C",X"C7",X"7B",X"C5",X"36",X"C4",X"B6",X"C4",X"7D",X"C6",X"1F",X"C9",X"48",X"CC",
		X"C7",X"CF",X"74",X"D3",X"38",X"D7",X"02",X"DB",X"C4",X"DE",X"7A",X"E2",X"1D",X"E6",X"A9",X"E9",
		X"1D",X"ED",X"79",X"F0",X"BC",X"F3",X"E3",X"F6",X"F2",X"F9",X"E6",X"FC",X"C5",X"FF",X"89",X"02",
		X"39",X"05",X"CC",X"07",X"50",X"0A",X"B7",X"0C",X"13",X"0F",X"4F",X"11",X"84",X"13",X"80",X"14",
		X"C3",X"13",X"01",X"12",X"80",X"0F",X"95",X"0C",X"5F",X"09",X"08",X"06",X"A0",X"02",X"35",X"FF",
		X"D3",X"FB",X"80",X"F8",X"3C",X"F5",X"10",X"F2",X"F8",X"EE",X"F9",X"EB",X"11",X"E9",X"43",X"E6",
		X"8A",X"E3",X"E9",X"E0",X"60",X"DE",X"EB",X"DB",X"8D",X"D9",X"44",X"D7",X"11",X"D5",X"EE",X"D2",
		X"E4",X"D0",X"E1",X"CE",X"3F",X"CD",X"55",X"CD",X"CC",X"CE",X"26",X"D1",X"14",X"D4",X"5D",X"D7",
		X"D9",X"DA",X"71",X"DE",X"11",X"E2",X"AE",X"E5",X"3D",X"E9",X"BE",X"EC",X"26",X"F0",X"7B",X"F3",
		X"B6",X"F6",X"D8",X"F9",X"E4",X"FC",X"D6",X"FF",X"AD",X"02",X"73",X"05",X"1A",X"08",X"B1",X"0A",
		X"2C",X"0D",X"97",X"0F",X"E8",X"11",X"2E",X"14",X"4F",X"16",X"77",X"18",X"97",X"19",X"EF",X"18",
		X"32",X"17",X"AF",X"14",X"BB",X"11",X"78",X"0E",X"12",X"0B",X"94",X"07",X"19",X"04",X"A0",X"00",
		X"3A",X"FD",X"E2",X"F9",X"A2",X"F6",X"78",X"F3",X"67",X"F0",X"6C",X"ED",X"8A",X"EA",X"C1",X"E7",
		X"0F",X"E5",X"74",X"E2",X"F2",X"DF",X"82",X"DD",X"2B",X"DB",X"E6",X"D8",X"B8",X"D6",X"9E",X"D4",
		X"92",X"D2",X"C4",X"D0",X"90",X"D0",X"DE",X"D1",X"12",X"D4",X"EA",X"D6",X"1D",X"DA",X"8E",X"DD",
		X"17",X"E1",X"B0",X"E4",X"41",X"E8",X"CB",X"EB",X"45",X"EF",X"AA",X"F2",X"F8",X"F5",X"30",X"F9",
		X"4D",X"FC",X"55",X"FF",X"40",X"02",X"16",X"05",X"D3",X"07",X"7C",X"0A",X"0C",X"0D",X"87",X"0F",
		X"EA",X"11",X"3C",X"14",X"76",X"16",X"A0",X"18",X"B2",X"1A",X"B6",X"1C",X"A6",X"1E",X"85",X"20",
		X"53",X"22",X"12",X"24",X"BF",X"25",X"5E",X"27",X"EE",X"28",X"70",X"2A",X"E2",X"2B",X"47",X"2D",
		X"A0",X"2E",X"EC",X"2F",X"2A",X"31",X"5D",X"32",X"83",X"33",X"A0",X"34",X"B2",X"35",X"B7",X"36",
		X"B3",X"37",X"A6",X"38",X"90",X"39",X"6E",X"3A",X"45",X"3B",X"0F",X"3C",X"D5",X"3C",X"92",X"3D",
		X"36",X"3E",X"6D",X"3D",X"14",X"3B",X"D4",X"37",X"F0",X"33",X"B3",X"2F",X"3F",X"2B",X"B4",X"26",
		X"25",X"22",X"A0",X"1D",X"2B",X"19",X"D0",X"14",X"8F",X"10",X"69",X"0C",X"64",X"08",X"7D",X"04",
		X"B6",X"00",X"0D",X"FD",X"83",X"F9",X"15",X"F6",X"C7",X"F2",X"92",X"EF",X"7C",X"EC",X"7B",X"E9",
		X"9C",X"E6",X"CD",X"E3",X"22",X"E1",X"7A",X"DE",X"78",X"DC",X"48",X"DC",X"5B",X"DD",X"47",X"DF",
		X"BF",X"E1",X"8D",X"E4",X"8E",X"E7",X"A9",X"EA",X"CE",X"ED",X"F0",X"F0",X"0B",X"F4",X"16",X"F7",
		X"10",X"FA",X"F6",X"FC",X"C7",X"FF",X"81",X"02",X"28",X"05",X"B8",X"07",X"37",X"0A",X"9B",X"0C",
		X"ED",X"0E",X"2A",X"11",X"57",X"13",X"6B",X"15",X"76",X"17",X"65",X"19",X"52",X"1B",X"C5",X"1C",
		X"74",X"1C",X"D5",X"1A",X"5B",X"18",X"53",X"15",X"F5",X"11",X"67",X"0E",X"C1",X"0A",X"16",X"07",
		X"6F",X"03",X"D7",X"FF",X"50",X"FC",X"E0",X"F8",X"87",X"F5",X"48",X"F2",X"21",X"EF",X"15",X"EC",
		X"20",X"E9",X"46",X"E6",X"82",X"E3",X"D9",X"E0",X"43",X"DE",X"C8",X"DB",X"60",X"D9",X"11",X"D7",
		X"D2",X"D4",X"B1",X"D2",X"92",X"D0",X"9B",X"CF",X"66",X"D0",X"39",X"D2",X"CE",X"D4",X"CF",X"D7",
		X"1E",X"DB",X"8D",X"DE",X"11",X"E2",X"93",X"E5",X"12",X"E9",X"7E",X"EC",X"DC",X"EF",X"22",X"F3",
		X"54",X"F6",X"6B",X"F9",X"6E",X"FC",X"56",X"FF",X"27",X"02",X"E0",X"04",X"84",X"07",X"0F",X"0A",
		X"88",X"0C",X"E9",X"0E",X"37",X"11",X"6F",X"13",X"96",X"15",X"A7",X"17",X"A8",X"19",X"96",X"1B",
		X"75",X"1D",X"40",X"1F",X"FD",X"20",X"A9",X"22",X"47",X"24",X"D4",X"25",X"54",X"27",X"C6",X"28",
		X"2D",X"2A",X"82",X"2B",X"CE",X"2C",X"0B",X"2E",X"3E",X"2F",X"65",X"30",X"81",X"31",X"90",X"32",
		X"9A",X"33",X"93",X"34",X"86",X"35",X"6E",X"36",X"4F",X"37",X"23",X"38",X"F3",X"38",X"B6",X"39",
		X"74",X"3A",X"26",X"3B",X"D7",X"3B",X"79",X"3C",X"1C",X"3D",X"AF",X"3D",X"46",X"3E",X"C9",X"3E",
		X"56",X"3F",X"C3",X"3F",X"6B",X"40",X"63",X"41",X"C5",X"41",X"34",X"42",X"90",X"42",X"F2",X"42",
		X"47",X"43",X"9B",X"43",X"E7",X"43",X"34",X"44",X"77",X"44",X"B9",X"44",X"F6",X"44",X"2F",X"45",
		X"63",X"45",X"96",X"45",X"C3",X"45",X"EE",X"45",X"15",X"46",X"38",X"46",X"57",X"46",X"76",X"46",
		X"90",X"46",X"A7",X"46",X"BB",X"46",X"CC",X"46",X"DC",X"46",X"EA",X"46",X"F3",X"46",X"FB",X"46",
		X"00",X"47",X"04",X"47",X"04",X"47",X"03",X"47",X"01",X"47",X"FC",X"46",X"F6",X"46",X"EC",X"46",
		X"E2",X"46",X"D7",X"46",X"C9",X"46",X"B9",X"46",X"A8",X"46",X"95",X"46",X"82",X"46",X"6D",X"46",
		X"56",X"46",X"3F",X"46",X"26",X"46",X"0B",X"46",X"F0",X"45",X"D2",X"45",X"B6",X"45",X"96",X"45",
		X"77",X"45",X"56",X"45",X"35",X"45",X"13",X"45",X"F1",X"44",X"CC",X"44",X"A7",X"44",X"81",X"44",
		X"5C",X"44",X"34",X"44",X"0C",X"44",X"E2",X"43",X"BB",X"43",X"90",X"43",X"68",X"43",X"3A",X"43",
		X"11",X"43",X"E3",X"42",X"B9",X"42",X"89",X"42",X"55",X"42",X"BE",X"40",X"97",X"3D",X"8A",X"39",
		X"D8",X"34",X"D3",X"2F",X"9A",X"2A",X"50",X"25",X"06",X"20",X"CD",X"1A",X"AA",X"15",X"A3",X"10",
		X"BE",X"0B",X"FC",X"06",X"5C",X"02",X"E2",X"FD",X"8D",X"F9",X"57",X"F5",X"48",X"F1",X"58",X"ED",
		X"8D",X"E9",X"E0",X"E5",X"56",X"E2",X"E7",X"DE",X"99",X"DB",X"63",X"D8",X"54",X"D5",X"4B",X"D2",
		X"E0",X"CF",X"4B",X"CF",X"06",X"D0",X"A5",X"D1",X"D1",X"D3",X"5F",X"D6",X"20",X"D9",X"02",X"DC",
		X"ED",X"DE",X"DD",X"E1",X"C4",X"E4",X"A1",X"E7",X"6D",X"EA",X"28",X"ED",X"CE",X"EF",X"64",X"F2",
		X"E3",X"F4",X"4F",X"F7",X"A6",X"F9",X"EE",X"FB",X"1E",X"FE",X"40",X"00",X"4C",X"02",X"4B",X"04",
		X"33",X"06",X"13",X"08",X"D8",X"09",X"97",X"0B",X"18",X"0C",X"E1",X"0A",X"AB",X"08",X"B8",X"05",
		X"5F",X"02",X"C0",X"FE",X"03",X"FB",X"35",X"F7",X"6E",X"F3",X"AD",X"EF",X"00",X"EC",X"67",X"E8",
		X"E8",X"E4",X"82",X"E1",X"35",X"DE",X"04",X"DB",X"ED",X"D7",X"F2",X"D4",X"11",X"D2",X"47",X"CF",
		X"96",X"CC",X"FF",X"C9",X"7F",X"C7",X"16",X"C5",X"BF",X"C2",X"85",X"C0",X"51",X"BE",X"88",X"BC",
		X"81",X"BC",X"DD",X"BD",X"1E",X"C0",X"F3",X"C2",X"25",X"C6",X"8D",X"C9",X"10",X"CD",X"9D",X"D0",
		X"28",X"D4",X"A8",X"D7",X"17",X"DB",X"73",X"DE",X"B9",X"E1",X"E6",X"E4",X"FE",X"E7",X"FD",X"EA",
		X"E5",X"ED",X"B6",X"F0",X"70",X"F3",X"11",X"F6",X"9F",X"F8",X"13",X"FB",X"7A",X"FD",X"C4",X"FF",
		X"03",X"02",X"23",X"04",X"45",X"06",X"57",X"07",X"9C",X"06",X"D2",X"04",X"3D",X"02",X"3D",X"FF",
		X"EC",X"FB",X"78",X"F8",X"ED",X"F4",X"67",X"F1",X"E4",X"ED",X"75",X"EA",X"12",X"E7",X"CB",X"E3",
		X"9A",X"E0",X"81",X"DD",X"7F",X"DA",X"9A",X"D7",X"CA",X"D4",X"14",X"D2",X"77",X"CF",X"EF",X"CC",
		X"7E",X"CA",X"25",X"C8",X"DF",X"C5",X"B0",X"C3",X"94",X"C1",X"8D",X"BF",X"98",X"BD",X"B6",X"BB",
		X"E4",X"B9",X"27",X"B8",X"78",X"B6",X"D9",X"B4",X"4D",X"B3",X"CD",X"B1",X"5E",X"B0",X"FC",X"AE",
		X"A9",X"AD",X"64",X"AC",X"2C",X"AB",X"00",X"AA",X"E0",X"A8",X"CC",X"A7",X"C4",X"A6",X"C8",X"A5",
		X"D8",X"A4",X"F0",X"A3",X"13",X"A3",X"41",X"A2",X"77",X"A1",X"B7",X"A0",X"01",X"A0",X"54",X"9F",
		X"AE",X"9E",X"10",X"9E",X"7A",X"9D",X"ED",X"9C",X"67",X"9C",X"E9",X"9B",X"70",X"9B",X"00",X"9B",
		X"95",X"9A",X"31",X"9A",X"D3",X"99",X"7B",X"99",X"28",X"99",X"DB",X"98",X"95",X"98",X"53",X"98",
		X"18",X"98",X"E0",X"97",X"AA",X"97",X"7D",X"97",X"52",X"97",X"2D",X"97",X"0B",X"97",X"EF",X"96",
		X"D3",X"96",X"C0",X"96",X"AD",X"96",X"9F",X"96",X"94",X"96",X"8C",X"96",X"87",X"96",X"86",X"96",
		X"88",X"96",X"8C",X"96",X"93",X"96",X"9E",X"96",X"AB",X"96",X"B9",X"96",X"CB",X"96",X"E0",X"96",
		X"F5",X"96",X"0F",X"97",X"29",X"97",X"47",X"97",X"63",X"97",X"86",X"97",X"A7",X"97",X"CE",X"97",
		X"F1",X"97",X"1B",X"98",X"42",X"98",X"71",X"98",X"9A",X"98",X"CB",X"98",X"F5",X"98",X"2D",X"99",
		X"4F",X"99",X"0D",X"9A",X"8C",X"9C",X"38",X"A0",X"AC",X"A4",X"94",X"A9",X"C3",X"AE",X"0F",X"B4",
		X"66",X"B9",X"B3",X"BE",X"EF",X"C3",X"0F",X"C9",X"13",X"CE",X"F4",X"D2",X"B3",X"D7",X"50",X"DC",
		X"C7",X"E0",X"19",X"E5",X"4D",X"E9",X"5C",X"ED",X"4A",X"F1",X"16",X"F5",X"C4",X"F8",X"53",X"FC",
		X"C0",X"FF",X"14",X"03",X"4B",X"06",X"66",X"09",X"66",X"0C",X"4E",X"0F",X"19",X"12",X"D0",X"14",
		X"6D",X"17",X"F3",X"19",X"63",X"1C",X"BD",X"1E",X"03",X"21",X"35",X"23",X"52",X"25",X"5C",X"27",
		X"54",X"29",X"3B",X"2B",X"0E",X"2D",X"D4",X"2E",X"85",X"30",X"2A",X"32",X"BD",X"33",X"44",X"35",
		X"B8",X"36",X"24",X"38",X"7D",X"39",X"CF",X"3A",X"0C",X"3C",X"46",X"3D",X"67",X"3E",X"8E",X"3F",
		X"87",X"3F",X"C9",X"3D",X"07",X"3B",X"8B",X"37",X"AB",X"33",X"85",X"2F",X"42",X"2B",X"F4",X"26",
		X"AA",X"22",X"6D",X"1E",X"48",X"1A",X"39",X"16",X"46",X"12",X"6D",X"0E",X"B3",X"0A",X"16",X"07",
		X"96",X"03",X"32",X"00",X"EA",X"FC",X"BE",X"F9",X"AE",X"F6",X"B7",X"F3",X"D8",X"F0",X"16",X"EE",
		X"69",X"EB",X"D6",X"E8",X"50",X"E6",X"29",X"E4",X"BC",X"E3",X"BF",X"E4",X"AA",X"E6",X"31",X"E9",
		X"16",X"EC",X"33",X"EF",X"6E",X"F2",X"B7",X"F5",X"FE",X"F8",X"39",X"FC",X"68",X"FF",X"83",X"02",
		X"8C",X"05",X"7E",X"08",X"5B",X"0B",X"1E",X"0E",X"CC",X"10",X"63",X"13",X"E7",X"15",X"50",X"18",
		X"AA",X"1A",X"EB",X"1C",X"1C",X"1F",X"34",X"21",X"42",X"23",X"30",X"25",X"23",X"27",X"18",X"28",
		X"3E",X"27",X"4C",X"25",X"92",X"22",X"66",X"1F",X"EA",X"1B",X"4C",X"18",X"96",X"14",X"E4",X"10",
		X"37",X"0D",X"9D",X"09",X"13",X"06",X"A1",X"02",X"47",X"FF",X"08",X"FC",X"E0",X"F8",X"D2",X"F5",
		X"DD",X"F2",X"02",X"F0",X"3C",X"ED",X"92",X"EA",X"FD",X"E7",X"7E",X"E5",X"15",X"E3",X"C3",X"E0",
		X"86",X"DE",X"57",X"DC",X"64",X"DA",X"0C",X"DA",X"3F",X"DB",X"5A",X"DD",X"21",X"E0",X"3F",X"E3",
		X"A2",X"E6",X"1A",X"EA",X"A9",X"ED",X"22",X"F1",X"8B",X"F4",X"01",X"F8",X"63",X"FB",X"AF",X"FE",
		X"E0",X"01",X"FD",X"04",X"00",X"08",X"EA",X"0A",X"BC",X"0D",X"76",X"10",X"1A",X"13",X"A8",X"15",
		X"1E",X"18",X"7D",X"1A",X"CB",X"1C",X"01",X"1F",X"27",X"21",X"36",X"23",X"36",X"25",X"21",X"27",
		X"FD",X"28",X"C5",X"2A",X"81",X"2C",X"28",X"2E",X"C2",X"2F",X"4E",X"31",X"C9",X"32",X"38",X"34",
		X"98",X"35",X"EC",X"36",X"32",X"38",X"6C",X"39",X"9A",X"3A",X"BD",X"3B",X"D4",X"3C",X"E0",X"3D",
		X"E1",X"3E",X"D7",X"3F",X"C5",X"40",X"A9",X"41",X"81",X"42",X"55",X"43",X"1A",X"44",X"DC",X"44",
		X"92",X"45",X"33",X"46",X"67",X"45",X"FE",X"42",X"A8",X"3F",X"A9",X"3B",X"4F",X"37",X"BB",X"32",
		X"13",X"2E",X"64",X"29",X"BE",X"24",X"2C",X"20",X"B2",X"1B",X"50",X"17",X"0F",X"13",X"EC",X"0E",
		X"EB",X"0A",X"08",X"07",X"43",X"03",X"A1",X"FF",X"18",X"FC",X"B2",X"F8",X"64",X"F5",X"38",X"F2",
		X"22",X"EF",X"2B",X"EC",X"47",X"E9",X"89",X"E6",X"CB",X"E3",X"B1",X"E1",X"72",X"E1",X"80",X"E2",
		X"6D",X"E4",X"E6",X"E6",X"BD",X"E9",X"C6",X"EC",X"ED",X"EF",X"1A",X"F3",X"49",X"F6",X"6C",X"F9",
		X"83",X"FC",X"86",X"FF",X"76",X"02",X"4F",X"05",X"14",X"08",X"C3",X"0A",X"5C",X"0D",X"DF",X"0F",
		X"4E",X"12",X"A7",X"14",X"ED",X"16",X"1E",X"19",X"3B",X"1B",X"45",X"1D",X"40",X"1F",X"27",X"21",
		X"FB",X"22",X"C2",X"24",X"76",X"26",X"1E",X"28",X"B3",X"29",X"3A",X"2B",X"B3",X"2C",X"20",X"2E",
		X"7F",X"2F",X"CF",X"30",X"13",X"32",X"4C",X"33",X"79",X"34",X"99",X"35",X"B0",X"36",X"B9",X"37",
		X"BA",X"38",X"B0",X"39",X"9D",X"3A",X"80",X"3B",X"59",X"3C",X"2B",X"3D",X"F2",X"3D",X"B2",X"3E",
		X"69",X"3F",X"19",X"40",X"C2",X"40",X"62",X"41",X"FA",X"41",X"8D",X"42",X"18",X"43",X"9E",X"43",
		X"1B",X"44",X"95",X"44",X"08",X"45",X"74",X"45",X"DC",X"45",X"3E",X"46",X"99",X"46",X"F0",X"46",
		X"43",X"47",X"91",X"47",X"D8",X"47",X"1F",X"48",X"5E",X"48",X"9C",X"48",X"D2",X"48",X"07",X"49",
		X"36",X"49",X"66",X"49",X"8C",X"49",X"B4",X"49",X"D3",X"49",X"F7",X"49",X"0A",X"4A",X"30",X"4A",
		X"47",X"49",X"A0",X"46",X"F8",X"42",X"93",X"3E",X"CD",X"39",X"C7",X"34",X"A9",X"2F",X"84",X"2A",
		X"6D",X"25",X"65",X"20",X"7B",X"1B",X"AD",X"16",X"01",X"12",X"78",X"0D",X"11",X"09",X"CF",X"04",
		X"AD",X"00",X"AE",X"FC",X"CF",X"F8",X"13",X"F5",X"75",X"F1",X"F7",X"ED",X"96",X"EA",X"54",X"E7",
		X"2C",X"E4",X"21",X"E1",X"32",X"DE",X"5A",X"DB",X"9E",X"D8",X"FA",X"D5",X"6C",X"D3",X"F6",X"D0",
		X"96",X"CE",X"4B",X"CC",X"18",X"CA",X"F6",X"C7",X"EA",X"C5",X"F0",X"C3",X"09",X"C2",X"33",X"C0",
		X"71",X"BE",X"BC",X"BC",X"19",X"BB",X"88",X"B9",X"02",X"B8",X"8F",X"B6",X"29",X"B5",X"D0",X"B3",
		X"87",X"B2",X"49",X"B1",X"18",X"B0",X"F4",X"AE",X"DD",X"AD",X"CF",X"AC",X"CE",X"AB",X"D8",X"AA",
		X"ED",X"A9",X"0A",X"A9",X"32",X"A8",X"67",X"A7",X"A2",X"A6",X"E5",X"A5",X"34",X"A5",X"88",X"A4",
		X"E6",X"A3",X"4C",X"A3",X"BB",X"A2",X"30",X"A2",X"AC",X"A1",X"30",X"A1",X"BB",X"A0",X"4B",X"A0",
		X"E3",X"9F",X"80",X"9F",X"23",X"9F",X"CD",X"9E",X"7A",X"9E",X"31",X"9E",X"EA",X"9D",X"A9",X"9D",
		X"6D",X"9D",X"34",X"9D",X"02",X"9D",X"D3",X"9C",X"A7",X"9C",X"84",X"9C",X"62",X"9C",X"43",X"9C",
		X"29",X"9C",X"15",X"9C",X"FF",X"9B",X"F1",X"9B",X"E5",X"9B",X"DE",X"9B",X"D7",X"9B",X"D5",X"9B",
		X"D4",X"9B",X"D6",X"9B",X"DD",X"9B",X"E5",X"9B",X"EF",X"9B",X"FE",X"9B",X"0E",X"9C",X"20",X"9C",
		X"35",X"9C",X"4B",X"9C",X"64",X"9C",X"7F",X"9C",X"9A",X"9C",X"BB",X"9C",X"D8",X"9C",X"FB",X"9C",
		X"20",X"9D",X"45",X"9D",X"6C",X"9D",X"94",X"9D",X"BE",X"9D",X"E9",X"9D",X"15",X"9E",X"43",X"9E",
		X"73",X"9E",X"A2",X"9E",X"D4",X"9E",X"07",X"9F",X"3A",X"9F",X"70",X"9F",X"A6",X"9F",X"DC",X"9F",
		X"16",X"A0",X"4C",X"A0",X"87",X"A0",X"BF",X"A0",X"FD",X"A0",X"36",X"A1",X"75",X"A1",X"B0",X"A1",
		X"F2",X"A1",X"32",X"A2",X"C9",X"A3",X"FE",X"A6",X"20",X"AB",X"E9",X"AF",X"0B",X"B5",X"63",X"BA",
		X"CB",X"BF",X"34",X"C5",X"8C",X"CA",X"D1",X"CF",X"F7",X"D4",X"FD",X"D9",X"E0",X"DE",X"9F",X"E3",
		X"3A",X"E8",X"B0",X"EC",X"01",X"F1",X"32",X"F5",X"3E",X"F9",X"28",X"FD",X"F3",X"00",X"9C",X"04",
		X"28",X"08",X"91",X"0B",X"E2",X"0E",X"10",X"12",X"33",X"15",X"C7",X"17",X"83",X"18",X"E5",X"17",
		X"5E",X"16",X"43",X"14",X"C8",X"11",X"13",X"0F",X"40",X"0C",X"5F",X"09",X"7C",X"06",X"A1",X"03",
		X"D1",X"00",X"12",X"FE",X"65",X"FB",X"C7",X"F8",X"40",X"F6",X"CC",X"F3",X"6B",X"F1",X"1F",X"EF",
		X"E8",X"EC",X"C2",X"EA",X"B1",X"E8",X"B0",X"E6",X"C3",X"E4",X"E3",X"E2",X"18",X"E1",X"5A",X"DF",
		X"AF",X"DD",X"11",X"DC",X"83",X"DA",X"02",X"D9",X"91",X"D7",X"2D",X"D6",X"D6",X"D4",X"8A",X"D3",
		X"4D",X"D2",X"1A",X"D1",X"F5",X"CF",X"D7",X"CE",X"C9",X"CD",X"C1",X"CC",X"C8",X"CB",X"D4",X"CA",
		X"EE",X"C9",X"0E",X"C9",X"39",X"C8",X"6A",X"C7",X"A9",X"C6",X"EA",X"C5",X"3A",X"C5",X"89",X"C4",
		X"E9",X"C3",X"45",X"C3",X"B9",X"C2",X"1A",X"C2",X"7B",X"C2",X"A4",X"C4",X"DA",X"C7",X"CD",X"CB",
		X"2B",X"D0",X"CF",X"D4",X"8D",X"D9",X"56",X"DE",X"15",X"E3",X"C7",X"E7",X"5F",X"EC",X"DA",X"F0",
		X"3A",X"F5",X"78",X"F9",X"98",X"FD",X"94",X"01",X"72",X"05",X"2E",X"09",X"CD",X"0C",X"4E",X"10",
		X"B0",X"13",X"F4",X"16",X"1E",X"1A",X"29",X"1D",X"1D",X"20",X"F5",X"22",X"B8",X"25",X"36",X"28",
		X"0C",X"29",X"52",X"28",X"AA",X"26",X"56",X"24",X"A1",X"21",X"A8",X"1E",X"92",X"1B",X"68",X"18",
		X"41",X"15",X"1C",X"12",X"09",X"0F",X"04",X"0C",X"13",X"09",X"35",X"06",X"70",X"03",X"BB",X"00",
		X"23",X"FE",X"99",X"FB",X"2A",X"F9",X"CA",X"F6",X"83",X"F4",X"4D",X"F2",X"2C",X"F0",X"1A",X"EE",
		X"21",X"EC",X"32",X"EA",X"5B",X"E8",X"8D",X"E6",X"D7",X"E4",X"29",X"E3",X"91",X"E1",X"FF",X"DF",
		X"87",X"DE",X"0F",X"DD",X"B5",X"DB",X"50",X"DA",X"31",X"D9",X"69",X"D8",X"30",X"D7",X"15",X"D6",
		X"FA",X"D4",X"F0",X"D3",X"EA",X"D2",X"F6",X"D1",X"06",X"D1",X"21",X"D0",X"43",X"CF",X"71",X"CE",
		X"A8",X"CD",X"E5",X"CC",X"29",X"CC",X"76",X"CB",X"CB",X"CA",X"28",X"CA",X"8A",X"C9",X"F6",X"C8",
		X"66",X"C8",X"DD",X"C7",X"5C",X"C7",X"DE",X"C6",X"67",X"C6",X"F7",X"C5",X"8A",X"C5",X"27",X"C5",
		X"C5",X"C4",X"6A",X"C4",X"11",X"C4",X"BF",X"C3",X"72",X"C3",X"28",X"C3",X"E2",X"C2",X"A3",X"C2",
		X"63",X"C2",X"2E",X"C2",X"F6",X"C1",X"C5",X"C1",X"95",X"C1",X"6D",X"C1",X"44",X"C1",X"22",X"C1",
		X"FE",X"C0",X"E2",X"C0",X"C4",X"C0",X"B0",X"C0",X"96",X"C0",X"88",X"C0",X"71",X"C0",X"6B",X"C0",
		X"56",X"C0",X"56",X"C0",X"43",X"C0",X"4E",X"C0",X"32",X"C0",X"7B",X"C0",X"4F",X"C1",X"43",X"C1",
		X"51",X"C1",X"51",X"C1",X"5F",X"C1",X"63",X"C1",X"73",X"C1",X"7D",X"C1",X"8C",X"C1",X"9B",X"C1",
		X"AC",X"C1",X"BD",X"C1",X"D2",X"C1",X"E6",X"C1",X"FC",X"C1",X"15",X"C2",X"2C",X"C2",X"47",X"C2",
		X"60",X"C2",X"7C",X"C2",X"97",X"C2",X"B5",X"C2",X"D3",X"C2",X"F4",X"C2",X"12",X"C3",X"32",X"C3",
		X"53",X"C3",X"75",X"C3",X"98",X"C3",X"BE",X"C3",X"E0",X"C3",X"06",X"C4",X"2A",X"C4",X"51",X"C4",
		X"75",X"C4",X"9E",X"C4",X"C5",X"C4",X"EE",X"C4",X"16",X"C5",X"40",X"C5",X"68",X"C5",X"93",X"C5",
		X"BD",X"C5",X"E8",X"C5",X"11",X"C6",X"3F",X"C6",X"69",X"C6",X"96",X"C6",X"C1",X"C6",X"F0",X"C6",
		X"1B",X"C7",X"49",X"C7",X"76",X"C7",X"A4",X"C7",X"D1",X"C7",X"FF",X"C7",X"2D",X"C8",X"5D",X"C8",
		X"8A",X"C8",X"BA",X"C8",X"E9",X"C8",X"18",X"C9",X"47",X"C9",X"78",X"C9",X"A6",X"C9",X"D7",X"C9",
		X"03",X"CA",X"35",X"CA",X"65",X"CA",X"95",X"CA",X"C5",X"CA",X"F6",X"CA",X"26",X"CB",X"57",X"CB",
		X"85",X"CB",X"B8",X"CB",X"E7",X"CB",X"18",X"CC",X"48",X"CC",X"77",X"CC",X"A8",X"CC",X"D8",X"CC",
		X"09",X"CD",X"3A",X"CD",X"6A",X"CD",X"9B",X"CD",X"CA",X"CD",X"FB",X"CD",X"2C",X"CE",X"5B",X"CE",
		X"8E",X"CE",X"BD",X"CE",X"EC",X"CE",X"1D",X"CF",X"4C",X"CF",X"7D",X"CF",X"AC",X"CF",X"DD",X"CF",
		X"0C",X"D0",X"3C",X"D0",X"6C",X"D0",X"9B",X"D0",X"CC",X"D0",X"FB",X"D0",X"2C",X"D1",X"5A",X"D1",
		X"8B",X"D1",X"BA",X"D1",X"E8",X"D1",X"15",X"D2",X"47",X"D2",X"75",X"D2",X"A5",X"D2",X"D3",X"D2",
		X"02",X"D3",X"2F",X"D3",X"60",X"D3",X"8D",X"D3",X"BC",X"D3",X"E7",X"D3",X"17",X"D4",X"43",X"D4",
		X"76",X"D4",X"9F",X"D4",X"D4",X"D4",X"F1",X"D4",X"E8",X"D5",X"96",X"D8",X"4C",X"DC",X"BB",X"E0",
		X"8B",X"E5",X"9D",X"EA",X"C5",X"EF",X"F6",X"F4",X"16",X"FA",X"25",X"FF",X"15",X"04",X"EA",X"08",
		X"9A",X"0D",X"2A",X"12",X"94",X"16",X"DA",X"1A",X"FE",X"1E",X"00",X"23",X"DD",X"26",X"9C",X"2A",
		X"36",X"2E",X"B5",X"31",X"12",X"35",X"53",X"38",X"77",X"3B",X"7E",X"3E",X"6B",X"41",X"3B",X"44",
		X"F3",X"46",X"90",X"49",X"18",X"4C",X"86",X"4E",X"DC",X"50",X"1F",X"53",X"4D",X"55",X"64",X"57",
		X"68",X"59",X"59",X"5B",X"34",X"5D",X"FE",X"5E",X"B9",X"60",X"5E",X"62",X"F6",X"63",X"7C",X"65",
		X"F5",X"66",X"5C",X"68",X"B6",X"69",X"FF",X"6A",X"3C",X"6C",X"6C",X"6D",X"8F",X"6E",X"A3",X"6F",
		X"AE",X"70",X"AC",X"71",X"9F",X"72",X"85",X"73",X"62",X"74",X"34",X"75",X"FB",X"75",X"B9",X"76",
		X"6E",X"77",X"18",X"78",X"BB",X"78",X"55",X"79",X"E8",X"79",X"71",X"7A",X"F4",X"7A",X"6C",X"7B",
		X"DE",X"7B",X"4A",X"7C",X"AE",X"7C",X"0C",X"7D",X"62",X"7D",X"B3",X"7D",X"FE",X"7D",X"44",X"7E",
		X"82",X"7E",X"BC",X"7E",X"F1",X"7E",X"21",X"7F",X"4A",X"7F",X"6F",X"7F",X"90",X"7F",X"AD",X"7F",
		X"C5",X"7F",X"D7",X"7F",X"E7",X"7F",X"F2",X"7F",X"F9",X"7F",X"FE",X"7F",X"FF",X"7F",X"FA",X"7F",
		X"F4",X"7F",X"EB",X"7F",X"DE",X"7F",X"CE",X"7F",X"BB",X"7F",X"A5",X"7F",X"8D",X"7F",X"72",X"7F",
		X"54",X"7F",X"34",X"7F",X"11",X"7F",X"EC",X"7E",X"C6",X"7E",X"9C",X"7E",X"71",X"7E",X"44",X"7E",
		X"14",X"7E",X"E3",X"7D",X"B0",X"7D",X"7B",X"7D",X"44",X"7D",X"0C",X"7D",X"D3",X"7C",X"98",X"7C",
		X"5B",X"7C",X"1E",X"7C",X"DF",X"7B",X"9E",X"7B",X"5E",X"7B",X"1C",X"7B",X"D7",X"7A",X"93",X"7A",
		X"4E",X"7A",X"04",X"7A",X"BD",X"79",X"73",X"79",X"29",X"79",X"DD",X"78",X"92",X"78",X"47",X"78",
		X"FA",X"77",X"AB",X"77",X"5D",X"77",X"0E",X"77",X"BE",X"76",X"6E",X"76",X"1C",X"76",X"CC",X"75",
		X"79",X"75",X"25",X"75",X"D3",X"74",X"80",X"74",X"2E",X"74",X"D8",X"73",X"82",X"73",X"2E",X"73",
		X"DA",X"72",X"82",X"72",X"2C",X"72",X"D4",X"71",X"80",X"71",X"27",X"71",X"D3",X"70",X"79",X"70",
		X"23",X"70",X"CB",X"6F",X"74",X"6F",X"1B",X"6F",X"C3",X"6E",X"69",X"6E",X"13",X"6E",X"B6",X"6D",
		X"65",X"6D",X"C9",X"6C",X"89",X"6A",X"FA",X"66",X"9B",X"62",X"BC",X"5D",X"92",X"58",X"42",X"53",
		X"E9",X"4D",X"93",X"48",X"51",X"43",X"26",X"3E",X"1B",X"39",X"2E",X"34",X"68",X"2F",X"C2",X"2A",
		X"40",X"26",X"E2",X"21",X"A8",X"1D",X"8F",X"19",X"97",X"15",X"C0",X"11",X"0C",X"0E",X"74",X"0A",
		X"FC",X"06",X"9F",X"03",X"63",X"00",X"3F",X"FD",X"37",X"FA",X"47",X"F7",X"73",X"F4",X"B6",X"F1",
		X"12",X"EF",X"83",X"EC",X"0C",X"EA",X"A9",X"E7",X"5F",X"E5",X"26",X"E3",X"02",X"E1",X"EF",X"DE",
		X"F3",X"DC",X"04",X"DB",X"2B",X"D9",X"5F",X"D7",X"A7",X"D5",X"FC",X"D3",X"63",X"D2",X"D6",X"D0",
		X"5B",X"CF",X"EA",X"CD",X"8C",X"CC",X"34",X"CB",X"F1",X"C9",X"B1",X"C8",X"8B",X"C7",X"59",X"C6",
		X"FB",X"C5",X"5F",X"C7",X"DD",X"C9",X"21",X"CD",X"D7",X"D0",X"D6",X"D4",X"F7",X"D8",X"27",X"DD",
		X"54",X"E1",X"78",X"E5",X"86",X"E9",X"81",X"ED",X"5F",X"F1",X"22",X"F5",X"CA",X"F8",X"55",X"FC",
		X"C4",X"FF",X"17",X"03",X"4C",X"06",X"69",X"09",X"6A",X"0C",X"53",X"0F",X"21",X"12",X"D9",X"14",
		X"74",X"17",X"FF",X"19",X"70",X"1C",X"B9",X"1E",X"81",X"1F",X"B7",X"1E",X"FF",X"1C",X"98",X"1A",
		X"CF",X"17",X"C3",X"14",X"9C",X"11",X"5F",X"0E",X"27",X"0B",X"F2",X"07",X"D0",X"04",X"BA",X"01",
		X"BD",X"FE",X"D1",X"FB",X"FD",X"F8",X"3E",X"F6",X"96",X"F3",X"02",X"F1",X"87",X"EE",X"21",X"EC",
		X"CF",X"E9",X"8E",X"E7",X"64",X"E5",X"4C",X"E3",X"48",X"E1",X"55",X"DF",X"73",X"DD",X"A4",X"DB",
		X"E4",X"D9",X"35",X"D8",X"95",X"D6",X"04",X"D5",X"82",X"D3",X"0E",X"D2",X"A7",X"D0",X"4E",X"CF",
		X"02",X"CE",X"C2",X"CC",X"8F",X"CB",X"66",X"CA",X"4B",X"C9",X"39",X"C8",X"31",X"C7",X"35",X"C6",
		X"44",X"C5",X"5C",X"C4",X"7D",X"C3",X"A7",X"C2",X"DA",X"C1",X"16",X"C1",X"59",X"C0",X"A7",X"BF",
		X"F8",X"BE",X"57",X"BE",X"BE",X"BD",X"69",X"BE",X"B5",X"C0",X"EE",X"C3",X"CF",X"C7",X"0C",X"CC",
		X"87",X"D0",X"15",X"D5",X"AC",X"D9",X"36",X"DE",X"B5",X"E2",X"17",X"E7",X"63",X"EB",X"8D",X"EF",
		X"9C",X"F3",X"8A",X"F7",X"5B",X"FB",X"0C",X"FF",X"9D",X"02",X"12",X"06",X"6B",X"09",X"A4",X"0C",
		X"C5",X"0F",X"C9",X"12",X"B5",X"15",X"85",X"18",X"3D",X"1B",X"DD",X"1D",X"67",X"20",X"D9",X"22",
		X"36",X"25",X"7D",X"27",X"B1",X"29",X"D1",X"2B",X"DD",X"2D",X"D6",X"2F",X"BC",X"31",X"93",X"33",
		X"58",X"35",X"0D",X"37",X"AF",X"38",X"44",X"3A",X"C7",X"3B",X"40",X"3D",X"A7",X"3E",X"04",X"40",
		X"50",X"41",X"91",X"42",X"C5",X"43",X"EE",X"44",X"07",X"46",X"1A",X"47",X"1A",X"48",X"1B",X"49",
		X"04",X"4A",X"F5",X"4A",X"C7",X"4A",X"E9",X"48",X"0A",X"46",X"77",X"42",X"7F",X"3E",X"44",X"3A",
		X"EF",X"35",X"8E",X"31",X"33",X"2D",X"E7",X"28",X"AF",X"24",X"91",X"20",X"8D",X"1C",X"A7",X"18",
		X"DC",X"14",X"30",X"11",X"A0",X"0D",X"30",X"0A",X"D9",X"06",X"9E",X"03",X"80",X"00",X"7E",X"FD",
		X"91",X"FA",X"BF",X"F7",X"04",X"F5",X"65",X"F2",X"D2",X"EF",X"99",X"ED",X"0E",X"ED",X"EF",X"ED",
		X"B6",X"EF",X"18",X"F2",X"D5",X"F4",X"CF",X"F7",X"E4",X"FA",X"06",X"FE",X"26",X"01",X"41",X"04",
		X"4A",X"07",X"46",X"0A",X"2B",X"0D",X"FD",X"0F",X"B8",X"12",X"5E",X"15",X"ED",X"17",X"6A",X"1A",
		X"CD",X"1C",X"20",X"1F",X"5B",X"21",X"83",X"23",X"98",X"25",X"9B",X"27",X"8A",X"29",X"6A",X"2B",
		X"36",X"2D",X"F4",X"2E",X"A0",X"30",X"3E",X"32",X"CB",X"33",X"4B",X"35",X"BA",X"36",X"1E",X"38",
		X"74",X"39",X"BC",X"3A",X"F9",X"3B",X"28",X"3D",X"4B",X"3E",X"65",X"3F",X"72",X"40",X"75",X"41",
		X"6D",X"42",X"5A",X"43",X"3F",X"44",X"1A",X"45",X"EB",X"45",X"B4",X"46",X"73",X"47",X"2A",X"48",
		X"D8",X"48",X"81",X"49",X"20",X"4A",X"BB",X"4A",X"2E",X"4B",X"1B",X"4A",X"93",X"47",X"29",X"44",
		X"28",X"40",X"D3",X"3B",X"4A",X"37",X"AF",X"32",X"0E",X"2E",X"7C",X"29",X"FC",X"24",X"92",X"20",
		X"45",X"1C",X"16",X"18",X"06",X"14",X"11",X"10",X"40",X"0C",X"8C",X"08",X"F7",X"04",X"7F",X"01",
		X"26",X"FE",X"E6",X"FA",X"C7",X"F7",X"BC",X"F4",X"D1",X"F1",X"F9",X"EE",X"45",X"EC",X"92",X"E9",
		X"A5",X"E7",X"87",X"E7",X"9A",X"E8",X"81",X"EA",X"E6",X"EC",X"A4",X"EF",X"8D",X"F2",X"92",X"F5",
		X"9E",X"F8",X"AA",X"FB",X"A9",X"FE",X"9B",X"01",X"7D",X"04",X"4A",X"07",X"05",X"0A",X"A9",X"0C",
		X"36",X"0F",X"B1",X"11",X"16",X"14",X"69",X"16",X"A4",X"18",X"D0",X"1A",X"E5",X"1C",X"EA",X"1E",
		X"D9",X"20",X"BD",X"22",X"87",X"24",X"3D",X"26",X"8B",X"26",X"40",X"25",X"03",X"23",X"1A",X"20",
		X"D0",X"1C",X"46",X"19",X"A0",X"15",X"EC",X"11",X"3D",X"0E",X"95",X"0A",X"02",X"07",X"81",X"03",
		X"18",X"00",X"C9",X"FC",X"92",X"F9",X"75",X"F6",X"70",X"F3",X"85",X"F0",X"B3",X"ED",X"F8",X"EA",
		X"54",X"E8",X"CA",X"E5",X"51",X"E3",X"F4",X"E0",X"A6",X"DE",X"75",X"DC",X"45",X"DA",X"A9",X"D8",
		X"D3",X"D8",X"41",X"DA",X"85",X"DC",X"50",X"DF",X"72",X"E2",X"C4",X"E5",X"2F",X"E9",X"9E",X"EC",
		X"0B",X"F0",X"6C",X"F3",X"BD",X"F6",X"F7",X"F9",X"1F",X"FD",X"2D",X"00",X"24",X"03",X"04",X"06",
		X"CD",X"08",X"7F",X"0B",X"1A",X"0E",X"A1",X"10",X"0E",X"13",X"69",X"15",X"AE",X"17",X"E0",X"19",
		X"FD",X"1B",X"09",X"1E",X"02",X"20",X"EA",X"21",X"BF",X"23",X"85",X"25",X"3B",X"27",X"E0",X"28",
		X"75",X"2A",X"FE",X"2B",X"75",X"2D",X"E2",X"2E",X"3F",X"30",X"90",X"31",X"D4",X"32",X"0D",X"34",
		X"37",X"35",X"5A",X"36",X"6D",X"37",X"79",X"38",X"77",X"39",X"6E",X"3A",X"5A",X"3B",X"3D",X"3C",
		X"15",X"3D",X"E6",X"3D",X"AC",X"3E",X"6D",X"3F",X"1F",X"40",X"D8",X"40",X"32",X"41",X"E3",X"3F",
		X"41",X"3D",X"CB",X"39",X"CC",X"35",X"7E",X"31",X"05",X"2D",X"7C",X"28",X"F0",X"23",X"73",X"1F",
		X"0A",X"1B",X"B8",X"16",X"82",X"12",X"69",X"0E",X"72",X"0A",X"96",X"06",X"DA",X"02",X"3C",X"FF",
		X"BD",X"FB",X"5B",X"F8",X"16",X"F5",X"E8",X"F1",X"DD",X"EE",X"E5",X"EB",X"0D",X"E9",X"48",X"E6",
		X"A7",X"E3",X"07",X"E1",X"7A",X"DF",X"B2",X"DF",X"FC",X"E0",X"0F",X"E3",X"93",X"E5",X"6A",X"E8",
		X"64",X"EB",X"7A",X"EE",X"90",X"F1",X"A5",X"F4",X"AD",X"F7",X"A8",X"FA",X"8F",X"FD",X"66",X"00",
		X"23",X"03",X"D0",X"05",X"64",X"08",X"E3",X"0A",X"4E",X"0D",X"A6",X"0F",X"E8",X"11",X"16",X"14",
		X"33",X"16",X"3D",X"18",X"35",X"1A",X"1A",X"1C",X"EE",X"1D",X"B4",X"1F",X"68",X"21",X"0D",X"23",
		X"A2",X"24",X"29",X"26",X"A3",X"27",X"0E",X"29",X"6D",X"2A",X"BE",X"2B",X"03",X"2D",X"3B",X"2E",
		X"68",X"2F",X"89",X"30",X"A0",X"31",X"AA",X"32",X"AD",X"33",X"A2",X"34",X"92",X"35",X"73",X"36",
		X"50",X"37",X"20",X"38",X"EC",X"38",X"AA",X"39",X"66",X"3A",X"12",X"3B",X"C2",X"3B",X"5B",X"3C",
		X"05",X"3D",X"E0",X"3C",X"FF",X"3A",X"02",X"38",X"49",X"34",X"20",X"30",X"B3",X"2B",X"26",X"27",
		X"8D",X"22",X"FB",X"1D",X"77",X"19",X"08",X"15",X"B6",X"10",X"7E",X"0C",X"65",X"08",X"6D",X"04",
		X"94",X"00",X"D7",X"FC",X"3B",X"F9",X"BD",X"F5",X"5D",X"F2",X"17",X"EF",X"F1",X"EB",X"E1",X"E8",
		X"F3",X"E5",X"15",X"E3",X"5F",X"E0",X"A7",X"DD",X"A9",X"DB",X"79",X"DB",X"80",X"DC",X"5F",X"DE",
		X"C0",X"E0",X"7A",X"E3",X"64",X"E6",X"69",X"E9",X"75",X"EC",X"80",X"EF",X"84",X"F2",X"78",X"F5",
		X"5B",X"F8",X"2D",X"FB",X"E9",X"FD",X"8F",X"00",X"22",X"03",X"A1",X"05",X"09",X"08",X"5E",X"0A",
		X"9F",X"0C",X"CC",X"0E",X"E7",X"10",X"EF",X"12",X"E6",X"14",X"CC",X"16",X"A1",X"18",X"65",X"1A",
		X"19",X"1C",X"BE",X"1D",X"54",X"1F",X"DC",X"20",X"55",X"22",X"BF",X"23",X"1F",X"25",X"70",X"26",
		X"B7",X"27",X"EF",X"28",X"1F",X"2A",X"3F",X"2B",X"58",X"2C",X"65",X"2D",X"69",X"2E",X"5F",X"2F",
		X"50",X"30",X"33",X"31",X"12",X"32",X"E4",X"32",X"B0",X"33",X"71",X"34",X"2E",X"35",X"DE",X"35",
		X"8F",X"36",X"2A",X"37",X"D6",X"37",X"05",X"38",X"81",X"36",X"BC",X"33",X"28",X"30",X"14",X"2C",
		X"B4",X"27",X"2D",X"23",X"95",X"1E",X"03",X"1A",X"7D",X"15",X"0D",X"11",X"B2",X"0C",X"77",X"08",
		X"59",X"04",X"5B",X"00",X"7B",X"FC",X"BA",X"F8",X"19",X"F5",X"98",X"F1",X"31",X"EE",X"E9",X"EA",
		X"BC",X"E7",X"AE",X"E4",X"B6",X"E1",X"DD",X"DE",X"17",X"DC",X"73",X"D9",X"D8",X"D6",X"6F",X"D5",
		X"C7",X"D5",X"22",X"D7",X"3F",X"D9",X"CA",X"DB",X"A5",X"DE",X"A1",X"E1",X"B6",X"E4",X"CF",X"E7",
		X"E3",X"EA",X"EC",X"ED",X"E7",X"F0",X"CE",X"F3",X"A2",X"F6",X"62",X"F9",X"0E",X"FC",X"A2",X"FE",
		X"21",X"01",X"8E",X"03",X"E5",X"05",X"29",X"08",X"59",X"0A",X"78",X"0C",X"81",X"0E",X"7D",X"10",
		X"62",X"12",X"42",X"14",X"C6",X"15",X"9F",X"15",X"15",X"14",X"AE",X"11",X"B1",X"0E",X"5F",X"0B",
		X"D7",X"07",X"37",X"04",X"8F",X"00",X"F0",X"FC",X"5A",X"F9",X"D8",X"F5",X"69",X"F2",X"14",X"EF",
		X"D6",X"EB",X"B3",X"E8",X"A8",X"E5",X"B8",X"E2",X"DE",X"DF",X"1F",X"DD",X"77",X"DA",X"E8",X"D7",
		X"6D",X"D5",X"0B",X"D3",X"BC",X"D0",X"84",X"CE",X"5E",X"CC",X"4D",X"CA",X"4D",X"C8",X"65",X"C6",
		X"8A",X"C4",X"C3",X"C2",X"0B",X"C1",X"65",X"BF",X"CD",X"BD",X"44",X"BC",X"CC",X"BA",X"61",X"B9",
		X"07",X"B8",X"B6",X"B6",X"77",X"B5",X"42",X"B4",X"18",X"B3",X"FC",X"B1",X"EC",X"B0",X"E7",X"AF",
		X"EB",X"AE",X"FD",X"AD",X"17",X"AD",X"3B",X"AC",X"69",X"AB",X"A0",X"AA",X"E0",X"A9",X"2B",X"A9",
		X"79",X"A8",X"F8",X"A7",X"FD",X"A8",X"7A",X"AB",X"D4",X"AE",X"C6",X"B2",X"0D",X"B7",X"88",X"BB",
		X"16",X"C0",X"A7",X"C4",X"2D",X"C9",X"A2",X"CD",X"FF",X"D1",X"3F",X"D6",X"65",X"DA",X"6D",X"DE",
		X"52",X"E2",X"1D",X"E6",X"CA",X"E9",X"58",X"ED",X"C9",X"F0",X"1C",X"F4",X"56",X"F7",X"71",X"FA",
		X"77",X"FD",X"5C",X"00",X"31",X"03",X"E3",X"05",X"94",X"08",X"77",X"0A",X"88",X"0A",X"70",X"09",
		X"84",X"07",X"1D",X"05",X"5F",X"02",X"76",X"FF",X"71",X"FC",X"67",X"F9",X"5D",X"F6",X"5E",X"F3",
		X"6E",X"F0",X"90",X"ED",X"C5",X"EA",X"0F",X"E8",X"6F",X"E5",X"E5",X"E2",X"6E",X"E0",X"0D",X"DE",
		X"C0",X"DB",X"8A",X"D9",X"65",X"D7",X"55",X"D5",X"55",X"D3",X"6B",X"D1",X"8E",X"CF",X"C5",X"CD",
		X"0B",X"CC",X"63",X"CA",X"CB",X"C8",X"41",X"C7",X"C7",X"C5",X"58",X"C4",X"FB",X"C2",X"A9",X"C1",
		X"63",X"C0",X"2C",X"BF",X"00",X"BE",X"E1",X"BC",X"CC",X"BB",X"C3",X"BA",X"C5",X"B9",X"D1",X"B8",
		X"E6",X"B7",X"06",X"B7",X"30",X"B6",X"64",X"B5",X"9F",X"B4",X"E2",X"B3",X"2F",X"B3",X"84",X"B2",
		X"E2",X"B1",X"46",X"B1",X"B1",X"B0",X"25",X"B0",X"9E",X"AF",X"1F",X"AF",X"A5",X"AE",X"33",X"AE",
		X"C7",X"AD",X"61",X"AD",X"01",X"AD",X"A5",X"AC",X"50",X"AC",X"FF",X"AB",X"B4",X"AB",X"6C",X"AB",
		X"2C",X"AB",X"EF",X"AA",X"B6",X"AA",X"7F",X"AA",X"50",X"AA",X"24",X"AA",X"FD",X"A9",X"D6",X"A9",
		X"B7",X"A9",X"97",X"A9",X"81",X"A9",X"67",X"A9",X"56",X"A9",X"43",X"A9",X"3B",X"A9",X"2E",X"A9",
		X"58",X"AA",X"1F",X"AD",X"D5",X"B0",X"35",X"B5",X"EE",X"B9",X"E2",X"BE",X"E6",X"C3",X"F1",X"C8",
		X"ED",X"CD",X"D7",X"D2",X"A5",X"D7",X"58",X"DC",X"E8",X"E0",X"59",X"E5",X"A5",X"E9",X"D2",X"ED",
		X"DC",X"F1",X"C9",X"F5",X"90",X"F9",X"3B",X"FD",X"C3",X"00",X"2F",X"04",X"7F",X"07",X"B4",X"0A",
		X"CB",X"0D",X"C9",X"10",X"AB",X"13",X"77",X"16",X"27",X"19",X"C2",X"1B",X"45",X"1E",X"B2",X"20",
		X"0A",X"23",X"4B",X"25",X"79",X"27",X"94",X"29",X"9B",X"2B",X"8D",X"2D",X"72",X"2F",X"42",X"31",
		X"05",X"33",X"B3",X"34",X"54",X"36",X"E4",X"37",X"67",X"39",X"DA",X"3A",X"41",X"3C",X"96",X"3D",
		X"E3",X"3E",X"1E",X"40",X"54",X"41",X"75",X"42",X"95",X"43",X"9B",X"44",X"AB",X"45",X"AC",X"45",
		X"F6",X"43",X"3C",X"41",X"C7",X"3D",X"EC",X"39",X"CC",X"35",X"90",X"31",X"46",X"2D",X"02",X"29",
		X"CA",X"24",X"A8",X"20",X"9B",X"1C",X"A9",X"18",X"D5",X"14",X"1D",X"11",X"82",X"0D",X"06",X"0A",
		X"A1",X"06",X"5C",X"03",X"32",X"00",X"22",X"FD",X"2C",X"FA",X"4F",X"F7",X"8B",X"F4",X"E0",X"F1",
		X"4B",X"EF",X"C7",X"EC",X"90",X"EA",X"FD",X"E9",X"E1",X"EA",X"AC",X"EC",X"14",X"EF",X"DB",X"F1",
		X"DC",X"F4",X"FD",X"F7",X"29",X"FB",X"55",X"FE",X"78",X"01",X"8E",X"04",X"92",X"07",X"83",X"0A",
		X"5D",X"0D",X"23",X"10",X"D3",X"12",X"6D",X"15",X"EE",X"17",X"5E",X"1A",X"B5",X"1C",X"FD",X"1E",
		X"2B",X"21",X"49",X"23",X"51",X"25",X"4D",X"27",X"2C",X"29",X"11",X"2B",X"11",X"2C",X"4C",X"2B",
		X"6B",X"29",X"C0",X"26",X"A4",X"23",X"36",X"20",X"A4",X"1C",X"FD",X"18",X"57",X"15",X"B5",X"11",
		X"24",X"0E",X"A5",X"0A",X"3E",X"07",X"EC",X"03",X"B6",X"00",X"98",X"FD",X"93",X"FA",X"A4",X"F7",
		X"CF",X"F4",X"14",X"F2",X"6C",X"EF",X"DE",X"EC",X"66",X"EA",X"04",X"E8",X"B6",X"E5",X"7C",X"E3",
		X"56",X"E1",X"5B",X"DF",X"E2",X"DE",X"F7",X"DF",X"F9",X"E1",X"A1",X"E4",X"A7",X"E7",X"F2",X"EA",
		X"55",X"EE",X"C7",X"F1",X"36",X"F5",X"9F",X"F8",X"F5",X"FB",X"3A",X"FF",X"66",X"02",X"81",X"05",
		X"81",X"08",X"69",X"0B",X"3B",X"0E",X"F5",X"10",X"98",X"13",X"24",X"16",X"9A",X"18",X"FB",X"1A",
		X"47",X"1D",X"7D",X"1F",X"A3",X"21",X"B2",X"23",X"A8",X"25",X"3C",X"26",X"2F",X"25",X"33",X"23",
		X"7F",X"20",X"6E",X"1D",X"17",X"1A",X"A4",X"16",X"1F",X"13",X"9F",X"0F",X"24",X"0C",X"BC",X"08",
		X"63",X"05",X"26",X"02",X"FA",X"FE",X"EB",X"FB",X"EF",X"F8",X"0F",X"F6",X"44",X"F3",X"93",X"F0",
		X"F7",X"ED",X"73",X"EB",X"03",X"E9",X"AA",X"E6",X"65",X"E4",X"35",X"E2",X"16",X"E0",X"0C",X"DE",
		X"14",X"DC",X"2C",X"DA",X"58",X"D8",X"93",X"D6",X"E1",X"D4",X"3B",X"D3",X"A7",X"D1",X"22",X"D0",
		X"AA",X"CE",X"40",X"CD",X"E4",X"CB",X"94",X"CA",X"52",X"C9",X"1B",X"C8",X"F2",X"C6",X"D3",X"C5",
		X"C0",X"C4",X"B6",X"C3",X"B9",X"C2",X"C4",X"C1",X"DD",X"C0",X"FA",X"BF",X"26",X"BF",X"55",X"BE",
		X"93",X"BD",X"D1",X"BC",X"24",X"BC",X"72",X"BB",X"E9",X"BB",X"0E",X"BE",X"27",X"C1",X"F3",X"C4",
		X"1D",X"C9",X"87",X"CD",X"0A",X"D2",X"96",X"D6",X"17",X"DB",X"8D",X"DF",X"E7",X"E3",X"2C",X"E8",
		X"50",X"EC",X"5B",X"F0",X"43",X"F4",X"0C",X"F8",X"B8",X"FB",X"46",X"FF",X"B5",X"02",X"0A",X"06",
		X"3F",X"09",X"5C",X"0C",X"5D",X"0F",X"44",X"12",X"11",X"15",X"C7",X"17",X"65",X"1A",X"ED",X"1C",
		X"5D",X"1F",X"B8",X"21",X"FE",X"23",X"2F",X"26",X"4B",X"28",X"56",X"2A",X"4E",X"2C",X"34",X"2E",
		X"09",X"30",X"CB",X"31",X"7F",X"33",X"21",X"35",X"B5",X"36",X"3B",X"38",X"B0",X"39",X"19",X"3B",
		X"73",X"3C",X"BE",X"3D",X"00",X"3F",X"34",X"40",X"5B",X"41",X"78",X"42",X"89",X"43",X"8E",X"44",
		X"8A",X"45",X"7B",X"46",X"60",X"47",X"3F",X"48",X"13",X"49",X"DE",X"49",X"9F",X"4A",X"59",X"4B",
		X"0A",X"4C",X"B1",X"4C",X"53",X"4D",X"EF",X"4D",X"81",X"4E",X"0B",X"4F",X"90",X"4F",X"0E",X"50",
		X"86",X"50",X"F7",X"50",X"61",X"51",X"C7",X"51",X"26",X"52",X"81",X"52",X"D6",X"52",X"23",X"53",
		X"6F",X"53",X"B6",X"53",X"F7",X"53",X"34",X"54",X"6C",X"54",X"A0",X"54",X"CF",X"54",X"FB",X"54",
		X"23",X"55",X"47",X"55",X"67",X"55",X"86",X"55",X"A0",X"55",X"B6",X"55",X"C8",X"55",X"D9",X"55",
		X"E8",X"55",X"F1",X"55",X"F8",X"55",X"FF",X"55",X"01",X"56",X"01",X"56",X"FE",X"55",X"F9",X"55",
		X"F2",X"55",X"E9",X"55",X"DE",X"55",X"D0",X"55",X"C0",X"55",X"B0",X"55",X"9B",X"55",X"88",X"55",
		X"70",X"55",X"59",X"55",X"3E",X"55",X"21",X"55",X"05",X"55",X"E6",X"54",X"C8",X"54",X"A6",X"54",
		X"84",X"54",X"60",X"54",X"3A",X"54",X"14",X"54",X"EC",X"53",X"C4",X"53",X"9A",X"53",X"70",X"53",
		X"45",X"53",X"19",X"53",X"EC",X"52",X"BC",X"52",X"8E",X"52",X"5E",X"52",X"2E",X"52",X"FE",X"51",
		X"CB",X"51",X"98",X"51",X"66",X"51",X"30",X"51",X"FC",X"50",X"C7",X"50",X"92",X"50",X"5C",X"50",
		X"24",X"50",X"ED",X"4F",X"B7",X"4F",X"7E",X"4F",X"47",X"4F",X"0D",X"4F",X"D4",X"4E",X"9B",X"4E",
		X"62",X"4E",X"27",X"4E",X"ED",X"4D",X"B0",X"4D",X"76",X"4D",X"39",X"4D",X"FE",X"4C",X"C2",X"4C",
		X"87",X"4C",X"48",X"4C",X"0F",X"4C",X"D0",X"4B",X"96",X"4B",X"56",X"4B",X"1C",X"4B",X"D7",X"4A",
		X"AA",X"4A",X"E9",X"49",X"73",X"47",X"D5",X"43",X"72",X"3F",X"9C",X"3A",X"82",X"35",X"4B",X"30",
		X"0A",X"2B",X"D4",X"25",X"B0",X"20",X"A6",X"1B",X"BA",X"16",X"F3",X"11",X"4A",X"0D",X"C6",X"08",
		X"66",X"04",X"28",X"00",X"0E",X"FC",X"17",X"F8",X"42",X"F4",X"8B",X"F0",X"F5",X"EC",X"7E",X"E9",
		X"24",X"E6",X"E8",X"E2",X"C8",X"DF",X"C4",X"DC",X"DB",X"D9",X"0B",X"D7",X"55",X"D4",X"B7",X"D1",
		X"30",X"CF",X"BF",X"CC",X"65",X"CA",X"21",X"C8",X"F1",X"C5",X"D6",X"C3",X"CE",X"C1",X"DB",X"BF",
		X"F8",X"BD",X"27",X"BC",X"68",X"BA",X"BB",X"B8",X"1D",X"B7",X"8F",X"B5",X"10",X"B4",X"A0",X"B2",
		X"3F",X"B1",X"EB",X"AF",X"A5",X"AE",X"6D",X"AD",X"3F",X"AC",X"1E",X"AB",X"0B",X"AA",X"02",X"A9",
		X"06",X"A8",X"12",X"A7",X"2B",X"A6",X"4C",X"A5",X"79",X"A4",X"AE",X"A3",X"EE",X"A2",X"36",X"A2",
		X"85",X"A1",X"DF",X"A0",X"41",X"A0",X"AA",X"9F",X"1C",X"9F",X"92",X"9E",X"13",X"9E",X"98",X"9D",
		X"27",X"9D",X"B9",X"9C",X"56",X"9C",X"F4",X"9B",X"9C",X"9B",X"46",X"9B",X"FB",X"9A",X"B0",X"9A",
		X"6E",X"9A",X"2B",X"9A",X"F9",X"99",X"B9",X"99",X"8B",X"9A",X"0C",X"9D",X"87",X"A0",X"B6",X"A4",
		X"45",X"A9",X"15",X"AE",X"F9",X"B2",X"E8",X"B7",X"C9",X"BC",X"9B",X"C1",X"52",X"C6",X"EF",X"CA",
		X"6C",X"CF",X"CB",X"D3",X"06",X"D8",X"23",X"DC",X"1E",X"E0",X"FB",X"E3",X"B6",X"E7",X"55",X"EB",
		X"D3",X"EE",X"35",X"F2",X"7A",X"F5",X"A5",X"F8",X"B4",X"FB",X"AC",X"FE",X"87",X"01",X"4A",X"04",
		X"F7",X"06",X"8B",X"09",X"0B",X"0C",X"75",X"0E",X"C8",X"10",X"08",X"13",X"33",X"15",X"4C",X"17",
		X"53",X"19",X"46",X"1B",X"29",X"1D",X"FB",X"1E",X"BC",X"20",X"6E",X"22",X"10",X"24",X"A4",X"25",
		X"27",X"27",X"9E",X"28",X"07",X"2A",X"62",X"2B",X"B0",X"2C",X"F2",X"2D",X"28",X"2F",X"55",X"30",
		X"71",X"31",X"86",X"32",X"8F",X"33",X"90",X"34",X"84",X"35",X"6E",X"36",X"52",X"37",X"2B",X"38",
		X"FA",X"38",X"C0",X"39",X"81",X"3A",X"38",X"3B",X"E7",X"3B",X"8F",X"3C",X"2F",X"3D",X"C7",X"3D",
		X"5A",X"3E",X"E6",X"3E",X"6B",X"3F",X"EA",X"3F",X"62",X"40",X"D6",X"40",X"44",X"41",X"AC",X"41",
		X"0E",X"42",X"6A",X"42",X"C3",X"42",X"16",X"43",X"65",X"43",X"AF",X"43",X"DA",X"43",X"89",X"42",
		X"BF",X"3F",X"15",X"3C",X"D4",X"37",X"42",X"33",X"7D",X"2E",X"A9",X"29",X"D0",X"24",X"07",X"20",
		X"51",X"1B",X"B6",X"16",X"39",X"12",X"DA",X"0D",X"9C",X"09",X"7D",X"05",X"83",X"01",X"A8",X"FD",
		X"EB",X"F9",X"4E",X"F6",X"D1",X"F2",X"70",X"EF",X"2F",X"EC",X"04",X"E9",X"FB",X"E5",X"06",X"E3",
		X"38",X"E0",X"69",X"DD",X"5C",X"DB",X"21",X"DB",X"18",X"DC",X"E6",X"DD",X"36",X"E0",X"DF",X"E2",
		X"B6",X"E5",X"AA",X"E8",X"A4",X"EB",X"A0",X"EE",X"92",X"F1",X"77",X"F4",X"4C",X"F7",X"0D",X"FA",
		X"BB",X"FC",X"55",X"FF",X"D9",X"01",X"4A",X"04",X"A5",X"06",X"F0",X"08",X"25",X"0B",X"49",X"0D",
		X"58",X"0F",X"56",X"11",X"43",X"13",X"1F",X"15",X"EA",X"16",X"A6",X"18",X"51",X"1A",X"EE",X"1B",
		X"7C",X"1D",X"FB",X"1E",X"70",X"20",X"D3",X"21",X"2B",X"23",X"77",X"24",X"B5",X"25",X"E8",X"26",
		X"12",X"28",X"2D",X"29",X"42",X"2A",X"48",X"2B",X"48",X"2C",X"3B",X"2D",X"26",X"2E",X"06",X"2F",
		X"E3",X"2F",X"AE",X"30",X"79",X"31",X"36",X"32",X"F0",X"32",X"9C",X"33",X"4A",X"34",X"E5",X"34",
		X"83",X"35",X"EF",X"34",X"B6",X"32",X"89",X"2F",X"AD",X"2B",X"72",X"27",X"FB",X"22",X"6D",X"1E",
		X"D5",X"19",X"4A",X"15",X"CC",X"10",X"69",X"0C",X"1F",X"08",X"F4",X"03",X"E4",X"FF",X"F8",X"FB",
		X"28",X"F8",X"78",X"F4",X"E8",X"F0",X"75",X"ED",X"1C",X"EA",X"E6",X"E6",X"C7",X"E3",X"C6",X"E0",
		X"DF",X"DD",X"10",X"DB",X"5B",X"D8",X"BF",X"D5",X"38",X"D3",X"C9",X"D0",X"71",X"CE",X"2B",X"CC",
		X"FF",X"C9",X"E4",X"C7",X"DD",X"C5",X"E8",X"C3",X"06",X"C2",X"36",X"C0",X"76",X"BE",X"C8",X"BC",
		X"2B",X"BB",X"9C",X"B9",X"1D",X"B8",X"AD",X"B6",X"4A",X"B5",X"F6",X"B3",X"AF",X"B2",X"77",X"B1",
		X"48",X"B0",X"28",X"AF",X"11",X"AE",X"09",X"AD",X"0A",X"AC",X"17",X"AB",X"2E",X"AA",X"4D",X"A9",
		X"79",X"A8",X"AE",X"A7",X"EC",X"A6",X"31",X"A6",X"81",X"A5",X"D8",X"A4",X"37",X"A4",X"A1",X"A3",
		X"0F",X"A3",X"86",X"A2",X"03",X"A2",X"88",X"A1",X"12",X"A1",X"A6",X"A0",X"3D",X"A0",X"DD",X"9F",
		X"80",X"9F",X"2B",X"9F",X"DB",X"9E",X"90",X"9E",X"49",X"9E",X"0A",X"9E",X"CE",X"9D",X"98",X"9D",
		X"65",X"9D",X"37",X"9D",X"07",X"9D",X"11",X"9D",X"AA",X"9E",X"A8",X"A1",X"80",X"A5",X"E9",X"A9",
		X"A0",X"AE",X"86",X"B3",X"78",X"B8",X"6D",X"BD",X"54",X"C2",X"25",X"C7",X"DA",X"CB",X"75",X"D0",
		X"EC",X"D4",X"44",X"D9",X"7A",X"DD",X"91",X"E1",X"87",X"E5",X"5D",X"E9",X"10",X"ED",X"AA",X"F0",
		X"21",X"F4",X"7E",X"F7",X"BD",X"FA",X"E3",X"FD",X"E9",X"00",X"D9",X"03",X"B0",X"06",X"6F",X"09",
		X"15",X"0C",X"A6",X"0E",X"1D",X"11",X"80",X"13",X"CF",X"15",X"0A",X"18",X"31",X"1A",X"45",X"1C",
		X"45",X"1E",X"35",X"20",X"12",X"22",X"DE",X"23",X"9B",X"25",X"47",X"27",X"E2",X"28",X"72",X"2A",
		X"F2",X"2B",X"62",X"2D",X"C5",X"2E",X"1E",X"30",X"68",X"31",X"A4",X"32",X"D6",X"33",X"FB",X"34",
		X"16",X"36",X"27",X"37",X"18",X"38",X"92",X"37",X"86",X"35",X"92",X"32",X"FF",X"2E",X"11",X"2B",
		X"EB",X"26",X"AF",X"22",X"6A",X"1E",X"30",X"1A",X"02",X"16",X"ED",X"11",X"EE",X"0D",X"0E",X"0A",
		X"46",X"06",X"9E",X"02",X"13",X"FF",X"A4",X"FB",X"50",X"F8",X"1B",X"F5",X"FE",X"F1",X"FE",X"EE",
		X"16",X"EC",X"49",X"E9",X"93",X"E6",X"F6",X"E3",X"6E",X"E1",X"00",X"DF",X"A4",X"DC",X"5F",X"DA",
		X"2E",X"D8",X"12",X"D6",X"06",X"D4",X"10",X"D2",X"2B",X"D0",X"57",X"CE",X"94",X"CC",X"E1",X"CA",
		X"3F",X"C9",X"AC",X"C7",X"28",X"C6",X"B3",X"C4",X"4D",X"C3",X"F3",X"C1",X"A8",X"C0",X"68",X"BF",
		X"34",X"BE",X"0F",X"BD",X"F2",X"BB",X"E2",X"BA",X"DD",X"B9",X"E5",X"B8",X"F6",X"B7",X"0D",X"B7",
		X"31",X"B6",X"60",X"B5",X"97",X"B4",X"D7",X"B3",X"1E",X"B3",X"6E",X"B2",X"C8",X"B1",X"27",X"B1",
		X"8F",X"B0",X"FC",X"AF",X"73",X"AF",X"EF",X"AE",X"74",X"AE",X"FE",X"AD",X"8E",X"AD",X"25",X"AD",
		X"C1",X"AC",X"63",X"AC",X"0B",X"AC",X"B6",X"AB",X"69",X"AB",X"1F",X"AB",X"DC",X"AA",X"9C",X"AA",
		X"61",X"AA",X"29",X"AA",X"F7",X"A9",X"C8",X"A9",X"9F",X"A9",X"79",X"A9",X"56",X"A9",X"38",X"A9",
		X"1B",X"A9",X"03",X"A9",X"ED",X"A8",X"DD",X"A8",X"CD",X"A8",X"C3",X"A8",X"B9",X"A8",X"B4",X"A8",
		X"B2",X"A8",X"B2",X"A8",X"B3",X"A8",X"B6",X"A8",X"BE",X"A8",X"C5",X"A8",X"D0",X"A8",X"DE",X"A8",
		X"ED",X"A8",X"FD",X"A8",X"11",X"A9",X"26",X"A9",X"3D",X"A9",X"55",X"A9",X"70",X"A9",X"8A",X"A9",
		X"A9",X"A9",X"C6",X"A9",X"E8",X"A9",X"08",X"AA",X"2D",X"AA",X"50",X"AA",X"75",X"AA",X"9C",X"AA",
		X"C5",X"AA",X"EC",X"AA",X"18",X"AB",X"41",X"AB",X"6D",X"AB",X"9C",X"AB",X"CA",X"AB",X"F8",X"AB",
		X"28",X"AC",X"59",X"AC",X"8B",X"AC",X"BB",X"AC",X"F0",X"AC",X"22",X"AD",X"57",X"AD",X"8C",X"AD",
		X"C3",X"AD",X"F7",X"AD",X"2F",X"AE",X"5F",X"AE",X"D4",X"AE",X"E3",X"B0",X"47",X"B4",X"7F",X"B8",
		X"3C",X"BD",X"46",X"C2",X"76",X"C7",X"B2",X"CC",X"E8",X"D1",X"0F",X"D7",X"1D",X"DC",X"0D",X"E1",
		X"DD",X"E5",X"8B",X"EA",X"16",X"EF",X"7D",X"F3",X"BF",X"F7",X"E2",X"FB",X"E0",X"FF",X"BE",X"03",
		X"7C",X"07",X"1B",X"0B",X"96",X"0E",X"F9",X"11",X"39",X"15",X"66",X"18",X"68",X"1B",X"68",X"1E",
		X"6A",X"20",X"A0",X"20",X"B8",X"1F",X"02",X"1E",X"D2",X"1B",X"4C",X"19",X"9E",X"16",X"D1",X"13",
		X"FD",X"10",X"2C",X"0E",X"65",X"0B",X"A5",X"08",X"F9",X"05",X"5C",X"03",X"D6",X"00",X"5D",X"FE",
		X"FD",X"FB",X"AE",X"F9",X"73",X"F7",X"4A",X"F5",X"35",X"F3",X"30",X"F1",X"3B",X"EF",X"5A",X"ED",
		X"8A",X"EB",X"C8",X"E9",X"17",X"E8",X"75",X"E6",X"E3",X"E4",X"5E",X"E3",X"E6",X"E1",X"7C",X"E0",
		X"20",X"DF",X"CF",X"DD",X"8B",X"DC",X"53",X"DB",X"27",X"DA",X"05",X"D9",X"EE",X"D7",X"E3",X"D6",
		X"E1",X"D5",X"E9",X"D4",X"FA",X"D3",X"15",X"D3",X"39",X"D2",X"65",X"D1",X"9B",X"D0",X"D9",X"CF",
		X"1E",X"CF",X"6B",X"CE",X"C0",X"CD",X"1C",X"CD",X"7D",X"CC",X"E6",X"CB",X"57",X"CB",X"CC",X"CA",
		X"4A",X"CA",X"CC",X"C9",X"54",X"C9",X"E2",X"C8",X"75",X"C8",X"0E",X"C8",X"AC",X"C7",X"51",X"C7",
		X"F9",X"C6",X"A4",X"C6",X"55",X"C6",X"0A",X"C6",X"C3",X"C5",X"80",X"C5",X"42",X"C5",X"07",X"C5",
		X"D0",X"C4",X"9E",X"C4",X"6B",X"C4",X"40",X"C4",X"18",X"C4",X"F2",X"C3",X"CD",X"C3",X"AE",X"C3",
		X"8F",X"C3",X"77",X"C3",X"69",X"C3",X"B7",X"C4",X"92",X"C7",X"4E",X"CB",X"AC",X"CF",X"5D",X"D4",
		X"45",X"D9",X"3D",X"DE",X"37",X"E3",X"23",X"E8",X"FC",X"EC",X"B9",X"F1",X"58",X"F6",X"D3",X"FA",
		X"32",X"FF",X"6B",X"03",X"84",X"07",X"7A",X"0B",X"51",X"0F",X"05",X"13",X"9D",X"16",X"14",X"1A",
		X"6D",X"1D",X"A8",X"20",X"C8",X"23",X"CD",X"26",X"B7",X"29",X"86",X"2C",X"3D",X"2F",X"D9",X"31",
		X"63",X"34",X"D2",X"36",X"2C",X"39",X"6F",X"3B",X"9D",X"3D",X"B8",X"3F",X"C0",X"41",X"B3",X"43",
		X"95",X"45",X"65",X"47",X"22",X"49",X"D0",X"4A",X"6D",X"4C",X"FB",X"4D",X"77",X"4F",X"E8",X"50",
		X"48",X"52",X"9B",X"53",X"DF",X"54",X"18",X"56",X"43",X"57",X"63",X"58",X"74",X"59",X"80",X"5A",
		X"76",X"5B",X"6B",X"5C",X"29",X"5C",X"3E",X"5A",X"5C",X"57",X"C7",X"53",X"D5",X"4F",X"9F",X"4B",
		X"4D",X"47",X"F2",X"42",X"9F",X"3E",X"57",X"3A",X"26",X"36",X"0C",X"32",X"0C",X"2E",X"28",X"2A",
		X"63",X"26",X"BB",X"22",X"2D",X"1F",X"BE",X"1B",X"6A",X"18",X"32",X"15",X"14",X"12",X"0E",X"0F",
		X"22",X"0C",X"53",X"09",X"94",X"06",X"F8",X"03",X"5F",X"01",X"E3",X"FF",X"27",X"00",X"77",X"01",
		X"8E",X"03",X"15",X"06",X"EB",X"08",X"E5",X"0B",X"F9",X"0E",X"0C",X"12",X"1E",X"15",X"22",X"18",
		X"19",X"1B",X"F9",X"1D",X"C9",X"20",X"7F",X"23",X"22",X"26",X"AE",X"28",X"28",X"2B",X"89",X"2D",
		X"D6",X"2F",X"0D",X"32",X"32",X"34",X"41",X"36",X"3F",X"38",X"2B",X"3A",X"04",X"3C",X"CD",X"3D",
		X"83",X"3F",X"2B",X"41",X"C2",X"42",X"49",X"44",X"C1",X"45",X"2B",X"47",X"89",X"48",X"D7",X"49",
		X"19",X"4B",X"4E",X"4C",X"75",X"4D",X"92",X"4E",X"A1",X"4F",X"A9",X"50",X"A2",X"51",X"93",X"52",
		X"77",X"53",X"55",X"54",X"24",X"55",X"F1",X"55",X"AC",X"56",X"66",X"57",X"10",X"58",X"BD",X"58",
		X"56",X"59",X"F1",X"59",X"77",X"5A",X"10",X"5B",X"CE",X"5A",X"CC",X"58",X"BA",X"55",X"E7",X"51",
		X"AB",X"4D",X"27",X"49",X"87",X"44",X"DA",X"3F",X"35",X"3B",X"9C",X"36",X"1C",X"32",X"B4",X"2D",
		X"6A",X"29",X"3E",X"25",X"31",X"21",X"43",X"1D",X"76",X"19",X"C3",X"15",X"32",X"12",X"BD",X"0E",
		X"66",X"0B",X"2B",X"08",X"0A",X"05",X"03",X"02",X"1A",X"FF",X"45",X"FC",X"8A",X"F9",X"FD",X"F6",
		X"FB",X"F5",X"87",X"F6",X"04",X"F8",X"2D",X"FA",X"B7",X"FC",X"85",X"FF",X"73",X"02",X"73",X"05",
		X"71",X"08",X"6B",X"0B",X"5A",X"0E",X"3A",X"11",X"04",X"14",X"BC",X"16",X"5F",X"19",X"EC",X"1B",
		X"67",X"1E",X"C9",X"20",X"19",X"23",X"55",X"25",X"7C",X"27",X"8E",X"29",X"93",X"2B",X"7E",X"2D",
		X"60",X"2F",X"24",X"31",X"EF",X"32",X"09",X"34",X"59",X"33",X"7D",X"31",X"CD",X"2E",X"A2",X"2B",
		X"27",X"28",X"80",X"24",X"C5",X"20",X"09",X"1D",X"52",X"19",X"AA",X"15",X"14",X"12",X"97",X"0E",
		X"2F",X"0B",X"E3",X"07",X"AE",X"04",X"93",X"01",X"91",X"FE",X"A9",X"FB",X"D9",X"F8",X"21",X"F6",
		X"80",X"F3",X"F5",X"F0",X"80",X"EE",X"22",X"EC",X"D8",X"E9",X"A2",X"E7",X"7E",X"E5",X"6F",X"E3",
		X"72",X"E1",X"87",X"DF",X"AC",X"DD",X"E4",X"DB",X"2B",X"DA",X"81",X"D8",X"E6",X"D6",X"5C",X"D5",
		X"E0",X"D3",X"70",X"D2",X"11",X"D1",X"BE",X"CF",X"75",X"CE",X"3A",X"CD",X"0D",X"CC",X"E7",X"CA",
		X"D1",X"C9",X"C3",X"C8",X"C1",X"C7",X"C7",X"C6",X"DB",X"C5",X"F6",X"C4",X"1A",X"C4",X"46",X"C3",
		X"7F",X"C2",X"BD",X"C1",X"05",X"C1",X"54",X"C0",X"A8",X"BF",X"08",X"BF",X"6D",X"BE",X"DA",X"BD",
		X"4D",X"BD",X"C8",X"BC",X"48",X"BC",X"CF",X"BB",X"5C",X"BB",X"ED",X"BA",X"87",X"BA",X"23",X"BA",
		X"C8",X"B9",X"6E",X"B9",X"1D",X"B9",X"CC",X"B8",X"85",X"B8",X"3D",X"B8",X"FF",X"B7",X"BF",X"B7",
		X"8A",X"B7",X"52",X"B7",X"26",X"B7",X"F4",X"B6",X"D2",X"B6",X"A4",X"B6",X"98",X"B7",X"33",X"BA",
		X"C4",X"BD",X"02",X"C2",X"9F",X"C6",X"77",X"CB",X"64",X"D0",X"58",X"D5",X"3E",X"DA",X"14",X"DF",
		X"CF",X"E3",X"6D",X"E8",X"E9",X"EC",X"46",X"F1",X"83",X"F5",X"9D",X"F9",X"97",X"FD",X"6F",X"01",
		X"27",X"05",X"BF",X"08",X"3A",X"0C",X"96",X"0F",X"D6",X"12",X"F9",X"15",X"04",X"19",X"EE",X"1B",
		X"CA",X"1E",X"43",X"21",X"06",X"22",X"60",X"21",X"D2",X"1F",X"AD",X"1D",X"26",X"1B",X"65",X"18",
		X"83",X"15",X"97",X"12",X"A5",X"0F",X"BC",X"0C",X"DD",X"09",X"10",X"07",X"54",X"04",X"AB",X"01",
		X"17",X"FF",X"96",X"FC",X"29",X"FA",X"D0",X"F7",X"8A",X"F5",X"5A",X"F3",X"3B",X"F1",X"2E",X"EF",
		X"31",X"ED",X"4C",X"EB",X"6F",X"E9",X"AF",X"E7",X"E8",X"E5",X"1C",X"E5",X"13",X"E6",X"1B",X"E8",
		X"E6",X"EA",X"20",X"EE",X"A4",X"F1",X"4B",X"F5",X"06",X"F9",X"BC",X"FC",X"6C",X"00",X"09",X"04",
		X"95",X"07",X"08",X"0B",X"63",X"0E",X"A4",X"11",X"CE",X"14",X"DC",X"17",X"D2",X"1A",X"AD",X"1D",
		X"6F",X"20",X"1A",X"23",X"AF",X"25",X"29",X"28",X"91",X"2A",X"E2",X"2C",X"1D",X"2F",X"49",X"31",
		X"38",X"33",X"91",X"33",X"6D",X"32",X"5F",X"30",X"AF",X"2D",X"A3",X"2A",X"57",X"27",X"F2",X"23",
		X"7E",X"20",X"0D",X"1D",X"A5",X"19",X"4C",X"16",X"07",X"13",X"D6",X"0F",X"BC",X"0C",X"B9",X"09",
		X"CD",X"06",X"FB",X"03",X"3F",X"01",X"98",X"FE",X"09",X"FC",X"8E",X"F9",X"2B",X"F7",X"D6",X"F4",
		X"9F",X"F2",X"70",X"F0",X"62",X"EE",X"4F",X"EC",X"06",X"EB",X"8B",X"EB",X"31",X"ED",X"A7",X"EF",
		X"96",X"F2",X"D8",X"F5",X"3F",X"F9",X"BF",X"FC",X"3F",X"00",X"BA",X"03",X"26",X"07",X"83",X"0A",
		X"C9",X"0D",X"F9",X"10",X"0F",X"14",X"0E",X"17",X"F4",X"19",X"C3",X"1C",X"78",X"1F",X"18",X"22",
		X"A0",X"24",X"13",X"27",X"6D",X"29",X"B5",X"2B",X"E5",X"2D",X"06",X"30",X"10",X"32",X"FB",X"33",
		X"75",X"34",X"56",X"33",X"48",X"31",X"8E",X"2E",X"70",X"2B",X"12",X"28",X"96",X"24",X"0E",X"21",
		X"86",X"1D",X"05",X"1A",X"97",X"16",X"39",X"13",X"F4",X"0F",X"C4",X"0C",X"AB",X"09",X"AB",X"06",
		X"C3",X"03",X"F4",X"00",X"3B",X"FE",X"9A",X"FB",X"0C",X"F9",X"99",X"F6",X"35",X"F4",X"EB",X"F1",
		X"B1",X"EF",X"91",X"ED",X"73",X"EB",X"EC",X"E9",X"30",X"EA",X"B0",X"EB",X"05",X"EE",X"DF",X"F0",
		X"0D",X"F4",X"6A",X"F7",X"DE",X"FA",X"57",X"FE",X"CA",X"01",X"33",X"05",X"88",X"08",X"C9",X"0B",
		X"F4",X"0E",X"07",X"12",X"03",X"15",X"E7",X"17",X"B0",X"1A",X"65",X"1D",X"00",X"20",X"87",X"22",
		X"F6",X"24",X"51",X"27",X"94",X"29",X"C5",X"2B",X"E1",X"2D",X"EA",X"2F",X"DF",X"31",X"C6",X"33",
		X"98",X"35",X"5A",X"37",X"0D",X"39",X"AD",X"3A",X"3F",X"3C",X"C3",X"3D",X"35",X"3F",X"9D",X"40",
		X"F3",X"41",X"41",X"43",X"7D",X"44",X"AF",X"45",X"D4",X"46",X"EF",X"47",X"FD",X"48",X"01",X"4A",
		X"F8",X"4A",X"E7",X"4B",X"CC",X"4C",X"A7",X"4D",X"76",X"4E",X"40",X"4F",X"FD",X"4F",X"B6",X"50",
		X"5F",X"51",X"11",X"52",X"5B",X"52",X"F6",X"50",X"44",X"4E",X"C1",X"4A",X"B5",X"46",X"5D",X"42",
		X"DA",X"3D",X"45",X"39",X"B3",X"34",X"2D",X"30",X"B7",X"2B",X"5E",X"27",X"1F",X"23",X"FC",X"1E",
		X"F9",X"1A",X"14",X"17",X"4F",X"13",X"A8",X"0F",X"1D",X"0C",X"B0",X"08",X"61",X"05",X"2C",X"02",
		X"14",X"FF",X"15",X"FC",X"32",X"F9",X"65",X"F6",X"B0",X"F3",X"14",X"F1",X"8F",X"EE",X"1E",X"EC",
		X"C4",X"E9",X"7F",X"E7",X"4D",X"E5",X"2F",X"E3",X"23",X"E1",X"2C",X"DF",X"44",X"DD",X"6D",X"DB",
		X"A9",X"D9",X"F3",X"D7",X"50",X"D6",X"B9",X"D4",X"32",X"D3",X"BA",X"D1",X"4D",X"D0",X"F0",X"CE",
		X"A0",X"CD",X"5B",X"CC",X"26",X"CB",X"FA",X"C9",X"DB",X"C8",X"C4",X"C7",X"BC",X"C6",X"BA",X"C5",
		X"C6",X"C4",X"D9",X"C3",X"F8",X"C2",X"1F",X"C2",X"50",X"C1",X"89",X"C0",X"CA",X"BF",X"14",X"BF",
		X"66",X"BE",X"BF",X"BD",X"1F",X"BD",X"88",X"BC",X"F7",X"BB",X"6C",X"BB",X"E9",X"BA",X"6B",X"BA",
		X"F5",X"B9",X"83",X"B9",X"19",X"B9",X"B2",X"B8",X"53",X"B8",X"F8",X"B7",X"A0",X"B7",X"50",X"B7",
		X"03",X"B7",X"BC",X"B6",X"7A",X"B6",X"38",X"B6",X"1A",X"B6",X"78",X"B7",X"4E",X"BA",X"01",X"BE",
		X"4E",X"C2",X"EB",X"C6",X"BA",X"CB",X"9A",X"D0",X"7B",X"D5",X"4E",X"DA",X"0D",X"DF",X"B1",X"E3",
		X"38",X"E8",X"9F",X"EC",X"E6",X"F0",X"0C",X"F5",X"10",X"F9",X"F5",X"FC",X"B7",X"00",X"5C",X"04",
		X"E0",X"07",X"4B",X"0B",X"94",X"0E",X"C4",X"11",X"D3",X"14",X"D2",X"17",X"A8",X"1A",X"7C",X"1D",
		X"8F",X"1F",X"D1",X"1F",X"DF",X"1E",X"18",X"1D",X"CE",X"1A",X"2C",X"18",X"5B",X"15",X"6E",X"12",
		X"7A",X"0F",X"84",X"0C",X"9A",X"09",X"B9",X"06",X"EB",X"03",X"2F",X"01",X"89",X"FE",X"F5",X"FB",
		X"76",X"F9",X"0B",X"F7",X"B4",X"F4",X"71",X"F2",X"40",X"F0",X"24",X"EE",X"18",X"EC",X"1F",X"EA",
		X"38",X"E8",X"63",X"E6",X"9B",X"E4",X"E6",X"E2",X"40",X"E1",X"AA",X"DF",X"20",X"DE",X"A4",X"DC",
		X"37",X"DB",X"D8",X"D9",X"83",X"D8",X"3F",X"D7",X"03",X"D6",X"D4",X"D4",X"B0",X"D3",X"9A",X"D2",
		X"8A",X"D1",X"88",X"D0",X"8D",X"CF",X"9F",X"CE",X"B9",X"CD",X"DD",X"CC",X"08",X"CC",X"3D",X"CB",
		X"78",X"CA",X"BF",X"C9",X"08",X"C9",X"60",X"C8",X"B8",X"C7",X"22",X"C7",X"7D",X"C6",X"5C",X"C6",
		X"F1",X"C7",X"C5",X"CA",X"61",X"CE",X"7E",X"D2",X"E6",X"D6",X"73",X"DB",X"0E",X"E0",X"A6",X"E4",
		X"30",X"E9",X"A7",X"ED",X"04",X"F2",X"43",X"F6",X"64",X"FA",X"68",X"FE",X"4A",X"02",X"0E",X"06",
		X"B2",X"09",X"38",X"0D",X"A1",X"10",X"EC",X"13",X"1B",X"17",X"30",X"1A",X"27",X"1D",X"07",X"20",
		X"CB",X"22",X"7A",X"25",X"0D",X"28",X"8D",X"2A",X"F4",X"2C",X"45",X"2F",X"82",X"31",X"AB",X"33",
		X"BF",X"35",X"C0",X"37",X"AF",X"39",X"8D",X"3B",X"57",X"3D",X"12",X"3F",X"BA",X"40",X"56",X"42",
		X"DD",X"43",X"5B",X"45",X"C6",X"46",X"28",X"48",X"75",X"49",X"BC",X"4A",X"F0",X"4B",X"1C",X"4D",
		X"39",X"4E",X"4D",X"4F",X"53",X"50",X"52",X"51",X"3F",X"52",X"30",X"53",X"C5",X"53",X"AE",X"52",
		X"41",X"50",X"FD",X"4C",X"2E",X"49",X"0D",X"45",X"BE",X"40",X"5C",X"3C",X"F8",X"37",X"9E",X"33",
		X"55",X"2F",X"24",X"2B",X"0D",X"27",X"12",X"23",X"35",X"1F",X"73",X"1B",X"D1",X"17",X"4A",X"14",
		X"DF",X"10",X"94",X"0D",X"5E",X"0A",X"47",X"07",X"4A",X"04",X"67",X"01",X"9B",X"FE",X"E8",X"FB",
		X"4C",X"F9",X"C6",X"F6",X"55",X"F4",X"FB",X"F1",X"B3",X"EF",X"80",X"ED",X"61",X"EB",X"56",X"E9",
		X"5A",X"E7",X"73",X"E5",X"9B",X"E3",X"D5",X"E1",X"1C",X"E0",X"76",X"DE",X"DC",X"DC",X"54",X"DB",
		X"D8",X"D9",X"6B",X"D8",X"08",X"D7",X"B8",X"D5",X"6F",X"D4",X"36",X"D3",X"07",X"D2",X"E4",X"D0",
		X"CC",X"CF",X"BD",X"CE",X"B9",X"CD",X"C3",X"CC",X"D0",X"CB",X"12",X"CB",X"E6",X"CB",X"2C",X"CE",
		X"4E",X"D1",X"09",X"D5",X"17",X"D9",X"59",X"DD",X"AE",X"E1",X"08",X"E6",X"58",X"EA",X"97",X"EE",
		X"BF",X"F2",X"CE",X"F6",X"C0",X"FA",X"94",X"FE",X"49",X"02",X"E5",X"05",X"60",X"09",X"BF",X"0C",
		X"00",X"10",X"27",X"13",X"32",X"16",X"25",X"19",X"FC",X"1B",X"BB",X"1E",X"62",X"21",X"F1",X"23",
		X"6A",X"26",X"CB",X"28",X"18",X"2B",X"50",X"2D",X"72",X"2F",X"85",X"31",X"81",X"33",X"6C",X"35",
		X"45",X"37",X"0E",X"39",X"C4",X"3A",X"6B",X"3C",X"01",X"3E",X"88",X"3F",X"01",X"41",X"6E",X"42",
		X"C9",X"43",X"17",X"45",X"5A",X"46",X"90",X"47",X"B7",X"48",X"D5",X"49",X"E6",X"4A",X"EC",X"4B",
		X"E8",X"4C",X"D8",X"4D",X"C2",X"4E",X"9E",X"4F",X"5E",X"50",X"B2",X"4F",X"7C",X"4D",X"5F",X"4A",
		X"9E",X"46",X"86",X"42",X"32",X"3E",X"CD",X"39",X"5C",X"35",X"FA",X"30",X"A2",X"2C",X"66",X"28",
		X"3D",X"24",X"36",X"20",X"49",X"1C",X"7B",X"18",X"CB",X"14",X"37",X"11",X"C0",X"0D",X"66",X"0A",
		X"27",X"07",X"05",X"04",X"FD",X"00",X"0F",X"FE",X"3A",X"FB",X"7D",X"F8",X"D4",X"F5",X"47",X"F3",
		X"CE",X"F0",X"6B",X"EE",X"1D",X"EC",X"E2",X"E9",X"BC",X"E7",X"A8",X"E5",X"A8",X"E3",X"BA",X"E1",
		X"DC",X"DF",X"0F",X"DE",X"53",X"DC",X"A7",X"DA",X"09",X"D9",X"7B",X"D7",X"FA",X"D5",X"89",X"D4",
		X"26",X"D3",X"CF",X"D1",X"84",X"D0",X"47",X"CF",X"15",X"CE",X"EE",X"CC",X"D5",X"CB",X"C3",X"CA",
		X"C1",X"C9",X"C0",X"C8",X"D5",X"C7",X"EF",X"C6",X"4C",X"C7",X"4B",X"C9",X"3C",X"CC",X"DB",X"CF",
		X"D7",X"D3",X"13",X"D8",X"64",X"DC",X"C1",X"E0",X"13",X"E5",X"59",X"E9",X"89",X"ED",X"A0",X"F1",
		X"99",X"F5",X"78",X"F9",X"37",X"FD",X"D9",X"00",X"5E",X"04",X"C5",X"07",X"11",X"0B",X"40",X"0E",
		X"53",X"11",X"4F",X"14",X"2E",X"17",X"F5",X"19",X"A4",X"1C",X"3B",X"1F",X"BB",X"21",X"25",X"24",
		X"79",X"26",X"B8",X"28",X"E2",X"2A",X"FA",X"2C",X"FE",X"2E",X"EE",X"30",X"CF",X"32",X"9E",X"34",
		X"5B",X"36",X"09",X"38",X"A5",X"39",X"34",X"3B",X"B2",X"3C",X"24",X"3E",X"84",X"3F",X"DA",X"40",
		X"22",X"42",X"5D",X"43",X"8A",X"44",X"AE",X"45",X"C5",X"46",X"D0",X"47",X"D2",X"48",X"C8",X"49",
		X"B3",X"4A",X"95",X"4B",X"6D",X"4C",X"3C",X"4D",X"01",X"4E",X"BE",X"4E",X"74",X"4F",X"20",X"50",
		X"C5",X"50",X"60",X"51",X"F5",X"51",X"84",X"52",X"0B",X"53",X"8B",X"53",X"04",X"54",X"78",X"54",
		X"E3",X"54",X"4B",X"55",X"AB",X"55",X"08",X"56",X"5B",X"56",X"AD",X"56",X"F7",X"56",X"3F",X"57",
		X"82",X"57",X"BE",X"57",X"F7",X"57",X"2A",X"58",X"5B",X"58",X"87",X"58",X"AF",X"58",X"D3",X"58",
		X"F5",X"58",X"10",X"59",X"2A",X"59",X"40",X"59",X"51",X"59",X"61",X"59",X"6D",X"59",X"77",X"59",
		X"7F",X"59",X"83",X"59",X"83",X"59",X"82",X"59",X"7F",X"59",X"78",X"59",X"6F",X"59",X"65",X"59",
		X"58",X"59",X"4A",X"59",X"39",X"59",X"25",X"59",X"11",X"59",X"F8",X"58",X"E1",X"58",X"C7",X"58",
		X"AC",X"58",X"8D",X"58",X"6F",X"58",X"4E",X"58",X"2D",X"58",X"09",X"58",X"E5",X"57",X"BE",X"57",
		X"98",X"57",X"6F",X"57",X"46",X"57",X"19",X"57",X"EF",X"56",X"C2",X"56",X"96",X"56",X"65",X"56",
		X"36",X"56",X"06",X"56",X"D5",X"55",X"A1",X"55",X"70",X"55",X"3A",X"55",X"09",X"55",X"D1",X"54",
		X"9E",X"54",X"63",X"54",X"33",X"54",X"F3",X"53",X"CC",X"53",X"EF",X"52",X"5C",X"50",X"AD",X"4C",
		X"40",X"48",X"67",X"43",X"4B",X"3E",X"17",X"39",X"D8",X"33",X"A7",X"2E",X"83",X"29",X"7F",X"24",
		X"98",X"1F",X"D1",X"1A",X"2D",X"16",X"AE",X"11",X"4F",X"0D",X"17",X"09",X"FE",X"04",X"0B",X"01",
		X"35",X"FD",X"82",X"F9",X"EB",X"F5",X"78",X"F2",X"1F",X"EF",X"E5",X"EB",X"C3",X"E8",X"C0",X"E5",
		X"E2",X"E2",X"75",X"E1",X"AA",X"E1",X"D9",X"E2",X"BD",X"E4",X"0B",X"E7",X"A0",X"E9",X"58",X"EC",
		X"27",X"EF",X"FA",X"F1",X"C9",X"F4",X"8C",X"F7",X"45",X"FA",X"EB",X"FC",X"80",X"FF",X"01",X"02",
		X"6F",X"04",X"CB",X"06",X"11",X"09",X"47",X"0B",X"66",X"0D",X"79",X"0F",X"74",X"11",X"61",X"13",
		X"3B",X"15",X"09",X"17",X"BF",X"18",X"77",X"1A",X"9E",X"1B",X"02",X"1B",X"2A",X"19",X"7B",X"16",
		X"4D",X"13",X"CB",X"0F",X"1C",X"0C",X"5A",X"08",X"94",X"04",X"D6",X"00",X"26",X"FD",X"89",X"F9",
		X"05",X"F6",X"98",X"F2",X"44",X"EF",X"0B",X"EC",X"ED",X"E8",X"E8",X"E5",X"FC",X"E2",X"2B",X"E0",
		X"70",X"DD",X"CF",X"DA",X"42",X"D8",X"CF",X"D5",X"71",X"D3",X"28",X"D1",X"F4",X"CE",X"D6",X"CC",
		X"C8",X"CA",X"CF",X"C8",X"E8",X"C6",X"13",X"C5",X"4E",X"C3",X"9C",X"C1",X"F8",X"BF",X"65",X"BE",
		X"E0",X"BC",X"6B",X"BB",X"02",X"BA",X"AA",X"B8",X"5E",X"B7",X"21",X"B6",X"ED",X"B4",X"CA",X"B3",
		X"AD",X"B2",X"A2",X"B1",X"9D",X"B0",X"A5",X"AF",X"B7",X"AE",X"D3",X"AD",X"F9",X"AC",X"29",X"AC",
		X"60",X"AB",X"A6",X"AA",X"E8",X"A9",X"88",X"A9",X"D8",X"AA",X"78",X"AD",X"EB",X"B0",X"E8",X"B4",
		X"33",X"B9",X"A9",X"BD",X"33",X"C2",X"BA",X"C6",X"39",X"CB",X"A3",X"CF",X"F5",X"D3",X"2D",X"D8",
		X"47",X"DC",X"42",X"E0",X"21",X"E4",X"DF",X"E7",X"81",X"EB",X"02",X"EF",X"6D",X"F2",X"B4",X"F5",
		X"E5",X"F8",X"F8",X"FB",X"F4",X"FE",X"D1",X"01",X"9E",X"04",X"47",X"07",X"ED",X"09",X"7F",X"0B",
		X"4A",X"0B",X"08",X"0A",X"FC",X"07",X"7F",X"05",X"B4",X"02",X"C3",X"FF",X"B6",X"FC",X"AA",X"F9",
		X"9E",X"F6",X"9F",X"F3",X"AE",X"F0",X"D1",X"ED",X"05",X"EB",X"52",X"E8",X"B1",X"E5",X"27",X"E3",
		X"B2",X"E0",X"54",X"DE",X"07",X"DC",X"D1",X"D9",X"AC",X"D7",X"9C",X"D5",X"9E",X"D3",X"B5",X"D1",
		X"D9",X"CF",X"11",X"CE",X"58",X"CC",X"B2",X"CA",X"18",X"C9",X"8D",X"C7",X"14",X"C6",X"A7",X"C4",
		X"4B",X"C3",X"F8",X"C1",X"B5",X"C0",X"7D",X"BF",X"51",X"BE",X"31",X"BD",X"1E",X"BC",X"14",X"BB",
		X"16",X"BA",X"23",X"B9",X"39",X"B8",X"58",X"B7",X"83",X"B6",X"B4",X"B5",X"F3",X"B4",X"34",X"B4",
		X"83",X"B3",X"D5",X"B2",X"36",X"B2",X"93",X"B1",X"08",X"B1",X"6B",X"B0",X"A1",X"B0",X"93",X"B2",
		X"9D",X"B5",X"66",X"B9",X"9E",X"BD",X"18",X"C2",X"B2",X"C6",X"5A",X"CB",X"F8",X"CF",X"8B",X"D4",
		X"06",X"D9",X"68",X"DD",X"AC",X"E1",X"D3",X"E5",X"DA",X"E9",X"C1",X"ED",X"8A",X"F1",X"34",X"F5",
		X"BE",X"F8",X"2E",X"FC",X"7E",X"FF",X"B4",X"02",X"CD",X"05",X"CE",X"08",X"B3",X"0B",X"81",X"0E",
		X"34",X"11",X"BD",X"13",X"C2",X"14",X"33",X"14",X"B6",X"12",X"87",X"10",X"F6",X"0D",X"22",X"0B",
		X"2D",X"08",X"25",X"05",X"1F",X"02",X"1D",X"FF",X"29",X"FC",X"43",X"F9",X"6F",X"F6",X"B0",X"F3",
		X"05",X"F1",X"6F",X"EE",X"F0",X"EB",X"84",X"E9",X"2C",X"E7",X"E9",X"E4",X"B9",X"E2",X"A2",X"E0",
		X"96",X"DE",X"A0",X"DC",X"B7",X"DA",X"EA",X"D8",X"18",X"D7",X"EF",X"D5",X"8E",X"D6",X"61",X"D8",
		X"06",X"DB",X"27",X"DE",X"9C",X"E1",X"38",X"E5",X"EF",X"E8",X"A3",X"EC",X"54",X"F0",X"F3",X"F3",
		X"83",X"F7",X"FB",X"FA",X"58",X"FE",X"9E",X"01",X"CC",X"04",X"E1",X"07",X"DC",X"0A",X"BB",X"0D",
		X"87",X"10",X"38",X"13",X"D1",X"15",X"56",X"18",X"C4",X"1A",X"1B",X"1D",X"60",X"1F",X"8F",X"21",
		X"AA",X"23",X"B3",X"25",X"A8",X"27",X"8E",X"29",X"61",X"2B",X"23",X"2D",X"D6",X"2E",X"79",X"30",
		X"0B",X"32",X"90",X"33",X"04",X"35",X"6D",X"36",X"C6",X"37",X"14",X"39",X"55",X"3A",X"8A",X"3B",
		X"B1",X"3C",X"CE",X"3D",X"DF",X"3E",X"E5",X"3F",X"E1",X"40",X"D3",X"41",X"BB",X"42",X"9A",X"43",
		X"6E",X"44",X"39",X"45",X"FC",X"45",X"B8",X"46",X"69",X"47",X"14",X"48",X"B6",X"48",X"50",X"49",
		X"E5",X"49",X"71",X"4A",X"F8",X"4A",X"78",X"4B",X"F1",X"4B",X"64",X"4C",X"D1",X"4C",X"39",X"4D",
		X"99",X"4D",X"F5",X"4D",X"4D",X"4E",X"9D",X"4E",X"EB",X"4E",X"32",X"4F",X"76",X"4F",X"B4",X"4F",
		X"F0",X"4F",X"24",X"50",X"57",X"50",X"86",X"50",X"AF",X"50",X"D7",X"50",X"F9",X"50",X"18",X"51",
		X"34",X"51",X"4C",X"51",X"63",X"51",X"75",X"51",X"85",X"51",X"93",X"51",X"9E",X"51",X"A4",X"51",
		X"A9",X"51",X"AB",X"51",X"AD",X"51",X"AB",X"51",X"A4",X"51",X"9E",X"51",X"96",X"51",X"8B",X"51",
		X"7E",X"51",X"6F",X"51",X"5F",X"51",X"4B",X"51",X"39",X"51",X"22",X"51",X"0C",X"51",X"F1",X"50",
		X"D7",X"50",X"BA",X"50",X"A4",X"50",X"48",X"50",X"50",X"4E",X"01",X"4B",X"E1",X"46",X"3A",X"42",
		X"46",X"3D",X"2B",X"38",X"03",X"33",X"DF",X"2D",X"CB",X"28",X"D1",X"23",X"F2",X"1E",X"32",X"1A",
		X"96",X"15",X"1B",X"11",X"C3",X"0C",X"8E",X"08",X"7C",X"04",X"8C",X"00",X"BC",X"FC",X"0E",X"F9",
		X"7A",X"F5",X"0A",X"F2",X"B2",X"EE",X"7D",X"EB",X"5E",X"E8",X"66",X"E5",X"6F",X"E2",X"78",X"E0",
		X"4F",X"E0",X"3F",X"E1",X"01",X"E3",X"39",X"E5",X"C8",X"E7",X"7F",X"EA",X"53",X"ED",X"2C",X"F0",
		X"07",X"F3",X"D6",X"F5",X"9B",X"F8",X"4E",X"FB",X"F1",X"FD",X"7D",X"00",X"F9",X"02",X"62",X"05",
		X"B5",X"07",X"F7",X"09",X"24",X"0C",X"40",X"0E",X"48",X"10",X"40",X"12",X"26",X"14",X"FA",X"15",
		X"C0",X"17",X"75",X"19",X"1A",X"1B",X"B1",X"1C",X"3B",X"1E",X"B5",X"1F",X"22",X"21",X"83",X"22",
		X"D4",X"23",X"1A",X"25",X"56",X"26",X"84",X"27",X"A9",X"28",X"C2",X"29",X"D0",X"2A",X"D2",X"2B",
		X"CE",X"2C",X"BD",X"2D",X"A4",X"2E",X"82",X"2F",X"57",X"30",X"24",X"31",X"E6",X"31",X"A2",X"32",
		X"58",X"33",X"05",X"34",X"AB",X"34",X"49",X"35",X"E1",X"35",X"71",X"36",X"FC",X"36",X"80",X"37",
		X"FE",X"37",X"75",X"38",X"E9",X"38",X"56",X"39",X"BF",X"39",X"21",X"3A",X"7F",X"3A",X"D7",X"3A",
		X"2C",X"3B",X"7A",X"3B",X"C7",X"3B",X"0D",X"3C",X"50",X"3C",X"8E",X"3C",X"CA",X"3C",X"FF",X"3C",
		X"36",X"3D",X"63",X"3D",X"92",X"3D",X"B9",X"3D",X"E2",X"3D",X"01",X"3E",X"25",X"3E",X"3B",X"3E",
		X"65",X"3E",X"00",X"3E",X"E2",X"3B",X"95",X"38",X"83",X"34",X"FB",X"2F",X"2A",X"2B",X"3B",X"26",
		X"3F",X"21",X"4D",X"1C",X"67",X"17",X"9D",X"12",X"EE",X"0D",X"60",X"09",X"F1",X"04",X"A6",X"00",
		X"7B",X"FC",X"72",X"F8",X"8C",X"F4",X"C4",X"F0",X"1F",X"ED",X"96",X"E9",X"2C",X"E6",X"DF",X"E2",
		X"B2",X"DF",X"9D",X"DC",X"A7",X"D9",X"C8",X"D6",X"05",X"D4",X"59",X"D1",X"C7",X"CE",X"4A",X"CC",
		X"E5",X"C9",X"94",X"C7",X"5A",X"C5",X"34",X"C3",X"23",X"C1",X"24",X"BF",X"38",X"BD",X"5E",X"BB",
		X"96",X"B9",X"DE",X"B7",X"39",X"B6",X"A2",X"B4",X"1E",X"B3",X"A5",X"B1",X"3D",X"B0",X"E2",X"AE",
		X"94",X"AD",X"55",X"AC",X"23",X"AB",X"FC",X"A9",X"E2",X"A8",X"D6",X"A7",X"D2",X"A6",X"D9",X"A5",
		X"ED",X"A4",X"0A",X"A4",X"32",X"A3",X"63",X"A2",X"9E",X"A1",X"E2",X"A0",X"2E",X"A0",X"83",X"9F",
		X"E1",X"9E",X"47",X"9E",X"B6",X"9D",X"2A",X"9D",X"A5",X"9C",X"2A",X"9C",X"B4",X"9B",X"46",X"9B",
		X"DE",X"9A",X"7C",X"9A",X"1E",X"9A",X"C9",X"99",X"79",X"99",X"2D",X"99",X"E8",X"98",X"A6",X"98",
		X"6C",X"98",X"35",X"98",X"04",X"98",X"D7",X"97",X"AC",X"97",X"89",X"97",X"68",X"97",X"4B",X"97",
		X"32",X"97",X"1D",X"97",X"0B",X"97",X"FE",X"96",X"F2",X"96",X"EB",X"96",X"E7",X"96",X"E6",X"96",
		X"E7",X"96",X"ED",X"96",X"F3",X"96",X"FD",X"96",X"0B",X"97",X"1A",X"97",X"2B",X"97",X"3F",X"97",
		X"54",X"97",X"6E",X"97",X"88",X"97",X"A6",X"97",X"C2",X"97",X"E5",X"97",X"01",X"98",X"56",X"98",
		X"42",X"9A",X"8E",X"9D",X"AC",X"A1",X"57",X"A6",X"50",X"AB",X"71",X"B0",X"A1",X"B5",X"CE",X"BA",
		X"EB",X"BF",X"F1",X"C4",X"D9",X"C9",X"A4",X"CE",X"4A",X"D3",X"D1",X"D7",X"34",X"DC",X"75",X"E0",
		X"93",X"E4",X"91",X"E8",X"6D",X"EC",X"2B",X"F0",X"C7",X"F3",X"46",X"F7",X"A7",X"FA",X"EE",X"FD",
		X"15",X"01",X"23",X"04",X"16",X"07",X"F0",X"09",X"B2",X"0C",X"5D",X"0F",X"F0",X"11",X"6D",X"14",
		X"D4",X"16",X"24",X"19",X"62",X"1B",X"8A",X"1D",X"A0",X"1F",X"A4",X"21",X"94",X"23",X"73",X"25",
		X"43",X"27",X"FF",X"28",X"AD",X"2A",X"4B",X"2C",X"DB",X"2D",X"5A",X"2F",X"CC",X"30",X"32",X"32",
		X"89",X"33",X"D5",X"34",X"11",X"36",X"41",X"37",X"67",X"38",X"83",X"39",X"93",X"3A",X"99",X"3B",
		X"91",X"3C",X"83",X"3D",X"69",X"3E",X"46",X"3F",X"19",X"40",X"E5",X"40",X"A8",X"41",X"63",X"42",
		X"14",X"43",X"BF",X"43",X"5F",X"44",X"FC",X"44",X"8F",X"45",X"1D",X"46",X"A2",X"46",X"25",X"47",
		X"9B",X"47",X"12",X"48",X"7D",X"48",X"E7",X"48",X"46",X"49",X"A7",X"49",X"F9",X"49",X"51",X"4A",
		X"98",X"4A",X"F2",X"4A",X"A3",X"4A",X"98",X"48",X"69",X"45",X"73",X"41",X"0C",X"3D",X"5E",X"38",
		X"8F",X"33",X"B6",X"2E",X"E4",X"29",X"20",X"25",X"74",X"20",X"E4",X"1B",X"73",X"17",X"20",X"13",
		X"EE",X"0E",X"DB",X"0A",X"EA",X"06",X"1A",X"03",X"6C",X"FF",X"DA",X"FB",X"66",X"F8",X"10",X"F5",
		X"D7",X"F1",X"B8",X"EE",X"B7",X"EB",X"CA",X"E8",X"FF",X"E5",X"4E",X"E3",X"00",X"E2",X"59",X"E2",
		X"AE",X"E3",X"B9",X"E5",X"2E",X"E8",X"EC",X"EA",X"CC",X"ED",X"C4",X"F0",X"BC",X"F3",X"B2",X"F6",
		X"99",X"F9",X"75",X"FC",X"3C",X"FF",X"F2",X"01",X"91",X"04",X"21",X"07",X"99",X"09",X"FE",X"0B",
		X"4E",X"0E",X"8A",X"10",X"B4",X"12",X"CB",X"14",X"CE",X"16",X"C1",X"18",X"A3",X"1A",X"73",X"1C",
		X"32",X"1E",X"E3",X"1F",X"83",X"21",X"15",X"23",X"98",X"24",X"10",X"26",X"77",X"27",X"D1",X"28",
		X"20",X"2A",X"61",X"2B",X"97",X"2C",X"C1",X"2D",X"E0",X"2E",X"F5",X"2F",X"FD",X"30",X"FD",X"31",
		X"F3",X"32",X"DE",X"33",X"BF",X"34",X"98",X"35",X"68",X"36",X"31",X"37",X"F0",X"37",X"A7",X"38",
		X"57",X"39",X"FF",X"39",X"A1",X"3A",X"3A",X"3B",X"CD",X"3B",X"5A",X"3C",X"E0",X"3C",X"5F",X"3D",
		X"D8",X"3D",X"4D",X"3E",X"BB",X"3E",X"23",X"3F",X"84",X"3F",X"E4",X"3F",X"3E",X"40",X"91",X"40",
		X"E0",X"40",X"2D",X"41",X"73",X"41",X"B5",X"41",X"F4",X"41",X"2D",X"42",X"66",X"42",X"98",X"42",
		X"C6",X"42",X"F1",X"42",X"1A",X"43",X"40",X"43",X"61",X"43",X"80",X"43",X"9B",X"43",X"B4",X"43",
		X"CA",X"43",X"DD",X"43",X"ED",X"43",X"FC",X"43",X"07",X"44",X"0F",X"44",X"16",X"44",X"1B",X"44",
		X"1E",X"44",X"1F",X"44",X"1D",X"44",X"1B",X"44",X"15",X"44",X"0E",X"44",X"04",X"44",X"FA",X"43",
		X"ED",X"43",X"E1",X"43",X"D1",X"43",X"C1",X"43",X"AD",X"43",X"9B",X"43",X"84",X"43",X"70",X"43",
		X"56",X"43",X"41",X"43",X"1F",X"43",X"13",X"43",X"17",X"42",X"6A",X"3F",X"B8",X"3B",X"52",X"37",
		X"89",X"32",X"80",X"2D",X"64",X"28",X"3E",X"23",X"26",X"1E",X"22",X"19",X"39",X"14",X"6D",X"0F",
		X"C4",X"0A",X"3B",X"06",X"D8",X"01",X"96",X"FD",X"79",X"F9",X"7C",X"F5",X"A0",X"F1",X"E5",X"ED",
		X"4A",X"EA",X"CE",X"E6",X"70",X"E3",X"31",X"E0",X"0E",X"DD",X"04",X"DA",X"16",X"D7",X"44",X"D4",
		X"89",X"D1",X"EA",X"CE",X"5F",X"CC",X"EC",X"C9",X"8E",X"C7",X"48",X"C5",X"16",X"C3",X"F9",X"C0",
		X"EF",X"BE",X"F8",X"BC",X"13",X"BB",X"43",X"B9",X"81",X"B7",X"D4",X"B5",X"34",X"B4",X"A6",X"B2",
		X"22",X"B1",X"B5",X"AF",X"4F",X"AE",X"FC",X"AC",X"B4",X"AB",X"7C",X"AA",X"4C",X"A9",X"30",X"A8",
		X"17",X"A7",X"16",X"A6",X"08",X"A5",X"C1",X"A4",X"3D",X"A6",X"D8",X"A8",X"3A",X"AC",X"10",X"B0",
		X"30",X"B4",X"73",X"B8",X"C7",X"BC",X"16",X"C1",X"5B",X"C5",X"8E",X"C9",X"AA",X"CD",X"AA",X"D1",
		X"8F",X"D5",X"57",X"D9",X"05",X"DD",X"93",X"E0",X"06",X"E4",X"5D",X"E7",X"99",X"EA",X"BB",X"ED",
		X"C1",X"F0",X"B0",X"F3",X"85",X"F6",X"42",X"F9",X"E8",X"FB",X"78",X"FE",X"F1",X"00",X"55",X"03",
		X"A5",X"05",X"E2",X"07",X"0B",X"0A",X"20",X"0C",X"23",X"0E",X"16",X"10",X"F6",X"11",X"C5",X"13",
		X"86",X"15",X"36",X"17",X"D7",X"18",X"6A",X"1A",X"EE",X"1B",X"66",X"1D",X"CE",X"1E",X"2C",X"20",
		X"7A",X"21",X"BE",X"22",X"F6",X"23",X"21",X"25",X"42",X"26",X"59",X"27",X"64",X"28",X"66",X"29",
		X"5E",X"2A",X"4D",X"2B",X"31",X"2C",X"0E",X"2D",X"E0",X"2D",X"AB",X"2E",X"6F",X"2F",X"28",X"30",
		X"DC",X"30",X"88",X"31",X"2D",X"32",X"CB",X"32",X"61",X"33",X"F3",X"33",X"7C",X"34",X"FE",X"34",
		X"7F",X"35",X"F7",X"35",X"69",X"36",X"D5",X"36",X"3E",X"37",X"9F",X"37",X"FE",X"37",X"56",X"38",
		X"AC",X"38",X"FB",X"38",X"46",X"39",X"8E",X"39",X"D0",X"39",X"11",X"3A",X"4B",X"3A",X"84",X"3A",
		X"B8",X"3A",X"E9",X"3A",X"16",X"3B",X"41",X"3B",X"67",X"3B",X"8C",X"3B",X"AD",X"3B",X"CB",X"3B",
		X"E5",X"3B",X"FC",X"3B",X"13",X"3C",X"25",X"3C",X"38",X"3C",X"48",X"3C",X"54",X"3C",X"5D",X"3C",
		X"65",X"3C",X"6C",X"3C",X"6F",X"3C",X"73",X"3C",X"71",X"3C",X"71",X"3C",X"6E",X"3C",X"69",X"3C",
		X"61",X"3C",X"5A",X"3C",X"4F",X"3C",X"44",X"3C",X"3A",X"3C",X"2B",X"3C",X"1B",X"3C",X"0B",X"3C",
		X"F7",X"3B",X"E7",X"3B",X"D1",X"3B",X"BD",X"3B",X"A6",X"3B",X"8E",X"3B",X"74",X"3B",X"5C",X"3B",
		X"43",X"3B",X"27",X"3B",X"0C",X"3B",X"EF",X"3A",X"D1",X"3A",X"B3",X"3A",X"93",X"3A",X"74",X"3A",
		X"52",X"3A",X"33",X"3A",X"0C",X"3A",X"F2",X"39",X"95",X"39",X"A4",X"37",X"56",X"34",X"37",X"30",
		X"8F",X"2B",X"9C",X"26",X"80",X"21",X"58",X"1C",X"35",X"17",X"23",X"12",X"27",X"0D",X"4C",X"08",
		X"8F",X"03",X"F5",X"FE",X"7C",X"FA",X"29",X"F6",X"F7",X"F1",X"EA",X"ED",X"FC",X"E9",X"33",X"E6",
		X"88",X"E2",X"FE",X"DE",X"93",X"DB",X"44",X"D8",X"13",X"D5",X"00",X"D2",X"04",X"CF",X"27",X"CC",
		X"61",X"C9",X"B8",X"C6",X"23",X"C4",X"A9",X"C1",X"42",X"BF",X"F4",X"BC",X"BA",X"BA",X"96",X"B8",
		X"84",X"B6",X"8A",X"B4",X"9F",X"B2",X"CA",X"B0",X"02",X"AF",X"4F",X"AD",X"AC",X"AB",X"19",X"AA",
		X"96",X"A8",X"21",X"A7",X"BB",X"A5",X"64",X"A4",X"1B",X"A3",X"E0",X"A1",X"B1",X"A0",X"90",X"9F",
		X"7A",X"9E",X"70",X"9D",X"70",X"9C",X"99",X"9B",X"47",X"9C",X"73",X"9E",X"83",X"A1",X"30",X"A5",
		X"34",X"A9",X"72",X"AD",X"C3",X"B1",X"1D",X"B6",X"6C",X"BA",X"AE",X"BE",X"DA",X"C2",X"EE",X"C6",
		X"E5",X"CA",X"C3",X"CE",X"80",X"D2",X"24",X"D6",X"AB",X"D9",X"16",X"DD",X"62",X"E0",X"97",X"E3",
		X"AF",X"E6",X"B0",X"E9",X"97",X"EC",X"67",X"EF",X"1C",X"F2",X"BE",X"F4",X"46",X"F7",X"BB",X"F9",
		X"1C",X"FC",X"67",X"FE",X"9E",X"00",X"C3",X"02",X"D5",X"04",X"D6",X"06",X"C5",X"08",X"A3",X"0A",
		X"70",X"0C",X"2F",X"0E",X"DD",X"0F",X"7D",X"11",X"0D",X"13",X"90",X"14",X"07",X"16",X"6E",X"17",
		X"CB",X"18",X"1A",X"1A",X"60",X"1B",X"96",X"1C",X"C3",X"1D",X"E3",X"1E",X"FC",X"1F",X"07",X"21",
		X"0A",X"22",X"03",X"23",X"F2",X"23",X"D8",X"24",X"B7",X"25",X"8B",X"26",X"59",X"27",X"1E",X"28",
		X"DB",X"28",X"90",X"29",X"3E",X"2A",X"E5",X"2A",X"86",X"2B",X"1F",X"2C",X"B2",X"2C",X"3E",X"2D",
		X"C6",X"2D",X"46",X"2E",X"C2",X"2E",X"36",X"2F",X"A8",X"2F",X"12",X"30",X"7A",X"30",X"DA",X"30",
		X"38",X"31",X"90",X"31",X"E3",X"31",X"34",X"32",X"7D",X"32",X"C5",X"32",X"08",X"33",X"48",X"33",
		X"83",X"33",X"BC",X"33",X"F1",X"33",X"23",X"34",X"50",X"34",X"7C",X"34",X"A3",X"34",X"C8",X"34",
		X"EA",X"34",X"0B",X"35",X"27",X"35",X"43",X"35",X"5A",X"35",X"70",X"35",X"83",X"35",X"94",X"35",
		X"A3",X"35",X"B0",X"35",X"BA",X"35",X"C4",X"35",X"C9",X"35",X"D1",X"35",X"D1",X"35",X"D6",X"35",
		X"D0",X"35",X"D4",X"35",X"B0",X"34",X"EA",X"31",X"31",X"2E",X"CD",X"29",X"10",X"25",X"1A",X"20",
		X"10",X"1B",X"02",X"16",X"03",X"11",X"16",X"0C",X"46",X"07",X"94",X"02",X"03",X"FE",X"95",X"F9",
		X"48",X"F5",X"1E",X"F1",X"18",X"ED",X"32",X"E9",X"6D",X"E5",X"CA",X"E1",X"42",X"DE",X"DC",X"DA",
		X"94",X"D7",X"68",X"D4",X"57",X"D1",X"67",X"CE",X"84",X"CB",X"0D",X"C9",X"52",X"C8",X"FB",X"C8",
		X"88",X"CA",X"AF",X"CC",X"37",X"CF",X"F8",X"D1",X"D8",X"D4",X"C8",X"D7",X"B8",X"DA",X"A2",X"DD",
		X"81",X"E0",X"52",X"E3",X"0D",X"E6",X"BA",X"E8",X"50",X"EB",X"D8",X"ED",X"47",X"F0",X"A6",X"F2",
		X"EF",X"F4",X"26",X"F7",X"49",X"F9",X"5E",X"FB",X"5E",X"FD",X"4F",X"FF",X"2C",X"01",X"FC",X"02",
		X"BB",X"04",X"6C",X"06",X"0E",X"08",X"A0",X"09",X"25",X"0B",X"A0",X"0C",X"0A",X"0E",X"68",X"0F",
		X"BB",X"10",X"02",X"12",X"3C",X"13",X"6D",X"14",X"92",X"15",X"AC",X"16",X"BB",X"17",X"C3",X"18",
		X"BE",X"19",X"B4",X"1A",X"9E",X"1B",X"80",X"1C",X"58",X"1D",X"2B",X"1E",X"F4",X"1E",X"B6",X"1F",
		X"6F",X"20",X"22",X"21",X"CE",X"21",X"74",X"22",X"12",X"23",X"AA",X"23",X"3C",X"24",X"C8",X"24",
		X"4D",X"25",X"D0",X"25",X"49",X"26",X"C0",X"26",X"30",X"27",X"9D",X"27",X"03",X"28",X"66",X"28",
		X"C2",X"28",X"1E",X"29",X"70",X"29",X"C3",X"29",X"0E",X"2A",X"59",X"2A",X"9B",X"2A",X"E0",X"2A",
		X"1D",X"2B",X"59",X"2B",X"8D",X"2B",X"C4",X"2B",X"F1",X"2B",X"26",X"2C",X"48",X"2C",X"83",X"2C",
		X"F3",X"2B",X"A9",X"29",X"4D",X"26",X"31",X"22",X"AD",X"1D",X"E3",X"18",X"FF",X"13",X"11",X"0F",
		X"2F",X"0A",X"5C",X"05",X"A3",X"00",X"09",X"FC",X"8D",X"F7",X"30",X"F3",X"F9",X"EE",X"E1",X"EA",
		X"EC",X"E6",X"17",X"E3",X"64",X"DF",X"CF",X"DB",X"5B",X"D8",X"02",X"D5",X"CC",X"D1",X"AE",X"CE",
		X"AD",X"CB",X"C6",X"C8",X"FA",X"C5",X"5A",X"C3",X"37",X"C2",X"B0",X"C2",X"1A",X"C4",X"36",X"C6",
		X"B9",X"C8",X"80",X"CB",X"6A",X"CE",X"69",X"D1",X"67",X"D4",X"65",X"D7",X"55",X"DA",X"39",X"DD",
		X"09",X"E0",X"C9",X"E2",X"72",X"E5",X"0B",X"E8",X"8C",X"EA",X"FC",X"EC",X"56",X"EF",X"9F",X"F1",
		X"D2",X"F3",X"F6",X"F5",X"05",X"F8",X"06",X"FA",X"F5",X"FB",X"D2",X"FD",X"9F",X"FF",X"5E",X"01",
		X"0C",X"03",X"AE",X"04",X"40",X"06",X"C6",X"07",X"3C",X"09",X"A8",X"0A",X"05",X"0C",X"58",X"0D",
		X"9E",X"0E",X"DA",X"0F",X"09",X"11",X"2F",X"12",X"4A",X"13",X"58",X"14",X"60",X"15",X"5E",X"16",
		X"52",X"17",X"3C",X"18",X"1F",X"19",X"FA",X"19",X"CC",X"1A",X"97",X"1B",X"58",X"1C",X"13",X"1D",
		X"C9",X"1D",X"75",X"1E",X"1C",X"1F",X"BB",X"1F",X"55",X"20",X"E8",X"20",X"75",X"21",X"FD",X"21",
		X"80",X"22",X"FB",X"22",X"72",X"23",X"E4",X"23",X"52",X"24",X"BA",X"24",X"1D",X"25",X"7D",X"25",
		X"D8",X"25",X"2F",X"26",X"82",X"26",X"CF",X"26",X"1A",X"27",X"62",X"27",X"A4",X"27",X"E6",X"27",
		X"23",X"28",X"5C",X"28",X"91",X"28",X"C4",X"28",X"F5",X"28",X"21",X"29",X"4E",X"29",X"74",X"29",
		X"9A",X"29",X"BD",X"29",X"DC",X"29",X"F9",X"29",X"15",X"2A",X"2C",X"2A",X"45",X"2A",X"5A",X"2A",
		X"6E",X"2A",X"7F",X"2A",X"8E",X"2A",X"9B",X"2A",X"A7",X"2A",X"B1",X"2A",X"B9",X"2A",X"BE",X"2A",
		X"C4",X"2A",X"C6",X"2A",X"C9",X"2A",X"C9",X"2A",X"CA",X"2A",X"C5",X"2A",X"C5",X"2A",X"BE",X"2A",
		X"BF",X"2A",X"7B",X"2A",X"99",X"28",X"62",X"25",X"5A",X"21",X"C9",X"1C",X"EE",X"17",X"EC",X"12",
		X"DD",X"0D",X"D2",X"08",X"D7",X"03",X"F6",X"FE",X"30",X"FA",X"8C",X"F5",X"09",X"F1",X"A8",X"EC",
		X"6A",X"E8",X"4F",X"E4",X"55",X"E0",X"7F",X"DC",X"C8",X"D8",X"32",X"D5",X"BC",X"D1",X"65",X"CE",
		X"28",X"CB",X"10",X"C8",X"09",X"C5",X"2C",X"C2",X"4F",X"BF",X"74",X"BD",X"64",X"BD",X"73",X"BE",
		X"4E",X"C0",X"A1",X"C2",X"4B",X"C5",X"1C",X"C8",X"0B",X"CB",X"FF",X"CD",X"F4",X"D0",X"DD",X"D3",
		X"BD",X"D6",X"89",X"D9",X"48",X"DC",X"F1",X"DE",X"86",X"E1",X"08",X"E4",X"78",X"E6",X"D4",X"E8",
		X"1C",X"EB",X"51",X"ED",X"75",X"EF",X"86",X"F1",X"87",X"F3",X"76",X"F5",X"55",X"F7",X"26",X"F9",
		X"C6",X"FA",X"D7",X"FA",X"6A",X"F9",X"18",X"F7",X"25",X"F4",X"D9",X"F0",X"52",X"ED",X"B5",X"E9",
		X"08",X"E6",X"66",X"E2",X"CD",X"DE",X"49",X"DB",X"D6",X"D7",X"82",X"D4",X"43",X"D1",X"1F",X"CE",
		X"13",X"CB",X"24",X"C8",X"4C",X"C5",X"8F",X"C2",X"E8",X"BF",X"5C",X"BD",X"E6",X"BA",X"88",X"B8",
		X"3D",X"B6",X"0A",X"B4",X"EA",X"B1",X"E0",X"AF",X"E8",X"AD",X"05",X"AC",X"31",X"AA",X"71",X"A8",
		X"C2",X"A6",X"25",X"A5",X"96",X"A3",X"18",X"A2",X"AA",X"A0",X"48",X"9F",X"F8",X"9D",X"B3",X"9C",
		X"7D",X"9B",X"55",X"9A",X"39",X"99",X"28",X"98",X"23",X"97",X"2B",X"96",X"3E",X"95",X"5A",X"94",
		X"84",X"93",X"B3",X"92",X"F0",X"91",X"34",X"91",X"84",X"90",X"DA",X"8F",X"3D",X"8F",X"B0",X"8E",
		X"86",X"8F",X"EC",X"91",X"3B",X"95",X"2D",X"99",X"7D",X"9D",X"02",X"A2",X"9F",X"A6",X"41",X"AB",
		X"D9",X"AF",X"61",X"B4",X"D2",X"B8",X"2A",X"BD",X"63",X"C1",X"7F",X"C5",X"7C",X"C9",X"5C",X"CD",
		X"20",X"D1",X"C0",X"D4",X"48",X"D8",X"B0",X"DB",X"00",X"DF",X"32",X"E2",X"4C",X"E5",X"47",X"E8",
		X"30",X"EB",X"F8",X"ED",X"BC",X"F0",X"E5",X"F2",X"44",X"F3",X"5E",X"F2",X"9D",X"F0",X"54",X"EE",
		X"B2",X"EB",X"DD",X"E8",X"ED",X"E5",X"F6",X"E2",X"FA",X"DF",X"0F",X"DD",X"2C",X"DA",X"60",X"D7",
		X"A3",X"D4",X"FC",X"D1",X"69",X"CF",X"ED",X"CC",X"87",X"CA",X"35",X"C8",X"F7",X"C5",X"CF",X"C3",
		X"B9",X"C1",X"B9",X"BF",X"C8",X"BD",X"EE",X"BB",X"1D",X"BA",X"6A",X"B8",X"BD",X"B6",X"50",X"B6",
		X"8E",X"B7",X"CA",X"B9",X"BD",X"BC",X"14",X"C0",X"B2",X"C3",X"6D",X"C7",X"3A",X"CB",X"03",X"CF",
		X"C3",X"D2",X"72",X"D6",X"0F",X"DA",X"92",X"DD",X"FE",X"E0",X"51",X"E4",X"8B",X"E7",X"AB",X"EA",
		X"B2",X"ED",X"A1",X"F0",X"74",X"F3",X"34",X"F6",X"DD",X"F8",X"6F",X"FB",X"E9",X"FD",X"51",X"00",
		X"9F",X"02",X"E7",X"04",X"C3",X"06",X"E5",X"06",X"B0",X"05",X"9B",X"03",X"F3",X"00",X"F5",X"FD",
		X"C1",X"FA",X"72",X"F7",X"1B",X"F4",X"C6",X"F0",X"7F",X"ED",X"45",X"EA",X"1E",X"E7",X"0F",X"E4",
		X"16",X"E1",X"35",X"DE",X"6B",X"DB",X"B9",X"D8",X"1F",X"D6",X"99",X"D3",X"2A",X"D1",X"D2",X"CE",
		X"8F",X"CC",X"5F",X"CA",X"47",X"C8",X"3B",X"C6",X"4E",X"C4",X"61",X"C2",X"83",X"C1",X"66",X"C2",
		X"51",X"C4",X"03",X"C7",X"1E",X"CA",X"88",X"CD",X"12",X"D1",X"B4",X"D4",X"52",X"D8",X"EB",X"DB",
		X"73",X"DF",X"ED",X"E2",X"4B",X"E6",X"97",X"E9",X"C9",X"EC",X"E3",X"EF",X"E2",X"F2",X"CC",X"F5",
		X"9C",X"F8",X"56",X"FB",X"FA",X"FD",X"87",X"00",X"FD",X"02",X"60",X"05",X"AC",X"07",X"E9",X"09",
		X"0D",X"0C",X"22",X"0E",X"24",X"10",X"16",X"12",X"F3",X"13",X"C3",X"15",X"80",X"17",X"2E",X"19",
		X"CD",X"1A",X"60",X"1C",X"E1",X"1D",X"58",X"1F",X"BC",X"20",X"1C",X"22",X"62",X"23",X"BE",X"24",
		X"46",X"26",X"6B",X"27",X"93",X"28",X"A7",X"29",X"B8",X"2A",X"B7",X"2B",X"B3",X"2C",X"A0",X"2D",
		X"8A",X"2E",X"60",X"2F",X"3C",X"30",X"FE",X"30",X"D4",X"31",X"CE",X"31",X"0A",X"30",X"2B",X"2D",
		X"88",X"29",X"78",X"25",X"1F",X"21",X"A9",X"1C",X"24",X"18",X"A7",X"13",X"34",X"0F",X"DB",X"0A",
		X"9A",X"06",X"75",X"02",X"6E",X"FE",X"88",X"FA",X"BD",X"F6",X"15",X"F3",X"89",X"EF",X"19",X"EC",
		X"C8",X"E8",X"94",X"E5",X"7B",X"E2",X"7F",X"DF",X"9A",X"DC",X"D2",X"D9",X"21",X"D7",X"88",X"D4",
		X"1C",X"D2",X"37",X"D1",X"E9",X"D1",X"8F",X"D3",X"E1",X"D5",X"9A",X"D8",X"96",X"DB",X"B0",X"DE",
		X"DE",X"E1",X"0C",X"E5",X"34",X"E8",X"4E",X"EB",X"5A",X"EE",X"50",X"F1",X"36",X"F4",X"02",X"F7",
		X"BB",X"F9",X"5E",X"FC",X"EB",X"FE",X"62",X"01",X"C6",X"03",X"15",X"06",X"51",X"08",X"79",X"0A",
		X"8F",X"0C",X"94",X"0E",X"86",X"10",X"66",X"12",X"36",X"14",X"F6",X"15",X"A8",X"17",X"48",X"19",
		X"DD",X"1A",X"61",X"1C",X"D8",X"1D",X"42",X"1F",X"9E",X"20",X"EE",X"21",X"34",X"23",X"6A",X"24",
		X"97",X"25",X"B7",X"26",X"CE",X"27",X"DB",X"28",X"DC",X"29",X"D5",X"2A",X"C4",X"2B",X"A9",X"2C",
		X"85",X"2D",X"59",X"2E",X"24",X"2F",X"E8",X"2F",X"A3",X"30",X"58",X"31",X"03",X"32",X"A8",X"32",
		X"46",X"33",X"DD",X"33",X"6F",X"34",X"F8",X"34",X"7D",X"35",X"FD",X"35",X"74",X"36",X"E7",X"36",
		X"54",X"37",X"BE",X"37",X"20",X"38",X"7E",X"38",X"D8",X"38",X"2E",X"39",X"7D",X"39",X"C9",X"39",
		X"11",X"3A",X"55",X"3A",X"93",X"3A",X"D1",X"3A",X"09",X"3B",X"3D",X"3B",X"6E",X"3B",X"9D",X"3B",
		X"C6",X"3B",X"EE",X"3B",X"11",X"3C",X"35",X"3C",X"51",X"3C",X"6F",X"3C",X"88",X"3C",X"9E",X"3C",
		X"B1",X"3C",X"C4",X"3C",X"D1",X"3C",X"E0",X"3C",X"E9",X"3C",X"F4",X"3C",X"F8",X"3C",X"FE",X"3C",
		X"FF",X"3C",X"01",X"3D",X"FF",X"3C",X"FE",X"3C",X"F7",X"3C",X"F2",X"3C",X"E9",X"3C",X"E1",X"3C",
		X"D5",X"3C",X"CA",X"3C",X"BB",X"3C",X"AF",X"3C",X"99",X"3C",X"92",X"3C",X"3A",X"3C",X"40",X"3A",
		X"EE",X"36",X"CC",X"32",X"24",X"2E",X"2D",X"29",X"13",X"24",X"EB",X"1E",X"C8",X"19",X"B4",X"14",
		X"BB",X"0F",X"DF",X"0A",X"23",X"06",X"89",X"01",X"14",X"FD",X"BD",X"F8",X"8D",X"F4",X"80",X"F0",
		X"93",X"EC",X"C8",X"E8",X"20",X"E5",X"92",X"E1",X"2A",X"DE",X"D8",X"DA",X"AB",X"D7",X"93",X"D4",
		X"A1",X"D1",X"B3",X"CE",X"D1",X"CC",X"C1",X"CC",X"CA",X"CD",X"A1",X"CF",X"F1",X"D1",X"95",X"D4",
		X"63",X"D7",X"4F",X"DA",X"3D",X"DD",X"2F",X"E0",X"14",X"E3",X"EE",X"E5",X"B8",X"E8",X"6F",X"EB",
		X"13",X"EE",X"A3",X"F0",X"20",X"F3",X"89",X"F5",X"DD",X"F7",X"20",X"FA",X"4F",X"FC",X"6C",X"FE",
		X"75",X"00",X"6F",X"02",X"57",X"04",X"30",X"06",X"FB",X"07",X"8D",X"09",X"8A",X"09",X"09",X"08",
		X"9F",X"05",X"98",X"02",X"35",X"FF",X"9B",X"FB",X"E6",X"F7",X"29",X"F4",X"71",X"F0",X"C4",X"EC",
		X"2A",X"E9",X"A8",X"E5",X"3D",X"E2",X"EB",X"DE",X"B4",X"DB",X"99",X"D8",X"94",X"D5",X"AD",X"D2",
		X"DD",X"CF",X"28",X"CD",X"88",X"CA",X"03",X"C8",X"90",X"C5",X"39",X"C3",X"F1",X"C0",X"CA",X"BE",
		X"A0",X"BC",X"47",X"BB",X"BF",X"BB",X"60",X"BD",X"D4",X"BF",X"C1",X"C2",X"03",X"C6",X"6D",X"C9",
		X"F1",X"CC",X"76",X"D0",X"F9",X"D3",X"6C",X"D7",X"D4",X"DA",X"21",X"DE",X"5D",X"E1",X"7F",X"E4",
		X"8B",X"E7",X"7E",X"EA",X"5B",X"ED",X"1F",X"F0",X"CF",X"F2",X"68",X"F5",X"EB",X"F7",X"57",X"FA",
		X"B3",X"FC",X"F5",X"FE",X"29",X"01",X"44",X"03",X"44",X"05",X"CB",X"05",X"BA",X"04",X"B6",X"02",
		X"06",X"00",X"F5",X"FC",X"A2",X"F9",X"32",X"F6",X"B1",X"F2",X"36",X"EF",X"C3",X"EB",X"62",X"E8",
		X"14",X"E5",X"DB",X"E1",X"BA",X"DE",X"B2",X"DB",X"C2",X"D8",X"EB",X"D5",X"2D",X"D3",X"87",X"D0",
		X"F8",X"CD",X"80",X"CB",X"1F",X"C9",X"D2",X"C6",X"9B",X"C4",X"76",X"C2",X"6D",X"C0",X"64",X"BE",
		X"F8",X"BC",X"5D",X"BD",X"FE",X"BE",X"78",X"C1",X"75",X"C4",X"CC",X"C7",X"4B",X"CB",X"E5",X"CE",
		X"84",X"D2",X"20",X"D6",X"AD",X"D9",X"2B",X"DD",X"93",X"E0",X"E4",X"E3",X"1D",X"E7",X"3D",X"EA",
		X"47",X"ED",X"38",X"F0",X"11",X"F3",X"D1",X"F5",X"7D",X"F8",X"11",X"FB",X"90",X"FD",X"F9",X"FF",
		X"4E",X"02",X"8D",X"04",X"BB",X"06",X"D6",X"08",X"E0",X"0A",X"D5",X"0C",X"BC",X"0E",X"90",X"10",
		X"57",X"12",X"0B",X"14",X"B0",X"15",X"47",X"17",X"D1",X"18",X"4C",X"1A",X"BB",X"1B",X"1C",X"1D",
		X"6F",X"1E",X"B7",X"1F",X"F4",X"20",X"23",X"22",X"49",X"23",X"65",X"24",X"74",X"25",X"7B",X"26",
		X"77",X"27",X"68",X"28",X"51",X"29",X"32",X"2A",X"09",X"2B",X"D8",X"2B",X"9E",X"2C",X"5C",X"2D",
		X"15",X"2E",X"C5",X"2E",X"6E",X"2F",X"0E",X"30",X"A9",X"30",X"3D",X"31",X"CB",X"31",X"53",X"32",
		X"D5",X"32",X"51",X"33",X"C6",X"33",X"37",X"34",X"A2",X"34",X"0A",X"35",X"6B",X"35",X"C7",X"35",
		X"1F",X"36",X"73",X"36",X"C2",X"36",X"0C",X"37",X"53",X"37",X"95",X"37",X"D4",X"37",X"11",X"38",
		X"48",X"38",X"7A",X"38",X"AC",X"38",X"DA",X"38",X"03",X"39",X"2B",X"39",X"50",X"39",X"73",X"39",
		X"8F",X"39",X"AB",X"39",X"C4",X"39",X"DA",X"39",X"EF",X"39",X"01",X"3A",X"0F",X"3A",X"1E",X"3A",
		X"2A",X"3A",X"32",X"3A",X"3A",X"3A",X"40",X"3A",X"42",X"3A",X"44",X"3A",X"45",X"3A",X"43",X"3A",
		X"3E",X"3A",X"39",X"3A",X"33",X"3A",X"2B",X"3A",X"20",X"3A",X"15",X"3A",X"0A",X"3A",X"FB",X"39",
		X"ED",X"39",X"DC",X"39",X"CB",X"39",X"B9",X"39",X"A4",X"39",X"92",X"39",X"7B",X"39",X"65",X"39",
		X"4C",X"39",X"35",X"39",X"1B",X"39",X"01",X"39",X"E6",X"38",X"CA",X"38",X"AF",X"38",X"91",X"38",
		X"73",X"38",X"55",X"38",X"34",X"38",X"15",X"38",X"F6",X"37",X"D4",X"37",X"B3",X"37",X"90",X"37",
		X"6D",X"37",X"4B",X"37",X"26",X"37",X"03",X"37",X"DE",X"36",X"B9",X"36",X"96",X"36",X"6E",X"36",
		X"48",X"36",X"22",X"36",X"FC",X"35",X"D2",X"35",X"AC",X"35",X"85",X"35",X"5E",X"35",X"34",X"35",
		X"0D",X"35",X"E3",X"34",X"BB",X"34",X"90",X"34",X"68",X"34",X"3F",X"34",X"15",X"34",X"EA",X"33",
		X"C2",X"33",X"96",X"33",X"6B",X"33",X"40",X"33",X"17",X"33",X"EB",X"32",X"C1",X"32",X"96",X"32",
		X"6B",X"32",X"3D",X"32",X"15",X"32",X"E9",X"31",X"BD",X"31",X"92",X"31",X"67",X"31",X"3A",X"31",
		X"10",X"31",X"E3",X"30",X"B9",X"30",X"8B",X"30",X"62",X"30",X"34",X"30",X"0A",X"30",X"DC",X"2F",
		X"B2",X"2F",X"85",X"2F",X"5A",X"2F",X"2C",X"2F",X"04",X"2F",X"D6",X"2E",X"AC",X"2E",X"7C",X"2E",
		X"59",X"2E",X"F6",X"2D",X"93",X"2B",X"DF",X"27",X"77",X"23",X"92",X"1E",X"73",X"19",X"31",X"14",
		X"EC",X"0E",X"AE",X"09",X"88",X"04",X"77",X"FF",X"8A",X"FA",X"BB",X"F5",X"13",X"F1",X"8D",X"EC",
		X"2C",X"E8",X"F0",X"E3",X"D7",X"DF",X"E0",X"DB",X"0E",X"D8",X"5C",X"D4",X"CA",X"D0",X"57",X"CD",
		X"01",X"CA",X"CC",X"C6",X"B0",X"C3",X"B6",X"C0",X"DB",X"BD",X"69",X"BC",X"AD",X"BC",X"F1",X"BD",
		X"F3",X"BF",X"5F",X"C2",X"1A",X"C5",X"F6",X"C7",X"ED",X"CA",X"E4",X"CD",X"DD",X"D0",X"C7",X"D3",
		X"A7",X"D6",X"74",X"D9",X"31",X"DC",X"DA",X"DE",X"71",X"E1",X"F1",X"E3",X"5F",X"E6",X"B8",X"E8",
		X"01",X"EB",X"33",X"ED",X"57",X"EF",X"68",X"F1",X"69",X"F3",X"57",X"F5",X"35",X"F7",X"03",X"F9",
		X"C2",X"FA",X"73",X"FC",X"15",X"FE",X"AA",X"FF",X"2F",X"01",X"A9",X"02",X"15",X"04",X"76",X"05",
		X"CA",X"06",X"12",X"08",X"4F",X"09",X"80",X"0A",X"A9",X"0B",X"C7",X"0C",X"DB",X"0D",X"E4",X"0E",
		X"E3",X"0F",X"D9",X"10",X"C9",X"11",X"AE",X"12",X"8C",X"13",X"61",X"14",X"2D",X"15",X"F4",X"15",
		X"B2",X"16",X"6A",X"17",X"1B",X"18",X"C6",X"18",X"68",X"19",X"07",X"1A",X"9C",X"1A",X"2E",X"1B",
		X"B9",X"1B",X"3F",X"1C",X"C0",X"1C",X"3B",X"1D",X"B0",X"1D",X"22",X"1E",X"8F",X"1E",X"F6",X"1E",
		X"5A",X"1F",X"BB",X"1F",X"15",X"20",X"6B",X"20",X"BD",X"20",X"0E",X"21",X"59",X"21",X"A2",X"21",
		X"E6",X"21",X"28",X"22",X"64",X"22",X"9F",X"22",X"D8",X"22",X"0C",X"23",X"3E",X"23",X"6C",X"23",
		X"98",X"23",X"C1",X"23",X"EA",X"23",X"0E",X"24",X"30",X"24",X"50",X"24",X"6F",X"24",X"8B",X"24",
		X"A5",X"24",X"BC",X"24",X"D3",X"24",X"E5",X"24",X"F8",X"24",X"08",X"25",X"17",X"25",X"23",X"25",
		X"30",X"25",X"38",X"25",X"41",X"25",X"48",X"25",X"4D",X"25",X"51",X"25",X"54",X"25",X"55",X"25",
		X"55",X"25",X"55",X"25",X"51",X"25",X"4E",X"25",X"4B",X"25",X"45",X"25",X"3E",X"25",X"37",X"25",
		X"2F",X"25",X"26",X"25",X"1B",X"25",X"11",X"25",X"05",X"25",X"F7",X"24",X"EB",X"24",X"DD",X"24",
		X"CD",X"24",X"BF",X"24",X"AE",X"24",X"9E",X"24",X"8E",X"24",X"7A",X"24",X"67",X"24",X"55",X"24",
		X"42",X"24",X"2D",X"24",X"19",X"24",X"02",X"24",X"EF",X"23",X"D7",X"23",X"C2",X"23",X"AB",X"23",
		X"95",X"23",X"7D",X"23",X"66",X"23",X"4D",X"23",X"33",X"23",X"1B",X"23",X"02",X"23",X"E8",X"22",
		X"CE",X"22",X"B5",X"22",X"9A",X"22",X"80",X"22",X"64",X"22",X"4A",X"22",X"2F",X"22",X"13",X"22",
		X"F8",X"21",X"DD",X"21",X"C0",X"21",X"A3",X"21",X"86",X"21",X"6C",X"21",X"4D",X"21",X"32",X"21",
		X"15",X"21",X"E5",X"20",X"45",X"1F",X"20",X"1C",X"18",X"18",X"75",X"13",X"7C",X"0E",X"54",X"09",
		X"1C",X"04",X"E6",X"FE",X"C1",X"F9",X"B2",X"F4",X"C2",X"EF",X"F2",X"EA",X"47",X"E6",X"BD",X"E1",
		X"58",X"DD",X"18",X"D9",X"F9",X"D4",X"01",X"D1",X"2A",X"CD",X"73",X"C9",X"DD",X"C5",X"6A",X"C2",
		X"12",X"BF",X"DC",X"BB",X"BE",X"B8",X"C5",X"B5",X"D2",X"B2",X"93",X"B0",X"2C",X"B0",X"0B",X"B1",
		X"CA",X"B2",X"14",X"B5",X"B9",X"B7",X"94",X"BA",X"8D",X"BD",X"8F",X"C0",X"95",X"C3",X"90",X"C6",
		X"84",X"C9",X"64",X"CC",X"34",X"CF",X"F1",X"D1",X"9A",X"D4",X"2E",X"D7",X"B2",X"D9",X"1F",X"DC",
		X"7C",X"DE",X"C2",X"E0",X"F9",X"E2",X"1B",X"E5",X"30",X"E7",X"2F",X"E9",X"22",X"EB",X"FE",X"EC",
		X"CE",X"EE",X"4A",X"EF",X"18",X"EE",X"EC",X"EB",X"06",X"E9",X"C1",X"E5",X"36",X"E2",X"8E",X"DE",
		X"D9",X"DA",X"25",X"D7",X"7D",X"D3",X"E9",X"CF",X"67",X"CC",X"00",X"C9",X"B1",X"C5",X"7E",X"C2",
		X"66",X"BF",X"67",X"BC",X"83",X"B9",X"B9",X"B6",X"0A",X"B4",X"6F",X"B1",X"F1",X"AE",X"86",X"AC",
		X"36",X"AA",X"F7",X"A7",X"D5",X"A5",X"B5",X"A3",X"16",X"A2",X"3E",X"A2",X"BF",X"A3",X"1F",X"A6",
		X"12",X"A9",X"5D",X"AC",X"DD",X"AF",X"77",X"B3",X"19",X"B7",X"B9",X"BA",X"4D",X"BE",X"D0",X"C1",
		X"41",X"C5",X"9B",X"C8",X"DE",X"CB",X"08",X"CF",X"1B",X"D2",X"17",X"D5",X"FC",X"D7",X"C8",X"DA",
		X"7F",X"DD",X"1F",X"E0",X"AB",X"E2",X"1F",X"E5",X"84",X"E7",X"CF",X"E9",X"0B",X"EC",X"34",X"EE",
		X"4C",X"F0",X"4F",X"F2",X"45",X"F4",X"27",X"F6",X"FD",X"F7",X"BF",X"F9",X"76",X"FB",X"1B",X"FD",
		X"B4",X"FE",X"3C",X"00",X"BB",X"01",X"2B",X"03",X"8F",X"04",X"E8",X"05",X"35",X"07",X"75",X"08",
		X"AB",X"09",X"D5",X"0A",X"F6",X"0B",X"0D",X"0D",X"1A",X"0E",X"1D",X"0F",X"19",X"10",X"09",X"11",
		X"F2",X"11",X"D0",X"12",X"AF",X"13",X"46",X"14",X"34",X"13",X"BC",X"10",X"66",X"0D",X"7F",X"09",
		X"45",X"05",X"DC",X"00",X"62",X"FC",X"E6",X"F7",X"74",X"F3",X"17",X"EF",X"D2",X"EA",X"AA",X"E6",
		X"A0",X"E2",X"B5",X"DE",X"E7",X"DA",X"39",X"D7",X"AA",X"D3",X"3C",X"D0",X"E8",X"CC",X"B7",X"C9",
		X"9D",X"C6",X"A2",X"C3",X"BD",X"C0",X"FB",X"BD",X"48",X"BB",X"BB",X"B8",X"2E",X"B6",X"9B",X"B4",
		X"DF",X"B4",X"41",X"B6",X"78",X"B8",X"25",X"BB",X"29",X"BE",X"53",X"C1",X"9B",X"C4",X"E3",X"C7",
		X"2C",X"CB",X"69",X"CE",X"98",X"D1",X"B2",X"D4",X"BA",X"D7",X"AD",X"DA",X"8B",X"DD",X"4F",X"E0",
		X"02",X"E3",X"9C",X"E5",X"25",X"E8",X"93",X"EA",X"F3",X"EC",X"3A",X"EF",X"75",X"F1",X"97",X"F3",
		X"AD",X"F5",X"AE",X"F7",X"81",X"F9",X"C1",X"F9",X"79",X"F8",X"3E",X"F6",X"65",X"F3",X"26",X"F0",
		X"B3",X"EC",X"1C",X"E9",X"80",X"E5",X"E5",X"E1",X"5A",X"DE",X"D8",X"DA",X"78",X"D7",X"20",X"D4",
		X"F6",X"D0",X"B4",X"CD",X"3F",X"CA",X"56",X"C7",X"7C",X"C4",X"C1",X"C1",X"18",X"BF",X"8B",X"BC",
		X"16",X"BA",X"B4",X"B7",X"6D",X"B5",X"35",X"B3",X"1D",X"B1",X"02",X"AF",X"AC",X"AD",X"31",X"AE",
		X"EA",X"AF",X"7C",X"B2",X"8E",X"B5",X"F4",X"B8",X"88",X"BC",X"34",X"C0",X"E2",X"C3",X"8E",X"C7",
		X"2A",X"CB",X"B8",X"CE",X"2D",X"D2",X"8E",X"D5",X"D6",X"D8",X"05",X"DC",X"1E",X"DF",X"1D",X"E2",
		X"04",X"E5",X"D4",X"E7",X"8D",X"EA",X"31",X"ED",X"BC",X"EF",X"34",X"F2",X"97",X"F4",X"E5",X"F6",
		X"20",X"F9",X"49",X"FB",X"5F",X"FD",X"62",X"FF",X"54",X"01",X"37",X"03",X"0A",X"05",X"CB",X"06",
		X"7D",X"08",X"22",X"0A",X"B8",X"0B",X"3E",X"0D",X"BB",X"0E",X"26",X"10",X"88",X"11",X"DB",X"12",
		X"25",X"14",X"61",X"15",X"92",X"16",X"B9",X"17",X"D5",X"18",X"E6",X"19",X"EF",X"1A",X"ED",X"1B",
		X"E2",X"1C",X"CE",X"1D",X"B1",X"1E",X"8A",X"1F",X"5D",X"20",X"27",X"21",X"EB",X"21",X"A5",X"22",
		X"5A",X"23",X"06",X"24",X"AC",X"24",X"4C",X"25",X"E6",X"25",X"78",X"26",X"04",X"27",X"8B",X"27",
		X"0C",X"28",X"86",X"28",X"FD",X"28",X"6E",X"29",X"DA",X"29",X"42",X"2A",X"A4",X"2A",X"03",X"2B",
		X"5A",X"2B",X"B1",X"2B",X"01",X"2C",X"4F",X"2C",X"98",X"2C",X"DE",X"2C",X"1E",X"2D",X"5E",X"2D",
		X"98",X"2D",X"D1",X"2D",X"04",X"2E",X"37",X"2E",X"65",X"2E",X"90",X"2E",X"B8",X"2E",X"DE",X"2E",
		X"00",X"2F",X"22",X"2F",X"40",X"2F",X"5B",X"2F",X"74",X"2F",X"8D",X"2F",X"A1",X"2F",X"B4",X"2F",
		X"C3",X"2F",X"D4",X"2F",X"DF",X"2F",X"EB",X"2F",X"F2",X"2F",X"FC",X"2F",X"00",X"30",X"07",X"30",
		X"06",X"30",X"0B",X"30",X"05",X"30",X"0D",X"30",X"BD",X"2F",X"BE",X"2D",X"66",X"2A",X"39",X"26",
		X"85",X"21",X"85",X"1C",X"5E",X"17",X"2A",X"12",X"FB",X"0C",X"DD",X"07",X"D9",X"02",X"F3",X"FD",
		X"2E",X"F9",X"8A",X"F4",X"0B",X"F0",X"B0",X"EB",X"78",X"E7",X"63",X"E3",X"72",X"DF",X"A1",X"DB",
		X"F3",X"D7",X"61",X"D4",X"F4",X"D0",X"A1",X"CD",X"72",X"CA",X"55",X"C7",X"62",X"C4",X"74",X"C1",
		X"A0",X"BF",X"A3",X"BF",X"C2",X"C0",X"B4",X"C2",X"1D",X"C5",X"DE",X"C7",X"C9",X"CA",X"CE",X"CD",
		X"D9",X"D0",X"E5",X"D3",X"E3",X"D6",X"D9",X"D9",X"BB",X"DC",X"8C",X"DF",X"47",X"E2",X"F2",X"E4",
		X"86",X"E7",X"05",X"EA",X"71",X"EC",X"C9",X"EE",X"0D",X"F1",X"41",X"F3",X"61",X"F5",X"70",X"F7",
		X"6B",X"F9",X"59",X"FB",X"33",X"FD",X"02",X"FF",X"BC",X"00",X"6A",X"02",X"08",X"04",X"9A",X"05",
		X"1E",X"07",X"94",X"08",X"FD",X"09",X"5C",X"0B",X"AC",X"0C",X"F1",X"0D",X"2C",X"0F",X"5B",X"10",
		X"7E",X"11",X"99",X"12",X"A9",X"13",X"AF",X"14",X"AD",X"15",X"A0",X"16",X"8C",X"17",X"6D",X"18",
		X"46",X"19",X"1A",X"1A",X"E4",X"1A",X"A6",X"1B",X"63",X"1C",X"16",X"1D",X"C4",X"1D",X"6A",X"1E",
		X"0A",X"1F",X"A3",X"1F",X"37",X"20",X"C6",X"20",X"4E",X"21",X"CF",X"21",X"4C",X"22",X"C4",X"22",
		X"38",X"23",X"A4",X"23",X"0E",X"24",X"74",X"24",X"D4",X"24",X"30",X"25",X"87",X"25",X"DA",X"25",
		X"2A",X"26",X"74",X"26",X"BF",X"26",X"02",X"27",X"44",X"27",X"80",X"27",X"BC",X"27",X"F3",X"27",
		X"26",X"28",X"58",X"28",X"87",X"28",X"B2",X"28",X"DA",X"28",X"01",X"29",X"24",X"29",X"47",X"29",
		X"65",X"29",X"81",X"29",X"9C",X"29",X"B5",X"29",X"CB",X"29",X"DE",X"29",X"F0",X"29",X"01",X"2A",
		X"10",X"2A",X"1D",X"2A",X"26",X"2A",X"31",X"2A",X"3B",X"2A",X"40",X"2A",X"45",X"2A",X"48",X"2A",
		X"4A",X"2A",X"49",X"2A",X"4A",X"2A",X"48",X"2A",X"44",X"2A",X"3F",X"2A",X"3C",X"2A",X"34",X"2A",
		X"2D",X"2A",X"24",X"2A",X"19",X"2A",X"0F",X"2A",X"04",X"2A",X"F7",X"29",X"EA",X"29",X"DC",X"29",
		X"CC",X"29",X"BC",X"29",X"AD",X"29",X"9B",X"29",X"89",X"29",X"77",X"29",X"63",X"29",X"50",X"29",
		X"3C",X"29",X"27",X"29",X"10",X"29",X"FB",X"28",X"E3",X"28",X"CC",X"28",X"B4",X"28",X"9C",X"28",
		X"84",X"28",X"69",X"28",X"50",X"28",X"36",X"28",X"1D",X"28",X"01",X"28",X"E7",X"27",X"CC",X"27",
		X"B0",X"27",X"93",X"27",X"77",X"27",X"5B",X"27",X"3F",X"27",X"21",X"27",X"06",X"27",X"E6",X"26",
		X"C9",X"26",X"AA",X"26",X"8D",X"26",X"6D",X"26",X"51",X"26",X"31",X"26",X"13",X"26",X"F2",X"25",
		X"D5",X"25",X"B2",X"25",X"99",X"25",X"6F",X"25",X"5B",X"25",X"22",X"24",X"35",X"21",X"4F",X"1D",
		X"B8",X"18",X"C2",X"13",X"90",X"0E",X"4D",X"09",X"05",X"04",X"CB",X"FE",X"A6",X"F9",X"A1",X"F4",
		X"BA",X"EF",X"F5",X"EA",X"56",X"E6",X"DC",X"E1",X"85",X"DD",X"53",X"D9",X"45",X"D5",X"5A",X"D1",
		X"91",X"CD",X"E8",X"C9",X"60",X"C6",X"F8",X"C2",X"B0",X"BF",X"82",X"BC",X"75",X"B9",X"7C",X"B6",
		X"E3",X"B3",X"0E",X"B3",X"B1",X"B3",X"44",X"B5",X"78",X"B7",X"10",X"BA",X"E6",X"BC",X"DD",X"BF",
		X"E5",X"C2",X"EF",X"C5",X"F6",X"C8",X"ED",X"CB",X"D9",X"CE",X"B0",X"D1",X"77",X"D4",X"2A",X"D7",
		X"CA",X"D9",X"53",X"DC",X"CC",X"DE",X"2C",X"E1",X"7E",X"E3",X"BB",X"E5",X"E6",X"E7",X"FE",X"E9",
		X"08",X"EC",X"FE",X"ED",X"E5",X"EF",X"BA",X"F1",X"84",X"F3",X"3B",X"F5",X"E5",X"F6",X"80",X"F8",
		X"10",X"FA",X"91",X"FB",X"06",X"FD",X"6E",X"FE",X"C8",X"FF",X"18",X"01",X"5D",X"02",X"96",X"03",
		X"C5",X"04",X"E9",X"05",X"04",X"07",X"15",X"08",X"1D",X"09",X"1A",X"0A",X"10",X"0B",X"FC",X"0B",
		X"E2",X"0C",X"BD",X"0D",X"91",X"0E",X"5F",X"0F",X"25",X"10",X"E2",X"10",X"9C",X"11",X"2B",X"12",
		X"27",X"11",X"A3",X"0E",X"3B",X"0B",X"37",X"07",X"DC",X"02",X"51",X"FE",X"B0",X"F9",X"0E",X"F5",
		X"77",X"F0",X"F3",X"EB",X"8B",X"E7",X"3E",X"E3",X"10",X"DF",X"03",X"DB",X"15",X"D7",X"4A",X"D3",
		X"9C",X"CF",X"11",X"CC",X"A0",X"C8",X"53",X"C5",X"1E",X"C2",X"0B",X"BF",X"0D",X"BC",X"33",X"B9",
		X"69",X"B6",X"C7",X"B3",X"24",X"B1",X"55",X"AF",X"64",X"AF",X"A8",X"B0",X"C5",X"B2",X"68",X"B5",
		X"61",X"B8",X"8A",X"BB",X"CD",X"BE",X"1A",X"C2",X"61",X"C5",X"A4",X"C8",X"D2",X"CB",X"F6",X"CE",
		X"FB",X"D1",X"FC",X"D4",X"C0",X"D7",X"3C",X"DA",X"00",X"DD",X"A3",X"DF",X"38",X"E2",X"B1",X"E4",
		X"1D",X"E7",X"70",X"E9",X"B3",X"EB",X"E0",X"ED",X"FE",X"EF",X"08",X"F2",X"03",X"F4",X"EA",X"F5",
		X"C4",X"F7",X"8F",X"F9",X"49",X"FB",X"F4",X"FC",X"92",X"FE",X"22",X"00",X"A2",X"01",X"17",X"03",
		X"80",X"04",X"DE",X"05",X"2C",X"07",X"73",X"08",X"AA",X"09",X"DA",X"0A",X"FE",X"0B",X"1A",X"0D",
		X"28",X"0E",X"31",X"0F",X"2C",X"10",X"22",X"11",X"0E",X"12",X"F1",X"12",X"CD",X"13",X"A0",X"14",
		X"6A",X"15",X"2F",X"16",X"EC",X"16",X"A1",X"17",X"50",X"18",X"F9",X"18",X"98",X"19",X"35",X"1A",
		X"CC",X"1A",X"5C",X"1B",X"E4",X"1B",X"69",X"1C",X"EA",X"1C",X"64",X"1D",X"D9",X"1D",X"4A",X"1E",
		X"B4",X"1E",X"1C",X"1F",X"7F",X"1F",X"DC",X"1F",X"39",X"20",X"8E",X"20",X"E1",X"20",X"2F",X"21",
		X"7A",X"21",X"C3",X"21",X"05",X"22",X"47",X"22",X"83",X"22",X"BD",X"22",X"F5",X"22",X"29",X"23",
		X"5B",X"23",X"8A",X"23",X"B7",X"23",X"DF",X"23",X"07",X"24",X"2A",X"24",X"4E",X"24",X"6D",X"24",
		X"8C",X"24",X"A8",X"24",X"C2",X"24",X"D8",X"24",X"EF",X"24",X"03",X"25",X"15",X"25",X"25",X"25",
		X"34",X"25",X"3F",X"25",X"4D",X"25",X"55",X"25",X"60",X"25",X"66",X"25",X"6C",X"25",X"6D",X"25",
		X"7B",X"25",X"29",X"25",X"1D",X"23",X"BD",X"1F",X"86",X"1B",X"CB",X"16",X"C3",X"11",X"95",X"0C",
		X"58",X"07",X"23",X"02",X"00",X"FD",X"F5",X"F7",X"07",X"F3",X"3C",X"EE",X"95",X"E9",X"13",X"E5",
		X"B1",X"E0",X"77",X"DC",X"5E",X"D8",X"6B",X"D4",X"97",X"D0",X"E8",X"CC",X"55",X"C9",X"E7",X"C5",
		X"92",X"C2",X"63",X"BF",X"44",X"BC",X"51",X"B9",X"66",X"B6",X"9D",X"B4",X"AF",X"B4",X"E0",X"B5",
		X"E2",X"B7",X"5A",X"BA",X"2A",X"BD",X"24",X"C0",X"37",X"C3",X"51",X"C6",X"6D",X"C9",X"7C",X"CC",
		X"7E",X"CF",X"70",X"D2",X"4E",X"D5",X"18",X"D8",X"D0",X"DA",X"72",X"DD",X"FE",X"DF",X"78",X"E2",
		X"DE",X"E4",X"30",X"E7",X"70",X"E9",X"9B",X"EB",X"B6",X"ED",X"BF",X"EF",X"B7",X"F1",X"A5",X"F3",
		X"4A",X"F5",X"43",X"F5",X"BD",X"F3",X"49",X"F1",X"38",X"EE",X"CB",X"EA",X"23",X"E7",X"63",X"E3",
		X"9A",X"DF",X"D8",X"DB",X"22",X"D8",X"80",X"D4",X"F6",X"D0",X"83",X"CD",X"29",X"CA",X"EC",X"C6",
		X"CB",X"C3",X"C1",X"C0",X"D6",X"BD",X"04",X"BB",X"4E",X"B8",X"AC",X"B5",X"25",X"B3",X"B2",X"B0",
		X"5B",X"AE",X"14",X"AC",X"EE",X"A9",X"C5",X"A7",X"84",X"A6",X"26",X"A7",X"EC",X"A8",X"8D",X"AB",
		X"A6",X"AE",X"15",X"B2",X"AA",X"B5",X"5B",X"B9",X"0D",X"BD",X"BC",X"C0",X"59",X"C4",X"E9",X"C7",
		X"61",X"CB",X"C4",X"CE",X"0E",X"D2",X"42",X"D5",X"59",X"D8",X"5D",X"DB",X"45",X"DE",X"18",X"E1",
		X"D4",X"E3",X"7A",X"E6",X"09",X"E9",X"84",X"EB",X"E7",X"ED",X"3A",X"F0",X"79",X"F2",X"A5",X"F4",
		X"BE",X"F6",X"C5",X"F8",X"BB",X"FA",X"A1",X"FC",X"78",X"FE",X"3C",X"00",X"F2",X"01",X"9B",X"03",
		X"34",X"05",X"BF",X"06",X"3D",X"08",X"AE",X"09",X"14",X"0B",X"6D",X"0C",X"BA",X"0D",X"FA",X"0E",
		X"30",X"10",X"5A",X"11",X"7B",X"12",X"8F",X"13",X"9D",X"14",X"A0",X"15",X"9A",X"16",X"88",X"17",
		X"73",X"18",X"4E",X"19",X"20",X"1A",X"8D",X"19",X"52",X"17",X"24",X"14",X"49",X"10",X"0A",X"0C",
		X"94",X"07",X"04",X"03",X"6D",X"FE",X"E2",X"F9",X"67",X"F5",X"05",X"F1",X"BF",X"EC",X"95",X"E8",
		X"8C",X"E4",X"A2",X"E0",X"D8",X"DC",X"2E",X"D9",X"A2",X"D5",X"37",X"D2",X"E8",X"CE",X"B8",X"CB",
		X"A4",X"C8",X"A8",X"C5",X"CD",X"C2",X"05",X"C0",X"60",X"BD",X"C0",X"BA",X"B4",X"B8",X"81",X"B8",
		X"A7",X"B9",X"B5",X"BB",X"54",X"BE",X"51",X"C1",X"82",X"C4",X"D3",X"C7",X"2A",X"CB",X"83",X"CE",
		X"D1",X"D1",X"13",X"D5",X"3E",X"D8",X"5A",X"DB",X"5E",X"DE",X"4F",X"E1",X"25",X"E4",X"E9",X"E6",
		X"96",X"E9",X"2C",X"EC",X"AD",X"EE",X"1B",X"F1",X"73",X"F3",X"BA",X"F5",X"EA",X"F7",X"0E",X"FA",
		X"13",X"FC",X"17",X"FE",X"DF",X"FE",X"E0",X"FD",X"D6",X"FB",X"0B",X"F9",X"D3",X"F5",X"53",X"F2",
		X"B2",X"EE",X"FF",X"EA",X"50",X"E7",X"A6",X"E3",X"12",X"E0",X"8F",X"DC",X"26",X"D9",X"D3",X"D5",
		X"9E",X"D2",X"7E",X"CF",X"7B",X"CC",X"96",X"C9",X"C6",X"C6",X"12",X"C4",X"73",X"C1",X"ED",X"BE",
		X"7D",X"BC",X"29",X"BA",X"E3",X"B7",X"B9",X"B5",X"99",X"B3",X"DC",X"B1",X"E4",X"B1",X"5A",X"B3",
		X"BC",X"B5",X"B7",X"B8",X"0F",X"BC",X"A1",X"BF",X"4E",X"C3",X"04",X"C7",X"B7",X"CA",X"60",X"CE",
		X"F8",X"D1",X"79",X"D5",X"E7",X"D8",X"3B",X"DC",X"76",X"DF",X"9A",X"E2",X"A5",X"E5",X"97",X"E8",
		X"72",X"EB",X"34",X"EE",X"E3",X"F0",X"76",X"F3",X"F9",X"F5",X"60",X"F8",X"BE",X"FA",X"F9",X"FC",
		X"38",X"FF",X"68",X"00",X"C5",X"FF",X"07",X"FE",X"79",X"FB",X"78",X"F8",X"26",X"F5",X"B0",X"F1",
		X"22",X"EE",X"96",X"EA",X"0E",X"E7",X"9A",X"E3",X"35",X"E0",X"E8",X"DC",X"B1",X"D9",X"97",X"D6",
		X"90",X"D3",X"A7",X"D0",X"D5",X"CD",X"1D",X"CB",X"7C",X"C8",X"F3",X"C5",X"82",X"C3",X"25",X"C1",
		X"DF",X"BE",X"AF",X"BC",X"92",X"BA",X"8B",X"B8",X"95",X"B6",X"B2",X"B4",X"E2",X"B2",X"23",X"B1",
		X"76",X"AF",X"D9",X"AD",X"4D",X"AC",X"D0",X"AA",X"62",X"A9",X"01",X"A8",X"B1",X"A6",X"6E",X"A5",
		X"39",X"A4",X"0E",X"A3",X"F3",X"A1",X"E1",X"A0",X"DE",X"9F",X"E3",X"9E",X"F7",X"9D",X"10",X"9D",
		X"3B",X"9C",X"69",X"9B",X"A7",X"9A",X"E7",X"99",X"38",X"99",X"87",X"98",X"F0",X"97",X"46",X"97",
		X"6B",X"97",X"61",X"99",X"7E",X"9C",X"66",X"A0",X"C3",X"A4",X"6C",X"A9",X"34",X"AE",X"0B",X"B3",
		X"DC",X"B7",X"A0",X"BC",X"4B",X"C1",X"DF",X"C5",X"53",X"CA",X"AB",X"CE",X"E1",X"D2",X"F7",X"D6",
		X"EB",X"DA",X"C4",X"DE",X"7A",X"E2",X"15",X"E6",X"8F",X"E9",X"F1",X"EC",X"32",X"F0",X"5B",X"F3",
		X"67",X"F6",X"5B",X"F9",X"35",X"FC",X"F8",X"FE",X"A1",X"01",X"37",X"04",X"B4",X"06",X"1E",X"09",
		X"71",X"0B",X"B3",X"0D",X"DD",X"0F",X"F7",X"11",X"FB",X"13",X"F3",X"15",X"D4",X"17",X"AB",X"19",
		X"69",X"1B",X"22",X"1D",X"BD",X"1E",X"69",X"20",X"37",X"22",X"AE",X"23",X"20",X"25",X"7F",X"26",
		X"D5",X"27",X"1B",X"29",X"59",X"2A",X"89",X"2B",X"AE",X"2C",X"C8",X"2D",X"D7",X"2E",X"DC",X"2F",
		X"D6",X"30",X"C7",X"31",X"B0",X"32",X"8C",X"33",X"63",X"34",X"30",X"35",X"F5",X"35",X"B3",X"36",
		X"66",X"37",X"15",X"38",X"BB",X"38",X"59",X"39",X"F1",X"39",X"82",X"3A",X"0E",X"3B",X"93",X"3B",
		X"11",X"3C",X"88",X"3C",X"FD",X"3C",X"6A",X"3D",X"D3",X"3D",X"34",X"3E",X"94",X"3E",X"EA",X"3E",
		X"42",X"3F",X"8C",X"3F",X"D9",X"3F",X"DA",X"3E",X"27",X"3C",X"7A",X"38",X"1A",X"34",X"5D",X"2F",
		X"61",X"2A",X"54",X"25",X"3D",X"20",X"36",X"1B",X"41",X"16",X"67",X"11",X"AB",X"0C",X"12",X"08",
		X"98",X"03",X"44",X"FF",X"10",X"FB",X"00",X"F7",X"11",X"F3",X"45",X"EF",X"95",X"EB",X"09",X"E8",
		X"99",X"E4",X"48",X"E1",X"13",X"DE",X"FD",X"DA",X"00",X"D8",X"20",X"D5",X"56",X"D2",X"A7",X"CF",
		X"11",X"CD",X"90",X"CA",X"28",X"C8",X"D9",X"C5",X"99",X"C3",X"72",X"C1",X"5F",X"BF",X"5E",X"BD",
		X"72",X"BB",X"97",X"B9",X"CF",X"B7",X"15",X"B6",X"70",X"B4",X"D8",X"B2",X"53",X"B1",X"DB",X"AF",
		X"74",X"AE",X"16",X"AD",X"CD",X"AB",X"8B",X"AA",X"5C",X"A9",X"33",X"A8",X"1F",X"A7",X"0C",X"A6",
		X"12",X"A5",X"0F",X"A4",X"2F",X"A4",X"19",X"A6",X"14",X"A9",X"D0",X"AC",X"F7",X"B0",X"67",X"B5",
		X"F3",X"B9",X"8F",X"BE",X"21",X"C3",X"A8",X"C7",X"18",X"CC",X"70",X"D0",X"AA",X"D4",X"C8",X"D8",
		X"C5",X"DC",X"A7",X"E0",X"6A",X"E4",X"0E",X"E8",X"94",X"EB",X"FB",X"EE",X"49",X"F2",X"7C",X"F5",
		X"92",X"F8",X"90",X"FB",X"74",X"FE",X"3C",X"01",X"F5",X"03",X"5B",X"06",X"00",X"07",X"22",X"06",
		X"53",X"04",X"DC",X"01",X"05",X"FF",X"ED",X"FB",X"B8",X"F8",X"75",X"F5",X"34",X"F2",X"F9",X"EE",
		X"CE",X"EB",X"B4",X"E8",X"B1",X"E5",X"C3",X"E2",X"EC",X"DF",X"2B",X"DD",X"83",X"DA",X"F2",X"D7",
		X"74",X"D5",X"0F",X"D3",X"BD",X"D0",X"84",X"CE",X"5A",X"CC",X"4A",X"CA",X"46",X"C8",X"60",X"C6",
		X"75",X"C4",X"7C",X"C3",X"62",X"C4",X"6E",X"C6",X"4F",X"C9",X"A7",X"CC",X"52",X"D0",X"22",X"D4",
		X"0A",X"D8",X"EF",X"DB",X"D1",X"DF",X"A0",X"E3",X"5B",X"E7",X"FD",X"EA",X"8B",X"EE",X"F9",X"F1",
		X"53",X"F5",X"8E",X"F8",X"B2",X"FB",X"BB",X"FE",X"A9",X"01",X"7F",X"04",X"3E",X"07",X"E7",X"09",
		X"78",X"0C",X"F1",X"0E",X"57",X"11",X"A6",X"13",X"E3",X"15",X"0C",X"18",X"21",X"1A",X"24",X"1C",
		X"15",X"1E",X"F3",X"1F",X"C3",X"21",X"81",X"23",X"30",X"25",X"CE",X"26",X"5E",X"28",X"E1",X"29",
		X"54",X"2B",X"BC",X"2C",X"14",X"2E",X"61",X"2F",X"A0",X"30",X"D5",X"31",X"FD",X"32",X"1A",X"34",
		X"2D",X"35",X"35",X"36",X"31",X"37",X"26",X"38",X"0D",X"39",X"F0",X"39",X"C4",X"3A",X"8A",X"3B",
		X"E0",X"3A",X"8E",X"38",X"47",X"35",X"50",X"31",X"FD",X"2C",X"6B",X"28",X"C4",X"23",X"14",X"1F",
		X"6E",X"1A",X"D9",X"15",X"5E",X"11",X"FC",X"0C",X"BB",X"08",X"99",X"04",X"96",X"00",X"B2",X"FC",
		X"EF",X"F8",X"4C",X"F5",X"C6",X"F1",X"61",X"EE",X"14",X"EB",X"E8",X"E7",X"D3",X"E4",X"E0",X"E1",
		X"FE",X"DE",X"42",X"DC",X"89",X"D9",X"6B",X"D7",X"31",X"D7",X"4D",X"D8",X"4F",X"DA",X"E3",X"DC",
		X"D7",X"DF",X"FD",X"E2",X"42",X"E6",X"8F",X"E9",X"DC",X"EC",X"1F",X"F0",X"53",X"F3",X"75",X"F6",
		X"83",X"F9",X"7A",X"FC",X"5B",X"FF",X"24",X"02",X"DA",X"04",X"77",X"07",X"FF",X"09",X"71",X"0C",
		X"D1",X"0E",X"19",X"11",X"4E",X"13",X"71",X"15",X"81",X"17",X"7E",X"19",X"6A",X"1B",X"45",X"1D",
		X"0D",X"1F",X"C8",X"20",X"72",X"22",X"0F",X"24",X"9A",X"25",X"19",X"27",X"88",X"28",X"EC",X"29",
		X"43",X"2B",X"8C",X"2C",X"C9",X"2D",X"FC",X"2E",X"21",X"30",X"3C",X"31",X"4A",X"32",X"51",X"33",
		X"4D",X"34",X"3E",X"35",X"26",X"36",X"06",X"37",X"DC",X"37",X"A9",X"38",X"6E",X"39",X"2B",X"3A",
		X"DF",X"3A",X"8D",X"3B",X"30",X"3C",X"D2",X"3C",X"67",X"3D",X"F8",X"3D",X"83",X"3E",X"08",X"3F",
		X"84",X"3F",X"FD",X"3F",X"6F",X"40",X"DB",X"40",X"43",X"41",X"A5",X"41",X"01",X"42",X"58",X"42",
		X"AB",X"42",X"FB",X"42",X"44",X"43",X"8C",X"43",X"CC",X"43",X"09",X"44",X"41",X"44",X"79",X"44",
		X"A8",X"44",X"DA",X"44",X"FF",X"44",X"2E",X"45",X"49",X"45",X"78",X"45",X"9E",X"44",X"FC",X"41",
		X"4D",X"3E",X"DF",X"39",X"0A",X"35",X"F0",X"2F",X"C2",X"2A",X"8A",X"25",X"5F",X"20",X"45",X"1B",
		X"49",X"16",X"69",X"11",X"AC",X"0C",X"12",X"08",X"9C",X"03",X"47",X"FF",X"19",X"FB",X"0A",X"F7",
		X"1E",X"F3",X"55",X"EF",X"AB",X"EB",X"20",X"E8",X"B5",X"E4",X"67",X"E1",X"38",X"DE",X"23",X"DB",
		X"2A",X"D8",X"4C",X"D5",X"87",X"D2",X"DB",X"CF",X"47",X"CD",X"CA",X"CA",X"65",X"C8",X"15",X"C6",
		X"DA",X"C3",X"B5",X"C1",X"A4",X"BF",X"A6",X"BD",X"BA",X"BB",X"E2",X"B9",X"1B",X"B8",X"65",X"B6",
		X"C1",X"B4",X"2C",X"B3",X"A6",X"B1",X"2F",X"B0",X"C8",X"AE",X"6F",X"AD",X"25",X"AC",X"E8",X"AA",
		X"B7",X"A9",X"92",X"A8",X"79",X"A7",X"6E",X"A6",X"6F",X"A5",X"78",X"A4",X"8C",X"A3",X"AE",X"A2",
		X"D8",X"A1",X"0D",X"A1",X"47",X"A0",X"90",X"9F",X"E0",X"9E",X"36",X"9E",X"96",X"9D",X"01",X"9D",
		X"71",X"9C",X"E8",X"9B",X"68",X"9B",X"EE",X"9A",X"7E",X"9A",X"10",X"9A",X"AB",X"99",X"4D",X"99",
		X"F3",X"98",X"A0",X"98",X"54",X"98",X"0C",X"98",X"C9",X"97",X"8B",X"97",X"56",X"97",X"21",X"97",
		X"F3",X"96",X"C6",X"96",X"A3",X"96",X"80",X"96",X"65",X"96",X"4C",X"96",X"35",X"96",X"23",X"96",
		X"17",X"96",X"0C",X"96",X"05",X"96",X"00",X"96",X"01",X"96",X"02",X"96",X"09",X"96",X"10",X"96",
		X"1C",X"96",X"29",X"96",X"3A",X"96",X"4B",X"96",X"62",X"96",X"78",X"96",X"93",X"96",X"AE",X"96",
		X"D0",X"96",X"EA",X"96",X"14",X"97",X"29",X"97",X"DB",X"97",X"5F",X"9A",X"17",X"9E",X"A0",X"A2",
		X"A0",X"A7",X"EB",X"AC",X"54",X"B2",X"C8",X"B7",X"34",X"BD",X"8F",X"C2",X"CB",X"C7",X"ED",X"CC",
		X"E7",X"D1",X"C6",X"D6",X"76",X"DB",X"11",X"E0",X"6B",X"E4",X"85",X"E8",X"BB",X"EC",X"C9",X"F0",
		X"B8",X"F4",X"84",X"F8",X"31",X"FC",X"BF",X"FF",X"2D",X"03",X"82",X"06",X"B3",X"09",X"CB",X"0C",
		X"77",X"0E",X"58",X"0E",X"2D",X"0D",X"37",X"0B",X"D1",X"08",X"18",X"06",X"3E",X"03",X"46",X"00",
		X"50",X"FD",X"56",X"FA",X"6B",X"F7",X"8D",X"F4",X"C3",X"F1",X"09",X"EF",X"66",X"EC",X"D5",X"E9",
		X"5C",X"E7",X"F6",X"E4",X"A7",X"E2",X"68",X"E0",X"42",X"DE",X"29",X"DC",X"27",X"DA",X"37",X"D8",
		X"59",X"D6",X"8B",X"D4",X"CE",X"D2",X"1F",X"D1",X"83",X"CF",X"F5",X"CD",X"77",X"CC",X"05",X"CB",
		X"A2",X"C9",X"4D",X"C8",X"06",X"C7",X"CA",X"C5",X"9B",X"C4",X"76",X"C3",X"5D",X"C2",X"51",X"C1",
		X"4F",X"C0",X"5A",X"BF",X"6A",X"BE",X"87",X"BD",X"AC",X"BC",X"DD",X"BB",X"15",X"BB",X"57",X"BA",
		X"9F",X"B9",X"F3",X"B8",X"4A",X"B8",X"B0",X"B7",X"12",X"B7",X"8A",X"B6",X"F7",X"B5",X"8D",X"B6",
		X"EC",X"B8",X"56",X"BC",X"7F",X"C0",X"0E",X"C5",X"E4",X"C9",X"D1",X"CE",X"C7",X"D3",X"B4",X"D8",
		X"94",X"DD",X"57",X"E2",X"00",X"E7",X"85",X"EB",X"EE",X"EF",X"32",X"F4",X"57",X"F8",X"59",X"FC",
		X"3B",X"00",X"FC",X"03",X"9E",X"07",X"21",X"0B",X"88",X"0E",X"D0",X"11",X"FE",X"14",X"0D",X"18",
		X"04",X"1B",X"DF",X"1D",X"A3",X"20",X"4E",X"23",X"E1",X"25",X"5D",X"28",X"C3",X"2A",X"14",X"2D",
		X"4E",X"2F",X"77",X"31",X"8A",X"33",X"8A",X"35",X"77",X"37",X"54",X"39",X"1F",X"3B",X"D9",X"3C",
		X"82",X"3E",X"1C",X"40",X"A6",X"41",X"21",X"43",X"8F",X"44",X"EF",X"45",X"40",X"47",X"84",X"48",
		X"BA",X"49",X"E8",X"4A",X"05",X"4C",X"1B",X"4D",X"22",X"4E",X"22",X"4F",X"14",X"50",X"FE",X"50",
		X"D9",X"51",X"B1",X"52",X"7D",X"53",X"3F",X"54",X"FA",X"54",X"AA",X"55",X"55",X"56",X"F5",X"56",
		X"90",X"57",X"21",X"58",X"AC",X"58",X"31",X"59",X"AE",X"59",X"23",X"5A",X"95",X"5A",X"FE",X"5A",
		X"63",X"5B",X"C0",X"5B",X"19",X"5C",X"6C",X"5C",X"BB",X"5C",X"02",X"5D",X"47",X"5D",X"85",X"5D",
		X"C1",X"5D",X"F6",X"5D",X"29",X"5E",X"55",X"5E",X"7F",X"5E",X"A5",X"5E",X"C7",X"5E",X"E2",X"5E",
		X"FF",X"5E",X"13",X"5F",X"29",X"5F",X"39",X"5F",X"45",X"5F",X"4F",X"5F",X"56",X"5F",X"5A",X"5F",
		X"5D",X"5F",X"5A",X"5F",X"5A",X"5F",X"50",X"5F",X"48",X"5F",X"3B",X"5F",X"32",X"5F",X"1E",X"5F",
		X"12",X"5F",X"FA",X"5E",X"EB",X"5E",X"CA",X"5E",X"C4",X"5E",X"FE",X"5D",X"69",X"5B",X"A1",X"57",
		X"10",X"53",X"09",X"4E",X"B8",X"48",X"4E",X"43",X"D7",X"3D",X"69",X"38",X"10",X"33",X"D3",X"2D",
		X"B4",X"28",X"B8",X"23",X"E0",X"1E",X"2B",X"1A",X"9D",X"15",X"32",X"11",X"EC",X"0C",X"C9",X"08",
		X"C7",X"04",X"E8",X"00",X"2B",X"FD",X"8E",X"F9",X"0C",X"F6",X"AD",X"F2",X"66",X"EF",X"41",X"EC",
		X"3E",X"E9",X"BF",X"E7",X"01",X"E8",X"4A",X"E9",X"55",X"EB",X"CD",X"ED",X"95",X"F0",X"80",X"F3",
		X"84",X"F6",X"88",X"F9",X"8B",X"FC",X"82",X"FF",X"6C",X"02",X"42",X"05",X"05",X"08",X"B5",X"0A",
		X"4F",X"0D",X"D5",X"0F",X"45",X"12",X"A2",X"14",X"E8",X"16",X"1E",X"19",X"3E",X"1B",X"4E",X"1D",
		X"47",X"1F",X"35",X"21",X"09",X"23",X"D5",X"24",X"4D",X"25",X"FE",X"23",X"A6",X"21",X"8C",X"1E",
		X"09",X"1B",X"3C",X"17",X"51",X"13",X"55",X"0F",X"5F",X"0B",X"6F",X"07",X"95",X"03",X"D1",X"FF",
		X"25",X"FC",X"94",X"F8",X"1E",X"F5",X"C2",X"F1",X"83",X"EE",X"5E",X"EB",X"54",X"E8",X"65",X"E5",
		X"8E",X"E2",X"D2",X"DF",X"2A",X"DD",X"A0",X"DA",X"27",X"D8",X"CC",X"D5",X"75",X"D3",X"93",X"D1",
		X"89",X"D1",X"ED",X"D2",X"3B",X"D5",X"24",X"D8",X"6B",X"DB",X"EC",X"DE",X"86",X"E2",X"2B",X"E6",
		X"CD",X"E9",X"64",X"ED",X"E9",X"F0",X"59",X"F4",X"B3",X"F7",X"F7",X"FA",X"1E",X"FE",X"2F",X"01",
		X"27",X"04",X"06",X"07",X"CD",X"09",X"7D",X"0C",X"16",X"0F",X"99",X"11",X"04",X"14",X"5D",X"16",
		X"A0",X"18",X"D0",X"1A",X"EC",X"1C",X"F4",X"1E",X"EB",X"20",X"D2",X"22",X"A6",X"24",X"69",X"26",
		X"1C",X"28",X"C1",X"29",X"55",X"2B",X"DE",X"2C",X"52",X"2E",X"BE",X"2F",X"1B",X"31",X"6B",X"32",
		X"AE",X"33",X"E5",X"34",X"0F",X"36",X"31",X"37",X"42",X"38",X"4F",X"39",X"4D",X"3A",X"44",X"3B",
		X"2D",X"3C",X"11",X"3D",X"E9",X"3D",X"BA",X"3E",X"7F",X"3F",X"44",X"40",X"C8",X"40",X"9B",X"3F",
		X"EF",X"3C",X"5F",X"39",X"30",X"35",X"AB",X"30",X"F2",X"2B",X"28",X"27",X"5A",X"22",X"9A",X"1D",
		X"EB",X"18",X"58",X"14",X"E1",X"0F",X"8C",X"0B",X"53",X"07",X"3D",X"03",X"46",X"FF",X"72",X"FB",
		X"BB",X"F7",X"26",X"F4",X"AD",X"F0",X"53",X"ED",X"17",X"EA",X"F5",X"E6",X"F0",X"E3",X"06",X"E1",
		X"35",X"DE",X"7A",X"DB",X"DB",X"D8",X"53",X"D6",X"E1",X"D3",X"87",X"D1",X"3F",X"CF",X"10",X"CD",
		X"F2",X"CA",X"E9",X"C8",X"F2",X"C6",X"0E",X"C5",X"3C",X"C3",X"7B",X"C1",X"CB",X"BF",X"2C",X"BE",
		X"9B",X"BC",X"19",X"BB",X"A8",X"B9",X"46",X"B8",X"F0",X"B6",X"A8",X"B5",X"6E",X"B4",X"3D",X"B3",
		X"1D",X"B2",X"05",X"B1",X"FB",X"AF",X"FA",X"AE",X"05",X"AE",X"32",X"AD",X"F0",X"AD",X"4B",X"B0",
		X"97",X"B3",X"8E",X"B7",X"E0",X"BB",X"70",X"C0",X"14",X"C5",X"C0",X"C9",X"63",X"CE",X"F5",X"D2",
		X"70",X"D7",X"CF",X"DB",X"0F",X"E0",X"33",X"E4",X"38",X"E8",X"1B",X"EC",X"E2",X"EF",X"88",X"F3",
		X"11",X"F7",X"7B",X"FA",X"CC",X"FD",X"FD",X"00",X"16",X"04",X"10",X"07",X"FA",X"09",X"BC",X"0C",
		X"7E",X"0F",X"83",X"11",X"9C",X"11",X"6E",X"10",X"5A",X"0E",X"BD",X"0B",X"C3",X"08",X"98",X"05",
		X"51",X"02",X"05",X"FF",X"B9",X"FB",X"78",X"F8",X"47",X"F5",X"28",X"F2",X"1F",X"EF",X"2C",X"EC",
		X"52",X"E9",X"8D",X"E6",X"E1",X"E3",X"4B",X"E1",X"CC",X"DE",X"60",X"DC",X"0D",X"DA",X"CB",X"D7",
		X"A2",X"D5",X"88",X"D3",X"85",X"D1",X"91",X"CF",X"B3",X"CD",X"E2",X"CB",X"26",X"CA",X"76",X"C8",
		X"DC",X"C6",X"4B",X"C5",X"D0",X"C3",X"5C",X"C2",X"FE",X"C0",X"A5",X"BF",X"61",X"BE",X"23",X"BD",
		X"FA",X"BB",X"D1",X"BA",X"C3",X"B9",X"AD",X"B8",X"C1",X"B7",X"95",X"B6",X"0C",X"B5",X"37",X"B4",
		X"54",X"B3",X"8B",X"B2",X"C0",X"B1",X"05",X"B1",X"4D",X"B0",X"A2",X"AF",X"FD",X"AE",X"61",X"AE",
		X"CB",X"AD",X"3D",X"AD",X"B7",X"AC",X"37",X"AC",X"BC",X"AB",X"4A",X"AB",X"DF",X"AA",X"77",X"AA",
		X"19",X"AA",X"BC",X"A9",X"69",X"A9",X"17",X"A9",X"CF",X"A8",X"87",X"A8",X"48",X"A8",X"0A",X"A8",
		X"D5",X"A7",X"A0",X"A7",X"74",X"A7",X"46",X"A7",X"23",X"A7",X"FE",X"A6",X"E2",X"A6",X"C4",X"A6",
		X"B2",X"A6",X"98",X"A6",X"8E",X"A6",X"76",X"A6",X"91",X"A7",X"71",X"AA",X"5C",X"AE",X"00",X"B3",
		X"09",X"B8",X"53",X"BD",X"B3",X"C2",X"17",X"C8",X"70",X"CD",X"B6",X"D2",X"DC",X"D7",X"E6",X"DC",
		X"CC",X"E1",X"8E",X"E6",X"2B",X"EB",X"A7",X"EF",X"FC",X"F3",X"2F",X"F8",X"3F",X"FC",X"2C",X"00",
		X"FA",X"03",X"A5",X"07",X"35",X"0B",X"A3",X"0E",X"F5",X"11",X"28",X"15",X"4A",X"18",X"04",X"1B",
		X"E9",X"1B",X"48",X"1B",X"B2",X"19",X"71",X"17",X"CD",X"14",X"E7",X"11",X"DF",X"0E",X"C9",X"0B",
		X"B2",X"08",X"A0",X"05",X"9C",X"02",X"A7",X"FF",X"C7",X"FC",X"FA",X"F9",X"42",X"F7",X"9F",X"F4",
		X"14",X"F2",X"9B",X"EF",X"39",X"ED",X"EB",X"EA",X"B1",X"E8",X"88",X"E6",X"75",X"E4",X"75",X"E2",
		X"86",X"E0",X"A8",X"DE",X"DB",X"DC",X"20",X"DB",X"74",X"D9",X"D6",X"D7",X"49",X"D6",X"C9",X"D4",
		X"59",X"D3",X"F6",X"D1",X"A1",X"D0",X"55",X"CF",X"1A",X"CE",X"E9",X"CC",X"C3",X"CB",X"AA",X"CA",
		X"9C",X"C9",X"99",X"C8",X"9F",X"C7",X"B0",X"C6",X"C9",X"C5",X"ED",X"C4",X"1A",X"C4",X"50",X"C3",
		X"8E",X"C2",X"D6",X"C1",X"24",X"C1",X"7A",X"C0",X"D9",X"BF",X"3E",X"BF",X"AB",X"BE",X"1F",X"BE",
		X"98",X"BD",X"1A",X"BD",X"A1",X"BC",X"2F",X"BC",X"C1",X"BB",X"58",X"BB",X"F7",X"BA",X"9B",X"BA",
		X"43",X"BA",X"F1",X"B9",X"A3",X"B9",X"5C",X"B9",X"15",X"B9",X"D5",X"B8",X"9B",X"B8",X"64",X"B8",
		X"2F",X"B8",X"00",X"B8",X"D4",X"B7",X"AD",X"B7",X"88",X"B7",X"67",X"B7",X"48",X"B7",X"2F",X"B7",
		X"17",X"B7",X"03",X"B7",X"F2",X"B6",X"E1",X"B6",X"D6",X"B6",X"CC",X"B6",X"C5",X"B6",X"C0",X"B6",
		X"BE",X"B6",X"BE",X"B6",X"C1",X"B6",X"C6",X"B6",X"CC",X"B6",X"D4",X"B6",X"DF",X"B6",X"EB",X"B6",
		X"FB",X"B6",X"0A",X"B7",X"1C",X"B7",X"2E",X"B7",X"44",X"B7",X"5A",X"B7",X"71",X"B7",X"8A",X"B7",
		X"A5",X"B7",X"BF",X"B7",X"DF",X"B7",X"FC",X"B7",X"1D",X"B8",X"4D",X"B8",X"EE",X"B9",X"37",X"BD",
		X"71",X"C1",X"56",X"C6",X"91",X"CB",X"05",X"D1",X"86",X"D6",X"0C",X"DC",X"7E",X"E1",X"DC",X"E6",
		X"19",X"EC",X"37",X"F1",X"2C",X"F6",X"02",X"FB",X"AB",X"FF",X"36",X"04",X"97",X"08",X"D8",X"0C",
		X"F2",X"10",X"EB",X"14",X"C1",X"18",X"77",X"1C",X"0A",X"20",X"81",X"23",X"D7",X"26",X"13",X"2A",
		X"31",X"2D",X"33",X"30",X"1A",X"33",X"E8",X"35",X"9C",X"38",X"37",X"3B",X"BA",X"3D",X"28",X"40",
		X"7E",X"42",X"BF",X"44",X"EA",X"46",X"01",X"49",X"05",X"4B",X"F6",X"4C",X"D3",X"4E",X"9F",X"50",
		X"5A",X"52",X"05",X"54",X"9C",X"55",X"26",X"57",X"A1",X"58",X"0A",X"5A",X"68",X"5B",X"B6",X"5C",
		X"F8",X"5D",X"29",X"5F",X"54",X"60",X"69",X"61",X"7A",X"62",X"3A",X"62",X"34",X"60",X"26",X"5D",
		X"59",X"59",X"23",X"55",X"A9",X"50",X"13",X"4C",X"70",X"47",X"D7",X"42",X"49",X"3E",X"D3",X"39",
		X"77",X"35",X"38",X"31",X"14",X"2D",X"12",X"29",X"2F",X"25",X"67",X"21",X"C1",X"1D",X"34",X"1A",
		X"CA",X"16",X"77",X"13",X"46",X"10",X"27",X"0D",X"2D",X"0A",X"3F",X"07",X"7A",X"04",X"BA",X"01",
		X"2D",X"00",X"80",X"00",X"F3",X"01",X"37",X"04",X"F4",X"06",X"04",X"0A",X"3C",X"0D",X"8C",X"10",
		X"DC",X"13",X"2B",X"17",X"6B",X"1A",X"9C",X"1D",X"B8",X"20",X"BE",X"23",X"AC",X"26",X"83",X"29",
		X"42",X"2C",X"EB",X"2E",X"7C",X"31",X"F9",X"33",X"5D",X"36",X"AC",X"38",X"E6",X"3A",X"09",X"3D",
		X"1E",X"3F",X"19",X"41",X"0C",X"43",X"AC",X"44",X"8C",X"44",X"E0",X"42",X"47",X"40",X"09",X"3D",
		X"69",X"39",X"92",X"35",X"9D",X"31",X"A0",X"2D",X"A7",X"29",X"BC",X"25",X"E2",X"21",X"20",X"1E",
		X"77",X"1A",X"E7",X"16",X"72",X"13",X"1A",X"10",X"DB",X"0C",X"B8",X"09",X"AB",X"06",X"BC",X"03",
		X"E3",X"00",X"25",X"FE",X"7A",X"FB",X"EE",X"F8",X"6A",X"F6",X"0F",X"F4",X"AC",X"F1",X"48",X"F0",
		X"CC",X"F0",X"7D",X"F2",X"09",X"F5",X"14",X"F8",X"74",X"FB",X"FC",X"FE",X"9B",X"02",X"3C",X"06",
		X"DA",X"09",X"65",X"0D",X"E2",X"10",X"46",X"14",X"94",X"17",X"C7",X"1A",X"E3",X"1D",X"E3",X"20",
		X"CD",X"23",X"9D",X"26",X"54",X"29",X"F3",X"2B",X"7B",X"2E",X"EA",X"30",X"48",X"33",X"8E",X"35",
		X"C1",X"37",X"DF",X"39",X"CE",X"3B",X"17",X"3C",X"BE",X"3A",X"67",X"38",X"61",X"35",X"F5",X"31",
		X"48",X"2E",X"7D",X"2A",X"A4",X"26",X"CD",X"22",X"02",X"1F",X"48",X"1B",X"A3",X"17",X"17",X"14",
		X"A3",X"10",X"48",X"0D",X"08",X"0A",X"E4",X"06",X"D6",X"03",X"E3",X"00",X"0A",X"FE",X"47",X"FB",
		X"9F",X"F8",X"09",X"F6",X"8F",X"F3",X"23",X"F1",X"D8",X"EE",X"89",X"EC",X"02",X"EB",X"65",X"EB",
		X"0C",X"ED",X"96",X"EF",X"A5",X"F2",X"0D",X"F6",X"A3",X"F9",X"53",X"FD",X"05",X"01",X"B3",X"04",
		X"53",X"08",X"E2",X"0B",X"57",X"0F",X"B8",X"12",X"FD",X"15",X"2A",X"19",X"39",X"1C",X"34",X"1F",
		X"13",X"22",X"DB",X"24",X"8A",X"27",X"20",X"2A",X"A0",X"2C",X"0A",X"2F",X"5E",X"31",X"9B",X"33",
		X"C8",X"35",X"DD",X"37",X"E1",X"39",X"D1",X"3B",X"B0",X"3D",X"7D",X"3F",X"39",X"41",X"E5",X"42",
		X"80",X"44",X"0A",X"46",X"88",X"47",X"F7",X"48",X"57",X"4A",X"A8",X"4B",X"EE",X"4C",X"25",X"4E",
		X"50",X"4F",X"6F",X"50",X"85",X"51",X"8C",X"52",X"8B",X"53",X"7A",X"54",X"66",X"55",X"41",X"56",
		X"16",X"57",X"DF",X"57",X"A3",X"58",X"5A",X"59",X"0E",X"5A",X"B3",X"5A",X"57",X"5B",X"E9",X"5B",
		X"7F",X"5C",X"04",X"5D",X"8B",X"5D",X"03",X"5E",X"7A",X"5E",X"E3",X"5E",X"52",X"5F",X"AC",X"5F",
		X"10",X"60",X"5C",X"60",X"B9",X"60",X"F6",X"60",X"50",X"61",X"75",X"61",X"FD",X"61",X"01",X"63",
		X"23",X"63",X"5C",X"63",X"82",X"63",X"AB",X"63",X"CC",X"63",X"E9",X"63",X"09",X"64",X"1B",X"64",
		X"35",X"64",X"12",X"63",X"27",X"60",X"35",X"5C",X"87",X"57",X"73",X"52",X"20",X"4D",X"B8",X"47",
		X"49",X"42",X"E7",X"3C",X"97",X"37",X"68",X"32",X"54",X"2D",X"66",X"28",X"9B",X"23",X"F4",X"1E",
		X"72",X"1A",X"13",X"16",X"D9",X"11",X"C0",X"0D",X"CC",X"09",X"F5",X"05",X"43",X"02",X"AB",X"FE",
		X"38",X"FB",X"DE",X"F7",X"A7",X"F4",X"7C",X"F1",X"C3",X"EE",X"E4",X"ED",X"90",X"EE",X"2E",X"F0",
		X"76",X"F2",X"22",X"F5",X"11",X"F8",X"1E",X"FB",X"3D",X"FE",X"5B",X"01",X"74",X"04",X"80",X"07",
		X"7D",X"0A",X"61",X"0D",X"36",X"10",X"F2",X"12",X"9C",X"15",X"2B",X"18",X"A9",X"1A",X"0F",X"1D",
		X"62",X"1F",X"9F",X"21",X"CB",X"23",X"DF",X"25",X"E6",X"27",X"D6",X"29",X"B6",X"2B",X"85",X"2D",
		X"45",X"2F",X"F3",X"30",X"91",X"32",X"20",X"34",X"A1",X"35",X"12",X"37",X"79",X"38",X"CE",X"39",
		X"1A",X"3B",X"56",X"3C",X"89",X"3D",X"AC",X"3E",X"C6",X"3F",X"D4",X"40",X"DB",X"41",X"D2",X"42",
		X"C2",X"43",X"A6",X"44",X"82",X"45",X"55",X"46",X"1D",X"47",X"DF",X"47",X"97",X"48",X"48",X"49",
		X"F1",X"49",X"8F",X"4A",X"2D",X"4B",X"95",X"4B",X"50",X"4A",X"7C",X"47",X"BB",X"43",X"57",X"3F",
		X"9B",X"3A",X"A9",X"35",X"A4",X"30",X"9B",X"2B",X"A3",X"26",X"BC",X"21",X"F2",X"1C",X"43",X"18",
		X"BB",X"13",X"4E",X"0F",X"08",X"0B",X"E1",X"06",X"DD",X"02",X"F8",X"FE",X"37",X"FB",X"94",X"F7",
		X"10",X"F4",X"A9",X"F0",X"61",X"ED",X"34",X"EA",X"26",X"E7",X"2F",X"E4",X"54",X"E1",X"90",X"DE",
		X"E9",X"DB",X"54",X"D9",X"DB",X"D6",X"74",X"D4",X"28",X"D2",X"EB",X"CF",X"C8",X"CD",X"B5",X"CB",
		X"B7",X"C9",X"CA",X"C7",X"F0",X"C5",X"28",X"C4",X"70",X"C2",X"C9",X"C0",X"32",X"BF",X"AA",X"BD",
		X"31",X"BC",X"C7",X"BA",X"6A",X"B9",X"1D",X"B8",X"DB",X"B6",X"A8",X"B5",X"7D",X"B4",X"65",X"B3",
		X"50",X"B2",X"4D",X"B1",X"63",X"B0",X"05",X"B1",X"53",X"B3",X"9F",X"B6",X"9A",X"BA",X"F7",X"BE",
		X"91",X"C3",X"44",X"C8",X"00",X"CD",X"B1",X"D1",X"53",X"D6",X"DC",X"DA",X"4B",X"DF",X"9A",X"E3",
		X"CB",X"E7",X"DD",X"EB",X"CD",X"EF",X"A1",X"F3",X"53",X"F7",X"E9",X"FA",X"5D",X"FE",X"B8",X"01",
		X"F3",X"04",X"18",X"08",X"1B",X"0B",X"0B",X"0E",X"D9",X"10",X"A1",X"13",X"BB",X"15",X"E2",X"15",
		X"B0",X"14",X"94",X"12",X"E6",X"0F",X"DA",X"0C",X"9C",X"09",X"3E",X"06",X"DA",X"02",X"75",X"FF",
		X"1F",X"FC",X"D6",X"F8",X"A2",X"F5",X"81",X"F2",X"7B",X"EF",X"8A",X"EC",X"B3",X"E9",X"F0",X"E6",
		X"48",X"E4",X"B3",X"E1",X"38",X"DF",X"D0",X"DC",X"80",X"DA",X"40",X"D8",X"1C",X"D6",X"02",X"D4",
		X"06",X"D2",X"16",X"D0",X"8B",X"CF",X"CC",X"D0",X"1C",X"D3",X"2F",X"D6",X"AD",X"D9",X"7A",X"DD",
		X"64",X"E1",X"61",X"E5",X"5B",X"E9",X"4A",X"ED",X"25",X"F1",X"F0",X"F4",X"9E",X"F8",X"35",X"FC",
		X"AD",X"FF",X"0B",X"03",X"51",X"06",X"7A",X"09",X"88",X"0C",X"7D",X"0F",X"5A",X"12",X"1B",X"15",
		X"CA",X"17",X"5A",X"1A",X"DD",X"1C",X"3D",X"1F",X"9C",X"21",X"7A",X"23",X"78",X"23",X"05",X"22",
		X"A3",X"1F",X"A6",X"1C",X"4B",X"19",X"B6",X"15",X"0B",X"12",X"52",X"0E",X"9D",X"0A",X"F6",X"06",
		X"62",X"03",X"E0",X"FF",X"7A",X"FC",X"29",X"F9",X"F4",X"F5",X"D5",X"F2",X"D3",X"EF",X"E9",X"EC",
		X"19",X"EA",X"60",X"E7",X"C1",X"E4",X"35",X"E2",X"C3",X"DF",X"63",X"DD",X"20",X"DB",X"E2",X"D8",
		X"03",X"D7",X"EF",X"D6",X"64",X"D8",X"CC",X"DA",X"D9",X"DD",X"47",X"E1",X"F3",X"E4",X"B9",X"E8",
		X"8B",X"EC",X"57",X"F0",X"1B",X"F4",X"C8",X"F7",X"63",X"FB",X"E4",X"FE",X"4D",X"02",X"9A",X"05",
		X"D0",X"08",X"E9",X"0B",X"EA",X"0E",X"CF",X"11",X"9F",X"14",X"54",X"17",X"F4",X"19",X"7C",X"1C",
		X"ED",X"1E",X"49",X"21",X"91",X"23",X"C3",X"25",X"E4",X"27",X"EE",X"29",X"E8",X"2B",X"CE",X"2D",
		X"A5",X"2F",X"68",X"31",X"1D",X"33",X"C1",X"34",X"56",X"36",X"DC",X"37",X"54",X"39",X"BC",X"3A",
		X"18",X"3C",X"66",X"3D",X"AA",X"3E",X"DD",X"3F",X"06",X"41",X"23",X"42",X"36",X"43",X"3D",X"44",
		X"39",X"45",X"2B",X"46",X"13",X"47",X"F0",X"47",X"C5",X"48",X"91",X"49",X"56",X"4A",X"0F",X"4B",
		X"C1",X"4B",X"6C",X"4C",X"0D",X"4D",X"AA",X"4D",X"3D",X"4E",X"C9",X"4E",X"4F",X"4F",X"CD",X"4F",
		X"46",X"50",X"B8",X"50",X"23",X"51",X"89",X"51",X"EB",X"51",X"45",X"52",X"9C",X"52",X"EC",X"52",
		X"38",X"53",X"7F",X"53",X"C0",X"53",X"FE",X"53",X"37",X"54",X"6D",X"54",X"9E",X"54",X"C9",X"54",
		X"F3",X"54",X"18",X"55",X"3A",X"55",X"58",X"55",X"73",X"55",X"8A",X"55",X"9D",X"55",X"AF",X"55",
		X"BD",X"55",X"CA",X"55",X"D0",X"55",X"D7",X"55",X"DB",X"55",X"DB",X"55",X"DA",X"55",X"D5",X"55",
		X"CF",X"55",X"C6",X"55",X"BC",X"55",X"B0",X"55",X"A0",X"55",X"90",X"55",X"7E",X"55",X"6A",X"55",
		X"52",X"55",X"3C",X"55",X"23",X"55",X"09",X"55",X"EB",X"54",X"CD",X"54",X"AF",X"54",X"8F",X"54",
		X"6C",X"54",X"4A",X"54",X"25",X"54",X"00",X"54",X"D9",X"53",X"B3",X"53",X"89",X"53",X"60",X"53",
		X"33",X"53",X"08",X"53",X"DC",X"52",X"B0",X"52",X"80",X"52",X"53",X"52",X"24",X"52",X"F1",X"51",
		X"C1",X"51",X"8E",X"51",X"5B",X"51",X"27",X"51",X"F6",X"50",X"C1",X"50",X"8C",X"50",X"57",X"50",
		X"1F",X"50",X"EA",X"4F",X"B4",X"4F",X"7B",X"4F",X"44",X"4F",X"0C",X"4F",X"D3",X"4E",X"9A",X"4E",
		X"60",X"4E",X"27",X"4E",X"ED",X"4D",X"B3",X"4D",X"78",X"4D",X"3C",X"4D",X"04",X"4D",X"C7",X"4C",
		X"8B",X"4C",X"51",X"4C",X"14",X"4C",X"D7",X"4B",X"9C",X"4B",X"60",X"4B",X"22",X"4B",X"E6",X"4A",
		X"A9",X"4A",X"6C",X"4A",X"2F",X"4A",X"F2",X"49",X"B4",X"49",X"77",X"49",X"3B",X"49",X"FC",X"48",
		X"BE",X"48",X"81",X"48",X"43",X"48",X"06",X"48",X"C8",X"47",X"89",X"47",X"4D",X"47",X"0D",X"47",
		X"D0",X"46",X"93",X"46",X"54",X"46",X"18",X"46",X"D9",X"45",X"9D",X"45",X"5E",X"45",X"20",X"45",
		X"E3",X"44",X"A6",X"44",X"68",X"44",X"2A",X"44",X"EC",X"43",X"B0",X"43",X"72",X"43",X"35",X"43",
		X"F8",X"42",X"BC",X"42",X"7F",X"42",X"40",X"42",X"05",X"42",X"C8",X"41",X"8B",X"41",X"4D",X"41",
		X"13",X"41",X"D6",X"40",X"9B",X"40",X"5D",X"40",X"22",X"40",X"E5",X"3F",X"AA",X"3F",X"6F",X"3F",
		X"33",X"3F",X"F7",X"3E",X"BC",X"3E",X"81",X"3E",X"46",X"3E",X"0C",X"3E",X"CF",X"3D",X"97",X"3D",
		X"59",X"3D",X"21",X"3D",X"E4",X"3C",X"AD",X"3C",X"6D",X"3C",X"94",X"3B",X"D1",X"38",X"91",X"34",
		X"B1",X"2F",X"51",X"2A",X"C2",X"24",X"0E",X"1F",X"60",X"19",X"B9",X"13",X"2D",X"0E",X"BC",X"08",
		X"71",X"03",X"49",X"FE",X"4A",X"F9",X"6E",X"F4",X"BC",X"EF",X"30",X"EB",X"CB",X"E6",X"87",X"E2",
		X"6B",X"DE",X"72",X"DA",X"9D",X"D6",X"E7",X"D2",X"56",X"CF",X"DF",X"CB",X"8D",X"C8",X"50",X"C5",
		X"64",X"C2",X"46",X"C1",X"CA",X"C1",X"50",X"C3",X"8B",X"C5",X"30",X"C8",X"1E",X"CB",X"2F",X"CE",
		X"55",X"D1",X"7A",X"D4",X"A1",X"D7",X"B5",X"DA",X"C0",X"DD",X"B2",X"E0",X"96",X"E3",X"62",X"E6",
		X"1B",X"E9",X"BE",X"EB",X"4C",X"EE",X"C4",X"F0",X"2A",X"F3",X"7A",X"F5",X"B9",X"F7",X"E1",X"F9",
		X"FC",X"FB",X"02",X"FE",X"F7",X"FF",X"DB",X"01",X"B0",X"03",X"73",X"05",X"2A",X"07",X"CF",X"08",
		X"67",X"0A",X"F1",X"0B",X"6D",X"0D",X"DC",X"0E",X"40",X"10",X"96",X"11",X"DF",X"12",X"1D",X"14",
		X"52",X"15",X"78",X"16",X"98",X"17",X"AA",X"18",X"B4",X"19",X"B4",X"1A",X"A9",X"1B",X"96",X"1C",
		X"7B",X"1D",X"57",X"1E",X"2A",X"1F",X"F7",X"1F",X"B8",X"20",X"77",X"21",X"2B",X"22",X"C3",X"22",
		X"CB",X"21",X"27",X"1F",X"8D",X"1B",X"42",X"17",X"9D",X"12",X"BC",X"0D",X"C7",X"08",X"CB",X"03",
		X"E1",X"FE",X"06",X"FA",X"48",X"F5",X"A6",X"F0",X"27",X"EC",X"C9",X"E7",X"8E",X"E3",X"75",X"DF",
		X"7F",X"DB",X"A9",X"D7",X"F6",X"D3",X"62",X"D0",X"EE",X"CC",X"97",X"C9",X"5F",X"C6",X"44",X"C3",
		X"47",X"C0",X"62",X"BD",X"99",X"BA",X"E8",X"B7",X"51",X"B5",X"D2",X"B2",X"6B",X"B0",X"19",X"AE",
		X"DF",X"AB",X"BB",X"A9",X"A9",X"A7",X"AC",X"A5",X"C3",X"A3",X"EC",X"A1",X"28",X"A0",X"75",X"9E",
		X"D4",X"9C",X"44",X"9B",X"C4",X"99",X"52",X"98",X"F1",X"96",X"9E",X"95",X"58",X"94",X"20",X"93",
		X"F7",X"91",X"D9",X"90",X"CA",X"8F",X"C6",X"8E",X"CD",X"8D",X"E0",X"8C",X"FE",X"8B",X"28",X"8B",
		X"5B",X"8A",X"98",X"89",X"E0",X"88",X"30",X"88",X"8B",X"87",X"ED",X"86",X"58",X"86",X"CA",X"85",
		X"46",X"85",X"CA",X"84",X"54",X"84",X"E7",X"83",X"81",X"83",X"20",X"83",X"C6",X"82",X"75",X"82",
		X"28",X"82",X"E2",X"81",X"A1",X"81",X"66",X"81",X"31",X"81",X"01",X"81",X"D5",X"80",X"AF",X"80",
		X"8F",X"80",X"72",X"80",X"5B",X"80",X"46",X"80",X"38",X"80",X"2D",X"80",X"22",X"80",X"20",X"80",
		X"21",X"80",X"24",X"80",X"2C",X"80",X"35",X"80",X"44",X"80",X"54",X"80",X"67",X"80",X"7E",X"80",
		X"97",X"80",X"B3",X"80",X"D2",X"80",X"F3",X"80",X"18",X"81",X"3C",X"81",X"68",X"81",X"90",X"81",
		X"C0",X"81",X"EA",X"81",X"1F",X"82",X"4C",X"82",X"89",X"82",X"B5",X"82",X"0F",X"84",X"3B",X"87",
		X"73",X"8B",X"6D",X"90",X"CA",X"95",X"6C",X"9B",X"21",X"A1",X"DD",X"A6",X"89",X"AC",X"22",X"B2",
		X"99",X"B7",X"F4",X"BC",X"27",X"C2",X"38",X"C7",X"21",X"CC",X"E4",X"D0",X"81",X"D5",X"FB",X"D9",
		X"4F",X"DE",X"81",X"E2",X"90",X"E6",X"7C",X"EA",X"49",X"EE",X"F6",X"F1",X"82",X"F5",X"F3",X"F8",
		X"45",X"FC",X"7B",X"FF",X"96",X"02",X"96",X"05",X"7D",X"08",X"4B",X"0B",X"00",X"0E",X"9C",X"10",
		X"23",X"13",X"96",X"15",X"F2",X"17",X"37",X"1A",X"6A",X"1C",X"8A",X"1E",X"96",X"20",X"90",X"22",
		X"78",X"24",X"50",X"26",X"15",X"28",X"CA",X"29",X"71",X"2B",X"08",X"2D",X"8F",X"2E",X"07",X"30",
		X"74",X"31",X"D2",X"32",X"22",X"34",X"69",X"35",X"7D",X"36",X"DD",X"35",X"A2",X"33",X"72",X"30",
		X"95",X"2C",X"5B",X"28",X"E7",X"23",X"5A",X"1F",X"C6",X"1A",X"3D",X"16",X"C3",X"11",X"63",X"0D",
		X"1C",X"09",X"F4",X"04",X"E8",X"00",X"FD",X"FC",X"31",X"F9",X"86",X"F5",X"F6",X"F1",X"87",X"EE",
		X"33",X"EB",X"FD",X"E7",X"E3",X"E4",X"E4",X"E1",X"FE",X"DE",X"33",X"DC",X"81",X"D9",X"E6",X"D6",
		X"62",X"D4",X"F8",X"D1",X"A1",X"CF",X"60",X"CD",X"33",X"CB",X"1A",X"C9",X"17",X"C7",X"24",X"C5",
		X"43",X"C3",X"77",X"C1",X"BA",X"BF",X"0E",X"BE",X"73",X"BC",X"E6",X"BA",X"68",X"B9",X"FA",X"B7",
		X"9B",X"B6",X"47",X"B5",X"02",X"B4",X"CD",X"B2",X"A0",X"B1",X"83",X"B0",X"6E",X"AF",X"68",X"AE",
		X"6A",X"AD",X"79",X"AC",X"91",X"AB",X"B3",X"AA",X"E0",X"A9",X"17",X"A9",X"56",X"A8",X"9E",X"A7",
		X"EF",X"A6",X"48",X"A6",X"AA",X"A5",X"14",X"A5",X"85",X"A4",X"FD",X"A3",X"7C",X"A3",X"04",X"A3",
		X"8F",X"A2",X"24",X"A2",X"BD",X"A1",X"5D",X"A1",X"04",X"A1",X"B0",X"A0",X"60",X"A0",X"18",X"A0",
		X"D2",X"9F",X"95",X"9F",X"58",X"9F",X"26",X"9F",X"F1",X"9E",X"CB",X"9E",X"92",X"9E",X"F3",X"9E",
		X"36",X"A1",X"C6",X"A4",X"31",X"A9",X"1E",X"AE",X"5C",X"B3",X"C0",X"B8",X"2D",X"BE",X"97",X"C3",
		X"EF",X"C8",X"2E",X"CE",X"4C",X"D3",X"49",X"D8",X"24",X"DD",X"DB",X"E1",X"6D",X"E6",X"DA",X"EA",
		X"23",X"EF",X"4B",X"F3",X"4F",X"F7",X"33",X"FB",X"F4",X"FE",X"97",X"02",X"19",X"06",X"7F",X"09",
		X"C8",X"0C",X"F6",X"0F",X"04",X"13",X"FB",X"15",X"D7",X"18",X"9C",X"1B",X"45",X"1E",X"D9",X"20",
		X"56",X"23",X"BE",X"25",X"0C",X"28",X"4A",X"2A",X"70",X"2C",X"86",X"2E",X"87",X"30",X"75",X"32",
		X"52",X"34",X"20",X"36",X"D8",X"37",X"86",X"39",X"1F",X"3B",X"AB",X"3C",X"26",X"3E",X"96",X"3F",
		X"F6",X"40",X"4B",X"42",X"8D",X"43",X"CB",X"44",X"F1",X"45",X"1E",X"47",X"D8",X"47",X"BD",X"46",
		X"2E",X"44",X"B5",X"40",X"A8",X"3C",X"42",X"38",X"AA",X"33",X"FF",X"2E",X"51",X"2A",X"AD",X"25",
		X"1F",X"21",X"A7",X"1C",X"4B",X"18",X"0F",X"14",X"F0",X"0F",X"F3",X"0B",X"14",X"08",X"57",X"04",
		X"B7",X"00",X"2F",X"FD",X"C1",X"F9",X"73",X"F6",X"3F",X"F3",X"29",X"F0",X"2A",X"ED",X"49",X"EA",
		X"7E",X"E7",X"CF",X"E4",X"33",X"E2",X"B2",X"DF",X"47",X"DD",X"F0",X"DA",X"B0",X"D8",X"82",X"D6",
		X"6A",X"D4",X"66",X"D2",X"72",X"D0",X"91",X"CE",X"C1",X"CC",X"03",X"CB",X"56",X"C9",X"B7",X"C7",
		X"29",X"C6",X"A9",X"C4",X"37",X"C3",X"D5",X"C1",X"81",X"C0",X"37",X"BF",X"FC",X"BD",X"CF",X"BC",
		X"AA",X"BB",X"93",X"BA",X"87",X"B9",X"86",X"B8",X"90",X"B7",X"A6",X"B6",X"C3",X"B5",X"EB",X"B4",
		X"1D",X"B4",X"56",X"B3",X"9B",X"B2",X"E6",X"B1",X"3A",X"B1",X"96",X"B0",X"F9",X"AF",X"65",X"AF",
		X"D7",X"AE",X"51",X"AE",X"D3",X"AD",X"5A",X"AD",X"E8",X"AC",X"7C",X"AC",X"17",X"AC",X"B5",X"AB",
		X"5B",X"AB",X"05",X"AB",X"B7",X"AA",X"6B",X"AA",X"25",X"AA",X"E4",X"A9",X"A9",X"A9",X"71",X"A9",
		X"3E",X"A9",X"0F",X"A9",X"E5",X"A8",X"BD",X"A8",X"9B",X"A8",X"7C",X"A8",X"5F",X"A8",X"46",X"A8",
		X"33",X"A8",X"20",X"A8",X"12",X"A8",X"07",X"A8",X"FE",X"A7",X"F8",X"A7",X"F5",X"A7",X"F6",X"A7",
		X"F8",X"A7",X"FC",X"A7",X"06",X"A8",X"0E",X"A8",X"1A",X"A8",X"29",X"A8",X"39",X"A8",X"4B",X"A8",
		X"5F",X"A8",X"77",X"A8",X"8C",X"A8",X"A6",X"A8",X"DB",X"A8",X"A8",X"AA",X"18",X"AE",X"7C",X"B2",
		X"89",X"B7",X"F0",X"BC",X"8A",X"C2",X"36",X"C8",X"E2",X"CD",X"7C",X"D3",X"FF",X"D8",X"61",X"DE",
		X"A2",X"E3",X"BD",X"E8",X"B2",X"ED",X"83",X"F2",X"2A",X"F7",X"AE",X"FB",X"0A",X"00",X"45",X"04",
		X"59",X"08",X"51",X"0C",X"1F",X"10",X"D4",X"13",X"61",X"17",X"D9",X"1A",X"23",X"1E",X"6C",X"21",
		X"E8",X"23",X"62",X"24",X"83",X"23",X"B3",X"21",X"50",X"1F",X"89",X"1C",X"8D",X"19",X"71",X"16",
		X"4B",X"13",X"21",X"10",X"01",X"0D",X"F0",X"09",X"F1",X"06",X"02",X"04",X"2B",X"01",X"67",X"FE",
		X"BC",X"FB",X"25",X"F9",X"A4",X"F6",X"37",X"F4",X"E0",X"F1",X"9B",X"EF",X"6D",X"ED",X"4F",X"EB",
		X"47",X"E9",X"4B",X"E7",X"69",X"E5",X"99",X"E3",X"43",X"E3",X"BA",X"E4",X"3E",X"E7",X"84",X"EA",
		X"35",X"EE",X"31",X"F2",X"48",X"F6",X"72",X"FA",X"93",X"FE",X"AC",X"02",X"AD",X"06",X"9D",X"0A",
		X"6E",X"0E",X"27",X"12",X"BE",X"15",X"3D",X"19",X"9B",X"1C",X"E1",X"1F",X"09",X"23",X"16",X"26",
		X"09",X"29",X"E2",X"2B",X"9F",X"2E",X"48",X"31",X"D7",X"33",X"4F",X"36",X"B0",X"38",X"FB",X"3A",
		X"33",X"3D",X"55",X"3F",X"62",X"41",X"5E",X"43",X"46",X"45",X"1E",X"47",X"E2",X"48",X"94",X"4A",
		X"38",X"4C",X"CB",X"4D",X"4E",X"4F",X"C3",X"50",X"29",X"52",X"82",X"53",X"CB",X"54",X"08",X"56",
		X"38",X"57",X"5C",X"58",X"72",X"59",X"7E",X"5A",X"7E",X"5B",X"72",X"5C",X"5E",X"5D",X"3F",X"5E",
		X"14",X"5F",X"E1",X"5F",X"A3",X"60",X"5D",X"61",X"0E",X"62",X"B8",X"62",X"57",X"63",X"F0",X"63",
		X"81",X"64",X"0A",X"65",X"8B",X"65",X"05",X"66",X"79",X"66",X"E7",X"66",X"4C",X"67",X"AE",X"67",
		X"07",X"68",X"5E",X"68",X"A8",X"68",X"F5",X"68",X"37",X"69",X"78",X"69",X"B0",X"69",X"E7",X"69",
		X"16",X"6A",X"44",X"6A",X"69",X"6A",X"8F",X"6A",X"A9",X"6A",X"CE",X"6A",X"9E",X"6A",X"A3",X"68",
		X"2E",X"65",X"CE",X"60",X"DA",X"5B",X"8F",X"56",X"16",X"51",X"90",X"4B",X"09",X"46",X"98",X"40",
		X"3C",X"3B",X"FF",X"35",X"E3",X"30",X"ED",X"2B",X"19",X"27",X"6D",X"22",X"E1",X"1D",X"7E",X"19",
		X"3C",X"15",X"1F",X"11",X"22",X"0D",X"49",X"09",X"8F",X"05",X"F6",X"01",X"7B",X"FE",X"1F",X"FB",
		X"DA",X"F7",X"B8",X"F4",X"AC",X"F1",X"BF",X"EE",X"E8",X"EB",X"2D",X"E9",X"86",X"E6",X"FB",X"E3",
		X"83",X"E1",X"23",X"DF",X"D7",X"DC",X"A1",X"DA",X"7D",X"D8",X"6F",X"D6",X"71",X"D4",X"88",X"D2",
		X"AE",X"D0",X"E8",X"CE",X"30",X"CD",X"8A",X"CB",X"F3",X"C9",X"6C",X"C8",X"F2",X"C6",X"88",X"C5",
		X"2A",X"C4",X"DB",X"C2",X"98",X"C1",X"63",X"C0",X"35",X"BF",X"3D",X"BE",X"FA",X"BE",X"57",X"C1",
		X"AC",X"C4",X"AD",X"C8",X"09",X"CD",X"A7",X"D1",X"55",X"D6",X"0E",X"DB",X"BB",X"DF",X"59",X"E4",
		X"DC",X"E8",X"45",X"ED",X"8E",X"F1",X"BB",X"F5",X"C5",X"F9",X"B1",X"FD",X"7A",X"01",X"27",X"05",
		X"B4",X"08",X"24",X"0C",X"76",X"0F",X"AD",X"12",X"C6",X"15",X"C5",X"18",X"AB",X"1B",X"76",X"1E",
		X"17",X"21",X"18",X"22",X"55",X"21",X"88",X"1F",X"F8",X"1C",X"FC",X"19",X"B3",X"16",X"4A",X"13",
		X"CB",X"0F",X"4E",X"0C",X"D4",X"08",X"6D",X"05",X"14",X"02",X"D6",X"FE",X"A9",X"FB",X"9A",X"F8",
		X"9F",X"F5",X"BB",X"F2",X"F0",X"EF",X"3F",X"ED",X"A4",X"EA",X"1F",X"E8",X"AF",X"E5",X"56",X"E3",
		X"11",X"E1",X"E2",X"DE",X"C3",X"DC",X"BB",X"DA",X"C1",X"D8",X"DD",X"D6",X"09",X"D5",X"46",X"D3",
		X"93",X"D1",X"EF",X"CF",X"5C",X"CE",X"D9",X"CC",X"64",X"CB",X"FA",X"C9",X"9F",X"C8",X"53",X"C7",
		X"12",X"C6",X"DD",X"C4",X"B6",X"C3",X"99",X"C2",X"8B",X"C1",X"82",X"C0",X"88",X"BF",X"95",X"BE",
		X"B0",X"BD",X"D0",X"BC",X"FF",X"BB",X"31",X"BB",X"73",X"BA",X"B4",X"B9",X"09",X"B9",X"5E",X"B8",
		X"17",X"B9",X"99",X"BB",X"28",X"BF",X"72",X"C3",X"24",X"C8",X"18",X"CD",X"21",X"D2",X"36",X"D7",
		X"40",X"DC",X"37",X"E1",X"13",X"E6",X"D5",X"EA",X"74",X"EF",X"F2",X"F3",X"4D",X"F8",X"87",X"FC",
		X"9D",X"00",X"92",X"04",X"67",X"08",X"1A",X"0C",X"AE",X"0F",X"23",X"13",X"7F",X"16",X"B6",X"19",
		X"D7",X"1C",X"D5",X"1F",X"CC",X"22",X"3A",X"25",X"B7",X"25",X"B9",X"24",X"C3",X"22",X"2D",X"20",
		X"32",X"1D",X"FA",X"19",X"A2",X"16",X"3E",X"13",X"D8",X"0F",X"7F",X"0C",X"33",X"09",X"FB",X"05",
		X"D5",X"02",X"C9",X"FF",X"D1",X"FC",X"F4",X"F9",X"2B",X"F7",X"7B",X"F4",X"E0",X"F1",X"5E",X"EF",
		X"ED",X"EC",X"98",X"EA",X"4F",X"E8",X"22",X"E6",X"01",X"E4",X"FE",X"E1",X"FB",X"DF",X"31",X"DF",
		X"4D",X"E0",X"8E",X"E2",X"A0",X"E5",X"28",X"E9",X"01",X"ED",X"FD",X"F0",X"0B",X"F5",X"1B",X"F9",
		X"1E",X"FD",X"0E",X"01",X"EC",X"04",X"AF",X"08",X"58",X"0C",X"E7",X"0F",X"55",X"13",X"AD",X"16",
		X"DF",X"19",X"13",X"1D",X"5B",X"20",X"45",X"23",X"20",X"26",X"DB",X"28",X"81",X"2B",X"0E",X"2E",
		X"86",X"30",X"E6",X"32",X"31",X"35",X"68",X"37",X"89",X"39",X"95",X"3B",X"91",X"3D",X"79",X"3F",
		X"50",X"41",X"14",X"43",X"C9",X"44",X"6C",X"46",X"FE",X"47",X"83",X"49",X"F9",X"4A",X"5E",X"4C",
		X"B9",X"4D",X"03",X"4F",X"41",X"50",X"73",X"51",X"98",X"52",X"B1",X"53",X"BE",X"54",X"BF",X"55",
		X"B5",X"56",X"A3",X"57",X"84",X"58",X"5B",X"59",X"2B",X"5A",X"F1",X"5A",X"AC",X"5B",X"5F",X"5C",
		X"0A",X"5D",X"AD",X"5D",X"47",X"5E",X"DB",X"5E",X"65",X"5F",X"EA",X"5F",X"66",X"60",X"DD",X"60",
		X"4D",X"61",X"B7",X"61",X"19",X"62",X"75",X"62",X"CD",X"62",X"1F",X"63",X"6A",X"63",X"B2",X"63",
		X"F5",X"63",X"32",X"64",X"69",X"64",X"9B",X"64",X"CA",X"64",X"F5",X"64",X"1A",X"65",X"3F",X"65",
		X"5D",X"65",X"59",X"65",X"B1",X"63",X"64",X"60",X"1F",X"5C",X"32",X"57",X"EA",X"51",X"6C",X"4C",
		X"D9",X"46",X"48",X"41",X"C6",X"3B",X"5B",X"36",X"0E",X"31",X"E3",X"2B",X"DC",X"26",X"F8",X"21",
		X"3C",X"1D",X"A5",X"18",X"31",X"14",X"E3",X"0F",X"B7",X"0B",X"B2",X"07",X"C8",X"03",X"06",X"00",
		X"5F",X"FC",X"DE",X"F8",X"70",X"F5",X"2E",X"F2",X"EE",X"EE",X"87",X"EC",X"24",X"EC",X"19",X"ED",
		X"00",X"EF",X"79",X"F1",X"54",X"F4",X"63",X"F7",X"93",X"FA",X"CC",X"FD",X"06",X"01",X"36",X"04",
		X"58",X"07",X"65",X"0A",X"60",X"0D",X"46",X"10",X"15",X"13",X"CF",X"15",X"6F",X"18",X"FB",X"1A",
		X"71",X"1D",X"D1",X"1F",X"1B",X"22",X"54",X"24",X"78",X"26",X"88",X"28",X"87",X"2A",X"73",X"2C",
		X"4C",X"2E",X"17",X"30",X"CC",X"31",X"77",X"33",X"0F",X"35",X"99",X"36",X"13",X"38",X"81",X"39",
		X"DF",X"3A",X"33",X"3C",X"75",X"3D",X"AF",X"3E",X"DA",X"3F",X"FC",X"40",X"0F",X"42",X"1B",X"43",
		X"18",X"44",X"0F",X"45",X"F7",X"45",X"DB",X"46",X"B0",X"47",X"80",X"48",X"41",X"49",X"01",X"4A",
		X"B2",X"4A",X"64",X"4B",X"02",X"4C",X"AC",X"4C",X"C9",X"4C",X"FC",X"4A",X"CD",X"47",X"BA",X"43",
		X"1B",X"3F",X"27",X"3A",X"0A",X"35",X"DB",X"2F",X"B2",X"2A",X"96",X"25",X"91",X"20",X"A9",X"1B",
		X"E2",X"16",X"3A",X"12",X"B7",X"0D",X"57",X"09",X"1B",X"05",X"00",X"01",X"08",X"FD",X"30",X"F9",
		X"7B",X"F5",X"E2",X"F1",X"6C",X"EE",X"0E",X"EB",X"D5",X"E7",X"B0",X"E4",X"B2",X"E1",X"C0",X"DE",
		X"2C",X"DD",X"85",X"DD",X"03",X"DF",X"54",X"E1",X"22",X"E4",X"45",X"E7",X"91",X"EA",X"F5",X"ED",
		X"5E",X"F1",X"C2",X"F4",X"18",X"F8",X"60",X"FB",X"92",X"FE",X"AE",X"01",X"B2",X"04",X"A1",X"07",
		X"78",X"0A",X"37",X"0D",X"E1",X"0F",X"72",X"12",X"EF",X"14",X"54",X"17",X"A7",X"19",X"E3",X"1B",
		X"0D",X"1E",X"20",X"20",X"2D",X"22",X"D0",X"23",X"8F",X"23",X"CB",X"21",X"0B",X"1F",X"AD",X"1B",
		X"ED",X"17",X"F2",X"13",X"DF",X"0F",X"C1",X"0B",X"AA",X"07",X"A4",X"03",X"AF",X"FF",X"D5",X"FB",
		X"13",X"F8",X"70",X"F4",X"E4",X"F0",X"78",X"ED",X"27",X"EA",X"F4",X"E6",X"D8",X"E3",X"DB",X"E0",
		X"F5",X"DD",X"2D",X"DB",X"78",X"D8",X"E3",X"D5",X"58",X"D3",X"F6",X"D0",X"90",X"CE",X"4E",X"CD",
		X"04",X"CE",X"ED",X"CF",X"B1",X"D2",X"F3",X"D5",X"8A",X"D9",X"4D",X"DD",X"28",X"E1",X"01",X"E5",
		X"D6",X"E8",X"9A",X"EC",X"4E",X"F0",X"E7",X"F3",X"6B",X"F7",X"D0",X"FA",X"1F",X"FE",X"52",X"01",
		X"6C",X"04",X"6C",X"07",X"53",X"0A",X"20",X"0D",X"D6",X"0F",X"72",X"12",X"FC",X"14",X"6E",X"17",
		X"C9",X"19",X"15",X"1C",X"1C",X"1E",X"5C",X"1E",X"F5",X"1C",X"8E",X"1A",X"76",X"17",X"F6",X"13",
		X"36",X"10",X"57",X"0C",X"6C",X"08",X"83",X"04",X"A8",X"00",X"DF",X"FC",X"2D",X"F9",X"92",X"F5",
		X"13",X"F2",X"AC",X"EE",X"63",X"EB",X"33",X"E8",X"22",X"E5",X"27",X"E2",X"48",X"DF",X"7F",X"DC",
		X"D2",X"D9",X"3A",X"D7",X"BE",X"D4",X"4F",X"D2",X"05",X"D0",X"B5",X"CD",X"4F",X"CC",X"E8",X"CC",
		X"C3",X"CE",X"84",X"D1",X"C8",X"D4",X"67",X"D8",X"34",X"DC",X"17",X"E0",X"FE",X"E3",X"E0",X"E7",
		X"B2",X"EB",X"6F",X"EF",X"13",X"F3",X"A1",X"F6",X"12",X"FA",X"69",X"FD",X"A4",X"00",X"C5",X"03",
		X"CC",X"06",X"B9",X"09",X"8D",X"0C",X"4A",X"0F",X"EB",X"11",X"77",X"14",X"EB",X"16",X"4C",X"19",
		X"93",X"1B",X"C9",X"1D",X"EA",X"1F",X"F7",X"21",X"F0",X"23",X"D9",X"25",X"AE",X"27",X"73",X"29",
		X"27",X"2B",X"CB",X"2C",X"5F",X"2E",X"E4",X"2F",X"5A",X"31",X"C1",X"32",X"1A",X"34",X"67",X"35",
		X"A5",X"36",X"D8",X"37",X"FE",X"38",X"19",X"3A",X"27",X"3B",X"2A",X"3C",X"24",X"3D",X"12",X"3E",
		X"F6",X"3E",X"CF",X"3F",X"A0",X"40",X"69",X"41",X"27",X"42",X"DC",X"42",X"89",X"43",X"2D",X"44",
		X"CB",X"44",X"61",X"45",X"EF",X"45",X"76",X"46",X"F6",X"46",X"6F",X"47",X"E1",X"47",X"4E",X"48",
		X"B3",X"48",X"15",X"49",X"6E",X"49",X"C3",X"49",X"12",X"4A",X"5E",X"4A",X"A1",X"4A",X"E3",X"4A",
		X"1D",X"4B",X"55",X"4B",X"86",X"4B",X"B7",X"4B",X"DE",X"4B",X"08",X"4C",X"22",X"4C",X"4F",X"4C",
		X"03",X"4C",X"E1",X"49",X"63",X"46",X"07",X"42",X"21",X"3D",X"ED",X"37",X"90",X"32",X"27",X"2D",
		X"C2",X"27",X"6F",X"22",X"37",X"1D",X"1D",X"18",X"23",X"13",X"50",X"0E",X"9F",X"09",X"12",X"05",
		X"AA",X"00",X"68",X"FC",X"49",X"F8",X"4B",X"F4",X"72",X"F0",X"B8",X"EC",X"1D",X"E9",X"A2",X"E5",
		X"46",X"E2",X"07",X"DF",X"E4",X"DB",X"DD",X"D8",X"F2",X"D5",X"21",X"D3",X"67",X"D0",X"C9",X"CD",
		X"3E",X"CB",X"D0",X"C8",X"75",X"C6",X"30",X"C4",X"FF",X"C1",X"E3",X"BF",X"DB",X"BD",X"E8",X"BB",
		X"05",X"BA",X"36",X"B8",X"77",X"B6",X"CC",X"B4",X"2B",X"B3",X"A1",X"B1",X"22",X"B0",X"B4",X"AE",
		X"53",X"AD",X"03",X"AC",X"BC",X"AA",X"86",X"A9",X"59",X"A8",X"3F",X"A7",X"2A",X"A6",X"26",X"A5",
		X"27",X"A4",X"3A",X"A3",X"51",X"A2",X"7A",X"A1",X"A4",X"A0",X"E2",X"9F",X"1D",X"9F",X"6E",X"9E",
		X"BD",X"9D",X"1E",X"9D",X"7C",X"9C",X"EF",X"9B",X"5B",X"9B",X"DF",X"9A",X"58",X"9A",X"F1",X"99",
		X"6E",X"99",X"22",X"99",X"70",X"98",X"3B",X"97",X"F7",X"96",X"9C",X"96",X"55",X"96",X"0E",X"96",
		X"CB",X"95",X"95",X"95",X"50",X"95",X"01",X"96",X"8B",X"98",X"30",X"9C",X"A0",X"A0",X"79",X"A5",
		X"9D",X"AA",X"D8",X"AF",X"23",X"B5",X"60",X"BA",X"8A",X"BF",X"9B",X"C4",X"8D",X"C9",X"5F",X"CE",
		X"0D",X"D3",X"98",X"D7",X"01",X"DC",X"46",X"E0",X"67",X"E4",X"66",X"E8",X"44",X"EC",X"03",X"F0",
		X"A0",X"F3",X"21",X"F7",X"82",X"FA",X"C7",X"FD",X"ED",X"00",X"FB",X"03",X"EB",X"06",X"C5",X"09",
		X"81",X"0C",X"2B",X"0F",X"B9",X"11",X"33",X"14",X"94",X"16",X"E3",X"18",X"19",X"1B",X"3E",X"1D",
		X"4D",X"1F",X"4D",X"21",X"36",X"23",X"12",X"25",X"D8",X"26",X"92",X"28",X"38",X"2A",X"D2",X"2B",
		X"57",X"2D",X"D4",X"2E",X"3B",X"30",X"9B",X"31",X"E6",X"32",X"2E",X"34",X"5E",X"35",X"8F",X"36",
		X"A4",X"37",X"C7",X"38",X"23",X"39",X"A6",X"37",X"F4",X"34",X"6F",X"31",X"6E",X"2D",X"1D",X"29",
		X"A9",X"24",X"23",X"20",X"A2",X"1B",X"2B",X"17",X"CA",X"12",X"80",X"0E",X"55",X"0A",X"45",X"06",
		X"56",X"02",X"82",X"FE",X"D1",X"FA",X"3C",X"F7",X"C7",X"F3",X"6F",X"F0",X"32",X"ED",X"0F",X"EA",
		X"0D",X"E7",X"1F",X"E4",X"50",X"E1",X"94",X"DE",X"F8",X"DB",X"78",X"D9",X"79",X"D8",X"2B",X"D9",
		X"DF",X"DA",X"4C",X"DD",X"25",X"E0",X"45",X"E3",X"86",X"E6",X"DD",X"E9",X"30",X"ED",X"7F",X"F0",
		X"C1",X"F3",X"EF",X"F6",X"09",X"FA",X"10",X"FD",X"FD",X"FF",X"D2",X"02",X"93",X"05",X"39",X"08",
		X"CD",X"0A",X"47",X"0D",X"AE",X"0F",X"FD",X"11",X"3D",X"14",X"62",X"16",X"7A",X"18",X"75",X"1A",
		X"73",X"1C",X"DA",X"1D",X"6A",X"1D",X"AE",X"1B",X"13",X"19",X"F0",X"15",X"73",X"12",X"C9",X"0E",
		X"05",X"0B",X"41",X"07",X"7E",X"03",X"CC",X"FF",X"2E",X"FC",X"A5",X"F8",X"35",X"F5",X"DE",X"F1",
		X"A1",X"EE",X"81",X"EB",X"77",X"E8",X"89",X"E5",X"B3",X"E2",X"F8",X"DF",X"52",X"DD",X"C5",X"DA",
		X"4C",X"D8",X"EE",X"D5",X"A0",X"D3",X"70",X"D1",X"4A",X"CF",X"6A",X"CE",X"4C",X"CF",X"33",X"D1",
		X"DC",X"D3",X"EE",X"D6",X"4C",X"DA",X"CA",X"DD",X"5C",X"E1",X"ED",X"E4",X"78",X"E8",X"F0",X"EB",
		X"58",X"EF",X"A9",X"F2",X"E3",X"F5",X"03",X"F9",X"0C",X"FC",X"FD",X"FE",X"D5",X"01",X"96",X"04",
		X"3C",X"07",X"CF",X"09",X"49",X"0C",X"B0",X"0E",X"FE",X"10",X"3B",X"13",X"5F",X"15",X"7D",X"17",
		X"30",X"19",X"23",X"19",X"B2",X"17",X"5F",X"15",X"77",X"12",X"34",X"0F",X"BF",X"0B",X"2C",X"08",
		X"96",X"04",X"00",X"01",X"79",X"FD",X"02",X"FA",X"9F",X"F6",X"55",X"F3",X"23",X"F0",X"0A",X"ED",
		X"0A",X"EA",X"23",X"E7",X"53",X"E4",X"9D",X"E1",X"FE",X"DE",X"77",X"DC",X"04",X"DA",X"A9",X"D7",
		X"64",X"D5",X"30",X"D3",X"11",X"D1",X"08",X"CF",X"10",X"CD",X"2A",X"CB",X"55",X"C9",X"93",X"C7",
		X"E1",X"C5",X"40",X"C4",X"AD",X"C2",X"2C",X"C1",X"B7",X"BF",X"50",X"BE",X"F8",X"BC",X"AD",X"BB",
		X"6F",X"BA",X"40",X"B9",X"19",X"B8",X"FF",X"B6",X"F3",X"B5",X"F0",X"B4",X"F8",X"B3",X"0C",X"B3",
		X"27",X"B2",X"4E",X"B1",X"7F",X"B0",X"B9",X"AF",X"FC",X"AE",X"47",X"AE",X"9A",X"AD",X"F5",X"AC",
		X"58",X"AC",X"C3",X"AB",X"35",X"AB",X"AF",X"AA",X"2E",X"AA",X"B7",X"A9",X"43",X"A9",X"D8",X"A8",
		X"73",X"A8",X"12",X"A8",X"B9",X"A7",X"65",X"A7",X"14",X"A7",X"CA",X"A6",X"86",X"A6",X"45",X"A6",
		X"0A",X"A6",X"D2",X"A5",X"A0",X"A5",X"72",X"A5",X"48",X"A5",X"22",X"A5",X"01",X"A5",X"E3",X"A4",
		X"C7",X"A4",X"B0",X"A4",X"9D",X"A4",X"8C",X"A4",X"7E",X"A4",X"74",X"A4",X"6F",X"A4",X"6A",X"A4",
		X"68",X"A4",X"69",X"A4",X"6E",X"A4",X"73",X"A4",X"7C",X"A4",X"88",X"A4",X"96",X"A4",X"A5",X"A4",
		X"B8",X"A4",X"CB",X"A4",X"E0",X"A4",X"F8",X"A4",X"12",X"A5",X"2E",X"A5",X"4B",X"A5",X"6A",X"A5",
		X"8B",X"A5",X"AC",X"A5",X"D0",X"A5",X"F4",X"A5",X"1B",X"A6",X"45",X"A6",X"6C",X"A6",X"97",X"A6",
		X"C2",X"A6",X"EF",X"A6",X"1E",X"A7",X"4C",X"A7",X"7B",X"A7",X"AC",X"A7",X"DE",X"A7",X"11",X"A8",
		X"44",X"A8",X"7A",X"A8",X"AF",X"A8",X"E5",X"A8",X"1B",X"A9",X"52",X"A9",X"8B",X"A9",X"C4",X"A9",
		X"FE",X"A9",X"3A",X"AA",X"74",X"AA",X"B0",X"AA",X"EA",X"AA",X"27",X"AB",X"63",X"AB",X"A1",X"AB",
		X"E0",X"AB",X"1E",X"AC",X"5D",X"AC",X"9B",X"AC",X"DB",X"AC",X"1C",X"AD",X"5B",X"AD",X"9B",X"AD",
		X"DD",X"AD",X"1C",X"AE",X"5E",X"AE",X"9F",X"AE",X"E3",X"AE",X"25",X"AF",X"67",X"AF",X"AA",X"AF",
		X"EC",X"AF",X"2E",X"B0",X"71",X"B0",X"B4",X"B0",X"F8",X"B0",X"3B",X"B1",X"7F",X"B1",X"C2",X"B1",
		X"06",X"B2",X"49",X"B2",X"8E",X"B2",X"D1",X"B2",X"14",X"B3",X"5A",X"B3",X"9E",X"B3",X"E3",X"B3",
		X"27",X"B4",X"6B",X"B4",X"AE",X"B4",X"F2",X"B4",X"36",X"B5",X"7B",X"B5",X"BF",X"B5",X"02",X"B6",
		X"46",X"B6",X"8A",X"B6",X"CF",X"B6",X"13",X"B7",X"56",X"B7",X"9B",X"B7",X"DF",X"B7",X"22",X"B8",
		X"65",X"B8",X"AB",X"B8",X"ED",X"B8",X"30",X"B9",X"75",X"B9",X"B7",X"B9",X"FB",X"B9",X"3C",X"BA",
		X"7F",X"BA",X"C2",X"BA",X"06",X"BB",X"47",X"BB",X"8B",X"BB",X"CD",X"BB",X"10",X"BC",X"51",X"BC",
		X"94",X"BC",X"D6",X"BC",X"19",X"BD",X"59",X"BD",X"9B",X"BD",X"DA",X"BD",X"1C",X"BE",X"5E",X"BE",
		X"A0",X"BE",X"E0",X"BE",X"23",X"BF",X"61",X"BF",X"A2",X"BF",X"E2",X"BF",X"23",X"C0",X"62",X"C0",
		X"A4",X"C0",X"E1",X"C0",X"25",X"C1",X"5A",X"C1",X"D9",X"C1",X"E4",X"C3",X"34",X"C7",X"4B",X"CB",
		X"DF",X"CF",X"BD",X"D4",X"BE",X"D9",X"CA",X"DE",X"D0",X"E3",X"C5",X"E8",X"A1",X"ED",X"5F",X"F2",
		X"FD",X"F6",X"7A",X"FB",X"D4",X"FF",X"0D",X"04",X"22",X"08",X"16",X"0C",X"E8",X"0F",X"99",X"13",
		X"2A",X"17",X"9D",X"1A",X"F1",X"1D",X"28",X"21",X"43",X"24",X"41",X"27",X"24",X"2A",X"EE",X"2C",
		X"9E",X"2F",X"38",X"32",X"B6",X"34",X"1F",X"37",X"70",X"39",X"B1",X"3B",X"D4",X"3D",X"EC",X"3F",
		X"E8",X"41",X"D8",X"43",X"AF",X"45",X"7A",X"47",X"2C",X"49",X"D7",X"4A",X"65",X"4C",X"F3",X"4D",
		X"5F",X"4F",X"D4",X"50",X"17",X"52",X"9F",X"53",X"8D",X"55",X"AF",X"56",X"E1",X"57",X"F2",X"58",
		X"03",X"5A",X"01",X"5B",X"FA",X"5B",X"E2",X"5C",X"C4",X"5D",X"97",X"5E",X"66",X"5F",X"26",X"60",
		X"E0",X"60",X"8E",X"61",X"36",X"62",X"D2",X"62",X"68",X"63",X"F5",X"63",X"7C",X"64",X"FA",X"64",
		X"72",X"65",X"E1",X"65",X"48",X"66",X"AC",X"66",X"07",X"67",X"5D",X"67",X"AD",X"67",X"F4",X"67",
		X"3B",X"68",X"77",X"68",X"B4",X"68",X"E5",X"68",X"18",X"69",X"3B",X"69",X"6F",X"69",X"F1",X"68",
		X"CB",X"66",X"9D",X"63",X"B3",X"5F",X"65",X"5B",X"D3",X"56",X"27",X"52",X"6F",X"4D",X"C0",X"48",
		X"1C",X"44",X"94",X"3F",X"25",X"3B",X"D2",X"36",X"9E",X"32",X"8A",X"2E",X"94",X"2A",X"C0",X"26",
		X"06",X"23",X"6E",X"1F",X"F0",X"1B",X"92",X"18",X"4D",X"15",X"26",X"12",X"18",X"0F",X"24",X"0C",
		X"49",X"09",X"87",X"06",X"DB",X"03",X"46",X"01",X"C8",X"FE",X"60",X"FC",X"0B",X"FA",X"CC",X"F7",
		X"A0",X"F5",X"87",X"F3",X"7E",X"F1",X"8B",X"EF",X"A7",X"ED",X"D4",X"EB",X"11",X"EA",X"5C",X"E8",
		X"BB",X"E6",X"25",X"E5",X"9F",X"E3",X"27",X"E2",X"BB",X"E0",X"5F",X"DF",X"0D",X"DE",X"C8",X"DC",
		X"90",X"DB",X"65",X"DA",X"42",X"D9",X"29",X"D8",X"20",X"D7",X"1C",X"D6",X"24",X"D5",X"35",X"D4",
		X"50",X"D3",X"74",X"D2",X"A1",X"D1",X"D6",X"D0",X"14",X"D0",X"59",X"CF",X"A6",X"CE",X"FA",X"CD",
		X"56",X"CD",X"BA",X"CC",X"23",X"CC",X"92",X"CB",X"0B",X"CB",X"87",X"CA",X"09",X"CA",X"92",X"C9",
		X"22",X"C9",X"B4",X"C8",X"50",X"C8",X"EC",X"C7",X"91",X"C7",X"39",X"C7",X"E7",X"C6",X"95",X"C6",
		X"50",X"C6",X"08",X"C6",X"E0",X"C6",X"38",X"C9",X"70",X"CC",X"44",X"D0",X"6C",X"D4",X"CB",X"D8",
		X"3B",X"DD",X"B3",X"E1",X"1C",X"E6",X"78",X"EA",X"B9",X"EE",X"E1",X"F2",X"EB",X"F6",X"D8",X"FA",
		X"A4",X"FE",X"53",X"02",X"E2",X"05",X"54",X"09",X"AB",X"0C",X"E1",X"0F",X"03",X"13",X"02",X"16",
		X"E9",X"18",X"B6",X"1B",X"6C",X"1E",X"04",X"21",X"93",X"23",X"B7",X"25",X"3F",X"26",X"85",X"25",
		X"FE",X"23",X"EC",X"21",X"86",X"1F",X"ED",X"1C",X"36",X"1A",X"78",X"17",X"B6",X"14",X"FE",X"11",
		X"4E",X"0F",X"AE",X"0C",X"20",X"0A",X"A2",X"07",X"39",X"05",X"DF",X"02",X"9D",X"00",X"6B",X"FE",
		X"4C",X"FC",X"3D",X"FA",X"42",X"F8",X"57",X"F6",X"7D",X"F4",X"B2",X"F2",X"F9",X"F0",X"4E",X"EF",
		X"B3",X"ED",X"23",X"EC",X"A5",X"EA",X"30",X"E9",X"CE",X"E7",X"73",X"E6",X"29",X"E5",X"E8",X"E3",
		X"B5",X"E2",X"8B",X"E1",X"6E",X"E0",X"5A",X"DF",X"51",X"DE",X"51",X"DD",X"5D",X"DC",X"70",X"DB",
		X"8E",X"DA",X"B3",X"D9",X"E1",X"D8",X"15",X"D8",X"55",X"D7",X"9A",X"D6",X"EB",X"D5",X"3E",X"D5",
		X"9B",X"D4",X"FC",X"D3",X"67",X"D3",X"D5",X"D2",X"76",X"D2",X"88",X"D3",X"E0",X"D5",X"FB",X"D8",
		X"97",X"DC",X"7C",X"E0",X"8D",X"E4",X"AB",X"E8",X"CD",X"EC",X"E2",X"F0",X"E5",X"F4",X"D2",X"F8",
		X"A6",X"FC",X"5C",X"00",X"F8",X"03",X"78",X"07",X"DC",X"0A",X"22",X"0E",X"4D",X"11",X"5C",X"14",
		X"52",X"17",X"2B",X"1A",X"EF",X"1C",X"97",X"1F",X"29",X"22",X"A5",X"24",X"08",X"27",X"57",X"29",
		X"91",X"2B",X"B5",X"2D",X"C6",X"2F",X"C4",X"31",X"B0",X"33",X"88",X"35",X"4F",X"37",X"05",X"39",
		X"AC",X"3A",X"42",X"3C",X"C8",X"3D",X"40",X"3F",X"AA",X"40",X"05",X"42",X"51",X"43",X"92",X"44",
		X"C5",X"45",X"EA",X"46",X"07",X"48",X"15",X"49",X"19",X"4A",X"0F",X"4B",X"FD",X"4B",X"E1",X"4C",
		X"BA",X"4D",X"8A",X"4E",X"50",X"4F",X"FA",X"4F",X"51",X"4F",X"50",X"4D",X"85",X"4A",X"2E",X"47",
		X"86",X"43",X"AF",X"3F",X"C5",X"3B",X"D5",X"37",X"ED",X"33",X"13",X"30",X"4E",X"2C",X"A0",X"28",
		X"0A",X"25",X"8E",X"21",X"2A",X"1E",X"E3",X"1A",X"B6",X"17",X"A0",X"14",X"A7",X"11",X"C6",X"0E",
		X"F9",X"0B",X"4A",X"09",X"AB",X"06",X"29",X"04",X"B5",X"01",X"60",X"FF",X"0D",X"FD",X"59",X"FB",
		X"3E",X"FB",X"2F",X"FC",X"E0",X"FD",X"02",X"00",X"72",X"02",X"09",X"05",X"B8",X"07",X"6D",X"0A",
		X"1F",X"0D",X"C8",X"0F",X"64",X"12",X"EF",X"14",X"6A",X"17",X"D0",X"19",X"24",X"1C",X"66",X"1E",
		X"92",X"20",X"AE",X"22",X"B3",X"24",X"A9",X"26",X"8E",X"28",X"60",X"2A",X"20",X"2C",X"D3",X"2D",
		X"72",X"2F",X"04",X"31",X"86",X"32",X"F9",X"33",X"60",X"35",X"B8",X"36",X"02",X"38",X"40",X"39",
		X"70",X"3A",X"96",X"3B",X"AE",X"3C",X"BD",X"3D",X"C1",X"3E",X"B9",X"3F",X"A6",X"40",X"8A",X"41",
		X"64",X"42",X"35",X"43",X"FB",X"43",X"BB",X"44",X"6F",X"45",X"21",X"46",X"C4",X"46",X"64",X"47",
		X"F8",X"47",X"89",X"48",X"0F",X"49",X"91",X"49",X"08",X"4A",X"87",X"4A",X"9D",X"4A",X"35",X"49",
		X"BA",X"46",X"8A",X"43",X"ED",X"3F",X"0D",X"3C",X"0E",X"38",X"FD",X"33",X"F3",X"2F",X"F1",X"2B",
		X"03",X"28",X"2B",X"24",X"6B",X"20",X"C7",X"1C",X"3A",X"19",X"CE",X"15",X"77",X"12",X"40",X"0F",
		X"22",X"0C",X"1E",X"09",X"30",X"06",X"5E",X"03",X"A3",X"00",X"01",X"FE",X"72",X"FB",X"FD",X"F8",
		X"9B",X"F6",X"4F",X"F4",X"15",X"F2",X"F1",X"EF",X"DD",X"ED",X"DE",X"EB",X"EE",X"E9",X"12",X"E8",
		X"43",X"E6",X"88",X"E4",X"DA",X"E2",X"3E",X"E1",X"AF",X"DF",X"30",X"DE",X"BC",X"DC",X"58",X"DB",
		X"FE",X"D9",X"B4",X"D8",X"74",X"D7",X"42",X"D6",X"19",X"D5",X"FE",X"D3",X"EB",X"D2",X"E6",X"D1",
		X"E6",X"D0",X"F6",X"CF",X"09",X"CF",X"2F",X"CE",X"4C",X"CD",X"41",X"CD",X"B1",X"CE",X"02",X"D1",
		X"F5",X"D3",X"3F",X"D7",X"C6",X"DA",X"65",X"DE",X"11",X"E2",X"B4",X"E5",X"50",X"E9",X"D7",X"EC",
		X"4D",X"F0",X"A7",X"F3",X"EE",X"F6",X"18",X"FA",X"2E",X"FD",X"24",X"00",X"05",X"03",X"CD",X"05",
		X"7F",X"08",X"17",X"0B",X"9A",X"0D",X"06",X"10",X"5F",X"12",X"A1",X"14",X"D1",X"16",X"EC",X"18",
		X"F5",X"1A",X"E9",X"1C",X"CF",X"1E",X"A0",X"20",X"63",X"22",X"14",X"24",X"B7",X"25",X"46",X"27",
		X"CD",X"28",X"41",X"2A",X"AA",X"2B",X"00",X"2D",X"53",X"2E",X"8E",X"2F",X"C6",X"30",X"EA",X"31",
		X"0B",X"33",X"15",X"34",X"24",X"35",X"11",X"36",X"2C",X"37",X"8A",X"38",X"60",X"39",X"3D",X"3A",
		X"06",X"3B",X"CD",X"3B",X"88",X"3C",X"3E",X"3D",X"E8",X"3D",X"8D",X"3E",X"2A",X"3F",X"BE",X"3F",
		X"4E",X"40",X"D6",X"40",X"55",X"41",X"CF",X"41",X"43",X"42",X"B1",X"42",X"1B",X"43",X"7C",X"43",
		X"DA",X"43",X"33",X"44",X"83",X"44",X"D2",X"44",X"1A",X"45",X"5F",X"45",X"9C",X"45",X"D8",X"45",
		X"0F",X"46",X"42",X"46",X"70",X"46",X"9C",X"46",X"C3",X"46",X"E8",X"46",X"06",X"47",X"16",X"47",
		X"F5",X"45",X"8E",X"43",X"69",X"40",X"BF",X"3C",X"D0",X"38",X"B4",X"34",X"8C",X"30",X"5F",X"2C",
		X"42",X"28",X"32",X"24",X"39",X"20",X"59",X"1C",X"97",X"18",X"ED",X"14",X"61",X"11",X"F1",X"0D",
		X"9D",X"0A",X"63",X"07",X"44",X"04",X"41",X"01",X"55",X"FE",X"86",X"FB",X"C9",X"F8",X"2B",X"F6",
		X"9A",X"F3",X"2D",X"F1",X"C0",X"EE",X"E1",X"EC",X"83",X"EC",X"31",X"ED",X"95",X"EE",X"69",X"F0",
		X"87",X"F2",X"D2",X"F4",X"31",X"F7",X"9A",X"F9",X"01",X"FC",X"64",X"FE",X"BA",X"00",X"01",X"03",
		X"3C",X"05",X"65",X"07",X"7E",X"09",X"86",X"0B",X"7E",X"0D",X"63",X"0F",X"39",X"11",X"FD",X"12",
		X"B3",X"14",X"58",X"16",X"F2",X"17",X"79",X"19",X"F7",X"1A",X"60",X"1C",X"BF",X"1D",X"0E",X"1E",
		X"00",X"1D",X"24",X"1B",X"B3",X"18",X"F4",X"15",X"FA",X"12",X"E9",X"0F",X"CA",X"0C",X"B3",X"09",
		X"9F",X"06",X"9E",X"03",X"AB",X"00",X"D0",X"FD",X"06",X"FB",X"53",X"F8",X"B3",X"F5",X"2C",X"F3",
		X"B6",X"F0",X"58",X"EE",X"0E",X"EC",X"D7",X"E9",X"B4",X"E7",X"A3",X"E5",X"A4",X"E3",X"B9",X"E1",
		X"DE",X"DF",X"13",X"DE",X"5B",X"DC",X"B2",X"DA",X"16",X"D9",X"8B",X"D7",X"0D",X"D6",X"9E",X"D4",
		X"3C",X"D3",X"E6",X"D1",X"9E",X"D0",X"62",X"CF",X"34",X"CE",X"10",X"CD",X"F7",X"CB",X"E9",X"CA",
		X"E7",X"C9",X"ED",X"C8",X"FE",X"C7",X"18",X"C7",X"3E",X"C6",X"69",X"C5",X"A1",X"C4",X"DA",X"C3",
		X"24",X"C3",X"71",X"C2",X"CA",X"C1",X"23",X"C1",X"8F",X"C0",X"F3",X"BF",X"36",X"C0",X"DD",X"C1",
		X"4F",X"C4",X"59",X"C7",X"B1",X"CA",X"40",X"CE",X"E4",X"D1",X"8F",X"D5",X"34",X"D9",X"D0",X"DC",
		X"54",X"E0",X"C8",X"E3",X"23",X"E7",X"66",X"EA",X"90",X"ED",X"A2",X"F0",X"99",X"F3",X"79",X"F6",
		X"43",X"F9",X"F3",X"FB",X"8D",X"FE",X"0F",X"01",X"7E",X"03",X"D7",X"05",X"1B",X"08",X"4C",X"0A",
		X"68",X"0C",X"73",X"0E",X"6D",X"10",X"54",X"12",X"28",X"14",X"EE",X"15",X"A4",X"17",X"4A",X"19",
		X"E1",X"1A",X"68",X"1C",X"E1",X"1D",X"4E",X"1F",X"AD",X"20",X"FE",X"21",X"44",X"23",X"7E",X"24",
		X"AA",X"25",X"CC",X"26",X"E3",X"27",X"F0",X"28",X"F4",X"29",X"E8",X"2A",X"D8",X"2B",X"B9",X"2C",
		X"99",X"2D",X"67",X"2E",X"35",X"2F",X"EF",X"2F",X"B6",X"30",X"C4",X"30",X"70",X"2F",X"3F",X"2D",
		X"73",X"2A",X"51",X"27",X"F8",X"23",X"87",X"20",X"0A",X"1D",X"90",X"19",X"20",X"16",X"C2",X"12",
		X"78",X"0F",X"43",X"0C",X"25",X"09",X"1F",X"06",X"30",X"03",X"5A",X"00",X"9A",X"FD",X"F2",X"FA",
		X"60",X"F8",X"E3",X"F5",X"7D",X"F3",X"2A",X"F1",X"ED",X"EE",X"C2",X"EC",X"AC",X"EA",X"A7",X"E8",
		X"B5",X"E6",X"D4",X"E4",X"03",X"E3",X"43",X"E1",X"94",X"DF",X"F4",X"DD",X"62",X"DC",X"DF",X"DA",
		X"68",X"D9",X"02",X"D8",X"A8",X"D6",X"5A",X"D5",X"18",X"D4",X"E4",X"D2",X"BA",X"D1",X"9D",X"D0",
		X"89",X"CF",X"81",X"CE",X"83",X"CD",X"8D",X"CC",X"A4",X"CB",X"C3",X"CA",X"EC",X"C9",X"1C",X"C9",
		X"56",X"C8",X"98",X"C7",X"E1",X"C6",X"33",X"C6",X"8A",X"C5",X"EC",X"C4",X"53",X"C4",X"C1",X"C3",
		X"38",X"C3",X"B1",X"C2",X"33",X"C2",X"BA",X"C1",X"48",X"C1",X"DB",X"C0",X"74",X"C0",X"11",X"C0",
		X"B6",X"BF",X"5E",X"BF",X"0B",X"BF",X"BD",X"BE",X"74",X"BE",X"2E",X"BE",X"ED",X"BD",X"AF",X"BD",
		X"77",X"BD",X"43",X"BD",X"0F",X"BD",X"E3",X"BC",X"B8",X"BC",X"92",X"BC",X"6E",X"BC",X"4F",X"BC",
		X"30",X"BC",X"19",X"BC",X"00",X"BC",X"EC",X"BB",X"DA",X"BB",X"CB",X"BB",X"BF",X"BB",X"B5",X"BB",
		X"AB",X"BB",X"A8",X"BB",X"A5",X"BB",X"A4",X"BB",X"A3",X"BB",X"A7",X"BB",X"AD",X"BB",X"B5",X"BB",
		X"BC",X"BB",X"C7",X"BB",X"D2",X"BB",X"E2",X"BB",X"F0",X"BB",X"02",X"BC",X"12",X"BC",X"28",X"BC",
		X"3A",X"BC",X"56",X"BC",X"64",X"BC",X"D0",X"BC",X"8D",X"BE",X"38",X"C1",X"80",X"C4",X"25",X"C8",
		X"01",X"CC",X"F5",X"CF",X"F1",X"D3",X"E8",X"D7",X"D1",X"DB",X"A6",X"DF",X"67",X"E3",X"0B",X"E7",
		X"97",X"EA",X"07",X"EE",X"5E",X"F1",X"97",X"F4",X"B8",X"F7",X"BE",X"FA",X"AB",X"FD",X"7C",X"00",
		X"3A",X"03",X"DC",X"05",X"6C",X"08",X"E0",X"0A",X"45",X"0D",X"8D",X"0F",X"CB",X"11",X"15",X"13",
		X"09",X"13",X"37",X"12",X"CF",X"10",X"14",X"0F",X"1C",X"0D",X"04",X"0B",X"DC",X"08",X"B1",X"06",
		X"88",X"04",X"66",X"02",X"4C",X"00",X"42",X"FE",X"45",X"FC",X"55",X"FA",X"74",X"F8",X"A5",X"F6",
		X"E5",X"F4",X"32",X"F3",X"8D",X"F1",X"F6",X"EF",X"6E",X"EE",X"F5",X"EC",X"89",X"EB",X"26",X"EA",
		X"D6",X"E8",X"87",X"E7",X"82",X"E6",X"C4",X"E6",X"0E",X"E8",X"FF",X"E9",X"5D",X"EC",X"FF",X"EE",
		X"C4",X"F1",X"9C",X"F4",X"79",X"F7",X"4F",X"FA",X"1C",X"FD",X"D9",X"FF",X"87",X"02",X"1F",X"05",
		X"A8",X"07",X"1B",X"0A",X"7A",X"0C",X"C5",X"0E",X"FB",X"10",X"20",X"13",X"33",X"15",X"31",X"17",
		X"22",X"19",X"FE",X"1A",X"C8",X"1C",X"84",X"1E",X"2F",X"20",X"CB",X"21",X"5A",X"23",X"D7",X"24",
		X"48",X"26",X"AA",X"27",X"01",X"29",X"4A",X"2A",X"87",X"2B",X"B7",X"2C",X"DC",X"2D",X"F5",X"2E",
		X"04",X"30",X"07",X"31",X"03",X"32",X"F1",X"32",X"D9",X"33",X"B5",X"34",X"88",X"35",X"54",X"36",
		X"16",X"37",X"CE",X"37",X"83",X"38",X"2B",X"39",X"CF",X"39",X"68",X"3A",X"02",X"3B",X"88",X"3B",
		X"1D",X"3C",X"11",X"3C",X"B8",X"3A",X"8F",X"38",X"D5",X"35",X"CA",X"32",X"8A",X"2F",X"33",X"2C",
		X"D1",X"28",X"73",X"25",X"1F",X"22",X"DC",X"1E",X"AB",X"1B",X"8F",X"18",X"89",X"15",X"9A",X"12",
		X"C1",X"0F",X"FF",X"0C",X"54",X"0A",X"BE",X"07",X"3E",X"05",X"D6",X"02",X"80",X"00",X"38",X"FE",
		X"05",X"FC",X"E3",X"F9",X"D3",X"F7",X"D6",X"F5",X"F9",X"F3",X"3C",X"F3",X"AD",X"F3",X"D3",X"F4",
		X"78",X"F6",X"69",X"F8",X"8C",X"FA",X"C6",X"FC",X"0C",X"FF",X"52",X"01",X"97",X"03",X"CF",X"05",
		X"FC",X"07",X"1A",X"0A",X"2A",X"0C",X"28",X"0E",X"16",X"10",X"F7",X"11",X"C6",X"13",X"85",X"15",
		X"34",X"17",X"D8",X"18",X"68",X"1A",X"ED",X"1B",X"60",X"1D",X"CD",X"1E",X"22",X"20",X"7D",X"21",
		X"59",X"22",X"E3",X"21",X"8B",X"20",X"96",X"1E",X"44",X"1C",X"B7",X"19",X"09",X"17",X"4B",X"14",
		X"8B",X"11",X"CF",X"0E",X"20",X"0C",X"7E",X"09",X"EC",X"06",X"6C",X"04",X"00",X"02",X"A7",X"FF",
		X"60",X"FD",X"2A",X"FB",X"08",X"F9",X"F8",X"F6",X"F9",X"F4",X"0B",X"F3",X"30",X"F1",X"63",X"EF",
		X"A8",X"ED",X"FA",X"EB",X"5D",X"EA",X"CD",X"E8",X"4C",X"E7",X"D8",X"E5",X"71",X"E4",X"18",X"E3",
		X"C9",X"E1",X"8B",X"E0",X"55",X"DF",X"2B",X"DE",X"0B",X"DD",X"F8",X"DB",X"ED",X"DA",X"EE",X"D9",
		X"F8",X"D8",X"0A",X"D8",X"28",X"D7",X"4E",X"D6",X"7A",X"D5",X"B3",X"D4",X"EF",X"D3",X"36",X"D3",
		X"83",X"D2",X"DA",X"D1",X"33",X"D1",X"9A",X"D0",X"00",X"D0",X"74",X"CF",X"E1",X"CE",X"A4",X"CE",
		X"A5",X"CF",X"92",X"D1",X"16",X"D4",X"F9",X"D6",X"15",X"DA",X"4F",X"DD",X"94",X"E0",X"D8",X"E3",
		X"13",X"E7",X"41",X"EA",X"5B",X"ED",X"62",X"F0",X"52",X"F3",X"30",X"F6",X"F3",X"F8",X"A0",X"FB",
		X"3A",X"FE",X"BD",X"00",X"29",X"03",X"82",X"05",X"C6",X"07",X"F7",X"09",X"14",X"0C",X"21",X"0E",
		X"18",X"10",X"01",X"12",X"D8",X"13",X"9D",X"15",X"53",X"17",X"FB",X"18",X"94",X"1A",X"1C",X"1C",
		X"95",X"1D",X"04",X"1F",X"62",X"20",X"B6",X"21",X"FB",X"22",X"38",X"24",X"65",X"25",X"8A",X"26",
		X"A1",X"27",X"AF",X"28",X"B2",X"29",X"AB",X"2A",X"9A",X"2B",X"80",X"2C",X"5C",X"2D",X"31",X"2E",
		X"FC",X"2E",X"C0",X"2F",X"79",X"30",X"2D",X"31",X"D5",X"31",X"7F",X"32",X"F1",X"32",X"39",X"32",
		X"81",X"30",X"31",X"2E",X"7B",X"2B",X"88",X"28",X"74",X"25",X"54",X"22",X"2F",X"1F",X"15",X"1C",
		X"04",X"19",X"08",X"16",X"1A",X"13",X"43",X"10",X"81",X"0D",X"D4",X"0A",X"3C",X"08",X"BA",X"05",
		X"4B",X"03",X"F2",X"00",X"AB",X"FE",X"79",X"FC",X"5A",X"FA",X"4C",X"F8",X"4F",X"F6",X"65",X"F4",
		X"8A",X"F2",X"C1",X"F0",X"09",X"EF",X"5E",X"ED",X"C4",X"EB",X"37",X"EA",X"B6",X"E8",X"46",X"E7",
		X"E1",X"E5",X"89",X"E4",X"3F",X"E3",X"FF",X"E1",X"CA",X"E0",X"A3",X"DF",X"85",X"DE",X"73",X"DD",
		X"6A",X"DC",X"6B",X"DB",X"75",X"DA",X"89",X"D9",X"A7",X"D8",X"CD",X"D7",X"FC",X"D6",X"34",X"D6",
		X"72",X"D5",X"B9",X"D4",X"08",X"D4",X"5D",X"D3",X"B9",X"D2",X"1D",X"D2",X"86",X"D1",X"F7",X"D0",
		X"6F",X"D0",X"EA",X"CF",X"6D",X"CF",X"F6",X"CE",X"84",X"CE",X"17",X"CE",X"B0",X"CD",X"4F",X"CD",
		X"EF",X"CC",X"96",X"CC",X"41",X"CC",X"F1",X"CB",X"A6",X"CB",X"5E",X"CB",X"1B",X"CB",X"DA",X"CA",
		X"9E",X"CA",X"66",X"CA",X"31",X"CA",X"01",X"CA",X"D1",X"C9",X"A6",X"C9",X"7F",X"C9",X"59",X"C9",
		X"38",X"C9",X"19",X"C9",X"FC",X"C8",X"E4",X"C8",X"CC",X"C8",X"B7",X"C8",X"A3",X"C8",X"94",X"C8",
		X"85",X"C8",X"7A",X"C8",X"70",X"C8",X"69",X"C8",X"63",X"C8",X"5F",X"C8",X"5E",X"C8",X"5E",X"C8",
		X"61",X"C8",X"62",X"C8",X"69",X"C8",X"6E",X"C8",X"76",X"C8",X"80",X"C8",X"8C",X"C8",X"97",X"C8",
		X"A5",X"C8",X"B3",X"C8",X"C2",X"C8",X"D5",X"C8",X"E5",X"C8",X"F9",X"C8",X"0F",X"C9",X"23",X"C9",
		X"3B",X"C9",X"52",X"C9",X"6B",X"C9",X"83",X"C9",X"9E",X"C9",X"B8",X"C9",X"D3",X"C9",X"EE",X"C9",
		X"0D",X"CA",X"2A",X"CA",X"4B",X"CA",X"68",X"CA",X"8B",X"CA",X"A9",X"CA",X"CB",X"CA",X"EA",X"CA",
		X"0D",X"CB",X"30",X"CB",X"54",X"CB",X"74",X"CB",X"9C",X"CB",X"BD",X"CB",X"E8",X"CB",X"04",X"CC",
		X"78",X"CC",X"18",X"CE",X"86",X"D0",X"7E",X"D3",X"C4",X"D6",X"3D",X"DA",X"CA",X"DD",X"5A",X"E1",
		X"E7",X"E4",X"68",X"E8",X"D7",X"EB",X"2F",X"EF",X"73",X"F2",X"9E",X"F5",X"B1",X"F8",X"AB",X"FB",
		X"8E",X"FE",X"56",X"01",X"0A",X"04",X"A4",X"06",X"2A",X"09",X"99",X"0B",X"F5",X"0D",X"3A",X"10",
		X"6B",X"12",X"8A",X"14",X"96",X"16",X"90",X"18",X"77",X"1A",X"4D",X"1C",X"14",X"1E",X"C9",X"1F",
		X"70",X"21",X"07",X"23",X"8F",X"24",X"08",X"26",X"75",X"27",X"D2",X"28",X"24",X"2A",X"67",X"2B",
		X"A2",X"2C",X"CE",X"2D",X"F0",X"2E",X"05",X"30",X"12",X"31",X"12",X"32",X"09",X"33",X"F6",X"33",
		X"DA",X"34",X"B3",X"35",X"85",X"36",X"4C",X"37",X"0F",X"38",X"C4",X"38",X"79",X"39",X"ED",X"39",
		X"40",X"39",X"AD",X"37",X"8C",X"35",X"0C",X"33",X"57",X"30",X"81",X"2D",X"9F",X"2A",X"BC",X"27",
		X"E0",X"24",X"0E",X"22",X"4B",X"1F",X"9A",X"1C",X"FB",X"19",X"6F",X"17",X"F4",X"14",X"92",X"12",
		X"3D",X"10",X"00",X"0E",X"D2",X"0B",X"B9",X"09",X"AE",X"07",X"BB",X"05",X"D0",X"03",X"FC",X"01",
		X"31",X"00",X"81",X"FE",X"D0",X"FC",X"D4",X"FB",X"06",X"FC",X"ED",X"FC",X"58",X"FE",X"0D",X"00",
		X"F7",X"01",X"FA",X"03",X"0C",X"06",X"1F",X"08",X"31",X"0A",X"39",X"0C",X"38",X"0E",X"28",X"10",
		X"0B",X"12",X"E0",X"13",X"A6",X"15",X"5E",X"17",X"04",X"19",X"A0",X"1A",X"2A",X"1C",X"A9",X"1D",
		X"18",X"1F",X"7D",X"20",X"D1",X"21",X"1E",X"23",X"55",X"24",X"91",X"25",X"35",X"26",X"B0",X"25",
		X"6E",X"24",X"A6",X"22",X"95",X"20",X"4E",X"1E",X"EE",X"1B",X"83",X"19",X"15",X"17",X"AD",X"14",
		X"4E",X"12",X"FD",X"0F",X"BA",X"0D",X"85",X"0B",X"63",X"09",X"4F",X"07",X"4F",X"05",X"5A",X"03",
		X"7A",X"01",X"A8",X"FF",X"E6",X"FD",X"32",X"FC",X"8F",X"FA",X"F7",X"F8",X"71",X"F7",X"F3",X"F5",
		X"86",X"F4",X"33",X"F3",X"DE",X"F2",X"8C",X"F3",X"D5",X"F4",X"8A",X"F6",X"80",X"F8",X"9C",X"FA",
		X"CD",X"FC",X"05",X"FF",X"3C",X"01",X"6B",X"03",X"94",X"05",X"AD",X"07",X"BA",X"09",X"B5",X"0B",
		X"A4",X"0D",X"80",X"0F",X"4F",X"11",X"0B",X"13",X"C0",X"14",X"5A",X"16",X"FD",X"17",X"B6",X"19",
		X"2E",X"1B",X"9A",X"1C",X"FD",X"1D",X"4A",X"1F",X"99",X"20",X"76",X"21",X"23",X"21",X"0C",X"20",
		X"6B",X"1E",X"77",X"1C",X"4D",X"1A",X"07",X"18",X"B1",X"15",X"5A",X"13",X"08",X"11",X"BB",X"0E",
		X"7F",X"0C",X"4E",X"0A",X"2A",X"08",X"17",X"06",X"15",X"04",X"23",X"02",X"3F",X"00",X"6E",X"FE",
		X"AB",X"FC",X"F7",X"FA",X"51",X"F9",X"B8",X"F7",X"2F",X"F6",X"B3",X"F4",X"45",X"F3",X"E2",X"F1",
		X"8C",X"F0",X"42",X"EF",X"04",X"EE",X"CF",X"EC",X"A9",X"EB",X"8B",X"EA",X"77",X"E9",X"6F",X"E8",
		X"6E",X"E7",X"77",X"E6",X"8A",X"E5",X"A6",X"E4",X"C9",X"E3",X"F8",X"E2",X"2B",X"E2",X"68",X"E1",
		X"AA",X"E0",X"F7",X"DF",X"49",X"DF",X"A1",X"DE",X"01",X"DE",X"66",X"DD",X"D4",X"DC",X"45",X"DC",
		X"BE",X"DB",X"3D",X"DB",X"C0",X"DA",X"48",X"DA",X"D6",X"D9",X"69",X"D9",X"02",X"D9",X"9F",X"D8",
		X"41",X"D8",X"E7",X"D7",X"90",X"D7",X"3F",X"D7",X"F1",X"D6",X"A7",X"D6",X"61",X"D6",X"1E",X"D6",
		X"E0",X"D5",X"A4",X"D5",X"6D",X"D5",X"36",X"D5",X"06",X"D5",X"D5",X"D4",X"AB",X"D4",X"81",X"D4",
		X"5C",X"D4",X"37",X"D4",X"18",X"D4",X"F8",X"D3",X"DD",X"D3",X"C2",X"D3",X"AE",X"D3",X"93",X"D3",
		X"31",X"D4",X"DA",X"D5",X"21",X"D8",X"D9",X"DA",X"C8",X"DD",X"DF",X"E0",X"02",X"E4",X"29",X"E7",
		X"48",X"EA",X"5C",X"ED",X"5B",X"F0",X"4C",X"F3",X"27",X"F6",X"ED",X"F8",X"9C",X"FB",X"38",X"FE",
		X"BD",X"00",X"2D",X"03",X"88",X"05",X"D0",X"07",X"06",X"0A",X"25",X"0C",X"32",X"0E",X"2E",X"10",
		X"1A",X"12",X"F3",X"13",X"BD",X"15",X"76",X"17",X"1F",X"19",X"BB",X"1A",X"46",X"1C",X"C2",X"1D",
		X"34",X"1F",X"96",X"20",X"EB",X"21",X"36",X"23",X"72",X"24",X"A2",X"25",X"C9",X"26",X"E4",X"27",
		X"F3",X"28",X"F9",X"29",X"F5",X"2A",X"E5",X"2B",X"CF",X"2C",X"AE",X"2D",X"85",X"2E",X"51",X"2F",
		X"19",X"30",X"D2",X"30",X"8B",X"31",X"36",X"32",X"E1",X"32",X"79",X"33",X"1A",X"34",X"22",X"34",
		X"13",X"33",X"5C",X"31",X"2F",X"2F",X"C1",X"2C",X"25",X"2A",X"76",X"27",X"C1",X"24",X"0E",X"22",
		X"62",X"1F",X"C4",X"1C",X"33",X"1A",X"B3",X"17",X"46",X"15",X"EB",X"12",X"A1",X"10",X"6A",X"0E",
		X"44",X"0C",X"32",X"0A",X"2E",X"08",X"3C",X"06",X"5B",X"04",X"8B",X"02",X"C9",X"00",X"17",X"FF",
		X"75",X"FD",X"DE",X"FB",X"6C",X"FA",X"F7",X"F9",X"70",X"FA",X"7A",X"FB",X"EB",X"FC",X"96",X"FE",
		X"66",X"00",X"49",X"02",X"37",X"04",X"23",X"06",X"0C",X"08",X"E9",X"09",X"BF",X"0B",X"85",X"0D",
		X"41",X"0F",X"ED",X"10",X"8E",X"12",X"20",X"14",X"A4",X"15",X"1C",X"17",X"86",X"18",X"E4",X"19",
		X"35",X"1B",X"79",X"1C",X"B2",X"1D",X"DF",X"1E",X"04",X"20",X"1A",X"21",X"29",X"22",X"2B",X"23",
		X"25",X"24",X"15",X"25",X"FD",X"25",X"D9",X"26",X"AE",X"27",X"7A",X"28",X"3F",X"29",X"FC",X"29",
		X"B0",X"2A",X"5F",X"2B",X"04",X"2C",X"A4",X"2C",X"3C",X"2D",X"CE",X"2D",X"59",X"2E",X"DF",X"2E",
		X"5F",X"2F",X"D8",X"2F",X"4B",X"30",X"BC",X"30",X"24",X"31",X"89",X"31",X"E7",X"31",X"43",X"32",
		X"99",X"32",X"E1",X"32",X"52",X"32",X"D1",X"30",X"C6",X"2E",X"57",X"2C",X"B3",X"29",X"EE",X"26",
		X"1C",X"24",X"49",X"21",X"7B",X"1E",X"B7",X"1B",X"03",X"19",X"60",X"16",X"D0",X"13",X"51",X"11",
		X"E5",X"0E",X"8E",X"0C",X"47",X"0A",X"13",X"08",X"F3",X"05",X"E4",X"03",X"E6",X"01",X"FA",X"FF",
		X"1F",X"FE",X"52",X"FC",X"96",X"FA",X"E9",X"F8",X"4B",X"F7",X"BA",X"F5",X"36",X"F4",X"C0",X"F2",
		X"58",X"F1",X"FC",X"EF",X"AC",X"EE",X"6A",X"ED",X"30",X"EC",X"01",X"EB",X"DF",X"E9",X"C8",X"E8",
		X"BB",X"E7",X"B6",X"E6",X"BA",X"E5",X"C9",X"E4",X"E0",X"E3",X"02",X"E3",X"28",X"E2",X"5B",X"E1",
		X"92",X"E0",X"D4",X"DF",X"1A",X"DF",X"6B",X"DE",X"C0",X"DD",X"1F",X"DD",X"80",X"DC",X"EC",X"DB",
		X"5A",X"DB",X"85",X"DB",X"AD",X"DC",X"65",X"DE",X"86",X"E0",X"DF",X"E2",X"5E",X"E5",X"EC",X"E7",
		X"80",X"EA",X"0D",X"ED",X"95",X"EF",X"0E",X"F2",X"79",X"F4",X"D3",X"F6",X"1C",X"F9",X"53",X"FB",
		X"79",X"FD",X"8B",X"FF",X"8F",X"01",X"80",X"03",X"62",X"05",X"32",X"07",X"F3",X"08",X"A5",X"0A",
		X"48",X"0C",X"DE",X"0D",X"63",X"0F",X"DC",X"10",X"49",X"12",X"A6",X"13",X"FA",X"14",X"40",X"16",
		X"7C",X"17",X"AA",X"18",X"CF",X"19",X"E8",X"1A",X"F7",X"1B",X"FC",X"1C",X"F9",X"1D",X"EB",X"1E",
		X"D3",X"1F",X"B3",X"20",X"8B",X"21",X"5A",X"22",X"22",X"23",X"E2",X"23",X"99",X"24",X"49",X"25",
		X"F2",X"25",X"94",X"26",X"2F",X"27",X"C4",X"27",X"54",X"28",X"DB",X"28",X"60",X"29",X"DD",X"29",
		X"54",X"2A",X"C7",X"2A",X"33",X"2B",X"9B",X"2B",X"FE",X"2B",X"5C",X"2C",X"B6",X"2C",X"0B",X"2D",
		X"5C",X"2D",X"A8",X"2D",X"F2",X"2D",X"37",X"2E",X"79",X"2E",X"B5",X"2E",X"EF",X"2E",X"24",X"2F",
		X"59",X"2F",X"88",X"2F",X"B4",X"2F",X"DF",X"2F",X"05",X"30",X"27",X"30",X"49",X"30",X"68",X"30",
		X"84",X"30",X"9D",X"30",X"B4",X"30",X"C9",X"30",X"DB",X"30",X"EA",X"30",X"F9",X"30",X"05",X"31",
		X"0F",X"31",X"16",X"31",X"1D",X"31",X"21",X"31",X"24",X"31",X"24",X"31",X"24",X"31",X"21",X"31",
		X"1E",X"31",X"18",X"31",X"10",X"31",X"08",X"31",X"01",X"31",X"F6",X"30",X"EB",X"30",X"DD",X"30",
		X"CF",X"30",X"BE",X"30",X"AF",X"30",X"9C",X"30",X"8A",X"30",X"74",X"30",X"69",X"30",X"E3",X"2F",
		X"62",X"2E",X"47",X"2C",X"C1",X"29",X"01",X"27",X"1A",X"24",X"27",X"21",X"30",X"1E",X"3F",X"1B",
		X"58",X"18",X"82",X"15",X"BC",X"12",X"09",X"10",X"6B",X"0D",X"E1",X"0A",X"68",X"08",X"07",X"06",
		X"B7",X"03",X"7B",X"01",X"54",X"FF",X"3D",X"FD",X"38",X"FB",X"44",X"F9",X"62",X"F7",X"8F",X"F5",
		X"CE",X"F3",X"1A",X"F2",X"77",X"F0",X"E0",X"EE",X"5A",X"ED",X"DF",X"EB",X"75",X"EA",X"13",X"E9",
		X"C1",X"E7",X"79",X"E6",X"3F",X"E5",X"0E",X"E4",X"EA",X"E2",X"CF",X"E1",X"C1",X"E0",X"B9",X"DF",
		X"C1",X"DE",X"CA",X"DD",X"E4",X"DC",X"FF",X"DB",X"2C",X"DB",X"56",X"DA",X"9B",X"D9",X"BC",X"D8",
		X"B1",X"D7",X"05",X"D7",X"55",X"D6",X"B4",X"D5",X"15",X"D5",X"84",X"D4",X"B6",X"D4",X"D2",X"D5",
		X"74",X"D7",X"75",X"D9",X"AB",X"DB",X"06",X"DE",X"6C",X"E0",X"D6",X"E2",X"3C",X"E5",X"9C",X"E7",
		X"EE",X"E9",X"34",X"EC",X"69",X"EE",X"90",X"F0",X"A5",X"F2",X"AB",X"F4",X"A1",X"F6",X"85",X"F8",
		X"5B",X"FA",X"20",X"FC",X"D7",X"FD",X"7D",X"FF",X"19",X"01",X"A0",X"02",X"22",X"04",X"90",X"05",
		X"FD",X"06",X"17",X"08",X"30",X"08",X"92",X"07",X"7C",X"06",X"15",X"05",X"7E",X"03",X"C9",X"01",
		X"07",X"00",X"40",X"FE",X"79",X"FC",X"B9",X"FA",X"01",X"F9",X"53",X"F7",X"B1",X"F5",X"1B",X"F4",
		X"91",X"F2",X"14",X"F1",X"A5",X"EF",X"3E",X"EE",X"E8",X"EC",X"9B",X"EB",X"5C",X"EA",X"26",X"E9",
		X"FC",X"E7",X"DB",X"E6",X"C8",X"E5",X"BC",X"E4",X"BA",X"E3",X"C2",X"E2",X"D4",X"E1",X"ED",X"E0",
		X"11",X"E0",X"3C",X"DF",X"71",X"DE",X"AA",X"DD",X"EE",X"DC",X"38",X"DC",X"8A",X"DB",X"E1",X"DA",
		X"42",X"DA",X"A9",X"D9",X"14",X"D9",X"86",X"D8",X"FE",X"D7",X"7C",X"D7",X"01",X"D7",X"89",X"D6",
		X"17",X"D6",X"AA",X"D5",X"43",X"D5",X"E0",X"D4",X"82",X"D4",X"26",X"D4",X"D4",X"D3",X"7D",X"D3",
		X"58",X"D3",X"1D",X"D4",X"9D",X"D5",X"92",X"D7",X"D4",X"D9",X"3E",X"DC",X"C2",X"DE",X"4F",X"E1",
		X"DC",X"E3",X"62",X"E6",X"DD",X"E8",X"47",X"EB",X"A4",X"ED",X"F3",X"EF",X"2E",X"F2",X"56",X"F4",
		X"70",X"F6",X"78",X"F8",X"6F",X"FA",X"55",X"FC",X"2C",X"FE",X"F3",X"FF",X"A8",X"01",X"53",X"03",
		X"EB",X"04",X"7A",X"06",X"F3",X"07",X"6E",X"09",X"55",X"0A",X"42",X"0A",X"9A",X"09",X"83",X"08",
		X"2D",X"07",X"AC",X"05",X"15",X"04",X"71",X"02",X"CA",X"00",X"24",X"FF",X"88",X"FD",X"F0",X"FB",
		X"64",X"FA",X"E1",X"F8",X"6A",X"F7",X"00",X"F6",X"A0",X"F4",X"4C",X"F3",X"03",X"F2",X"C4",X"F0",
		X"93",X"EF",X"6B",X"EE",X"4D",X"ED",X"3B",X"EC",X"30",X"EB",X"31",X"EA",X"37",X"E9",X"60",X"E8",
		X"65",X"E8",X"34",X"E9",X"7E",X"EA",X"1E",X"EC",X"EF",X"ED",X"DD",X"EF",X"DA",X"F1",X"DC",X"F3",
		X"D9",X"F5",X"D2",X"F7",X"C1",X"F9",X"A5",X"FB",X"7A",X"FD",X"42",X"FF",X"FB",X"00",X"A9",X"02",
		X"49",X"04",X"DB",X"05",X"5E",X"07",X"D6",X"08",X"3F",X"0A",X"9E",X"0B",X"EE",X"0C",X"36",X"0E",
		X"6F",X"0F",X"9F",X"10",X"C3",X"11",X"DF",X"12",X"ED",X"13",X"F5",X"14",X"F1",X"15",X"E6",X"16",
		X"CE",X"17",X"B3",X"18",X"89",X"19",X"5D",X"1A",X"26",X"1B",X"E8",X"1B",X"A2",X"1C",X"54",X"1D",
		X"02",X"1E",X"A6",X"1E",X"45",X"1F",X"DE",X"1F",X"70",X"20",X"FD",X"20",X"83",X"21",X"03",X"22",
		X"80",X"22",X"F6",X"22",X"68",X"23",X"D3",X"23",X"3B",X"24",X"9E",X"24",X"F3",X"24",X"86",X"24",
		X"4A",X"23",X"93",X"21",X"87",X"1F",X"50",X"1D",X"F7",X"1A",X"95",X"18",X"30",X"16",X"D2",X"13",
		X"7C",X"11",X"31",X"0F",X"F6",X"0C",X"CA",X"0A",X"AE",X"08",X"A2",X"06",X"A7",X"04",X"BC",X"02",
		X"DF",X"00",X"15",X"FF",X"58",X"FD",X"A8",X"FB",X"0B",X"FA",X"78",X"F8",X"F6",X"F6",X"7D",X"F5",
		X"17",X"F4",X"B3",X"F2",X"A7",X"F1",X"8D",X"F1",X"18",X"F2",X"16",X"F3",X"59",X"F4",X"C9",X"F5",
		X"55",X"F7",X"ED",X"F8",X"8A",X"FA",X"27",X"FC",X"BE",X"FD",X"4E",X"FF",X"D4",X"00",X"4E",X"02",
		X"BF",X"03",X"25",X"05",X"80",X"06",X"CF",X"07",X"14",X"09",X"4C",X"0A",X"7B",X"0B",X"9F",X"0C",
		X"B8",X"0D",X"C9",X"0E",X"CF",X"0F",X"CD",X"10",X"C1",X"11",X"AB",X"12",X"8D",X"13",X"67",X"14",
		X"3B",X"15",X"05",X"16",X"C9",X"16",X"83",X"17",X"38",X"18",X"E4",X"18",X"8C",X"19",X"2C",X"1A",
		X"C7",X"1A",X"5B",X"1B",X"E9",X"1B",X"70",X"1C",X"F3",X"1C",X"72",X"1D",X"E9",X"1D",X"5C",X"1E",
		X"CA",X"1E",X"34",X"1F",X"9A",X"1F",X"FA",X"1F",X"57",X"20",X"AE",X"20",X"03",X"21",X"50",X"21",
		X"A3",X"21",X"BD",X"21",X"FA",X"20",X"8C",X"1F",X"B5",X"1D",X"99",X"1B",X"56",X"19",X"02",X"17",
		X"A1",X"14",X"44",X"12",X"EC",X"0F",X"A1",X"0D",X"60",X"0B",X"2F",X"09",X"0E",X"07",X"FE",X"04",
		X"FB",X"02",X"0C",X"01",X"2C",X"FF",X"5B",X"FD",X"99",X"FB",X"E6",X"F9",X"42",X"F8",X"AC",X"F6",
		X"24",X"F5",X"AA",X"F3",X"3A",X"F2",X"DE",X"F0",X"84",X"EF",X"BE",X"EE",X"DC",X"EE",X"85",X"EF",
		X"90",X"F0",X"D4",X"F1",X"40",X"F3",X"C0",X"F4",X"4B",X"F6",X"D9",X"F7",X"64",X"F9",X"E9",X"FA",
		X"67",X"FC",X"DD",X"FD",X"48",X"FF",X"A6",X"00",X"FA",X"01",X"45",X"03",X"84",X"04",X"BA",X"05",
		X"E5",X"06",X"06",X"08",X"1C",X"09",X"29",X"0A",X"2D",X"0B",X"27",X"0C",X"18",X"0D",X"03",X"0E",
		X"C8",X"0E",X"BA",X"0E",X"F5",X"0D",X"BF",X"0C",X"3B",X"0B",X"8B",X"09",X"C1",X"07",X"EC",X"05",
		X"13",X"04",X"3B",X"02",X"69",X"00",X"A1",X"FE",X"E4",X"FC",X"33",X"FB",X"90",X"F9",X"F8",X"F7",
		X"6D",X"F6",X"EE",X"F4",X"7E",X"F3",X"1A",X"F2",X"C1",X"F0",X"75",X"EF",X"33",X"EE",X"FC",X"EC",
		X"D3",X"EB",X"B0",X"EA",X"9E",X"E9",X"8B",X"E8",X"EE",X"E7",X"37",X"E8",X"08",X"E9",X"40",X"EA",
		X"B0",X"EB",X"4A",X"ED",X"F6",X"EE",X"AC",X"F0",X"64",X"F2",X"19",X"F4",X"C7",X"F5",X"6D",X"F7",
		X"08",X"F9",X"97",X"FA",X"1C",X"FC",X"94",X"FD",X"02",X"FF",X"62",X"00",X"B8",X"01",X"02",X"03",
		X"41",X"04",X"75",X"05",X"9F",X"06",X"BF",X"07",X"D3",X"08",X"DF",X"09",X"E2",X"0A",X"DB",X"0B",
		X"CD",X"0C",X"B5",X"0D",X"94",X"0E",X"6C",X"0F",X"3A",X"10",X"03",X"11",X"C3",X"11",X"7D",X"12",
		X"31",X"13",X"DC",X"13",X"81",X"14",X"21",X"15",X"BA",X"15",X"4E",X"16",X"DC",X"16",X"64",X"17",
		X"E7",X"17",X"64",X"18",X"DD",X"18",X"50",X"19",X"BF",X"19",X"29",X"1A",X"8E",X"1A",X"EE",X"1A",
		X"4D",X"1B",X"A5",X"1B",X"FB",X"1B",X"4C",X"1C",X"9C",X"1C",X"E3",X"1C",X"2B",X"1D",X"6E",X"1D",
		X"AD",X"1D",X"EA",X"1D",X"26",X"1E",X"5B",X"1E",X"8E",X"1E",X"C0",X"1E",X"EF",X"1E",X"1A",X"1F",
		X"44",X"1F",X"6A",X"1F",X"90",X"1F",X"B0",X"1F",X"D3",X"1F",X"EE",X"1F",X"0E",X"20",X"1F",X"20",
		X"4E",X"20",X"A9",X"20",X"B7",X"20",X"CE",X"20",X"D9",X"20",X"F0",X"20",X"C4",X"20",X"C2",X"1F",
		X"2A",X"1E",X"32",X"1C",X"FE",X"19",X"A7",X"17",X"41",X"15",X"D5",X"12",X"6C",X"10",X"0C",X"0E",
		X"B7",X"0B",X"70",X"09",X"37",X"07",X"0E",X"05",X"F8",X"02",X"F1",X"00",X"FC",X"FE",X"16",X"FD",
		X"42",X"FB",X"7A",X"F9",X"C4",X"F7",X"1A",X"F6",X"81",X"F4",X"F5",X"F2",X"76",X"F1",X"05",X"F0",
		X"A1",X"EE",X"48",X"ED",X"FE",X"EB",X"BD",X"EA",X"8A",X"E9",X"60",X"E8",X"41",X"E7",X"2D",X"E6",
		X"22",X"E5",X"21",X"E4",X"2B",X"E3",X"3C",X"E2",X"56",X"E1",X"79",X"E0",X"A6",X"DF",X"DA",X"DE",
		X"15",X"DE",X"58",X"DD",X"A3",X"DC",X"F6",X"DB",X"4D",X"DB",X"AD",X"DA",X"13",X"DA",X"80",X"D9",
		X"F2",X"D8",X"6B",X"D8",X"E7",X"D7",X"6C",X"D7",X"F4",X"D6",X"83",X"D6",X"16",X"D6",X"B0",X"D5",
		X"4C",X"D5",X"ED",X"D4",X"93",X"D4",X"3D",X"D4",X"EC",X"D3",X"9F",X"D3",X"56",X"D3",X"11",X"D3",
		X"CE",X"D2",X"91",X"D2",X"55",X"D2",X"1D",X"D2",X"E8",X"D1",X"B8",X"D1",X"8B",X"D1",X"5F",X"D1",
		X"36",X"D1",X"11",X"D1",X"EF",X"D0",X"CE",X"D0",X"AF",X"D0",X"95",X"D0",X"7C",X"D0",X"66",X"D0",
		X"51",X"D0",X"3F",X"D0",X"2F",X"D0",X"21",X"D0",X"15",X"D0",X"09",X"D0",X"01",X"D0",X"FC",X"CF",
		X"F5",X"CF",X"F2",X"CF",X"F0",X"CF",X"F0",X"CF",X"F1",X"CF",X"F4",X"CF",X"F9",X"CF",X"FD",X"CF",
		X"03",X"D0",X"0D",X"D0",X"15",X"D0",X"1E",X"D0",X"29",X"D0",X"37",X"D0",X"45",X"D0",X"53",X"D0",
		X"62",X"D0",X"73",X"D0",X"86",X"D0",X"95",X"D0",X"BE",X"D0",X"A0",X"D1",X"2A",X"D3",X"16",X"D5",
		X"47",X"D7",X"99",X"D9",X"02",X"DC",X"6F",X"DE",X"DA",X"E0",X"3F",X"E3",X"99",X"E5",X"E4",X"E7",
		X"21",X"EA",X"4E",X"EC",X"6C",X"EE",X"77",X"F0",X"75",X"F2",X"62",X"F4",X"3E",X"F6",X"0C",X"F8",
		X"C9",X"F9",X"78",X"FB",X"19",X"FD",X"AD",X"FE",X"32",X"00",X"AB",X"01",X"17",X"03",X"75",X"04",
		X"CA",X"05",X"11",X"07",X"4E",X"08",X"7F",X"09",X"A7",X"0A",X"C2",X"0B",X"D4",X"0C",X"DE",X"0D",
		X"DE",X"0E",X"D5",X"0F",X"C2",X"10",X"A7",X"11",X"85",X"12",X"59",X"13",X"26",X"14",X"EC",X"14",
		X"AA",X"15",X"60",X"16",X"10",X"17",X"B9",X"17",X"5D",X"18",X"F9",X"18",X"91",X"19",X"22",X"1A",
		X"AC",X"1A",X"32",X"1B",X"B2",X"1B",X"22",X"1C",X"EA",X"1B",X"FD",X"1A",X"A7",X"19",X"06",X"18",
		X"3D",X"16",X"58",X"14",X"6D",X"12",X"7C",X"10",X"8F",X"0E",X"A9",X"0C",X"CD",X"0A",X"FC",X"08",
		X"39",X"07",X"83",X"05",X"D8",X"03",X"3C",X"02",X"AC",X"00",X"2A",X"FF",X"B6",X"FD",X"4B",X"FC",
		X"EF",X"FA",X"9D",X"F9",X"57",X"F8",X"1D",X"F7",X"ED",X"F5",X"C8",X"F4",X"AD",X"F3",X"9B",X"F2",
		X"94",X"F1",X"96",X"F0",X"A0",X"EF",X"B5",X"EE",X"D0",X"ED",X"F5",X"EC",X"20",X"EC",X"55",X"EB",
		X"91",X"EA",X"D4",X"E9",X"1E",X"E9",X"6E",X"E8",X"C7",X"E7",X"24",X"E7",X"87",X"E6",X"F2",X"E5",
		X"63",X"E5",X"D9",X"E4",X"55",X"E4",X"D4",X"E3",X"5A",X"E3",X"E4",X"E2",X"75",X"E2",X"09",X"E2",
		X"A1",X"E1",X"41",X"E1",X"E2",X"E0",X"1C",X"E1",X"0B",X"E2",X"67",X"E3",X"11",X"E5",X"E2",X"E6",
		X"CE",X"E8",X"C5",X"EA",X"BE",X"EC",X"B6",X"EE",X"A6",X"F0",X"8C",X"F2",X"68",X"F4",X"33",X"F6",
		X"F4",X"F7",X"A8",X"F9",X"4E",X"FB",X"E5",X"FC",X"71",X"FE",X"EF",X"FF",X"5F",X"01",X"C4",X"02",
		X"1E",X"04",X"6B",X"05",X"AD",X"06",X"E4",X"07",X"10",X"09",X"33",X"0A",X"4A",X"0B",X"57",X"0C",
		X"5C",X"0D",X"57",X"0E",X"4A",X"0F",X"33",X"10",X"15",X"11",X"EE",X"11",X"C0",X"12",X"8A",X"13",
		X"4B",X"14",X"06",X"15",X"B9",X"15",X"66",X"16",X"0F",X"17",X"AE",X"17",X"48",X"18",X"DE",X"18",
		X"6B",X"19",X"F5",X"19",X"78",X"1A",X"F6",X"1A",X"6E",X"1B",X"E2",X"1B",X"52",X"1C",X"BC",X"1C",
		X"23",X"1D",X"83",X"1D",X"E2",X"1D",X"3A",X"1E",X"8F",X"1E",X"E3",X"1E",X"2F",X"1F",X"79",X"1F",
		X"C1",X"1F",X"03",X"20",X"44",X"20",X"81",X"20",X"BB",X"20",X"F1",X"20",X"25",X"21",X"55",X"21",
		X"84",X"21",X"B0",X"21",X"DA",X"21",X"00",X"22",X"24",X"22",X"46",X"22",X"65",X"22",X"83",X"22",
		X"9E",X"22",X"B7",X"22",X"CF",X"22",X"E5",X"22",X"F8",X"22",X"0A",X"23",X"1A",X"23",X"28",X"23",
		X"35",X"23",X"41",X"23",X"4B",X"23",X"53",X"23",X"58",X"23",X"5E",X"23",X"63",X"23",X"67",X"23",
		X"68",X"23",X"66",X"23",X"67",X"23",X"65",X"23",X"63",X"23",X"5E",X"23",X"58",X"23",X"53",X"23",
		X"4C",X"23",X"44",X"23",X"3C",X"23",X"30",X"23",X"27",X"23",X"1B",X"23",X"10",X"23",X"01",X"23",
		X"FA",X"22",X"90",X"22",X"6A",X"21",X"D5",X"1F",X"F2",X"1D",X"E4",X"1B",X"BC",X"19",X"8A",X"17",
		X"54",X"15",X"24",X"13",X"FB",X"10",X"DF",X"0E",X"CF",X"0C",X"CE",X"0A",X"DB",X"08",X"F8",X"06",
		X"22",X"05",X"5E",X"03",X"A6",X"01",X"FE",X"FF",X"63",X"FE",X"D7",X"FC",X"58",X"FB",X"E4",X"F9",
		X"7F",X"F8",X"25",X"F7",X"D7",X"F5",X"94",X"F4",X"5E",X"F3",X"31",X"F2",X"10",X"F1",X"F8",X"EF",
		X"E9",X"EE",X"E5",X"ED",X"EB",X"EC",X"F9",X"EB",X"10",X"EB",X"30",X"EA",X"57",X"E9",X"85",X"E8",
		X"BF",X"E7",X"FD",X"E6",X"43",X"E6",X"8E",X"E5",X"E3",X"E4",X"3E",X"E4",X"9E",X"E3",X"06",X"E3",
		X"73",X"E2",X"E6",X"E1",X"60",X"E1",X"DC",X"E0",X"62",X"E0",X"E8",X"DF",X"78",X"DF",X"06",X"DF",
		X"E1",X"DE",X"79",X"DF",X"8C",X"E0",X"F1",X"E1",X"87",X"E3",X"3E",X"E5",X"01",X"E7",X"CD",X"E8",
		X"97",X"EA",X"5D",X"EC",X"1B",X"EE",X"CE",X"EF",X"76",X"F1",X"15",X"F3",X"A4",X"F4",X"2A",X"F6",
		X"A2",X"F7",X"10",X"F9",X"71",X"FA",X"C8",X"FB",X"11",X"FD",X"51",X"FE",X"85",X"FF",X"AE",X"00",
		X"CD",X"01",X"E4",X"02",X"F0",X"03",X"F5",X"04",X"F0",X"05",X"E1",X"06",X"CB",X"07",X"AC",X"08",
		X"85",X"09",X"59",X"0A",X"22",X"0B",X"E5",X"0B",X"A2",X"0C",X"57",X"0D",X"05",X"0E",X"AF",X"0E",
		X"50",X"0F",X"ED",X"0F",X"83",X"10",X"15",X"11",X"9E",X"11",X"27",X"12",X"A5",X"12",X"26",X"13",
		X"97",X"13",X"17",X"14",X"B2",X"14",X"18",X"15",X"81",X"15",X"E1",X"15",X"40",X"16",X"9A",X"16",
		X"F1",X"16",X"42",X"17",X"92",X"17",X"DD",X"17",X"25",X"18",X"6B",X"18",X"AD",X"18",X"EB",X"18",
		X"27",X"19",X"5F",X"19",X"97",X"19",X"CA",X"19",X"FB",X"19",X"29",X"1A",X"55",X"1A",X"7F",X"1A",
		X"A5",X"1A",X"CC",X"1A",X"EF",X"1A",X"10",X"1B",X"2E",X"1B",X"4B",X"1B",X"67",X"1B",X"7F",X"1B",
		X"97",X"1B",X"AD",X"1B",X"C0",X"1B",X"D3",X"1B",X"E5",X"1B",X"F3",X"1B",X"00",X"1C",X"0D",X"1C",
		X"19",X"1C",X"23",X"1C",X"2C",X"1C",X"31",X"1C",X"39",X"1C",X"3D",X"1C",X"40",X"1C",X"43",X"1C",
		X"46",X"1C",X"47",X"1C",X"46",X"1C",X"45",X"1C",X"42",X"1C",X"40",X"1C",X"3C",X"1C",X"37",X"1C",
		X"32",X"1C",X"2B",X"1C",X"24",X"1C",X"1B",X"1C",X"14",X"1C",X"0B",X"1C",X"01",X"1C",X"F6",X"1B",
		X"EB",X"1B",X"DF",X"1B",X"D3",X"1B",X"C6",X"1B",X"B9",X"1B",X"AC",X"1B",X"9D",X"1B",X"8F",X"1B",
		X"80",X"1B",X"6F",X"1B",X"60",X"1B",X"4F",X"1B",X"3F",X"1B",X"2D",X"1B",X"1C",X"1B",X"0A",X"1B",
		X"F8",X"1A",X"E6",X"1A",X"D2",X"1A",X"C0",X"1A",X"AD",X"1A",X"98",X"1A",X"84",X"1A",X"70",X"1A",
		X"5E",X"1A",X"34",X"1A",X"6C",X"19",X"16",X"18",X"6B",X"16",X"8A",X"14",X"8B",X"12",X"7C",X"10",
		X"68",X"0E",X"57",X"0C",X"4B",X"0A",X"4A",X"08",X"53",X"06",X"6B",X"04",X"91",X"02",X"C4",X"00",
		X"06",X"FF",X"56",X"FD",X"B5",X"FB",X"21",X"FA",X"9A",X"F8",X"20",X"F7",X"B4",X"F5",X"52",X"F4",
		X"FF",X"F2",X"B6",X"F1",X"7A",X"F0",X"49",X"EF",X"20",X"EE",X"04",X"ED",X"F1",X"EB",X"E8",X"EA",
		X"EA",X"E9",X"F4",X"E8",X"07",X"E8",X"22",X"E7",X"47",X"E6",X"73",X"E5",X"A7",X"E4",X"E2",X"E3",
		X"25",X"E3",X"6F",X"E2",X"C3",X"E1",X"19",X"E1",X"7A",X"E0",X"DE",X"DF",X"48",X"DF",X"B9",X"DE",
		X"31",X"DE",X"AD",X"DD",X"30",X"DD",X"B7",X"DC",X"43",X"DC",X"D5",X"DB",X"6B",X"DB",X"06",X"DB",
		X"B0",X"DA",X"ED",X"DA",X"C2",X"DB",X"EF",X"DC",X"5C",X"DE",X"EA",X"DF",X"8F",X"E1",X"3C",X"E3",
		X"EC",X"E4",X"97",X"E6",X"3E",X"E8",X"DC",X"E9",X"72",X"EB",X"FB",X"EC",X"7B",X"EE",X"ED",X"EF",
		X"55",X"F1",X"B3",X"F2",X"05",X"F4",X"4B",X"F5",X"87",X"F6",X"BA",X"F7",X"E2",X"F8",X"00",X"FA",
		X"16",X"FB",X"22",X"FC",X"24",X"FD",X"1F",X"FE",X"10",X"FF",X"F9",X"FF",X"D9",X"00",X"B3",X"01",
		X"87",X"02",X"51",X"03",X"14",X"04",X"D2",X"04",X"88",X"05",X"39",X"06",X"E3",X"06",X"88",X"07",
		X"24",X"08",X"BD",X"08",X"51",X"09",X"DE",X"09",X"67",X"0A",X"EA",X"0A",X"69",X"0B",X"E3",X"0B",
		X"59",X"0C",X"CA",X"0C",X"34",X"0D",X"9F",X"0D",X"03",X"0E",X"64",X"0E",X"C0",X"0E",X"16",X"0F",
		X"EC",X"0E",X"26",X"0E",X"05",X"0D",X"A4",X"0B",X"20",X"0A",X"86",X"08",X"E4",X"06",X"3D",X"05",
		X"9B",X"03",X"FD",X"01",X"6A",X"00",X"E0",X"FE",X"60",X"FD",X"ED",X"FB",X"83",X"FA",X"24",X"F9",
		X"D3",X"F7",X"8C",X"F6",X"50",X"F5",X"1E",X"F4",X"F8",X"F2",X"DB",X"F1",X"C9",X"F0",X"C1",X"EF",
		X"C0",X"EE",X"CB",X"ED",X"D9",X"EC",X"1B",X"EC",X"09",X"EC",X"72",X"EC",X"30",X"ED",X"21",X"EE",
		X"35",X"EF",X"5B",X"F0",X"8C",X"F1",X"BF",X"F2",X"F5",X"F3",X"24",X"F5",X"4E",X"F6",X"72",X"F7",
		X"8F",X"F8",X"A3",X"F9",X"B1",X"FA",X"B5",X"FB",X"AF",X"FC",X"A3",X"FD",X"90",X"FE",X"72",X"FF",
		X"50",X"00",X"22",X"01",X"F2",X"01",X"B6",X"02",X"78",X"03",X"30",X"04",X"E6",X"04",X"29",X"05",
		X"CC",X"04",X"0F",X"04",X"0E",X"03",X"E6",X"01",X"A1",X"00",X"53",X"FF",X"FF",X"FD",X"AB",X"FC",
		X"5A",X"FB",X"10",X"FA",X"CE",X"F8",X"93",X"F7",X"60",X"F6",X"38",X"F5",X"19",X"F4",X"04",X"F3",
		X"F8",X"F1",X"F6",X"F0",X"FB",X"EF",X"09",X"EF",X"20",X"EE",X"3F",X"ED",X"68",X"EC",X"97",X"EB",
		X"D0",X"EA",X"0B",X"EA",X"69",X"E9",X"66",X"E9",X"E7",X"E9",X"B9",X"EA",X"C1",X"EB",X"EA",X"EC",
		X"28",X"EE",X"6F",X"EF",X"BB",X"F0",X"04",X"F2",X"4A",X"F3",X"8B",X"F4",X"C1",X"F5",X"F0",X"F6",
		X"18",X"F8",X"36",X"F9",X"4E",X"FA",X"5A",X"FB",X"60",X"FC",X"5A",X"FD",X"50",X"FE",X"3C",X"FF",
		X"1E",X"00",X"F9",X"00",X"CF",X"01",X"9B",X"02",X"61",X"03",X"20",X"04",X"DA",X"04",X"8B",X"05",
		X"38",X"06",X"DE",X"06",X"7E",X"07",X"19",X"08",X"AD",X"08",X"3C",X"09",X"C8",X"09",X"4C",X"0A",
		X"CD",X"0A",X"49",X"0B",X"C0",X"0B",X"34",X"0C",X"A1",X"0C",X"0B",X"0D",X"71",X"0D",X"D3",X"0D",
		X"32",X"0E",X"8C",X"0E",X"E3",X"0E",X"38",X"0F",X"87",X"0F",X"D3",X"0F",X"1F",X"10",X"65",X"10",
		X"AA",X"10",X"DE",X"10",X"84",X"10",X"A6",X"0F",X"77",X"0E",X"15",X"0D",X"92",X"0B",X"FE",X"09",
		X"63",X"08",X"CA",X"06",X"32",X"05",X"A2",X"03",X"1B",X"02",X"9D",X"00",X"2A",X"FF",X"C2",X"FD",
		X"64",X"FC",X"12",X"FB",X"CB",X"F9",X"8E",X"F8",X"5E",X"F7",X"36",X"F6",X"18",X"F5",X"06",X"F4",
		X"FC",X"F2",X"FB",X"F1",X"05",X"F1",X"15",X"F0",X"31",X"EF",X"51",X"EE",X"7C",X"ED",X"AE",X"EC",
		X"E7",X"EB",X"28",X"EB",X"71",X"EA",X"BF",X"E9",X"14",X"E9",X"70",X"E8",X"D2",X"E7",X"3A",X"E7",
		X"A9",X"E6",X"1C",X"E6",X"96",X"E5",X"14",X"E5",X"98",X"E4",X"20",X"E4",X"AD",X"E3",X"42",X"E3",
		X"D8",X"E2",X"74",X"E2",X"14",X"E2",X"B7",X"E1",X"5F",X"E1",X"0B",X"E1",X"BB",X"E0",X"6D",X"E0",
		X"2A",X"E0",X"64",X"E0",X"29",X"E1",X"40",X"E2",X"8F",X"E3",X"FF",X"E4",X"82",X"E6",X"0A",X"E8",
		X"99",X"E9",X"23",X"EB",X"A7",X"EC",X"24",X"EE",X"99",X"EF",X"02",X"F1",X"62",X"F2",X"B5",X"F3",
		X"02",X"F5",X"41",X"F6",X"79",X"F7",X"A5",X"F8",X"C7",X"F9",X"DF",X"FA",X"F1",X"FB",X"F7",X"FC",
		X"F5",X"FD",X"EA",X"FE",X"D7",X"FF",X"BB",X"00",X"99",X"01",X"70",X"02",X"3E",X"03",X"05",X"04",
		X"C5",X"04",X"80",X"05",X"33",X"06",X"E0",X"06",X"89",X"07",X"27",X"08",X"C2",X"08",X"59",X"09",
		X"E9",X"09",X"74",X"0A",X"FB",X"0A",X"7C",X"0B",X"FA",X"0B",X"6F",X"0C",X"E4",X"0C",X"51",X"0D",
		X"BE",X"0D",X"20",X"0E",X"8F",X"0E",X"0D",X"0F",X"66",X"0F",X"C0",X"0F",X"14",X"10",X"68",X"10",
		X"B4",X"10",X"01",X"11",X"47",X"11",X"8D",X"11",X"CD",X"11",X"0E",X"12",X"4A",X"12",X"83",X"12",
		X"BA",X"12",X"EE",X"12",X"22",X"13",X"51",X"13",X"7F",X"13",X"AA",X"13",X"D3",X"13",X"FA",X"13",
		X"20",X"14",X"42",X"14",X"65",X"14",X"83",X"14",X"A2",X"14",X"BD",X"14",X"D8",X"14",X"F0",X"14",
		X"0A",X"15",X"1B",X"15",X"36",X"15",X"ED",X"14",X"17",X"14",X"EC",X"12",X"83",X"11",X"F9",X"0F",
		X"5B",X"0E",X"B5",X"0C",X"0E",X"0B",X"6B",X"09",X"CC",X"07",X"38",X"06",X"AC",X"04",X"2E",X"03",
		X"B7",X"01",X"4F",X"00",X"F1",X"FE",X"A0",X"FD",X"57",X"FC",X"1A",X"FB",X"E8",X"F9",X"C1",X"F8",
		X"A1",X"F7",X"8E",X"F6",X"83",X"F5",X"82",X"F4",X"89",X"F3",X"99",X"F2",X"B3",X"F1",X"D3",X"F0",
		X"FE",X"EF",X"2F",X"EF",X"66",X"EE",X"A7",X"ED",X"EE",X"EC",X"3B",X"EC",X"8F",X"EB",X"EA",X"EA",
		X"4A",X"EA",X"B1",X"E9",X"1F",X"E9",X"90",X"E8",X"08",X"E8",X"84",X"E7",X"08",X"E7",X"8F",X"E6",
		X"1D",X"E6",X"AD",X"E5",X"44",X"E5",X"DB",X"E4",X"7C",X"E4",X"1C",X"E4",X"C4",X"E3",X"6D",X"E3",
		X"1D",X"E3",X"CB",X"E2",X"C4",X"E2",X"53",X"E3",X"3A",X"E4",X"63",X"E5",X"AD",X"E6",X"12",X"E8",
		X"7F",X"E9",X"F1",X"EA",X"62",X"EC",X"CF",X"ED",X"35",X"EF",X"93",X"F0",X"E7",X"F1",X"33",X"F3",
		X"76",X"F4",X"AE",X"F5",X"DC",X"F6",X"01",X"F8",X"1E",X"F9",X"2F",X"FA",X"38",X"FB",X"39",X"FC",
		X"31",X"FD",X"22",X"FE",X"0A",X"FF",X"E9",X"FF",X"C1",X"00",X"89",X"01",X"CE",X"01",X"94",X"01",
		X"0C",X"01",X"4E",X"00",X"6F",X"FF",X"7B",X"FE",X"7F",X"FD",X"7C",X"FC",X"7A",X"FB",X"79",X"FA",
		X"7F",X"F9",X"87",X"F8",X"99",X"F7",X"AF",X"F6",X"CD",X"F5",X"F5",X"F4",X"22",X"F4",X"55",X"F3",
		X"91",X"F2",X"D4",X"F1",X"1E",X"F1",X"6C",X"F0",X"C2",X"EF",X"1E",X"EF",X"81",X"EE",X"E9",X"ED",
		X"56",X"ED",X"C8",X"EC",X"43",X"EC",X"C0",X"EB",X"43",X"EB",X"CB",X"EA",X"58",X"EA",X"E9",X"E9",
		X"7F",X"E9",X"19",X"E9",X"B8",X"E8",X"59",X"E8",X"00",X"E8",X"A8",X"E7",X"55",X"E7",X"08",X"E7",
		X"BC",X"E6",X"74",X"E6",X"2F",X"E6",X"ED",X"E5",X"B0",X"E5",X"74",X"E5",X"3B",X"E5",X"06",X"E5",
		X"D2",X"E4",X"A2",X"E4",X"73",X"E4",X"47",X"E4",X"1F",X"E4",X"F6",X"E3",X"D2",X"E3",X"AF",X"E3",
		X"8F",X"E3",X"72",X"E3",X"55",X"E3",X"39",X"E3",X"21",X"E3",X"0B",X"E3",X"F5",X"E2",X"E0",X"E2",
		X"CE",X"E2",X"BF",X"E2",X"AF",X"E2",X"A3",X"E2",X"97",X"E2",X"8C",X"E2",X"83",X"E2",X"7A",X"E2",
		X"73",X"E2",X"6E",X"E2",X"69",X"E2",X"64",X"E2",X"64",X"E2",X"62",X"E2",X"62",X"E2",X"64",X"E2",
		X"65",X"E2",X"68",X"E2",X"6A",X"E2",X"6F",X"E2",X"75",X"E2",X"7B",X"E2",X"82",X"E2",X"89",X"E2",
		X"92",X"E2",X"9B",X"E2",X"A5",X"E2",X"AD",X"E2",X"B9",X"E2",X"C5",X"E2",X"D1",X"E2",X"DD",X"E2",
		X"EB",X"E2",X"F8",X"E2",X"06",X"E3",X"18",X"E3",X"25",X"E3",X"35",X"E3",X"45",X"E3",X"55",X"E3",
		X"66",X"E3",X"78",X"E3",X"89",X"E3",X"9C",X"E3",X"AD",X"E3",X"C0",X"E3",X"D4",X"E3",X"E8",X"E3",
		X"FC",X"E3",X"0F",X"E4",X"23",X"E4",X"38",X"E4",X"4C",X"E4",X"62",X"E4",X"78",X"E4",X"8C",X"E4",
		X"A1",X"E4",X"B8",X"E4",X"CE",X"E4",X"E4",X"E4",X"FC",X"E4",X"12",X"E5",X"28",X"E5",X"3F",X"E5",
		X"57",X"E5",X"6E",X"E5",X"86",X"E5",X"9C",X"E5",X"B4",X"E5",X"CC",X"E5",X"E4",X"E5",X"FA",X"E5",
		X"14",X"E6",X"2C",X"E6",X"44",X"E6",X"5D",X"E6",X"74",X"E6",X"8E",X"E6",X"A5",X"E6",X"BE",X"E6",
		X"D7",X"E6",X"F0",X"E6",X"08",X"E7",X"20",X"E7",X"39",X"E7",X"53",X"E7",X"6B",X"E7",X"84",X"E7",
		X"9B",X"E7",X"B6",X"E7",X"CF",X"E7",X"E8",X"E7",X"00",X"E8",X"1B",X"E8",X"33",X"E8",X"4D",X"E8",
		X"63",X"E8",X"7F",X"E8",X"94",X"E8",X"F4",X"E8",X"D4",X"E9",X"02",X"EB",X"67",X"EC",X"E7",X"ED",
		X"79",X"EF",X"12",X"F1",X"AC",X"F2",X"42",X"F4",X"D0",X"F5",X"5A",X"F7",X"D5",X"F8",X"47",X"FA",
		X"B0",X"FB",X"0B",X"FD",X"60",X"FE",X"A6",X"FF",X"E3",X"00",X"14",X"02",X"3D",X"03",X"5C",X"04",
		X"71",X"05",X"7B",X"06",X"7E",X"07",X"77",X"08",X"65",X"09",X"51",X"0A",X"24",X"0B",X"7B",X"0B",
		X"5E",X"0B",X"FE",X"0A",X"6A",X"0A",X"B9",X"09",X"F6",X"08",X"29",X"08",X"58",X"07",X"83",X"06",
		X"B1",X"05",X"E2",X"04",X"16",X"04",X"50",X"03",X"8F",X"02",X"D5",X"01",X"20",X"01",X"6F",X"00",
		X"C8",X"FF",X"24",X"FF",X"84",X"FE",X"EC",X"FD",X"57",X"FD",X"C9",X"FC",X"3F",X"FC",X"BB",X"FB",
		X"3A",X"FB",X"BE",X"FA",X"47",X"FA",X"D5",X"F9",X"66",X"F9",X"FB",X"F8",X"95",X"F8",X"33",X"F8",
		X"D2",X"F7",X"77",X"F7",X"1E",X"F7",X"CA",X"F6",X"79",X"F6",X"29",X"F6",X"DF",X"F5",X"97",X"F5",
		X"51",X"F5",X"10",X"F5",X"CF",X"F4",X"91",X"F4",X"57",X"F4",X"1E",X"F4",X"E8",X"F3",X"B4",X"F3",
		X"83",X"F3",X"55",X"F3",X"27",X"F3",X"FC",X"F2",X"D4",X"F2",X"B0",X"F2",X"F8",X"F2",X"B1",X"F3",
		X"AB",X"F4",X"D2",X"F5",X"14",X"F7",X"63",X"F8",X"B8",X"F9",X"10",X"FB",X"63",X"FC",X"B1",X"FD",
		X"F7",X"FE",X"35",X"00",X"6A",X"01",X"96",X"02",X"BA",X"03",X"D3",X"04",X"E3",X"05",X"EC",X"06",
		X"EA",X"07",X"E1",X"08",X"CE",X"09",X"B5",X"0A",X"92",X"0B",X"69",X"0C",X"35",X"0D",X"FD",X"0D",
		X"BE",X"0E",X"75",X"0F",X"29",X"10",X"D4",X"10",X"7A",X"11",X"19",X"12",X"B4",X"12",X"47",X"13",
		X"D5",X"13",X"5F",X"14",X"E4",X"14",X"62",X"15",X"DC",X"15",X"51",X"16",X"C2",X"16",X"2D",X"17",
		X"96",X"17",X"F7",X"17",X"59",X"18",X"B4",X"18",X"0C",X"19",X"61",X"19",X"B0",X"19",X"FD",X"19",
		X"45",X"1A",X"8D",X"1A",X"D0",X"1A",X"10",X"1B",X"4E",X"1B",X"88",X"1B",X"BF",X"1B",X"F6",X"1B",
		X"25",X"1C",X"57",X"1C",X"83",X"1C",X"AF",X"1C",X"D6",X"1C",X"FD",X"1C",X"20",X"1D",X"44",X"1D",
		X"63",X"1D",X"82",X"1D",X"9E",X"1D",X"B9",X"1D",X"CF",X"1D",X"E9",X"1D",X"FC",X"1D",X"13",X"1E",
		X"20",X"1E",X"37",X"1E",X"3C",X"1E",X"62",X"1E",X"AD",X"1E",X"B3",X"1E",X"BE",X"1E",X"C8",X"1E",
		X"B7",X"1E",X"2B",X"1E",X"46",X"1D",X"28",X"1C",X"E3",X"1A",X"8C",X"19",X"2B",X"18",X"C5",X"16",
		X"60",X"15",X"01",X"14",X"A6",X"12",X"54",X"11",X"0B",X"10",X"CB",X"0E",X"94",X"0D",X"66",X"0C",
		X"43",X"0B",X"28",X"0A",X"15",X"09",X"0C",X"08",X"0C",X"07",X"15",X"06",X"24",X"05",X"3C",X"04",
		X"5C",X"03",X"83",X"02",X"B3",X"01",X"E8",X"00",X"25",X"00",X"69",X"FF",X"B4",X"FE",X"03",X"FE",
		X"59",X"FD",X"B5",X"FC",X"16",X"FC",X"7F",X"FB",X"EC",X"FA",X"5E",X"FA",X"D4",X"F9",X"50",X"F9",
		X"D0",X"F8",X"56",X"F8",X"E0",X"F7",X"6D",X"F7",X"01",X"F7",X"96",X"F6",X"30",X"F6",X"CE",X"F5",
		X"70",X"F5",X"15",X"F5",X"BE",X"F4",X"6B",X"F4",X"1B",X"F4",X"CD",X"F3",X"83",X"F3",X"3C",X"F3",
		X"F8",X"F2",X"B7",X"F2",X"78",X"F2",X"3B",X"F2",X"01",X"F2",X"CB",X"F1",X"95",X"F1",X"64",X"F1",
		X"33",X"F1",X"05",X"F1",X"D9",X"F0",X"AF",X"F0",X"87",X"F0",X"61",X"F0",X"3D",X"F0",X"1C",X"F0",
		X"FB",X"EF",X"DC",X"EF",X"BF",X"EF",X"A4",X"EF",X"89",X"EF",X"71",X"EF",X"58",X"EF",X"44",X"EF",
		X"30",X"EF",X"1C",X"EF",X"0C",X"EF",X"FA",X"EE",X"EB",X"EE",X"DD",X"EE",X"D0",X"EE",X"C5",X"EE",
		X"BA",X"EE",X"AF",X"EE",X"A7",X"EE",X"9D",X"EE",X"97",X"EE",X"91",X"EE",X"8B",X"EE",X"86",X"EE",
		X"84",X"EE",X"80",X"EE",X"7E",X"EE",X"7C",X"EE",X"7D",X"EE",X"7C",X"EE",X"7D",X"EE",X"7E",X"EE",
		X"81",X"EE",X"81",X"EE",X"87",X"EE",X"89",X"EE",X"8F",X"EE",X"8F",X"EE",X"BF",X"EE",X"64",X"EF",
		X"54",X"F0",X"76",X"F1",X"B4",X"F2",X"05",X"F4",X"5A",X"F5",X"B4",X"F6",X"0B",X"F8",X"5C",X"F9",
		X"A8",X"FA",X"EA",X"FB",X"25",X"FD",X"54",X"FE",X"7D",X"FF",X"9C",X"00",X"B1",X"01",X"BE",X"02",
		X"C1",X"03",X"BC",X"04",X"AE",X"05",X"98",X"06",X"7B",X"07",X"55",X"08",X"28",X"09",X"F3",X"09",
		X"B8",X"0A",X"74",X"0B",X"2D",X"0C",X"DC",X"0C",X"85",X"0D",X"2A",X"0E",X"CA",X"0E",X"60",X"0F",
		X"F4",X"0F",X"80",X"10",X"09",X"11",X"8C",X"11",X"08",X"12",X"83",X"12",X"F8",X"12",X"67",X"13",
		X"D2",X"13",X"3A",X"14",X"9E",X"14",X"FD",X"14",X"59",X"15",X"B1",X"15",X"03",X"16",X"56",X"16",
		X"A3",X"16",X"EE",X"16",X"35",X"17",X"79",X"17",X"BA",X"17",X"F7",X"17",X"34",X"18",X"6C",X"18",
		X"A1",X"18",X"D6",X"18",X"04",X"19",X"34",X"19",X"60",X"19",X"89",X"19",X"B2",X"19",X"D7",X"19",
		X"FA",X"19",X"1C",X"1A",X"3B",X"1A",X"59",X"1A",X"75",X"1A",X"90",X"1A",X"A8",X"1A",X"BF",X"1A",
		X"D4",X"1A",X"E9",X"1A",X"FA",X"1A",X"0C",X"1B",X"1B",X"1B",X"29",X"1B",X"37",X"1B",X"40",X"1B",
		X"4C",X"1B",X"54",X"1B",X"5C",X"1B",X"64",X"1B",X"6A",X"1B",X"6E",X"1B",X"73",X"1B",X"77",X"1B",
		X"77",X"1B",X"77",X"1B",X"79",X"1B",X"77",X"1B",X"75",X"1B",X"73",X"1B",X"70",X"1B",X"6E",X"1B",
		X"67",X"1B",X"62",X"1B",X"5C",X"1B",X"56",X"1B",X"4F",X"1B",X"46",X"1B",X"3C",X"1B",X"34",X"1B",
		X"2B",X"1B",X"21",X"1B",X"18",X"1B",X"0C",X"1B",X"01",X"1B",X"F5",X"1A",X"E8",X"1A",X"DD",X"1A",
		X"CE",X"1A",X"C0",X"1A",X"B3",X"1A",X"A5",X"1A",X"96",X"1A",X"87",X"1A",X"78",X"1A",X"68",X"1A",
		X"59",X"1A",X"47",X"1A",X"37",X"1A",X"27",X"1A",X"15",X"1A",X"04",X"1A",X"F2",X"19",X"E1",X"19",
		X"CE",X"19",X"BD",X"19",X"A9",X"19",X"98",X"19",X"84",X"19",X"73",X"19",X"5C",X"19",X"4D",X"19",
		X"FF",X"18",X"47",X"18",X"51",X"17",X"31",X"16",X"F9",X"14",X"B3",X"13",X"69",X"12",X"1D",X"11",
		X"D4",X"0F",X"91",X"0E",X"54",X"0D",X"1E",X"0C",X"F2",X"0A",X"CE",X"09",X"B1",X"08",X"A0",X"07",
		X"97",X"06",X"93",X"05",X"9C",X"04",X"AA",X"03",X"C2",X"02",X"E1",X"01",X"08",X"01",X"36",X"00",
		X"6A",X"FF",X"A7",X"FE",X"E9",X"FD",X"33",X"FD",X"82",X"FC",X"D7",X"FB",X"33",X"FB",X"95",X"FA",
		X"FB",X"F9",X"68",X"F9",X"D8",X"F8",X"4F",X"F8",X"CB",X"F7",X"4B",X"F7",X"D1",X"F6",X"59",X"F6",
		X"E7",X"F5",X"7B",X"F5",X"10",X"F5",X"AB",X"F4",X"48",X"F4",X"EB",X"F3",X"8E",X"F3",X"37",X"F3",
		X"E5",X"F2",X"94",X"F2",X"46",X"F2",X"FD",X"F1",X"B4",X"F1",X"72",X"F1",X"2D",X"F1",X"1A",X"F1",
		X"73",X"F1",X"0E",X"F2",X"D7",X"F2",X"BB",X"F3",X"B0",X"F4",X"AC",X"F5",X"AD",X"F6",X"AE",X"F7",
		X"AB",X"F8",X"A3",X"F9",X"96",X"FA",X"83",X"FB",X"67",X"FC",X"47",X"FD",X"20",X"FE",X"F0",X"FE",
		X"BC",X"FF",X"7E",X"00",X"3C",X"01",X"F3",X"01",X"A3",X"02",X"4F",X"03",X"F4",X"03",X"93",X"04",
		X"2C",X"05",X"C2",X"05",X"4C",X"06",X"7D",X"06",X"51",X"06",X"EB",X"05",X"5F",X"05",X"BB",X"04",
		X"09",X"04",X"4E",X"03",X"91",X"02",X"D5",X"01",X"18",X"01",X"60",X"00",X"AC",X"FF",X"FD",X"FE",
		X"52",X"FE",X"AD",X"FD",X"0C",X"FD",X"70",X"FC",X"DD",X"FB",X"4C",X"FB",X"BE",X"FA",X"37",X"FA",
		X"B4",X"F9",X"39",X"F9",X"BF",X"F8",X"49",X"F8",X"DB",X"F7",X"6F",X"F7",X"05",X"F7",X"A2",X"F6",
		X"40",X"F6",X"E3",X"F5",X"89",X"F5",X"33",X"F5",X"DF",X"F4",X"91",X"F4",X"44",X"F4",X"FB",X"F3",
		X"B5",X"F3",X"70",X"F3",X"30",X"F3",X"F2",X"F2",X"B6",X"F2",X"7D",X"F2",X"46",X"F2",X"11",X"F2",
		X"E0",X"F1",X"B0",X"F1",X"81",X"F1",X"57",X"F1",X"2D",X"F1",X"06",X"F1",X"E0",X"F0",X"BC",X"F0",
		X"98",X"F0",X"77",X"F0",X"59",X"F0",X"3E",X"F0",X"20",X"F0",X"07",X"F0",X"ED",X"EF",X"D6",X"EF",
		X"C2",X"EF",X"AD",X"EF",X"98",X"EF",X"87",X"EF",X"77",X"EF",X"67",X"EF",X"59",X"EF",X"4B",X"EF",
		X"3E",X"EF",X"34",X"EF",X"28",X"EF",X"20",X"EF",X"17",X"EF",X"0F",X"EF",X"0A",X"EF",X"03",X"EF",
		X"FE",X"EE",X"F9",X"EE",X"F6",X"EE",X"F5",X"EE",X"F2",X"EE",X"EF",X"EE",X"EF",X"EE",X"F0",X"EE",
		X"F1",X"EE",X"F1",X"EE",X"F4",X"EE",X"F7",X"EE",X"FA",X"EE",X"FC",X"EE",X"01",X"EF",X"04",X"EF",
		X"0B",X"EF",X"10",X"EF",X"17",X"EF",X"1C",X"EF",X"24",X"EF",X"2B",X"EF",X"31",X"EF",X"39",X"EF",
		X"42",X"EF",X"4A",X"EF",X"53",X"EF",X"5D",X"EF",X"66",X"EF",X"6F",X"EF",X"7A",X"EF",X"83",X"EF",
		X"91",X"EF",X"BB",X"EF",X"4B",X"F0",X"2B",X"F1",X"25",X"F2",X"3D",X"F3",X"5B",X"F4",X"82",X"F5",
		X"A5",X"F6",X"C8",X"F7",X"E6",X"F8",X"FE",X"F9",X"0F",X"FB",X"15",X"FC",X"18",X"FD",X"12",X"FE",
		X"03",X"FF",X"ED",X"FF",X"D0",X"00",X"A9",X"01",X"7E",X"02",X"4A",X"03",X"0F",X"04",X"CD",X"04",
		X"86",X"05",X"38",X"06",X"E6",X"06",X"89",X"07",X"2A",X"08",X"C5",X"08",X"59",X"09",X"EA",X"09",
		X"74",X"0A",X"F9",X"0A",X"7B",X"0B",X"F6",X"0B",X"6E",X"0C",X"E1",X"0C",X"50",X"0D",X"BA",X"0D",
		X"21",X"0E",X"84",X"0E",X"E2",X"0E",X"3F",X"0F",X"96",X"0F",X"EC",X"0F",X"3C",X"10",X"8A",X"10",
		X"D5",X"10",X"1D",X"11",X"60",X"11",X"A3",X"11",X"E1",X"11",X"1E",X"12",X"59",X"12",X"90",X"12",
		X"C5",X"12",X"F8",X"12",X"28",X"13",X"57",X"13",X"83",X"13",X"AB",X"13",X"D4",X"13",X"F9",X"13",
		X"1D",X"14",X"40",X"14",X"60",X"14",X"80",X"14",X"9C",X"14",X"B7",X"14",X"D1",X"14",X"E9",X"14",
		X"02",X"15",X"16",X"15",X"2A",X"15",X"3C",X"15",X"4F",X"15",X"5F",X"15",X"6D",X"15",X"7B",X"15",
		X"88",X"15",X"95",X"15",X"9E",X"15",X"A9",X"15",X"B1",X"15",X"B8",X"15",X"BE",X"15",X"C5",X"15",
		X"CA",X"15",X"CD",X"15",X"D0",X"15",X"D3",X"15",X"D5",X"15",X"D6",X"15",X"D7",X"15",X"D7",X"15",
		X"D4",X"15",X"D4",X"15",X"D0",X"15",X"CD",X"15",X"CA",X"15",X"C6",X"15",X"C1",X"15",X"BD",X"15",
		X"B6",X"15",X"B1",X"15",X"AA",X"15",X"A1",X"15",X"9A",X"15",X"92",X"15",X"8A",X"15",X"82",X"15",
		X"79",X"15",X"6E",X"15",X"65",X"15",X"5A",X"15",X"51",X"15",X"44",X"15",X"39",X"15",X"2E",X"15",
		X"22",X"15",X"15",X"15",X"0A",X"15",X"FD",X"14",X"F1",X"14",X"E4",X"14",X"D7",X"14",X"C9",X"14",
		X"BC",X"14",X"AC",X"14",X"9F",X"14",X"91",X"14",X"82",X"14",X"73",X"14",X"65",X"14",X"55",X"14",
		X"47",X"14",X"38",X"14",X"29",X"14",X"1A",X"14",X"09",X"14",X"FA",X"13",X"E9",X"13",X"D9",X"13",
		X"C8",X"13",X"B9",X"13",X"A8",X"13",X"98",X"13",X"87",X"13",X"78",X"13",X"65",X"13",X"56",X"13",
		X"45",X"13",X"35",X"13",X"23",X"13",X"13",X"13",X"02",X"13",X"F2",X"12",X"DF",X"12",X"CE",X"12",
		X"BE",X"12",X"AC",X"12",X"9A",X"12",X"8B",X"12",X"78",X"12",X"69",X"12",X"56",X"12",X"44",X"12",
		X"33",X"12",X"23",X"12",X"11",X"12",X"FF",X"11",X"EE",X"11",X"DD",X"11",X"CB",X"11",X"B9",X"11",
		X"A8",X"11",X"96",X"11",X"85",X"11",X"74",X"11",X"62",X"11",X"50",X"11",X"40",X"11",X"2F",X"11",
		X"1D",X"11",X"0C",X"11",X"FA",X"10",X"E9",X"10",X"D9",X"10",X"C7",X"10",X"B5",X"10",X"A4",X"10",
		X"92",X"10",X"81",X"10",X"70",X"10",X"5F",X"10",X"4D",X"10",X"3D",X"10",X"2C",X"10",X"1B",X"10",
		X"0A",X"10",X"F8",X"0F",X"E8",X"0F",X"D8",X"0F",X"C7",X"0F",X"B6",X"0F",X"A5",X"0F",X"93",X"0F",
		X"82",X"0F",X"72",X"0F",X"62",X"0F",X"52",X"0F",X"40",X"0F",X"30",X"0F",X"1E",X"0F",X"0E",X"0F",
		X"FE",X"0E",X"EE",X"0E",X"DD",X"0E",X"CD",X"0E",X"BD",X"0E",X"AB",X"0E",X"9D",X"0E",X"8C",X"0E",
		X"7C",X"0E",X"6C",X"0E",X"5C",X"0E",X"4C",X"0E",X"3D",X"0E",X"2C",X"0E",X"1C",X"0E",X"0C",X"0E",
		X"FC",X"0D",X"ED",X"0D",X"DC",X"0D",X"CE",X"0D",X"BD",X"0D",X"B0",X"0D",X"9E",X"0D",X"8F",X"0D",
		X"80",X"0D",X"71",X"0D",X"61",X"0D",X"52",X"0D",X"42",X"0D",X"32",X"0D",X"23",X"0D",X"16",X"0D",
		X"06",X"0D",X"F6",X"0C",X"E6",X"0C",X"D9",X"0C",X"CA",X"0C",X"BC",X"0C",X"AC",X"0C",X"9D",X"0C",
		X"8D",X"0C",X"80",X"0C",X"71",X"0C",X"62",X"0C",X"52",X"0C",X"45",X"0C",X"36",X"0C",X"28",X"0C",
		X"1A",X"0C",X"0C",X"0C",X"FD",X"0B",X"F0",X"0B",X"E1",X"0B",X"D3",X"0B",X"C6",X"0B",X"B7",X"0B",
		X"A8",X"0B",X"9C",X"0B",X"8B",X"0B",X"81",X"0B",X"4E",X"0B",X"CC",X"0A",X"17",X"0A",X"44",X"09",
		X"5C",X"08",X"69",X"07",X"72",X"06",X"7B",X"05",X"85",X"04",X"93",X"03",X"A6",X"02",X"C0",X"01",
		X"DF",X"00",X"06",X"00",X"36",X"FF",X"69",X"FE",X"A3",X"FD",X"E3",X"FC",X"2B",X"FC",X"79",X"FB",
		X"CC",X"FA",X"26",X"FA",X"85",X"F9",X"E9",X"F8",X"56",X"F8",X"C5",X"F7",X"3A",X"F7",X"B5",X"F6",
		X"34",X"F6",X"B7",X"F5",X"3F",X"F5",X"CD",X"F4",X"5D",X"F4",X"F1",X"F3",X"89",X"F3",X"27",X"F3",
		X"C9",X"F2",X"6E",X"F2",X"14",X"F2",X"C1",X"F1",X"6E",X"F1",X"20",X"F1",X"D5",X"F0",X"8D",X"F0",
		X"49",X"F0",X"05",X"F0",X"C7",X"EF",X"8B",X"EF",X"50",X"EF",X"18",X"EF",X"E3",X"EE",X"B1",X"EE",
		X"80",X"EE",X"54",X"EE",X"25",X"EE",X"15",X"EE",X"53",X"EE",X"C8",X"EE",X"61",X"EF",X"0E",X"F0",
		X"C8",X"F0",X"8C",X"F1",X"4F",X"F2",X"14",X"F3",X"D5",X"F3",X"95",X"F4",X"4F",X"F5",X"06",X"F6",
		X"B5",X"F6",X"63",X"F7",X"0B",X"F8",X"AB",X"F8",X"48",X"F9",X"E0",X"F9",X"73",X"FA",X"00",X"FB",
		X"8A",X"FB",X"0F",X"FC",X"90",X"FC",X"0D",X"FD",X"85",X"FD",X"F8",X"FD",X"68",X"FE",X"9A",X"FE",
		X"83",X"FE",X"41",X"FE",X"DF",X"FD",X"6E",X"FD",X"EF",X"FC",X"6A",X"FC",X"E2",X"FB",X"5B",X"FB",
		X"D4",X"FA",X"50",X"FA",X"CF",X"F9",X"51",X"F9",X"D6",X"F8",X"60",X"F8",X"EE",X"F7",X"80",X"F7",
		X"14",X"F7",X"AF",X"F6",X"4C",X"F6",X"ED",X"F5",X"90",X"F5",X"37",X"F5",X"E2",X"F4",X"90",X"F4",
		X"43",X"F4",X"F6",X"F3",X"AE",X"F3",X"69",X"F3",X"24",X"F3",X"E4",X"F2",X"A8",X"F2",X"6D",X"F2",
		X"34",X"F2",X"FE",X"F1",X"CA",X"F1",X"98",X"F1",X"69",X"F1",X"3B",X"F1",X"11",X"F1",X"E7",X"F0",
		X"C0",X"F0",X"9A",X"F0",X"77",X"F0",X"53",X"F0",X"35",X"F0",X"15",X"F0",X"F9",X"EF",X"DD",X"EF",
		X"C3",X"EF",X"AB",X"EF",X"94",X"EF",X"7D",X"EF",X"68",X"EF",X"55",X"EF",X"72",X"EF",X"D6",X"EF",
		X"62",X"F0",X"0D",X"F1",X"C7",X"F1",X"8A",X"F2",X"53",X"F3",X"1D",X"F4",X"E5",X"F4",X"AB",X"F5",
		X"6B",X"F6",X"28",X"F7",X"DF",X"F7",X"92",X"F8",X"3E",X"F9",X"E7",X"F9",X"8B",X"FA",X"27",X"FB",
		X"C1",X"FB",X"55",X"FC",X"E1",X"FC",X"6C",X"FD",X"F2",X"FD",X"71",X"FE",X"EC",X"FE",X"66",X"FF",
		X"DB",X"FF",X"4C",X"00",X"BB",X"00",X"25",X"01",X"8A",X"01",X"EE",X"01",X"4D",X"02",X"A9",X"02",
		X"01",X"03",X"57",X"03",X"AC",X"03",X"FA",X"03",X"46",X"04",X"91",X"04",X"D9",X"04",X"1D",X"05",
		X"60",X"05",X"9F",X"05",X"DD",X"05",X"19",X"06",X"52",X"06",X"88",X"06",X"BE",X"06",X"F0",X"06",
		X"21",X"07",X"4F",X"07",X"7D",X"07",X"A9",X"07",X"D2",X"07",X"F9",X"07",X"20",X"08",X"44",X"08",
		X"67",X"08",X"8A",X"08",X"AA",X"08",X"C8",X"08",X"E6",X"08",X"01",X"09",X"1D",X"09",X"36",X"09",
		X"4E",X"09",X"66",X"09",X"7C",X"09",X"92",X"09",X"A5",X"09",X"B9",X"09",X"CA",X"09",X"DB",X"09",
		X"EC",X"09",X"FB",X"09",X"0A",X"0A",X"16",X"0A",X"23",X"0A",X"2F",X"0A",X"3B",X"0A",X"46",X"0A",
		X"49",X"0A",X"10",X"0A",X"9C",X"09",X"06",X"09",X"58",X"08",X"9F",X"07",X"DD",X"06",X"1A",X"06",
		X"58",X"05",X"95",X"04",X"D8",X"03",X"1F",X"03",X"6B",X"02",X"BB",X"01",X"11",X"01",X"6B",X"00",
		X"CD",X"FF",X"32",X"FF",X"9C",X"FE",X"0C",X"FE",X"81",X"FD",X"FA",X"FC",X"78",X"FC",X"FA",X"FB",
		X"82",X"FB",X"0C",X"FB",X"9C",X"FA",X"30",X"FA",X"C7",X"F9",X"62",X"F9",X"02",X"F9",X"A5",X"F8",
		X"4A",X"F8",X"F2",X"F7",X"9F",X"F7",X"4E",X"F7",X"01",X"F7",X"B7",X"F6",X"6E",X"F6",X"2A",X"F6",
		X"E7",X"F5",X"A9",X"F5",X"6C",X"F5",X"31",X"F5",X"FA",X"F4",X"C3",X"F4",X"8F",X"F4",X"5F",X"F4",
		X"2E",X"F4",X"02",X"F4",X"D6",X"F3",X"AD",X"F3",X"84",X"F3",X"61",X"F3",X"3A",X"F3",X"2C",X"F3",
		X"61",X"F3",X"C6",X"F3",X"48",X"F4",X"DB",X"F4",X"7D",X"F5",X"22",X"F6",X"CB",X"F6",X"75",X"F7",
		X"1C",X"F8",X"BE",X"F8",X"5F",X"F9",X"FA",X"F9",X"92",X"FA",X"25",X"FB",X"B3",X"FB",X"3D",X"FC",
		X"C6",X"FC",X"47",X"FD",X"C4",X"FD",X"3C",X"FE",X"B2",X"FE",X"25",X"FF",X"92",X"FF",X"FB",X"FF",
		X"61",X"00",X"C4",X"00",X"24",X"01",X"7F",X"01",X"DA",X"01",X"30",X"02",X"82",X"02",X"D1",X"02",
		X"20",X"03",X"6A",X"03",X"B2",X"03",X"F8",X"03",X"39",X"04",X"79",X"04",X"B8",X"04",X"F3",X"04",
		X"2C",X"05",X"64",X"05",X"9A",X"05",X"CE",X"05",X"FE",X"05",X"2E",X"06",X"5C",X"06",X"89",X"06",
		X"B2",X"06",X"DA",X"06",X"00",X"07",X"27",X"07",X"4A",X"07",X"6D",X"07",X"8D",X"07",X"AD",X"07",
		X"CC",X"07",X"E8",X"07",X"03",X"08",X"1E",X"08",X"37",X"08",X"50",X"08",X"67",X"08",X"7C",X"08",
		X"92",X"08",X"A6",X"08",X"B7",X"08",X"CC",X"08",X"DB",X"08",X"EC",X"08",X"FB",X"08",X"09",X"09",
		X"16",X"09",X"25",X"09",X"30",X"09",X"3D",X"09",X"46",X"09",X"50",X"09",X"59",X"09",X"62",X"09",
		X"6A",X"09",X"73",X"09",X"55",X"09",X"FA",X"08",X"7D",X"08",X"E5",X"07",X"44",X"07",X"96",X"06",
		X"E8",X"05",X"37",X"05",X"89",X"04",X"DE",X"03",X"34",X"03",X"92",X"02",X"F1",X"01",X"57",X"01",
		X"C1",X"00",X"30",X"00",X"A4",X"FF",X"1D",X"FF",X"99",X"FE",X"1B",X"FE",X"A0",X"FD",X"2A",X"FD",
		X"B8",X"FC",X"4A",X"FC",X"DF",X"FB",X"78",X"FB",X"16",X"FB",X"B6",X"FA",X"5C",X"FA",X"02",X"FA",
		X"AF",X"F9",X"5C",X"F9",X"0D",X"F9",X"C1",X"F8",X"78",X"F8",X"32",X"F8",X"EF",X"F7",X"AE",X"F7",
		X"6E",X"F7",X"34",X"F7",X"F7",X"F6",X"C2",X"F6",X"8C",X"F6",X"59",X"F6",X"29",X"F6",X"FA",X"F5",
		X"CC",X"F5",X"A1",X"F5",X"77",X"F5",X"51",X"F5",X"2B",X"F5",X"07",X"F5",X"E4",X"F4",X"C6",X"F4",
		X"A4",X"F4",X"A1",X"F4",X"DC",X"F4",X"3B",X"F5",X"B3",X"F5",X"3A",X"F6",X"C8",X"F6",X"5F",X"F7",
		X"F6",X"F7",X"8B",X"F8",X"1F",X"F9",X"B1",X"F9",X"40",X"FA",X"CA",X"FA",X"51",X"FB",X"D3",X"FB",
		X"51",X"FC",X"CC",X"FC",X"43",X"FD",X"B6",X"FD",X"25",X"FE",X"91",X"FE",X"F9",X"FE",X"5E",X"FF",
		X"BE",X"FF",X"1D",X"00",X"77",X"00",X"CF",X"00",X"21",X"01",X"74",X"01",X"C1",X"01",X"10",X"02",
		X"59",X"02",X"9E",X"02",X"E3",X"02",X"25",X"03",X"65",X"03",X"A4",X"03",X"DE",X"03",X"16",X"04",
		X"4B",X"04",X"82",X"04",X"B5",X"04",X"E7",X"04",X"14",X"05",X"42",X"05",X"6F",X"05",X"97",X"05",
		X"C0",X"05",X"E5",X"05",X"0C",X"06",X"2F",X"06",X"51",X"06",X"74",X"06",X"93",X"06",X"B2",X"06",
		X"BB",X"06",X"8A",X"06",X"36",X"06",X"C6",X"05",X"49",X"05",X"C0",X"04",X"35",X"04",X"A7",X"03",
		X"1A",X"03",X"90",X"02",X"06",X"02",X"81",X"01",X"FF",X"00",X"80",X"00",X"06",X"00",X"91",X"FF",
		X"1D",X"FF",X"AF",X"FE",X"44",X"FE",X"DD",X"FD",X"79",X"FD",X"18",X"FD",X"BD",X"FC",X"62",X"FC",
		X"0B",X"FC",X"B7",X"FB",X"67",X"FB",X"1C",X"FB",X"FD",X"FA",X"11",X"FB",X"45",X"FB",X"90",X"FB",
		X"E5",X"FB",X"43",X"FC",X"A7",X"FC",X"0D",X"FD",X"70",X"FD",X"D8",X"FD",X"38",X"FE",X"9A",X"FE",
		X"F8",X"FE",X"55",X"FF",X"AD",X"FF",X"04",X"00",X"58",X"00",X"A7",X"00",X"F5",X"00",X"41",X"01",
		X"8B",X"01",X"D0",X"01",X"14",X"02",X"56",X"02",X"96",X"02",X"D2",X"02",X"0E",X"03",X"3A",X"03",
		X"2F",X"03",X"FB",X"02",X"B0",X"02",X"53",X"02",X"EC",X"01",X"80",X"01",X"11",X"01",X"A2",X"00",
		X"35",X"00",X"CA",X"FF",X"5F",X"FF",X"F7",X"FE",X"93",X"FE",X"30",X"FE",X"D3",X"FD",X"76",X"FD",
		X"1E",X"FD",X"C7",X"FC",X"76",X"FC",X"26",X"FC",X"DB",X"FB",X"91",X"FB",X"49",X"FB",X"06",X"FB",
		X"C3",X"FA",X"83",X"FA",X"46",X"FA",X"0A",X"FA",X"D2",X"F9",X"9B",X"F9",X"68",X"F9",X"35",X"F9",
		X"05",X"F9",X"D8",X"F8",X"AC",X"F8",X"81",X"F8",X"57",X"F8",X"30",X"F8",X"0B",X"F8",X"E6",X"F7",
		X"C5",X"F7",X"A5",X"F7",X"85",X"F7",X"68",X"F7",X"4B",X"F7",X"30",X"F7",X"16",X"F7",X"FC",X"F6",
		X"E5",X"F6",X"CE",X"F6",X"B9",X"F6",X"A5",X"F6",X"91",X"F6",X"80",X"F6",X"6F",X"F6",X"5F",X"F6",
		X"4F",X"F6",X"42",X"F6",X"35",X"F6",X"27",X"F6",X"1D",X"F6",X"12",X"F6",X"07",X"F6",X"FF",X"F5",
		X"F5",X"F5",X"EE",X"F5",X"E6",X"F5",X"DF",X"F5",X"D9",X"F5",X"D4",X"F5",X"CF",X"F5",X"CB",X"F5",
		X"C8",X"F5",X"C4",X"F5",X"C0",X"F5",X"C0",X"F5",X"BD",X"F5",X"C0",X"F5",X"B7",X"F5",X"A1",X"F5",
		X"A4",X"F5",X"A2",X"F5",X"A4",X"F5",X"A4",X"F5",X"A7",X"F5",X"A8",X"F5",X"AD",X"F5",X"AF",X"F5",
		X"B2",X"F5",X"B4",X"F5",X"B9",X"F5",X"BD",X"F5",X"C1",X"F5",X"C7",X"F5",X"CB",X"F5",X"D1",X"F5",
		X"D6",X"F5",X"DC",X"F5",X"E1",X"F5",X"E8",X"F5",X"EE",X"F5",X"F5",X"F5",X"FC",X"F5",X"03",X"F6",
		X"09",X"F6",X"11",X"F6",X"17",X"F6",X"1E",X"F6",X"27",X"F6",X"34",X"F6",X"6B",X"F6",X"CB",X"F6",
		X"40",X"F7",X"C7",X"F7",X"57",X"F8",X"E8",X"F8",X"7C",X"F9",X"11",X"FA",X"A2",X"FA",X"31",X"FB",
		X"BD",X"FB",X"46",X"FC",X"CB",X"FC",X"4A",X"FD",X"C8",X"FD",X"42",X"FE",X"B6",X"FE",X"28",X"FF",
		X"95",X"FF",X"FE",X"FF",X"64",X"00",X"C7",X"00",X"26",X"01",X"83",X"01",X"DC",X"01",X"32",X"02",
		X"84",X"02",X"C3",X"02",X"CE",X"02",X"B8",X"02",X"8D",X"02",X"57",X"02",X"15",X"02",X"CD",X"01",
		X"85",X"01",X"3C",X"01",X"F1",X"00",X"A8",X"00",X"60",X"00",X"19",X"00",X"D7",X"FF",X"95",X"FF",
		X"53",X"FF",X"16",X"FF",X"DA",X"FE",X"A0",X"FE",X"69",X"FE",X"34",X"FE",X"00",X"FE",X"CE",X"FD",
		X"9E",X"FD",X"6E",X"FD",X"42",X"FD",X"18",X"FD",X"F1",X"FC",X"F0",X"FC",X"17",X"FD",X"57",X"FD",
		X"AA",X"FD",X"05",X"FE",X"69",X"FE",X"CC",X"FE",X"32",X"FF",X"97",X"FF",X"FA",X"FF",X"5B",X"00",
		X"BA",X"00",X"17",X"01",X"72",X"01",X"C8",X"01",X"1E",X"02",X"6E",X"02",X"BD",X"02",X"09",X"03",
		X"52",X"03",X"99",X"03",X"DE",X"03",X"22",X"04",X"60",X"04",X"9D",X"04",X"D8",X"04",X"10",X"05",
		X"48",X"05",X"7C",X"05",X"B2",X"05",X"E1",X"05",X"11",X"06",X"3F",X"06",X"69",X"06",X"94",X"06",
		X"BD",X"06",X"E3",X"06",X"08",X"07",X"2C",X"07",X"4E",X"07",X"6E",X"07",X"90",X"07",X"AE",X"07",
		X"CB",X"07",X"E7",X"07",X"02",X"08",X"19",X"08",X"32",X"08",X"4A",X"08",X"60",X"08",X"76",X"08",
		X"89",X"08",X"9C",X"08",X"AF",X"08",X"B7",X"08",X"94",X"08",X"52",X"08",X"FB",X"07",X"9A",X"07",
		X"2E",X"07",X"C0",X"06",X"51",X"06",X"E0",X"05",X"73",X"05",X"07",X"05",X"9C",X"04",X"36",X"04",
		X"D1",X"03",X"71",X"03",X"11",X"03",X"B7",X"02",X"5F",X"02",X"09",X"02",X"B5",X"01",X"67",X"01",
		X"18",X"01",X"CF",X"00",X"87",X"00",X"43",X"00",X"00",X"00",X"C1",X"FF",X"82",X"FF",X"60",X"FF",
		X"68",X"FF",X"87",X"FF",X"B9",X"FF",X"F5",X"FF",X"38",X"00",X"7F",X"00",X"C8",X"00",X"12",X"01",
		X"5B",X"01",X"A3",X"01",X"EA",X"01",X"2E",X"02",X"71",X"02",X"B2",X"02",X"F0",X"02",X"2D",X"03",
		X"67",X"03",X"A0",X"03",X"D6",X"03",X"0B",X"04",X"3E",X"04",X"6E",X"04",X"9D",X"04",X"CA",X"04",
		X"F6",X"04",X"20",X"05",X"43",X"05",X"3F",X"05",X"1A",X"05",X"E1",X"04",X"9A",X"04",X"4E",X"04",
		X"FA",X"03",X"A6",X"03",X"4F",X"03",X"FA",X"02",X"A5",X"02",X"54",X"02",X"04",X"02",X"B6",X"01",
		X"6A",X"01",X"21",X"01",X"D9",X"00",X"95",X"00",X"52",X"00",X"13",X"00",X"D5",X"FF",X"99",X"FF",
		X"60",X"FF",X"29",X"FF",X"F2",X"FE",X"C0",X"FE",X"8F",X"FE",X"5F",X"FE",X"31",X"FE",X"05",X"FE",
		X"D9",X"FD",X"B0",X"FD",X"88",X"FD",X"64",X"FD",X"3E",X"FD",X"1C",X"FD",X"FA",X"FC",X"DA",X"FC",
		X"BA",X"FC",X"9E",X"FC",X"80",X"FC",X"64",X"FC",X"4B",X"FC",X"32",X"FC",X"19",X"FC",X"02",X"FC",
		X"ED",X"FB",X"D8",X"FB",X"C4",X"FB",X"B2",X"FB",X"9E",X"FB",X"8D",X"FB",X"7C",X"FB",X"6C",X"FB",
		X"5E",X"FB",X"50",X"FB",X"42",X"FB",X"36",X"FB",X"29",X"FB",X"1E",X"FB",X"13",X"FB",X"08",X"FB",
		X"00",X"FB",X"F6",X"FA",X"EE",X"FA",X"E6",X"FA",X"DF",X"FA",X"D8",X"FA",X"D1",X"FA",X"CC",X"FA",
		X"C7",X"FA",X"C3",X"FA",X"BE",X"FA",X"B9",X"FA",X"B7",X"FA",X"B3",X"FA",X"B1",X"FA",X"B0",X"FA",
		X"AE",X"FA",X"AB",X"FA",X"A9",X"FA",X"AA",X"FA",X"A9",X"FA",X"A8",X"FA",X"A8",X"FA",X"A8",X"FA",
		X"A8",X"FA",X"AA",X"FA",X"AA",X"FA",X"AC",X"FA",X"AD",X"FA",X"AE",X"FA",X"B1",X"FA",X"B3",X"FA",
		X"B4",X"FA",X"B7",X"FA",X"BB",X"FA",X"BE",X"FA",X"C1",X"FA",X"C4",X"FA",X"C7",X"FA",X"CC",X"FA",
		X"D0",X"FA",X"D3",X"FA",X"D8",X"FA",X"DB",X"FA",X"E0",X"FA",X"E4",X"FA",X"E9",X"FA",X"EE",X"FA",
		X"F5",X"FA",X"16",X"FB",X"56",X"FB",X"A8",X"FB",X"05",X"FC",X"69",X"FC",X"D4",X"FC",X"3C",X"FD",
		X"A5",X"FD",X"0D",X"FE",X"74",X"FE",X"D9",X"FE",X"3A",X"FF",X"98",X"FF",X"F4",X"FF",X"4B",X"00",
		X"A3",X"00",X"F5",X"00",X"47",X"01",X"95",X"01",X"E0",X"01",X"29",X"02",X"6E",X"02",X"B3",X"02",
		X"F4",X"02",X"32",X"03",X"6F",X"03",X"AA",X"03",X"E3",X"03",X"1A",X"04",X"4D",X"04",X"81",X"04",
		X"B2",X"04",X"E0",X"04",X"0F",X"05",X"39",X"05",X"63",X"05",X"8C",X"05",X"B2",X"05",X"D7",X"05",
		X"FB",X"05",X"1F",X"06",X"3F",X"06",X"60",X"06",X"7E",X"06",X"9C",X"06",X"B7",X"06",X"D1",X"06",
		X"EC",X"06",X"05",X"07",X"1C",X"07",X"33",X"07",X"48",X"07",X"5D",X"07",X"71",X"07",X"84",X"07",
		X"80",X"07",X"5D",X"07",X"29",X"07",X"E6",X"06",X"9E",X"06",X"50",X"06",X"02",X"06",X"B2",X"05",
		X"63",X"05",X"16",X"05",X"C7",X"04",X"7E",X"04",X"34",X"04",X"EE",X"03",X"A9",X"03",X"67",X"03",
		X"26",X"03",X"E8",X"02",X"AC",X"02",X"73",X"02",X"3B",X"02",X"04",X"02",X"D0",X"01",X"9D",X"01",
		X"6D",X"01",X"3E",X"01",X"0F",X"01",X"EA",X"00",X"E2",X"00",X"F3",X"00",X"14",X"01",X"3F",X"01",
		X"71",X"01",X"A6",X"01",X"DE",X"01",X"15",X"02",X"4C",X"02",X"83",X"02",X"B8",X"02",X"EB",X"02",
		X"20",X"03",X"50",X"03",X"80",X"03",X"AE",X"03",X"DB",X"03",X"06",X"04",X"30",X"04",X"58",X"04",
		X"7E",X"04",X"A3",X"04",X"C6",X"04",X"E9",X"04",X"0B",X"05",X"2A",X"05",X"48",X"05",X"66",X"05",
		X"81",X"05",X"9D",X"05",X"B7",X"05",X"D0",X"05",X"E7",X"05",X"FF",X"05",X"14",X"06",X"2A",X"06",
		X"3D",X"06",X"51",X"06",X"62",X"06",X"75",X"06",X"84",X"06",X"93",X"06",X"A3",X"06",X"B1",X"06",
		X"BF",X"06",X"CC",X"06",X"D7",X"06",X"E4",X"06",X"EF",X"06",X"F9",X"06",X"04",X"07",X"11",X"07",
		X"2A",X"07",X"2F",X"07",X"35",X"07",X"1F",X"07",X"F3",X"06",X"B8",X"06",X"75",X"06",X"2C",X"06",
		X"DD",X"05",X"91",X"05",X"44",X"05",X"F8",X"04",X"AC",X"04",X"64",X"04",X"1B",X"04",X"D5",X"03",
		X"92",X"03",X"51",X"03",X"10",X"03",X"D4",X"02",X"99",X"02",X"5E",X"02",X"29",X"02",X"F3",X"01",
		X"BF",X"01",X"8D",X"01",X"5D",X"01",X"2E",X"01",X"02",X"01",X"D7",X"00",X"AE",X"00",X"86",X"00",
		X"5E",X"00",X"39",X"00",X"15",X"00",X"F4",X"FF",X"D3",X"FF",X"B2",X"FF",X"94",X"FF",X"76",X"FF",
		X"5A",X"FF",X"3F",X"FF",X"25",X"FF",X"0B",X"FF",X"F4",X"FE",X"DB",X"FE",X"C5",X"FE",X"AF",X"FE",
		X"9B",X"FE",X"86",X"FE",X"73",X"FE",X"63",X"FE",X"50",X"FE",X"40",X"FE",X"32",X"FE",X"21",X"FE",
		X"13",X"FE",X"05",X"FE",X"F8",X"FD",X"EC",X"FD",X"E0",X"FD",X"D5",X"FD",X"C8",X"FD",X"BF",X"FD",
		X"B6",X"FD",X"AA",X"FD",X"A4",X"FD",X"9B",X"FD",X"95",X"FD",X"8D",X"FD",X"87",X"FD",X"80",X"FD",
		X"7A",X"FD",X"75",X"FD",X"71",X"FD",X"6C",X"FD",X"67",X"FD",X"63",X"FD",X"5F",X"FD",X"5C",X"FD",
		X"59",X"FD",X"56",X"FD",X"54",X"FD",X"51",X"FD",X"4F",X"FD",X"4E",X"FD",X"4C",X"FD",X"4B",X"FD",
		X"4A",X"FD",X"4A",X"FD",X"48",X"FD",X"49",X"FD",X"48",X"FD",X"49",X"FD",X"48",X"FD",X"49",X"FD",
		X"4A",X"FD",X"4B",X"FD",X"4D",X"FD",X"4E",X"FD",X"50",X"FD",X"53",X"FD",X"53",X"FD",X"55",X"FD",
		X"57",X"FD",X"59",X"FD",X"5B",X"FD",X"5F",X"FD",X"60",X"FD",X"63",X"FD",X"68",X"FD",X"6A",X"FD",
		X"72",X"FD",X"92",X"FD",X"C2",X"FD",X"FD",X"FD",X"3F",X"FE",X"82",X"FE",X"C9",X"FE",X"10",X"FF",
		X"55",X"FF",X"9B",X"FF",X"DF",X"FF",X"20",X"00",X"5F",X"00",X"9E",X"00",X"DA",X"00",X"15",X"01",
		X"4E",X"01",X"85",X"01",X"BA",X"01",X"EC",X"01",X"1F",X"02",X"4F",X"02",X"7C",X"02",X"A9",X"02",
		X"D3",X"02",X"FD",X"02",X"25",X"03",X"4A",X"03",X"62",X"03",X"62",X"03",X"55",X"03",X"3F",X"03",
		X"22",X"03",X"02",X"03",X"E0",X"02",X"BC",X"02",X"9A",X"02",X"77",X"02",X"55",X"02",X"33",X"02",
		X"11",X"02",X"F0",X"01",X"D1",X"01",X"B3",X"01",X"97",X"01",X"7A",X"01",X"5E",X"01",X"45",X"01",
		X"2B",X"01",X"13",X"01",X"FC",X"00",X"E5",X"00",X"D0",X"00",X"BA",X"00",X"A6",X"00",X"96",X"00",
		X"9A",X"00",X"AF",X"00",X"CF",X"00",X"F5",X"00",X"1E",X"01",X"4A",X"01",X"77",X"01",X"A5",X"01",
		X"D3",X"01",X"FD",X"01",X"29",X"02",X"53",X"02",X"7D",X"02",X"A4",X"02",X"CB",X"02",X"F0",X"02",
		X"14",X"03",X"37",X"03",X"57",X"03",X"78",X"03",X"97",X"03",X"B5",X"03",X"D2",X"03",X"ED",X"03",
		X"09",X"04",X"21",X"04",X"3A",X"04",X"47",X"04",X"41",X"04",X"2D",X"04",X"12",X"04",X"F2",X"03",
		X"CE",X"03",X"A8",X"03",X"82",X"03",X"5B",X"03",X"36",X"03",X"0F",X"03",X"EC",X"02",X"C7",X"02",
		X"A4",X"02",X"83",X"02",X"61",X"02",X"42",X"02",X"23",X"02",X"06",X"02",X"E9",X"01",X"CE",X"01",
		X"B5",X"01",X"9B",X"01",X"81",X"01",X"6A",X"01",X"53",X"01",X"3C",X"01",X"28",X"01",X"27",X"01",
		X"34",X"01",X"4B",X"01",X"68",X"01",X"88",X"01",X"AC",X"01",X"D1",X"01",X"F6",X"01",X"1B",X"02",
		X"3D",X"02",X"63",X"02",X"83",X"02",X"A6",X"02",X"C6",X"02",X"E5",X"02",X"03",X"03",X"21",X"03",
		X"3D",X"03",X"57",X"03",X"71",X"03",X"8A",X"03",X"A4",X"03",X"BA",X"03",X"D1",X"03",X"E6",X"03",
		X"FA",X"03",X"0E",X"04",X"1A",X"04",X"15",X"04",X"04",X"04",X"EA",X"03",X"CE",X"03",X"AD",X"03",
		X"8C",X"03",X"6A",X"03",X"48",X"03",X"23",X"03",X"00",X"03",X"DE",X"02",X"BF",X"02",X"9F",X"02",
		X"81",X"02",X"64",X"02",X"47",X"02",X"2A",X"02",X"10",X"02",X"F7",X"01",X"DD",X"01",X"C4",X"01",
		X"AE",X"01",X"98",X"01",X"82",X"01",X"6E",X"01",X"5B",X"01",X"48",X"01",X"43",X"01",X"4B",X"01",
		X"5F",X"01",X"76",X"01",X"91",X"01",X"B0",X"01",X"CE",X"01",X"EC",X"01",X"0C",X"02",X"2B",X"02",
		X"48",X"02",X"66",X"02",X"83",X"02",X"9E",X"02",X"B9",X"02",X"D4",X"02",X"EC",X"02",X"03",X"03",
		X"1B",X"03",X"30",X"03",X"47",X"03",X"5A",X"03",X"6E",X"03",X"81",X"03",X"93",X"03",X"A4",X"03",
		X"B7",X"03",X"C2",X"03",X"BF",X"03",X"AF",X"03",X"9C",X"03",X"83",X"03",X"67",X"03",X"49",X"03",
		X"29",X"03",X"0D",X"03",X"EF",X"02",X"D2",X"02",X"B6",X"02",X"99",X"02",X"7E",X"02",X"64",X"02",
		X"4B",X"02",X"32",X"02",X"1A",X"02",X"02",X"02",X"EC",X"01",X"D9",X"01",X"C4",X"01",X"B0",X"01",
		X"9A",X"01",X"89",X"01",X"78",X"01",X"67",X"01",X"56",X"01",X"47",X"01",X"38",X"01",X"28",X"01",
		X"1A",X"01",X"0D",X"01",X"00",X"01",X"F4",X"00",X"E9",X"00",X"DD",X"00",X"D4",X"00",X"C8",X"00",
		X"BE",X"00",X"B4",X"00",X"AB",X"00",X"A3",X"00",X"9B",X"00",X"92",X"00",X"8B",X"00",X"85",X"00",
		X"7E",X"00",X"77",X"00",X"71",X"00",X"6B",X"00",X"66",X"00",X"60",X"00",X"5B",X"00",X"56",X"00",
		X"55",X"00",X"5F",X"00",X"71",X"00",X"8C",X"00",X"A7",X"00",X"C5",X"00",X"E6",X"00",X"04",X"01",
		X"24",X"01",X"45",X"01",X"62",X"01",X"81",X"01",X"9E",X"01",X"BA",X"01",X"D5",X"01",X"F0",X"01",
		X"09",X"02",X"23",X"02",X"3B",X"02",X"51",X"02",X"66",X"02",X"7D",X"02",X"91",X"02",X"A5",X"02",
		X"B8",X"02",X"CB",X"02",X"DB",X"02",X"EC",X"02",X"FB",X"02",X"0B",X"03",X"1A",X"03",X"27",X"03",
		X"35",X"03",X"43",X"03",X"50",X"03",X"5B",X"03",X"67",X"03",X"72",X"03",X"7B",X"03",X"87",X"03",
		X"90",X"03",X"99",X"03",X"A0",X"03",X"A9",X"03",X"AF",X"03",X"B8",X"03",X"BE",X"03",X"C4",X"03",
		X"CC",X"03",X"D1",X"03",X"D6",X"03",X"DC",X"03",X"E1",X"03",X"E6",X"03",X"EA",X"03",X"ED",X"03",
		X"F3",X"03",X"F5",X"03",X"F8",X"03",X"FC",X"03",X"FE",X"03",X"00",X"04",X"02",X"04",X"05",X"04",
		X"06",X"04",X"08",X"04",X"0A",X"04",X"0B",X"04",X"0C",X"04",X"0C",X"04",X"0E",X"04",X"0E",X"04",
		X"0D",X"04",X"0D",X"04",X"0E",X"04",X"0E",X"04",X"0E",X"04",X"0E",X"04",X"0C",X"04",X"0B",X"04",
		X"0C",X"04",X"09",X"04",X"09",X"04",X"05",X"04",X"F7",X"03",X"E6",X"03",X"D8",X"03",X"BF",X"03",
		X"A5",X"03",X"8B",X"03",X"71",X"03",X"56",X"03",X"3E",X"03",X"24",X"03",X"0D",X"03",X"F5",X"02",
		X"DE",X"02",X"C9",X"02",X"B3",X"02",X"9E",X"02",X"89",X"02",X"76",X"02",X"64",X"02",X"51",X"02",
		X"42",X"02",X"30",X"02",X"1F",X"02",X"11",X"02",X"02",X"02",X"F3",X"01",X"E6",X"01",X"DF",X"01",
		X"E0",X"01",X"E4",X"01",X"EB",X"01",X"F5",X"01",X"FE",X"01",X"09",X"02",X"14",X"02",X"1F",X"02",
		X"2A",X"02",X"35",X"02",X"3F",X"02",X"47",X"02",X"53",X"02",X"5B",X"02",X"64",X"02",X"6C",X"02",
		X"73",X"02",X"7C",X"02",X"84",X"02",X"8B",X"02",X"91",X"02",X"98",X"02",X"9E",X"02",X"A3",X"02",
		X"A8",X"02",X"AF",X"02",X"B2",X"02",X"AD",X"02",X"A5",X"02",X"9A",X"02",X"8E",X"02",X"82",X"02",
		X"72",X"02",X"64",X"02",X"57",X"02",X"47",X"02",X"3A",X"02",X"2D",X"02",X"1F",X"02",X"13",X"02",
		X"07",X"02",X"FB",X"01",X"F1",X"01",X"E6",X"01",X"DA",X"01",X"D1",X"01",X"C7",X"01",X"BD",X"01",
		X"B5",X"01",X"AC",X"01",X"A4",X"01",X"9C",X"01",X"95",X"01",X"8D",X"01",X"87",X"01",X"80",X"01",
		X"7A",X"01",X"75",X"01",X"6F",X"01",X"6A",X"01",X"63",X"01",X"5F",X"01",X"59",X"01",X"54",X"01",
		X"52",X"01",X"4E",X"01",X"49",X"01",X"46",X"01",X"43",X"01",X"41",X"01",X"3E",X"01",X"3C",X"01",
		X"39",X"01",X"36",X"01",X"34",X"01",X"30",X"01",X"2F",X"01",X"2E",X"01",X"2C",X"01",X"2B",X"01",
		X"29",X"01",X"29",X"01",X"27",X"01",X"26",X"01",X"26",X"01",X"25",X"01",X"25",X"01",X"24",X"01",
		X"23",X"01",X"21",X"01",X"22",X"01",X"23",X"01",X"23",X"01",X"24",X"01",X"23",X"01",X"23",X"01",
		X"23",X"01",X"25",X"01",X"25",X"01",X"26",X"01",X"27",X"01",X"27",X"01",X"29",X"01",X"29",X"01",
		X"29",X"01",X"2A",X"01",X"2C",X"01",X"2D",X"01",X"2D",X"01",X"2F",X"01",X"31",X"01",X"32",X"01",
		X"33",X"01",X"35",X"01",X"35",X"01",X"37",X"01",X"38",X"01",X"3B",X"01",X"3C",X"01",X"3E",X"01",
		X"3F",X"01",X"41",X"01",X"43",X"01",X"43",X"01",X"47",X"01",X"49",X"01",X"49",X"01",X"4D",X"01",
		X"4D",X"01",X"4F",X"01",X"52",X"01",X"53",X"01",X"54",X"01",X"57",X"01",X"59",X"01",X"5A",X"01",
		X"5D",X"01",X"61",X"01",X"61",X"01",X"64",X"01",X"66",X"01",X"68",X"01",X"6A",X"01",X"6C",X"01",
		X"6E",X"01",X"70",X"01",X"73",X"01",X"75",X"01",X"76",X"01",X"78",X"01",X"7B",X"01",X"7D",X"01",
		X"7F",X"01",X"81",X"01",X"82",X"01",X"87",X"01",X"89",X"01",X"89",X"01",X"8C",X"01",X"90",X"01",
		X"91",X"01",X"93",X"01",X"95",X"01",X"98",X"01",X"9A",X"01",X"9D",X"01",X"A0",X"01",X"A1",X"01",
		X"A4",X"01",X"A6",X"01",X"A8",X"01",X"A9",X"01",X"AC",X"01",X"AF",X"01",X"B1",X"01",X"B2",X"01",
		X"B4",X"01",X"B7",X"01",X"B9",X"01",X"BD",X"01",X"BF",X"01",X"C1",X"01",X"C1",X"01",X"C5",X"01",
		X"C6",X"01",X"C9",X"01",X"CC",X"01",X"CE",X"01",X"D1",X"01",X"D2",X"01",X"D5",X"01",X"D7",X"01",
		X"D9",X"01",X"DB",X"01",X"DD",X"01",X"DF",X"01",X"E2",X"01",X"E4",X"01",X"E6",X"01",X"E8",X"01",
		X"EA",X"01",X"EC",X"01",X"EE",X"01",X"F1",X"01",X"F3",X"01",X"F5",X"01",X"F7",X"01",X"F9",X"01",
		X"FB",X"01",X"FC",X"01",X"00",X"02",X"02",X"02",X"03",X"02",X"06",X"02",X"09",X"02",X"0A",X"02",
		X"0B",X"02",X"0D",X"02",X"10",X"02",X"12",X"02",X"14",X"02",X"16",X"02",X"19",X"02",X"1B",X"02",
		X"1C",X"02",X"1D",X"02",X"21",X"02",X"21",X"02",X"24",X"02",X"26",X"02",X"29",X"02",X"2A",X"02",
		X"2B",X"02",X"2E",X"02",X"30",X"02",X"33",X"02",X"34",X"02",X"35",X"02",X"38",X"02",X"39",X"02",
		X"3B",X"02",X"3C",X"02",X"3F",X"02",X"41",X"02",X"42",X"02",X"45",X"02",X"47",X"02",X"47",X"02",
		X"4B",X"02",X"4D",X"02",X"4D",X"02",X"4E",X"02",X"52",X"02",X"53",X"02",X"56",X"02",X"57",X"02",
		X"59",X"02",X"5C",X"02",X"5D",X"02",X"5E",X"02",X"60",X"02",X"61",X"02",X"63",X"02",X"66",X"02",
		X"66",X"02",X"6A",X"02",X"6C",X"02",X"6D",X"02",X"6F",X"02",X"70",X"02",X"72",X"02",X"74",X"02",
		X"74",X"02",X"77",X"02",X"78",X"02",X"7B",X"02",X"7C",X"02",X"7E",X"02",X"7F",X"02",X"80",X"02",
		X"82",X"02",X"83",X"02",X"85",X"02",X"87",X"02",X"89",X"02",X"8A",X"02",X"8C",X"02",X"8D",X"02",
		X"8F",X"02",X"91",X"02",X"91",X"02",X"94",X"02",X"95",X"02",X"97",X"02",X"99",X"02",X"9A",X"02",
		X"9C",X"02",X"9E",X"02",X"9F",X"02",X"A1",X"02",X"A2",X"02",X"A3",X"02",X"A5",X"02",X"A7",X"02",
		X"A8",X"02",X"A9",X"02",X"AC",X"02",X"AD",X"02",X"AE",X"02",X"AF",X"02",X"B1",X"02",X"B3",X"02",
		X"B3",X"02",X"B5",X"02",X"B5",X"02",X"B8",X"02",X"B8",X"02",X"BC",X"02",X"BC",X"02",X"BD",X"02",
		X"BE",X"02",X"C0",X"02",X"C1",X"02",X"C3",X"02",X"C4",X"02",X"C4",X"02",X"C6",X"02",X"C9",X"02",
		X"C9",X"02",X"CC",X"02",X"CC",X"02",X"CF",X"02",X"CE",X"02",X"D1",X"02",X"D2",X"02",X"D3",X"02",
		X"D5",X"02",X"D7",X"02",X"D7",X"02",X"D8",X"02",X"DA",X"02",X"DA",X"02",X"DC",X"02",X"DD",X"02",
		X"DF",X"02",X"E0",X"02",X"E1",X"02",X"E1",X"02",X"E2",X"02",X"E5",X"02",X"E5",X"02",X"E7",X"02",
		X"E8",X"02",X"EA",X"02",X"EB",X"02",X"ED",X"02",X"EE",X"02",X"ED",X"02",X"F0",X"02",X"F0",X"02",
		X"F1",X"02",X"F2",X"02",X"F4",X"02",X"F5",X"02",X"F6",X"02",X"F6",X"02",X"F8",X"02",X"FA",X"02",
		X"FB",X"02",X"FC",X"02",X"FD",X"02",X"FE",X"02",X"FF",X"02",X"00",X"03",X"01",X"03",X"02",X"03",
		X"04",X"03",X"05",X"03",X"07",X"03",X"07",X"03",X"09",X"03",X"09",X"03",X"09",X"03",X"0A",X"03",
		X"0D",X"03",X"0E",X"03",X"0E",X"03",X"11",X"03",X"10",X"03",X"11",X"03",X"13",X"03",X"13",X"03",
		X"13",X"03",X"15",X"03",X"17",X"03",X"17",X"03",X"18",X"03",X"19",X"03",X"1A",X"03",X"1C",X"03",
		X"1C",X"03",X"1E",X"03",X"1E",X"03",X"21",X"03",X"21",X"03",X"22",X"03",X"22",X"03",X"23",X"03",
		X"24",X"03",X"27",X"03",X"2E",X"03",X"2F",X"03",X"2F",X"03",X"31",X"03",X"32",X"03",X"33",X"03",
		X"33",X"03",X"34",X"03",X"35",X"03",X"36",X"03",X"37",X"03",X"38",X"03",X"3A",X"03",X"3B",X"03",
		X"3A",X"03",X"3A",X"03",X"3C",X"03",X"3D",X"03",X"3F",X"03",X"3D",X"03",X"3E",X"03",X"40",X"03",
		X"41",X"03",X"42",X"03",X"42",X"03",X"44",X"03",X"44",X"03",X"46",X"03",X"44",X"03",X"47",X"03",
		X"47",X"03",X"49",X"03",X"4A",X"03",X"4A",X"03",X"4A",X"03",X"4B",X"03",X"4C",X"03",X"4D",X"03",
		X"4D",X"03",X"50",X"03",X"4F",X"03",X"51",X"03",X"51",X"03",X"52",X"03",X"51",X"03",X"53",X"03",
		X"53",X"03",X"54",X"03",X"56",X"03",X"55",X"03",X"57",X"03",X"57",X"03",X"58",X"03",X"59",X"03",
		X"58",X"03",X"5B",X"03",X"5A",X"03",X"5B",X"03",X"5D",X"03",X"5E",X"03",X"5F",X"03",X"5F",X"03",
		X"5F",X"03",X"60",X"03",X"61",X"03",X"61",X"03",X"62",X"03",X"61",X"03",X"64",X"03",X"64",X"03",
		X"64",X"03",X"65",X"03",X"66",X"03",X"66",X"03",X"68",X"03",X"67",X"03",X"69",X"03",X"6A",X"03",
		X"69",X"03",X"6A",X"03",X"6A",X"03",X"6B",X"03",X"6C",X"03",X"6C",X"03",X"6D",X"03",X"6E",X"03",
		X"6D",X"03",X"6E",X"03",X"70",X"03",X"70",X"03",X"71",X"03",X"72",X"03",X"71",X"03",X"71",X"03",
		X"71",X"03",X"74",X"03",X"74",X"03",X"75",X"03",X"75",X"03",X"75",X"03",X"75",X"03",X"77",X"03",
		X"77",X"03",X"77",X"03",X"78",X"03",X"78",X"03",X"79",X"03",X"7B",X"03",X"7A",X"03",X"7C",X"03",
		X"7B",X"03",X"7D",X"03",X"7D",X"03",X"7D",X"03",X"7E",X"03",X"7D",X"03",X"7F",X"03",X"7E",X"03",
		X"7F",X"03",X"80",X"03",X"80",X"03",X"81",X"03",X"80",X"03",X"81",X"03",X"81",X"03",X"82",X"03",
		X"82",X"03",X"82",X"03",X"85",X"03",X"83",X"03",X"85",X"03",X"85",X"03",X"86",X"03",X"86",X"03",
		X"87",X"03",X"88",X"03",X"88",X"03",X"89",X"03",X"88",X"03",X"89",X"03",X"8B",X"03",X"89",X"03",
		X"8B",X"03",X"8B",X"03",X"8B",X"03",X"8A",X"03",X"8C",X"03",X"8C",X"03",X"8C",X"03",X"8E",X"03",
		X"8E",X"03",X"8F",X"03",X"8D",X"03",X"90",X"03",X"8F",X"03",X"8E",X"03",X"8F",X"03",X"90",X"03",
		X"91",X"03",X"90",X"03",X"91",X"03",X"92",X"03",X"93",X"03",X"92",X"03",X"94",X"03",X"92",X"03",
		X"94",X"03",X"94",X"03",X"94",X"03",X"95",X"03",X"95",X"03",X"95",X"03",X"95",X"03",X"96",X"03",
		X"96",X"03",X"96",X"03",X"97",X"03",X"97",X"03",X"96",X"03",X"97",X"03",X"96",X"03",X"97",X"03",
		X"99",X"03",X"98",X"03",X"98",X"03",X"99",X"03",X"9A",X"03",X"99",X"03",X"9B",X"03",X"9B",X"03",
		X"9B",X"03",X"9D",X"03",X"9C",X"03",X"9D",X"03",X"9C",X"03",X"9E",X"03",X"9D",X"03",X"9C",X"03",
		X"9E",X"03",X"9D",X"03",X"9E",X"03",X"9E",X"03",X"9F",X"03",X"9F",X"03",X"9E",X"03",X"9E",X"03",
		X"9F",X"03",X"A0",X"03",X"A0",X"03",X"A0",X"03",X"A1",X"03",X"A1",X"03",X"A1",X"03",X"A2",X"03",
		X"A1",X"03",X"A3",X"03",X"A2",X"03",X"A3",X"03",X"A2",X"03",X"A3",X"03",X"A3",X"03",X"A3",X"03",
		X"A4",X"03",X"A3",X"03",X"A5",X"03",X"A3",X"03",X"A2",X"03",X"A5",X"03",X"A5",X"03",X"A5",X"03",
		X"A6",X"03",X"A6",X"03",X"A4",X"03",X"A5",X"03",X"A6",X"03",X"A5",X"03",X"A5",X"03",X"A7",X"03",
		X"A7",X"03",X"A8",X"03",X"A7",X"03",X"A7",X"03",X"A7",X"03",X"A7",X"03",X"A7",X"03",X"A8",X"03",
		X"A8",X"03",X"A7",X"03",X"A9",X"03",X"A8",X"03",X"A8",X"03",X"A9",X"03",X"A9",X"03",X"A8",X"03",
		X"A9",X"03",X"A9",X"03",X"AA",X"03",X"AA",X"03",X"AA",X"03",X"AA",X"03",X"AA",X"03",X"AA",X"03",
		X"AA",X"03",X"AA",X"03",X"AC",X"03",X"AB",X"03",X"AB",X"03",X"AB",X"03",X"AC",X"03",X"AB",X"03",
		X"AB",X"03",X"AA",X"03",X"AC",X"03",X"AA",X"03",X"AC",X"03",X"AC",X"03",X"AC",X"03",X"AC",X"03",
		X"AC",X"03",X"AC",X"03",X"AD",X"03",X"AD",X"03",X"AD",X"03",X"AD",X"03",X"AD",X"03",X"AC",X"03",
		X"AD",X"03",X"AD",X"03",X"AD",X"03",X"AC",X"03",X"AE",X"03",X"AD",X"03",X"AE",X"03",X"AE",X"03",
		X"AE",X"03",X"AF",X"03",X"AE",X"03",X"AD",X"03",X"AE",X"03",X"AE",X"03",X"AE",X"03",X"AE",X"03",
		X"AE",X"03",X"AF",X"03",X"AF",X"03",X"AF",X"03",X"AF",X"03",X"AF",X"03",X"AE",X"03",X"AE",X"03",
		X"AF",X"03",X"AF",X"03",X"AF",X"03",X"AF",X"03",X"B0",X"03",X"B0",X"03",X"AF",X"03",X"AE",X"03",
		X"AF",X"03",X"AF",X"03",X"AF",X"03",X"B0",X"03",X"AF",X"03",X"AF",X"03",X"AF",X"03",X"AE",X"03",
		X"B1",X"03",X"B0",X"03",X"B0",X"03",X"B0",X"03",X"AF",X"03",X"B0",X"03",X"B0",X"03",X"B1",X"03",
		X"B0",X"03",X"B1",X"03",X"B0",X"03",X"AF",X"03",X"AF",X"03",X"B1",X"03",X"B0",X"03",X"B0",X"03",
		X"B0",X"03",X"B1",X"03",X"B1",X"03",X"B0",X"03",X"B0",X"03",X"B1",X"03",X"B0",X"03",X"B0",X"03",
		X"B0",X"03",X"AF",X"03",X"B0",X"03",X"AF",X"03",X"AF",X"03",X"AF",X"03",X"B0",X"03",X"B0",X"03",
		X"B0",X"03",X"AF",X"03",X"AF",X"03",X"B1",X"03",X"B0",X"03",X"B0",X"03",X"B1",X"03",X"B0",X"03",
		X"B0",X"03",X"B0",X"03",X"B1",X"03",X"B0",X"03",X"B0",X"03",X"B0",X"03",X"B0",X"03",X"B0",X"03",
		X"B0",X"03",X"AF",X"03",X"B1",X"03",X"AF",X"03",X"B0",X"03",X"B0",X"03",X"AE",X"03",X"AF",X"03",
		X"AF",X"03",X"AF",X"03",X"AF",X"03",X"AF",X"03",X"AF",X"03",X"AE",X"03",X"AE",X"03",X"AE",X"03",
		X"AF",X"03",X"AF",X"03",X"B0",X"03",X"AF",X"03",X"AF",X"03",X"AF",X"03",X"AF",X"03",X"AF",X"03",
		X"AF",X"03",X"AF",X"03",X"AD",X"03",X"AE",X"03",X"AE",X"03",X"AE",X"03",X"AF",X"03",X"AD",X"03",
		X"AD",X"03",X"AE",X"03",X"AE",X"03",X"AD",X"03",X"AE",X"03",X"AE",X"03",X"AE",X"03",X"AE",X"03",
		X"AD",X"03",X"AD",X"03",X"AD",X"03",X"AD",X"03",X"AD",X"03",X"AD",X"03",X"AE",X"03",X"AD",X"03",
		X"AB",X"03",X"AC",X"03",X"AD",X"03",X"AC",X"03",X"AB",X"03",X"AC",X"03",X"AC",X"03",X"AC",X"03",
		X"AC",X"03",X"AB",X"03",X"AC",X"03",X"AC",X"03",X"AC",X"03",X"AD",X"03",X"AB",X"03",X"AB",X"03",
		X"AA",X"03",X"AC",X"03",X"AC",X"03",X"AC",X"03",X"AB",X"03",X"AB",X"03",X"AB",X"03",X"A9",X"03",
		X"A9",X"03",X"AB",X"03",X"A9",X"03",X"A9",X"03",X"AB",X"03",X"AA",X"03",X"AA",X"03",X"AB",X"03",
		X"AB",X"03",X"A9",X"03",X"AA",X"03",X"A9",X"03",X"A9",X"03",X"A9",X"03",X"A8",X"03",X"AA",X"03",
		X"A8",X"03",X"A7",X"03",X"A9",X"03",X"A7",X"03",X"A9",X"03",X"A8",X"03",X"AA",X"03",X"A7",X"03",
		X"A7",X"03",X"A8",X"03",X"A8",X"03",X"A8",X"03",X"A7",X"03",X"A6",X"03",X"A6",X"03",X"A6",X"03",
		X"A6",X"03",X"A6",X"03",X"A6",X"03",X"A6",X"03",X"A5",X"03",X"A8",X"03",X"A5",X"03",X"A5",X"03",
		X"A5",X"03",X"A5",X"03",X"A5",X"03",X"A6",X"03",X"A5",X"03",X"A5",X"03",X"A4",X"03",X"A4",X"03",
		X"A4",X"03",X"A4",X"03",X"A3",X"03",X"A4",X"03",X"A3",X"03",X"A3",X"03",X"A2",X"03",X"A3",X"03",
		X"A4",X"03",X"A2",X"03",X"A2",X"03",X"A2",X"03",X"A3",X"03",X"A3",X"03",X"A2",X"03",X"A2",X"03",
		X"A2",X"03",X"A0",X"03",X"A2",X"03",X"A1",X"03",X"A1",X"03",X"A2",X"03",X"A1",X"03",X"A0",X"03",
		X"A0",X"03",X"A0",X"03",X"A0",X"03",X"A0",X"03",X"9F",X"03",X"9F",X"03",X"9F",X"03",X"9F",X"03",
		X"A0",X"03",X"A0",X"03",X"9E",X"03",X"9E",X"03",X"9E",X"03",X"9F",X"03",X"9D",X"03",X"9D",X"03",
		X"9D",X"03",X"9D",X"03",X"9D",X"03",X"9D",X"03",X"9D",X"03",X"9B",X"03",X"9B",X"03",X"9C",X"03",
		X"9B",X"03",X"9B",X"03",X"9C",X"03",X"9B",X"03",X"9A",X"03",X"9A",X"03",X"9B",X"03",X"9B",X"03",
		X"9A",X"03",X"9A",X"03",X"9A",X"03",X"99",X"03",X"99",X"03",X"98",X"03",X"98",X"03",X"99",X"03",
		X"99",X"03",X"99",X"03",X"98",X"03",X"98",X"03",X"98",X"03",X"97",X"03",X"98",X"03",X"96",X"03",
		X"97",X"03",X"97",X"03",X"98",X"03",X"98",X"03",X"96",X"03",X"96",X"03",X"96",X"03",X"96",X"03",
		X"97",X"03",X"95",X"03",X"95",X"03",X"95",X"03",X"93",X"03",X"95",X"03",X"93",X"03",X"94",X"03",
		X"93",X"03",X"94",X"03",X"93",X"03",X"93",X"03",X"93",X"03",X"93",X"03",X"93",X"03",X"92",X"03",
		X"92",X"03",X"92",X"03",X"93",X"03",X"92",X"03",X"91",X"03",X"91",X"03",X"91",X"03",X"92",X"03",
		X"91",X"03",X"91",X"03",X"92",X"03",X"90",X"03",X"90",X"03",X"8E",X"03",X"8F",X"03",X"8F",X"03",
		X"8F",X"03",X"8E",X"03",X"8F",X"03",X"8E",X"03",X"8E",X"03",X"8E",X"03",X"8D",X"03",X"8D",X"03",
		X"8C",X"03",X"8D",X"03",X"8D",X"03",X"8C",X"03",X"8D",X"03",X"8B",X"03",X"8C",X"03",X"8A",X"03",
		X"8B",X"03",X"8B",X"03",X"8C",X"03",X"8A",X"03",X"8A",X"03",X"8A",X"03",X"8A",X"03",X"88",X"03",
		X"89",X"03",X"88",X"03",X"89",X"03",X"89",X"03",X"89",X"03",X"88",X"03",X"88",X"03",X"87",X"03",
		X"87",X"03",X"87",X"03",X"88",X"03",X"86",X"03",X"86",X"03",X"87",X"03",X"86",X"03",X"86",X"03",
		X"85",X"03",X"86",X"03",X"86",X"03",X"85",X"03",X"84",X"03",X"83",X"03",X"84",X"03",X"84",X"03",
		X"83",X"03",X"83",X"03",X"83",X"03",X"82",X"03",X"83",X"03",X"82",X"03",X"83",X"03",X"82",X"03",
		X"82",X"03",X"80",X"03",X"81",X"03",X"81",X"03",X"81",X"03",X"80",X"03",X"81",X"03",X"7F",X"03",
		X"80",X"03",X"7F",X"03",X"80",X"03",X"7F",X"03",X"7F",X"03",X"7F",X"03",X"7E",X"03",X"7E",X"03",
		X"7C",X"03",X"7C",X"03",X"7C",X"03",X"7D",X"03",X"7B",X"03",X"7D",X"03",X"7B",X"03",X"7B",X"03",
		X"7B",X"03",X"7B",X"03",X"7C",X"03",X"7B",X"03",X"7A",X"03",X"7A",X"03",X"7A",X"03",X"7A",X"03",
		X"79",X"03",X"79",X"03",X"78",X"03",X"79",X"03",X"78",X"03",X"79",X"03",X"78",X"03",X"77",X"03",
		X"77",X"03",X"77",X"03",X"77",X"03",X"75",X"03",X"75",X"03",X"76",X"03",X"76",X"03",X"76",X"03",
		X"75",X"03",X"76",X"03",X"76",X"03",X"74",X"03",X"74",X"03",X"74",X"03",X"73",X"03",X"73",X"03",
		X"73",X"03",X"73",X"03",X"72",X"03",X"71",X"03",X"72",X"03",X"72",X"03",X"72",X"03",X"71",X"03",
		X"71",X"03",X"70",X"03",X"70",X"03",X"70",X"03",X"71",X"03",X"70",X"03",X"70",X"03",X"6F",X"03",
		X"6F",X"03",X"6E",X"03",X"6D",X"03",X"6E",X"03",X"6D",X"03",X"6C",X"03",X"6D",X"03",X"6E",X"03",
		X"6C",X"03",X"6B",X"03",X"6C",X"03",X"6A",X"03",X"6B",X"03",X"6B",X"03",X"6B",X"03",X"6A",X"03",
		X"6A",X"03",X"6B",X"03",X"6B",X"03",X"6A",X"03",X"68",X"03",X"68",X"03",X"69",X"03",X"68",X"03",
		X"67",X"03",X"67",X"03",X"68",X"03",X"67",X"03",X"67",X"03",X"67",X"03",X"67",X"03",X"66",X"03",
		X"67",X"03",X"65",X"03",X"65",X"03",X"65",X"03",X"64",X"03",X"64",X"03",X"63",X"03",X"64",X"03",
		X"63",X"03",X"63",X"03",X"63",X"03",X"63",X"03",X"62",X"03",X"62",X"03",X"62",X"03",X"61",X"03",
		X"60",X"03",X"61",X"03",X"60",X"03",X"5F",X"03",X"60",X"03",X"61",X"03",X"5E",X"03",X"5F",X"03",
		X"60",X"03",X"5F",X"03",X"5F",X"03",X"5E",X"03",X"5D",X"03",X"5E",X"03",X"5D",X"03",X"5D",X"03",
		X"5D",X"03",X"5D",X"03",X"5C",X"03",X"5C",X"03",X"5C",X"03",X"5A",X"03",X"5B",X"03",X"5C",X"03",
		X"5A",X"03",X"5A",X"03",X"5B",X"03",X"5B",X"03",X"58",X"03",X"59",X"03",X"59",X"03",X"57",X"03",
		X"57",X"03",X"58",X"03",X"56",X"03",X"57",X"03",X"57",X"03",X"57",X"03",X"57",X"03",X"57",X"03",
		X"57",X"03",X"57",X"03",X"56",X"03",X"54",X"03",X"54",X"03",X"54",X"03",X"55",X"03",X"53",X"03",
		X"54",X"03",X"53",X"03",X"52",X"03",X"52",X"03",X"51",X"03",X"52",X"03",X"50",X"03",X"50",X"03",
		X"50",X"03",X"52",X"03",X"51",X"03",X"4F",X"03",X"4F",X"03",X"4F",X"03",X"4F",X"03",X"4F",X"03",
		X"4F",X"03",X"4F",X"03",X"4D",X"03",X"4E",X"03",X"4E",X"03",X"4D",X"03",X"4D",X"03",X"4D",X"03",
		X"4C",X"03",X"4C",X"03",X"4C",X"03",X"4C",X"03",X"4C",X"03",X"4B",X"03",X"4B",X"03",X"49",X"03",
		X"4B",X"03",X"4A",X"03",X"49",X"03",X"49",X"03",X"48",X"03",X"49",X"03",X"48",X"03",X"48",X"03",
		X"48",X"03",X"48",X"03",X"47",X"03",X"47",X"03",X"46",X"03",X"45",X"03",X"44",X"03",X"45",X"03",
		X"45",X"03",X"45",X"03",X"43",X"03",X"49",X"03",X"4C",X"03",X"4D",X"03",X"4B",X"03",X"4A",X"03",
		X"4B",X"03",X"4B",X"03",X"4A",X"03",X"49",X"03",X"4B",X"03",X"49",X"03",X"4A",X"03",X"49",X"03",
		X"49",X"03",X"48",X"03",X"4A",X"03",X"48",X"03",X"46",X"03",X"47",X"03",X"47",X"03",X"46",X"03",
		X"46",X"03",X"46",X"03",X"45",X"03",X"45",X"03",X"45",X"03",X"44",X"03",X"45",X"03",X"43",X"03",
		X"44",X"03",X"44",X"03",X"43",X"03",X"43",X"03",X"44",X"03",X"42",X"03",X"43",X"03",X"41",X"03",
		X"41",X"03",X"41",X"03",X"41",X"03",X"40",X"03",X"40",X"03",X"40",X"03",X"40",X"03",X"3F",X"03",
		X"3F",X"03",X"3F",X"03",X"3E",X"03",X"3E",X"03",X"3E",X"03",X"3E",X"03",X"3C",X"03",X"3E",X"03",
		X"3C",X"03",X"3C",X"03",X"3C",X"03",X"3C",X"03",X"3B",X"03",X"3B",X"03",X"3B",X"03",X"3B",X"03",
		X"3A",X"03",X"39",X"03",X"39",X"03",X"38",X"03",X"3A",X"03",X"38",X"03",X"39",X"03",X"38",X"03",
		X"37",X"03",X"37",X"03",X"38",X"03",X"36",X"03",X"36",X"03",X"36",X"03",X"35",X"03",X"35",X"03",
		X"34",X"03",X"35",X"03",X"34",X"03",X"34",X"03",X"34",X"03",X"33",X"03",X"34",X"03",X"34",X"03",
		X"32",X"03",X"32",X"03",X"32",X"03",X"32",X"03",X"31",X"03",X"31",X"03",X"31",X"03",X"30",X"03",
		X"30",X"03",X"31",X"03",X"2E",X"03",X"2F",X"03",X"2E",X"03",X"2E",X"03",X"2F",X"03",X"2D",X"03",
		X"2E",X"03",X"2E",X"03",X"2D",X"03",X"2D",X"03",X"2B",X"03",X"2C",X"03",X"2C",X"03",X"2A",X"03",
		X"2B",X"03",X"2B",X"03",X"2A",X"03",X"2A",X"03",X"2A",X"03",X"2A",X"03",X"2A",X"03",X"28",X"03",
		X"29",X"03",X"28",X"03",X"29",X"03",X"28",X"03",X"28",X"03",X"27",X"03",X"27",X"03",X"25",X"03",
		X"24",X"03",X"25",X"03",X"25",X"03",X"24",X"03",X"24",X"03",X"24",X"03",X"24",X"03",X"25",X"03",
		X"23",X"03",X"24",X"03",X"22",X"03",X"22",X"03",X"22",X"03",X"21",X"03",X"21",X"03",X"22",X"03",
		X"22",X"03",X"21",X"03",X"20",X"03",X"20",X"03",X"20",X"03",X"20",X"03",X"1F",X"03",X"20",X"03",
		X"1F",X"03",X"1E",X"03",X"1E",X"03",X"1E",X"03",X"1D",X"03",X"1D",X"03",X"1D",X"03",X"1E",X"03",
		X"1C",X"03",X"1B",X"03",X"1B",X"03",X"1B",X"03",X"1A",X"03",X"1B",X"03",X"19",X"03",X"1A",X"03",
		X"1A",X"03",X"18",X"03",X"19",X"03",X"19",X"03",X"18",X"03",X"18",X"03",X"18",X"03",X"18",X"03",
		X"16",X"03",X"17",X"03",X"16",X"03",X"16",X"03",X"17",X"03",X"16",X"03",X"14",X"03",X"15",X"03",
		X"16",X"03",X"14",X"03",X"14",X"03",X"13",X"03",X"13",X"03",X"13",X"03",X"13",X"03",X"13",X"03",
		X"13",X"03",X"12",X"03",X"11",X"03",X"11",X"03",X"12",X"03",X"10",X"03",X"0F",X"03",X"10",X"03",
		X"0F",X"03",X"0F",X"03",X"0F",X"03",X"0F",X"03",X"0E",X"03",X"0E",X"03",X"0F",X"03",X"0C",X"03",
		X"0D",X"03",X"0E",X"03",X"0B",X"03",X"0B",X"03",X"0C",X"03",X"0B",X"03",X"0B",X"03",X"0B",X"03",
		X"0A",X"03",X"0A",X"03",X"0B",X"03",X"09",X"03",X"09",X"03",X"09",X"03",X"09",X"03",X"08",X"03",
		X"09",X"03",X"08",X"03",X"07",X"03",X"07",X"03",X"08",X"03",X"07",X"03",X"06",X"03",X"08",X"03",
		X"05",X"03",X"05",X"03",X"05",X"03",X"04",X"03",X"03",X"03",X"04",X"03",X"05",X"03",X"04",X"03",
		X"03",X"03",X"04",X"03",X"04",X"03",X"03",X"03",X"02",X"03",X"03",X"03",X"01",X"03",X"02",X"03",
		X"00",X"03",X"00",X"03",X"00",X"03",X"FF",X"02",X"00",X"03",X"FE",X"02",X"FE",X"02",X"FD",X"02",
		X"FE",X"02",X"FE",X"02",X"FE",X"02",X"FD",X"02",X"FD",X"02",X"FC",X"02",X"FD",X"02",X"FD",X"02",
		X"FC",X"02",X"FA",X"02",X"FC",X"02",X"FB",X"02",X"FB",X"02",X"FA",X"02",X"FA",X"02",X"F9",X"02",
		X"FA",X"02",X"FA",X"02",X"F8",X"02",X"F9",X"02",X"F8",X"02",X"F7",X"02",X"F7",X"02",X"F8",X"02",
		X"F6",X"02",X"F6",X"02",X"F5",X"02",X"F5",X"02",X"F5",X"02",X"F5",X"02",X"F5",X"02",X"F3",X"02",
		X"F4",X"02",X"F4",X"02",X"F4",X"02",X"F2",X"02",X"F4",X"02",X"F3",X"02",X"F2",X"02",X"F2",X"02",
		X"F2",X"02",X"F1",X"02",X"F1",X"02",X"F1",X"02",X"F1",X"02",X"F0",X"02",X"EF",X"02",X"EF",X"02",
		X"EE",X"02",X"F0",X"02",X"EF",X"02",X"EF",X"02",X"EE",X"02",X"EE",X"02",X"ED",X"02",X"EE",X"02",
		X"EC",X"02",X"EC",X"02",X"ED",X"02",X"EC",X"02",X"EC",X"02",X"EB",X"02",X"EA",X"02",X"EA",X"02",
		X"EA",X"02",X"E9",X"02",X"E9",X"02",X"E8",X"02",X"EA",X"02",X"EA",X"02",X"E8",X"02",X"E8",X"02",
		X"E8",X"02",X"E8",X"02",X"E7",X"02",X"E7",X"02",X"E6",X"02",X"E6",X"02",X"E7",X"02",X"E6",X"02",
		X"E5",X"02",X"E5",X"02",X"E5",X"02",X"E4",X"02",X"E4",X"02",X"E5",X"02",X"E3",X"02",X"E3",X"02",
		X"E3",X"02",X"E1",X"02",X"E2",X"02",X"E3",X"02",X"E2",X"02",X"E0",X"02",X"E1",X"02",X"E1",X"02",
		X"E0",X"02",X"E0",X"02",X"E0",X"02",X"DE",X"02",X"DE",X"02",X"DE",X"02",X"DE",X"02",X"DC",X"02",
		X"DE",X"02",X"DE",X"02",X"DD",X"02",X"DD",X"02",X"DD",X"02",X"DC",X"02",X"DD",X"02",X"DC",X"02",
		X"DC",X"02",X"DA",X"02",X"DC",X"02",X"DB",X"02",X"DA",X"02",X"D9",X"02",X"D9",X"02",X"D9",X"02",
		X"D9",X"02",X"D9",X"02",X"D8",X"02",X"D7",X"02",X"D8",X"02",X"D7",X"02",X"D6",X"02",X"D8",X"02",
		X"D6",X"02",X"D7",X"02",X"D7",X"02",X"D6",X"02",X"D6",X"02",X"D5",X"02",X"D6",X"02",X"D4",X"02",
		X"D3",X"02",X"D3",X"02",X"D3",X"02",X"D3",X"02",X"D3",X"02",X"D2",X"02",X"D1",X"02",X"D3",X"02",
		X"D2",X"02",X"D2",X"02",X"D0",X"02",X"D0",X"02",X"D0",X"02",X"D0",X"02",X"D1",X"02",X"CF",X"02",
		X"D0",X"02",X"D0",X"02",X"CF",X"02",X"CF",X"02",X"CF",X"02",X"CE",X"02",X"CD",X"02",X"CE",X"02",
		X"CD",X"02",X"CD",X"02",X"CC",X"02",X"CC",X"02",X"CB",X"02",X"CB",X"02",X"CB",X"02",X"CB",X"02",
		X"CA",X"02",X"CA",X"02",X"C9",X"02",X"C9",X"02",X"CA",X"02",X"C9",X"02",X"C8",X"02",X"C8",X"02",
		X"C7",X"02",X"C6",X"02",X"C7",X"02",X"C6",X"02",X"C8",X"02",X"C6",X"02",X"C6",X"02",X"C6",X"02",
		X"C7",X"02",X"C5",X"02",X"C6",X"02",X"C4",X"02",X"C9",X"02",X"CB",X"02",X"CA",X"02",X"CB",X"02",
		X"CB",X"02",X"CA",X"02",X"C9",X"02",X"CA",X"02",X"CA",X"02",X"C9",X"02",X"C8",X"02",X"C7",X"02",
		X"C7",X"02",X"C8",X"02",X"C6",X"02",X"C7",X"02",X"C7",X"02",X"C5",X"02",X"C5",X"02",X"C4",X"02",
		X"C6",X"02",X"C5",X"02",X"C6",X"02",X"C4",X"02",X"C4",X"02",X"C5",X"02",X"C3",X"02",X"C3",X"02",
		X"C3",X"02",X"C2",X"02",X"C2",X"02",X"C2",X"02",X"C2",X"02",X"C1",X"02",X"C1",X"02",X"C3",X"02",
		X"C0",X"02",X"C0",X"02",X"BF",X"02",X"C1",X"02",X"BE",X"02",X"BE",X"02",X"BF",X"02",X"BE",X"02",
		X"BF",X"02",X"BE",X"02",X"BE",X"02",X"BD",X"02",X"BD",X"02",X"BC",X"02",X"BD",X"02",X"BD",X"02",
		X"BB",X"02",X"BB",X"02",X"BB",X"02",X"BB",X"02",X"BA",X"02",X"B9",X"02",X"BA",X"02",X"B9",X"02",
		X"B9",X"02",X"B9",X"02",X"B9",X"02",X"B8",X"02",X"B8",X"02",X"B8",X"02",X"B7",X"02",X"B7",X"02",
		X"B6",X"02",X"B6",X"02",X"B6",X"02",X"B6",X"02",X"B6",X"02",X"B5",X"02",X"B5",X"02",X"B4",X"02",
		X"B4",X"02",X"B4",X"02",X"B3",X"02",X"B3",X"02",X"B3",X"02",X"B3",X"02",X"B3",X"02",X"B3",X"02",
		X"B2",X"02",X"B3",X"02",X"B3",X"02",X"AF",X"02",X"B2",X"02",X"B1",X"02",X"B0",X"02",X"B0",X"02",
		X"B0",X"02",X"AE",X"02",X"AF",X"02",X"AF",X"02",X"AF",X"02",X"AE",X"02",X"AE",X"02",X"AE",X"02",
		X"AE",X"02",X"AD",X"02",X"AD",X"02",X"AC",X"02",X"AB",X"02",X"AB",X"02",X"AC",X"02",X"AC",X"02",
		X"AB",X"02",X"AC",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"A9",X"02",X"A8",X"02",X"A9",X"02",
		X"A9",X"02",X"A8",X"02",X"A8",X"02",X"A8",X"02",X"A7",X"02",X"A7",X"02",X"A6",X"02",X"A6",X"02",
		X"A6",X"02",X"A8",X"02",X"A6",X"02",X"A5",X"02",X"A5",X"02",X"A5",X"02",X"A4",X"02",X"A4",X"02",
		X"A3",X"02",X"A3",X"02",X"A3",X"02",X"A3",X"02",X"A3",X"02",X"A2",X"02",X"A1",X"02",X"A3",X"02",
		X"A1",X"02",X"A1",X"02",X"A0",X"02",X"A1",X"02",X"9F",X"02",X"A0",X"02",X"A0",X"02",X"9F",X"02",
		X"9F",X"02",X"9F",X"02",X"A0",X"02",X"9D",X"02",X"9E",X"02",X"9F",X"02",X"9D",X"02",X"9C",X"02",
		X"9D",X"02",X"9E",X"02",X"9C",X"02",X"9D",X"02",X"9C",X"02",X"9B",X"02",X"9A",X"02",X"9B",X"02",
		X"9A",X"02",X"9A",X"02",X"9B",X"02",X"9A",X"02",X"98",X"02",X"99",X"02",X"99",X"02",X"9A",X"02",
		X"97",X"02",X"99",X"02",X"97",X"02",X"97",X"02",X"97",X"02",X"98",X"02",X"96",X"02",X"95",X"02",
		X"96",X"02",X"97",X"02",X"95",X"02",X"95",X"02",X"94",X"02",X"94",X"02",X"94",X"02",X"94",X"02",
		X"94",X"02",X"94",X"02",X"93",X"02",X"93",X"02",X"91",X"02",X"92",X"02",X"93",X"02",X"92",X"02",
		X"91",X"02",X"92",X"02",X"91",X"02",X"90",X"02",X"90",X"02",X"8F",X"02",X"90",X"02",X"8E",X"02",
		X"8F",X"02",X"8F",X"02",X"8E",X"02",X"8F",X"02",X"8E",X"02",X"8D",X"02",X"8E",X"02",X"8E",X"02",
		X"8D",X"02",X"8C",X"02",X"8C",X"02",X"8C",X"02",X"8C",X"02",X"8C",X"02",X"8A",X"02",X"8B",X"02",
		X"8A",X"02",X"8B",X"02",X"8A",X"02",X"89",X"02",X"88",X"02",X"89",X"02",X"89",X"02",X"88",X"02",
		X"87",X"02",X"88",X"02",X"87",X"02",X"86",X"02",X"88",X"02",X"88",X"02",X"87",X"02",X"86",X"02",
		X"86",X"02",X"85",X"02",X"85",X"02",X"84",X"02",X"86",X"02",X"84",X"02",X"84",X"02",X"84",X"02",
		X"84",X"02",X"82",X"02",X"83",X"02",X"82",X"02",X"83",X"02",X"81",X"02",X"81",X"02",X"80",X"02",
		X"81",X"02",X"82",X"02",X"83",X"02",X"81",X"02",X"80",X"02",X"81",X"02",X"80",X"02",X"7F",X"02",
		X"80",X"02",X"7F",X"02",X"7E",X"02",X"7E",X"02",X"7F",X"02",X"7D",X"02",X"7D",X"02",X"7D",X"02",
		X"7E",X"02",X"7D",X"02",X"7C",X"02",X"7E",X"02",X"7B",X"02",X"7D",X"02",X"7B",X"02",X"7C",X"02",
		X"7B",X"02",X"7A",X"02",X"7A",X"02",X"7B",X"02",X"7A",X"02",X"78",X"02",X"79",X"02",X"79",X"02",
		X"79",X"02",X"79",X"02",X"78",X"02",X"78",X"02",X"77",X"02",X"78",X"02",X"77",X"02",X"76",X"02",
		X"75",X"02",X"75",X"02",X"74",X"02",X"74",X"02",X"75",X"02",X"75",X"02",X"75",X"02",X"73",X"02",
		X"75",X"02",X"75",X"02",X"73",X"02",X"72",X"02",X"74",X"02",X"72",X"02",X"73",X"02",X"72",X"02",
		X"73",X"02",X"71",X"02",X"71",X"02",X"71",X"02",X"70",X"02",X"70",X"02",X"71",X"02",X"70",X"02",
		X"6D",X"02",X"6E",X"02",X"6F",X"02",X"6F",X"02",X"6E",X"02",X"6E",X"02",X"6F",X"02",X"6F",X"02",
		X"6D",X"02",X"6D",X"02",X"6C",X"02",X"6C",X"02",X"6B",X"02",X"6C",X"02",X"6B",X"02",X"6A",X"02",
		X"6B",X"02",X"6B",X"02",X"6C",X"02",X"6A",X"02",X"6A",X"02",X"6B",X"02",X"69",X"02",X"69",X"02",
		X"69",X"02",X"68",X"02",X"67",X"02",X"68",X"02",X"68",X"02",X"68",X"02",X"68",X"02",X"66",X"02",
		X"66",X"02",X"67",X"02",X"66",X"02",X"67",X"02",X"66",X"02",X"64",X"02",X"64",X"02",X"66",X"02",
		X"64",X"02",X"64",X"02",X"64",X"02",X"63",X"02",X"64",X"02",X"62",X"02",X"63",X"02",X"62",X"02",
		X"63",X"02",X"62",X"02",X"62",X"02",X"61",X"02",X"62",X"02",X"61",X"02",X"61",X"02",X"60",X"02",
		X"61",X"02",X"60",X"02",X"5F",X"02",X"5E",X"02",X"5F",X"02",X"60",X"02",X"60",X"02",X"5D",X"02",
		X"5E",X"02",X"5E",X"02",X"5E",X"02",X"5C",X"02",X"5D",X"02",X"5C",X"02",X"5C",X"02",X"5B",X"02",
		X"5C",X"02",X"5D",X"02",X"5A",X"02",X"5A",X"02",X"5A",X"02",X"5A",X"02",X"5A",X"02",X"5A",X"02",
		X"5A",X"02",X"59",X"02",X"59",X"02",X"5A",X"02",X"59",X"02",X"58",X"02",X"57",X"02",X"58",X"02",
		X"58",X"02",X"58",X"02",X"57",X"02",X"57",X"02",X"57",X"02",X"57",X"02",X"56",X"02",X"57",X"02",
		X"55",X"02",X"56",X"02",X"56",X"02",X"54",X"02",X"54",X"02",X"55",X"02",X"54",X"02",X"55",X"02",
		X"53",X"02",X"54",X"02",X"54",X"02",X"54",X"02",X"53",X"02",X"53",X"02",X"52",X"02",X"53",X"02",
		X"50",X"02",X"52",X"02",X"51",X"02",X"51",X"02",X"50",X"02",X"50",X"02",X"4F",X"02",X"50",X"02",
		X"4F",X"02",X"50",X"02",X"4E",X"02",X"4E",X"02",X"4E",X"02",X"52",X"02",X"54",X"02",X"52",X"02",
		X"53",X"02",X"53",X"02",X"53",X"02",X"51",X"02",X"53",X"02",X"53",X"02",X"51",X"02",X"51",X"02",
		X"51",X"02",X"50",X"02",X"4F",X"02",X"4F",X"02",X"50",X"02",X"4F",X"02",X"4F",X"02",X"4F",X"02",
		X"4E",X"02",X"4E",X"02",X"4E",X"02",X"50",X"02",X"4E",X"02",X"4D",X"02",X"4D",X"02",X"4D",X"02",
		X"4C",X"02",X"4C",X"02",X"4C",X"02",X"4C",X"02",X"4B",X"02",X"4A",X"02",X"4B",X"02",X"4A",X"02",
		X"4A",X"02",X"4A",X"02",X"4B",X"02",X"4A",X"02",X"47",X"02",X"48",X"02",X"49",X"02",X"48",X"02",
		X"48",X"02",X"48",X"02",X"48",X"02",X"47",X"02",X"46",X"02",X"47",X"02",X"48",X"02",X"46",X"02",
		X"45",X"02",X"45",X"02",X"47",X"02",X"45",X"02",X"44",X"02",X"45",X"02",X"44",X"02",X"44",X"02",
		X"43",X"02",X"43",X"02",X"45",X"02",X"43",X"02",X"43",X"02",X"43",X"02",X"43",X"02",X"42",X"02",
		X"42",X"02",X"42",X"02",X"42",X"02",X"41",X"02",X"40",X"02",X"41",X"02",X"41",X"02",X"41",X"02",
		X"40",X"02",X"41",X"02",X"3F",X"02",X"3F",X"02",X"3F",X"02",X"3E",X"02",X"3D",X"02",X"3E",X"02",
		X"3E",X"02",X"3E",X"02",X"3E",X"02",X"3D",X"02",X"3E",X"02",X"3D",X"02",X"3C",X"02",X"3C",X"02",
		X"3C",X"02",X"3B",X"02",X"3B",X"02",X"3B",X"02",X"3A",X"02",X"3A",X"02",X"3A",X"02",X"3A",X"02",
		X"3A",X"02",X"3A",X"02",X"38",X"02",X"39",X"02",X"3A",X"02",X"38",X"02",X"38",X"02",X"38",X"02",
		X"38",X"02",X"38",X"02",X"37",X"02",X"38",X"02",X"38",X"02",X"35",X"02",X"36",X"02",X"36",X"02",
		X"36",X"02",X"35",X"02",X"36",X"02",X"35",X"02",X"37",X"02",X"34",X"02",X"34",X"02",X"34",X"02",
		X"34",X"02",X"34",X"02",X"33",X"02",X"33",X"02",X"33",X"02",X"34",X"02",X"33",X"02",X"32",X"02",
		X"33",X"02",X"31",X"02",X"31",X"02",X"31",X"02",X"31",X"02",X"30",X"02",X"31",X"02",X"30",X"02",
		X"31",X"02",X"2F",X"02",X"2F",X"02",X"2F",X"02",X"2F",X"02",X"2E",X"02",X"2E",X"02",X"2E",X"02",
		X"2E",X"02",X"2E",X"02",X"2C",X"02",X"2D",X"02",X"2D",X"02",X"2C",X"02",X"2C",X"02",X"2B",X"02",
		X"2D",X"02",X"2C",X"02",X"2B",X"02",X"2A",X"02",X"2C",X"02",X"2B",X"02",X"2A",X"02",X"2A",X"02",
		X"2A",X"02",X"29",X"02",X"29",X"02",X"29",X"02",X"2A",X"02",X"28",X"02",X"27",X"02",X"27",X"02",
		X"28",X"02",X"28",X"02",X"28",X"02",X"27",X"02",X"27",X"02",X"27",X"02",X"25",X"02",X"26",X"02",
		X"26",X"02",X"26",X"02",X"25",X"02",X"26",X"02",X"26",X"02",X"24",X"02",X"23",X"02",X"24",X"02",
		X"24",X"02",X"24",X"02",X"23",X"02",X"23",X"02",X"24",X"02",X"23",X"02",X"22",X"02",X"22",X"02",
		X"22",X"02",X"22",X"02",X"21",X"02",X"20",X"02",X"21",X"02",X"21",X"02",X"1F",X"02",X"21",X"02",
		X"20",X"02",X"20",X"02",X"1E",X"02",X"1F",X"02",X"20",X"02",X"1F",X"02",X"1F",X"02",X"1D",X"02",
		X"1D",X"02",X"1E",X"02",X"1D",X"02",X"1C",X"02",X"1D",X"02",X"1D",X"02",X"1D",X"02",X"1B",X"02",
		X"1C",X"02",X"1C",X"02",X"1B",X"02",X"1B",X"02",X"1B",X"02",X"1A",X"02",X"1B",X"02",X"1A",X"02",
		X"1C",X"02",X"1A",X"02",X"1A",X"02",X"19",X"02",X"1A",X"02",X"19",X"02",X"19",X"02",X"18",X"02",
		X"17",X"02",X"18",X"02",X"18",X"02",X"18",X"02",X"17",X"02",X"17",X"02",X"17",X"02",X"16",X"02",
		X"16",X"02",X"17",X"02",X"17",X"02",X"16",X"02",X"15",X"02",X"16",X"02",X"14",X"02",X"14",X"02",
		X"14",X"02",X"14",X"02",X"14",X"02",X"15",X"02",X"13",X"02",X"13",X"02",X"14",X"02",X"12",X"02",
		X"12",X"02",X"11",X"02",X"12",X"02",X"11",X"02",X"11",X"02",X"10",X"02",X"11",X"02",X"10",X"02",
		X"10",X"02",X"10",X"02",X"10",X"02",X"10",X"02",X"11",X"02",X"0F",X"02",X"0F",X"02",X"0F",X"02",
		X"0F",X"02",X"0D",X"02",X"0D",X"02",X"0F",X"02",X"0D",X"02",X"0C",X"02",X"0D",X"02",X"0D",X"02",
		X"0C",X"02",X"0C",X"02",X"0B",X"02",X"0B",X"02",X"0B",X"02",X"0C",X"02",X"0B",X"02",X"0A",X"02",
		X"0B",X"02",X"0B",X"02",X"0B",X"02",X"0A",X"02",X"0A",X"02",X"0A",X"02",X"0A",X"02",X"08",X"02",
		X"09",X"02",X"09",X"02",X"08",X"02",X"07",X"02",X"09",X"02",X"08",X"02",X"09",X"02",X"07",X"02",
		X"08",X"02",X"07",X"02",X"07",X"02",X"07",X"02",X"07",X"02",X"08",X"02",X"07",X"02",X"06",X"02",
		X"05",X"02",X"05",X"02",X"05",X"02",X"04",X"02",X"03",X"02",X"04",X"02",X"04",X"02",X"04",X"02",
		X"02",X"02",X"03",X"02",X"03",X"02",X"03",X"02",X"01",X"02",X"02",X"02",X"01",X"02",X"01",X"02",
		X"01",X"02",X"00",X"02",X"00",X"02",X"01",X"02",X"00",X"02",X"FF",X"01",X"00",X"02",X"01",X"02",
		X"00",X"02",X"FF",X"01",X"FF",X"01",X"FF",X"01",X"00",X"02",X"FF",X"01",X"FE",X"01",X"FF",X"01",
		X"FF",X"01",X"FF",X"01",X"FE",X"01",X"FD",X"01",X"FD",X"01",X"FD",X"01",X"FC",X"01",X"FC",X"01",
		X"FC",X"01",X"FC",X"01",X"FC",X"01",X"FA",X"01",X"FD",X"01",X"FB",X"01",X"FA",X"01",X"FA",X"01",
		X"FA",X"01",X"FA",X"01",X"FB",X"01",X"F9",X"01",X"FA",X"01",X"F8",X"01",X"F9",X"01",X"F9",X"01",
		X"F9",X"01",X"F9",X"01",X"F8",X"01",X"F9",X"01",X"F8",X"01",X"F7",X"01",X"F7",X"01",X"F7",X"01",
		X"F6",X"01",X"F6",X"01",X"F6",X"01",X"F6",X"01",X"F6",X"01",X"F4",X"01",X"F5",X"01",X"F5",X"01",
		X"F5",X"01",X"F5",X"01",X"F4",X"01",X"F4",X"01",X"F4",X"01",X"F4",X"01",X"F3",X"01",X"F3",X"01",
		X"F4",X"01",X"F3",X"01",X"F2",X"01",X"F1",X"01",X"F3",X"01",X"F2",X"01",X"F2",X"01",X"F1",X"01",
		X"F1",X"01",X"F2",X"01",X"F1",X"01",X"F0",X"01",X"F0",X"01",X"F0",X"01",X"F0",X"01",X"EE",X"01",
		X"EF",X"01",X"F0",X"01",X"EE",X"01",X"F0",X"01",X"EF",X"01",X"EE",X"01",X"EF",X"01",X"EE",X"01",
		X"EE",X"01",X"ED",X"01",X"ED",X"01",X"ED",X"01",X"EC",X"01",X"EC",X"01",X"EB",X"01",X"EC",X"01",
		X"EC",X"01",X"ED",X"01",X"EB",X"01",X"EB",X"01",X"EB",X"01",X"EA",X"01",X"EB",X"01",X"EA",X"01",
		X"EA",X"01",X"E9",X"01",X"EA",X"01",X"E8",X"01",X"E9",X"01",X"E9",X"01",X"EC",X"01",X"EE",X"01",
		X"EB",X"01",X"ED",X"01",X"EC",X"01",X"ED",X"01",X"EB",X"01",X"EC",X"01",X"EB",X"01",X"EA",X"01",
		X"EA",X"01",X"EB",X"01",X"EB",X"01",X"EC",X"01",X"EA",X"01",X"EA",X"01",X"EA",X"01",X"E9",X"01",
		X"E9",X"01",X"E9",X"01",X"E9",X"01",X"E9",X"01",X"E9",X"01",X"E8",X"01",X"E9",X"01",X"E9",X"01",
		X"E8",X"01",X"E9",X"01",X"E8",X"01",X"E6",X"01",X"E6",X"01",X"E7",X"01",X"E6",X"01",X"E5",X"01",
		X"E7",X"01",X"E8",X"01",X"E7",X"01",X"E5",X"01",X"E4",X"01",X"E5",X"01",X"E5",X"01",X"E4",X"01",
		X"E4",X"01",X"E5",X"01",X"E4",X"01",X"E4",X"01",X"E2",X"01",X"E3",X"01",X"E2",X"01",X"E2",X"01",
		X"E1",X"01",X"E3",X"01",X"E2",X"01",X"E2",X"01",X"E2",X"01",X"E2",X"01",X"E2",X"01",X"E2",X"01",
		X"E1",X"01",X"E0",X"01",X"E0",X"01",X"E0",X"01",X"E0",X"01",X"E0",X"01",X"DF",X"01",X"DF",X"01",
		X"DF",X"01",X"E0",X"01",X"DF",X"01",X"DD",X"01",X"DE",X"01",X"DE",X"01",X"DD",X"01",X"DD",X"01",
		X"DD",X"01",X"DE",X"01",X"DD",X"01",X"DC",X"01",X"DD",X"01",X"DC",X"01",X"DC",X"01",X"DB",X"01",
		X"DC",X"01",X"DB",X"01",X"DB",X"01",X"DA",X"01",X"DB",X"01",X"DA",X"01",X"D9",X"01",X"DA",X"01",
		X"DA",X"01",X"DA",X"01",X"D9",X"01",X"D9",X"01",X"D8",X"01",X"D9",X"01",X"D8",X"01",X"D8",X"01",
		X"DA",X"01",X"D8",X"01",X"D7",X"01",X"D8",X"01",X"D7",X"01",X"D6",X"01",X"D7",X"01",X"D7",X"01",
		X"D7",X"01",X"D5",X"01",X"D6",X"01",X"D6",X"01",X"D6",X"01",X"D5",X"01",X"D6",X"01",X"D5",X"01",
		X"D5",X"01",X"D5",X"01",X"D3",X"01",X"D4",X"01",X"D5",X"01",X"D4",X"01",X"D4",X"01",X"D2",X"01",
		X"D4",X"01",X"D2",X"01",X"D1",X"01",X"D2",X"01",X"D2",X"01",X"D2",X"01",X"D0",X"01",X"D1",X"01",
		X"D1",X"01",X"D1",X"01",X"D1",X"01",X"D0",X"01",X"D0",X"01",X"D0",X"01",X"D0",X"01",X"D0",X"01",
		X"CF",X"01",X"D1",X"01",X"CE",X"01",X"CF",X"01",X"CF",X"01",X"CF",X"01",X"CE",X"01",X"CE",X"01",
		X"CE",X"01",X"CF",X"01",X"CE",X"01",X"CC",X"01",X"CD",X"01",X"CD",X"01",X"CD",X"01",X"CD",X"01",
		X"CD",X"01",X"CC",X"01",X"CC",X"01",X"CB",X"01",X"CC",X"01",X"CB",X"01",X"CA",X"01",X"CB",X"01",
		X"CB",X"01",X"C9",X"01",X"CA",X"01",X"CA",X"01",X"CA",X"01",X"CA",X"01",X"CA",X"01",X"C9",X"01",
		X"CA",X"01",X"C9",X"01",X"C9",X"01",X"C8",X"01",X"C7",X"01",X"C7",X"01",X"C8",X"01",X"C7",X"01",
		X"C7",X"01",X"C7",X"01",X"C6",X"01",X"C6",X"01",X"C7",X"01",X"C5",X"01",X"C6",X"01",X"C6",X"01",
		X"C7",X"01",X"C5",X"01",X"C5",X"01",X"C6",X"01",X"C5",X"01",X"C5",X"01",X"C4",X"01",X"C3",X"01",
		X"C5",X"01",X"C5",X"01",X"C4",X"01",X"C4",X"01",X"C3",X"01",X"C3",X"01",X"C1",X"01",X"C3",X"01",
		X"C3",X"01",X"C2",X"01",X"C2",X"01",X"C3",X"01",X"C2",X"01",X"C1",X"01",X"C0",X"01",X"C0",X"01",
		X"C0",X"01",X"C1",X"01",X"BF",X"01",X"C0",X"01",X"C2",X"01",X"C0",X"01",X"C1",X"01",X"C0",X"01",
		X"BE",X"01",X"C0",X"01",X"C1",X"01",X"BF",X"01",X"BD",X"01",X"BF",X"01",X"BE",X"01",X"BE",X"01",
		X"BD",X"01",X"BE",X"01",X"BD",X"01",X"BE",X"01",X"BD",X"01",X"BD",X"01",X"BC",X"01",X"BB",X"01",
		X"BC",X"01",X"BB",X"01",X"BC",X"01",X"BA",X"01",X"BB",X"01",X"BB",X"01",X"BA",X"01",X"BB",X"01",
		X"BA",X"01",X"BA",X"01",X"BB",X"01",X"BA",X"01",X"BA",X"01",X"B9",X"01",X"B9",X"01",X"B8",X"01",
		X"B9",X"01",X"B9",X"01",X"B8",X"01",X"B9",X"01",X"B7",X"01",X"B8",X"01",X"B8",X"01",X"B6",X"01",
		X"B7",X"01",X"B8",X"01",X"B7",X"01",X"B8",X"01",X"B5",X"01",X"B6",X"01",X"B5",X"01",X"B7",X"01",
		X"B5",X"01",X"B5",X"01",X"B6",X"01",X"B5",X"01",X"B6",X"01",X"B4",X"01",X"B4",X"01",X"B4",X"01",
		X"B4",X"01",X"B4",X"01",X"B3",X"01",X"B3",X"01",X"B4",X"01",X"B2",X"01",X"B3",X"01",X"B2",X"01",
		X"B3",X"01",X"B2",X"01",X"B2",X"01",X"B3",X"01",X"B2",X"01",X"B1",X"01",X"B1",X"01",X"B1",X"01",
		X"B2",X"01",X"B2",X"01",X"B2",X"01",X"B0",X"01",X"B0",X"01",X"B0",X"01",X"B1",X"01",X"B0",X"01",
		X"AE",X"01",X"AF",X"01",X"AE",X"01",X"AE",X"01",X"AF",X"01",X"AE",X"01",X"AF",X"01",X"AE",X"01",
		X"AE",X"01",X"AD",X"01",X"AD",X"01",X"AD",X"01",X"AC",X"01",X"AC",X"01",X"AE",X"01",X"AC",X"01",
		X"AC",X"01",X"AC",X"01",X"AC",X"01",X"AB",X"01",X"AC",X"01",X"AB",X"01",X"AC",X"01",X"AA",X"01",
		X"AC",X"01",X"AA",X"01",X"AA",X"01",X"AA",X"01",X"AB",X"01",X"A9",X"01",X"A8",X"01",X"AA",X"01",
		X"A9",X"01",X"AA",X"01",X"A8",X"01",X"A8",X"01",X"A8",X"01",X"A8",X"01",X"A8",X"01",X"A9",X"01",
		X"A8",X"01",X"A7",X"01",X"A6",X"01",X"A6",X"01",X"A6",X"01",X"A7",X"01",X"A6",X"01",X"A7",X"01",
		X"A6",X"01",X"A7",X"01",X"A7",X"01",X"A5",X"01",X"A4",X"01",X"A4",X"01",X"A5",X"01",X"A5",X"01",
		X"A5",X"01",X"A5",X"01",X"A5",X"01",X"A5",X"01",X"A4",X"01",X"A4",X"01",X"A5",X"01",X"A3",X"01",
		X"A3",X"01",X"A3",X"01",X"A3",X"01",X"A2",X"01",X"A2",X"01",X"A2",X"01",X"A3",X"01",X"A2",X"01",
		X"A1",X"01",X"A0",X"01",X"A1",X"01",X"A1",X"01",X"A1",X"01",X"A0",X"01",X"A0",X"01",X"A1",X"01",
		X"9F",X"01",X"9F",X"01",X"9F",X"01",X"9E",X"01",X"9E",X"01",X"9F",X"01",X"9F",X"01",X"9F",X"01",
		X"9F",X"01",X"9E",X"01",X"9F",X"01",X"9D",X"01",X"9D",X"01",X"9C",X"01",X"9D",X"01",X"9D",X"01",
		X"9D",X"01",X"9D",X"01",X"9D",X"01",X"9C",X"01",X"9C",X"01",X"9B",X"01",X"9B",X"01",X"9B",X"01",
		X"9B",X"01",X"9C",X"01",X"9C",X"01",X"9C",X"01",X"9B",X"01",X"99",X"01",X"9A",X"01",X"99",X"01",
		X"9B",X"01",X"9A",X"01",X"9B",X"01",X"99",X"01",X"99",X"01",X"98",X"01",X"99",X"01",X"99",X"01",
		X"99",X"01",X"98",X"01",X"99",X"01",X"98",X"01",X"98",X"01",X"98",X"01",X"96",X"01",X"98",X"01",
		X"97",X"01",X"97",X"01",X"96",X"01",X"94",X"01",X"96",X"01",X"98",X"01",X"96",X"01",X"97",X"01",
		X"96",X"01",X"95",X"01",X"95",X"01",X"95",X"01",X"95",X"01",X"94",X"01",X"92",X"01",X"97",X"01",
		X"9A",X"01",X"99",X"01",X"98",X"01",X"98",X"01",X"97",X"01",X"98",X"01",X"97",X"01",X"97",X"01",
		X"97",X"01",X"96",X"01",X"97",X"01",X"96",X"01",X"96",X"01",X"97",X"01",X"96",X"01",X"95",X"01",
		X"94",X"01",X"96",X"01",X"96",X"01",X"95",X"01",X"94",X"01",X"93",X"01",X"95",X"01",X"94",X"01",
		X"94",X"01",X"92",X"01",X"93",X"01",X"94",X"01",X"93",X"01",X"93",X"01",X"93",X"01",X"92",X"01",
		X"92",X"01",X"93",X"01",X"90",X"01",X"91",X"01",X"91",X"01",X"91",X"01",X"91",X"01",X"91",X"01",
		X"91",X"01",X"90",X"01",X"90",X"01",X"91",X"01",X"90",X"01",X"90",X"01",X"90",X"01",X"90",X"01",
		X"8F",X"01",X"8F",X"01",X"90",X"01",X"8F",X"01",X"8F",X"01",X"8F",X"01",X"8F",X"01",X"8E",X"01",
		X"8E",X"01",X"8E",X"01",X"8E",X"01",X"8C",X"01",X"8D",X"01",X"8D",X"01",X"8E",X"01",X"8D",X"01",
		X"8D",X"01",X"8C",X"01",X"8B",X"01",X"8C",X"01",X"8C",X"01",X"8C",X"01",X"8B",X"01",X"8B",X"01",
		X"8B",X"01",X"8C",X"01",X"8A",X"01",X"8B",X"01",X"8A",X"01",X"8A",X"01",X"89",X"01",X"8B",X"01",
		X"89",X"01",X"89",X"01",X"88",X"01",X"8A",X"01",X"89",X"01",X"88",X"01",X"88",X"01",X"89",X"01",
		X"88",X"01",X"89",X"01",X"88",X"01",X"89",X"01",X"88",X"01",X"87",X"01",X"87",X"01",X"88",X"01",
		X"87",X"01",X"85",X"01",X"84",X"01",X"87",X"01",X"86",X"01",X"86",X"01",X"87",X"01",X"85",X"01",
		X"85",X"01",X"85",X"01",X"84",X"01",X"86",X"01",X"86",X"01",X"84",X"01",X"84",X"01",X"84",X"01",
		X"84",X"01",X"84",X"01",X"82",X"01",X"82",X"01",X"84",X"01",X"82",X"01",X"85",X"01",X"84",X"01",
		X"82",X"01",X"83",X"01",X"82",X"01",X"82",X"01",X"82",X"01",X"83",X"01",X"82",X"01",X"83",X"01",
		X"81",X"01",X"80",X"01",X"81",X"01",X"81",X"01",X"80",X"01",X"7F",X"01",X"80",X"01",X"81",X"01",
		X"81",X"01",X"81",X"01",X"7F",X"01",X"80",X"01",X"7F",X"01",X"7F",X"01",X"7F",X"01",X"7D",X"01",
		X"7E",X"01",X"7E",X"01",X"7E",X"01",X"7D",X"01",X"7E",X"01",X"7D",X"01",X"7D",X"01",X"7D",X"01",
		X"7D",X"01",X"7D",X"01",X"7C",X"01",X"7B",X"01",X"7B",X"01",X"7C",X"01",X"7C",X"01",X"7C",X"01",
		X"7C",X"01",X"7B",X"01",X"7B",X"01",X"7B",X"01",X"7B",X"01",X"7B",X"01",X"7A",X"01",X"79",X"01",
		X"7A",X"01",X"7A",X"01",X"7B",X"01",X"7C",X"01",X"78",X"01",X"7A",X"01",X"79",X"01",X"79",X"01",
		X"78",X"01",X"7A",X"01",X"78",X"01",X"78",X"01",X"79",X"01",X"78",X"01",X"77",X"01",X"77",X"01",
		X"76",X"01",X"76",X"01",X"77",X"01",X"76",X"01",X"78",X"01",X"78",X"01",X"76",X"01",X"75",X"01",
		X"76",X"01",X"76",X"01",X"77",X"01",X"76",X"01",X"75",X"01",X"75",X"01",X"75",X"01",X"75",X"01",
		X"75",X"01",X"75",X"01",X"74",X"01",X"73",X"01",X"75",X"01",X"73",X"01",X"73",X"01",X"74",X"01",
		X"73",X"01",X"72",X"01",X"73",X"01",X"74",X"01",X"73",X"01",X"72",X"01",X"72",X"01",X"72",X"01",
		X"72",X"01",X"72",X"01",X"73",X"01",X"71",X"01",X"71",X"01",X"71",X"01",X"71",X"01",X"71",X"01",
		X"70",X"01",X"72",X"01",X"71",X"01",X"70",X"01",X"71",X"01",X"70",X"01",X"70",X"01",X"6F",X"01",
		X"70",X"01",X"70",X"01",X"6F",X"01",X"6E",X"01",X"6F",X"01",X"6D",X"01",X"6F",X"01",X"6E",X"01",
		X"6D",X"01",X"6E",X"01",X"6E",X"01",X"6E",X"01",X"6E",X"01",X"6D",X"01",X"6C",X"01",X"6C",X"01",
		X"6D",X"01",X"6D",X"01",X"6C",X"01",X"6B",X"01",X"6C",X"01",X"6C",X"01",X"6C",X"01",X"6B",X"01",
		X"6B",X"01",X"6B",X"01",X"6B",X"01",X"6B",X"01",X"6B",X"01",X"6B",X"01",X"69",X"01",X"6A",X"01",
		X"6A",X"01",X"6A",X"01",X"6A",X"01",X"69",X"01",X"68",X"01",X"68",X"01",X"69",X"01",X"69",X"01",
		X"69",X"01",X"69",X"01",X"68",X"01",X"68",X"01",X"67",X"01",X"66",X"01",X"68",X"01",X"68",X"01",
		X"66",X"01",X"67",X"01",X"67",X"01",X"68",X"01",X"67",X"01",X"67",X"01",X"66",X"01",X"65",X"01",
		X"67",X"01",X"67",X"01",X"66",X"01",X"66",X"01",X"65",X"01",X"65",X"01",X"66",X"01",X"65",X"01",
		X"65",X"01",X"64",X"01",X"65",X"01",X"64",X"01",X"64",X"01",X"63",X"01",X"64",X"01",X"65",X"01",
		X"65",X"01",X"64",X"01",X"63",X"01",X"62",X"01",X"63",X"01",X"63",X"01",X"63",X"01",X"63",X"01",
		X"63",X"01",X"62",X"01",X"62",X"01",X"62",X"01",X"62",X"01",X"62",X"01",X"60",X"01",X"61",X"01",
		X"60",X"01",X"61",X"01",X"60",X"01",X"60",X"01",X"60",X"01",X"60",X"01",X"5F",X"01",X"5F",X"01",
		X"61",X"01",X"60",X"01",X"5F",X"01",X"5E",X"01",X"5E",X"01",X"5F",X"01",X"5E",X"01",X"5F",X"01",
		X"5E",X"01",X"5E",X"01",X"5D",X"01",X"5E",X"01",X"5F",X"01",X"5F",X"01",X"5E",X"01",X"5D",X"01",
		X"5D",X"01",X"5D",X"01",X"5D",X"01",X"5D",X"01",X"5C",X"01",X"5B",X"01",X"5C",X"01",X"5D",X"01",
		X"5D",X"01",X"5C",X"01",X"5B",X"01",X"5A",X"01",X"5A",X"01",X"5A",X"01",X"5B",X"01",X"5B",X"01",
		X"5B",X"01",X"5A",X"01",X"5A",X"01",X"5A",X"01",X"5B",X"01",X"5A",X"01",X"5B",X"01",X"5A",X"01",
		X"59",X"01",X"5A",X"01",X"58",X"01",X"5A",X"01",X"59",X"01",X"58",X"01",X"58",X"01",X"58",X"01",
		X"58",X"01",X"59",X"01",X"57",X"01",X"58",X"01",X"58",X"01",X"57",X"01",X"56",X"01",X"56",X"01",
		X"55",X"01",X"58",X"01",X"56",X"01",X"56",X"01",X"56",X"01",X"56",X"01",X"56",X"01",X"56",X"01",
		X"56",X"01",X"55",X"01",X"55",X"01",X"56",X"01",X"56",X"01",X"56",X"01",X"56",X"01",X"54",X"01",
		X"54",X"01",X"54",X"01",X"55",X"01",X"54",X"01",X"53",X"01",X"53",X"01",X"53",X"01",X"53",X"01",
		X"53",X"01",X"53",X"01",X"53",X"01",X"54",X"01",X"53",X"01",X"52",X"01",X"52",X"01",X"53",X"01",
		X"51",X"01",X"52",X"01",X"53",X"01",X"51",X"01",X"51",X"01",X"50",X"01",X"51",X"01",X"52",X"01",
		X"50",X"01",X"50",X"01",X"50",X"01",X"50",X"01",X"51",X"01",X"51",X"01",X"52",X"01",X"50",X"01",
		X"4F",X"01",X"4F",X"01",X"50",X"01",X"4F",X"01",X"50",X"01",X"50",X"01",X"4F",X"01",X"4C",X"01",
		X"50",X"01",X"52",X"01",X"51",X"01",X"52",X"01",X"51",X"01",X"52",X"01",X"53",X"01",X"50",X"01",
		X"50",X"01",X"50",X"01",X"50",X"01",X"50",X"01",X"4F",X"01",X"51",X"01",X"4F",X"01",X"4F",X"01",
		X"4F",X"01",X"4F",X"01",X"4F",X"01",X"4F",X"01",X"4F",X"01",X"4F",X"01",X"4D",X"01",X"4F",X"01",
		X"4E",X"01",X"4E",X"01",X"4F",X"01",X"4E",X"01",X"4D",X"01",X"4E",X"01",X"4C",X"01",X"4D",X"01",
		X"4D",X"01",X"4C",X"01",X"4D",X"01",X"4B",X"01",X"4D",X"01",X"4C",X"01",X"4B",X"01",X"4C",X"01",
		X"4C",X"01",X"4B",X"01",X"4B",X"01",X"4A",X"01",X"4B",X"01",X"4B",X"01",X"4A",X"01",X"49",X"01",
		X"49",X"01",X"4A",X"01",X"4B",X"01",X"49",X"01",X"4A",X"01",X"4B",X"01",X"4A",X"01",X"49",X"01",
		X"49",X"01",X"49",X"01",X"49",X"01",X"49",X"01",X"49",X"01",X"49",X"01",X"48",X"01",X"48",X"01",
		X"48",X"01",X"47",X"01",X"48",X"01",X"48",X"01",X"46",X"01",X"46",X"01",X"47",X"01",X"48",X"01",
		X"48",X"01",X"46",X"01",X"47",X"01",X"46",X"01",X"45",X"01",X"46",X"01",X"46",X"01",X"47",X"01",
		X"46",X"01",X"46",X"01",X"45",X"01",X"44",X"01",X"45",X"01",X"45",X"01",X"45",X"01",X"43",X"01",
		X"44",X"01",X"45",X"01",X"45",X"01",X"44",X"01",X"44",X"01",X"45",X"01",X"43",X"01",X"43",X"01",
		X"42",X"01",X"41",X"01",X"44",X"01",X"43",X"01",X"43",X"01",X"42",X"01",X"42",X"01",X"42",X"01",
		X"41",X"01",X"41",X"01",X"42",X"01",X"41",X"01",X"41",X"01",X"41",X"01",X"41",X"01",X"41",X"01",
		X"41",X"01",X"41",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"41",X"01",X"41",X"01",X"40",X"01",
		X"41",X"01",X"40",X"01",X"3E",X"01",X"3F",X"01",X"3F",X"01",X"3E",X"01",X"3F",X"01",X"3F",X"01",
		X"3E",X"01",X"3F",X"01",X"3E",X"01",X"3E",X"01",X"3D",X"01",X"3E",X"01",X"3E",X"01",X"3E",X"01",
		X"3D",X"01",X"3D",X"01",X"3D",X"01",X"3D",X"01",X"3E",X"01",X"3C",X"01",X"3B",X"01",X"3B",X"01",
		X"3C",X"01",X"3C",X"01",X"3C",X"01",X"3B",X"01",X"3D",X"01",X"3C",X"01",X"3A",X"01",X"3B",X"01",
		X"3B",X"01",X"3B",X"01",X"3B",X"01",X"3B",X"01",X"3A",X"01",X"3B",X"01",X"3B",X"01",X"39",X"01",
		X"3B",X"01",X"3A",X"01",X"3A",X"01",X"39",X"01",X"3A",X"01",X"37",X"01",X"39",X"01",X"39",X"01",
		X"3A",X"01",X"39",X"01",X"39",X"01",X"38",X"01",X"37",X"01",X"38",X"01",X"37",X"01",X"37",X"01",
		X"37",X"01",X"37",X"01",X"37",X"01",X"36",X"01",X"36",X"01",X"37",X"01",X"37",X"01",X"37",X"01",
		X"37",X"01",X"36",X"01",X"37",X"01",X"35",X"01",X"36",X"01",X"36",X"01",X"35",X"01",X"37",X"01",
		X"35",X"01",X"34",X"01",X"35",X"01",X"34",X"01",X"35",X"01",X"36",X"01",X"35",X"01",X"34",X"01",
		X"34",X"01",X"34",X"01",X"35",X"01",X"33",X"01",X"34",X"01",X"34",X"01",X"33",X"01",X"33",X"01",
		X"33",X"01",X"33",X"01",X"33",X"01",X"32",X"01",X"33",X"01",X"32",X"01",X"31",X"01",X"32",X"01",
		X"32",X"01",X"32",X"01",X"32",X"01",X"31",X"01",X"31",X"01",X"31",X"01",X"30",X"01",X"30",X"01",
		X"31",X"01",X"30",X"01",X"33",X"01",X"30",X"01",X"31",X"01",X"30",X"01",X"2F",X"01",X"2F",X"01",
		X"30",X"01",X"31",X"01",X"2E",X"01",X"30",X"01",X"30",X"01",X"2F",X"01",X"30",X"01",X"2F",X"01",
		X"2F",X"01",X"2F",X"01",X"2F",X"01",X"2D",X"01",X"2E",X"01",X"2E",X"01",X"2E",X"01",X"2F",X"01",
		X"2E",X"01",X"2C",X"01",X"2E",X"01",X"2D",X"01",X"2E",X"01",X"2D",X"01",X"2D",X"01",X"2E",X"01",
		X"2D",X"01",X"2C",X"01",X"2C",X"01",X"2C",X"01",X"2D",X"01",X"2C",X"01",X"2D",X"01",X"2C",X"01",
		X"2A",X"01",X"2B",X"01",X"2C",X"01",X"29",X"01",X"2B",X"01",X"2B",X"01",X"2B",X"01",X"2A",X"01",
		X"29",X"01",X"29",X"01",X"2A",X"01",X"2A",X"01",X"2B",X"01",X"29",X"01",X"29",X"01",X"29",X"01",
		X"29",X"01",X"29",X"01",X"2A",X"01",X"28",X"01",X"29",X"01",X"2B",X"01",X"28",X"01",X"28",X"01",
		X"28",X"01",X"29",X"01",X"27",X"01",X"27",X"01",X"26",X"01",X"28",X"01",X"28",X"01",X"28",X"01",
		X"26",X"01",X"27",X"01",X"28",X"01",X"27",X"01",X"27",X"01",X"26",X"01",X"26",X"01",X"26",X"01",
		X"25",X"01",X"25",X"01",X"26",X"01",X"25",X"01",X"26",X"01",X"25",X"01",X"24",X"01",X"27",X"01",
		X"26",X"01",X"24",X"01",X"25",X"01",X"25",X"01",X"24",X"01",X"23",X"01",X"24",X"01",X"24",X"01",
		X"24",X"01",X"24",X"01",X"24",X"01",X"26",X"01",X"23",X"01",X"23",X"01",X"23",X"01",X"22",X"01",
		X"23",X"01",X"23",X"01",X"24",X"01",X"22",X"01",X"22",X"01",X"22",X"01",X"23",X"01",X"22",X"01",
		X"22",X"01",X"22",X"01",X"22",X"01",X"21",X"01",X"22",X"01",X"20",X"01",X"21",X"01",X"21",X"01",
		X"21",X"01",X"21",X"01",X"21",X"01",X"20",X"01",X"1F",X"01",X"20",X"01",X"20",X"01",X"22",X"01",
		X"20",X"01",X"20",X"01",X"1F",X"01",X"20",X"01",X"21",X"01",X"1F",X"01",X"20",X"01",X"20",X"01",
		X"1F",X"01",X"1F",X"01",X"1E",X"01",X"1E",X"01",X"1E",X"01",X"1E",X"01",X"1E",X"01",X"1E",X"01",
		X"1D",X"01",X"1D",X"01",X"1D",X"01",X"1D",X"01",X"1E",X"01",X"1D",X"01",X"1D",X"01",X"1D",X"01",
		X"1D",X"01",X"1C",X"01",X"1B",X"01",X"1B",X"01",X"1B",X"01",X"1D",X"01",X"1C",X"01",X"1C",X"01",
		X"1C",X"01",X"1C",X"01",X"1C",X"01",X"1C",X"01",X"1B",X"01",X"1D",X"01",X"1B",X"01",X"1C",X"01",
		X"1B",X"01",X"1A",X"01",X"1A",X"01",X"1A",X"01",X"1A",X"01",X"19",X"01",X"19",X"01",X"1A",X"01",
		X"19",X"01",X"1A",X"01",X"19",X"01",X"19",X"01",X"19",X"01",X"18",X"01",X"18",X"01",X"18",X"01",
		X"18",X"01",X"17",X"01",X"18",X"01",X"18",X"01",X"16",X"01",X"19",X"01",X"18",X"01",X"18",X"01",
		X"17",X"01",X"17",X"01",X"17",X"01",X"17",X"01",X"17",X"01",X"16",X"01",X"17",X"01",X"18",X"01",
		X"16",X"01",X"15",X"01",X"16",X"01",X"16",X"01",X"16",X"01",X"16",X"01",X"17",X"01",X"17",X"01",
		X"14",X"01",X"15",X"01",X"15",X"01",X"16",X"01",X"15",X"01",X"15",X"01",X"14",X"01",X"16",X"01",
		X"14",X"01",X"16",X"01",X"17",X"01",X"16",X"01",X"17",X"01",X"18",X"01",X"16",X"01",X"15",X"01",
		X"16",X"01",X"16",X"01",X"16",X"01",X"16",X"01",X"16",X"01",X"16",X"01",X"14",X"01",X"15",X"01",
		X"15",X"01",X"14",X"01",X"15",X"01",X"14",X"01",X"15",X"01",X"15",X"01",X"14",X"01",X"14",X"01",
		X"14",X"01",X"14",X"01",X"15",X"01",X"15",X"01",X"15",X"01",X"14",X"01",X"13",X"01",X"14",X"01",
		X"13",X"01",X"11",X"01",X"12",X"01",X"13",X"01",X"14",X"01",X"13",X"01",X"12",X"01",X"12",X"01",
		X"12",X"01",X"12",X"01",X"13",X"01",X"12",X"01",X"12",X"01",X"12",X"01",X"11",X"01",X"12",X"01",
		X"12",X"01",X"10",X"01",X"11",X"01",X"10",X"01",X"12",X"01",X"10",X"01",X"11",X"01",X"10",X"01",
		X"10",X"01",X"11",X"01",X"10",X"01",X"10",X"01",X"10",X"01",X"10",X"01",X"0F",X"01",X"0F",X"01",
		X"0F",X"01",X"0F",X"01",X"10",X"01",X"10",X"01",X"10",X"01",X"0F",X"01",X"0F",X"01",X"0E",X"01",
		X"0E",X"01",X"0F",X"01",X"0F",X"01",X"0F",X"01",X"0D",X"01",X"0E",X"01",X"0E",X"01",X"0D",X"01",
		X"0D",X"01",X"0D",X"01",X"0D",X"01",X"0E",X"01",X"0D",X"01",X"0C",X"01",X"0D",X"01",X"0C",X"01",
		X"0B",X"01",X"0A",X"01",X"0B",X"01",X"0C",X"01",X"0B",X"01",X"0D",X"01",X"0D",X"01",X"0B",X"01",
		X"0B",X"01",X"0A",X"01",X"0B",X"01",X"0B",X"01",X"0B",X"01",X"0B",X"01",X"0A",X"01",X"0B",X"01",
		X"0A",X"01",X"0A",X"01",X"0B",X"01",X"09",X"01",X"0A",X"01",X"0A",X"01",X"09",X"01",X"09",X"01",
		X"0A",X"01",X"09",X"01",X"09",X"01",X"09",X"01",X"09",X"01",X"09",X"01",X"09",X"01",X"08",X"01",
		X"09",X"01",X"08",X"01",X"08",X"01",X"08",X"01",X"07",X"01",X"07",X"01",X"07",X"01",X"07",X"01",
		X"07",X"01",X"07",X"01",X"06",X"01",X"07",X"01",X"08",X"01",X"07",X"01",X"07",X"01",X"07",X"01",
		X"06",X"01",X"07",X"01",X"06",X"01",X"06",X"01",X"05",X"01",X"06",X"01",X"06",X"01",X"07",X"01",
		X"06",X"01",X"05",X"01",X"04",X"01",X"04",X"01",X"05",X"01",X"05",X"01",X"05",X"01",X"06",X"01",
		X"05",X"01",X"04",X"01",X"05",X"01",X"03",X"01",X"03",X"01",X"05",X"01",X"04",X"01",X"04",X"01",
		X"03",X"01",X"04",X"01",X"04",X"01",X"02",X"01",X"03",X"01",X"03",X"01",X"02",X"01",X"04",X"01",
		X"02",X"01",X"04",X"01",X"02",X"01",X"02",X"01",X"03",X"01",X"01",X"01",X"03",X"01",X"01",X"01",
		X"01",X"01",X"02",X"01",X"02",X"01",X"00",X"01",X"01",X"01",X"02",X"01",X"00",X"01",X"02",X"01",
		X"01",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",
		X"01",X"01",X"00",X"01",X"00",X"01",X"FF",X"00",X"00",X"01",X"FF",X"00",X"00",X"01",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"00",X"01",X"FF",X"00",X"FE",X"00",X"FE",X"00",X"FF",X"00",X"FD",X"00",
		X"FE",X"00",X"FE",X"00",X"FE",X"00",X"FE",X"00",X"FE",X"00",X"FE",X"00",X"FD",X"00",X"FD",X"00",
		X"FC",X"00",X"FD",X"00",X"FE",X"00",X"FE",X"00",X"FD",X"00",X"FE",X"00",X"FD",X"00",X"FC",X"00",
		X"FC",X"00",X"FB",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",X"FB",X"00",X"FA",X"00",
		X"FB",X"00",X"FC",X"00",X"FB",X"00",X"FB",X"00",X"FB",X"00",X"FC",X"00",X"FA",X"00",X"FB",X"00",
		X"FA",X"00",X"FA",X"00",X"FB",X"00",X"FA",X"00",X"FA",X"00",X"FA",X"00",X"FB",X"00",X"FA",X"00",
		X"F9",X"00",X"F9",X"00",X"FA",X"00",X"F9",X"00",X"F8",X"00",X"F9",X"00",X"F9",X"00",X"F9",X"00",
		X"F9",X"00",X"F7",X"00",X"F8",X"00",X"F8",X"00",X"F8",X"00",X"FA",X"00",X"F8",X"00",X"F8",X"00",
		X"F9",X"00",X"F8",X"00",X"F7",X"00",X"F7",X"00",X"F7",X"00",X"F8",X"00",X"F7",X"00",X"F7",X"00",
		X"F7",X"00",X"F7",X"00",X"F7",X"00",X"F7",X"00",X"F6",X"00",X"F6",X"00",X"F6",X"00",X"F5",X"00",
		X"F6",X"00",X"F5",X"00",X"F7",X"00",X"F7",X"00",X"F4",X"00",X"F5",X"00",X"F4",X"00",X"F4",X"00",
		X"F4",X"00",X"F5",X"00",X"F6",X"00",X"F5",X"00",X"F5",X"00",X"F4",X"00",X"F3",X"00",X"F4",X"00",
		X"F4",X"00",X"F5",X"00",X"F4",X"00",X"F4",X"00",X"F4",X"00",X"F4",X"00",X"F3",X"00",X"F3",X"00",
		X"F3",X"00",X"F3",X"00",X"F4",X"00",X"F2",X"00",X"F4",X"00",X"F3",X"00",X"F4",X"00",X"F2",X"00",
		X"F1",X"00",X"F2",X"00",X"F2",X"00",X"F2",X"00",X"F2",X"00",X"F2",X"00",X"F3",X"00",X"F1",X"00",
		X"F1",X"00",X"F2",X"00",X"F2",X"00",X"F2",X"00",X"F1",X"00",X"F1",X"00",X"F1",X"00",X"F0",X"00",
		X"F2",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"EE",X"00",X"F0",X"00",X"F1",X"00",
		X"F1",X"00",X"F2",X"00",X"EF",X"00",X"EF",X"00",X"EF",X"00",X"F0",X"00",X"EF",X"00",X"EF",X"00",
		X"EE",X"00",X"F0",X"00",X"EF",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",
		X"EE",X"00",X"EF",X"00",X"EE",X"00",X"EF",X"00",X"EE",X"00",X"EC",X"00",X"ED",X"00",X"EE",X"00",
		X"ED",X"00",X"EE",X"00",X"ED",X"00",X"EC",X"00",X"EE",X"00",X"ED",X"00",X"EC",X"00",X"EC",X"00",
		X"EB",X"00",X"EC",X"00",X"EC",X"00",X"EC",X"00",X"EB",X"00",X"EB",X"00",X"EC",X"00",X"EC",X"00",
		X"EB",X"00",X"EA",X"00",X"EA",X"00",X"ED",X"00",X"EB",X"00",X"EB",X"00",X"EB",X"00",X"EB",X"00",
		X"EB",X"00",X"EA",X"00",X"EA",X"00",X"E9",X"00",X"E9",X"00",X"EA",X"00",X"EB",X"00",X"EA",X"00",
		X"EB",X"00",X"EA",X"00",X"EA",X"00",X"E9",X"00",X"E8",X"00",X"E9",X"00",X"E9",X"00",X"E9",X"00",
		X"E9",X"00",X"E9",X"00",X"E9",X"00",X"E9",X"00",X"E8",X"00",X"E9",X"00",X"E8",X"00",X"E8",X"00",
		X"E8",X"00",X"E9",X"00",X"E8",X"00",X"E8",X"00",X"E8",X"00",X"E7",X"00",X"E7",X"00",X"E7",X"00",
		X"E6",X"00",X"E7",X"00",X"E7",X"00",X"E6",X"00",X"E7",X"00",X"E7",X"00",X"E7",X"00",X"E6",X"00",
		X"E6",X"00",X"E7",X"00",X"E5",X"00",X"E7",X"00",X"E6",X"00",X"E6",X"00",X"E5",X"00",X"E6",X"00",
		X"E5",X"00",X"E4",X"00",X"E6",X"00",X"E5",X"00",X"E5",X"00",X"E5",X"00",X"E5",X"00",X"E5",X"00",
		X"E5",X"00",X"E4",X"00",X"E6",X"00",X"E7",X"00",X"E7",X"00",X"E6",X"00",X"E6",X"00",X"E5",X"00",
		X"E6",X"00",X"E5",X"00",X"E6",X"00",X"E6",X"00",X"E7",X"00",X"E7",X"00",X"E5",X"00",X"E5",X"00",
		X"E3",X"00",X"E4",X"00",X"E5",X"00",X"E5",X"00",X"E5",X"00",X"E6",X"00",X"E5",X"00",X"E5",X"00",
		X"E3",X"00",X"E4",X"00",X"E5",X"00",X"E4",X"00",X"E4",X"00",X"E4",X"00",X"E4",X"00",X"E5",X"00",
		X"E4",X"00",X"E4",X"00",X"E3",X"00",X"E3",X"00",X"E3",X"00",X"E2",X"00",X"E3",X"00",X"E3",X"00",
		X"E3",X"00",X"E4",X"00",X"E2",X"00",X"E2",X"00",X"E3",X"00",X"E3",X"00",X"E2",X"00",X"E3",X"00",
		X"E2",X"00",X"E3",X"00",X"E2",X"00",X"E2",X"00",X"E2",X"00",X"E2",X"00",X"E0",X"00",X"E2",X"00",
		X"E1",X"00",X"E0",X"00",X"E2",X"00",X"E1",X"00",X"E1",X"00",X"E1",X"00",X"E0",X"00",X"DF",X"00",
		X"E1",X"00",X"E1",X"00",X"E0",X"00",X"E0",X"00",X"E1",X"00",X"E0",X"00",X"E0",X"00",X"E0",X"00",
		X"DE",X"00",X"DF",X"00",X"DF",X"00",X"DF",X"00",X"DE",X"00",X"DF",X"00",X"E0",X"00",X"DF",X"00",
		X"E0",X"00",X"DF",X"00",X"DF",X"00",X"DE",X"00",X"DE",X"00",X"DD",X"00",X"DE",X"00",X"DE",X"00",
		X"DE",X"00",X"DE",X"00",X"DE",X"00",X"DE",X"00",X"DD",X"00",X"DC",X"00",X"DC",X"00",X"DD",X"00",
		X"DB",X"00",X"DC",X"00",X"DC",X"00",X"DB",X"00",X"DD",X"00",X"DD",X"00",X"DC",X"00",X"DB",X"00",
		X"DB",X"00",X"DB",X"00",X"DC",X"00",X"DC",X"00",X"DC",X"00",X"DC",X"00",X"DD",X"00",X"DC",X"00",
		X"DC",X"00",X"DB",X"00",X"DA",X"00",X"DB",X"00",X"DB",X"00",X"DC",X"00",X"DB",X"00",X"DC",X"00",
		X"DC",X"00",X"DC",X"00",X"DA",X"00",X"DA",X"00",X"DB",X"00",X"DB",X"00",X"D9",X"00",X"D9",X"00",
		X"DA",X"00",X"DA",X"00",X"DB",X"00",X"DA",X"00",X"DA",X"00",X"DB",X"00",X"DA",X"00",X"D9",X"00",
		X"D9",X"00",X"D9",X"00",X"D9",X"00",X"D9",X"00",X"DA",X"00",X"D9",X"00",X"D8",X"00",X"D8",X"00",
		X"D8",X"00",X"D7",X"00",X"D8",X"00",X"D8",X"00",X"D7",X"00",X"D8",X"00",X"D8",X"00",X"D8",X"00",
		X"D8",X"00",X"D6",X"00",X"D7",X"00",X"D7",X"00",X"D8",X"00",X"D7",X"00",X"D8",X"00",X"D7",X"00",
		X"D8",X"00",X"D8",X"00",X"D7",X"00",X"D5",X"00",X"D5",X"00",X"D5",X"00",X"D6",X"00",X"D6",X"00",
		X"D6",X"00",X"D6",X"00",X"D6",X"00",X"D6",X"00",X"D6",X"00",X"D4",X"00",X"D5",X"00",X"D5",X"00",
		X"D5",X"00",X"D5",X"00",X"D5",X"00",X"D5",X"00",X"D5",X"00",X"D5",X"00",X"D4",X"00",X"D5",X"00",
		X"D4",X"00",X"D4",X"00",X"D5",X"00",X"D4",X"00",X"D4",X"00",X"D2",X"00",X"D4",X"00",X"D4",X"00",
		X"D4",X"00",X"D4",X"00",X"D4",X"00",X"D5",X"00",X"D3",X"00",X"D2",X"00",X"D3",X"00",X"D3",X"00",
		X"D2",X"00",X"D2",X"00",X"D2",X"00",X"D3",X"00",X"D2",X"00",X"D2",X"00",X"D2",X"00",X"D2",X"00",
		X"D0",X"00",X"D2",X"00",X"D2",X"00",X"D2",X"00",X"D2",X"00",X"D2",X"00",X"D2",X"00",X"D2",X"00",
		X"D1",X"00",X"D0",X"00",X"D1",X"00",X"D1",X"00",X"D2",X"00",X"D0",X"00",X"D1",X"00",X"D1",X"00",
		X"D1",X"00",X"D0",X"00",X"D1",X"00",X"D0",X"00",X"D0",X"00",X"D0",X"00",X"D0",X"00",X"D1",X"00",
		X"CF",X"00",X"CF",X"00",X"D1",X"00",X"CF",X"00",X"CF",X"00",X"D0",X"00",X"CE",X"00",X"CF",X"00",
		X"CF",X"00",X"CF",X"00",X"CF",X"00",X"CF",X"00",X"CF",X"00",X"CE",X"00",X"CF",X"00",X"CE",X"00",
		X"CE",X"00",X"CD",X"00",X"CD",X"00",X"CD",X"00",X"CE",X"00",X"CD",X"00",X"CE",X"00",X"CD",X"00",
		X"CD",X"00",X"CD",X"00",X"CD",X"00",X"CC",X"00",X"CC",X"00",X"CD",X"00",X"CD",X"00",X"CD",X"00",
		X"CE",X"00",X"CE",X"00",X"CE",X"00",X"CD",X"00",X"CB",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",
		X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CD",X"00",
		X"CB",X"00",X"CB",X"00",X"CA",X"00",X"CB",X"00",X"CB",X"00",X"CB",X"00",X"CC",X"00",X"CB",X"00",
		X"CC",X"00",X"CB",X"00",X"CA",X"00",X"CA",X"00",X"C9",X"00",X"CA",X"00",X"CA",X"00",X"CA",X"00",
		X"CA",X"00",X"C9",X"00",X"CB",X"00",X"CB",X"00",X"C8",X"00",X"C9",X"00",X"C9",X"00",X"C8",X"00",
		X"C9",X"00",X"C8",X"00",X"C8",X"00",X"C8",X"00",X"C9",X"00",X"C9",X"00",X"C8",X"00",X"C8",X"00",
		X"C8",X"00",X"C9",X"00",X"C8",X"00",X"C9",X"00",X"C7",X"00",X"CA",X"00",X"C8",X"00",X"C7",X"00",
		X"C8",X"00",X"C8",X"00",X"C8",X"00",X"C7",X"00",X"C7",X"00",X"C7",X"00",X"C7",X"00",X"C5",X"00",
		X"C6",X"00",X"C6",X"00",X"C7",X"00",X"C7",X"00",X"C7",X"00",X"C5",X"00",X"C7",X"00",X"C6",X"00",
		X"C7",X"00",X"C6",X"00",X"C5",X"00",X"C7",X"00",X"C6",X"00",X"C6",X"00",X"C6",X"00",X"C6",X"00",
		X"C6",X"00",X"C5",X"00",X"C5",X"00",X"C5",X"00",X"C4",X"00",X"C6",X"00",X"C5",X"00",X"C5",X"00",
		X"C5",X"00",X"C4",X"00",X"C5",X"00",X"C5",X"00",X"C4",X"00",X"C3",X"00",X"C4",X"00",X"C4",X"00",
		X"C4",X"00",X"C4",X"00",X"C4",X"00",X"C4",X"00",X"C5",X"00",X"C4",X"00",X"C2",X"00",X"C3",X"00",
		X"C3",X"00",X"C3",X"00",X"C4",X"00",X"C4",X"00",X"C3",X"00",X"C2",X"00",X"C4",X"00",X"C3",X"00",
		X"C4",X"00",X"C4",X"00",X"C2",X"00",X"C2",X"00",X"C1",X"00",X"C2",X"00",X"C2",X"00",X"C2",X"00",
		X"C2",X"00",X"C1",X"00",X"C3",X"00",X"C2",X"00",X"C3",X"00",X"C0",X"00",X"C1",X"00",X"C1",X"00",
		X"C0",X"00",X"C2",X"00",X"C0",X"00",X"C1",X"00",X"C0",X"00",X"C0",X"00",X"C1",X"00",X"C0",X"00",
		X"C1",X"00",X"BF",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C1",X"00",X"C1",X"00",X"C1",X"00",
		X"C0",X"00",X"C0",X"00",X"C0",X"00",X"BF",X"00",X"BF",X"00",X"BF",X"00",X"BF",X"00",X"BF",X"00",
		X"C0",X"00",X"BF",X"00",X"BF",X"00",X"C0",X"00",X"BF",X"00",X"BF",X"00",X"BE",X"00",X"BF",X"00",
		X"BE",X"00",X"BE",X"00",X"BF",X"00",X"C0",X"00",X"BE",X"00",X"BE",X"00",X"BE",X"00",X"BE",X"00",
		X"BD",X"00",X"BD",X"00",X"BD",X"00",X"BD",X"00",X"BC",X"00",X"BE",X"00",X"BE",X"00",X"BE",X"00",
		X"BD",X"00",X"BD",X"00",X"BD",X"00",X"BF",X"00",X"C1",X"00",X"C0",X"00",X"BF",X"00",X"BE",X"00",
		X"BF",X"00",X"BF",X"00",X"BD",X"00",X"BE",X"00",X"BE",X"00",X"BE",X"00",X"BE",X"00",X"BE",X"00",
		X"BE",X"00",X"BC",X"00",X"BC",X"00",X"BD",X"00",X"BC",X"00",X"BD",X"00",X"BD",X"00",X"BD",X"00",
		X"BE",X"00",X"BD",X"00",X"BD",X"00",X"BD",X"00",X"BD",X"00",X"BC",X"00",X"BC",X"00",X"BC",X"00",
		X"BB",X"00",X"BC",X"00",X"BD",X"00",X"BC",X"00",X"BC",X"00",X"BC",X"00",X"BC",X"00",X"BC",X"00",
		X"BC",X"00",X"BB",X"00",X"BB",X"00",X"BA",X"00",X"BA",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",
		X"BB",X"00",X"BB",X"00",X"BC",X"00",X"BB",X"00",X"BA",X"00",X"BA",X"00",X"BA",X"00",X"BA",X"00",
		X"BC",X"00",X"BA",X"00",X"BA",X"00",X"BA",X"00",X"BC",X"00",X"BA",X"00",X"B9",X"00",X"BA",X"00",
		X"B9",X"00",X"B9",X"00",X"B8",X"00",X"B9",X"00",X"BA",X"00",X"B9",X"00",X"BA",X"00",X"B9",X"00",
		X"B8",X"00",X"B9",X"00",X"B9",X"00",X"B9",X"00",X"B8",X"00",X"B9",X"00",X"B8",X"00",X"B9",X"00",
		X"B8",X"00",X"B9",X"00",X"B8",X"00",X"B7",X"00",X"B8",X"00",X"B7",X"00",X"B8",X"00",X"B8",X"00",
		X"B7",X"00",X"B8",X"00",X"B7",X"00",X"B7",X"00",X"B6",X"00",X"B7",X"00",X"B6",X"00",X"B7",X"00",
		X"B7",X"00",X"B7",X"00",X"B7",X"00",X"B6",X"00",X"B7",X"00",X"B6",X"00",X"B6",X"00",X"B6",X"00",
		X"B6",X"00",X"B5",X"00",X"B7",X"00",X"B5",X"00",X"B6",X"00",X"B6",X"00",X"B6",X"00",X"B5",X"00",
		X"B5",X"00",X"B5",X"00",X"B6",X"00",X"B4",X"00",X"B6",X"00",X"B4",X"00",X"B5",X"00",X"B5",X"00",
		X"B5",X"00",X"B4",X"00",X"B5",X"00",X"B4",X"00",X"B4",X"00",X"B4",X"00",X"B4",X"00",X"B3",X"00",
		X"B4",X"00",X"B3",X"00",X"B3",X"00",X"B3",X"00",X"B5",X"00",X"B4",X"00",X"B5",X"00",X"B4",X"00",
		X"B4",X"00",X"B3",X"00",X"B3",X"00",X"B3",X"00",X"B4",X"00",X"B4",X"00",X"B3",X"00",X"B3",X"00",
		X"B3",X"00",X"B2",X"00",X"B3",X"00",X"B2",X"00",X"B2",X"00",X"B2",X"00",X"B3",X"00",X"B1",X"00",
		X"B2",X"00",X"B1",X"00",X"B2",X"00",X"B3",X"00",X"B2",X"00",X"B3",X"00",X"B2",X"00",X"B2",X"00",
		X"B2",X"00",X"AF",X"00",X"B0",X"00",X"B1",X"00",X"B0",X"00",X"B0",X"00",X"B2",X"00",X"B0",X"00",
		X"B0",X"00",X"B1",X"00",X"B2",X"00",X"B1",X"00",X"B1",X"00",X"B0",X"00",X"B0",X"00",X"B1",X"00",
		X"AE",X"00",X"B0",X"00",X"AF",X"00",X"B0",X"00",X"B0",X"00",X"AF",X"00",X"B1",X"00",X"B0",X"00",
		X"AF",X"00",X"B0",X"00",X"B0",X"00",X"AE",X"00",X"AF",X"00",X"B0",X"00",X"AE",X"00",X"AF",X"00",
		X"AF",X"00",X"AF",X"00",X"AF",X"00",X"AF",X"00",X"B0",X"00",X"AF",X"00",X"AE",X"00",X"AD",X"00",
		X"AE",X"00",X"AD",X"00",X"AE",X"00",X"AE",X"00",X"AE",X"00",X"AF",X"00",X"AE",X"00",X"AE",X"00",
		X"AF",X"00",X"AE",X"00",X"AE",X"00",X"AD",X"00",X"AD",X"00",X"AD",X"00",X"AD",X"00",X"AD",X"00",
		X"AE",X"00",X"AD",X"00",X"AD",X"00",X"AD",X"00",X"AD",X"00",X"AC",X"00",X"AD",X"00",X"AD",X"00",
		X"AC",X"00",X"AD",X"00",X"AB",X"00",X"AC",X"00",X"AC",X"00",X"AC",X"00",X"AC",X"00",X"AD",X"00",
		X"AD",X"00",X"AC",X"00",X"AC",X"00",X"AC",X"00",X"AB",X"00",X"AC",X"00",X"AB",X"00",X"AA",X"00",
		X"AB",X"00",X"AB",X"00",X"AA",X"00",X"AB",X"00",X"AB",X"00",X"AA",X"00",X"AB",X"00",X"AB",X"00",
		X"AA",X"00",X"AA",X"00",X"AB",X"00",X"A9",X"00",X"AA",X"00",X"AA",X"00",X"A9",X"00",X"AA",X"00",
		X"AA",X"00",X"AB",X"00",X"A9",X"00",X"A9",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"A9",X"00",
		X"AA",X"00",X"A8",X"00",X"A9",X"00",X"A8",X"00",X"A8",X"00",X"A9",X"00",X"A9",X"00",X"A8",X"00",
		X"A8",X"00",X"A8",X"00",X"A9",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"00",X"A6",X"00",
		X"A7",X"00",X"A9",X"00",X"A7",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"00",X"A7",X"00",X"A8",X"00",
		X"A8",X"00",X"A7",X"00",X"A7",X"00",X"A7",X"00",X"A6",X"00",X"A7",X"00",X"A7",X"00",X"A8",X"00",
		X"A7",X"00",X"A7",X"00",X"A7",X"00",X"A7",X"00",X"A8",X"00",X"A7",X"00",X"A6",X"00",X"A7",X"00",
		X"A6",X"00",X"A6",X"00",X"A6",X"00",X"A6",X"00",X"A7",X"00",X"A6",X"00",X"A6",X"00",X"A6",X"00",
		X"A7",X"00",X"A5",X"00",X"A5",X"00",X"A3",X"00",X"A6",X"00",X"A5",X"00",X"A4",X"00",X"A5",X"00",
		X"A6",X"00",X"A4",X"00",X"A5",X"00",X"A5",X"00",X"A4",X"00",X"A6",X"00",X"A6",X"00",X"A5",X"00",
		X"A4",X"00",X"A5",X"00",X"A4",X"00",X"A5",X"00",X"A4",X"00",X"A4",X"00",X"A5",X"00",X"A4",X"00",
		X"A3",X"00",X"A4",X"00",X"A3",X"00",X"A4",X"00",X"A4",X"00",X"A4",X"00",X"A2",X"00",X"A3",X"00",
		X"A4",X"00",X"A3",X"00",X"A3",X"00",X"A3",X"00",X"A3",X"00",X"A3",X"00",X"A3",X"00",X"A3",X"00",
		X"A3",X"00",X"A2",X"00",X"A1",X"00",X"A3",X"00",X"A1",X"00",X"A2",X"00",X"A2",X"00",X"A3",X"00",
		X"A4",X"00",X"A2",X"00",X"A2",X"00",X"A2",X"00",X"A1",X"00",X"A2",X"00",X"A2",X"00",X"A2",X"00",
		X"A3",X"00",X"A2",X"00",X"A1",X"00",X"A1",X"00",X"A2",X"00",X"A0",X"00",X"A1",X"00",X"A1",X"00",
		X"A1",X"00",X"A1",X"00",X"9F",X"00",X"A1",X"00",X"A1",X"00",X"A1",X"00",X"A0",X"00",X"A0",X"00",
		X"A1",X"00",X"A1",X"00",X"A0",X"00",X"9F",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A1",X"00",
		X"A0",X"00",X"A0",X"00",X"A1",X"00",X"A0",X"00",X"A0",X"00",X"9F",X"00",X"9F",X"00",X"9F",X"00",
		X"9F",X"00",X"9E",X"00",X"A0",X"00",X"9F",X"00",X"9F",X"00",X"A0",X"00",X"9E",X"00",X"9F",X"00",
		X"A0",X"00",X"9F",X"00",X"9F",X"00",X"9D",X"00",X"9E",X"00",X"9E",X"00",X"9E",X"00",X"9D",X"00",
		X"9E",X"00",X"9D",X"00",X"9C",X"00",X"9E",X"00",X"9D",X"00",X"9D",X"00",X"9E",X"00",X"9D",X"00",
		X"9C",X"00",X"9D",X"00",X"9C",X"00",X"9D",X"00",X"9D",X"00",X"9C",X"00",X"9E",X"00",X"9D",X"00",
		X"9D",X"00",X"9C",X"00",X"9E",X"00",X"9D",X"00",X"9E",X"00",X"9D",X"00",X"9C",X"00",X"9C",X"00",
		X"9C",X"00",X"9C",X"00",X"9C",X"00",X"9D",X"00",X"9C",X"00",X"9C",X"00",X"9C",X"00",X"9B",X"00",
		X"9C",X"00",X"9D",X"00",X"9C",X"00",X"9E",X"00",X"9C",X"00",X"9C",X"00",X"9D",X"00",X"9C",X"00",
		X"9C",X"00",X"9C",X"00",X"9B",X"00",X"9B",X"00",X"9B",X"00",X"9C",X"00",X"9A",X"00",X"9C",X"00",
		X"9B",X"00",X"9B",X"00",X"9B",X"00",X"9A",X"00",X"9B",X"00",X"9B",X"00",X"99",X"00",X"9A",X"00",
		X"9B",X"00",X"99",X"00",X"9A",X"00",X"9A",X"00",X"9B",X"00",X"9A",X"00",X"9A",X"00",X"9C",X"00",
		X"99",X"00",X"9A",X"00",X"9A",X"00",X"9B",X"00",X"9B",X"00",X"99",X"00",X"99",X"00",X"99",X"00",
		X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",
		X"99",X"00",X"98",X"00",X"99",X"00",X"98",X"00",X"98",X"00",X"98",X"00",X"98",X"00",X"9A",X"00",
		X"98",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"96",X"00",X"99",X"00",X"99",X"00",X"97",X"00",
		X"98",X"00",X"97",X"00",X"98",X"00",X"97",X"00",X"96",X"00",X"98",X"00",X"97",X"00",X"97",X"00",
		X"96",X"00",X"96",X"00",X"96",X"00",X"98",X"00",X"97",X"00",X"97",X"00",X"97",X"00",X"96",X"00",
		X"96",X"00",X"96",X"00",X"97",X"00",X"97",X"00",X"96",X"00",X"96",X"00",X"97",X"00",X"96",X"00",
		X"96",X"00",X"96",X"00",X"96",X"00",X"96",X"00",X"96",X"00",X"96",X"00",X"96",X"00",X"95",X"00",
		X"94",X"00",X"95",X"00",X"95",X"00",X"95",X"00",X"94",X"00",X"95",X"00",X"95",X"00",X"95",X"00",
		X"95",X"00",X"94",X"00",X"96",X"00",X"95",X"00",X"95",X"00",X"94",X"00",X"94",X"00",X"92",X"00",
		X"94",X"00",X"94",X"00",X"96",X"00",X"94",X"00",X"94",X"00",X"94",X"00",X"93",X"00",X"94",X"00",
		X"94",X"00",X"94",X"00",X"94",X"00",X"93",X"00",X"93",X"00",X"93",X"00",X"93",X"00",X"91",X"00",
		X"93",X"00",X"92",X"00",X"92",X"00",X"93",X"00",X"92",X"00",X"92",X"00",X"92",X"00",X"93",X"00",
		X"93",X"00",X"94",X"00",X"92",X"00",X"94",X"00",X"92",X"00",X"92",X"00",X"93",X"00",X"92",X"00",
		X"92",X"00",X"92",X"00",X"92",X"00",X"92",X"00",X"92",X"00",X"93",X"00",X"92",X"00",X"92",X"00",
		X"92",X"00",X"92",X"00",X"91",X"00",X"91",X"00",X"90",X"00",X"90",X"00",X"90",X"00",X"91",X"00",
		X"92",X"00",X"92",X"00",X"91",X"00",X"91",X"00",X"91",X"00",X"91",X"00",X"91",X"00",X"91",X"00",
		X"92",X"00",X"91",X"00",X"90",X"00",X"90",X"00",X"90",X"00",X"8F",X"00",X"90",X"00",X"90",X"00",
		X"90",X"00",X"91",X"00",X"8F",X"00",X"90",X"00",X"90",X"00",X"90",X"00",X"90",X"00",X"90",X"00",
		X"90",X"00",X"8F",X"00",X"8F",X"00",X"8D",X"00",X"8E",X"00",X"8F",X"00",X"8F",X"00",X"8E",X"00",
		X"8F",X"00",X"8F",X"00",X"90",X"00",X"8F",X"00",X"8F",X"00",X"90",X"00",X"8F",X"00",X"8F",X"00",
		X"8F",X"00",X"8E",X"00",X"8E",X"00",X"8F",X"00",X"8E",X"00",X"8D",X"00",X"8E",X"00",X"8E",X"00",
		X"8E",X"00",X"8E",X"00",X"8F",X"00",X"8E",X"00",X"8E",X"00",X"8F",X"00",X"8E",X"00",X"8E",X"00",
		X"8C",X"00",X"8D",X"00",X"8D",X"00",X"8D",X"00",X"8D",X"00",X"8D",X"00",X"8C",X"00",X"8C",X"00",
		X"8D",X"00",X"8D",X"00",X"8D",X"00",X"8E",X"00",X"8D",X"00",X"8D",X"00",X"8E",X"00",X"8C",X"00",
		X"8C",X"00",X"8C",X"00",X"8C",X"00",X"8C",X"00",X"8C",X"00",X"8C",X"00",X"8C",X"00",X"8D",X"00",
		X"8C",X"00",X"8C",X"00",X"8C",X"00",X"8D",X"00",X"8C",X"00",X"8C",X"00",X"8B",X"00",X"8B",X"00",
		X"8A",X"00",X"8B",X"00",X"8C",X"00",X"8B",X"00",X"8B",X"00",X"8B",X"00",X"8A",X"00",X"8C",X"00",
		X"8B",X"00",X"8A",X"00",X"8B",X"00",X"8B",X"00",X"8B",X"00",X"8A",X"00",X"8A",X"00",X"8C",X"00",
		X"8B",X"00",X"89",X"00",X"8A",X"00",X"8A",X"00",X"8B",X"00",X"8A",X"00",X"8A",X"00",X"8A",X"00",
		X"8A",X"00",X"8A",X"00",X"8A",X"00",X"8B",X"00",X"8A",X"00",X"8A",X"00",X"89",X"00",X"89",X"00",
		X"8A",X"00",X"89",X"00",X"89",X"00",X"89",X"00",X"89",X"00",X"8A",X"00",X"8A",X"00",X"89",X"00",
		X"89",X"00",X"89",X"00",X"89",X"00",X"89",X"00",X"89",X"00",X"89",X"00",X"89",X"00",X"88",X"00",
		X"89",X"00",X"88",X"00",X"89",X"00",X"88",X"00",X"89",X"00",X"88",X"00",X"88",X"00",X"87",X"00",
		X"88",X"00",X"87",X"00",X"88",X"00",X"87",X"00",X"87",X"00",X"88",X"00",X"89",X"00",X"88",X"00",
		X"87",X"00",X"87",X"00",X"87",X"00",X"87",X"00",X"87",X"00",X"86",X"00",X"87",X"00",X"87",X"00",
		X"87",X"00",X"87",X"00",X"86",X"00",X"87",X"00",X"88",X"00",X"86",X"00",X"87",X"00",X"86",X"00",
		X"86",X"00",X"85",X"00",X"86",X"00",X"87",X"00",X"86",X"00",X"85",X"00",X"87",X"00",X"86",X"00",
		X"86",X"00",X"85",X"00",X"85",X"00",X"86",X"00",X"86",X"00",X"86",X"00",X"85",X"00",X"85",X"00",
		X"85",X"00",X"85",X"00",X"86",X"00",X"85",X"00",X"85",X"00",X"86",X"00",X"84",X"00",X"85",X"00",
		X"85",X"00",X"84",X"00",X"85",X"00",X"84",X"00",X"84",X"00",X"84",X"00",X"85",X"00",X"85",X"00",
		X"85",X"00",X"85",X"00",X"84",X"00",X"84",X"00",X"84",X"00",X"84",X"00",X"84",X"00",X"85",X"00",
		X"83",X"00",X"85",X"00",X"85",X"00",X"84",X"00",X"83",X"00",X"86",X"00",X"83",X"00",X"84",X"00",
		X"84",X"00",X"83",X"00",X"83",X"00",X"82",X"00",X"83",X"00",X"82",X"00",X"82",X"00",X"83",X"00",
		X"83",X"00",X"83",X"00",X"83",X"00",X"84",X"00",X"82",X"00",X"83",X"00",X"84",X"00",X"83",X"00",
		X"83",X"00",X"83",X"00",X"82",X"00",X"82",X"00",X"81",X"00",X"81",X"00",X"82",X"00",X"81",X"00",
		X"82",X"00",X"82",X"00",X"82",X"00",X"82",X"00",X"82",X"00",X"81",X"00",X"81",X"00",X"83",X"00",
		X"83",X"00",X"82",X"00",X"83",X"00",X"81",X"00",X"81",X"00",X"82",X"00",X"81",X"00",X"81",X"00",
		X"81",X"00",X"82",X"00",X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",
		X"81",X"00",X"81",X"00",X"81",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"81",X"00",
		X"80",X"00",X"81",X"00",X"80",X"00",X"7F",X"00",X"7F",X"00",X"7F",X"00",X"7F",X"00",X"7F",X"00",
		X"7F",X"00",X"80",X"00",X"7F",X"00",X"80",X"00",X"80",X"00",X"7F",X"00",X"7F",X"00",X"7F",X"00",
		X"80",X"00",X"7F",X"00",X"7F",X"00",X"7F",X"00",X"7F",X"00",X"7E",X"00",X"7F",X"00",X"7E",X"00",
		X"7F",X"00",X"80",X"00",X"7F",X"00",X"80",X"00",X"7E",X"00",X"80",X"00",X"7D",X"00",X"7E",X"00",
		X"7E",X"00",X"7E",X"00",X"7D",X"00",X"7E",X"00",X"7C",X"00",X"7F",X"00",X"7E",X"00",X"7E",X"00",
		X"7E",X"00",X"7E",X"00",X"7E",X"00",X"7E",X"00",X"7E",X"00",X"7E",X"00",X"7E",X"00",X"7D",X"00",
		X"7D",X"00",X"7E",X"00",X"7D",X"00",X"7D",X"00",X"7D",X"00",X"7D",X"00",X"7C",X"00",X"7D",X"00",
		X"7D",X"00",X"7D",X"00",X"7D",X"00",X"7D",X"00",X"7D",X"00",X"7C",X"00",X"7D",X"00",X"7D",X"00",
		X"7C",X"00",X"7D",X"00",X"7C",X"00",X"7C",X"00",X"7D",X"00",X"7D",X"00",X"7C",X"00",X"7C",X"00",
		X"7C",X"00",X"7C",X"00",X"7B",X"00",X"7C",X"00",X"7C",X"00",X"7E",X"00",X"7C",X"00",X"7B",X"00",
		X"7C",X"00",X"7C",X"00",X"7B",X"00",X"7B",X"00",X"7B",X"00",X"7B",X"00",X"7A",X"00",X"7B",X"00",
		X"7A",X"00",X"7B",X"00",X"7B",X"00",X"7B",X"00",X"7B",X"00",X"7B",X"00",X"7B",X"00",X"7B",X"00",
		X"7B",X"00",X"7B",X"00",X"7B",X"00",X"7B",X"00",X"7C",X"00",X"7B",X"00",X"7A",X"00",X"7A",X"00",
		X"78",X"00",X"7A",X"00",X"79",X"00",X"7B",X"00",X"7A",X"00",X"7A",X"00",X"7A",X"00",X"7B",X"00",
		X"7B",X"00",X"7B",X"00",X"7A",X"00",X"7B",X"00",X"7B",X"00",X"79",X"00",X"79",X"00",X"79",X"00",
		X"78",X"00",X"7A",X"00",X"79",X"00",X"78",X"00",X"79",X"00",X"7A",X"00",X"78",X"00",X"79",X"00",
		X"79",X"00",X"7A",X"00",X"79",X"00",X"78",X"00",X"79",X"00",X"7A",X"00",X"79",X"00",X"7A",X"00",
		X"7A",X"00",X"78",X"00",X"79",X"00",X"79",X"00",X"77",X"00",X"77",X"00",X"79",X"00",X"78",X"00",
		X"77",X"00",X"79",X"00",X"79",X"00",X"78",X"00",X"78",X"00",X"78",X"00",X"77",X"00",X"78",X"00",
		X"78",X"00",X"78",X"00",X"78",X"00",X"78",X"00",X"77",X"00",X"77",X"00",X"76",X"00",X"76",X"00",
		X"76",X"00",X"77",X"00",X"78",X"00",X"76",X"00",X"77",X"00",X"77",X"00",X"77",X"00",X"77",X"00",
		X"76",X"00",X"77",X"00",X"76",X"00",X"78",X"00",X"77",X"00",X"75",X"00",X"75",X"00",X"75",X"00",
		X"75",X"00",X"76",X"00",X"76",X"00",X"76",X"00",X"76",X"00",X"76",X"00",X"76",X"00",X"75",X"00",
		X"75",X"00",X"75",X"00",X"76",X"00",X"76",X"00",X"76",X"00",X"77",X"00",X"76",X"00",X"76",X"00",
		X"75",X"00",X"76",X"00",X"76",X"00",X"76",X"00",X"75",X"00",X"75",X"00",X"75",X"00",X"75",X"00",
		X"75",X"00",X"75",X"00",X"76",X"00",X"76",X"00",X"75",X"00",X"76",X"00",X"76",X"00",X"75",X"00",
		X"75",X"00",X"75",X"00",X"75",X"00",X"74",X"00",X"74",X"00",X"75",X"00",X"74",X"00",X"73",X"00",
		X"74",X"00",X"75",X"00",X"73",X"00",X"75",X"00",X"75",X"00",X"74",X"00",X"73",X"00",X"73",X"00",
		X"73",X"00",X"74",X"00",X"73",X"00",X"74",X"00",X"74",X"00",X"73",X"00",X"73",X"00",X"73",X"00",
		X"74",X"00",X"73",X"00",X"73",X"00",X"73",X"00",X"73",X"00",X"73",X"00",X"73",X"00",X"75",X"00",
		X"73",X"00",X"71",X"00",X"73",X"00",X"73",X"00",X"73",X"00",X"74",X"00",X"73",X"00",X"73",X"00",
		X"73",X"00",X"72",X"00",X"72",X"00",X"72",X"00",X"72",X"00",X"72",X"00",X"72",X"00",X"73",X"00",
		X"71",X"00",X"71",X"00",X"71",X"00",X"71",X"00",X"72",X"00",X"71",X"00",X"72",X"00",X"72",X"00",
		X"72",X"00",X"73",X"00",X"72",X"00",X"72",X"00",X"71",X"00",X"71",X"00",X"70",X"00",X"70",X"00",
		X"70",X"00",X"70",X"00",X"71",X"00",X"70",X"00",X"71",X"00",X"72",X"00",X"72",X"00",X"71",X"00",
		X"71",X"00",X"73",X"00",X"71",X"00",X"71",X"00",X"72",X"00",X"72",X"00",X"71",X"00",X"71",X"00",
		X"70",X"00",X"70",X"00",X"70",X"00",X"70",X"00",X"70",X"00",X"70",X"00",X"70",X"00",X"70",X"00",
		X"6F",X"00",X"6F",X"00",X"71",X"00",X"6F",X"00",X"70",X"00",X"71",X"00",X"70",X"00",X"70",X"00",
		X"70",X"00",X"6F",X"00",X"70",X"00",X"70",X"00",X"70",X"00",X"6E",X"00",X"6D",X"00",X"6E",X"00",
		X"6E",X"00",X"6E",X"00",X"6F",X"00",X"6F",X"00",X"6F",X"00",X"6E",X"00",X"6F",X"00",X"6F",X"00",
		X"6F",X"00",X"6F",X"00",X"6F",X"00",X"71",X"00",X"6F",X"00",X"6E",X"00",X"6F",X"00",X"6F",X"00",
		X"6E",X"00",X"6F",X"00",X"6D",X"00",X"6E",X"00",X"6E",X"00",X"6E",X"00",X"6E",X"00",X"6E",X"00",
		X"6F",X"00",X"6E",X"00",X"6E",X"00",X"6D",X"00",X"6F",X"00",X"6E",X"00",X"6D",X"00",X"6F",X"00",
		X"6E",X"00",X"6E",X"00",X"6D",X"00",X"6D",X"00",X"6C",X"00",X"6D",X"00",X"6D",X"00",X"6D",X"00",
		X"6C",X"00",X"6E",X"00",X"6D",X"00",X"6D",X"00",X"6E",X"00",X"6E",X"00",X"6E",X"00",X"6C",X"00",
		X"6D",X"00",X"6D",X"00",X"6C",X"00",X"6D",X"00",X"6B",X"00",X"6D",X"00",X"6D",X"00",X"6D",X"00",
		X"6B",X"00",X"6B",X"00",X"6D",X"00",X"6D",X"00",X"6C",X"00",X"6C",X"00",X"6D",X"00",X"6C",X"00",
		X"6C",X"00",X"6C",X"00",X"6C",X"00",X"6C",X"00",X"6C",X"00",X"6C",X"00",X"6C",X"00",X"6D",X"00",
		X"6C",X"00",X"6B",X"00",X"6D",X"00",X"6B",X"00",X"6A",X"00",X"6B",X"00",X"6C",X"00",X"6A",X"00",
		X"6B",X"00",X"6B",X"00",X"6D",X"00",X"6C",X"00",X"6D",X"00",X"6C",X"00",X"6B",X"00",X"6B",X"00",
		X"6B",X"00",X"6B",X"00",X"6A",X"00",X"6B",X"00",X"6C",X"00",X"6B",X"00",X"6C",X"00",X"6A",X"00",
		X"6A",X"00",X"69",X"00",X"69",X"00",X"69",X"00",X"6A",X"00",X"69",X"00",X"6A",X"00",X"69",X"00",
		X"69",X"00",X"6B",X"00",X"69",X"00",X"69",X"00",X"6B",X"00",X"69",X"00",X"69",X"00",X"6B",X"00",
		X"68",X"00",X"6A",X"00",X"69",X"00",X"6A",X"00",X"69",X"00",X"69",X"00",X"69",X"00",X"6A",X"00",
		X"69",X"00",X"69",X"00",X"6A",X"00",X"6B",X"00",X"68",X"00",X"69",X"00",X"6A",X"00",X"68",X"00",
		X"69",X"00",X"69",X"00",X"6A",X"00",X"69",X"00",X"6A",X"00",X"69",X"00",X"68",X"00",X"6A",X"00",
		X"69",X"00",X"69",X"00",X"67",X"00",X"69",X"00",X"68",X"00",X"69",X"00",X"68",X"00",X"68",X"00",
		X"67",X"00",X"68",X"00",X"6A",X"00",X"69",X"00",X"68",X"00",X"68",X"00",X"67",X"00",X"68",X"00",
		X"67",X"00",X"68",X"00",X"68",X"00",X"68",X"00",X"68",X"00",X"68",X"00",X"68",X"00",X"68",X"00",
		X"67",X"00",X"67",X"00",X"67",X"00",X"67",X"00",X"66",X"00",X"68",X"00",X"68",X"00",X"67",X"00",
		X"67",X"00",X"67",X"00",X"67",X"00",X"67",X"00",X"68",X"00",X"67",X"00",X"67",X"00",X"68",X"00",
		X"67",X"00",X"68",X"00",X"68",X"00",X"67",X"00",X"67",X"00",X"65",X"00",X"65",X"00",X"67",X"00",
		X"66",X"00",X"67",X"00",X"68",X"00",X"67",X"00",X"68",X"00",X"66",X"00",X"66",X"00",X"66",X"00",
		X"66",X"00",X"67",X"00",X"67",X"00",X"67",X"00",X"67",X"00",X"66",X"00",X"66",X"00",X"66",X"00",
		X"66",X"00",X"66",X"00",X"65",X"00",X"64",X"00",X"65",X"00",X"65",X"00",X"65",X"00",X"64",X"00",
		X"65",X"00",X"65",X"00",X"65",X"00",X"65",X"00",X"65",X"00",X"66",X"00",X"66",X"00",X"65",X"00",
		X"65",X"00",X"65",X"00",X"65",X"00",X"65",X"00",X"65",X"00",X"65",X"00",X"65",X"00",X"64",X"00",
		X"64",X"00",X"63",X"00",X"64",X"00",X"65",X"00",X"63",X"00",X"64",X"00",X"64",X"00",X"63",X"00",
		X"65",X"00",X"65",X"00",X"65",X"00",X"64",X"00",X"64",X"00",X"64",X"00",X"63",X"00",X"64",X"00",
		X"64",X"00",X"64",X"00",X"64",X"00",X"65",X"00",X"64",X"00",X"62",X"00",X"63",X"00",X"63",X"00",
		X"63",X"00",X"63",X"00",X"62",X"00",X"63",X"00",X"63",X"00",X"63",X"00",X"63",X"00",X"64",X"00",
		X"63",X"00",X"62",X"00",X"61",X"00",X"63",X"00",X"63",X"00",X"63",X"00",X"63",X"00",X"63",X"00",
		X"62",X"00",X"64",X"00",X"64",X"00",X"61",X"00",X"63",X"00",X"61",X"00",X"61",X"00",X"60",X"00",
		X"62",X"00",X"62",X"00",X"61",X"00",X"62",X"00",X"62",X"00",X"64",X"00",X"62",X"00",X"64",X"00",
		X"63",X"00",X"62",X"00",X"62",X"00",X"62",X"00",X"62",X"00",X"63",X"00",X"61",X"00",X"63",X"00",
		X"62",X"00",X"61",X"00",X"61",X"00",X"61",X"00",X"61",X"00",X"61",X"00",X"61",X"00",X"61",X"00",
		X"61",X"00",X"61",X"00",X"62",X"00",X"61",X"00",X"61",X"00",X"60",X"00",X"61",X"00",X"61",X"00",
		X"61",X"00",X"61",X"00",X"61",X"00",X"61",X"00",X"61",X"00",X"60",X"00",X"61",X"00",X"61",X"00",
		X"61",X"00",X"60",X"00",X"60",X"00",X"5F",X"00",X"61",X"00",X"60",X"00",X"60",X"00",X"60",X"00",
		X"60",X"00",X"61",X"00",X"61",X"00",X"60",X"00",X"5F",X"00",X"60",X"00",X"5F",X"00",X"61",X"00",
		X"61",X"00",X"60",X"00",X"61",X"00",X"61",X"00",X"61",X"00",X"5F",X"00",X"62",X"00",X"60",X"00",
		X"5E",X"00",X"60",X"00",X"5F",X"00",X"5F",X"00",X"5F",X"00",X"5F",X"00",X"5E",X"00",X"5E",X"00",
		X"5F",X"00",X"5F",X"00",X"60",X"00",X"5E",X"00",X"5F",X"00",X"5F",X"00",X"5F",X"00",X"5E",X"00",
		X"60",X"00",X"5E",X"00",X"61",X"00",X"60",X"00",X"5E",X"00",X"5F",X"00",X"5F",X"00",X"60",X"00",
		X"5E",X"00",X"5E",X"00",X"5E",X"00",X"5F",X"00",X"5E",X"00",X"5E",X"00",X"5E",X"00",X"5C",X"00",
		X"5D",X"00",X"5D",X"00",X"5F",X"00",X"5E",X"00",X"5E",X"00",X"5E",X"00",X"5E",X"00",X"5E",X"00",
		X"5F",X"00",X"5F",X"00",X"5D",X"00",X"5E",X"00",X"5E",X"00",X"5E",X"00",X"5D",X"00",X"5D",X"00",
		X"5D",X"00",X"5E",X"00",X"5D",X"00",X"5F",X"00",X"5E",X"00",X"5E",X"00",X"5E",X"00",X"5D",X"00",
		X"5E",X"00",X"5C",X"00",X"5E",X"00",X"5D",X"00",X"5D",X"00",X"5B",X"00",X"5D",X"00",X"5C",X"00",
		X"5D",X"00",X"5C",X"00",X"5D",X"00",X"5D",X"00",X"5C",X"00",X"5C",X"00",X"5D",X"00",X"5C",X"00",
		X"5B",X"00",X"5C",X"00",X"5B",X"00",X"5D",X"00",X"5B",X"00",X"5B",X"00",X"5D",X"00",X"5B",X"00",
		X"5D",X"00",X"5C",X"00",X"5C",X"00",X"5D",X"00",X"5D",X"00",X"5C",X"00",X"5C",X"00",X"5B",X"00",
		X"5C",X"00",X"5D",X"00",X"5C",X"00",X"5D",X"00",X"5A",X"00",X"5B",X"00",X"5B",X"00",X"5B",X"00",
		X"5B",X"00",X"5C",X"00",X"5B",X"00",X"5B",X"00",X"5A",X"00",X"5B",X"00",X"5B",X"00",X"5B",X"00",
		X"5C",X"00",X"5B",X"00",X"5A",X"00",X"5D",X"00",X"5B",X"00",X"5B",X"00",X"5B",X"00",X"5B",X"00",
		X"5A",X"00",X"5A",X"00",X"5A",X"00",X"5B",X"00",X"5B",X"00",X"5A",X"00",X"5A",X"00",X"5A",X"00",
		X"5B",X"00",X"5A",X"00",X"5A",X"00",X"5A",X"00",X"5A",X"00",X"5A",X"00",X"5A",X"00",X"5B",X"00",
		X"5A",X"00",X"5A",X"00",X"5B",X"00",X"5A",X"00",X"5A",X"00",X"5B",X"00",X"5A",X"00",X"5A",X"00",
		X"5A",X"00",X"5A",X"00",X"5A",X"00",X"5A",X"00",X"5A",X"00",X"59",X"00",X"58",X"00",X"59",X"00",
		X"59",X"00",X"59",X"00",X"59",X"00",X"59",X"00",X"59",X"00",X"59",X"00",X"59",X"00",X"58",X"00",
		X"58",X"00",X"59",X"00",X"59",X"00",X"59",X"00",X"59",X"00",X"58",X"00",X"59",X"00",X"58",X"00",
		X"58",X"00",X"5A",X"00",X"58",X"00",X"5A",X"00",X"59",X"00",X"59",X"00",X"59",X"00",X"58",X"00",
		X"58",X"00",X"58",X"00",X"57",X"00",X"58",X"00",X"58",X"00",X"58",X"00",X"58",X"00",X"58",X"00",
		X"57",X"00",X"56",X"00",X"58",X"00",X"58",X"00",X"57",X"00",X"58",X"00",X"58",X"00",X"58",X"00",
		X"57",X"00",X"58",X"00",X"59",X"00",X"59",X"00",X"58",X"00",X"58",X"00",X"58",X"00",X"58",X"00",
		X"57",X"00",X"57",X"00",X"57",X"00",X"57",X"00",X"57",X"00",X"57",X"00",X"58",X"00",X"58",X"00",
		X"58",X"00",X"57",X"00",X"58",X"00",X"57",X"00",X"57",X"00",X"55",X"00",X"57",X"00",X"57",X"00",
		X"57",X"00",X"57",X"00",X"58",X"00",X"57",X"00",X"58",X"00",X"58",X"00",X"57",X"00",X"58",X"00",
		X"56",X"00",X"58",X"00",X"55",X"00",X"57",X"00",X"56",X"00",X"56",X"00",X"56",X"00",X"56",X"00",
		X"56",X"00",X"55",X"00",X"55",X"00",X"56",X"00",X"57",X"00",X"56",X"00",X"57",X"00",X"55",X"00",
		X"56",X"00",X"56",X"00",X"55",X"00",X"56",X"00",X"56",X"00",X"56",X"00",X"56",X"00",X"57",X"00",
		X"56",X"00",X"56",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",
		X"56",X"00",X"56",X"00",X"53",X"00",X"56",X"00",X"54",X"00",X"54",X"00",X"56",X"00",X"56",X"00",
		X"54",X"00",X"55",X"00",X"56",X"00",X"55",X"00",X"54",X"00",X"55",X"00",X"55",X"00",X"55",X"00",
		X"55",X"00",X"55",X"00",X"56",X"00",X"54",X"00",X"54",X"00",X"54",X"00",X"54",X"00",X"54",X"00",
		X"54",X"00",X"55",X"00",X"55",X"00",X"54",X"00",X"54",X"00",X"53",X"00",X"54",X"00",X"54",X"00",
		X"55",X"00",X"54",X"00",X"54",X"00",X"54",X"00",X"53",X"00",X"54",X"00",X"55",X"00",X"54",X"00",
		X"54",X"00",X"55",X"00",X"55",X"00",X"54",X"00",X"53",X"00",X"53",X"00",X"53",X"00",X"53",X"00",
		X"52",X"00",X"53",X"00",X"53",X"00",X"52",X"00",X"52",X"00",X"53",X"00",X"54",X"00",X"53",X"00",
		X"53",X"00",X"53",X"00",X"54",X"00",X"53",X"00",X"53",X"00",X"53",X"00",X"53",X"00",X"53",X"00",
		X"52",X"00",X"53",X"00",X"52",X"00",X"53",X"00",X"53",X"00",X"54",X"00",X"52",X"00",X"53",X"00",
		X"52",X"00",X"52",X"00",X"53",X"00",X"53",X"00",X"52",X"00",X"52",X"00",X"52",X"00",X"52",X"00",
		X"52",X"00",X"51",X"00",X"53",X"00",X"52",X"00",X"52",X"00",X"53",X"00",X"51",X"00",X"51",X"00",
		X"52",X"00",X"51",X"00",X"52",X"00",X"52",X"00",X"52",X"00",X"52",X"00",X"51",X"00",X"51",X"00",
		X"52",X"00",X"52",X"00",X"52",X"00",X"52",X"00",X"51",X"00",X"51",X"00",X"52",X"00",X"50",X"00",
		X"51",X"00",X"51",X"00",X"50",X"00",X"51",X"00",X"51",X"00",X"52",X"00",X"51",X"00",X"50",X"00",
		X"50",X"00",X"51",X"00",X"50",X"00",X"50",X"00",X"52",X"00",X"50",X"00",X"50",X"00",X"50",X"00",
		X"51",X"00",X"52",X"00",X"51",X"00",X"52",X"00",X"51",X"00",X"50",X"00",X"51",X"00",X"51",X"00",
		X"50",X"00",X"4F",X"00",X"4F",X"00",X"51",X"00",X"4F",X"00",X"50",X"00",X"51",X"00",X"50",X"00",
		X"50",X"00",X"50",X"00",X"4F",X"00",X"50",X"00",X"4F",X"00",X"4F",X"00",X"4F",X"00",X"50",X"00",
		X"51",X"00",X"50",X"00",X"51",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"51",X"00",
		X"50",X"00",X"4E",X"00",X"4E",X"00",X"4E",X"00",X"4F",X"00",X"4F",X"00",X"4E",X"00",X"4E",X"00",
		X"4F",X"00",X"4F",X"00",X"4F",X"00",X"50",X"00",X"4F",X"00",X"4F",X"00",X"4F",X"00",X"50",X"00",
		X"50",X"00",X"50",X"00",X"4E",X"00",X"51",X"00",X"4E",X"00",X"4E",X"00",X"4E",X"00",X"4F",X"00",
		X"50",X"00",X"50",X"00",X"50",X"00",X"4F",X"00",X"4E",X"00",X"4F",X"00",X"4E",X"00",X"4E",X"00",
		X"4F",X"00",X"4E",X"00",X"4E",X"00",X"4E",X"00",X"4E",X"00",X"4E",X"00",X"4E",X"00",X"4E",X"00",
		X"4E",X"00",X"4E",X"00",X"4F",X"00",X"4F",X"00",X"50",X"00",X"4F",X"00",X"4D",X"00",X"4E",X"00",
		X"4E",X"00",X"4F",X"00",X"4D",X"00",X"4D",X"00",X"4F",X"00",X"4D",X"00",X"4E",X"00",X"4E",X"00",
		X"4E",X"00",X"4D",X"00",X"4D",X"00",X"4D",X"00",X"4D",X"00",X"4E",X"00",X"4D",X"00",X"4D",X"00",
		X"4C",X"00",X"4D",X"00",X"4C",X"00",X"4C",X"00",X"4E",X"00",X"4D",X"00",X"4D",X"00",X"4D",X"00",
		X"4D",X"00",X"4E",X"00",X"4D",X"00",X"4D",X"00",X"4D",X"00",X"4D",X"00",X"4D",X"00",X"4C",X"00",
		X"4D",X"00",X"4D",X"00",X"4F",X"00",X"4D",X"00",X"4D",X"00",X"4D",X"00",X"4C",X"00",X"4C",X"00",
		X"4B",X"00",X"4B",X"00",X"4B",X"00",X"4C",X"00",X"4B",X"00",X"4C",X"00",X"4C",X"00",X"4D",X"00",
		X"4C",X"00",X"4D",X"00",X"4D",X"00",X"4D",X"00",X"4C",X"00",X"4D",X"00",X"4C",X"00",X"4C",X"00",
		X"4C",X"00",X"4C",X"00",X"4C",X"00",X"4B",X"00",X"4B",X"00",X"4C",X"00",X"4B",X"00",X"4C",X"00",
		X"4B",X"00",X"4D",X"00",X"4B",X"00",X"4C",X"00",X"4B",X"00",X"4A",X"00",X"4B",X"00",X"4C",X"00",
		X"4B",X"00",X"4B",X"00",X"4B",X"00",X"4B",X"00",X"4B",X"00",X"4B",X"00",X"4A",X"00",X"4A",X"00",
		X"4C",X"00",X"4A",X"00",X"4B",X"00",X"4A",X"00",X"4B",X"00",X"4A",X"00",X"4C",X"00",X"4B",X"00",
		X"4D",X"00",X"4A",X"00",X"4C",X"00",X"4C",X"00",X"4A",X"00",X"4B",X"00",X"4C",X"00",X"49",X"00",
		X"4A",X"00",X"4A",X"00",X"4A",X"00",X"49",X"00",X"4A",X"00",X"4B",X"00",X"4B",X"00",X"4A",X"00",
		X"4B",X"00",X"4B",X"00",X"4A",X"00",X"4A",X"00",X"49",X"00",X"4B",X"00",X"4A",X"00",X"4A",X"00",
		X"49",X"00",X"49",X"00",X"4A",X"00",X"4B",X"00",X"4A",X"00",X"4A",X"00",X"4A",X"00",X"4B",X"00",
		X"4A",X"00",X"4A",X"00",X"4B",X"00",X"B0",X"B0",X"E9",X"FF",X"BD",X"FE",X"DA",X"FB",X"14",X"FA",
		X"9A",X"F8",X"63",X"F5",X"DE",X"F4",X"D2",X"F3",X"85",X"F2",X"7E",X"EF",X"23",X"EE",X"4E",X"ED",
		X"5A",X"EB",X"D2",X"E9",X"F7",X"E7",X"E8",X"E4",X"3D",X"E3",X"7C",X"E1",X"63",X"E0",X"95",X"E0",
		X"7A",X"E0",X"2D",X"E0",X"A3",X"E2",X"9C",X"E2",X"0B",X"E3",X"C3",X"E3",X"B1",X"E5",X"46",X"E6",
		X"33",X"E7",X"1A",X"E9",X"61",X"E9",X"7E",X"EA",X"AF",X"E9",X"58",X"EC",X"30",X"EC",X"38",X"EC",
		X"9E",X"EC",X"AE",X"EE",X"2F",X"EF",X"14",X"EF",X"22",X"F0",X"C1",X"F0",X"A8",X"F1",X"40",X"F2",
		X"12",X"F4",X"9F",X"F5",X"0E",X"F6",X"04",X"F7",X"2C",X"F6",X"F7",X"F6",X"C0",X"F7",X"4E",X"FA",
		X"C6",X"F9",X"A4",X"FA",X"71",X"FB",X"4D",X"FC",X"CD",X"FE",X"82",X"FE",X"41",X"01",X"15",X"02",
		X"F0",X"03",X"40",X"06",X"DA",X"09",X"1F",X"0C",X"33",X"0E",X"F5",X"11",X"B9",X"14",X"3D",X"19",
		X"7C",X"1D",X"87",X"1F",X"2D",X"17",X"67",X"0D",X"7E",X"03",X"CF",X"F7",X"4D",X"ED",X"52",X"E2",
		X"21",X"E5",X"B1",X"EA",X"B9",X"F1",X"32",X"F7",X"D8",X"FC",X"3D",X"05",X"D6",X"0A",X"69",X"13",
		X"83",X"1A",X"C3",X"1D",X"43",X"0E",X"BF",X"FD",X"91",X"EB",X"D9",X"E2",X"1E",X"EB",X"39",X"F4",
		X"35",X"FE",X"93",X"08",X"B9",X"10",X"2D",X"1B",X"B2",X"18",X"F6",X"02",X"37",X"EE",X"C4",X"E2",
		X"54",X"EF",X"C6",X"F6",X"8D",X"02",X"3E",X"0C",X"FD",X"15",X"DC",X"1C",X"A0",X"0C",X"C1",X"F6",
		X"6C",X"E5",X"A0",X"E9",X"48",X"F5",X"CE",X"FC",X"9B",X"09",X"83",X"11",X"A2",X"1C",X"F1",X"16",
		X"51",X"01",X"47",X"EB",X"D6",X"E4",X"00",X"F1",X"B3",X"F9",X"C5",X"04",X"DC",X"0D",X"3A",X"18",
		X"13",X"1C",X"29",X"0A",X"62",X"F3",X"76",X"E4",X"2D",X"EB",X"8B",X"F5",X"33",X"FE",X"B6",X"09",
		X"51",X"11",X"EF",X"1C",X"58",X"14",X"89",X"FF",X"7C",X"E8",X"51",X"E5",X"7C",X"F1",X"46",X"FA",
		X"56",X"04",X"70",X"0D",X"E5",X"19",X"56",X"1C",X"5B",X"09",X"6F",X"F4",X"0C",X"E4",X"BA",X"E9",
		X"77",X"F4",X"86",X"FE",X"8A",X"09",X"29",X"11",X"48",X"1D",X"45",X"16",X"37",X"FF",X"BD",X"E9",
		X"BF",X"E4",X"6E",X"EF",X"98",X"F8",X"39",X"03",X"A3",X"0D",X"E9",X"18",X"7C",X"1D",X"5D",X"0A",
		X"D5",X"F4",X"E3",X"E3",X"8A",X"E9",X"BF",X"F4",X"9A",X"FD",X"BC",X"08",X"12",X"10",X"A7",X"1C",
		X"CA",X"15",X"DE",X"01",X"45",X"EB",X"4E",X"E2",X"DF",X"EF",X"9D",X"F8",X"43",X"02",X"1C",X"0B",
		X"EC",X"15",X"5A",X"1D",X"84",X"0F",X"F1",X"F7",X"23",X"E5",X"55",X"E7",X"7D",X"F3",X"D6",X"FC",
		X"33",X"07",X"94",X"0E",X"D7",X"1A",X"76",X"1A",X"4A",X"05",X"BB",X"EF",X"B2",X"E2",X"E1",X"EB",
		X"2E",X"F7",X"37",X"FF",X"5B",X"0A",X"BD",X"13",X"AA",X"1D",X"93",X"12",X"55",X"FD",X"78",X"E8",
		X"CC",X"E3",X"AF",X"F0",X"70",X"F8",X"14",X"04",X"13",X"0C",X"F0",X"18",X"03",X"1D",X"E4",X"0A",
		X"E6",X"F5",X"B2",X"E3",X"99",X"E9",X"8C",X"F4",X"73",X"FC",X"76",X"08",X"CB",X"0E",X"FF",X"1C",
		X"BF",X"18",X"88",X"04",X"FE",X"ED",X"3C",X"E2",X"E8",X"ED",X"51",X"F7",X"49",X"01",X"1F",X"0A",
		X"1E",X"14",X"F4",X"1E",X"5A",X"12",X"FB",X"FC",X"6B",X"E7",X"7E",X"E4",X"E0",X"F0",X"F5",X"F8",
		X"1E",X"04",X"87",X"0C",X"C3",X"18",X"89",X"1C",X"A6",X"0C",X"7B",X"F7",X"E0",X"E3",X"DE",X"E7",
		X"53",X"F4",X"34",X"FC",X"96",X"07",X"44",X"0E",X"E5",X"1B",X"99",X"1A",X"3B",X"07",X"F9",X"F1",
		X"1E",X"E4",X"D1",X"EA",X"87",X"F5",X"57",X"FF",X"94",X"09",X"0E",X"11",X"3C",X"1C",X"83",X"16",
		X"27",X"01",X"FC",X"EB",X"C9",X"E3",X"B5",X"ED",X"AD",X"F7",X"BC",X"01",X"CC",X"09",X"3D",X"14",
		X"71",X"1E",X"F6",X"12",X"E5",X"FD",X"4C",X"E9",X"FC",X"E3",X"EE",X"EF",X"38",X"F9",X"68",X"04",
		X"88",X"0C",X"8B",X"16",X"54",X"1E",X"38",X"0F",X"66",X"F8",X"EF",X"E4",X"29",X"E6",X"C8",X"F2",
		X"81",X"F9",X"82",X"05",X"84",X"0E",X"F1",X"18",X"A9",X"1B",X"72",X"0A",X"54",X"F4",X"F1",X"E3",
		X"C2",X"E8",X"64",X"F3",X"DC",X"FC",X"35",X"07",X"C3",X"0E",X"DB",X"1B",X"11",X"1A",X"68",X"07",
		X"55",X"F2",X"DE",X"E1",X"85",X"EA",X"C5",X"F4",X"96",X"FD",X"49",X"08",X"66",X"0F",X"CA",X"1C",
		X"86",X"19",X"BE",X"05",X"E6",X"EF",X"1E",X"E4",X"CB",X"EB",X"95",X"F5",X"A4",X"FF",X"8C",X"09",
		X"1B",X"11",X"A3",X"1D",X"51",X"16",X"D8",X"02",X"DA",X"ED",X"99",X"E3",X"CF",X"EC",X"97",X"F6",
		X"9B",X"FF",X"F8",X"08",X"2C",X"12",X"D4",X"1D",X"4E",X"15",X"AC",X"00",X"E0",X"EC",X"B8",X"E3",
		X"D2",X"EE",X"72",X"F6",X"67",X"00",X"9A",X"0A",X"66",X"12",X"19",X"1D",X"00",X"14",X"49",X"FF",
		X"3D",X"EA",X"0D",X"E3",X"D7",X"ED",X"CC",X"F7",X"44",X"00",X"69",X"0A",X"61",X"14",X"28",X"1E",
		X"15",X"14",X"7E",X"FF",X"0E",X"E9",X"27",X"E4",X"B8",X"EE",X"60",X"F7",X"61",X"01",X"DC",X"09",
		X"23",X"14",X"C2",X"1D",X"84",X"14",X"B9",X"FF",X"BB",X"E9",X"56",X"E4",X"D3",X"EE",X"25",X"F7",
		X"EC",X"01",X"47",X"0B",X"49",X"14",X"61",X"1E",X"F6",X"14",X"1A",X"FF",X"24",X"EB",X"6F",X"E4",
		X"02",X"EE",X"5A",X"F7",X"8E",X"01",X"EE",X"09",X"C6",X"13",X"06",X"1E",X"8A",X"14",X"33",X"01",
		X"BF",X"EB",X"A2",X"E2",X"CE",X"ED",X"CB",X"F6",X"4B",X"FF",X"85",X"09",X"BA",X"12",X"11",X"1D",
		X"3D",X"15",X"21",X"02",X"81",X"ED",X"E8",X"E3",X"5C",X"ED",X"DB",X"F6",X"B1",X"FF",X"A4",X"08",
		X"3A",X"11",X"A4",X"1D",X"B3",X"17",X"0B",X"03",X"1A",X"EE",X"4F",X"E3",X"79",X"EB",X"75",X"F4",
		X"D6",X"FD",X"A7",X"08",X"F1",X"0F",X"F3",X"1B",X"66",X"1A",X"7C",X"06",X"EA",X"F0",X"96",X"E2",
		X"C6",X"EA",X"47",X"F3",X"9F",X"FC",X"1B",X"06",X"97",X"0F",X"E0",X"1A",X"63",X"1B",X"0D",X"08",
		X"1A",X"F4",X"0F",X"E3",X"3D",X"E9",X"44",X"F3",X"54",X"FC",X"D5",X"05",X"F3",X"0D",X"6D",X"18",
		X"F0",X"1C",X"E0",X"0C",X"8B",X"F8",X"BC",X"E4",X"90",X"E7",X"DD",X"F0",X"29",X"FA",X"53",X"03",
		X"E2",X"0C",X"BC",X"16",X"93",X"1E",X"30",X"10",X"66",X"FC",X"8E",X"E7",X"81",X"E4",X"C9",X"EE",
		X"51",X"F7",X"1F",X"01",X"86",X"0B",X"2B",X"14",X"B6",X"1E",X"59",X"15",X"5D",X"FF",X"80",X"EC",
		X"71",X"E2",X"BB",X"EC",X"01",X"F6",X"28",X"FF",X"C1",X"07",X"47",X"11",X"63",X"1C",X"CA",X"19",
		X"1B",X"04",X"48",X"F1",X"DB",X"E2",X"FD",X"E9",X"1E",X"F3",X"7E",X"FD",X"7C",X"05",X"89",X"10",
		X"37",X"18",X"80",X"1D",X"E2",X"0A",X"35",X"F8",X"4F",X"E4",X"DB",X"E6",X"49",X"F0",X"40",X"FA",
		X"C1",X"03",X"B9",X"0D",X"58",X"15",X"24",X"1E",X"1B",X"10",X"25",X"FD",X"C0",X"E8",X"11",X"E4",
		X"A1",X"EE",X"2A",X"F7",X"9E",X"00",X"E3",X"09",X"74",X"12",X"E9",X"1B",X"4D",X"18",X"23",X"02",
		X"95",X"EF",X"9A",X"E2",X"47",X"EC",X"C2",X"F3",X"2F",X"FD",X"B1",X"05",X"A4",X"0F",X"81",X"19",
		X"55",X"1C",X"F4",X"09",X"2B",X"F7",X"43",X"E3",X"04",X"E7",X"28",X"F0",X"D8",X"F9",X"37",X"02",
		X"75",X"0C",X"90",X"15",X"F6",X"1E",X"2F",X"12",X"98",X"FD",X"2D",X"EA",X"D0",X"E2",X"2C",X"EE",
		X"DD",X"F5",X"8B",X"FF",X"9D",X"09",X"3B",X"11",X"D6",X"1B",X"C1",X"19",X"DD",X"05",X"9C",X"F3",
		X"CE",X"E1",X"93",X"E9",X"6F",X"F2",X"0A",X"FC",X"95",X"04",X"1D",X"0E",X"7D",X"17",X"3A",X"1F",
		X"17",X"0F",X"36",X"FC",X"B6",X"E6",X"E8",X"E4",X"C5",X"EE",X"B2",X"F7",X"93",X"00",X"34",X"0A",
		X"18",X"13",X"01",X"1C",X"FB",X"17",X"FF",X"02",X"B7",X"F0",X"87",X"E2",X"4A",X"EB",X"6A",X"F3",
		X"80",X"FD",X"B3",X"04",X"22",X"0F",X"ED",X"16",X"A2",X"1E",X"4C",X"0D",X"54",X"FA",X"BE",X"E5",
		X"16",X"E5",X"BA",X"EF",X"25",X"F7",X"51",X"00",X"7E",X"09",X"DF",X"11",X"78",X"1C",X"E1",X"18",
		X"9C",X"04",X"F5",X"F0",X"1C",X"E2",X"F2",X"EA",X"3E",X"F2",X"D5",X"FC",X"38",X"04",X"1E",X"0F",
		X"3D",X"16",X"B5",X"1E",X"2F",X"0F",X"0E",X"FC",X"FC",X"E7",X"D6",X"E3",X"92",X"EE",X"A5",X"F6",
		X"39",X"00",X"31",X"08",X"32",X"11",X"9C",X"1B",X"F4",X"1A",X"AD",X"06",X"AC",X"F3",X"0F",X"E3",
		X"E1",X"E8",X"E9",X"F0",X"69",X"FA",X"BA",X"02",X"74",X"0C",X"B6",X"15",X"3F",X"1E",X"B2",X"12",
		X"98",X"FF",X"47",X"EB",X"FB",X"E2",X"3E",X"ED",X"79",X"F4",X"9B",X"FE",X"55",X"07",X"5C",X"0F",
		X"69",X"18",X"ED",X"1C",X"C1",X"0B",X"4C",X"F9",X"E6",X"E4",X"1F",X"E6",X"30",X"F0",X"69",X"F8",
		X"6D",X"00",X"C9",X"09",X"D2",X"11",X"4F",X"1C",X"70",X"18",X"D1",X"04",X"CD",X"F2",X"0B",X"E2",
		X"E6",X"E8",X"66",X"F1",X"E8",X"FA",X"0A",X"03",X"14",X"0D",X"E9",X"15",X"D8",X"1E",X"08",X"13",
		X"94",X"FE",X"EC",X"EB",X"0A",X"E3",X"20",X"ED",X"20",X"F4",X"3D",X"FE",X"F7",X"05",X"DB",X"0F",
		X"95",X"18",X"63",X"1D",X"E8",X"0C",X"8A",X"FA",X"9C",X"E6",X"42",X"E4",X"E9",X"EE",X"24",X"F6",
		X"D2",X"FF",X"6E",X"09",X"54",X"11",X"02",X"1B",X"F5",X"1B",X"E1",X"06",X"6A",X"F6",X"46",X"E4",
		X"E0",X"E6",X"BF",X"EF",X"E9",X"F9",X"FB",X"01",X"78",X"0A",X"D0",X"12",X"AA",X"1D",X"06",X"18",
		X"A9",X"04",X"EE",X"F1",X"93",X"E2",X"5F",X"E9",X"C9",X"F1",X"DD",X"FB",X"2F",X"03",X"33",X"0C",
		X"32",X"14",X"C1",X"1E",X"40",X"14",X"DD",X"00",X"9A",X"ED",X"92",X"E1",X"4C",X"EB",X"3A",X"F3",
		X"AE",X"FC",X"62",X"05",X"A7",X"0E",X"B6",X"16",X"E3",X"1E",X"DC",X"10",X"52",X"FE",X"46",X"EB",
		X"23",X"E3",X"56",X"EC",X"DF",X"F3",X"6E",X"FD",X"96",X"06",X"56",X"0F",X"77",X"17",X"4E",X"1E",
		X"B5",X"0D",X"CB",X"FB",X"A7",X"E8",X"35",X"E3",X"AB",X"ED",X"48",X"F5",X"00",X"FF",X"15",X"07",
		X"B4",X"0F",X"8E",X"19",X"89",X"1D",X"F9",X"0C",X"01",X"FB",X"05",X"E7",X"A3",X"E4",X"A5",X"EE",
		X"AA",X"F6",X"69",X"FF",X"E8",X"06",X"A7",X"10",X"23",X"19",X"62",X"1D",X"EC",X"0B",X"2E",X"F9",
		X"19",X"E6",X"2C",X"E5",X"F5",X"EE",X"58",X"F6",X"C0",X"FF",X"C5",X"07",X"EE",X"0F",X"8D",X"19",
		X"EE",X"1C",X"53",X"0A",X"B3",X"F8",X"1D",X"E6",X"73",X"E5",X"F9",X"EE",X"3F",X"F7",X"41",X"FF",
		X"6A",X"08",X"23",X"10",X"5D",X"19",X"40",X"1D",X"70",X"0B",X"DE",X"F9",X"D6",X"E5",X"2B",X"E4",
		X"1B",X"EE",X"20",X"F7",X"72",X"FF",X"A6",X"07",X"15",X"11",X"1B",X"19",X"8B",X"1C",X"45",X"0B",
		X"B9",X"F9",X"47",X"E7",X"F2",X"E3",X"83",X"EE",X"6C",X"F6",X"7C",X"FF",X"9F",X"07",X"A5",X"0F",
		X"E5",X"18",X"26",X"1D",X"F8",X"0C",X"17",X"FC",X"48",X"E8",X"0F",X"E3",X"D9",X"EC",X"51",X"F5",
		X"DA",X"FE",X"B3",X"06",X"FC",X"0E",X"C6",X"17",X"12",X"1E",X"DE",X"0E",X"D3",X"FC",X"CD",X"E9",
		X"41",X"E2",X"E3",X"EB",X"C1",X"F3",X"EB",X"FD",X"38",X"05",X"C6",X"0D",X"AA",X"15",X"15",X"1E",
		X"88",X"11",X"07",X"00",X"9B",X"EC",X"14",X"E2",X"8E",X"EA",X"8F",X"F2",X"26",X"FC",X"98",X"03",
		X"32",X"0D",X"EA",X"13",X"7A",X"1D",X"09",X"15",X"4A",X"03",X"7F",X"F0",X"ED",X"E1",X"7D",X"E8",
		X"94",X"F1",X"1A",X"FA",X"AD",X"01",X"98",X"0B",X"8A",X"12",X"26",X"1D",X"BA",X"19",X"72",X"05",
		X"75",X"F4",X"69",X"E3",X"4F",X"E7",X"1C",X"F0",X"B7",X"F8",X"96",X"00",X"EA",X"08",X"CD",X"11",
		X"3D",X"1A",X"4E",X"1C",X"80",X"0A",X"C5",X"F8",X"EA",X"E6",X"6E",X"E4",X"B2",X"ED",X"F4",X"F4",
		X"A1",X"FE",X"8F",X"06",X"43",X"0F",X"EB",X"17",X"EF",X"1E",X"69",X"10",X"BA",X"FE",X"69",X"EB",
		X"4B",X"E2",X"7A",X"EB",X"18",X"F3",X"CF",X"FC",X"47",X"04",X"B7",X"0C",X"0C",X"14",X"34",X"1E",
		X"4A",X"16",X"B9",X"02",X"98",X"F1",X"D6",X"E2",X"81",X"E7",X"E2",X"F0",X"AA",X"F9",X"C3",X"01",
		X"7E",X"0A",X"DC",X"11",X"A4",X"1A",X"4B",X"1B",X"A4",X"08",X"E5",X"F8",X"47",X"E5",X"DE",X"E4",
		X"68",X"EE",X"83",X"F5",X"1E",X"FF",X"F0",X"06",X"A2",X"0F",X"AC",X"17",X"9D",X"1E",X"57",X"10",
		X"88",X"FE",X"C6",X"EC",X"4F",X"E2",X"C2",X"EA",X"CA",X"F1",X"A4",X"FB",X"6E",X"03",X"CC",X"0B",
		X"93",X"13",X"BA",X"1C",X"32",X"18",X"B5",X"05",X"0A",X"F5",X"92",X"E3",X"45",X"E6",X"BC",X"EE",
		X"85",X"F7",X"3F",X"00",X"9C",X"07",X"C2",X"0F",X"3A",X"18",X"58",X"1D",X"E7",X"0D",X"99",X"FC",
		X"B9",X"EA",X"1B",X"E2",X"22",X"EB",X"F4",X"F2",X"82",X"FC",X"2A",X"04",X"AB",X"0C",X"71",X"13",
		X"FF",X"1C",X"54",X"17",X"2D",X"05",X"EF",X"F3",X"DA",X"E2",X"0E",X"E6",X"37",X"EF",X"EE",X"F7",
		X"34",X"00",X"B8",X"07",X"A8",X"0F",X"3D",X"18",X"7C",X"1D",X"B6",X"0E",X"A0",X"FD",X"89",X"EA",
		X"96",X"E1",X"E4",X"EA",X"37",X"F2",X"3C",X"FB",X"A5",X"02",X"B0",X"0B",X"D7",X"12",X"93",X"1D",
		X"AE",X"19",X"25",X"06",X"D0",X"F5",X"E9",X"E3",X"A4",X"E5",X"15",X"EF",X"62",X"F6",X"51",X"FE",
		X"97",X"06",X"9C",X"0F",X"51",X"17",X"3A",X"1E",X"80",X"11",X"CC",X"00",X"CE",X"EE",X"1D",X"E2",
		X"57",X"E9",X"14",X"F1",X"0F",X"FA",X"FA",X"01",X"38",X"0A",X"70",X"11",X"E8",X"1A",X"D6",X"1C",
		X"32",X"0B",X"AB",X"FA",X"45",X"E8",X"EA",X"E2",X"0D",X"ED",X"FF",X"F3",X"70",X"FC",X"70",X"03",
		X"BA",X"0C",X"1D",X"14",X"69",X"1D",X"CA",X"18",X"8D",X"05",X"AF",X"F4",X"B8",X"E3",X"DC",X"E5",
		X"7C",X"EE",X"E5",X"F6",X"D2",X"FE",X"0B",X"06",X"20",X"0F",X"95",X"16",X"3A",X"1E",X"EE",X"12",
		X"99",X"00",X"B8",X"EF",X"AA",X"E1",X"44",X"E8",X"AE",X"F0",X"2D",X"F8",X"B6",X"00",X"E6",X"08",
		X"08",X"10",X"37",X"19",X"D1",X"1D",X"3B",X"0E",X"1F",X"FE",X"4B",X"EB",X"E4",X"E1",X"2C",X"EA",
		X"62",X"F2",X"00",X"FB",X"CF",X"01",X"7B",X"0A",X"8F",X"12",X"71",X"1B",X"AB",X"1C",X"6C",X"0A",
		X"9B",X"FA",X"CE",X"E7",X"EE",X"E2",X"81",X"EC",X"25",X"F3",X"DB",X"FC",X"30",X"03",X"65",X"0C",
		X"B0",X"13",X"4E",X"1C",X"05",X"1A",X"91",X"07",X"54",X"F7",X"B1",X"E5",X"05",X"E4",X"E9",X"EC",
		X"A2",X"F4",X"3D",X"FD",X"14",X"04",X"E3",X"0C",X"92",X"14",X"7C",X"1D",X"66",X"17",X"1F",X"06",
		X"21",X"F6",X"01",X"E5",X"27",X"E5",X"F1",X"ED",X"B9",X"F5",X"2D",X"FE",X"16",X"05",X"2C",X"0E",
		X"65",X"14",X"FE",X"1D",X"88",X"16",X"CF",X"04",X"E5",X"F4",X"AB",X"E3",X"B4",X"E5",X"10",X"EF",
		X"BE",X"F5",X"ED",X"FD",X"FA",X"05",X"93",X"0E",X"29",X"15",X"2F",X"1E",X"97",X"15",X"1D",X"04",
		X"10",X"F4",X"28",X"E3",X"44",X"E5",X"D0",X"EE",X"F5",X"F5",X"EF",X"FD",X"28",X"06",X"8C",X"0E",
		X"CE",X"15",X"5A",X"1D",X"84",X"16",X"09",X"04",X"7F",X"F4",X"0B",X"E3",X"2F",X"E5",X"E9",X"EE",
		X"28",X"F6",X"4A",X"FE",X"1C",X"05",X"97",X"0D",X"1C",X"15",X"3E",X"1E",X"8E",X"17",X"67",X"05",
		X"A4",X"F5",X"72",X"E4",X"DD",X"E4",X"31",X"EE",X"CD",X"F4",X"E3",X"FD",X"52",X"05",X"88",X"0D",
		X"23",X"14",X"D5",X"1D",X"0A",X"19",X"DF",X"06",X"6C",X"F7",X"78",X"E5",X"C8",X"E3",X"C7",X"EC",
		X"07",X"F4",X"40",X"FC",X"D9",X"03",X"72",X"0C",X"46",X"13",X"A5",X"1C",X"CB",X"1A",X"3A",X"09",
		X"DB",X"F9",X"6B",X"E7",X"54",X"E2",X"CE",X"EB",X"95",X"F2",X"93",X"FB",X"AF",X"02",X"94",X"0A",
		X"D6",X"11",X"98",X"1A",X"35",X"1D",X"47",X"0C",X"25",X"FC",X"09",X"EB",X"72",X"E2",X"C5",X"E9",
		X"7C",X"F1",X"F9",X"F9",X"B6",X"01",X"45",X"09",X"64",X"10",X"63",X"18",X"DB",X"1D",X"DA",X"10",
		X"88",X"FF",X"81",X"EE",X"3E",X"E2",X"DC",X"E7",X"3A",X"F0",X"06",X"F8",X"CB",X"FF",X"39",X"07",
		X"7C",X"0E",X"29",X"16",X"92",X"1D",X"46",X"15",X"D3",X"03",X"B8",X"F3",X"7C",X"E3",X"97",X"E5",
		X"60",X"EE",X"12",X"F5",X"70",X"FD",X"10",X"05",X"62",X"0C",X"A4",X"13",X"C5",X"1C",X"4C",X"1A",
		X"E3",X"08",X"28",X"F9",X"EA",X"E7",X"21",X"E3",X"DA",X"EB",X"AF",X"F2",X"9C",X"FA",X"33",X"02",
		X"82",X"09",X"73",X"11",X"E2",X"19",X"D3",X"1D",X"F1",X"0E",X"C5",X"FE",X"0A",X"EE",X"83",X"E2",
		X"37",X"E8",X"89",X"EF",X"92",X"F7",X"58",X"FF",X"5B",X"06",X"60",X"0E",X"E8",X"15",X"9A",X"1E",
		X"E0",X"16",X"EB",X"04",X"67",X"F6",X"22",X"E5",X"A7",X"E4",X"B2",X"EC",X"5B",X"F4",X"B6",X"FB",
		X"43",X"03",X"78",X"0B",X"0D",X"12",X"A9",X"1A",X"70",X"1C",X"C0",X"0C",X"A0",X"FD",X"42",X"EC",
		X"AA",X"E1",X"53",X"E9",X"A9",X"F0",X"E0",X"F7",X"A8",X"FF",X"09",X"07",X"D6",X"0E",X"0D",X"16",
		X"CA",X"1D",X"1C",X"16",X"18",X"04",X"20",X"F5",X"11",X"E4",X"03",X"E4",X"20",X"ED",X"77",X"F4",
		X"DC",X"FB",X"6B",X"03",X"FF",X"0A",X"74",X"12",X"E4",X"1A",X"C6",X"1C",X"EC",X"0D",X"DF",X"FD",
		X"77",X"ED",X"CC",X"E1",X"3C",X"E8",X"0F",X"F0",X"73",X"F7",X"2C",X"FF",X"74",X"06",X"4D",X"0E",
		X"D6",X"14",X"79",X"1D",X"2A",X"18",X"74",X"06",X"6A",X"F8",X"35",X"E6",X"2A",X"E3",X"86",X"EB",
		X"D3",X"F2",X"D2",X"FA",X"70",X"01",X"32",X"09",X"60",X"10",X"61",X"18",X"5D",X"1E",X"46",X"12",
		X"40",X"01",X"CC",X"F1",X"4B",X"E3",X"39",X"E6",X"36",X"EE",X"0B",X"F5",X"37",X"FD",X"53",X"04",
		X"83",X"0B",X"AA",X"12",X"E3",X"1A",X"EA",X"1C",X"AE",X"0C",X"6F",X"FD",X"DD",X"EC",X"16",X"E2",
		X"BD",X"E8",X"E9",X"EF",X"04",X"F7",X"B3",X"FE",X"DF",X"05",X"29",X"0E",X"07",X"15",X"82",X"1D",
		X"99",X"19",X"22",X"08",X"40",X"FA",X"1D",X"E8",X"FE",X"E1",X"52",X"EA",X"B5",X"F1",X"F4",X"F8",
		X"FE",X"00",X"B2",X"07",X"82",X"0F",X"5F",X"16",X"2D",X"1E",X"85",X"16",X"4C",X"05",X"85",X"F6",
		X"94",X"E5",X"BE",X"E3",X"31",X"EC",X"DD",X"F2",X"32",X"FA",X"69",X"01",X"17",X"09",X"8E",X"10",
		X"C8",X"17",X"57",X"1E",X"E0",X"13",X"75",X"03",X"79",X"F4",X"89",X"E4",X"9F",X"E4",X"38",X"ED",
		X"E0",X"F3",X"36",X"FB",X"38",X"02",X"01",X"0A",X"8B",X"11",X"BD",X"18",X"44",X"1E",X"76",X"12",
		X"4E",X"01",X"BF",X"F2",X"83",X"E3",X"0F",X"E5",X"62",X"ED",X"B5",X"F4",X"B1",X"FB",X"D4",X"02",
		X"B1",X"0A",X"F0",X"11",X"58",X"19",X"34",X"1E",X"50",X"11",X"2B",X"01",X"16",X"F2",X"8F",X"E2",
		X"8B",X"E5",X"D8",X"ED",X"8E",X"F4",X"AD",X"FB",X"37",X"03",X"89",X"0A",X"A2",X"11",X"43",X"19",
		X"E3",X"1D",X"57",X"11",X"90",X"01",X"92",X"F2",X"A7",X"E3",X"88",X"E5",X"89",X"ED",X"8E",X"F4",
		X"AE",X"FB",X"88",X"02",X"5C",X"0A",X"9B",X"11",X"C7",X"18",X"D8",X"1D",X"B0",X"12",X"8B",X"02",
		X"6A",X"F3",X"77",X"E3",X"91",X"E4",X"9F",X"EC",X"4E",X"F3",X"89",X"FB",X"08",X"02",X"93",X"09",
		X"80",X"10",X"F7",X"17",X"0E",X"1E",X"A1",X"14",X"43",X"04",X"66",X"F5",X"22",X"E5",X"B1",X"E3",
		X"08",X"EC",X"C9",X"F2",X"3E",X"FA",X"EC",X"00",X"7B",X"08",X"45",X"0F",X"5A",X"16",X"78",X"1E",
		X"DA",X"17",X"A2",X"06",X"9A",X"F8",X"45",X"E7",X"60",X"E2",X"5F",X"EA",X"85",X"F1",X"AE",X"F8",
		X"FA",X"FF",X"EC",X"06",X"07",X"0E",X"D7",X"14",X"BD",X"1C",X"CD",X"1A",X"6F",X"0A",X"06",X"FC",
		X"6C",X"EB",X"A4",X"E1",X"37",X"E8",X"D1",X"EF",X"7B",X"F6",X"92",X"FD",X"00",X"05",X"F2",X"0B",
		X"C2",X"12",X"D6",X"1A",X"F0",X"1C",X"DA",X"0E",X"B0",X"FF",X"D9",X"F0",X"4E",X"E2",X"97",X"E5",
		X"70",X"ED",X"7A",X"F4",X"E4",X"FB",X"88",X"02",X"7A",X"09",X"DD",X"10",X"D0",X"17",X"3D",X"1E",
		X"07",X"15",X"AB",X"04",X"E8",X"F6",X"D8",X"E5",X"23",X"E3",X"1E",X"EB",X"D9",X"F1",X"AB",X"F8",
		X"C0",X"FF",X"B1",X"06",X"FF",X"0D",X"91",X"14",X"92",X"1C",X"2C",X"1B",X"93",X"0A",X"CC",X"FC",
		X"72",X"EC",X"24",X"E2",X"4B",X"E7",X"94",X"EE",X"A8",X"F5",X"13",X"FD",X"82",X"03",X"E6",X"0A",
		X"7D",X"11",X"30",X"19",X"30",X"1E",X"6A",X"12",X"96",X"02",X"AB",X"F4",X"4F",X"E5",X"CA",X"E3",
		X"84",X"EB",X"4D",X"F2",X"C2",X"F9",X"8C",X"00",X"A7",X"07",X"A8",X"0E",X"69",X"15",X"F9",X"1C",
		X"D4",X"1A",X"8B",X"0A",X"8D",X"FC",X"C3",X"EC",X"09",X"E2",X"38",X"E7",X"B0",X"EE",X"63",X"F5",
		X"A8",X"FC",X"5F",X"03",X"98",X"0A",X"45",X"11",X"8E",X"18",X"3C",X"1E",X"70",X"14",X"3D",X"04",
		X"AF",X"F6",X"3F",X"E6",X"9B",X"E2",X"59",X"EA",X"59",X"F1",X"EB",X"F7",X"54",X"FF",X"02",X"06",
		X"04",X"0D",X"77",X"13",X"9F",X"1B",X"24",X"1D",X"6F",X"0E",X"8D",X"FF",X"1A",X"F1",X"33",X"E3",
		X"08",X"E5",X"E7",X"EC",X"59",X"F3",X"A8",X"FA",X"0A",X"01",X"81",X"08",X"6B",X"0F",X"27",X"16",
		X"45",X"1D",X"74",X"19",X"45",X"09",X"C8",X"FB",X"CD",X"EB",X"DC",X"E1",X"81",X"E7",X"B5",X"EE",
		X"2A",X"F5",X"8A",X"FC",X"C0",X"02",X"39",X"0A",X"C7",X"10",X"8F",X"17",X"25",X"1E",X"8B",X"16",
		X"40",X"06",X"DA",X"F8",X"4B",X"E8",X"55",X"E2",X"2F",X"E9",X"1E",X"F0",X"DA",X"F6",X"F2",X"FD",
		X"6E",X"04",X"57",X"0B",X"37",X"12",X"2C",X"19",X"1D",X"1E",X"B0",X"13",X"8C",X"03",X"54",X"F6",
		X"97",X"E6",X"13",X"E3",X"FC",X"E9",X"E0",X"F0",X"D5",X"F7",X"7F",X"FE",X"FC",X"04",X"76",X"0C",
		X"7D",X"12",X"64",X"1A",X"45",X"1E",X"1F",X"12",X"B2",X"02",X"39",X"F5",X"9C",X"E5",X"48",X"E3",
		X"94",X"EA",X"1C",X"F1",X"3C",X"F8",X"E0",X"FE",X"65",X"05",X"86",X"0C",X"C1",X"12",X"5B",X"1A",
		X"4C",X"1D",X"84",X"11",X"51",X"02",X"C9",X"F4",X"45",X"E5",X"2F",X"E3",X"9B",X"EA",X"1D",X"F1",
		X"36",X"F8",X"2F",X"FF",X"B0",X"05",X"6F",X"0C",X"B9",X"12",X"7A",X"1A",X"38",X"1E",X"00",X"12",
		X"8F",X"02",X"52",X"F5",X"A6",X"E5",X"9C",X"E2",X"5E",X"EA",X"0D",X"F1",X"C5",X"F7",X"39",X"FE",
		X"30",X"05",X"E4",X"0B",X"36",X"12",X"58",X"19",X"D5",X"1D",X"4C",X"13",X"4C",X"04",X"DB",X"F6",
		X"27",X"E7",X"75",X"E2",X"6F",X"E9",X"1F",X"F0",X"0A",X"F7",X"8C",X"FD",X"FE",X"03",X"E1",X"0A",
		X"89",X"11",X"2A",X"18",X"38",X"1E",X"B2",X"15",X"B9",X"06",X"1A",X"F9",X"E1",X"E9",X"E4",X"E1",
		X"FC",X"E7",X"79",X"EE",X"8B",X"F5",X"26",X"FC",X"CC",X"02",X"5F",X"09",X"12",X"10",X"37",X"16",
		X"8F",X"1D",X"09",X"19",X"F0",X"09",X"6E",X"FC",X"F8",X"ED",X"2A",X"E2",X"D3",X"E5",X"34",X"ED",
		X"7D",X"F3",X"61",X"FA",X"D5",X"00",X"AA",X"07",X"59",X"0E",X"A6",X"14",X"DF",X"1B",X"79",X"1C",
		X"F6",X"0E",X"E6",X"00",X"04",X"F3",X"B1",X"E4",X"1B",X"E3",X"45",X"EB",X"31",X"F1",X"19",X"F8",
		X"43",X"FE",X"85",X"05",X"9D",X"0B",X"5B",X"12",X"F4",X"18",X"9D",X"1E",X"C9",X"14",X"0B",X"06",
		X"A7",X"F8",X"73",X"E9",X"51",X"E1",X"70",X"E8",X"89",X"EE",X"93",X"F5",X"BB",X"FB",X"B4",X"02",
		X"C7",X"08",X"90",X"0F",X"78",X"15",X"3F",X"1D",X"AD",X"1A",X"3C",X"0C",X"D3",X"FE",X"BD",X"F0",
		X"5B",X"E3",X"0A",X"E4",X"CB",X"EB",X"C6",X"F1",X"B9",X"F8",X"1D",X"FF",X"DA",X"05",X"EE",X"0B",
		X"BF",X"12",X"32",X"19",X"DA",X"1E",X"5C",X"14",X"B9",X"05",X"CF",X"F8",X"D5",X"E9",X"40",X"E1",
		X"E1",X"E7",X"29",X"EE",X"05",X"F5",X"FC",X"FA",X"15",X"02",X"3E",X"08",X"0F",X"0F",X"AB",X"14",
		X"7D",X"1C",X"1B",X"1C",X"5B",X"0E",X"8D",X"00",X"16",X"F3",X"C3",X"E4",X"BB",X"E2",X"96",X"EA",
		X"2F",X"F0",X"84",X"F7",X"85",X"FD",X"4A",X"04",X"54",X"0A",X"6B",X"11",X"14",X"17",X"4F",X"1E",
		X"9C",X"18",X"09",X"0A",X"BD",X"FC",X"CE",X"EE",X"40",X"E2",X"1C",X"E5",X"45",X"EC",X"7F",X"F2",
		X"3A",X"F9",X"4A",X"FF",X"E6",X"05",X"50",X"0C",X"93",X"12",X"DC",X"18",X"99",X"1E",X"18",X"15",
		X"75",X"06",X"BC",X"F9",X"4D",X"EB",X"68",X"E1",X"04",X"E7",X"8C",X"ED",X"E6",X"F3",X"30",X"FA",
		X"B7",X"00",X"F1",X"06",X"80",X"0D",X"8E",X"13",X"94",X"1A",X"29",X"1E",X"8A",X"12",X"8B",X"04",
		X"A0",X"F7",X"29",X"E9",X"CA",X"E1",X"F1",X"E7",X"22",X"EE",X"BA",X"F4",X"F2",X"FA",X"9E",X"01",
		X"A3",X"07",X"54",X"0E",X"2C",X"14",X"25",X"1B",X"4E",X"1D",X"9C",X"11",X"AE",X"03",X"CE",X"F6",
		X"41",X"E8",X"2C",X"E1",X"82",X"E8",X"4E",X"EE",X"15",X"F5",X"26",X"FB",X"D7",X"01",X"B8",X"07",
		X"4F",X"0E",X"2C",X"14",X"1F",X"1B",X"9C",X"1D",X"7D",X"11",X"A1",X"03",X"D3",X"F6",X"BD",X"E8",
		X"83",X"E1",X"1F",X"E8",X"06",X"EE",X"C1",X"F4",X"E5",X"FA",X"76",X"01",X"71",X"07",X"01",X"0E",
		X"AE",X"13",X"95",X"1A",X"68",X"1E",X"C3",X"12",X"C9",X"04",X"01",X"F8",X"E7",X"E9",X"8C",X"E1",
		X"2F",X"E7",X"75",X"ED",X"CB",X"F3",X"0C",X"FA",X"7C",X"00",X"B2",X"06",X"F2",X"0C",X"0E",X"13",
		X"44",X"19",X"CF",X"1E",X"16",X"15",X"29",X"07",X"6D",X"FA",X"A1",X"EC",X"04",X"E2",X"89",X"E5",
		X"90",X"EC",X"5A",X"F2",X"FA",X"F8",X"D5",X"FE",X"6A",X"05",X"30",X"0B",X"DF",X"11",X"53",X"17",
		X"46",X"1E",X"87",X"18",X"A2",X"0A",X"E3",X"FD",X"93",X"F0",X"78",X"E3",X"60",X"E3",X"01",X"EB",
		X"5A",X"F0",X"27",X"F7",X"C4",X"FC",X"82",X"03",X"14",X"09",X"E9",X"0F",X"58",X"15",X"84",X"1C",
		X"32",X"1C",X"63",X"0F",X"12",X"02",X"84",X"F5",X"89",X"E7",X"D0",X"E1",X"76",X"E8",X"22",X"EE",
		X"D0",X"F4",X"8A",X"FA",X"FE",X"00",X"DE",X"06",X"37",X"0D",X"37",X"13",X"79",X"19",X"92",X"1E",
		X"89",X"15",X"CE",X"07",X"46",X"FB",X"C8",X"ED",X"E9",X"E1",X"A5",X"E4",X"E6",X"EB",X"4B",X"F1",
		X"1C",X"F8",X"9A",X"FD",X"49",X"04",X"D5",X"09",X"98",X"10",X"A5",X"15",X"3E",X"1D",X"21",X"1C",
		X"C3",X"0E",X"CC",X"01",X"3D",X"F5",X"60",X"E7",X"8F",X"E1",X"5B",X"E8",X"EF",X"ED",X"60",X"F4",
		X"5A",X"FA",X"91",X"00",X"94",X"06",X"97",X"0C",X"C2",X"12",X"7F",X"18",X"BF",X"1E",X"8F",X"17",
		X"87",X"09",X"3D",X"FD",X"12",X"F0",X"85",X"E3",X"42",X"E3",X"D4",X"EA",X"E0",X"EF",X"A9",X"F6",
		X"0C",X"FC",X"B3",X"02",X"21",X"08",X"D6",X"0E",X"29",X"14",X"08",X"1B",X"0B",X"1E",X"71",X"13",
		X"F6",X"05",X"B5",X"F9",X"48",X"EC",X"C3",X"E1",X"3D",X"E5",X"14",X"EC",X"9C",X"F1",X"19",X"F8",
		X"87",X"FD",X"19",X"04",X"88",X"09",X"24",X"10",X"4F",X"15",X"78",X"1C",X"99",X"1C",X"AF",X"10",
		X"99",X"03",X"7A",X"F7",X"CE",X"E9",X"A4",X"E1",X"80",X"E6",X"EF",X"EC",X"84",X"F2",X"F9",X"F8",
		X"5D",X"FE",X"FC",X"04",X"43",X"0A",X"FF",X"10",X"E0",X"15",X"58",X"1D",X"00",X"1C",X"5C",X"0F",
		X"6A",X"02",X"5A",X"F6",X"C6",X"E8",X"9C",X"E1",X"1C",X"E7",X"33",X"ED",X"E1",X"F2",X"2F",X"F9",
		X"C3",X"FE",X"1B",X"05",X"6F",X"0A",X"19",X"11",X"EF",X"15",X"51",X"1D",X"24",X"1C",X"4B",X"0F",
		X"A0",X"02",X"80",X"F6",X"12",X"E9",X"55",X"E1",X"F1",X"E6",X"DA",X"EC",X"B2",X"F2",X"D6",X"F8",
		X"73",X"FE",X"9C",X"04",X"1F",X"0A",X"7A",X"10",X"9D",X"15",X"A0",X"1C",X"27",X"1D",X"98",X"10",
		X"1C",X"04",X"D3",X"F7",X"DF",X"EA",X"7F",X"E1",X"FD",X"E5",X"1B",X"EC",X"DD",X"F1",X"D2",X"F7",
		X"8F",X"FD",X"8E",X"03",X"3F",X"09",X"37",X"0F",X"CD",X"14",X"12",X"1B",X"1C",X"1E",X"4F",X"13",
		X"BF",X"06",X"58",X"FA",X"03",X"EE",X"83",X"E2",X"40",X"E4",X"C9",X"EA",X"5A",X"F0",X"5C",X"F6",
		X"18",X"FC",X"F0",X"01",X"C3",X"07",X"75",X"0D",X"62",X"13",X"DD",X"18",X"A4",X"1E",X"85",X"17",
		X"74",X"0A",X"53",X"FE",X"32",X"F2",X"43",X"E5",X"00",X"E2",X"FA",X"E8",X"15",X"EE",X"6C",X"F4",
		X"CE",X"F9",X"E1",X"FF",X"70",X"05",X"4B",X"0B",X"0D",X"11",X"98",X"16",X"E7",X"1C",X"42",X"1C",
		X"88",X"0F",X"C0",X"03",X"3E",X"F7",X"0A",X"EB",X"FE",X"E0",X"FB",X"E5",X"8E",X"EB",X"A5",X"F1",
		X"18",X"F7",X"2A",X"FD",X"90",X"02",X"9E",X"08",X"FA",X"0D",X"0A",X"14",X"5D",X"19",X"BC",X"1E",
		X"83",X"16",X"10",X"0A",X"C2",X"FD",X"18",X"F2",X"02",X"E5",X"E2",X"E1",X"DE",X"E8",X"E9",X"ED",
		X"22",X"F4",X"7C",X"F9",X"7A",X"FF",X"F0",X"04",X"C9",X"0A",X"5B",X"10",X"F8",X"15",X"F6",X"1B",
		X"8B",X"1D",X"A8",X"11",X"F2",X"05",X"7B",X"F9",X"CE",X"ED",X"28",X"E2",X"4F",X"E4",X"57",X"EA",
		X"07",X"F0",X"A1",X"F5",X"76",X"FB",X"EB",X"00",X"D2",X"06",X"20",X"0C",X"2F",X"12",X"29",X"17",
		X"E2",X"1D",X"77",X"1B",X"89",X"0E",X"0A",X"03",X"CD",X"F6",X"D2",X"EA",X"3B",X"E1",X"CC",X"E5",
		X"61",X"EB",X"40",X"F1",X"AA",X"F6",X"90",X"FC",X"E4",X"01",X"D0",X"07",X"0C",X"0D",X"10",X"13",
		X"0D",X"18",X"60",X"1E",X"D3",X"19",X"0E",X"0D",X"7C",X"01",X"88",X"F5",X"5E",X"E9",X"49",X"E1",
		X"74",X"E6",X"D6",X"EB",X"BC",X"F1",X"10",X"F7",X"F0",X"FC",X"3D",X"02",X"1A",X"08",X"53",X"0D",
		X"44",X"13",X"44",X"18",X"6C",X"1E",X"9B",X"19",X"EE",X"0C",X"76",X"01",X"8D",X"F5",X"87",X"E9",
		X"43",X"E1",X"4F",X"E6",X"A9",X"EB",X"89",X"F1",X"CE",X"F6",X"AC",X"FC",X"E3",X"01",X"C3",X"07",
		X"E1",X"0C",X"E0",X"12",X"B1",X"17",X"45",X"1E",X"F1",X"1A",X"27",X"0E",X"EA",X"02",X"E9",X"F6",
		X"3F",X"EB",X"31",X"E1",X"4B",X"E5",X"F1",X"EA",X"8D",X"F0",X"FB",X"F5",X"A0",X"FB",X"FB",X"00",
		X"A3",X"06",X"E9",X"0B",X"A4",X"11",X"B2",X"16",X"E2",X"1C",X"D3",X"1C",X"05",X"11",X"B5",X"05",
		X"BA",X"F9",X"70",X"EE",X"E9",X"E2",X"74",X"E3",X"A6",X"E9",X"D0",X"EE",X"89",X"F4",X"D9",X"F9",
		X"73",X"FF",X"C9",X"04",X"56",X"0A",X"AC",X"0F",X"26",X"15",X"98",X"1A",X"C5",X"1E",X"8B",X"15",
		X"C6",X"09",X"1B",X"FE",X"E1",X"F2",X"A5",X"E6",X"87",X"E1",X"81",X"E7",X"7D",X"EC",X"5B",X"F2",
		X"73",X"F7",X"37",X"FD",X"4E",X"02",X"0E",X"08",X"12",X"0D",X"E5",X"12",X"AC",X"17",X"FB",X"1D",
		X"5A",X"1B",X"2E",X"0F",X"1C",X"04",X"58",X"F8",X"19",X"ED",X"4D",X"E2",X"F9",X"E3",X"F8",X"E9",
		X"1D",X"EF",X"B9",X"F4",X"F6",X"F9",X"7F",X"FF",X"B9",X"04",X"3C",X"0A",X"6B",X"0F",X"EC",X"14",
		X"1B",X"1A",X"C2",X"1E",X"E0",X"16",X"04",X"0B",X"B0",X"FF",X"79",X"F4",X"98",X"E8",X"FC",X"E0",
		X"57",X"E6",X"79",X"EB",X"19",X"F1",X"3F",X"F6",X"CD",X"FB",X"F4",X"00",X"77",X"06",X"98",X"0B",
		X"1C",X"11",X"1C",X"16",X"EE",X"1B",X"2B",X"1E",X"B1",X"13",X"7A",X"08",X"ED",X"FC",X"0C",X"F2",
		X"13",X"E6",X"98",X"E1",X"8E",X"E7",X"72",X"EC",X"25",X"F2",X"28",X"F7",X"C0",X"FC",X"C8",X"01",
		X"54",X"07",X"53",X"0C",X"E8",X"11",X"B8",X"16",X"BF",X"1C",X"98",X"1D",X"50",X"12",X"72",X"07",
		X"D1",X"FB",X"26",X"F1",X"37",X"E5",X"DC",X"E1",X"E3",X"E7",X"BF",X"EC",X"5D",X"F2",X"65",X"F7",
		X"E1",X"FC",X"F0",X"01",X"5E",X"07",X"68",X"0C",X"DA",X"11",X"BE",X"16",X"8A",X"1C",X"A2",X"1D",
		X"B9",X"12",X"EB",X"07",X"56",X"FC",X"DF",X"F1",X"B1",X"E5",X"5A",X"E1",X"81",X"E7",X"42",X"EC",
		X"DE",X"F1",X"D7",X"F6",X"48",X"FC",X"52",X"01",X"AC",X"06",X"BB",X"0B",X"0B",X"11",X"0A",X"16",
		X"81",X"1B",X"C0",X"1E",X"F9",X"14",X"CC",X"09",X"AC",X"FE",X"E5",X"F3",X"5C",X"E8",X"44",X"E1",
		X"09",X"E6",X"2F",X"EB",X"7C",X"F0",X"A2",X"F5",X"DA",X"FA",X"06",X"00",X"29",X"05",X"5E",X"0A",
		X"69",X"0F",X"B0",X"14",X"92",X"19",X"CC",X"1E",X"11",X"19",X"1F",X"0D",X"B9",X"02",X"60",X"F7",
		X"CC",X"EC",X"40",X"E2",X"AD",X"E3",X"67",X"E9",X"58",X"EE",X"A8",X"F3",X"B1",X"F8",X"EF",X"FD",
		X"F4",X"02",X"31",X"08",X"24",X"0D",X"71",X"12",X"2C",X"17",X"F5",X"1C",X"CF",X"1D",X"74",X"12",
		X"1B",X"08",X"B3",X"FC",X"86",X"F2",X"B2",X"E6",X"23",X"E1",X"AC",X"E6",X"88",X"EB",X"DA",X"F0",
		X"D7",X"F5",X"07",X"FB",X"12",X"00",X"2B",X"05",X"3F",X"0A",X"3F",X"0F",X"63",X"14",X"3B",X"19",
		X"79",X"1E",X"36",X"1A",X"6E",X"0E",X"50",X"04",X"F9",X"F8",X"DB",X"EE",X"8F",X"E3",X"8F",X"E2",
		X"4A",X"E8",X"18",X"ED",X"59",X"F2",X"50",X"F7",X"6F",X"FC",X"6E",X"01",X"7D",X"06",X"7E",X"0B",
		X"81",X"10",X"7F",X"15",X"85",X"1A",X"C8",X"1E",X"CC",X"17",X"6D",X"0C",X"24",X"02",X"29",X"F7",
		X"D1",X"EC",X"6A",X"E2",X"62",X"E3",X"07",X"E9",X"CE",X"ED",X"02",X"F3",X"ED",X"F7",X"02",X"FD",
		X"F4",X"01",X"FB",X"06",X"EB",X"0B",X"E8",X"10",X"D3",X"15",X"D9",X"1A",X"D0",X"1E",X"55",X"17",
		X"11",X"0C",X"E4",X"01",X"F6",X"F6",X"CC",X"EC",X"12",X"E2",X"41",X"E3",X"FB",X"E8",X"A3",X"ED",
		X"DA",X"F2",X"AE",X"F7",X"C5",X"FC",X"A0",X"01",X"A3",X"06",X"84",X"0B",X"77",X"10",X"5D",X"15",
		X"41",X"1A",X"D1",X"1E",X"C3",X"18",X"64",X"0D",X"7B",X"03",X"79",X"F8",X"9E",X"EE",X"8D",X"E3",
		X"60",X"E2",X"09",X"E8",X"AC",X"EC",X"CF",X"F1",X"A5",X"F6",X"A2",X"FB",X"84",X"00",X"69",X"05",
		X"58",X"0A",X"23",X"0F",X"27",X"14",X"B8",X"18",X"26",X"1E",X"D2",X"1B",X"91",X"10",X"CD",X"06",
		X"D4",X"FB",X"1D",X"F2",X"DA",X"E6",X"31",X"E1",X"1A",X"E6",X"EE",X"EA",X"E3",X"EF",X"C7",X"F4",
		X"A8",X"F9",X"8C",X"FE",X"60",X"03",X"47",X"08",X"0B",X"0D",X"F7",X"11",X"A2",X"16",X"BB",X"1B",
		X"A2",X"1E",X"2A",X"16",X"72",X"0B",X"65",X"01",X"E1",X"F6",X"E5",X"EC",X"A0",X"E2",X"01",X"E3",
		X"7D",X"E8",X"0F",X"ED",X"18",X"F2",X"D6",X"F6",X"BC",X"FB",X"88",X"00",X"55",X"05",X"2E",X"0A",
		X"E0",X"0E",X"D0",X"13",X"49",X"18",X"A5",X"1D",X"D9",X"1C",X"38",X"12",X"6A",X"08",X"DA",X"FD",
		X"0C",X"F4",X"64",X"E9",X"65",X"E1",X"98",X"E4",X"B4",X"E9",X"61",X"EE",X"49",X"F3",X"04",X"F8",
		X"DA",X"FC",X"9B",X"01",X"5B",X"06",X"27",X"0B",X"CD",X"0F",X"B0",X"14",X"1F",X"19",X"51",X"1E",
		X"A1",X"1B",X"A3",X"10",X"16",X"07",X"86",X"FC",X"ED",X"F2",X"3A",X"E8",X"50",X"E1",X"18",X"E5",
		X"08",X"EA",X"BF",X"EE",X"8C",X"F3",X"49",X"F8",X"04",X"FD",X"C6",X"01",X"6D",X"06",X"3B",X"0B",
		X"C7",X"0F",X"AE",X"14",X"FC",X"18",X"50",X"1E",X"EA",X"1B",X"2E",X"11",X"A2",X"07",X"42",X"FD",
		X"A5",X"F3",X"35",X"E9",X"65",X"E1",X"83",X"E4",X"81",X"E9",X"21",X"EE",X"E6",X"F2",X"97",X"F7",
		X"45",X"FC",X"FF",X"00",X"99",X"05",X"5E",X"0A",X"DB",X"0E",X"B8",X"13",X"FC",X"17",X"49",X"1D",
		X"A0",X"1D",X"DA",X"13",X"08",X"0A",X"11",X"00",X"30",X"F6",X"66",X"EC",X"B5",X"E2",X"C2",X"E2",
		X"31",X"E8",X"75",X"EC",X"6F",X"F1",X"DE",X"F5",X"B7",X"FA",X"2F",X"FF",X"F6",X"03",X"6F",X"08",
		X"2D",X"0D",X"A1",X"11",X"5D",X"16",X"C7",X"1A",X"15",X"1F",X"D8",X"18",X"46",X"0E",X"E9",X"04",
		X"B7",X"FA",X"6C",X"F1",X"E9",X"E6",X"0E",X"E1",X"9B",X"E5",X"11",X"EA",X"DC",X"EE",X"5A",X"F3",
		X"15",X"F8",X"92",X"FC",X"45",X"01",X"B8",X"05",X"6C",X"0A",X"CF",X"0E",X"90",X"13",X"CB",X"17",
		X"D9",X"1C",X"40",X"1E",X"19",X"15",X"49",X"0B",X"AB",X"01",X"D4",X"F7",X"75",X"EE",X"3F",X"E4",
		X"AA",X"E1",X"0B",X"E7",X"1A",X"EB",X"1C",X"F0",X"52",X"F4",X"34",X"F9",X"74",X"FD",X"49",X"02",
		X"80",X"06",X"57",X"0B",X"7D",X"0F",X"65",X"14",X"55",X"18",X"B1",X"1D",X"7B",X"1D",X"D9",X"13",
		X"4B",X"0A",X"B7",X"00",X"04",X"F7",X"BD",X"ED",X"B3",X"E3",X"C4",X"E1",X"45",X"E7",X"3D",X"EB",
		X"36",X"F0",X"5E",X"F4",X"36",X"F9",X"66",X"FD",X"2F",X"02",X"5D",X"06",X"24",X"0B",X"43",X"0F",
		X"1A",X"14",X"03",X"18",X"41",X"1D",X"1F",X"1E",X"FD",X"14",X"60",X"0B",X"07",X"02",X"4D",X"F8",
		X"43",X"EF",X"0B",X"E5",X"28",X"E1",X"5B",X"E6",X"6B",X"EA",X"36",X"EF",X"75",X"F3",X"1B",X"F8",
		X"69",X"FC",X"FB",X"00",X"4C",X"05",X"D1",X"09",X"23",X"0E",X"9C",X"12",X"EE",X"16",X"69",X"1B",
		X"F2",X"1E",X"92",X"18",X"8C",X"0E",X"82",X"05",X"D5",X"FB",X"C6",X"F2",X"09",X"E9",X"7D",X"E1",
		X"EF",X"E3",X"D7",X"E8",X"FC",X"EC",X"AC",X"F1",X"DA",X"F5",X"82",X"FA",X"A6",X"FE",X"4E",X"03",
		X"65",X"07",X"11",X"0C",X"12",X"10",X"D3",X"14",X"9E",X"18",X"C6",X"1D",X"65",X"1D",X"48",X"14",
		X"E5",X"0A",X"C4",X"01",X"3F",X"F8",X"66",X"EF",X"7B",X"E5",X"43",X"E1",X"CF",X"E5",X"16",X"EA",
		X"83",X"EE",X"E9",X"F2",X"36",X"F7",X"AD",X"FB",X"DF",X"FF",X"65",X"04",X"7A",X"08",X"17",X"0D",
		X"04",X"11",X"C5",X"15",X"67",X"19",X"BD",X"1E",X"68",X"1C",X"91",X"12",X"94",X"09",X"64",X"00",
		X"1A",X"F7",X"4B",X"EE",X"87",X"E4",X"76",X"E1",X"43",X"E6",X"56",X"EA",X"D3",X"EE",X"15",X"F3",
		X"6A",X"F7",X"C0",X"FB",X"F7",X"FF",X"5D",X"04",X"77",X"08",X"F1",X"0C",X"E9",X"10",X"85",X"15",
		X"37",X"19",X"5D",X"1E",X"09",X"1D",X"71",X"13",X"95",X"0A",X"70",X"01",X"58",X"F8",X"83",X"EF",
		X"04",X"E6",X"1A",X"E1",X"6D",X"E5",X"86",X"E9",X"F8",X"ED",X"20",X"F2",X"7B",X"F6",X"AC",X"FA",
		X"F6",X"FE",X"2C",X"03",X"66",X"07",X"9D",X"0B",X"CB",X"0F",X"07",X"14",X"1C",X"18",X"85",X"1C",
		X"CE",X"1E",X"FC",X"16",X"DA",X"0D",X"E6",X"04",X"FB",X"FB",X"06",X"F3",X"22",X"EA",X"D0",X"E1",
		X"17",X"E3",X"CB",X"E7",X"D0",X"EB",X"2D",X"F0",X"4E",X"F4",X"94",X"F8",X"BE",X"FC",X"EE",X"00",
		X"22",X"05",X"3E",X"09",X"7C",X"0D",X"7D",X"11",X"D9",X"15",X"97",X"19",X"73",X"1E",X"07",X"1D",
		X"5B",X"13",X"F3",X"0A",X"CA",X"01",X"2B",X"F9",X"46",X"F0",X"59",X"E7",X"C8",X"E0",X"A4",X"E4",
		X"A3",X"E8",X"0E",X"ED",X"01",X"F1",X"64",X"F5",X"52",X"F9",X"B0",X"FD",X"98",X"01",X"F1",X"05",
		X"D0",X"09",X"2E",X"0E",X"F6",X"11",X"68",X"16",X"FD",X"19",X"C6",X"1E",X"3B",X"1C",X"D4",X"12",
		X"5F",X"0A",X"7B",X"01",X"D5",X"F8",X"2F",X"F0",X"3E",X"E7",X"BD",X"E0",X"84",X"E4",X"8A",X"E8",
		X"D2",X"EC",X"CC",X"F0",X"0D",X"F5",X"02",X"F9",X"3E",X"FD",X"2E",X"01",X"64",X"05",X"4C",X"09",
		X"84",X"0D",X"5A",X"11",X"A1",X"15",X"4B",X"19",X"EE",X"1D",X"AB",X"1D",X"E8",X"14",X"7B",X"0C",
		X"AB",X"03",X"3C",X"FB",X"7F",X"F2",X"12",X"EA",X"D8",X"E1",X"C7",X"E2",X"67",X"E7",X"33",X"EB",
		X"79",X"EF",X"60",X"F3",X"91",X"F7",X"79",X"FB",X"A1",X"FF",X"84",X"03",X"AB",X"07",X"84",X"0B",
		X"AA",X"0F",X"78",X"13",X"A2",X"17",X"60",X"1B",X"32",X"1F",X"F7",X"19",X"03",X"11",X"9E",X"08",
		X"1C",X"00",X"8C",X"F7",X"4E",X"EF",X"5D",X"E6",X"CE",X"E0",X"AE",X"E4",X"93",X"E8",X"B8",X"EC",
		X"A3",X"F0",X"B6",X"F4",X"A8",X"F8",X"AC",X"FC",X"9E",X"00",X"97",X"04",X"8C",X"08",X"78",X"0C",
		X"6C",X"10",X"50",X"14",X"3E",X"18",X"30",X"1C",X"1C",X"1F",X"A5",X"18",X"01",X"10",X"A1",X"07",
		X"50",X"FF",X"CE",X"F6",X"BC",X"EE",X"DE",X"E5",X"F0",X"E0",X"CD",X"E4",X"A1",X"E8",X"B7",X"EC",
		X"98",X"F0",X"98",X"F4",X"80",X"F8",X"70",X"FC",X"5B",X"00",X"3E",X"04",X"2C",X"08",X"02",X"0C",
		X"F5",X"0F",X"B9",X"13",X"B6",X"17",X"5F",X"1B",X"51",X"1F",X"84",X"1A",X"A4",X"11",X"A8",X"09",
		X"30",X"01",X"17",X"F9",X"C6",X"F0",X"90",X"E8",X"27",X"E1",X"4B",X"E3",X"78",X"E7",X"47",X"EB",
		X"3F",X"EF",X"18",X"F3",X"04",X"F7",X"DD",X"FA",X"C2",X"FE",X"93",X"02",X"75",X"06",X"3F",X"0A",
		X"21",X"0E",X"DC",X"11",X"C8",X"15",X"61",X"19",X"92",X"1D",X"58",X"1E",X"63",X"16",X"5E",X"0E",
		X"04",X"06",X"18",X"FE",X"BB",X"F5",X"FA",X"ED",X"51",X"E5",X"DE",X"E0",X"DB",X"E4",X"8B",X"E8",
		X"88",X"EC",X"46",X"F0",X"2F",X"F4",X"F4",X"F7",X"D0",X"FB",X"96",X"FF",X"63",X"03",X"2C",X"07",
		X"EE",X"0A",X"BD",X"0E",X"6C",X"12",X"4A",X"16",X"CD",X"19",X"FC",X"1D",X"0D",X"1E",X"B3",X"15",
		X"FA",X"0D",X"A4",X"05",X"ED",X"FD",X"9D",X"F5",X"09",X"EE",X"73",X"E5",X"F8",X"E0",X"99",X"E4",
		X"54",X"E8",X"30",X"EC",X"F0",X"EF",X"BD",X"F3",X"7D",X"F7",X"42",X"FB",X"01",X"FF",X"BB",X"02",
		X"79",X"06",X"2C",X"0A",X"E8",X"0D",X"92",X"11",X"4F",X"15",X"E8",X"18",X"C1",X"1C",X"2C",X"1F",
		X"93",X"18",X"5C",X"10",X"9A",X"08",X"95",X"00",X"D5",X"F8",X"DA",X"F0",X"23",X"E9",X"A2",X"E1",
		X"96",X"E2",X"C5",X"E6",X"50",X"EA",X"2B",X"EE",X"D1",X"F1",X"92",X"F5",X"42",X"F9",X"F5",X"FC",
		X"A6",X"00",X"4B",X"04",X"00",X"08",X"98",X"0B",X"55",X"0F",X"D4",X"12",X"A4",X"16",X"FA",X"19",
		X"1D",X"1E",X"13",X"1E",X"10",X"16",X"79",X"0E",X"85",X"06",X"E3",X"FE",X"08",X"F7",X"6D",X"EF",
		X"8A",X"E7",X"F1",X"E0",X"42",X"E3",X"38",X"E7",X"C8",X"EA",X"86",X"EE",X"24",X"F2",X"D1",X"F5",
		X"73",X"F9",X"14",X"FD",X"B8",X"00",X"4E",X"04",X"F3",X"07",X"7C",X"0B",X"28",X"0F",X"A0",X"12",
		X"54",X"16",X"AB",X"19",X"A1",X"1D",X"96",X"1E",X"57",X"17",X"A2",X"0F",X"00",X"08",X"50",X"00",
		X"C7",X"F8",X"0F",X"F1",X"AC",X"E9",X"E3",X"E1",X"00",X"E2",X"42",X"E6",X"88",X"E9",X"65",X"ED",
		X"CD",X"F0",X"91",X"F4",X"02",X"F8",X"B5",X"FB",X"28",X"FF",X"D3",X"02",X"42",X"06",X"E9",X"09",
		X"52",X"0D",X"F7",X"10",X"54",X"14",X"04",X"18",X"3F",X"1B",X"0E",X"1F",X"2A",X"1C",X"10",X"14",
		X"D7",X"0C",X"19",X"05",X"C9",X"FD",X"22",X"F6",X"DD",X"EE",X"22",X"E7",X"07",X"E1",X"33",X"E3",
		X"04",X"E7",X"6E",X"EA",X"19",X"EE",X"8B",X"F1",X"29",X"F5",X"98",X"F8",X"30",X"FC",X"9B",X"FF",
		X"2F",X"03",X"93",X"06",X"27",X"0A",X"81",X"0D",X"18",X"11",X"60",X"14",X"05",X"18",X"28",X"1B",
		X"02",X"1F",X"89",X"1C",X"A0",X"14",X"81",X"0D",X"EC",X"05",X"B1",X"FE",X"3F",X"F7",X"FC",X"EF",
		X"9F",X"E8",X"B5",X"E1",X"3E",X"E2",X"4A",X"E6",X"75",X"E9",X"34",X"ED",X"77",X"F0",X"22",X"F4",
		X"6A",X"F7",X"0A",X"FB",X"50",X"FE",X"E8",X"01",X"2C",X"05",X"BF",X"08",X"FE",X"0B",X"8C",X"0F",
		X"C4",X"12",X"53",X"16",X"7A",X"19",X"2C",X"1D",X"0F",X"1F",X"24",X"19",X"90",X"11",X"80",X"0A",
		X"14",X"03",X"07",X"FC",X"A2",X"F4",X"AE",X"ED",X"26",X"E6",X"D3",X"E0",X"70",X"E3",X"0D",X"E7",
		X"61",X"EA",X"E4",X"ED",X"38",X"F1",X"B5",X"F4",X"06",X"F8",X"7B",X"FB",X"C9",X"FE",X"39",X"02",
		X"84",X"05",X"EE",X"08",X"34",X"0C",X"99",X"0F",X"DB",X"12",X"3B",X"16",X"77",X"19",X"E6",X"1C",
		X"37",X"1F",X"C4",X"19",X"57",X"12",X"5A",X"0B",X"29",X"04",X"20",X"FD",X"05",X"F6",X"FC",X"EE",
		X"EC",X"E7",X"55",X"E1",X"64",X"E2",X"2A",X"E6",X"52",X"E9",X"D4",X"EC",X"12",X"F0",X"81",X"F3",
		X"C4",X"F6",X"25",X"FA",X"6B",X"FD",X"BE",X"00",X"07",X"04",X"50",X"07",X"9C",X"0A",X"D9",X"0D",
		X"29",X"11",X"54",X"14",X"B4",X"17",X"B5",X"1A",X"63",X"1E",X"2E",X"1E",X"F2",X"16",X"29",X"10",
		X"04",X"09",X"2D",X"02",X"25",X"FB",X"48",X"F4",X"5D",X"ED",X"5C",X"E6",X"98",X"E0",X"2D",X"E3",
		X"8A",X"E6",X"DC",X"E9",X"1E",X"ED",X"70",X"F0",X"AC",X"F3",X"FA",X"F6",X"32",X"FA",X"7B",X"FD",
		X"AE",X"00",X"F2",X"03",X"21",X"07",X"61",X"0A",X"8B",X"0D",X"C8",X"10",X"EA",X"13",X"2A",X"17",
		X"34",X"1A",X"A6",X"1D",X"FA",X"1E",X"BD",X"18",X"E8",X"11",X"FB",X"0A",X"43",X"04",X"56",X"FD",
		X"B6",X"F6",X"BB",X"EF",X"49",X"E9",X"0D",X"E2",X"5F",X"E1",X"4A",X"E5",X"28",X"E8",X"A6",X"EB",
		X"A9",X"EE",X"0B",X"F2",X"18",X"F5",X"6C",X"F8",X"7B",X"FB",X"C6",X"FE",X"D3",X"01",X"17",X"05",
		X"21",X"08",X"62",X"0B",X"66",X"0E",X"A5",X"11",X"9D",X"14",X"E6",X"17",X"C0",X"1A",X"4B",X"1E",
		X"74",X"1E",X"C2",X"17",X"36",X"11",X"5E",X"0A",X"D5",X"03",X"0A",X"FD",X"90",X"F6",X"BF",X"EF",
		X"68",X"E9",X"75",X"E2",X"52",X"E1",X"EF",X"E4",X"D8",X"E7",X"2E",X"EB",X"34",X"EE",X"71",X"F1",
		X"7F",X"F4",X"B0",X"F7",X"C1",X"FA",X"E7",X"FD",X"F8",X"00",X"14",X"04",X"24",X"07",X"3A",X"0A",
		X"4B",X"0D",X"54",X"10",X"6A",X"13",X"65",X"16",X"82",X"19",X"6A",X"1C",X"68",X"1F",X"C5",X"1B",
		X"AD",X"14",X"6C",X"0E",X"AB",X"07",X"53",X"01",X"AE",X"FA",X"56",X"F4",X"BE",X"ED",X"68",X"E7",
		X"3B",X"E1",X"28",X"E2",X"8D",X"E5",X"85",X"E8",X"AF",X"EB",X"B5",X"EE",X"D0",X"F1",X"DA",X"F4",
		X"EB",X"F7",X"F4",X"FA",X"FE",X"FD",X"03",X"01",X"07",X"04",X"0B",X"07",X"09",X"0A",X"0C",X"0D",
		X"00",X"10",X"07",X"13",X"EB",X"15",X"FF",X"18",X"BE",X"1B",X"0B",X"1F",X"64",X"1D",X"69",X"16",
		X"60",X"10",X"B2",X"09",X"96",X"03",X"FD",X"FC",X"EC",X"F6",X"52",X"F0",X"62",X"EA",X"87",X"E3",
		X"B5",X"E0",X"FE",X"E3",X"D9",X"E6",X"F9",X"E9",X"E9",X"EC",X"F9",X"EF",X"EC",X"F2",X"F0",X"F5",
		X"E0",X"F8",X"E2",X"FB",X"D0",X"FE",X"CA",X"01",X"B2",X"04",X"AB",X"07",X"8C",X"0A",X"84",X"0D",
		X"5E",X"10",X"59",X"13",X"23",X"16",X"2B",X"19",X"D2",X"1B",X"10",X"1F",X"6B",X"1D",X"BE",X"16",
		X"C5",X"10",X"54",X"0A",X"4B",X"04",X"F3",X"FD",X"ED",X"F7",X"9A",X"F1",X"AA",X"EB",X"34",X"E5",
		X"95",X"E0",X"EF",X"E2",X"F7",X"E5",X"E1",X"E8",X"D6",X"EB",X"C0",X"EE",X"B1",X"F1",X"96",X"F4",
		X"81",X"F7",X"61",X"FA",X"4B",X"FD",X"26",X"00",X"0C",X"03",X"E1",X"05",X"C4",X"08",X"93",X"0B",
		X"77",X"0E",X"3C",X"11",X"23",X"14",X"D8",X"16",X"CC",X"19",X"62",X"1C",X"7B",X"1F",X"A8",X"1C",
		X"FC",X"15",X"39",X"10",X"EC",X"09",X"11",X"04",X"DF",X"FD",X"01",X"F8",X"DE",X"F1",X"09",X"EC",
		X"DC",X"E5",X"CE",X"E0",X"62",X"E2",X"86",X"E5",X"3D",X"E8",X"3A",X"EB",X"F8",X"ED",X"EA",X"F0",
		X"AA",X"F3",X"95",X"F6",X"52",X"F9",X"36",X"FC",X"F1",X"FE",X"CD",X"01",X"88",X"04",X"5F",X"07",
		X"17",X"0A",X"E9",X"0C",X"9E",X"0F",X"69",X"12",X"1C",X"15",X"E4",X"17",X"8F",X"1A",X"61",X"1D",
		X"69",X"1F",X"08",X"1B",X"D5",X"14",X"0F",X"0F",X"11",X"09",X"44",X"03",X"58",X"FD",X"8D",X"F7",
		X"AC",X"F1",X"EA",X"EB",X"05",X"E6",X"E3",X"E0",X"2B",X"E2",X"39",X"E5",X"E2",X"E7",X"C2",X"EA",
		X"77",X"ED",X"49",X"F0",X"03",X"F3",X"C9",X"F5",X"84",X"F8",X"43",X"FB",X"FD",X"FD",X"B5",X"00",
		X"6D",X"03",X"1C",X"06",X"D6",X"08",X"7D",X"0B",X"38",X"0E",X"D6",X"10",X"93",X"13",X"24",X"16",
		X"EB",X"18",X"5D",X"1B",X"5F",X"1E",X"16",X"1F",X"5C",X"19",X"B1",X"13",X"E0",X"0D",X"38",X"08",
		X"75",X"02",X"D1",X"FC",X"1C",X"F7",X"7D",X"F1",X"D2",X"EB",X"34",X"E6",X"FF",X"E0",X"E3",X"E1",
		X"F0",X"E4",X"77",X"E7",X"4D",X"EA",X"E4",X"EC",X"AF",X"EF",X"43",X"F2",X"08",X"F5",X"9B",X"F7",
		X"5B",X"FA",X"EB",X"FC",X"A6",X"FF",X"2F",X"02",X"E7",X"04",X"6D",X"07",X"25",X"0A",X"A2",X"0C",
		X"5A",X"0F",X"CF",X"11",X"89",X"14",X"F1",X"16",X"B7",X"19",X"FB",X"1B",X"05",X"1F",X"46",X"1E",
		X"56",X"18",X"F9",X"12",X"42",X"0D",X"D5",X"07",X"36",X"02",X"CB",X"FC",X"33",X"F7",X"D3",X"F1",
		X"3F",X"EC",X"F1",X"E6",X"6A",X"E1",X"5F",X"E1",X"61",X"E4",X"CC",X"E6",X"90",X"E9",X"13",X"EC",
		X"C4",X"EE",X"4C",X"F1",X"F3",X"F3",X"7A",X"F6",X"19",X"F9",X"A0",X"FB",X"3A",X"FE",X"C0",X"00",
		X"53",X"03",X"D6",X"05",X"60",X"08",X"E6",X"0A",X"6B",X"0D",X"EF",X"0F",X"6B",X"12",X"F2",X"14",
		X"5F",X"17",X"F2",X"19",X"40",X"1C",X"0C",X"1F",X"24",X"1E",X"69",X"18",X"45",X"13",X"B0",X"0D",
		X"81",X"08",X"FE",X"02",X"D1",X"FD",X"59",X"F8",X"37",X"F3",X"BC",X"ED",X"B9",X"E8",X"10",X"E3",
		X"90",X"E0",X"38",X"E3",X"A6",X"E5",X"44",X"E8",X"BD",X"EA",X"50",X"ED",X"C9",X"EF",X"54",X"F2",
		X"CE",X"F4",X"54",X"F7",X"C9",X"F9",X"4A",X"FC",X"BC",X"FE",X"3B",X"01",X"A6",X"03",X"23",X"06",
		X"89",X"08",X"06",X"0B",X"67",X"0D",X"E0",X"0F",X"3B",X"12",X"B6",X"14",X"06",X"17",X"85",X"19",
		X"C0",X"1B",X"69",X"1E",X"1D",X"1F",X"44",X"1A",X"03",X"15",X"D8",X"0F",X"9F",X"0A",X"82",X"05",
		X"4C",X"00",X"3F",X"FB",X"07",X"F6",X"0D",X"F1",X"CC",X"EB",X"F8",X"E6",X"81",X"E1",X"ED",X"E0",
		X"DF",X"E3",X"12",X"E6",X"B0",X"E8",X"02",X"EB",X"87",X"ED",X"E3",X"EF",X"5C",X"F2",X"BC",X"F4",
		X"2A",X"F7",X"8C",X"F9",X"F1",X"FB",X"53",X"FE",X"B2",X"00",X"12",X"03",X"6A",X"05",X"C9",X"07",
		X"1B",X"0A",X"7D",X"0C",X"C3",X"0E",X"29",X"11",X"65",X"13",X"CF",X"15",X"FC",X"17",X"73",X"1A",
		X"7D",X"1C",X"39",X"1F",X"42",X"1E",X"F0",X"18",X"1C",X"14",X"00",X"0F",X"16",X"0A",X"13",X"05",
		X"25",X"00",X"37",X"FB",X"45",X"F6",X"6A",X"F1",X"6F",X"EC",X"B5",X"E7",X"8C",X"E2",X"8E",X"E0",
		X"25",X"E3",X"52",X"E5",X"D2",X"E7",X"0F",X"EA",X"7E",X"EC",X"BF",X"EE",X"25",X"F1",X"68",X"F3",
		X"C7",X"F5",X"08",X"F8",X"61",X"FA",X"A2",X"FC",X"F4",X"FE",X"32",X"01",X"81",X"03",X"BC",X"05",
		X"06",X"08",X"3F",X"0A",X"83",X"0C",X"BA",X"0E",X"FC",X"10",X"2E",X"13",X"6D",X"15",X"99",X"17",
		X"DB",X"19",X"F8",X"1B",X"5A",X"1E",X"6A",X"1F",X"05",X"1B",X"38",X"16",X"60",X"11",X"A4",X"0C",
		X"D0",X"07",X"1F",X"03",X"50",X"FE",X"AB",X"F9",X"DD",X"F4",X"49",X"F0",X"74",X"EB",X"FD",X"E6",
		X"FD",X"E1",X"9A",X"E0",X"37",X"E3",X"48",X"E5",X"AE",X"E7",X"D3",X"E9",X"26",X"EC",X"53",X"EE",
		X"9C",X"F0",X"CA",X"F2",X"0D",X"F5",X"3A",X"F7",X"77",X"F9",X"A1",X"FB",X"D9",X"FD",X"03",X"00",
		X"34",X"02",X"5B",X"04",X"89",X"06",X"AE",X"08",X"D8",X"0A",X"F9",X"0C",X"1E",X"0F",X"3E",X"11",
		X"5F",X"13",X"7C",X"15",X"9A",X"17",X"B3",X"19",X"CB",X"1B",X"EA",X"1D",X"A3",X"1F",X"45",X"1C",
		X"73",X"17",X"FB",X"12",X"51",X"0E",X"D4",X"09",X"35",X"05",X"BF",X"00",X"27",X"FC",X"BB",X"F7",
		X"27",X"F3",X"C7",X"EE",X"30",X"EA",X"EA",X"E5",X"3F",X"E1",X"E7",X"E0",X"65",X"E3",X"62",X"E5",
		X"A7",X"E7",X"B9",X"E9",X"ED",X"EB",X"05",X"EE",X"2F",X"F0",X"47",X"F2",X"6B",X"F4",X"85",X"F6",
		X"A1",X"F8",X"B8",X"FA",X"D0",X"FC",X"E7",X"FE",X"F8",X"00",X"0B",X"03",X"19",X"05",X"2D",X"07",
		X"35",X"09",X"46",X"0B",X"4A",X"0D",X"5B",X"0F",X"56",X"11",X"67",X"13",X"5C",X"15",X"71",X"17",
		X"57",X"19",X"78",X"1B",X"44",X"1D",X"85",X"1F",X"EA",X"1D",X"2C",X"19",X"FC",X"14",X"81",X"10",
		X"3F",X"0C",X"DA",X"07",X"94",X"03",X"3F",X"FF",X"FA",X"FA",X"B3",X"F6",X"6C",X"F2",X"36",X"EE",
		X"E7",X"E9",X"CC",X"E5",X"6C",X"E1",X"B7",X"E0",X"18",X"E3",X"F7",X"E4",X"26",X"E7",X"16",X"E9",
		X"38",X"EB",X"2C",X"ED",X"45",X"EF",X"3B",X"F1",X"4B",X"F3",X"40",X"F5",X"4B",X"F7",X"41",X"F9",
		X"45",X"FB",X"3A",X"FD",X"39",X"FF",X"2B",X"01",X"24",X"03",X"18",X"05",X"0D",X"07",X"FB",X"08",
		X"EC",X"0A",X"DB",X"0C",X"C7",X"0E",X"B4",X"10",X"9A",X"12",X"86",X"14",X"64",X"16",X"53",X"18",
		X"2B",X"1A",X"1A",X"1C",X"EA",X"1D",X"B1",X"1F",X"09",X"1D",X"9D",X"18",X"9F",X"14",X"68",X"10",
		X"5D",X"0C",X"37",X"08",X"2D",X"04",X"15",X"00",X"0C",X"FC",X"FE",X"F7",X"F9",X"F3",X"F2",X"EF",
		X"F3",X"EB",X"F8",X"E7",X"F2",X"E3",X"75",X"E0",X"6B",X"E1",X"85",X"E3",X"63",X"E5",X"60",X"E7",
		X"43",X"E9",X"3B",X"EB",X"1D",X"ED",X"10",X"EF",X"EF",X"F0",X"DE",X"F2",X"BB",X"F4",X"A7",X"F6",
		X"80",X"F8",X"69",X"FA",X"3E",X"FC",X"24",X"FE",X"F5",X"FF",X"DA",X"01",X"A6",X"03",X"87",X"05",
		X"53",X"07",X"33",X"09",X"F8",X"0A",X"D6",X"0C",X"96",X"0E",X"73",X"10",X"2F",X"12",X"09",X"14",
		X"C1",X"15",X"9C",X"17",X"4A",X"19",X"2C",X"1B",X"C9",X"1C",X"C8",X"1E",X"6D",X"1F",X"D5",X"1B",
		X"E7",X"17",X"0B",X"14",X"26",X"10",X"53",X"0C",X"71",X"08",X"A7",X"04",X"C8",X"00",X"09",X"FD",
		X"2F",X"F9",X"77",X"F5",X"A1",X"F1",X"F6",X"ED",X"1C",X"EA",X"88",X"E6",X"89",X"E2",X"1D",X"E0",
		X"E7",X"E1",X"B1",X"E3",X"8B",X"E5",X"58",X"E7",X"2A",X"E9",X"F8",X"EA",X"C4",X"EC",X"90",X"EE",
		X"58",X"F0",X"22",X"F2",X"E5",X"F3",X"AD",X"F5",X"6C",X"F7",X"34",X"F9",X"EF",X"FA",X"B4",X"FC",
		X"6A",X"FE",X"2B",X"00",X"DF",X"01",X"9E",X"03",X"50",X"05",X"0B",X"07",X"B9",X"08",X"73",X"0A",
		X"1E",X"0C",X"D4",X"0D",X"7C",X"0F",X"2E",X"11",X"D4",X"12",X"83",X"14",X"29",X"16",X"D4",X"17",
		X"75",X"19",X"1E",X"1B",X"BC",X"1C",X"69",X"1E",X"B1",X"1F",X"F7",X"1C",X"29",X"19",X"A3",X"15",
		X"F6",X"11",X"6C",X"0E",X"C9",X"0A",X"45",X"07",X"A8",X"03",X"2B",X"00",X"95",X"FC",X"1D",X"F9",
		X"8B",X"F5",X"1C",X"F2",X"8E",X"EE",X"29",X"EB",X"98",X"E7",X"47",X"E4",X"B7",X"E0",X"A9",X"E0",
		X"A6",X"E2",X"34",X"E4",X"FD",X"E5",X"9A",X"E7",X"58",X"E9",X"FA",X"EA",X"AE",X"EC",X"4F",X"EE",
		X"FF",X"EF",X"A0",X"F1",X"4D",X"F3",X"E9",X"F4",X"91",X"F6",X"2E",X"F8",X"D1",X"F9",X"6A",X"FB",
		X"0D",X"FD",X"A3",X"FE",X"42",X"00",X"D5",X"01",X"72",X"03",X"02",X"05",X"9B",X"06",X"28",X"08",
		X"BF",X"09",X"49",X"0B",X"DF",X"0C",X"65",X"0E",X"F9",X"0F",X"7B",X"11",X"0D",X"13",X"8B",X"14",
		X"1B",X"16",X"94",X"17",X"24",X"19",X"97",X"1A",X"2C",X"1C",X"8D",X"1D",X"43",X"1F",X"16",X"1F",
		X"A4",X"1B",X"67",X"18",X"01",X"15",X"C0",X"11",X"63",X"0E",X"25",X"0B",X"D3",X"07",X"97",X"04",
		X"4B",X"01",X"18",X"FE",X"D0",X"FA",X"A3",X"F7",X"61",X"F4",X"3D",X"F1",X"F9",X"ED",X"E1",X"EA",
		X"9A",X"E7",X"9D",X"E4",X"2E",X"E1",X"33",X"E0",X"0B",X"E2",X"71",X"E3",X"1B",X"E5",X"94",X"E6",
		X"30",X"E8",X"AB",X"E9",X"40",X"EB",X"BC",X"EC",X"4B",X"EE",X"C6",X"EF",X"52",X"F1",X"CC",X"F2",
		X"53",X"F4",X"CB",X"F5",X"4E",X"F7",X"C5",X"F8",X"46",X"FA",X"B8",X"FB",X"36",X"FD",X"A9",X"FE",
		X"22",X"00",X"90",X"01",X"08",X"03",X"75",X"04",X"E8",X"05",X"52",X"07",X"C3",X"08",X"2C",X"0A",
		X"99",X"0B",X"FF",X"0C",X"6A",X"0E",X"CD",X"0F",X"35",X"11",X"94",X"12",X"FC",X"13",X"58",X"15",
		X"BC",X"16",X"17",X"18",X"79",X"19",X"CE",X"1A",X"32",X"1C",X"7E",X"1D",X"F4",X"1E",X"84",X"1F",
		X"D3",X"1C",X"C5",X"19",X"C2",X"16",X"C2",X"13",X"C1",X"10",X"C6",X"0D",X"CC",X"0A",X"D9",X"07",
		X"E3",X"04",X"F5",X"01",X"06",X"FF",X"1F",X"FC",X"34",X"F9",X"52",X"F6",X"6C",X"F3",X"90",X"F0",
		X"B0",X"ED",X"DB",X"EA",X"FD",X"E7",X"31",X"E5",X"48",X"E2",X"15",X"E0",X"0F",X"E1",X"88",X"E2",
		X"E9",X"E3",X"52",X"E5",X"B6",X"E6",X"1A",X"E8",X"7B",X"E9",X"DD",X"EA",X"3C",X"EC",X"9A",X"ED",
		X"F6",X"EE",X"54",X"F0",X"AD",X"F1",X"06",X"F3",X"5E",X"F4",X"B4",X"F5",X"0A",X"F7",X"5D",X"F8",
		X"B0",X"F9",X"00",X"FB",X"52",X"FC",X"9E",X"FD",X"EE",X"FE",X"36",X"00",X"83",X"01",X"CB",X"02",
		X"15",X"04",X"5B",X"05",X"A3",X"06",X"E4",X"07",X"2B",X"09",X"6A",X"0A",X"AE",X"0B",X"EA",X"0C",
		X"2D",X"0E",X"65",X"0F",X"A6",X"10",X"DB",X"11",X"1A",X"13",X"4D",X"14",X"8A",X"15",X"B7",X"16",
		X"F4",X"17",X"1E",X"19",X"5B",X"1A",X"7E",X"1B",X"BF",X"1C",X"D6",X"1D",X"2F",X"1F",X"81",X"1F",
		X"ED",X"1C",X"45",X"1A",X"96",X"17",X"F2",X"14",X"4C",X"12",X"AC",X"0F",X"0D",X"0D",X"71",X"0A",
		X"D6",X"07",X"3D",X"05",X"AB",X"02",X"17",X"00",X"8C",X"FD",X"FB",X"FA",X"75",X"F8",X"EA",X"F5",
		X"68",X"F3",X"E2",X"F0",X"67",X"EE",X"E6",X"EB",X"6E",X"E9",X"F1",X"E6",X"84",X"E4",X"00",X"E2",
		X"F7",X"DF",X"C9",X"E0",X"19",X"E2",X"4B",X"E3",X"8D",X"E4",X"C0",X"E5",X"FC",X"E6",X"2C",X"E8",
		X"65",X"E9",X"97",X"EA",X"CD",X"EB",X"FB",X"EC",X"2F",X"EE",X"5A",X"EF",X"8B",X"F0",X"B4",X"F1",
		X"E3",X"F2",X"0A",X"F4",X"37",X"F5",X"5B",X"F6",X"85",X"F7",X"A8",X"F8",X"CE",X"F9",X"EF",X"FA",
		X"13",X"FC",X"30",X"FD",X"52",X"FE",X"6E",X"FF",X"8D",X"00",X"A7",X"01",X"C4",X"02",X"DC",X"03",
		X"F5",X"04",X"0B",X"06",X"23",X"07",X"35",X"08",X"4A",X"09",X"5C",X"0A",X"6D",X"0B",X"7D",X"0C",
		X"8D",X"0D",X"9A",X"0E",X"A7",X"0F",X"B5",X"10",X"C0",X"11",X"C8",X"12",X"D0",X"13",X"D8",X"14",
		X"DD",X"15",X"E3",X"16",X"E6",X"17",X"E8",X"18",X"EB",X"19",X"EA",X"1A",X"E9",X"1B",X"E7",X"1C",
		X"E4",X"1D",X"E4",X"1E",X"AD",X"1F",X"0D",X"1E",X"AE",X"1B",X"79",X"19",X"33",X"17",X"FC",X"14",
		X"BB",X"12",X"88",X"10",X"4E",X"0E",X"1E",X"0C",X"EA",X"09",X"BF",X"07",X"8F",X"05",X"6A",X"03",
		X"3E",X"01",X"1E",X"FF",X"F8",X"FC",X"DC",X"FA",X"BA",X"F8",X"A2",X"F6",X"86",X"F4",X"73",X"F2",
		X"5C",X"F0",X"4C",X"EE",X"37",X"EC",X"31",X"EA",X"1E",X"E8",X"1E",X"E6",X"0D",X"E4",X"1A",X"E2",
		X"08",X"E0",X"36",X"E0",X"6A",X"E1",X"5B",X"E2",X"70",X"E3",X"6A",X"E4",X"77",X"E5",X"73",X"E6",
		X"7B",X"E7",X"76",X"E8",X"7B",X"E9",X"74",X"EA",X"75",X"EB",X"6E",X"EC",X"6D",X"ED",X"62",X"EE",
		X"5F",X"EF",X"55",X"F0",X"4F",X"F1",X"41",X"F2",X"38",X"F3",X"2A",X"F4",X"1D",X"F5",X"0D",X"F6",
		X"01",X"F7",X"ED",X"F7",X"DD",X"F8",X"C7",X"F9",X"B5",X"FA",X"9F",X"FB",X"8A",X"FC",X"71",X"FD",
		X"5A",X"FE",X"40",X"FF",X"27",X"00",X"07",X"01",X"ED",X"01",X"CE",X"02",X"B0",X"03",X"8F",X"04",
		X"70",X"05",X"4B",X"06",X"2B",X"07",X"05",X"08",X"E0",X"08",X"BB",X"09",X"94",X"0A",X"6B",X"0B",
		X"42",X"0C",X"17",X"0D",X"EE",X"0D",X"C0",X"0E",X"94",X"0F",X"63",X"10",X"36",X"11",X"04",X"12",
		X"D3",X"12",X"9F",X"13",X"6E",X"14",X"37",X"15",X"03",X"16",X"CB",X"16",X"97",X"17",X"5B",X"18",
		X"26",X"19",X"E6",X"19",X"AF",X"1A",X"6E",X"1B",X"35",X"1C",X"EF",X"1C",X"BB",X"1D",X"6B",X"1E",
		X"46",X"1F",X"82",X"1F",X"D1",X"1D",X"0E",X"1C",X"4E",X"1A",X"90",X"18",X"D6",X"16",X"19",X"15",
		X"64",X"13",X"AA",X"11",X"F8",X"0F",X"44",X"0E",X"9B",X"0C",X"EA",X"0A",X"4A",X"09",X"97",X"07",
		X"00",X"06",X"40",X"04",X"AE",X"02",X"9C",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"1B",X"00",X"A0",X"01",
		X"7E",X"04",X"26",X"08",X"53",X"0C",X"B9",X"10",X"3A",X"15",X"AA",X"19",X"FE",X"1D",X"1A",X"22",
		X"FE",X"25",X"93",X"29",X"E7",X"2C",X"DB",X"2F",X"90",X"32",X"CE",X"34",X"81",X"37",X"37",X"3B",
		X"C8",X"3E",X"52",X"42",X"B6",X"45",X"0C",X"49",X"43",X"4C",X"6A",X"4F",X"6E",X"52",X"68",X"55",
		X"37",X"58",X"08",X"5B",X"1D",X"5D",X"7D",X"5D",X"BF",X"5C",X"3B",X"5B",X"38",X"59",X"E2",X"56",
		X"5D",X"54",X"BD",X"51",X"13",X"4F",X"66",X"4C",X"C0",X"49",X"23",X"47",X"95",X"44",X"13",X"42",
		X"A2",X"3F",X"42",X"3D",X"F4",X"3A",X"B5",X"38",X"89",X"36",X"6A",X"34",X"5F",X"32",X"5F",X"30",
		X"75",X"2E",X"94",X"2C",X"C5",X"2A",X"01",X"29",X"50",X"27",X"B3",X"25",X"66",X"25",X"99",X"26",
		X"AC",X"28",X"61",X"2B",X"6E",X"2E",X"B5",X"31",X"17",X"35",X"83",X"38",X"E9",X"3B",X"46",X"3F",
		X"8F",X"42",X"C4",X"45",X"E1",X"48",X"E6",X"4B",X"D3",X"4E",X"A7",X"51",X"60",X"54",X"01",X"57",
		X"8D",X"59",X"FD",X"5B",X"58",X"5E",X"9A",X"60",X"CA",X"62",X"E1",X"64",X"E8",X"66",X"D1",X"68",
		X"BB",X"6A",X"17",X"6C",X"C6",X"6B",X"45",X"6A",X"F8",X"67",X"2D",X"65",X"0E",X"62",X"C4",X"5E",
		X"61",X"5B",X"F8",X"57",X"91",X"54",X"35",X"51",X"E9",X"4D",X"AE",X"4A",X"88",X"47",X"78",X"44",
		X"7C",X"41",X"97",X"3E",X"C6",X"3B",X"0D",X"39",X"67",X"36",X"D8",X"33",X"5A",X"31",X"F2",X"2E",
		X"99",X"2C",X"59",X"2A",X"25",X"28",X"0A",X"26",X"F8",X"23",X"0E",X"23",X"BE",X"23",X"5C",X"25",
		X"A7",X"27",X"56",X"2A",X"45",X"2D",X"50",X"30",X"71",X"33",X"8D",X"36",X"A2",X"39",X"A5",X"3C",
		X"9C",X"3F",X"7B",X"42",X"45",X"45",X"F6",X"47",X"93",X"4A",X"17",X"4D",X"87",X"4F",X"DE",X"51",
		X"1F",X"54",X"4C",X"56",X"64",X"58",X"68",X"5A",X"58",X"5C",X"32",X"5E",X"FE",X"5F",X"B5",X"61",
		X"5D",X"63",X"F2",X"64",X"78",X"66",X"EA",X"67",X"50",X"69",X"A6",X"6A",X"F0",X"6B",X"2A",X"6D",
		X"56",X"6E",X"76",X"6F",X"86",X"70",X"8D",X"71",X"87",X"72",X"74",X"73",X"59",X"74",X"30",X"75",
		X"FE",X"75",X"C2",X"76",X"7A",X"77",X"2A",X"78",X"CE",X"78",X"6B",X"79",X"00",X"7A",X"8D",X"7A",
		X"10",X"7B",X"8D",X"7B",X"00",X"7C",X"6B",X"7C",X"D1",X"7C",X"2E",X"7D",X"85",X"7D",X"D6",X"7D",
		X"21",X"7E",X"65",X"7E",X"A3",X"7E",X"DD",X"7E",X"0E",X"7F",X"3E",X"7F",X"64",X"7F",X"89",X"7F",
		X"A7",X"7F",X"C0",X"7F",X"D5",X"7F",X"E5",X"7F",X"F2",X"7F",X"F8",X"7F",X"FD",X"7F",X"FD",X"7F",
		X"FA",X"7F",X"F2",X"7F",X"E9",X"7F",X"DA",X"7F",X"C9",X"7F",X"B5",X"7F",X"9C",X"7F",X"82",X"7F",
		X"65",X"7F",X"44",X"7F",X"23",X"7F",X"FB",X"7E",X"D5",X"7E",X"A9",X"7E",X"7E",X"7E",X"4D",X"7E",
		X"1D",X"7E",X"E9",X"7D",X"B6",X"7D",X"7C",X"7D",X"45",X"7D",X"0B",X"7D",X"CF",X"7C",X"8F",X"7C",
		X"52",X"7C",X"0D",X"7C",X"CD",X"7B",X"86",X"7B",X"43",X"7B",X"F8",X"7A",X"B4",X"7A",X"66",X"7A",
		X"22",X"7A",X"CD",X"79",X"91",X"79",X"91",X"78",X"F7",X"75",X"59",X"72",X"0C",X"6E",X"5D",X"69",
		X"70",X"64",X"6D",X"5F",X"62",X"5A",X"61",X"55",X"71",X"50",X"9C",X"4B",X"E2",X"46",X"49",X"42",
		X"CE",X"3D",X"74",X"39",X"3E",X"35",X"25",X"31",X"2C",X"2D",X"56",X"29",X"9C",X"25",X"01",X"22",
		X"84",X"1E",X"23",X"1B",X"DE",X"17",X"B4",X"14",X"A3",X"11",X"AD",X"0E",X"E1",X"0B",X"84",X"0A",
		X"A7",X"0A",X"AE",X"0B",X"5B",X"0D",X"6A",X"0F",X"B9",X"11",X"28",X"14",X"AB",X"16",X"2F",X"19",
		X"B1",X"1B",X"2A",X"1E",X"95",X"20",X"EF",X"22",X"38",X"25",X"72",X"27",X"98",X"29",X"AB",X"2B",
		X"AC",X"2D",X"9E",X"2F",X"79",X"31",X"47",X"33",X"00",X"35",X"AF",X"36",X"47",X"38",X"D8",X"39",
		X"4C",X"3B",X"C9",X"3C",X"A6",X"3D",X"D9",X"3C",X"EC",X"3A",X"3B",X"38",X"12",X"35",X"9E",X"31",
		X"02",X"2E",X"54",X"2A",X"A3",X"26",X"FB",X"22",X"60",X"1F",X"D7",X"1B",X"64",X"18",X"09",X"15",
		X"C7",X"11",X"9C",X"0E",X"8C",X"0B",X"93",X"08",X"B1",X"05",X"E8",X"02",X"36",X"00",X"9B",X"FD",
		X"14",X"FB",X"A6",X"F8",X"45",X"F6",X"05",X"F4",X"C3",X"F1",X"03",X"F0",X"EC",X"EF",X"0D",X"F1",
		X"FB",X"F2",X"6D",X"F5",X"32",X"F8",X"24",X"FB",X"2E",X"FE",X"40",X"01",X"51",X"04",X"55",X"07",
		X"4D",X"0A",X"30",X"0D",X"02",X"10",X"BD",X"12",X"63",X"15",X"F4",X"17",X"70",X"1A",X"D4",X"1C",
		X"24",X"1F",X"60",X"21",X"87",X"23",X"9D",X"25",X"9E",X"27",X"8F",X"29",X"6C",X"2B",X"37",X"2D",
		X"F3",X"2E",X"9E",X"30",X"38",X"32",X"C4",X"33",X"40",X"35",X"AD",X"36",X"0E",X"38",X"62",X"39",
		X"A7",X"3A",X"DF",X"3B",X"0D",X"3D",X"2C",X"3E",X"42",X"3F",X"4B",X"40",X"49",X"41",X"3E",X"42",
		X"28",X"43",X"07",X"44",X"DD",X"44",X"AB",X"45",X"6D",X"46",X"29",X"47",X"DC",X"47",X"86",X"48",
		X"28",X"49",X"C3",X"49",X"56",X"4A",X"E0",X"4A",X"66",X"4B",X"E3",X"4B",X"5B",X"4C",X"CC",X"4C",
		X"37",X"4D",X"9B",X"4D",X"FA",X"4D",X"54",X"4E",X"A6",X"4E",X"F6",X"4E",X"3E",X"4F",X"84",X"4F",
		X"C2",X"4F",X"FE",X"4F",X"33",X"50",X"68",X"50",X"95",X"50",X"BF",X"50",X"E6",X"50",X"08",X"51",
		X"24",X"51",X"41",X"51",X"55",X"51",X"6D",X"51",X"7A",X"51",X"8F",X"51",X"90",X"51",X"A6",X"51",
		X"DA",X"50",X"71",X"4E",X"13",X"4B",X"09",X"47",X"A1",X"42",X"FB",X"3D",X"3F",X"39",X"7B",X"34",
		X"C4",X"2F",X"1B",X"2B",X"8A",X"26",X"15",X"22",X"BF",X"1D",X"87",X"19",X"70",X"15",X"76",X"11",
		X"9E",X"0D",X"E5",X"09",X"4B",X"06",X"CC",X"02",X"6E",X"FF",X"29",X"FC",X"01",X"F9",X"F4",X"F5",
		X"00",X"F3",X"25",X"F0",X"62",X"ED",X"D8",X"EA",X"D4",X"E9",X"3C",X"EA",X"84",X"EB",X"68",X"ED",
		X"AC",X"EF",X"2B",X"F2",X"C9",X"F4",X"77",X"F7",X"28",X"FA",X"D5",X"FC",X"74",X"FF",X"07",X"02",
		X"8A",X"04",X"FA",X"06",X"58",X"09",X"A3",X"0B",X"DD",X"0D",X"02",X"10",X"17",X"12",X"17",X"14",
		X"06",X"16",X"E5",X"17",X"B5",X"19",X"6E",X"1B",X"20",X"1D",X"B6",X"1E",X"54",X"20",X"35",X"21",
		X"68",X"20",X"89",X"1E",X"E9",X"1B",X"D9",X"18",X"81",X"15",X"02",X"12",X"72",X"0E",X"E1",X"0A",
		X"55",X"07",X"DC",X"03",X"74",X"00",X"21",X"FD",X"E5",X"F9",X"C2",X"F6",X"B5",X"F3",X"C3",X"F0",
		X"E8",X"ED",X"24",X"EB",X"79",X"E8",X"E5",X"E5",X"65",X"E3",X"FD",X"E0",X"A6",X"DE",X"6B",X"DC",
		X"3C",X"DA",X"25",X"D8",X"2A",X"D6",X"90",X"D5",X"73",X"D6",X"3A",X"D8",X"A6",X"DA",X"6D",X"DD",
		X"74",X"E0",X"95",X"E3",X"C6",X"E6",X"F6",X"E9",X"1F",X"ED",X"39",X"F0",X"42",X"F3",X"37",X"F6",
		X"18",X"F9",X"E4",X"FB",X"99",X"FE",X"36",X"01",X"BF",X"03",X"34",X"06",X"91",X"08",X"DD",X"0A",
		X"11",X"0D",X"35",X"0F",X"43",X"11",X"44",X"13",X"2A",X"15",X"11",X"17",X"68",X"18",X"11",X"18",
		X"90",X"16",X"46",X"14",X"82",X"11",X"6C",X"0E",X"2E",X"0B",X"D8",X"07",X"7F",X"04",X"2A",X"01",
		X"E4",X"FD",X"AA",X"FA",X"87",X"F7",X"78",X"F4",X"80",X"F1",X"A0",X"EE",X"D5",X"EB",X"21",X"E9",
		X"85",X"E6",X"FF",X"E3",X"8E",X"E1",X"33",X"DF",X"EB",X"DC",X"B8",X"DA",X"99",X"D8",X"8C",X"D6",
		X"92",X"D4",X"AA",X"D2",X"D1",X"D0",X"0A",X"CF",X"55",X"CD",X"AE",X"CB",X"15",X"CA",X"8D",X"C8",
		X"13",X"C7",X"A6",X"C5",X"48",X"C4",X"F6",X"C2",X"B1",X"C1",X"79",X"C0",X"4B",X"BF",X"2B",X"BE",
		X"15",X"BD",X"0A",X"BC",X"09",X"BB",X"13",X"BA",X"26",X"B9",X"45",X"B8",X"69",X"B7",X"99",X"B6",
		X"D2",X"B5",X"11",X"B5",X"5B",X"B4",X"AC",X"B3",X"05",X"B3",X"65",X"B2",X"CC",X"B1",X"3A",X"B1",
		X"AF",X"B0",X"2B",X"B0",X"AD",X"AF",X"35",X"AF",X"C3",X"AE",X"58",X"AE",X"F1",X"AD",X"91",X"AD",
		X"34",X"AD",X"DE",X"AC",X"8B",X"AC",X"40",X"AC",X"F7",X"AB",X"B4",X"AB",X"74",X"AB",X"39",X"AB",
		X"03",X"AB",X"CF",X"AA",X"A1",X"AA",X"73",X"AA",X"4C",X"AA",X"27",X"AA",X"06",X"AA",X"E9",X"A9",
		X"CF",X"A9",X"B6",X"A9",X"A3",X"A9",X"91",X"A9",X"82",X"A9",X"76",X"A9",X"6D",X"A9",X"64",X"A9",
		X"5F",X"A9",X"5C",X"A9",X"5D",X"A9",X"5F",X"A9",X"64",X"A9",X"69",X"A9",X"72",X"A9",X"7C",X"A9",
		X"89",X"A9",X"96",X"A9",X"A5",X"A9",X"B5",X"A9",X"C8",X"A9",X"DC",X"A9",X"F3",X"A9",X"0A",X"AA",
		X"24",X"AA",X"3D",X"AA",X"5A",X"AA",X"71",X"AA",X"BD",X"AA",X"86",X"AC",X"99",X"AF",X"76",X"B3",
		X"D5",X"B7",X"7D",X"BC",X"4B",X"C1",X"26",X"C6",X"FE",X"CA",X"C8",X"CF",X"7A",X"D4",X"12",X"D9",
		X"8C",X"DD",X"E5",X"E1",X"1F",X"E6",X"36",X"EA",X"2F",X"EE",X"06",X"F2",X"BE",X"F5",X"58",X"F9",
		X"D1",X"FC",X"2F",X"00",X"6D",X"03",X"94",X"06",X"98",X"09",X"8D",X"0C",X"59",X"0F",X"24",X"12",
		X"11",X"14",X"49",X"14",X"6F",X"13",X"D0",X"11",X"BC",X"0F",X"57",X"0D",X"CA",X"0A",X"22",X"08",
		X"73",X"05",X"C2",X"02",X"1D",X"00",X"82",X"FD",X"F6",X"FA",X"7C",X"F8",X"12",X"F6",X"BC",X"F3",
		X"77",X"F1",X"44",X"EF",X"23",X"ED",X"17",X"EB",X"1A",X"E9",X"2F",X"E7",X"54",X"E5",X"8A",X"E3",
		X"D0",X"E1",X"24",X"E0",X"88",X"DE",X"FA",X"DC",X"7A",X"DB",X"07",X"DA",X"A2",X"D8",X"4A",X"D7",
		X"FF",X"D5",X"C0",X"D4",X"89",X"D3",X"62",X"D2",X"44",X"D1",X"31",X"D0",X"27",X"CF",X"2B",X"CE",
		X"34",X"CD",X"4A",X"CC",X"66",X"CB",X"8C",X"CA",X"BA",X"C9",X"F2",X"C8",X"30",X"C8",X"78",X"C7",
		X"C5",X"C6",X"1E",X"C6",X"77",X"C5",X"DF",X"C4",X"45",X"C4",X"BC",X"C3",X"24",X"C3",X"2C",X"C3",
		X"D7",X"C4",X"97",X"C7",X"13",X"CB",X"FD",X"CE",X"2A",X"D3",X"77",X"D7",X"D1",X"DB",X"27",X"E0",
		X"6E",X"E4",X"A1",X"E8",X"BB",X"EC",X"BB",X"F0",X"9E",X"F4",X"63",X"F8",X"09",X"FC",X"93",X"FF",
		X"FD",X"02",X"4E",X"06",X"81",X"09",X"99",X"0C",X"98",X"0F",X"7A",X"12",X"46",X"15",X"F5",X"17",
		X"91",X"1A",X"11",X"1D",X"79",X"1F",X"94",X"20",X"20",X"20",X"C0",X"1E",X"B4",X"1C",X"46",X"1A",
		X"93",X"17",X"C3",X"14",X"DA",X"11",X"F5",X"0E",X"10",X"0C",X"3A",X"09",X"6E",X"06",X"B7",X"03",
		X"10",X"01",X"7E",X"FE",X"00",X"FC",X"96",X"F9",X"3D",X"F7",X"FA",X"F4",X"C7",X"F2",X"AC",X"F0",
		X"9D",X"EE",X"A4",X"EC",X"B8",X"EA",X"DF",X"E8",X"17",X"E7",X"5E",X"E5",X"B3",X"E3",X"19",X"E2",
		X"8B",X"E0",X"0D",X"DF",X"9C",X"DD",X"39",X"DC",X"E1",X"DA",X"95",X"D9",X"55",X"D8",X"23",X"D7",
		X"F8",X"D5",X"DE",X"D4",X"C9",X"D3",X"C0",X"D2",X"C1",X"D1",X"CD",X"D0",X"E0",X"CF",X"FE",X"CE",
		X"23",X"CE",X"53",X"CD",X"89",X"CC",X"C6",X"CB",X"0E",X"CB",X"5C",X"CA",X"AF",X"C9",X"0C",X"C9",
		X"70",X"C8",X"D7",X"C7",X"49",X"C7",X"BF",X"C6",X"3A",X"C6",X"BB",X"C5",X"43",X"C5",X"D2",X"C4",
		X"63",X"C4",X"FB",X"C3",X"98",X"C3",X"38",X"C3",X"E2",X"C2",X"8C",X"C2",X"3A",X"C2",X"ED",X"C1",
		X"A5",X"C1",X"5F",X"C1",X"1F",X"C1",X"E2",X"C0",X"AA",X"C0",X"73",X"C0",X"41",X"C0",X"11",X"C0",
		X"E7",X"BF",X"BD",X"BF",X"99",X"BF",X"75",X"BF",X"54",X"BF",X"38",X"BF",X"1C",X"BF",X"04",X"BF",
		X"EE",X"BE",X"DA",X"BE",X"CA",X"BE",X"BB",X"BE",X"AF",X"BE",X"A4",X"BE",X"9C",X"BE",X"97",X"BE",
		X"91",X"BE",X"8B",X"BE",X"8C",X"BE",X"8D",X"BE",X"91",X"BE",X"94",X"BE",X"99",X"BE",X"A1",X"BE",
		X"AA",X"BE",X"B2",X"BE",X"BE",X"BE",X"CA",X"BE",X"D7",X"BE",X"E7",X"BE",X"F9",X"BE",X"05",X"BF",
		X"3E",X"BF",X"E9",X"C0",X"E7",X"C3",X"B0",X"C7",X"01",X"CC",X"9A",X"D0",X"5D",X"D5",X"2A",X"DA",
		X"F8",X"DE",X"B5",X"E3",X"5C",X"E8",X"E8",X"EC",X"58",X"F1",X"A5",X"F5",X"D4",X"F9",X"E1",X"FD",
		X"CD",X"01",X"97",X"05",X"45",X"09",X"D3",X"0C",X"41",X"10",X"93",X"13",X"C6",X"16",X"DD",X"19",
		X"DC",X"1C",X"BE",X"1F",X"88",X"22",X"37",X"25",X"CF",X"27",X"51",X"2A",X"BA",X"2C",X"0E",X"2F",
		X"4D",X"31",X"77",X"33",X"8D",X"35",X"91",X"37",X"7E",X"39",X"5D",X"3B",X"28",X"3D",X"E2",X"3E",
		X"8C",X"40",X"26",X"42",X"AE",X"43",X"2A",X"45",X"95",X"46",X"F2",X"47",X"43",X"49",X"86",X"4A",
		X"BB",X"4B",X"E4",X"4C",X"FF",X"4D",X"11",X"4F",X"13",X"50",X"11",X"51",X"FE",X"51",X"D4",X"52",
		X"4C",X"52",X"53",X"50",X"7E",X"4D",X"0E",X"4A",X"49",X"46",X"4F",X"42",X"3F",X"3E",X"27",X"3A",
		X"16",X"36",X"15",X"32",X"26",X"2E",X"4E",X"2A",X"91",X"26",X"EC",X"22",X"62",X"1F",X"F7",X"1B",
		X"A3",X"18",X"6D",X"15",X"4D",X"12",X"4A",X"0F",X"5D",X"0C",X"8A",X"09",X"CD",X"06",X"2C",X"04",
		X"98",X"01",X"25",X"FF",X"B3",X"FC",X"E0",X"FA",X"BE",X"FA",X"C3",X"FB",X"95",X"FD",X"E2",X"FF",
		X"83",X"02",X"4E",X"05",X"33",X"08",X"21",X"0B",X"09",X"0E",X"E9",X"10",X"BC",X"13",X"7C",X"16",
		X"2A",X"19",X"C3",X"1B",X"49",X"1E",X"B7",X"20",X"15",X"23",X"5A",X"25",X"8D",X"27",X"AB",X"29",
		X"B9",X"2B",X"B1",X"2D",X"9B",X"2F",X"6E",X"31",X"34",X"33",X"E4",X"34",X"86",X"36",X"F1",X"36",
		X"CB",X"35",X"BB",X"33",X"01",X"31",X"E9",X"2D",X"91",X"2A",X"1D",X"27",X"9B",X"23",X"1A",X"20",
		X"A1",X"1C",X"3B",X"19",X"E3",X"15",X"A4",X"12",X"78",X"0F",X"67",X"0C",X"6B",X"09",X"89",X"06",
		X"BC",X"03",X"06",X"01",X"69",X"FE",X"E1",X"FB",X"6D",X"F9",X"0E",X"F7",X"C4",X"F4",X"8E",X"F2",
		X"69",X"F0",X"57",X"EE",X"57",X"EC",X"6A",X"EA",X"8D",X"E8",X"C0",X"E6",X"04",X"E5",X"56",X"E3",
		X"B7",X"E1",X"27",X"E0",X"A5",X"DE",X"31",X"DD",X"CA",X"DB",X"70",X"DA",X"21",X"D9",X"DF",X"D7",
		X"AA",X"D6",X"7F",X"D5",X"5E",X"D4",X"4A",X"D3",X"40",X"D2",X"3F",X"D1",X"47",X"D0",X"5B",X"CF",
		X"75",X"CE",X"99",X"CD",X"C7",X"CC",X"FC",X"CB",X"37",X"CB",X"7E",X"CA",X"CA",X"C9",X"1E",X"C9",
		X"79",X"C8",X"DA",X"C7",X"44",X"C7",X"B3",X"C6",X"28",X"C6",X"A5",X"C5",X"24",X"C5",X"AC",X"C4",
		X"38",X"C4",X"CB",X"C3",X"61",X"C3",X"FE",X"C2",X"9E",X"C2",X"45",X"C2",X"EF",X"C1",X"9D",X"C1",
		X"50",X"C1",X"08",X"C1",X"C3",X"C0",X"82",X"C0",X"45",X"C0",X"0C",X"C0",X"D6",X"BF",X"A4",X"BF",
		X"6F",X"BF",X"78",X"BF",X"02",X"C1",X"D5",X"C3",X"70",X"C7",X"8F",X"CB",X"F9",X"CF",X"8A",X"D4",
		X"26",X"D9",X"C4",X"DD",X"51",X"E2",X"CA",X"E6",X"2A",X"EB",X"6E",X"EF",X"93",X"F3",X"99",X"F7",
		X"7F",X"FB",X"45",X"FF",X"ED",X"02",X"75",X"06",X"DF",X"09",X"2D",X"0D",X"60",X"10",X"73",X"13",
		X"72",X"16",X"4E",X"19",X"1C",X"1C",X"C3",X"1E",X"68",X"21",X"28",X"23",X"32",X"23",X"32",X"22",
		X"6E",X"20",X"37",X"1E",X"B1",X"1B",X"03",X"19",X"3B",X"16",X"70",X"13",X"A2",X"10",X"DF",X"0D",
		X"27",X"0B",X"82",X"08",X"EA",X"05",X"69",X"03",X"F7",X"00",X"9B",X"FE",X"51",X"FC",X"1B",X"FA",
		X"F6",X"F7",X"E3",X"F5",X"E1",X"F3",X"F1",X"F1",X"10",X"F0",X"3F",X"EE",X"81",X"EC",X"D1",X"EA",
		X"2F",X"E9",X"9C",X"E7",X"17",X"E6",X"9F",X"E4",X"34",X"E3",X"D6",X"E1",X"86",X"E0",X"40",X"DF",
		X"07",X"DE",X"D7",X"DC",X"B5",X"DB",X"9B",X"DA",X"8C",X"D9",X"87",X"D8",X"8E",X"D7",X"9B",X"D6",
		X"B3",X"D5",X"D2",X"D4",X"FD",X"D3",X"2B",X"D3",X"65",X"D2",X"A4",X"D1",X"F0",X"D0",X"3C",X"D0",
		X"97",X"CF",X"EF",X"CE",X"5B",X"CE",X"B7",X"CD",X"BA",X"CD",X"60",X"CF",X"19",X"D2",X"8C",X"D5",
		X"6B",X"D9",X"90",X"DD",X"D1",X"E1",X"21",X"E6",X"68",X"EA",X"A6",X"EE",X"CC",X"F2",X"DC",X"F6",
		X"D0",X"FA",X"A8",X"FE",X"5F",X"02",X"FB",X"05",X"7B",X"09",X"DE",X"0C",X"22",X"10",X"4C",X"13",
		X"5B",X"16",X"4C",X"19",X"26",X"1C",X"E7",X"1E",X"8F",X"21",X"1F",X"24",X"98",X"26",X"FB",X"28",
		X"47",X"2B",X"7F",X"2D",X"A4",X"2F",X"B4",X"31",X"B2",X"33",X"9B",X"35",X"74",X"37",X"3A",X"39",
		X"F0",X"3A",X"95",X"3C",X"2C",X"3E",X"B1",X"3F",X"29",X"41",X"90",X"42",X"EC",X"43",X"3A",X"45",
		X"79",X"46",X"AB",X"47",X"D3",X"48",X"EE",X"49",X"FD",X"4A",X"00",X"4C",X"F8",X"4C",X"E6",X"4D",
		X"CB",X"4E",X"A5",X"4F",X"76",X"50",X"3B",X"51",X"FA",X"51",X"AF",X"52",X"5A",X"53",X"FE",X"53",
		X"9B",X"54",X"2F",X"55",X"BC",X"55",X"41",X"56",X"BF",X"56",X"39",X"57",X"A9",X"57",X"15",X"58",
		X"78",X"58",X"D7",X"58",X"30",X"59",X"83",X"59",X"D0",X"59",X"17",X"5A",X"5C",X"5A",X"99",X"5A",
		X"D3",X"5A",X"08",X"5B",X"37",X"5B",X"65",X"5B",X"8D",X"5B",X"AE",X"5B",X"D1",X"5B",X"EB",X"5B",
		X"04",X"5C",X"18",X"5C",X"2A",X"5C",X"38",X"5C",X"43",X"5C",X"49",X"5C",X"4F",X"5C",X"4F",X"5C",
		X"4F",X"5C",X"49",X"5C",X"44",X"5C",X"39",X"5C",X"2E",X"5C",X"20",X"5C",X"10",X"5C",X"FC",X"5B",
		X"E7",X"5B",X"CF",X"5B",X"B7",X"5B",X"9D",X"5B",X"80",X"5B",X"61",X"5B",X"41",X"5B",X"1E",X"5B",
		X"FC",X"5A",X"D6",X"5A",X"AF",X"5A",X"87",X"5A",X"5D",X"5A",X"32",X"5A",X"07",X"5A",X"D8",X"59",
		X"A9",X"59",X"78",X"59",X"48",X"59",X"15",X"59",X"E4",X"58",X"AE",X"58",X"79",X"58",X"43",X"58",
		X"0C",X"58",X"D3",X"57",X"9C",X"57",X"62",X"57",X"28",X"57",X"EC",X"56",X"B1",X"56",X"74",X"56",
		X"38",X"56",X"FA",X"55",X"BD",X"55",X"7B",X"55",X"40",X"55",X"D6",X"54",X"F5",X"52",X"C2",X"4F",
		X"CB",X"4B",X"4E",X"47",X"8A",X"42",X"9C",X"3D",X"A4",X"38",X"AD",X"33",X"C9",X"2E",X"F9",X"29",
		X"46",X"25",X"B0",X"20",X"3C",X"1C",X"E6",X"17",X"B5",X"13",X"A3",X"0F",X"B3",X"0B",X"E0",X"07",
		X"31",X"04",X"9D",X"00",X"2A",X"FD",X"D1",X"F9",X"97",X"F6",X"78",X"F3",X"74",X"F0",X"89",X"ED",
		X"B6",X"EA",X"FB",X"E7",X"5C",X"E5",X"CF",X"E2",X"5C",X"E0",X"FD",X"DD",X"B3",X"DB",X"7D",X"D9",
		X"5B",X"D7",X"4D",X"D5",X"52",X"D3",X"66",X"D1",X"8E",X"CF",X"C6",X"CD",X"0D",X"CC",X"67",X"CA",
		X"CE",X"C8",X"44",X"C7",X"CB",X"C5",X"5E",X"C4",X"FE",X"C2",X"AC",X"C1",X"67",X"C0",X"2E",X"BF",
		X"01",X"BE",X"E2",X"BC",X"C8",X"BB",X"BF",X"BA",X"D1",X"B9",X"45",X"BA",X"2B",X"BC",X"E8",X"BE",
		X"40",X"C2",X"EB",X"C5",X"CD",X"C9",X"C1",X"CD",X"C0",X"D1",X"B5",X"D5",X"9E",X"D9",X"71",X"DD",
		X"30",X"E1",X"D3",X"E4",X"5D",X"E8",X"CB",X"EB",X"1F",X"EF",X"57",X"F2",X"77",X"F5",X"7B",X"F8",
		X"67",X"FB",X"38",X"FE",X"F1",X"00",X"94",X"03",X"22",X"06",X"96",X"08",X"FA",X"0A",X"43",X"0D",
		X"7C",X"0F",X"A0",X"11",X"B2",X"13",X"AF",X"15",X"9D",X"17",X"78",X"19",X"44",X"1B",X"FD",X"1C",
		X"A9",X"1E",X"43",X"20",X"CF",X"21",X"4E",X"23",X"BE",X"24",X"21",X"26",X"76",X"27",X"BE",X"28",
		X"FA",X"29",X"2A",X"2B",X"4E",X"2C",X"68",X"2D",X"77",X"2E",X"7C",X"2F",X"75",X"30",X"67",X"31",
		X"4B",X"32",X"2A",X"33",X"FA",X"33",X"C3",X"34",X"52",X"34",X"5C",X"32",X"86",X"2F",X"0C",X"2C",
		X"3E",X"28",X"34",X"24",X"16",X"20",X"ED",X"1B",X"D0",X"17",X"BE",X"13",X"C3",X"0F",X"DD",X"0B",
		X"16",X"08",X"65",X"04",X"D5",X"00",X"5F",X"FD",X"06",X"FA",X"C7",X"F6",X"A4",X"F3",X"9A",X"F0",
		X"AB",X"ED",X"D6",X"EA",X"17",X"E8",X"71",X"E5",X"E3",X"E2",X"6A",X"E0",X"07",X"DE",X"B9",X"DB",
		X"7F",X"D9",X"5B",X"D7",X"47",X"D5",X"49",X"D3",X"5B",X"D1",X"7F",X"CF",X"B4",X"CD",X"FB",X"CB",
		X"4F",X"CA",X"B4",X"C8",X"29",X"C7",X"AB",X"C5",X"3A",X"C4",X"DB",X"C2",X"86",X"C1",X"3F",X"C0",
		X"02",X"BF",X"D6",X"BD",X"B1",X"BC",X"9B",X"BB",X"8D",X"BA",X"8D",X"B9",X"91",X"B8",X"AA",X"B7",
		X"C0",X"B6",X"EC",X"B5",X"11",X"B5",X"48",X"B5",X"13",X"B7",X"CD",X"B9",X"32",X"BD",X"F5",X"C0",
		X"F7",X"C4",X"0F",X"C9",X"33",X"CD",X"51",X"D1",X"65",X"D5",X"5F",X"D9",X"44",X"DD",X"11",X"E1",
		X"C0",X"E4",X"56",X"E8",X"CE",X"EB",X"2C",X"EF",X"6E",X"F2",X"94",X"F5",X"9E",X"F8",X"91",X"FB",
		X"6B",X"FE",X"2D",X"01",X"D5",X"03",X"6A",X"06",X"E2",X"08",X"50",X"0B",X"69",X"0D",X"E9",X"0D",
		X"14",X"0D",X"69",X"0B",X"2B",X"09",X"95",X"06",X"CB",X"03",X"E3",X"00",X"F3",X"FD",X"00",X"FB",
		X"15",X"F8",X"38",X"F5",X"6A",X"F2",X"B1",X"EF",X"09",X"ED",X"77",X"EA",X"F7",X"E7",X"8E",X"E5",
		X"38",X"E3",X"F9",X"E0",X"CA",X"DE",X"AE",X"DC",X"A6",X"DA",X"B0",X"D8",X"C9",X"D6",X"F5",X"D4",
		X"33",X"D3",X"7F",X"D1",X"DB",X"CF",X"47",X"CE",X"C0",X"CC",X"4A",X"CB",X"E0",X"C9",X"83",X"C8",
		X"33",X"C7",X"F3",X"C5",X"BB",X"C4",X"90",X"C3",X"70",X"C2",X"5C",X"C1",X"53",X"C0",X"55",X"BF",
		X"5F",X"BE",X"74",X"BD",X"90",X"BC",X"BB",X"BB",X"E9",X"BA",X"24",X"BA",X"66",X"B9",X"AF",X"B8",
		X"00",X"B8",X"5C",X"B7",X"BB",X"B6",X"23",X"B6",X"91",X"B5",X"09",X"B5",X"83",X"B4",X"07",X"B4",
		X"8E",X"B3",X"1F",X"B3",X"B0",X"B2",X"4B",X"B2",X"E9",X"B1",X"8F",X"B1",X"37",X"B1",X"E8",X"B0",
		X"9B",X"B0",X"53",X"B0",X"0D",X"B0",X"CF",X"AF",X"93",X"AF",X"5D",X"AF",X"28",X"AF",X"FC",X"AE",
		X"CE",X"AE",X"A8",X"AE",X"81",X"AE",X"62",X"AE",X"40",X"AE",X"2A",X"AE",X"0D",X"AE",X"FF",X"AD",
		X"DE",X"AD",X"68",X"AE",X"93",X"B0",X"C9",X"B3",X"B5",X"B7",X"09",X"BC",X"9E",X"C0",X"4C",X"C5",
		X"06",X"CA",X"B5",X"CE",X"57",X"D3",X"DE",X"D7",X"4B",X"DC",X"9B",X"E0",X"CE",X"E4",X"DC",X"E8",
		X"CF",X"EC",X"A1",X"F0",X"55",X"F4",X"E7",X"F7",X"5E",X"FB",X"B5",X"FE",X"F3",X"01",X"14",X"05",
		X"1A",X"08",X"05",X"0B",X"D8",X"0D",X"90",X"10",X"27",X"13",X"64",X"14",X"16",X"14",X"E1",X"12",
		X"FF",X"10",X"BD",X"0E",X"38",X"0C",X"93",X"09",X"D7",X"06",X"1C",X"04",X"62",X"01",X"B6",X"FE",
		X"14",X"FC",X"83",X"F9",X"03",X"F7",X"99",X"F4",X"3E",X"F2",X"F7",X"EF",X"C3",X"ED",X"A2",X"EB",
		X"91",X"E9",X"93",X"E7",X"A4",X"E5",X"CB",X"E3",X"FF",X"E1",X"43",X"E0",X"98",X"DE",X"FC",X"DC",
		X"6C",X"DB",X"EE",X"D9",X"7A",X"D8",X"15",X"D7",X"BD",X"D5",X"71",X"D4",X"32",X"D3",X"FF",X"D1",
		X"D7",X"D0",X"B8",X"CF",X"A6",X"CE",X"9E",X"CD",X"A0",X"CC",X"AC",X"CB",X"C1",X"CA",X"E0",X"C9",
		X"07",X"C9",X"37",X"C8",X"70",X"C7",X"AF",X"C6",X"F7",X"C5",X"46",X"C5",X"9E",X"C4",X"FD",X"C3",
		X"61",X"C3",X"CD",X"C2",X"41",X"C2",X"B9",X"C1",X"39",X"C1",X"BE",X"C0",X"48",X"C0",X"D9",X"BF",
		X"6F",X"BF",X"09",X"BF",X"AA",X"BE",X"4E",X"BE",X"F8",X"BD",X"A6",X"BD",X"58",X"BD",X"0E",X"BD",
		X"CA",X"BC",X"88",X"BC",X"4D",X"BC",X"14",X"BC",X"DE",X"BB",X"AC",X"BB",X"7E",X"BB",X"53",X"BB",
		X"2B",X"BB",X"05",X"BB",X"E3",X"BA",X"C5",X"BA",X"AB",X"BA",X"91",X"BA",X"7A",X"BA",X"67",X"BA",
		X"55",X"BA",X"47",X"BA",X"3A",X"BA",X"2F",X"BA",X"27",X"BA",X"22",X"BA",X"1D",X"BA",X"1C",X"BA",
		X"1B",X"BA",X"1E",X"BA",X"22",X"BA",X"27",X"BA",X"2D",X"BA",X"35",X"BA",X"3F",X"BA",X"4C",X"BA",
		X"58",X"BA",X"68",X"BA",X"76",X"BA",X"8A",X"BA",X"9A",X"BA",X"B0",X"BA",X"C2",X"BA",X"DC",X"BA",
		X"EF",X"BA",X"0E",X"BB",X"1B",X"BB",X"19",X"BC",X"AB",X"BE",X"2C",X"C2",X"58",X"C6",X"DB",X"CA",
		X"99",X"CF",X"69",X"D4",X"41",X"D9",X"0C",X"DE",X"C2",X"E2",X"62",X"E7",X"E4",X"EB",X"46",X"F0",
		X"87",X"F4",X"A8",X"F8",X"A9",X"FC",X"89",X"00",X"47",X"04",X"E9",X"07",X"68",X"0B",X"CE",X"0E",
		X"11",X"12",X"3D",X"15",X"47",X"18",X"40",X"1B",X"11",X"1E",X"E0",X"20",X"CE",X"22",X"08",X"23",
		X"2E",X"22",X"92",X"20",X"80",X"1E",X"1D",X"1C",X"90",X"19",X"EA",X"16",X"39",X"14",X"89",X"11",
		X"E4",X"0E",X"48",X"0C",X"BC",X"09",X"3F",X"07",X"D5",X"04",X"7C",X"02",X"37",X"00",X"05",X"FE",
		X"E2",X"FB",X"D2",X"F9",X"D3",X"F7",X"E7",X"F5",X"07",X"F4",X"39",X"F2",X"7C",X"F0",X"CD",X"EE",
		X"2C",X"ED",X"B3",X"EB",X"A3",X"EB",X"02",X"ED",X"3E",X"EF",X"13",X"F2",X"3F",X"F5",X"A3",X"F8",
		X"1E",X"FC",X"A4",X"FF",X"26",X"03",X"9B",X"06",X"FE",X"09",X"4F",X"0D",X"88",X"10",X"AA",X"13",
		X"B0",X"16",X"A2",X"19",X"78",X"1C",X"38",X"1F",X"DF",X"21",X"70",X"24",X"E9",X"26",X"4C",X"29",
		X"9A",X"2B",X"D4",X"2D",X"F7",X"2F",X"09",X"32",X"07",X"34",X"F3",X"35",X"CB",X"37",X"94",X"39",
		X"4A",X"3B",X"F2",X"3C",X"87",X"3E",X"10",X"40",X"87",X"41",X"F1",X"42",X"4D",X"44",X"9A",X"45",
		X"DD",X"46",X"0F",X"48",X"38",X"49",X"53",X"4A",X"63",X"4B",X"67",X"4C",X"60",X"4D",X"50",X"4E",
		X"36",X"4F",X"0F",X"50",X"E2",X"50",X"A7",X"51",X"68",X"52",X"1B",X"53",X"CC",X"53",X"6E",X"54",
		X"07",X"55",X"5F",X"54",X"36",X"52",X"30",X"4F",X"8B",X"4B",X"8E",X"47",X"5B",X"43",X"13",X"3F",
		X"C3",X"3A",X"7D",X"36",X"45",X"32",X"23",X"2E",X"1A",X"2A",X"2C",X"26",X"58",X"22",X"A3",X"1E",
		X"0A",X"1B",X"8B",X"17",X"2B",X"14",X"E4",X"10",X"BD",X"0D",X"A9",X"0A",X"B6",X"07",X"D5",X"04",
		X"12",X"02",X"60",X"FF",X"CE",X"FC",X"3F",X"FA",X"34",X"F8",X"D7",X"F7",X"B2",X"F8",X"5D",X"FA",
		X"8C",X"FC",X"11",X"FF",X"C4",X"01",X"94",X"04",X"6D",X"07",X"43",X"0A",X"13",X"0D",X"D5",X"0F",
		X"88",X"12",X"27",X"15",X"B2",X"17",X"2A",X"1A",X"8F",X"1C",X"DD",X"1E",X"1A",X"21",X"42",X"23",
		X"57",X"25",X"59",X"27",X"4B",X"29",X"28",X"2B",X"F8",X"2C",X"B2",X"2E",X"5F",X"30",X"FB",X"31",
		X"89",X"33",X"07",X"35",X"78",X"36",X"DA",X"37",X"2E",X"39",X"76",X"3A",X"B1",X"3B",X"DE",X"3C",
		X"03",X"3E",X"18",X"3F",X"24",X"40",X"24",X"41",X"1B",X"42",X"07",X"43",X"EA",X"43",X"C2",X"44",
		X"91",X"45",X"57",X"46",X"16",X"47",X"CA",X"47",X"78",X"48",X"1B",X"49",X"BA",X"49",X"4E",X"4A",
		X"DD",X"4A",X"62",X"4B",X"EB",X"4B",X"28",X"4C",X"D5",X"4A",X"3F",X"48",X"E2",X"44",X"01",X"41",
		X"D5",X"3C",X"7F",X"38",X"1B",X"34",X"B5",X"2F",X"5C",X"2B",X"16",X"27",X"E7",X"22",X"D2",X"1E",
		X"DB",X"1A",X"FE",X"16",X"40",X"13",X"A0",X"0F",X"1C",X"0C",X"B7",X"08",X"6C",X"05",X"3D",X"02",
		X"27",X"FF",X"2E",X"FC",X"4B",X"F9",X"85",X"F6",X"D0",X"F3",X"3C",X"F1",X"AB",X"EE",X"11",X"ED",
		X"23",X"ED",X"3D",X"EE",X"15",X"F0",X"5A",X"F2",X"EE",X"F4",X"A5",X"F7",X"77",X"FA",X"4A",X"FD",
		X"1E",X"00",X"E3",X"02",X"9E",X"05",X"47",X"08",X"DF",X"0A",X"63",X"0D",X"D4",X"0F",X"2F",X"12",
		X"7A",X"14",X"AC",X"16",X"D1",X"18",X"DF",X"1A",X"DC",X"1C",X"C6",X"1E",X"A0",X"20",X"69",X"22",
		X"22",X"24",X"CC",X"25",X"65",X"27",X"F0",X"28",X"6D",X"2A",X"DB",X"2B",X"39",X"2D",X"8F",X"2E",
		X"D3",X"2F",X"0F",X"31",X"3C",X"32",X"60",X"33",X"76",X"34",X"83",X"35",X"84",X"36",X"7C",X"37",
		X"68",X"38",X"4B",X"39",X"25",X"3A",X"F7",X"3A",X"BE",X"3B",X"80",X"3C",X"34",X"3D",X"E7",X"3D",
		X"8B",X"3E",X"30",X"3F",X"C4",X"3F",X"5B",X"40",X"DD",X"40",X"72",X"41",X"4D",X"41",X"85",X"3F",
		X"B2",X"3C",X"26",X"39",X"32",X"35",X"FC",X"30",X"A6",X"2C",X"45",X"28",X"EA",X"23",X"9B",X"1F",
		X"63",X"1B",X"41",X"17",X"3D",X"13",X"54",X"0F",X"88",X"0B",X"DA",X"07",X"4A",X"04",X"D5",X"00",
		X"7F",X"FD",X"44",X"FA",X"24",X"F7",X"1D",X"F4",X"33",X"F1",X"5F",X"EE",X"A5",X"EB",X"02",X"E9",
		X"76",X"E6",X"01",X"E4",X"A0",X"E1",X"56",X"DF",X"1E",X"DD",X"FB",X"DA",X"EB",X"D8",X"EF",X"D6",
		X"02",X"D5",X"28",X"D3",X"5E",X"D1",X"A6",X"CF",X"FD",X"CD",X"63",X"CC",X"D9",X"CA",X"5C",X"C9",
		X"ED",X"C7",X"8D",X"C6",X"3A",X"C5",X"F4",X"C3",X"BA",X"C2",X"8B",X"C1",X"69",X"C0",X"53",X"BF",
		X"46",X"BE",X"43",X"BD",X"4C",X"BC",X"5F",X"BB",X"7C",X"BA",X"A1",X"B9",X"D1",X"B8",X"08",X"B8",
		X"48",X"B7",X"90",X"B6",X"E1",X"B5",X"39",X"B5",X"98",X"B4",X"FF",X"B3",X"6D",X"B3",X"E3",X"B2",
		X"5E",X"B2",X"DF",X"B1",X"67",X"B1",X"F5",X"B0",X"8A",X"B0",X"24",X"B0",X"C2",X"AF",X"68",X"AF",
		X"11",X"AF",X"BF",X"AE",X"74",X"AE",X"2B",X"AE",X"E9",X"AD",X"AA",X"AD",X"6F",X"AD",X"38",X"AD",
		X"06",X"AD",X"D7",X"AC",X"AC",X"AC",X"85",X"AC",X"61",X"AC",X"41",X"AC",X"24",X"AC",X"09",X"AC",
		X"F2",X"AB",X"DF",X"AB",X"CF",X"AB",X"BF",X"AB",X"B6",X"AB",X"AC",X"AB",X"A6",X"AB",X"A2",X"AB",
		X"9E",X"AB",X"A0",X"AB",X"A3",X"AB",X"A7",X"AB",X"AF",X"AB",X"B8",X"AB",X"C3",X"AB",X"D1",X"AB",
		X"DF",X"AB",X"EE",X"AB",X"03",X"AC",X"15",X"AC",X"2A",X"AC",X"41",X"AC",X"59",X"AC",X"72",X"AC",
		X"8D",X"AC",X"AA",X"AC",X"C9",X"AC",X"E6",X"AC",X"07",X"AD",X"28",X"AD",X"4B",X"AD",X"6E",X"AD",
		X"93",X"AD",X"B7",X"AD",X"DD",X"AD",X"04",X"AE",X"2D",X"AE",X"54",X"AE",X"7E",X"AE",X"A8",X"AE",
		X"D6",X"AE",X"00",X"AF",X"2F",X"AF",X"5A",X"AF",X"8B",X"AF",X"B4",X"AF",X"EB",X"AF",X"11",X"B0",
		X"2C",X"B1",X"DD",X"B3",X"78",X"B7",X"BA",X"BB",X"52",X"C0",X"27",X"C5",X"0B",X"CA",X"F5",X"CE",
		X"D1",X"D3",X"9D",X"D8",X"4C",X"DD",X"E0",X"E1",X"50",X"E6",X"A4",X"EA",X"D5",X"EE",X"E7",X"F2",
		X"D5",X"F6",X"A4",X"FA",X"54",X"FE",X"E4",X"01",X"55",X"05",X"A9",X"08",X"E1",X"0B",X"FD",X"0E",
		X"FE",X"11",X"E5",X"14",X"B2",X"17",X"67",X"1A",X"04",X"1D",X"8C",X"1F",X"F9",X"21",X"53",X"24",
		X"97",X"26",X"C7",X"28",X"E0",X"2A",X"E8",X"2C",X"E2",X"2E",X"C3",X"30",X"96",X"32",X"56",X"34",
		X"07",X"36",X"A6",X"37",X"38",X"39",X"B9",X"3A",X"2C",X"3C",X"8F",X"3D",X"E8",X"3E",X"30",X"40",
		X"70",X"41",X"9B",X"42",X"C5",X"43",X"D8",X"44",X"EC",X"45",X"E4",X"46",X"EC",X"47",X"1D",X"48",
		X"AB",X"46",X"33",X"44",X"04",X"41",X"6B",X"3D",X"8D",X"39",X"92",X"35",X"87",X"31",X"80",X"2D",
		X"86",X"29",X"9B",X"25",X"C7",X"21",X"0B",X"1E",X"6B",X"1A",X"E3",X"16",X"7A",X"13",X"28",X"10",
		X"F3",X"0C",X"D5",X"09",X"D4",X"06",X"E9",X"03",X"1A",X"01",X"61",X"FE",X"C3",X"FB",X"31",X"F9",
		X"C4",X"F6",X"52",X"F4",X"99",X"F2",X"92",X"F2",X"A8",X"F3",X"89",X"F5",X"DE",X"F7",X"88",X"FA",
		X"5B",X"FD",X"42",X"00",X"32",X"03",X"20",X"06",X"03",X"09",X"D9",X"0B",X"9C",X"0E",X"4D",X"11",
		X"EC",X"13",X"72",X"16",X"E5",X"18",X"45",X"1B",X"8F",X"1D",X"C6",X"1F",X"EA",X"21",X"FA",X"23",
		X"F6",X"25",X"E4",X"27",X"BC",X"29",X"86",X"2B",X"3D",X"2D",X"DC",X"2E",X"2F",X"2F",X"FC",X"2D",
		X"E4",X"2B",X"2A",X"29",X"14",X"26",X"BF",X"22",X"50",X"1F",X"D3",X"1B",X"5A",X"18",X"EA",X"14",
		X"88",X"11",X"39",X"0E",X"02",X"0B",X"E1",X"07",X"D7",X"04",X"E4",X"01",X"0A",X"FF",X"46",X"FC",
		X"99",X"F9",X"04",X"F7",X"81",X"F4",X"18",X"F2",X"BF",X"EF",X"7F",X"ED",X"4D",X"EB",X"37",X"E9",
		X"22",X"E7",X"94",X"E5",X"AF",X"E5",X"FD",X"E6",X"17",X"E9",X"B0",X"EB",X"9C",X"EE",X"B3",X"F1",
		X"E2",X"F4",X"17",X"F8",X"49",X"FB",X"6D",X"FE",X"84",X"01",X"88",X"04",X"77",X"07",X"50",X"0A",
		X"13",X"0D",X"C0",X"0F",X"57",X"12",X"D5",X"14",X"42",X"17",X"98",X"19",X"DB",X"1B",X"07",X"1E",
		X"23",X"20",X"27",X"22",X"22",X"24",X"FE",X"25",X"D5",X"27",X"87",X"28",X"9C",X"27",X"C4",X"25",
		X"3C",X"23",X"52",X"20",X"23",X"1D",X"D7",X"19",X"7A",X"16",X"1F",X"13",X"C9",X"0F",X"86",X"0C",
		X"4E",X"09",X"31",X"06",X"25",X"03",X"32",X"00",X"56",X"FD",X"92",X"FA",X"E1",X"F7",X"4A",X"F5",
		X"C6",X"F2",X"59",X"F0",X"00",X"EE",X"BD",X"EB",X"8A",X"E9",X"6E",X"E7",X"62",X"E5",X"69",X"E3",
		X"81",X"E1",X"AA",X"DF",X"E3",X"DD",X"2E",X"DC",X"88",X"DA",X"F0",X"D8",X"67",X"D7",X"ED",X"D5",
		X"80",X"D4",X"1F",X"D3",X"CC",X"D1",X"85",X"D0",X"4B",X"CF",X"1C",X"CE",X"F9",X"CC",X"E1",X"CB",
		X"D5",X"CA",X"CF",X"C9",X"D8",X"C8",X"E6",X"C7",X"02",X"C7",X"23",X"C6",X"50",X"C5",X"83",X"C4",
		X"C4",X"C3",X"02",X"C3",X"59",X"C2",X"A0",X"C1",X"D8",X"C1",X"AC",X"C3",X"77",X"C6",X"F3",X"C9",
		X"CF",X"CD",X"EB",X"D1",X"1E",X"D6",X"61",X"DA",X"98",X"DE",X"C4",X"E2",X"D9",X"E6",X"DB",X"EA",
		X"BC",X"EE",X"85",X"F2",X"2D",X"F6",X"BC",X"F9",X"2C",X"FD",X"82",X"00",X"BB",X"03",X"D7",X"06",
		X"D9",X"09",X"C5",X"0C",X"95",X"0F",X"4C",X"12",X"EB",X"14",X"75",X"17",X"E8",X"19",X"44",X"1C",
		X"8B",X"1E",X"BE",X"20",X"DE",X"22",X"EA",X"24",X"E5",X"26",X"CA",X"28",X"A2",X"2A",X"67",X"2C",
		X"1A",X"2E",X"BF",X"2F",X"53",X"31",X"D9",X"32",X"51",X"34",X"BB",X"35",X"16",X"37",X"65",X"38",
		X"A7",X"39",X"DC",X"3A",X"06",X"3C",X"21",X"3D",X"35",X"3E",X"3A",X"3F",X"38",X"40",X"28",X"41",
		X"10",X"42",X"EF",X"42",X"C4",X"43",X"8E",X"44",X"51",X"45",X"0C",X"46",X"BD",X"46",X"68",X"47",
		X"09",X"48",X"A5",X"48",X"36",X"49",X"C4",X"49",X"48",X"4A",X"C7",X"4A",X"3E",X"4B",X"B0",X"4B",
		X"1C",X"4C",X"83",X"4C",X"E2",X"4C",X"3D",X"4D",X"92",X"4D",X"E2",X"4D",X"2E",X"4E",X"73",X"4E",
		X"B7",X"4E",X"F2",X"4E",X"2E",X"4F",X"5F",X"4F",X"92",X"4F",X"BC",X"4F",X"D4",X"4F",X"97",X"4E",
		X"EC",X"4B",X"6C",X"48",X"58",X"44",X"F5",X"3F",X"63",X"3B",X"BE",X"36",X"17",X"32",X"7F",X"2D",
		X"F6",X"28",X"88",X"24",X"36",X"20",X"FF",X"1B",X"EA",X"17",X"F3",X"13",X"1C",X"10",X"60",X"0C",
		X"C8",X"08",X"4B",X"05",X"EC",X"01",X"A9",X"FE",X"82",X"FB",X"72",X"F8",X"81",X"F5",X"A3",X"F2",
		X"E7",X"EF",X"30",X"ED",X"1A",X"EB",X"B8",X"EA",X"80",X"EB",X"17",X"ED",X"2E",X"EF",X"99",X"F1",
		X"31",X"F4",X"E6",X"F6",X"A1",X"F9",X"5E",X"FC",X"12",X"FF",X"BC",X"01",X"53",X"04",X"DC",X"06",
		X"51",X"09",X"B5",X"0B",X"02",X"0E",X"3E",X"10",X"68",X"12",X"80",X"14",X"84",X"16",X"79",X"18",
		X"58",X"1A",X"2A",X"1C",X"EA",X"1D",X"9C",X"1F",X"3A",X"21",X"CB",X"22",X"23",X"23",X"EE",X"21",
		X"D1",X"1F",X"0A",X"1D",X"E6",X"19",X"83",X"16",X"05",X"13",X"79",X"0F",X"F3",X"0B",X"72",X"08",
		X"03",X"05",X"A7",X"01",X"64",X"FE",X"34",X"FB",X"20",X"F8",X"23",X"F5",X"3D",X"F2",X"6E",X"EF",
		X"BA",X"EC",X"1A",X"EA",X"93",X"E7",X"20",X"E5",X"C2",X"E2",X"7B",X"E0",X"46",X"DE",X"25",X"DC",
		X"19",X"DA",X"1D",X"D8",X"34",X"D6",X"5C",X"D4",X"96",X"D2",X"DD",X"D0",X"37",X"CF",X"9E",X"CD",
		X"17",X"CC",X"9B",X"CA",X"30",X"C9",X"D0",X"C7",X"80",X"C6",X"38",X"C5",X"01",X"C4",X"D5",X"C2",
		X"B3",X"C1",X"9D",X"C0",X"92",X"BF",X"91",X"BE",X"9C",X"BD",X"B0",X"BC",X"CC",X"BB",X"F2",X"BA",
		X"24",X"BA",X"5B",X"B9",X"9D",X"B8",X"E6",X"B7",X"37",X"B7",X"90",X"B6",X"F1",X"B5",X"56",X"B5",
		X"C7",X"B4",X"3C",X"B4",X"B9",X"B3",X"3A",X"B3",X"C4",X"B2",X"52",X"B2",X"E8",X"B1",X"81",X"B1",
		X"22",X"B1",X"C7",X"B0",X"71",X"B0",X"1E",X"B0",X"D4",X"AF",X"8C",X"AF",X"49",X"AF",X"0B",X"AF",
		X"D0",X"AE",X"98",X"AE",X"67",X"AE",X"39",X"AE",X"0F",X"AE",X"E6",X"AD",X"C6",X"AD",X"9E",X"AD",
		X"B7",X"AD",X"52",X"AF",X"34",X"B2",X"E0",X"B5",X"0E",X"BA",X"83",X"BE",X"24",X"C3",X"D2",X"C7",
		X"7D",X"CC",X"1A",X"D1",X"A3",X"D5",X"12",X"DA",X"64",X"DE",X"97",X"E2",X"AD",X"E6",X"A1",X"EA",
		X"77",X"EE",X"2E",X"F2",X"C7",X"F5",X"41",X"F9",X"9F",X"FC",X"DE",X"FF",X"03",X"03",X"0D",X"06",
		X"FD",X"08",X"D2",X"0B",X"90",X"0E",X"36",X"11",X"C5",X"13",X"3C",X"16",X"A0",X"18",X"ED",X"1A",
		X"27",X"1D",X"4A",X"1F",X"5E",X"21",X"5C",X"23",X"49",X"25",X"23",X"27",X"EF",X"28",X"A6",X"2A",
		X"50",X"2C",X"E9",X"2D",X"75",X"2F",X"F0",X"30",X"60",X"32",X"BE",X"33",X"11",X"35",X"58",X"36",
		X"91",X"37",X"BE",X"38",X"E1",X"39",X"F7",X"3A",X"02",X"3C",X"02",X"3D",X"F9",X"3D",X"CC",X"3E",
		X"30",X"3E",X"2B",X"3C",X"53",X"39",X"E4",X"35",X"25",X"32",X"32",X"2E",X"2C",X"2A",X"1C",X"26",
		X"19",X"22",X"21",X"1E",X"40",X"1A",X"73",X"16",X"C4",X"12",X"2D",X"0F",X"B4",X"0B",X"53",X"08",
		X"0F",X"05",X"E4",X"01",X"D5",X"FE",X"E0",X"FB",X"02",X"F9",X"3E",X"F6",X"90",X"F3",X"FA",X"F0",
		X"78",X"EE",X"10",X"EC",X"C6",X"E9",X"D5",X"E8",X"6A",X"E9",X"E6",X"EA",X"09",X"ED",X"8C",X"EF",
		X"4E",X"F2",X"2F",X"F5",X"22",X"F8",X"15",X"FB",X"03",X"FE",X"E3",X"00",X"B4",X"03",X"72",X"06",
		X"20",X"09",X"B7",X"0B",X"3A",X"0E",X"A9",X"10",X"03",X"13",X"4A",X"15",X"7C",X"17",X"9C",X"19",
		X"A6",X"1B",X"A3",X"1D",X"88",X"1F",X"63",X"21",X"26",X"23",X"E8",X"24",X"1F",X"26",X"AC",X"25",
		X"0D",X"24",X"A4",X"21",X"C2",X"1E",X"8F",X"1B",X"31",X"18",X"C0",X"14",X"4A",X"11",X"DA",X"0D",
		X"74",X"0A",X"22",X"07",X"E4",X"03",X"BD",X"00",X"AE",X"FD",X"B4",X"FA",X"D2",X"F7",X"09",X"F5",
		X"55",X"F2",X"BA",X"EF",X"33",X"ED",X"C3",X"EA",X"67",X"E8",X"21",X"E6",X"EE",X"E3",X"D0",X"E1",
		X"C2",X"DF",X"C9",X"DD",X"DE",X"DB",X"09",X"DA",X"42",X"D8",X"8D",X"D6",X"E4",X"D4",X"4E",X"D3",
		X"C4",X"D1",X"4A",X"D0",X"DB",X"CE",X"7E",X"CD",X"2A",X"CC",X"E6",X"CA",X"AB",X"C9",X"7F",X"C8",
		X"5B",X"C7",X"45",X"C6",X"37",X"C5",X"36",X"C4",X"3F",X"C3",X"53",X"C2",X"6C",X"C1",X"93",X"C0",
		X"BE",X"BF",X"F8",X"BE",X"35",X"BE",X"81",X"BD",X"C5",X"BC",X"68",X"BC",X"9D",X"BD",X"0F",X"C0",
		X"49",X"C3",X"02",X"C7",X"08",X"CB",X"34",X"CF",X"70",X"D3",X"AD",X"D7",X"DF",X"DB",X"FE",X"DF",
		X"06",X"E4",X"F7",X"E7",X"C9",X"EB",X"82",X"EF",X"1A",X"F3",X"99",X"F6",X"FB",X"F9",X"3F",X"FD",
		X"67",X"00",X"78",X"03",X"6E",X"06",X"49",X"09",X"0C",X"0C",X"B8",X"0E",X"4C",X"11",X"CA",X"13",
		X"31",X"16",X"84",X"18",X"C2",X"1A",X"EB",X"1C",X"01",X"1F",X"06",X"21",X"F5",X"22",X"D5",X"24",
		X"A4",X"26",X"62",X"28",X"0F",X"2A",X"AE",X"2B",X"3E",X"2D",X"BD",X"2E",X"2F",X"30",X"94",X"31",
		X"EA",X"32",X"34",X"34",X"72",X"35",X"A1",X"36",X"C6",X"37",X"E1",X"38",X"EF",X"39",X"F5",X"3A",
		X"EB",X"3B",X"DC",X"3C",X"C0",X"3D",X"A1",X"3E",X"49",X"3F",X"6F",X"3E",X"3E",X"3C",X"40",X"39",
		X"B6",X"35",X"DC",X"31",X"D2",X"2D",X"B6",X"29",X"96",X"25",X"80",X"21",X"79",X"1D",X"8A",X"19",
		X"AF",X"15",X"F1",X"11",X"4F",X"0E",X"C7",X"0A",X"5C",X"07",X"0C",X"04",X"D8",X"00",X"BF",X"FD",
		X"BC",X"FA",X"D6",X"F7",X"08",X"F5",X"52",X"F2",X"B2",X"EF",X"2B",X"ED",X"B8",X"EA",X"5E",X"E8",
		X"14",X"E6",X"DF",X"E3",X"BE",X"E1",X"B2",X"DF",X"B5",X"DD",X"CD",X"DB",X"F4",X"D9",X"2C",X"D8",
		X"73",X"D6",X"CD",X"D4",X"33",X"D3",X"A8",X"D1",X"2D",X"D0",X"C1",X"CE",X"5F",X"CD",X"0D",X"CC",
		X"C8",X"CA",X"8D",X"C9",X"5E",X"C8",X"3D",X"C7",X"24",X"C6",X"17",X"C5",X"15",X"C4",X"1D",X"C3",
		X"2E",X"C2",X"4B",X"C1",X"6E",X"C0",X"9D",X"BF",X"D2",X"BE",X"12",X"BE",X"58",X"BD",X"A8",X"BC",
		X"FD",X"BB",X"5C",X"BB",X"C1",X"BA",X"2E",X"BA",X"A1",X"B9",X"1C",X"B9",X"9A",X"B8",X"21",X"B8",
		X"AB",X"B7",X"3F",X"B7",X"D5",X"B6",X"74",X"B6",X"14",X"B6",X"BE",X"B5",X"67",X"B5",X"1B",X"B5",
		X"CE",X"B4",X"8B",X"B4",X"46",X"B4",X"0E",X"B4",X"CF",X"B3",X"A1",X"B3",X"5F",X"B3",X"B9",X"B3",
		X"B0",X"B5",X"BE",X"B8",X"86",X"BC",X"B9",X"C0",X"32",X"C5",X"C7",X"C9",X"68",X"CE",X"01",X"D3",
		X"8D",X"D7",X"00",X"DC",X"5B",X"E0",X"98",X"E4",X"B7",X"E8",X"B6",X"EC",X"97",X"F0",X"58",X"F4",
		X"FC",X"F7",X"80",X"FB",X"E7",X"FE",X"30",X"02",X"5F",X"05",X"72",X"08",X"6E",X"0B",X"49",X"0E",
		X"12",X"11",X"BC",X"13",X"50",X"16",X"9D",X"17",X"54",X"17",X"1F",X"16",X"3A",X"14",X"F4",X"11",
		X"66",X"0F",X"B7",X"0C",X"F2",X"09",X"2F",X"07",X"68",X"04",X"B2",X"01",X"07",X"FF",X"6E",X"FC",
		X"E6",X"F9",X"72",X"F7",X"0E",X"F5",X"C0",X"F2",X"82",X"F0",X"58",X"EE",X"41",X"EC",X"3D",X"EA",
		X"47",X"E8",X"66",X"E6",X"95",X"E4",X"D2",X"E2",X"20",X"E1",X"7D",X"DF",X"E8",X"DD",X"64",X"DC",
		X"EA",X"DA",X"80",X"D9",X"24",X"D8",X"D2",X"D6",X"8F",X"D5",X"56",X"D4",X"29",X"D3",X"07",X"D2",
		X"F2",X"D0",X"E4",X"CF",X"E3",X"CE",X"EA",X"CD",X"FD",X"CC",X"18",X"CC",X"3C",X"CB",X"67",X"CA",
		X"9E",X"C9",X"D9",X"C8",X"21",X"C8",X"6C",X"C7",X"C2",X"C6",X"1B",X"C6",X"83",X"C5",X"E7",X"C4",
		X"5D",X"C4",X"CC",X"C3",X"48",X"C4",X"57",X"C6",X"51",X"C9",X"F6",X"CC",X"F4",X"D0",X"2E",X"D5",
		X"7F",X"D9",X"DA",X"DD",X"27",X"E2",X"6C",X"E6",X"95",X"EA",X"A9",X"EE",X"9E",X"F2",X"77",X"F6",
		X"35",X"FA",X"D2",X"FD",X"54",X"01",X"B7",X"04",X"FD",X"07",X"2A",X"0B",X"3A",X"0E",X"32",X"11",
		X"0D",X"14",X"D2",X"16",X"7D",X"19",X"10",X"1C",X"8F",X"1E",X"F4",X"20",X"46",X"23",X"82",X"25",
		X"AC",X"27",X"C0",X"29",X"C2",X"2B",X"B0",X"2D",X"8F",X"2F",X"5A",X"31",X"14",X"33",X"C1",X"34",
		X"5D",X"36",X"E7",X"37",X"64",X"39",X"D3",X"3A",X"35",X"3C",X"87",X"3D",X"CD",X"3E",X"07",X"40",
		X"36",X"41",X"54",X"42",X"6D",X"43",X"73",X"44",X"75",X"45",X"67",X"46",X"57",X"47",X"2F",X"48",
		X"14",X"49",X"17",X"49",X"77",X"47",X"DA",X"44",X"87",X"41",X"D1",X"3D",X"D6",X"39",X"C1",X"35",
		X"9E",X"31",X"82",X"2D",X"70",X"29",X"71",X"25",X"88",X"21",X"BA",X"1D",X"07",X"1A",X"70",X"16",
		X"F2",X"12",X"91",X"0F",X"4B",X"0C",X"22",X"09",X"10",X"06",X"19",X"03",X"3B",X"00",X"77",X"FD",
		X"C7",X"FA",X"2F",X"F8",X"AE",X"F5",X"42",X"F3",X"EC",X"F0",X"A9",X"EE",X"79",X"EC",X"5E",X"EA",
		X"54",X"E8",X"5C",X"E6",X"76",X"E4",X"A1",X"E2",X"DD",X"E0",X"29",X"DF",X"83",X"DD",X"ED",X"DB",
		X"65",X"DA",X"EA",X"D8",X"7E",X"D7",X"1F",X"D6",X"CE",X"D4",X"89",X"D3",X"4E",X"D2",X"20",X"D1",
		X"FD",X"CF",X"E5",X"CE",X"D8",X"CD",X"D5",X"CC",X"DC",X"CB",X"ED",X"CA",X"07",X"CA",X"2B",X"C9",
		X"57",X"C8",X"8C",X"C7",X"C8",X"C6",X"0E",X"C6",X"5B",X"C5",X"AF",X"C4",X"0B",X"C4",X"6D",X"C3",
		X"D7",X"C2",X"47",X"C2",X"BE",X"C1",X"3B",X"C1",X"BF",X"C0",X"47",X"C0",X"D6",X"BF",X"6A",X"BF",
		X"03",X"BF",X"A1",X"BE",X"47",X"BE",X"EE",X"BD",X"9C",X"BD",X"4D",X"BD",X"03",X"BD",X"BE",X"BC",
		X"7B",X"BC",X"40",X"BC",X"06",X"BC",X"D0",X"BB",X"9D",X"BB",X"71",X"BB",X"45",X"BB",X"1C",X"BB",
		X"F8",X"BA",X"D6",X"BA",X"B8",X"BA",X"9D",X"BA",X"83",X"BA",X"6E",X"BA",X"5A",X"BA",X"4A",X"BA",
		X"3B",X"BA",X"30",X"BA",X"25",X"BA",X"1E",X"BA",X"19",X"BA",X"18",X"BA",X"13",X"BA",X"16",X"BA",
		X"17",X"BA",X"1E",X"BA",X"21",X"BA",X"2C",X"BA",X"33",X"BA",X"42",X"BA",X"4F",X"BA",X"80",X"BB",
		X"34",X"BE",X"C8",X"C1",X"F9",X"C5",X"7E",X"CA",X"36",X"CF",X"00",X"D4",X"CC",X"D8",X"8B",X"DD",
		X"39",X"E2",X"CB",X"E6",X"41",X"EB",X"97",X"EF",X"CD",X"F3",X"E3",X"F7",X"D8",X"FB",X"AB",X"FF",
		X"61",X"03",X"F6",X"06",X"71",X"0A",X"C8",X"0D",X"06",X"11",X"26",X"14",X"2D",X"17",X"19",X"1A",
		X"EB",X"1C",X"A4",X"1F",X"45",X"22",X"CD",X"24",X"41",X"27",X"9E",X"29",X"E5",X"2B",X"17",X"2E",
		X"37",X"30",X"41",X"32",X"3A",X"34",X"20",X"36",X"F2",X"37",X"B5",X"39",X"68",X"3B",X"09",X"3D",
		X"9C",X"3E",X"1E",X"40",X"93",X"41",X"F9",X"42",X"51",X"44",X"9C",X"45",X"D9",X"46",X"09",X"48",
		X"2E",X"49",X"47",X"4A",X"55",X"4B",X"56",X"4C",X"4E",X"4D",X"3B",X"4E",X"1E",X"4F",X"F6",X"4F",
		X"C6",X"50",X"8D",X"51",X"4A",X"52",X"FC",X"52",X"AA",X"53",X"4E",X"54",X"EA",X"54",X"7D",X"55",
		X"0C",X"56",X"90",X"56",X"0F",X"57",X"86",X"57",X"F9",X"57",X"65",X"58",X"CB",X"58",X"29",X"59",
		X"83",X"59",X"D6",X"59",X"27",X"5A",X"6F",X"5A",X"B3",X"5A",X"F1",X"5A",X"2C",X"5B",X"60",X"5B",
		X"98",X"5B",X"95",X"5B",X"12",X"5A",X"42",X"57",X"A7",X"53",X"86",X"4F",X"1D",X"4B",X"88",X"46",
		X"E6",X"41",X"43",X"3D",X"AD",X"38",X"2D",X"34",X"C5",X"2F",X"77",X"2B",X"48",X"27",X"37",X"23",
		X"46",X"1F",X"72",X"1B",X"BF",X"17",X"28",X"14",X"B0",X"10",X"52",X"0D",X"12",X"0A",X"EE",X"06",
		X"E2",X"03",X"F1",X"00",X"1B",X"FE",X"5A",X"FB",X"B3",X"F8",X"20",X"F6",X"A6",X"F3",X"3F",X"F1",
		X"EE",X"EE",X"B1",X"EC",X"89",X"EA",X"72",X"E8",X"6E",X"E6",X"7A",X"E4",X"9B",X"E2",X"CB",X"E0",
		X"0A",X"DF",X"58",X"DD",X"BA",X"DB",X"26",X"DA",X"A4",X"D8",X"2E",X"D7",X"C7",X"D5",X"6B",X"D4",
		X"1E",X"D3",X"DC",X"D1",X"A6",X"D0",X"7C",X"CF",X"5B",X"CE",X"47",X"CD",X"3D",X"CC",X"40",X"CB",
		X"49",X"CA",X"5E",X"C9",X"7B",X"C8",X"A1",X"C7",X"D1",X"C6",X"08",X"C6",X"4A",X"C5",X"92",X"C4",
		X"E0",X"C3",X"39",X"C3",X"97",X"C2",X"FB",X"C1",X"67",X"C1",X"DB",X"C0",X"54",X"C0",X"D5",X"BF",
		X"59",X"BF",X"E6",X"BE",X"76",X"BE",X"0C",X"BE",X"A8",X"BD",X"48",X"BD",X"EF",X"BC",X"9A",X"BC",
		X"4A",X"BC",X"FD",X"BB",X"B5",X"BB",X"72",X"BB",X"32",X"BB",X"F8",X"BA",X"C0",X"BA",X"8B",X"BA",
		X"5D",X"BA",X"30",X"BA",X"06",X"BA",X"DF",X"B9",X"BD",X"B9",X"9E",X"B9",X"81",X"B9",X"68",X"B9",
		X"51",X"B9",X"3D",X"B9",X"2C",X"B9",X"1C",X"B9",X"10",X"B9",X"04",X"B9",X"FD",X"B8",X"F6",X"B8",
		X"F2",X"B8",X"F0",X"B8",X"F2",X"B8",X"F4",X"B8",X"F9",X"B8",X"FE",X"B8",X"06",X"B9",X"10",X"B9",
		X"1A",X"B9",X"28",X"B9",X"35",X"B9",X"44",X"B9",X"56",X"B9",X"69",X"B9",X"7D",X"B9",X"90",X"B9",
		X"A6",X"B9",X"BE",X"B9",X"D8",X"B9",X"F0",X"B9",X"0D",X"BA",X"27",X"BA",X"45",X"BA",X"64",X"BA",
		X"82",X"BA",X"A1",X"BA",X"C2",X"BA",X"E2",X"BA",X"04",X"BB",X"28",X"BB",X"4C",X"BB",X"70",X"BB",
		X"96",X"BB",X"BB",X"BB",X"E2",X"BB",X"08",X"BC",X"30",X"BC",X"58",X"BC",X"81",X"BC",X"AA",X"BC",
		X"D4",X"BC",X"FF",X"BC",X"29",X"BD",X"54",X"BD",X"7F",X"BD",X"AB",X"BD",X"D7",X"BD",X"05",X"BE",
		X"30",X"BE",X"5F",X"BE",X"8C",X"BE",X"BB",X"BE",X"E8",X"BE",X"18",X"BF",X"46",X"BF",X"76",X"BF",
		X"A3",X"BF",X"D4",X"BF",X"02",X"C0",X"34",X"C0",X"62",X"C0",X"99",X"C0",X"C1",X"C0",X"F9",X"C1",
		X"BE",X"C4",X"65",X"C8",X"AF",X"CC",X"4B",X"D1",X"20",X"D6",X"01",X"DB",X"EA",X"DF",X"C3",X"E4",
		X"8B",X"E9",X"35",X"EE",X"C2",X"F2",X"30",X"F7",X"7E",X"FB",X"A7",X"FF",X"B1",X"03",X"98",X"07",
		X"62",X"0B",X"0A",X"0F",X"94",X"12",X"FE",X"15",X"4B",X"19",X"7C",X"1C",X"8F",X"1F",X"8A",X"22",
		X"69",X"25",X"2F",X"28",X"DC",X"2A",X"70",X"2D",X"ED",X"2F",X"55",X"32",X"A5",X"34",X"E2",X"36",
		X"08",X"39",X"1C",X"3B",X"1C",X"3D",X"08",X"3F",X"E1",X"40",X"AD",X"42",X"65",X"44",X"0B",X"46",
		X"A2",X"47",X"2B",X"49",X"A2",X"4A",X"0D",X"4C",X"67",X"4D",X"B5",X"4E",X"F4",X"4F",X"2B",X"51",
		X"4E",X"52",X"6D",X"53",X"77",X"54",X"82",X"55",X"72",X"56",X"6E",X"57",X"7D",X"57",X"EA",X"55",
		X"5C",X"53",X"19",X"50",X"72",X"4C",X"89",X"48",X"82",X"44",X"6D",X"40",X"5F",X"3C",X"5B",X"38",
		X"6B",X"34",X"8E",X"30",X"CB",X"2C",X"22",X"29",X"95",X"25",X"20",X"22",X"CB",X"1E",X"8A",X"1B",
		X"69",X"18",X"5F",X"15",X"6D",X"12",X"95",X"0F",X"D4",X"0C",X"29",X"0A",X"96",X"07",X"18",X"05",
		X"B0",X"02",X"5C",X"00",X"1C",X"FE",X"EE",X"FB",X"D3",X"F9",X"CC",X"F7",X"D4",X"F5",X"EF",X"F3",
		X"19",X"F2",X"54",X"F0",X"9E",X"EE",X"F9",X"EC",X"5E",X"EB",X"D7",X"E9",X"5A",X"E8",X"ED",X"E6",
		X"88",X"E5",X"35",X"E4",X"EA",X"E2",X"AE",X"E1",X"7A",X"E0",X"56",X"DF",X"37",X"DE",X"27",X"DD",
		X"1E",X"DC",X"23",X"DB",X"29",X"DA",X"47",X"D9",X"53",X"D8",X"1D",X"D8",X"8D",X"D9",X"0B",X"DC",
		X"3F",X"DF",X"DF",X"E2",X"C6",X"E6",X"CA",X"EA",X"DD",X"EE",X"EC",X"F2",X"F0",X"F6",X"DF",X"FA",
		X"B8",X"FE",X"76",X"02",X"1C",X"06",X"A4",X"09",X"12",X"0D",X"60",X"10",X"96",X"13",X"B1",X"16",
		X"AF",X"19",X"94",X"1C",X"60",X"1F",X"13",X"22",X"B0",X"24",X"32",X"27",X"A1",X"29",X"F8",X"2B",
		X"2D",X"2E",X"01",X"2F",X"52",X"2E",X"BF",X"2C",X"88",X"2A",X"F1",X"27",X"17",X"25",X"25",X"22",
		X"1B",X"1F",X"16",X"1C",X"13",X"19",X"1F",X"16",X"38",X"13",X"67",X"10",X"A5",X"0D",X"FB",X"0A",
		X"62",X"08",X"E1",X"05",X"70",X"03",X"16",X"01",X"CF",X"FE",X"9B",X"FC",X"7A",X"FA",X"6B",X"F8",
		X"6C",X"F6",X"81",X"F4",X"A4",X"F2",X"DB",X"F0",X"1D",X"EF",X"72",X"ED",X"D3",X"EB",X"43",X"EA",
		X"C2",X"E8",X"4F",X"E7",X"E7",X"E5",X"8C",X"E4",X"3F",X"E3",X"FB",X"E1",X"C6",X"E0",X"9C",X"DF",
		X"7B",X"DE",X"65",X"DD",X"58",X"DC",X"57",X"DB",X"5F",X"DA",X"70",X"D9",X"8B",X"D8",X"AD",X"D7",
		X"DA",X"D6",X"0C",X"D6",X"4A",X"D5",X"89",X"D4",X"D7",X"D3",X"26",X"D3",X"84",X"D2",X"E4",X"D1",
		X"6E",X"D2",X"81",X"D4",X"74",X"D7",X"0D",X"DB",X"FD",X"DE",X"26",X"E3",X"61",X"E7",X"A8",X"EB",
		X"E3",X"EF",X"10",X"F4",X"26",X"F8",X"22",X"FC",X"04",X"00",X"C8",X"03",X"70",X"07",X"FA",X"0A",
		X"67",X"0E",X"B7",X"11",X"ED",X"14",X"04",X"18",X"04",X"1B",X"E7",X"1D",X"B4",X"20",X"63",X"23",
		X"02",X"26",X"7E",X"28",X"F4",X"2A",X"53",X"2C",X"0D",X"2C",X"CA",X"2A",X"D0",X"28",X"6C",X"26",
		X"BE",X"23",X"EA",X"20",X"03",X"1E",X"18",X"1B",X"2F",X"18",X"52",X"15",X"82",X"12",X"C3",X"0F",
		X"16",X"0D",X"7D",X"0A",X"F5",X"07",X"84",X"05",X"25",X"03",X"DA",X"00",X"A2",X"FE",X"7D",X"FC",
		X"6A",X"FA",X"67",X"F8",X"78",X"F6",X"97",X"F4",X"CA",X"F2",X"06",X"F1",X"8A",X"EF",X"9E",X"EF",
		X"05",X"F1",X"41",X"F3",X"07",X"F6",X"23",X"F9",X"70",X"FC",X"D4",X"FF",X"40",X"03",X"A8",X"06",
		X"03",X"0A",X"4F",X"0D",X"84",X"10",X"A5",X"13",X"AC",X"16",X"9E",X"19",X"76",X"1C",X"39",X"1F",
		X"E0",X"21",X"75",X"24",X"EF",X"26",X"59",X"29",X"A7",X"2B",X"E3",X"2D",X"08",X"30",X"1F",X"32",
		X"1A",X"34",X"16",X"36",X"2F",X"37",X"9A",X"36",X"FE",X"34",X"A3",X"32",X"DD",X"2F",X"C9",X"2C",
		X"95",X"29",X"4A",X"26",X"FE",X"22",X"B4",X"1F",X"7B",X"1C",X"4F",X"19",X"39",X"16",X"36",X"13",
		X"4A",X"10",X"72",X"0D",X"B4",X"0A",X"09",X"08",X"75",X"05",X"F6",X"02",X"8D",X"00",X"36",X"FE",
		X"F5",X"FB",X"C5",X"F9",X"AC",X"F7",X"A0",X"F5",X"A6",X"F3",X"DA",X"F1",X"83",X"F1",X"99",X"F2",
		X"8C",X"F4",X"17",X"F7",X"FD",X"F9",X"1A",X"FD",X"53",X"00",X"95",X"03",X"D6",X"06",X"0E",X"0A",
		X"36",X"0D",X"4C",X"10",X"4D",X"13",X"37",X"16",X"0B",X"19",X"C7",X"1B",X"6F",X"1E",X"FC",X"20",
		X"77",X"23",X"D7",X"25",X"29",X"28",X"61",X"2A",X"88",X"2C",X"97",X"2E",X"9A",X"30",X"81",X"32",
		X"6A",X"34",X"A1",X"35",X"25",X"35",X"92",X"33",X"39",X"31",X"6B",X"2E",X"4E",X"2B",X"0B",X"28",
		X"B2",X"24",X"55",X"21",X"FD",X"1D",X"B3",X"1A",X"78",X"17",X"53",X"14",X"3F",X"11",X"45",X"0E",
		X"5F",X"0B",X"91",X"08",X"D8",X"05",X"38",X"03",X"AA",X"00",X"36",X"FE",X"D4",X"FB",X"88",X"F9",
		X"4C",X"F7",X"28",X"F5",X"12",X"F3",X"12",X"F1",X"29",X"EF",X"90",X"EE",X"7E",X"EF",X"51",X"F1",
		X"CA",X"F3",X"9E",X"F6",X"B3",X"F9",X"E3",X"FC",X"21",X"00",X"5C",X"03",X"93",X"06",X"B8",X"09",
		X"CD",X"0C",X"CB",X"0F",X"B4",X"12",X"87",X"15",X"45",X"18",X"EA",X"1A",X"79",X"1D",X"F3",X"1F",
		X"57",X"22",X"A5",X"24",X"DE",X"26",X"05",X"29",X"15",X"2B",X"19",X"2D",X"01",X"2F",X"E8",X"30",
		X"4C",X"32",X"01",X"32",X"87",X"30",X"41",X"2E",X"7D",X"2B",X"69",X"28",X"27",X"25",X"D0",X"21",
		X"73",X"1E",X"19",X"1B",X"CD",X"17",X"8F",X"14",X"67",X"11",X"51",X"0E",X"54",X"0B",X"6D",X"08",
		X"9C",X"05",X"E1",X"02",X"3E",X"00",X"B0",X"FD",X"37",X"FB",X"D1",X"F8",X"85",X"F6",X"47",X"F4",
		X"22",X"F2",X"09",X"F0",X"0A",X"EE",X"13",X"EC",X"43",X"EB",X"0E",X"EC",X"C9",X"ED",X"33",X"F0",
		X"FF",X"F2",X"10",X"F6",X"3D",X"F9",X"7D",X"FC",X"B9",X"FF",X"F1",X"02",X"1A",X"06",X"32",X"09",
		X"34",X"0C",X"24",X"0F",X"FB",X"11",X"BC",X"14",X"65",X"17",X"FB",X"19",X"79",X"1C",X"E0",X"1E",
		X"33",X"21",X"6F",X"23",X"9B",X"25",X"B1",X"27",X"B6",X"29",X"A4",X"2B",X"8D",X"2D",X"16",X"2F",
		X"02",X"2F",X"A7",X"2D",X"7A",X"2B",X"C5",X"28",X"BB",X"25",X"7F",X"22",X"2C",X"1F",X"D2",X"1B",
		X"78",X"18",X"2C",X"15",X"ED",X"11",X"C5",X"0E",X"AF",X"0B",X"B0",X"08",X"C8",X"05",X"F5",X"02",
		X"3D",X"00",X"96",X"FD",X"08",X"FB",X"8E",X"F8",X"2A",X"F6",X"DB",X"F3",X"A0",X"F1",X"75",X"EF",
		X"61",X"ED",X"5C",X"EB",X"6B",X"E9",X"89",X"E7",X"BC",X"E5",X"FA",X"E3",X"4A",X"E2",X"A9",X"E0",
		X"18",X"DF",X"92",X"DD",X"1C",X"DC",X"B4",X"DA",X"59",X"D9",X"08",X"D8",X"C7",X"D6",X"8F",X"D5",
		X"64",X"D4",X"42",X"D3",X"2F",X"D2",X"22",X"D1",X"23",X"D0",X"2A",X"CF",X"3E",X"CE",X"59",X"CD",
		X"7E",X"CC",X"AB",X"CB",X"E1",X"CA",X"1E",X"CA",X"67",X"C9",X"AF",X"C8",X"2D",X"C8",X"23",X"C9",
		X"73",X"CB",X"90",X"CE",X"3D",X"D2",X"36",X"D6",X"5D",X"DA",X"96",X"DE",X"D2",X"E2",X"03",X"E7",
		X"23",X"EB",X"2A",X"EF",X"1D",X"F3",X"F0",X"F6",X"A8",X"FA",X"42",X"FE",X"C0",X"01",X"21",X"05",
		X"67",X"08",X"91",X"0B",X"A0",X"0E",X"95",X"11",X"6F",X"14",X"32",X"17",X"DC",X"19",X"6E",X"1C",
		X"EA",X"1E",X"4E",X"21",X"A0",X"23",X"DC",X"25",X"03",X"28",X"16",X"2A",X"18",X"2C",X"07",X"2E",
		X"E4",X"2F",X"AB",X"31",X"68",X"33",X"13",X"35",X"AD",X"36",X"38",X"38",X"B5",X"39",X"21",X"3B",
		X"81",X"3C",X"D4",X"3D",X"1A",X"3F",X"52",X"40",X"7F",X"41",X"A0",X"42",X"B5",X"43",X"BE",X"44",
		X"BD",X"45",X"B3",X"46",X"9B",X"47",X"7E",X"48",X"53",X"49",X"0F",X"4A",X"70",X"49",X"5D",X"47",
		X"73",X"44",X"F1",X"40",X"1A",X"3D",X"0D",X"39",X"EE",X"34",X"C5",X"30",X"A7",X"2C",X"97",X"28",
		X"9E",X"24",X"B9",X"20",X"F1",X"1C",X"41",X"19",X"B0",X"15",X"39",X"12",X"DF",X"0E",X"A1",X"0B",
		X"7B",X"08",X"70",X"05",X"7F",X"02",X"A6",X"FF",X"E7",X"FC",X"3D",X"FA",X"AB",X"F7",X"2E",X"F5",
		X"C8",X"F2",X"75",X"F0",X"38",X"EE",X"0D",X"EC",X"F6",X"E9",X"F1",X"E7",X"FF",X"E5",X"1D",X"E4",
		X"4C",X"E2",X"8A",X"E0",X"DA",X"DE",X"38",X"DD",X"A4",X"DB",X"20",X"DA",X"AA",X"D8",X"41",X"D7",
		X"E7",X"D5",X"97",X"D4",X"55",X"D3",X"1E",X"D2",X"F1",X"D0",X"D4",X"CF",X"BE",X"CE",X"B3",X"CD",
		X"B1",X"CC",X"BE",X"CB",X"CD",X"CA",X"EF",X"C9",X"15",X"C9",X"70",X"C9",X"51",X"CB",X"18",X"CE",
		X"81",X"D1",X"41",X"D5",X"3C",X"D9",X"4C",X"DD",X"66",X"E1",X"7B",X"E5",X"7F",X"E9",X"6D",X"ED",
		X"45",X"F1",X"04",X"F5",X"A5",X"F8",X"2D",X"FC",X"96",X"FF",X"E6",X"02",X"19",X"06",X"33",X"09",
		X"30",X"0C",X"15",X"0F",X"E1",X"11",X"95",X"14",X"2F",X"17",X"B8",X"19",X"22",X"1C",X"86",X"1E",
		X"75",X"20",X"BA",X"20",X"C0",X"1F",X"F5",X"1D",X"A2",X"1B",X"F9",X"18",X"1F",X"16",X"2A",X"13",
		X"2D",X"10",X"31",X"0D",X"3B",X"0A",X"56",X"07",X"7F",X"04",X"BC",X"01",X"0B",X"FF",X"6F",X"FC",
		X"E9",X"F9",X"78",X"F7",X"17",X"F5",X"CF",X"F2",X"96",X"F0",X"73",X"EE",X"61",X"EC",X"63",X"EA",
		X"73",X"E8",X"99",X"E6",X"C5",X"E4",X"43",X"E3",X"55",X"E3",X"B7",X"E4",X"EB",X"E6",X"AB",X"E9",
		X"BE",X"EC",X"04",X"F0",X"63",X"F3",X"C7",X"F6",X"28",X"FA",X"7D",X"FD",X"C1",X"00",X"F3",X"03",
		X"0E",X"07",X"13",X"0A",X"FE",X"0C",X"D4",X"0F",X"91",X"12",X"39",X"15",X"C8",X"17",X"44",X"1A",
		X"A6",X"1C",X"F5",X"1E",X"2F",X"21",X"58",X"23",X"6A",X"25",X"6C",X"27",X"59",X"29",X"37",X"2B",
		X"02",X"2D",X"BE",X"2E",X"67",X"30",X"03",X"32",X"8F",X"33",X"0B",X"35",X"7A",X"36",X"DB",X"37",
		X"2E",X"39",X"76",X"3A",X"B0",X"3B",X"DD",X"3C",X"FE",X"3D",X"16",X"3F",X"20",X"40",X"22",X"41",
		X"17",X"42",X"02",X"43",X"E6",X"43",X"BD",X"44",X"8C",X"45",X"54",X"46",X"11",X"47",X"C8",X"47",
		X"73",X"48",X"1B",X"49",X"99",X"49",X"A5",X"48",X"53",X"46",X"2F",X"43",X"79",X"3F",X"76",X"3B",
		X"3F",X"37",X"FA",X"32",X"AE",X"2E",X"6F",X"2A",X"3D",X"26",X"26",X"22",X"24",X"1E",X"41",X"1A",
		X"78",X"16",X"CC",X"12",X"3E",X"0F",X"CB",X"0B",X"74",X"08",X"39",X"05",X"1A",X"02",X"15",X"FF",
		X"28",X"FC",X"57",X"F9",X"9B",X"F6",X"F7",X"F3",X"69",X"F1",X"F3",X"EE",X"92",X"EC",X"44",X"EA",
		X"0C",X"E8",X"E8",X"E5",X"D5",X"E3",X"D7",X"E1",X"E8",X"DF",X"0C",X"DE",X"42",X"DC",X"84",X"DA",
		X"D9",X"D8",X"3D",X"D7",X"AE",X"D5",X"30",X"D4",X"BD",X"D2",X"5A",X"D1",X"03",X"D0",X"BA",X"CE",
		X"7B",X"CD",X"4A",X"CC",X"24",X"CB",X"09",X"CA",X"F9",X"C8",X"F4",X"C7",X"F9",X"C6",X"07",X"C6",
		X"21",X"C5",X"40",X"C4",X"6A",X"C3",X"9F",X"C2",X"DA",X"C1",X"1F",X"C1",X"6A",X"C0",X"BD",X"BF",
		X"1A",X"BF",X"7D",X"BE",X"E5",X"BD",X"56",X"BD",X"CC",X"BC",X"4B",X"BC",X"CE",X"BB",X"57",X"BB",
		X"E6",X"BA",X"7A",X"BA",X"15",X"BA",X"B5",X"B9",X"5A",X"B9",X"03",X"B9",X"B3",X"B8",X"65",X"B8",
		X"1D",X"B8",X"D8",X"B7",X"99",X"B7",X"5E",X"B7",X"25",X"B7",X"F2",X"B6",X"C2",X"B6",X"96",X"B6",
		X"6B",X"B6",X"47",X"B6",X"24",X"B6",X"06",X"B6",X"EA",X"B5",X"D0",X"B5",X"B9",X"B5",X"A8",X"B5",
		X"96",X"B5",X"89",X"B5",X"7E",X"B5",X"73",X"B5",X"6C",X"B5",X"68",X"B5",X"67",X"B5",X"65",X"B5",
		X"66",X"B5",X"6C",X"B5",X"6F",X"B5",X"78",X"B5",X"7F",X"B5",X"8E",X"B5",X"98",X"B5",X"AB",X"B5",
		X"B8",X"B5",X"E4",X"B6",X"97",X"B9",X"2B",X"BD",X"5D",X"C1",X"E2",X"C5",X"9E",X"CA",X"6B",X"CF",
		X"3C",X"D4",X"FF",X"D8",X"B0",X"DD",X"45",X"E2",X"C1",X"E6",X"19",X"EB",X"54",X"EF",X"6D",X"F3",
		X"69",X"F7",X"41",X"FB",X"FA",X"FE",X"92",X"02",X"0F",X"06",X"6D",X"09",X"B0",X"0C",X"D3",X"0F",
		X"DD",X"12",X"CD",X"15",X"A3",X"18",X"61",X"1B",X"06",X"1E",X"93",X"20",X"0A",X"23",X"6B",X"25",
		X"B6",X"27",X"ED",X"29",X"0E",X"2C",X"1E",X"2E",X"1A",X"30",X"04",X"32",X"DA",X"33",X"A4",X"35",
		X"57",X"37",X"FF",X"38",X"94",X"3A",X"1B",X"3C",X"93",X"3D",X"FF",X"3E",X"59",X"40",X"A9",X"41",
		X"E8",X"42",X"1F",X"44",X"45",X"45",X"66",X"46",X"72",X"47",X"7E",X"48",X"71",X"49",X"6D",X"4A",
		X"6E",X"4A",X"CF",X"48",X"3E",X"46",X"F9",X"42",X"52",X"3F",X"6D",X"3B",X"6A",X"37",X"5B",X"33",
		X"51",X"2F",X"52",X"2B",X"68",X"27",X"92",X"23",X"D8",X"1F",X"35",X"1C",X"AE",X"18",X"43",X"15",
		X"F3",X"11",X"BC",X"0E",X"A0",X"0B",X"9E",X"08",X"B6",X"05",X"E5",X"02",X"2C",X"00",X"8C",X"FD",
		X"FF",X"FA",X"8B",X"F8",X"26",X"F6",X"07",X"F4",X"71",X"F3",X"3C",X"F4",X"E4",X"F5",X"20",X"F8",
		X"B5",X"FA",X"83",X"FD",X"6A",X"00",X"60",X"03",X"54",X"06",X"42",X"09",X"21",X"0C",X"F1",X"0E",
		X"AD",X"11",X"57",X"14",X"EB",X"16",X"6B",X"19",X"D5",X"1B",X"2C",X"1E",X"6F",X"20",X"9C",X"22",
		X"B7",X"24",X"BE",X"26",X"B4",X"28",X"98",X"2A",X"69",X"2C",X"2B",X"2E",X"DC",X"2F",X"80",X"31",
		X"11",X"33",X"94",X"34",X"07",X"36",X"6F",X"37",X"C6",X"38",X"14",X"3A",X"52",X"3B",X"86",X"3C",
		X"AB",X"3D",X"C6",X"3E",X"D8",X"3F",X"DC",X"40",X"D4",X"41",X"C5",X"42",X"A9",X"43",X"84",X"44",
		X"54",X"45",X"1C",X"46",X"DB",X"46",X"8E",X"47",X"3D",X"48",X"E2",X"48",X"7D",X"49",X"15",X"4A",
		X"A1",X"4A",X"27",X"4B",X"A6",X"4B",X"1E",X"4C",X"91",X"4C",X"FB",X"4C",X"60",X"4D",X"BF",X"4D",
		X"19",X"4E",X"6B",X"4E",X"B9",X"4E",X"03",X"4F",X"45",X"4F",X"85",X"4F",X"BE",X"4F",X"F3",X"4F",
		X"24",X"50",X"4F",X"50",X"78",X"50",X"9B",X"50",X"BB",X"50",X"D6",X"50",X"F0",X"50",X"04",X"51",
		X"15",X"51",X"23",X"51",X"2C",X"51",X"35",X"51",X"39",X"51",X"3C",X"51",X"3A",X"51",X"35",X"51",
		X"2E",X"51",X"25",X"51",X"19",X"51",X"0A",X"51",X"FB",X"50",X"E7",X"50",X"D2",X"50",X"BD",X"50",
		X"A4",X"50",X"88",X"50",X"6B",X"50",X"4C",X"50",X"2D",X"50",X"0A",X"50",X"E7",X"4F",X"C1",X"4F",
		X"9A",X"4F",X"71",X"4F",X"48",X"4F",X"1C",X"4F",X"F0",X"4E",X"C3",X"4E",X"95",X"4E",X"65",X"4E",
		X"34",X"4E",X"FF",X"4D",X"CD",X"4D",X"99",X"4D",X"64",X"4D",X"2D",X"4D",X"F7",X"4C",X"BE",X"4C",
		X"86",X"4C",X"4C",X"4C",X"12",X"4C",X"D7",X"4B",X"9B",X"4B",X"5F",X"4B",X"22",X"4B",X"E3",X"4A",
		X"A5",X"4A",X"65",X"4A",X"27",X"4A",X"E5",X"49",X"A5",X"49",X"65",X"49",X"24",X"49",X"E3",X"48",
		X"A1",X"48",X"5C",X"48",X"1C",X"48",X"D4",X"47",X"9B",X"47",X"FE",X"46",X"D5",X"44",X"8B",X"41",
		X"8A",X"3D",X"19",X"39",X"68",X"34",X"97",X"2F",X"BE",X"2A",X"EB",X"25",X"2A",X"21",X"82",X"1C",
		X"F3",X"17",X"85",X"13",X"35",X"0F",X"06",X"0B",X"F7",X"06",X"09",X"03",X"3D",X"FF",X"90",X"FB",
		X"FE",X"F7",X"90",X"F4",X"3B",X"F1",X"06",X"EE",X"E7",X"EA",X"EB",X"E7",X"FD",X"E4",X"39",X"E2",
		X"7A",X"DF",X"D6",X"DD",X"C7",X"DD",X"AB",X"DE",X"42",X"E0",X"40",X"E2",X"87",X"E4",X"F0",X"E6",
		X"72",X"E9",X"F8",X"EB",X"7F",X"EE",X"FA",X"F0",X"6B",X"F3",X"CD",X"F5",X"1F",X"F8",X"5F",X"FA",
		X"8F",X"FC",X"AE",X"FE",X"B8",X"00",X"B2",X"02",X"9C",X"04",X"76",X"06",X"3D",X"08",X"F7",X"09",
		X"A0",X"0B",X"3C",X"0D",X"C4",X"0E",X"49",X"10",X"81",X"11",X"38",X"11",X"AF",X"0F",X"5F",X"0D",
		X"8A",X"0A",X"67",X"07",X"14",X"04",X"AE",X"00",X"43",X"FD",X"DD",X"F9",X"81",X"F6",X"3A",X"F3",
		X"05",X"F0",X"E9",X"EC",X"E1",X"E9",X"F2",X"E6",X"19",X"E4",X"5B",X"E1",X"B1",X"DE",X"20",X"DC",
		X"A6",X"D9",X"40",X"D7",X"F0",X"D4",X"B5",X"D2",X"8C",X"D0",X"7B",X"CE",X"76",X"CC",X"AB",X"CA",
		X"4C",X"CA",X"44",X"CB",X"0A",X"CD",X"63",X"CF",X"0F",X"D2",X"F1",X"D4",X"ED",X"D7",X"F5",X"DA",
		X"F9",X"DD",X"F9",X"E0",X"E7",X"E3",X"C8",X"E6",X"93",X"E9",X"4C",X"EC",X"EF",X"EE",X"80",X"F1",
		X"F8",X"F3",X"5F",X"F6",X"B0",X"F8",X"EE",X"FA",X"19",X"FD",X"32",X"FF",X"36",X"01",X"2B",X"03",
		X"0E",X"05",X"E1",X"06",X"A1",X"08",X"54",X"0A",X"F6",X"0B",X"8A",X"0D",X"0F",X"0F",X"88",X"10",
		X"F1",X"11",X"4E",X"13",X"9D",X"14",X"E2",X"15",X"1B",X"17",X"47",X"18",X"67",X"19",X"7E",X"1A",
		X"8A",X"1B",X"8B",X"1C",X"81",X"1D",X"71",X"1E",X"54",X"1F",X"2F",X"20",X"03",X"21",X"CD",X"21",
		X"8D",X"22",X"47",X"23",X"FB",X"23",X"A8",X"24",X"48",X"25",X"E5",X"25",X"7A",X"26",X"09",X"27",
		X"90",X"27",X"15",X"28",X"90",X"28",X"08",X"29",X"78",X"29",X"E3",X"29",X"48",X"2A",X"AC",X"2A",
		X"04",X"2B",X"5E",X"2B",X"B0",X"2B",X"FF",X"2B",X"46",X"2C",X"8C",X"2C",X"CE",X"2C",X"0C",X"2D",
		X"43",X"2D",X"7B",X"2D",X"AB",X"2D",X"DB",X"2D",X"05",X"2E",X"2F",X"2E",X"50",X"2E",X"76",X"2E",
		X"8E",X"2E",X"B7",X"2E",X"60",X"2E",X"89",X"2C",X"A9",X"29",X"1D",X"26",X"29",X"22",X"F9",X"1D",
		X"AD",X"19",X"54",X"15",X"02",X"11",X"C0",X"0C",X"93",X"08",X"7F",X"04",X"87",X"00",X"AC",X"FC",
		X"ED",X"F8",X"4B",X"F5",X"C9",X"F1",X"61",X"EE",X"1A",X"EB",X"EB",X"E7",X"DA",X"E4",X"E1",X"E1",
		X"06",X"DF",X"3F",X"DC",X"95",X"D9",X"FE",X"D6",X"85",X"D4",X"1B",X"D2",X"D8",X"D0",X"0C",X"D1",
		X"20",X"D2",X"D8",X"D3",X"EB",X"D5",X"42",X"D8",X"B8",X"DA",X"43",X"DD",X"CF",X"DF",X"5A",X"E2",
		X"DC",X"E4",X"4E",X"E7",X"B6",X"E9",X"0B",X"EC",X"50",X"EE",X"81",X"F0",X"A5",X"F2",X"B3",X"F4",
		X"B3",X"F6",X"9F",X"F8",X"7D",X"FA",X"4A",X"FC",X"08",X"FE",X"B5",X"FF",X"57",X"01",X"E4",X"02",
		X"70",X"04",X"9C",X"05",X"4A",X"05",X"D8",X"03",X"AA",X"01",X"04",X"FF",X"15",X"FC",X"FD",X"F8",
		X"D0",X"F5",X"A0",X"F2",X"75",X"EF",X"58",X"EC",X"48",X"E9",X"4E",X"E6",X"66",X"E3",X"96",X"E0",
		X"DC",X"DD",X"3A",X"DB",X"AC",X"D8",X"35",X"D6",X"D2",X"D3",X"87",X"D1",X"4E",X"CF",X"2C",X"CD",
		X"19",X"CB",X"1F",X"C9",X"30",X"C7",X"5A",X"C5",X"8A",X"C3",X"AA",X"C2",X"49",X"C3",X"CB",X"C4",
		X"F4",X"C6",X"77",X"C9",X"3D",X"CC",X"21",X"CF",X"18",X"D2",X"0B",X"D5",X"FE",X"D7",X"E2",X"DA",
		X"B8",X"DD",X"7C",X"E0",X"2B",X"E3",X"C8",X"E5",X"52",X"E8",X"C7",X"EA",X"27",X"ED",X"74",X"EF",
		X"AF",X"F1",X"D5",X"F3",X"EB",X"F5",X"EC",X"F7",X"DE",X"F9",X"BF",X"FB",X"90",X"FD",X"4F",X"FF",
		X"01",X"01",X"A1",X"02",X"35",X"04",X"BC",X"05",X"34",X"07",X"9D",X"08",X"FC",X"09",X"4B",X"0B",
		X"90",X"0C",X"C9",X"0D",X"F8",X"0E",X"1A",X"10",X"33",X"11",X"41",X"12",X"45",X"13",X"3F",X"14",
		X"30",X"15",X"17",X"16",X"F7",X"16",X"CC",X"17",X"99",X"18",X"5F",X"19",X"1D",X"1A",X"D3",X"1A",
		X"82",X"1B",X"2A",X"1C",X"C9",X"1C",X"65",X"1D",X"F9",X"1D",X"86",X"1E",X"0E",X"1F",X"8F",X"1F",
		X"0A",X"20",X"80",X"20",X"F1",X"20",X"5C",X"21",X"C3",X"21",X"23",X"22",X"80",X"22",X"D9",X"22",
		X"2D",X"23",X"7B",X"23",X"C7",X"23",X"0E",X"24",X"52",X"24",X"91",X"24",X"CD",X"24",X"05",X"25",
		X"39",X"25",X"6B",X"25",X"9B",X"25",X"C5",X"25",X"EE",X"25",X"11",X"26",X"34",X"26",X"54",X"26",
		X"71",X"26",X"8B",X"26",X"A4",X"26",X"B9",X"26",X"CE",X"26",X"DB",X"26",X"EC",X"26",X"F7",X"26",
		X"01",X"27",X"0A",X"27",X"11",X"27",X"15",X"27",X"19",X"27",X"19",X"27",X"1B",X"27",X"18",X"27",
		X"15",X"27",X"0E",X"27",X"09",X"27",X"FF",X"26",X"F8",X"26",X"EA",X"26",X"E1",X"26",X"D1",X"26",
		X"C7",X"26",X"B1",X"26",X"AC",X"26",X"20",X"26",X"22",X"24",X"3E",X"21",X"AB",X"1D",X"F8",X"19",
		X"EB",X"15",X"A4",X"11",X"62",X"0D",X"21",X"09",X"F4",X"04",X"D9",X"00",X"DB",X"FC",X"F5",X"F8",
		X"2E",X"F5",X"81",X"F1",X"F5",X"ED",X"86",X"EA",X"32",X"E7",X"FB",X"E3",X"E0",X"E0",X"E1",X"DD",
		X"F9",X"DA",X"2D",X"D8",X"78",X"D5",X"DD",X"D2",X"58",X"D0",X"EB",X"CD",X"99",X"CB",X"70",X"CA",
		X"A6",X"CA",X"AE",X"CB",X"50",X"CD",X"47",X"CF",X"7E",X"D1",X"CF",X"D3",X"36",X"D6",X"9E",X"D8",
		X"05",X"DB",X"61",X"DD",X"B4",X"DF",X"F7",X"E1",X"2D",X"E4",X"50",X"E6",X"66",X"E8",X"68",X"EA",
		X"5D",X"EC",X"40",X"EE",X"16",X"F0",X"D8",X"F1",X"8F",X"F3",X"35",X"F5",X"D0",X"F6",X"59",X"F8",
		X"D7",X"F9",X"48",X"FB",X"AB",X"FC",X"01",X"FE",X"4E",X"FF",X"8C",X"00",X"C1",X"01",X"EA",X"02",
		X"0A",X"04",X"1E",X"05",X"2A",X"06",X"2A",X"07",X"23",X"08",X"12",X"09",X"F8",X"09",X"D6",X"0A",
		X"AD",X"0B",X"7A",X"0C",X"40",X"0D",X"FE",X"0D",X"B5",X"0E",X"66",X"0F",X"0F",X"10",X"B1",X"10",
		X"4E",X"11",X"E3",X"11",X"72",X"12",X"FD",X"12",X"81",X"13",X"FF",X"13",X"79",X"14",X"EE",X"14",
		X"5D",X"15",X"C8",X"15",X"2D",X"16",X"8E",X"16",X"EB",X"16",X"44",X"17",X"99",X"17",X"E9",X"17",
		X"35",X"18",X"7D",X"18",X"C3",X"18",X"04",X"19",X"44",X"19",X"7D",X"19",X"B5",X"19",X"E9",X"19",
		X"1B",X"1A",X"49",X"1A",X"76",X"1A",X"9D",X"1A",X"C6",X"1A",X"E9",X"1A",X"0B",X"1B",X"27",X"1B",
		X"4B",X"1B",X"2D",X"1B",X"BD",X"19",X"3A",X"17",X"10",X"14",X"77",X"10",X"A2",X"0C",X"AD",X"08",
		X"AD",X"04",X"B0",X"00",X"C1",X"FC",X"E3",X"F8",X"1E",X"F5",X"71",X"F1",X"DE",X"ED",X"68",X"EA",
		X"0F",X"E7",X"CD",X"E3",X"AA",X"E0",X"A1",X"DD",X"B1",X"DA",X"DC",X"D7",X"20",X"D5",X"7A",X"D2",
		X"ED",X"CF",X"79",X"CD",X"19",X"CB",X"D0",X"C8",X"9A",X"C6",X"7A",X"C4",X"6D",X"C2",X"72",X"C0",
		X"8B",X"BE",X"B5",X"BC",X"F1",X"BA",X"3F",X"B9",X"9C",X"B7",X"08",X"B6",X"85",X"B4",X"0F",X"B3",
		X"A9",X"B1",X"50",X"B0",X"05",X"AF",X"C7",X"AD",X"97",X"AC",X"73",X"AB",X"5B",X"AA",X"4D",X"A9",
		X"4C",X"A8",X"54",X"A7",X"68",X"A6",X"88",X"A5",X"AF",X"A4",X"E1",X"A3",X"1C",X"A3",X"5F",X"A2",
		X"AD",X"A1",X"02",X"A1",X"5F",X"A0",X"C6",X"9F",X"32",X"9F",X"A6",X"9E",X"23",X"9E",X"A6",X"9D",
		X"2E",X"9D",X"C0",X"9C",X"57",X"9C",X"F4",X"9B",X"98",X"9B",X"40",X"9B",X"ED",X"9A",X"A1",X"9A",
		X"59",X"9A",X"1A",X"9A",X"DD",X"99",X"A3",X"99",X"70",X"99",X"41",X"99",X"18",X"99",X"F0",X"98",
		X"CF",X"98",X"B0",X"98",X"96",X"98",X"8D",X"98",X"A4",X"99",X"F1",X"9B",X"EE",X"9E",X"68",X"A2",
		X"22",X"A6",X"08",X"AA",X"FA",X"AD",X"EF",X"B1",X"D7",X"B5",X"B3",X"B9",X"77",X"BD",X"25",X"C1",
		X"B8",X"C4",X"35",X"C8",X"96",X"CB",X"DC",X"CE",X"0A",X"D2",X"1D",X"D5",X"17",X"D8",X"FA",X"DA",
		X"C4",X"DD",X"78",X"E0",X"13",X"E3",X"9A",X"E5",X"0B",X"E8",X"68",X"EA",X"B2",X"EC",X"E6",X"EE",
		X"0B",X"F1",X"1C",X"F3",X"18",X"F5",X"06",X"F7",X"E2",X"F8",X"B1",X"FA",X"6D",X"FC",X"1C",X"FE",
		X"BA",X"FF",X"49",X"01",X"CD",X"02",X"42",X"04",X"AB",X"05",X"04",X"07",X"57",X"08",X"99",X"09",
		X"D3",X"0A",X"FD",X"0B",X"21",X"0D",X"38",X"0E",X"46",X"0F",X"48",X"10",X"44",X"11",X"32",X"12",
		X"1C",X"13",X"F7",X"13",X"CE",X"14",X"A2",X"14",X"33",X"13",X"06",X"11",X"55",X"0E",X"58",X"0B",
		X"2B",X"08",X"ED",X"04",X"A5",X"01",X"64",X"FE",X"2F",X"FB",X"09",X"F8",X"F6",X"F4",X"FA",X"F1",
		X"12",X"EF",X"42",X"EC",X"88",X"E9",X"E6",X"E6",X"59",X"E4",X"E1",X"E1",X"81",X"DF",X"33",X"DD",
		X"FC",X"DA",X"D6",X"D8",X"C7",X"D6",X"C7",X"D4",X"DE",X"D2",X"FA",X"D0",X"79",X"CF",X"52",X"CF",
		X"31",X"D0",X"BB",X"D1",X"B5",X"D3",X"F5",X"D5",X"5C",X"D8",X"D7",X"DA",X"5A",X"DD",X"DD",X"DF",
		X"58",X"E2",X"C7",X"E4",X"28",X"E7",X"7A",X"E9",X"BB",X"EB",X"EC",X"ED",X"0B",X"F0",X"19",X"F2",
		X"16",X"F4",X"04",X"F6",X"E0",X"F7",X"AD",X"F9",X"69",X"FB",X"18",X"FD",X"B5",X"FE",X"49",X"00",
		X"C6",X"01",X"44",X"03",X"E3",X"03",X"30",X"03",X"B5",X"01",X"AA",X"FF",X"4E",X"FD",X"B7",X"FA",
		X"0A",X"F8",X"4E",X"F5",X"96",X"F2",X"DE",X"EF",X"38",X"ED",X"9F",X"EA",X"19",X"E8",X"A3",X"E5",
		X"44",X"E3",X"F3",X"E0",X"B9",X"DE",X"8F",X"DC",X"7B",X"DA",X"76",X"D8",X"87",X"D6",X"A6",X"D4",
		X"D9",X"D2",X"1B",X"D1",X"6C",X"CF",X"CB",X"CD",X"3E",X"CC",X"BE",X"CA",X"4B",X"C9",X"E8",X"C7",
		X"90",X"C6",X"45",X"C5",X"07",X"C4",X"D7",X"C2",X"B0",X"C1",X"96",X"C0",X"87",X"BF",X"84",X"BE",
		X"88",X"BD",X"9B",X"BC",X"B2",X"BB",X"D9",X"BA",X"05",X"BA",X"3C",X"B9",X"78",X"B8",X"C0",X"B7",
		X"0E",X"B7",X"67",X"B6",X"C4",X"B5",X"2D",X"B5",X"97",X"B4",X"10",X"B4",X"85",X"B3",X"0E",X"B3",
		X"8A",X"B2",X"B6",X"B2",X"2E",X"B4",X"76",X"B6",X"4B",X"B9",X"6F",X"BC",X"CA",X"BF",X"38",X"C3",
		X"B0",X"C6",X"25",X"CA",X"8E",X"CD",X"E3",X"D0",X"29",X"D4",X"58",X"D7",X"71",X"DA",X"72",X"DD",
		X"5C",X"E0",X"2F",X"E3",X"EB",X"E5",X"93",X"E8",X"23",X"EB",X"9C",X"ED",X"03",X"F0",X"53",X"F2",
		X"92",X"F4",X"BD",X"F6",X"D3",X"F8",X"DA",X"FA",X"B9",X"FC",X"6C",X"FD",X"F8",X"FC",X"D3",X"FB",
		X"31",X"FA",X"45",X"F8",X"27",X"F6",X"F3",X"F3",X"B4",X"F1",X"74",X"EF",X"38",X"ED",X"07",X"EB",
		X"E2",X"E8",X"CB",X"E6",X"C2",X"E4",X"CB",X"E2",X"E2",X"E0",X"0A",X"DF",X"44",X"DD",X"89",X"DB",
		X"E3",X"D9",X"46",X"D8",X"BE",X"D6",X"3D",X"D5",X"D1",X"D3",X"6C",X"D2",X"1C",X"D1",X"C8",X"CF",
		X"01",X"CF",X"8D",X"CF",X"F5",X"D0",X"F6",X"D2",X"52",X"D5",X"EB",X"D7",X"9F",X"DA",X"66",X"DD",
		X"2C",X"E0",X"EE",X"E2",X"A3",X"E5",X"4B",X"E8",X"E3",X"EA",X"67",X"ED",X"DA",X"EF",X"3B",X"F2",
		X"86",X"F4",X"C1",X"F6",X"E6",X"F8",X"FD",X"FA",X"FF",X"FC",X"F4",X"FE",X"D3",X"00",X"A7",X"02",
		X"66",X"04",X"19",X"06",X"B9",X"07",X"47",X"09",X"CD",X"09",X"21",X"09",X"C2",X"07",X"E1",X"05",
		X"BD",X"03",X"60",X"01",X"E9",X"FE",X"66",X"FC",X"E4",X"F9",X"67",X"F7",X"F7",X"F4",X"94",X"F2",
		X"41",X"F0",X"FF",X"ED",X"CD",X"EB",X"AF",X"E9",X"A1",X"E7",X"A4",X"E5",X"B9",X"E3",X"DF",X"E1",
		X"15",X"E0",X"5C",X"DE",X"B1",X"DC",X"18",X"DB",X"87",X"D9",X"0F",X"D8",X"94",X"D6",X"84",X"D5",
		X"C3",X"D5",X"EE",X"D6",X"B7",X"D8",X"E4",X"DA",X"50",X"DD",X"DD",X"DF",X"7E",X"E2",X"1F",X"E5",
		X"BE",X"E7",X"55",X"EA",X"DD",X"EC",X"56",X"EF",X"BF",X"F1",X"15",X"F4",X"5B",X"F6",X"8F",X"F8",
		X"AE",X"FA",X"BD",X"FC",X"BB",X"FE",X"A7",X"00",X"83",X"02",X"4E",X"04",X"0B",X"06",X"B8",X"07",
		X"55",X"09",X"E4",X"0A",X"65",X"0C",X"DB",X"0D",X"41",X"0F",X"9B",X"10",X"E8",X"11",X"2B",X"13",
		X"5F",X"14",X"8B",X"15",X"A9",X"16",X"C2",X"17",X"CA",X"18",X"CC",X"19",X"C4",X"1A",X"B3",X"1B",
		X"96",X"1C",X"73",X"1D",X"45",X"1E",X"12",X"1F",X"D4",X"1F",X"90",X"20",X"44",X"21",X"F1",X"21",
		X"96",X"22",X"36",X"23",X"CC",X"23",X"60",X"24",X"E8",X"24",X"76",X"25",X"BE",X"25",X"D1",X"24",
		X"F0",X"22",X"72",X"20",X"95",X"1D",X"7C",X"1A",X"43",X"17",X"00",X"14",X"BC",X"10",X"81",X"0D",
		X"52",X"0A",X"39",X"07",X"31",X"04",X"40",X"01",X"65",X"FE",X"9E",X"FB",X"F0",X"F8",X"57",X"F6",
		X"D4",X"F3",X"64",X"F1",X"0D",X"EF",X"C9",X"EC",X"99",X"EA",X"79",X"E8",X"71",X"E6",X"74",X"E4",
		X"92",X"E2",X"B2",X"E0",X"96",X"DF",X"C0",X"DF",X"AF",X"E0",X"2F",X"E2",X"FE",X"E3",X"0B",X"E6",
		X"32",X"E8",X"6B",X"EA",X"A5",X"EC",X"E0",X"EE",X"10",X"F1",X"37",X"F3",X"4D",X"F5",X"58",X"F7",
		X"53",X"F9",X"41",X"FB",X"1B",X"FD",X"E8",X"FE",X"A5",X"00",X"55",X"02",X"F5",X"03",X"88",X"05",
		X"0B",X"07",X"83",X"08",X"ED",X"09",X"4B",X"0B",X"9C",X"0C",X"E0",X"0D",X"1A",X"0F",X"48",X"10",
		X"6D",X"11",X"85",X"12",X"94",X"13",X"98",X"14",X"93",X"15",X"84",X"16",X"6D",X"17",X"4D",X"18",
		X"25",X"19",X"F4",X"19",X"BB",X"1A",X"7A",X"1B",X"33",X"1C",X"E1",X"1C",X"8C",X"1D",X"2D",X"1E",
		X"CB",X"1E",X"5E",X"1F",X"F0",X"1F",X"76",X"20",X"FC",X"20",X"76",X"21",X"F3",X"21",X"60",X"22",
		X"D9",X"22",X"C0",X"22",X"6C",X"21",X"51",X"1F",X"AF",X"1C",X"C1",X"19",X"A0",X"16",X"69",X"13",
		X"29",X"10",X"EF",X"0C",X"BF",X"09",X"A0",X"06",X"91",X"03",X"98",X"00",X"B6",X"FD",X"EA",X"FA",
		X"32",X"F8",X"90",X"F5",X"06",X"F3",X"91",X"F0",X"2F",X"EE",X"E3",X"EB",X"AB",X"E9",X"87",X"E7",
		X"75",X"E5",X"76",X"E3",X"88",X"E1",X"AC",X"DF",X"E0",X"DD",X"23",X"DC",X"77",X"DA",X"DB",X"D8",
		X"4C",X"D7",X"CE",X"D5",X"5D",X"D4",X"F9",X"D2",X"A3",X"D1",X"59",X"D0",X"1C",X"CF",X"EC",X"CD",
		X"C4",X"CC",X"AA",X"CB",X"99",X"CA",X"95",X"C9",X"98",X"C8",X"A8",X"C7",X"C0",X"C6",X"E2",X"C5",
		X"0D",X"C5",X"42",X"C4",X"7D",X"C3",X"BF",X"C2",X"0E",X"C2",X"60",X"C1",X"BB",X"C0",X"1D",X"C0",
		X"88",X"BF",X"F9",X"BE",X"6F",X"BE",X"EC",X"BD",X"70",X"BD",X"FB",X"BC",X"8A",X"BC",X"1F",X"BC",
		X"B9",X"BB",X"5A",X"BB",X"FE",X"BA",X"A9",X"BA",X"59",X"BA",X"0B",X"BA",X"C3",X"B9",X"80",X"B9",
		X"40",X"B9",X"06",X"B9",X"CE",X"B8",X"9B",X"B8",X"6A",X"B8",X"3E",X"B8",X"14",X"B8",X"F1",X"B7",
		X"CC",X"B7",X"B2",X"B7",X"8D",X"B7",X"B9",X"B7",X"11",X"B9",X"44",X"BB",X"05",X"BE",X"1B",X"C1",
		X"65",X"C4",X"CA",X"C7",X"33",X"CB",X"9E",X"CE",X"FA",X"D1",X"49",X"D5",X"85",X"D8",X"AA",X"DB",
		X"B9",X"DE",X"B3",X"E1",X"97",X"E4",X"5F",X"E7",X"15",X"EA",X"B3",X"EC",X"3B",X"EF",X"AE",X"F1",
		X"0E",X"F4",X"58",X"F6",X"90",X"F8",X"B2",X"FA",X"C8",X"FC",X"C2",X"FE",X"B7",X"00",X"D9",X"01",
		X"CB",X"01",X"07",X"01",X"BE",X"FF",X"2B",X"FE",X"5F",X"FC",X"7B",X"FA",X"85",X"F8",X"8D",X"F6",
		X"96",X"F4",X"A7",X"F2",X"C2",X"F0",X"E9",X"EE",X"1A",X"ED",X"5E",X"EB",X"AD",X"E9",X"0A",X"E8",
		X"74",X"E6",X"ED",X"E4",X"73",X"E3",X"08",X"E2",X"A7",X"E0",X"53",X"DF",X"0C",X"DE",X"D2",X"DC",
		X"A2",X"DB",X"7D",X"DA",X"63",X"D9",X"53",X"D8",X"4F",X"D7",X"53",X"D6",X"61",X"D5",X"78",X"D4",
		X"99",X"D3",X"C3",X"D2",X"F5",X"D1",X"2F",X"D1",X"71",X"D0",X"BB",X"CF",X"0D",X"CF",X"64",X"CE",
		X"C3",X"CD",X"29",X"CD",X"97",X"CC",X"09",X"CC",X"84",X"CB",X"03",X"CB",X"89",X"CA",X"12",X"CA",
		X"A3",X"C9",X"36",X"C9",X"D5",X"C8",X"70",X"C8",X"1B",X"C8",X"B9",X"C7",X"FA",X"C7",X"63",X"C9",
		X"7D",X"CB",X"19",X"CE",X"F7",X"D0",X"04",X"D4",X"22",X"D7",X"48",X"DA",X"69",X"DD",X"7F",X"E0",
		X"85",X"E3",X"7A",X"E6",X"5A",X"E9",X"26",X"EC",X"DB",X"EE",X"7D",X"F1",X"09",X"F4",X"81",X"F6",
		X"E3",X"F8",X"32",X"FB",X"6D",X"FD",X"93",X"FF",X"A9",X"01",X"AC",X"03",X"9D",X"05",X"7E",X"07",
		X"4E",X"09",X"0F",X"0B",X"BE",X"0C",X"60",X"0E",X"F3",X"0F",X"77",X"11",X"EF",X"12",X"59",X"14",
		X"B5",X"15",X"05",X"17",X"4A",X"18",X"81",X"19",X"AD",X"1A",X"D0",X"1B",X"E8",X"1C",X"F4",X"1D",
		X"F8",X"1E",X"EF",X"1F",X"E0",X"20",X"C5",X"21",X"A2",X"22",X"77",X"23",X"43",X"24",X"07",X"25",
		X"C3",X"25",X"77",X"26",X"25",X"27",X"CA",X"27",X"69",X"28",X"02",X"29",X"95",X"29",X"1F",X"2A",
		X"A6",X"2A",X"23",X"2B",X"9D",X"2B",X"10",X"2C",X"80",X"2C",X"EA",X"2C",X"4E",X"2D",X"AE",X"2D",
		X"09",X"2E",X"60",X"2E",X"B1",X"2E",X"FD",X"2E",X"46",X"2F",X"8B",X"2F",X"CD",X"2F",X"09",X"30",
		X"43",X"30",X"78",X"30",X"AB",X"30",X"DB",X"30",X"08",X"31",X"30",X"31",X"54",X"31",X"78",X"31",
		X"98",X"31",X"B5",X"31",X"D1",X"31",X"E8",X"31",X"FE",X"31",X"11",X"32",X"20",X"32",X"30",X"32",
		X"3B",X"32",X"46",X"32",X"4D",X"32",X"54",X"32",X"57",X"32",X"5C",X"32",X"5B",X"32",X"5B",X"32",
		X"56",X"32",X"54",X"32",X"4B",X"32",X"45",X"32",X"3B",X"32",X"32",X"32",X"24",X"32",X"18",X"32",
		X"07",X"32",X"FC",X"31",X"E5",X"31",X"DE",X"31",X"7A",X"31",X"FE",X"2F",X"B8",X"2D",X"F9",X"2A",
		X"DC",X"27",X"E3",X"24",X"AF",X"21",X"41",X"1E",X"EC",X"1A",X"94",X"17",X"57",X"14",X"27",X"11",
		X"12",X"0E",X"0F",X"0B",X"27",X"08",X"51",X"05",X"97",X"02",X"ED",X"FF",X"60",X"FD",X"E3",X"FA",
		X"7D",X"F8",X"2C",X"F6",X"EF",X"F3",X"C4",X"F1",X"AD",X"EF",X"A9",X"ED",X"B5",X"EB",X"D5",X"E9",
		X"03",X"E8",X"41",X"E6",X"90",X"E4",X"EE",X"E2",X"5B",X"E1",X"D5",X"DF",X"5F",X"DE",X"F5",X"DC",
		X"98",X"DB",X"49",X"DA",X"05",X"D9",X"CC",X"D7",X"A1",X"D6",X"80",X"D5",X"69",X"D4",X"5D",X"D3",
		X"5C",X"D2",X"64",X"D1",X"77",X"D0",X"93",X"CF",X"B5",X"CE",X"E3",X"CD",X"18",X"CD",X"57",X"CC",
		X"9A",X"CB",X"EB",X"CA",X"39",X"CA",X"C9",X"C9",X"71",X"CA",X"F3",X"CB",X"FF",X"CD",X"64",X"D0",
		X"FC",X"D2",X"B2",X"D5",X"74",X"D8",X"37",X"DB",X"F4",X"DD",X"A7",X"E0",X"4B",X"E3",X"DE",X"E5",
		X"5C",X"E8",X"CD",X"EA",X"28",X"ED",X"72",X"EF",X"A9",X"F1",X"CF",X"F3",X"E1",X"F5",X"E2",X"F7",
		X"D2",X"F9",X"B2",X"FB",X"82",X"FD",X"42",X"FF",X"F1",X"00",X"94",X"02",X"28",X"04",X"AE",X"05",
		X"26",X"07",X"93",X"08",X"F0",X"09",X"44",X"0B",X"8A",X"0C",X"C6",X"0D",X"F5",X"0E",X"1B",X"10",
		X"35",X"11",X"46",X"12",X"4B",X"13",X"49",X"14",X"3B",X"15",X"27",X"16",X"08",X"17",X"E2",X"17",
		X"B2",X"18",X"7B",X"19",X"3C",X"1A",X"F7",X"1A",X"A9",X"1B",X"54",X"1C",X"F8",X"1C",X"97",X"1D",
		X"2E",X"1E",X"C2",X"1E",X"2F",X"1F",X"99",X"1E",X"1D",X"1D",X"18",X"1B",X"B3",X"18",X"1A",X"16",
		X"5F",X"13",X"9C",X"10",X"D4",X"0D",X"16",X"0B",X"61",X"08",X"BB",X"05",X"24",X"03",X"A2",X"00",
		X"32",X"FE",X"D6",X"FB",X"8B",X"F9",X"53",X"F7",X"2F",X"F5",X"1D",X"F3",X"1C",X"F1",X"2B",X"EF",
		X"4D",X"ED",X"7E",X"EB",X"C1",X"E9",X"11",X"E8",X"72",X"E6",X"E2",X"E4",X"5D",X"E3",X"E9",X"E1",
		X"80",X"E0",X"26",X"DF",X"D7",X"DD",X"94",X"DC",X"5D",X"DB",X"34",X"DA",X"13",X"D9",X"FD",X"D7",
		X"F3",X"D6",X"F2",X"D5",X"FB",X"D4",X"0B",X"D4",X"27",X"D3",X"4C",X"D2",X"79",X"D1",X"AF",X"D0",
		X"EC",X"CF",X"31",X"CF",X"7F",X"CE",X"D3",X"CD",X"2E",X"CD",X"93",X"CC",X"FB",X"CB",X"6B",X"CB",
		X"E0",X"CA",X"5D",X"CA",X"DF",X"C9",X"66",X"C9",X"F4",X"C8",X"85",X"C8",X"1E",X"C8",X"BA",X"C7",
		X"5E",X"C7",X"05",X"C7",X"B0",X"C6",X"61",X"C6",X"15",X"C6",X"CE",X"C5",X"8A",X"C5",X"49",X"C5",
		X"0E",X"C5",X"D5",X"C4",X"A0",X"C4",X"71",X"C4",X"41",X"C4",X"17",X"C4",X"F1",X"C3",X"CB",X"C3",
		X"AA",X"C3",X"8E",X"C3",X"71",X"C3",X"59",X"C3",X"42",X"C3",X"2D",X"C3",X"1D",X"C3",X"0D",X"C3",
		X"FF",X"C2",X"F7",X"C2",X"ED",X"C2",X"E7",X"C2",X"E0",X"C2",X"DF",X"C2",X"DE",X"C2",X"DF",X"C2",
		X"E2",X"C2",X"E7",X"C2",X"ED",X"C2",X"F5",X"C2",X"FD",X"C2",X"06",X"C3",X"15",X"C3",X"22",X"C3",
		X"2F",X"C3",X"40",X"C3",X"51",X"C3",X"63",X"C3",X"78",X"C3",X"8C",X"C3",X"A0",X"C3",X"B8",X"C3",
		X"D1",X"C3",X"E8",X"C3",X"01",X"C4",X"1D",X"C4",X"38",X"C4",X"54",X"C4",X"71",X"C4",X"90",X"C4",
		X"AE",X"C4",X"CD",X"C4",X"ED",X"C4",X"0D",X"C5",X"2E",X"C5",X"51",X"C5",X"74",X"C5",X"95",X"C5",
		X"BA",X"C5",X"DD",X"C5",X"03",X"C6",X"28",X"C6",X"4E",X"C6",X"72",X"C6",X"9A",X"C6",X"BF",X"C6",
		X"E9",X"C6",X"0E",X"C7",X"3A",X"C7",X"5E",X"C7",X"31",X"C8",X"05",X"CA",X"6C",X"CC",X"39",X"CF",
		X"3B",X"D2",X"63",X"D5",X"92",X"D8",X"C5",X"DB",X"F0",X"DE",X"0D",X"E2",X"18",X"E5",X"11",X"E8",
		X"F5",X"EA",X"C4",X"ED",X"7C",X"F0",X"1F",X"F3",X"AC",X"F5",X"24",X"F8",X"89",X"FA",X"D7",X"FC",
		X"14",X"FF",X"3C",X"01",X"55",X"03",X"58",X"05",X"4C",X"07",X"2D",X"09",X"02",X"0B",X"98",X"0C",
		X"27",X"0D",X"DA",X"0C",X"05",X"0C",X"D2",X"0A",X"65",X"09",X"D4",X"07",X"30",X"06",X"84",X"04",
		X"D6",X"02",X"2A",X"01",X"87",X"FF",X"EB",X"FD",X"5A",X"FC",X"D3",X"FA",X"59",X"F9",X"EB",X"F7",
		X"89",X"F6",X"32",X"F5",X"E5",X"F3",X"A7",X"F2",X"70",X"F1",X"46",X"F0",X"22",X"EF",X"0F",X"EE",
		X"00",X"ED",X"01",X"EC",X"00",X"EB",X"96",X"EA",X"39",X"EB",X"7C",X"EC",X"32",X"EE",X"2B",X"F0",
		X"50",X"F2",X"87",X"F4",X"CB",X"F6",X"0A",X"F9",X"46",X"FB",X"77",X"FD",X"9D",X"FF",X"B2",X"01",
		X"BB",X"03",X"B2",X"05",X"9C",X"07",X"74",X"09",X"3E",X"0B",X"F7",X"0C",X"A2",X"0E",X"3F",X"10",
		X"CE",X"11",X"4B",X"13",X"C0",X"14",X"25",X"16",X"7D",X"17",X"CA",X"18",X"0B",X"1A",X"40",X"1B",
		X"69",X"1C",X"88",X"1D",X"9B",X"1E",X"A6",X"1F",X"A5",X"20",X"9B",X"21",X"87",X"22",X"6C",X"23",
		X"45",X"24",X"19",X"25",X"E3",X"25",X"A5",X"26",X"5F",X"27",X"12",X"28",X"BC",X"28",X"61",X"29",
		X"FF",X"29",X"97",X"2A",X"26",X"2B",X"B0",X"2B",X"33",X"2C",X"B3",X"2C",X"29",X"2D",X"9F",X"2D",
		X"07",X"2E",X"7B",X"2E",X"76",X"2E",X"6C",X"2D",X"BC",X"2B",X"9A",X"29",X"34",X"27",X"A6",X"24",
		X"04",X"22",X"5A",X"1F",X"B4",X"1C",X"14",X"1A",X"84",X"17",X"00",X"15",X"8E",X"12",X"2A",X"10",
		X"DD",X"0D",X"9D",X"0B",X"72",X"09",X"58",X"07",X"50",X"05",X"56",X"03",X"70",X"01",X"99",X"FF",
		X"D2",X"FD",X"18",X"FC",X"70",X"FA",X"D3",X"F8",X"48",X"F7",X"D1",X"F5",X"37",X"F5",X"88",X"F5",
		X"68",X"F6",X"AD",X"F7",X"2D",X"F9",X"D5",X"FA",X"8E",X"FC",X"54",X"FE",X"19",X"00",X"DB",X"01",
		X"95",X"03",X"45",X"05",X"EB",X"06",X"84",X"08",X"13",X"0A",X"92",X"0B",X"08",X"0D",X"70",X"0E",
		X"CD",X"0F",X"1B",X"11",X"5F",X"12",X"97",X"13",X"C7",X"14",X"E8",X"15",X"02",X"17",X"0D",X"18",
		X"19",X"19",X"CA",X"19",X"76",X"19",X"6D",X"18",X"EA",X"16",X"1E",X"15",X"22",X"13",X"0C",X"11",
		X"EC",X"0E",X"C9",X"0C",X"A8",X"0A",X"91",X"08",X"83",X"06",X"83",X"04",X"93",X"02",X"AE",X"00",
		X"DB",X"FE",X"15",X"FD",X"5C",X"FB",X"B4",X"F9",X"18",X"F8",X"8B",X"F6",X"09",X"F5",X"98",X"F3",
		X"2F",X"F2",X"D7",X"F0",X"88",X"EF",X"4B",X"EE",X"12",X"ED",X"99",X"EC",X"11",X"ED",X"1C",X"EE",
		X"8B",X"EF",X"3D",X"F1",X"FA",X"F2",X"D7",X"F4",X"D3",X"F6",X"C6",X"F8",X"B9",X"FA",X"A0",X"FC",
		X"80",X"FE",X"50",X"00",X"14",X"02",X"CC",X"03",X"77",X"05",X"11",X"07",X"9F",X"08",X"20",X"0A",
		X"96",X"0B",X"FD",X"0C",X"57",X"0E",X"A6",X"0F",X"E9",X"10",X"22",X"12",X"4C",X"13",X"72",X"14",
		X"59",X"15",X"3F",X"15",X"68",X"14",X"0F",X"13",X"68",X"11",X"8D",X"0F",X"98",X"0D",X"94",X"0B",
		X"8C",X"09",X"88",X"07",X"87",X"05",X"93",X"03",X"AA",X"01",X"CF",X"FF",X"01",X"FE",X"41",X"FC",
		X"90",X"FA",X"EB",X"F8",X"55",X"F7",X"CC",X"F5",X"50",X"F4",X"E0",X"F2",X"7F",X"F1",X"27",X"F0",
		X"DE",X"EE",X"9E",X"ED",X"6F",X"EC",X"41",X"EB",X"B3",X"EA",X"22",X"EB",X"26",X"EC",X"97",X"ED",
		X"45",X"EF",X"1D",X"F1",X"08",X"F3",X"02",X"F5",X"F7",X"F6",X"EC",X"F8",X"D4",X"FA",X"B7",X"FC",
		X"8A",X"FE",X"50",X"00",X"0A",X"02",X"B6",X"03",X"54",X"05",X"E6",X"06",X"68",X"08",X"DF",X"09",
		X"48",X"0B",X"A5",X"0C",X"F7",X"0D",X"3C",X"0F",X"76",X"10",X"A4",X"11",X"C8",X"12",X"E2",X"13",
		X"F0",X"14",X"F6",X"15",X"F1",X"16",X"E4",X"17",X"CE",X"18",X"AE",X"19",X"87",X"1A",X"56",X"1B",
		X"21",X"1C",X"E0",X"1C",X"99",X"1D",X"4A",X"1E",X"F7",X"1E",X"98",X"1F",X"37",X"20",X"CD",X"20",
		X"5F",X"21",X"E8",X"21",X"70",X"22",X"EE",X"22",X"68",X"23",X"DC",X"23",X"4D",X"24",X"B5",X"24",
		X"1D",X"25",X"7B",X"25",X"E0",X"25",X"CA",X"25",X"BA",X"24",X"13",X"23",X"02",X"21",X"B6",X"1E",
		X"43",X"1C",X"C0",X"19",X"35",X"17",X"B1",X"14",X"32",X"12",X"BF",X"0F",X"5B",X"0D",X"09",X"0B",
		X"C4",X"08",X"93",X"06",X"73",X"04",X"65",X"02",X"65",X"00",X"78",X"FE",X"9B",X"FC",X"CD",X"FA",
		X"10",X"F9",X"61",X"F7",X"BE",X"F5",X"2C",X"F4",X"A8",X"F2",X"32",X"F1",X"C5",X"EF",X"69",X"EE",
		X"17",X"ED",X"D1",X"EB",X"98",X"EA",X"67",X"E9",X"44",X"E8",X"2A",X"E7",X"1C",X"E6",X"16",X"E5",
		X"1A",X"E4",X"27",X"E3",X"3D",X"E2",X"5A",X"E1",X"84",X"E0",X"B3",X"DF",X"E9",X"DE",X"28",X"DE",
		X"6E",X"DD",X"BD",X"DC",X"13",X"DC",X"6D",X"DB",X"D0",X"DA",X"35",X"DA",X"A7",X"D9",X"19",X"D9",
		X"98",X"D8",X"10",X"D8",X"E9",X"D7",X"B7",X"D8",X"23",X"DA",X"FF",X"DB",X"1C",X"DE",X"61",X"E0",
		X"BC",X"E2",X"1D",X"E5",X"7C",X"E7",X"D7",X"E9",X"25",X"EC",X"67",X"EE",X"98",X"F0",X"BC",X"F2",
		X"CF",X"F4",X"D3",X"F6",X"C5",X"F8",X"A8",X"FA",X"7B",X"FC",X"3D",X"FE",X"F1",X"FF",X"98",X"01",
		X"2E",X"03",X"B9",X"04",X"36",X"06",X"A6",X"07",X"06",X"09",X"5A",X"0A",X"EC",X"0A",X"9A",X"0A",
		X"C4",X"09",X"8B",X"08",X"1B",X"07",X"85",X"05",X"DC",X"03",X"2A",X"02",X"79",X"00",X"C9",X"FE",
		X"22",X"FD",X"82",X"FB",X"EF",X"F9",X"64",X"F8",X"E6",X"F6",X"74",X"F5",X"0F",X"F4",X"B5",X"F2",
		X"66",X"F1",X"22",X"F0",X"EA",X"EE",X"BC",X"ED",X"9A",X"EC",X"81",X"EB",X"73",X"EA",X"6D",X"E9",
		X"73",X"E8",X"80",X"E7",X"97",X"E6",X"B4",X"E5",X"DE",X"E4",X"0D",X"E4",X"44",X"E3",X"82",X"E2",
		X"C9",X"E1",X"15",X"E1",X"6C",X"E0",X"C6",X"DF",X"26",X"DF",X"8E",X"DE",X"FB",X"DD",X"6E",X"DD",
		X"EA",X"DC",X"67",X"DC",X"EC",X"DB",X"75",X"DB",X"05",X"DB",X"96",X"DA",X"32",X"DA",X"CD",X"D9",
		X"6F",X"D9",X"14",X"D9",X"C0",X"D8",X"68",X"D8",X"43",X"D8",X"00",X"D9",X"6E",X"DA",X"4F",X"DC",
		X"76",X"DE",X"C9",X"E0",X"31",X"E3",X"A2",X"E5",X"13",X"E8",X"7E",X"EA",X"DC",X"EC",X"2F",X"EF",
		X"70",X"F1",X"A5",X"F3",X"C7",X"F5",X"D9",X"F7",X"DB",X"F9",X"CB",X"FB",X"AB",X"FD",X"7D",X"FF",
		X"3D",X"01",X"F1",X"02",X"93",X"04",X"28",X"06",X"AF",X"07",X"2B",X"09",X"95",X"0A",X"FC",X"0B",
		X"D3",X"0C",X"BD",X"0C",X"13",X"0C",X"05",X"0B",X"B7",X"09",X"3F",X"08",X"B3",X"06",X"19",X"05",
		X"7F",X"03",X"E5",X"01",X"53",X"00",X"C6",X"FE",X"47",X"FD",X"CF",X"FB",X"61",X"FA",X"00",X"F9",
		X"AB",X"F7",X"5F",X"F6",X"1F",X"F5",X"E9",X"F3",X"BE",X"F2",X"9E",X"F1",X"87",X"F0",X"79",X"EF",
		X"77",X"EE",X"7E",X"ED",X"8B",X"EC",X"A2",X"EB",X"C3",X"EA",X"EA",X"E9",X"1B",X"E9",X"51",X"E8",
		X"91",X"E7",X"D7",X"E6",X"25",X"E6",X"79",X"E5",X"D4",X"E4",X"35",X"E4",X"9D",X"E3",X"0A",X"E3",
		X"7E",X"E2",X"F5",X"E1",X"73",X"E1",X"F6",X"E0",X"7E",X"E0",X"0D",X"E0",X"9E",X"DF",X"35",X"DF",
		X"D0",X"DE",X"70",X"DE",X"15",X"DE",X"BD",X"DD",X"6A",X"DD",X"19",X"DD",X"CD",X"DC",X"84",X"DC",
		X"3F",X"DC",X"00",X"DC",X"BF",X"DB",X"84",X"DB",X"4D",X"DB",X"17",X"DB",X"E5",X"DA",X"B7",X"DA",
		X"88",X"DA",X"5F",X"DA",X"37",X"DA",X"12",X"DA",X"F0",X"D9",X"D0",X"D9",X"B3",X"D9",X"96",X"D9",
		X"7D",X"D9",X"64",X"D9",X"4F",X"D9",X"3C",X"D9",X"2A",X"D9",X"1A",X"D9",X"0C",X"D9",X"FE",X"D8",
		X"F3",X"D8",X"EB",X"D8",X"E3",X"D8",X"DC",X"D8",X"D7",X"D8",X"D3",X"D8",X"D1",X"D8",X"D0",X"D8",
		X"D0",X"D8",X"D2",X"D8",X"D4",X"D8",X"D8",X"D8",X"DD",X"D8",X"E2",X"D8",X"E9",X"D8",X"F1",X"D8",
		X"F9",X"D8",X"04",X"D9",X"0E",X"D9",X"19",X"D9",X"25",X"D9",X"33",X"D9",X"42",X"D9",X"4F",X"D9",
		X"5E",X"D9",X"6E",X"D9",X"7F",X"D9",X"91",X"D9",X"A1",X"D9",X"B4",X"D9",X"C7",X"D9",X"DD",X"D9",
		X"EF",X"D9",X"05",X"DA",X"19",X"DA",X"2E",X"DA",X"45",X"DA",X"5C",X"DA",X"73",X"DA",X"8A",X"DA",
		X"A2",X"DA",X"BC",X"DA",X"D4",X"DA",X"ED",X"DA",X"05",X"DB",X"20",X"DB",X"39",X"DB",X"53",X"DB",
		X"6E",X"DB",X"89",X"DB",X"A2",X"DB",X"BF",X"DB",X"DA",X"DB",X"F6",X"DB",X"11",X"DC",X"30",X"DC",
		X"4A",X"DC",X"67",X"DC",X"84",X"DC",X"A0",X"DC",X"BE",X"DC",X"DB",X"DC",X"F8",X"DC",X"16",X"DD",
		X"33",X"DD",X"51",X"DD",X"6F",X"DD",X"8D",X"DD",X"AA",X"DD",X"CA",X"DD",X"E7",X"DD",X"05",X"DE",
		X"23",X"DE",X"44",X"DE",X"61",X"DE",X"7F",X"DE",X"9D",X"DE",X"BE",X"DE",X"DB",X"DE",X"FB",X"DE",
		X"1A",X"DF",X"39",X"DF",X"57",X"DF",X"76",X"DF",X"90",X"DF",X"DE",X"DF",X"02",X"E1",X"C1",X"E2",
		X"E8",X"E4",X"47",X"E7",X"D3",X"E9",X"42",X"EC",X"CE",X"EE",X"72",X"F1",X"03",X"F4",X"8D",X"F6",
		X"03",X"F9",X"6B",X"FB",X"BF",X"FD",X"03",X"00",X"32",X"02",X"53",X"04",X"60",X"06",X"5D",X"08",
		X"47",X"0A",X"21",X"0C",X"EC",X"0D",X"A7",X"0F",X"52",X"11",X"EE",X"12",X"7E",X"14",X"FC",X"15",
		X"73",X"17",X"55",X"18",X"57",X"18",X"D3",X"17",X"ED",X"16",X"CE",X"15",X"86",X"14",X"2A",X"13",
		X"C3",X"11",X"5A",X"10",X"ED",X"0E",X"89",X"0D",X"2B",X"0C",X"D4",X"0A",X"86",X"09",X"41",X"08",
		X"05",X"07",X"D4",X"05",X"AC",X"04",X"8E",X"03",X"7A",X"02",X"6D",X"01",X"6A",X"00",X"70",X"FF",
		X"80",X"FE",X"95",X"FD",X"B3",X"FC",X"D7",X"FB",X"23",X"FB",X"3C",X"FB",X"08",X"FC",X"41",X"FD",
		X"C3",X"FE",X"6D",X"00",X"35",X"02",X"07",X"04",X"DB",X"05",X"AD",X"07",X"78",X"09",X"3C",X"0B",
		X"F1",X"0C",X"9B",X"0E",X"39",X"10",X"CB",X"11",X"4D",X"13",X"C5",X"14",X"2F",X"16",X"8D",X"17",
		X"DC",X"18",X"23",X"1A",X"5C",X"1B",X"8B",X"1C",X"AF",X"1D",X"C9",X"1E",X"D4",X"1F",X"DE",X"20",
		X"72",X"21",X"2B",X"21",X"58",X"20",X"21",X"1F",X"B6",X"1D",X"20",X"1C",X"7A",X"1A",X"C8",X"18",
		X"17",X"17",X"67",X"15",X"BD",X"13",X"1C",X"12",X"85",X"10",X"F7",X"0E",X"77",X"0D",X"01",X"0C",
		X"96",X"0A",X"36",X"09",X"E3",X"07",X"99",X"06",X"5D",X"05",X"2A",X"04",X"00",X"03",X"E0",X"01",
		X"CA",X"00",X"BE",X"FF",X"BB",X"FE",X"BF",X"FD",X"CE",X"FC",X"E4",X"FB",X"02",X"FB",X"28",X"FA",
		X"56",X"F9",X"8B",X"F8",X"C8",X"F7",X"0A",X"F7",X"53",X"F6",X"A4",X"F5",X"FA",X"F4",X"58",X"F4",
		X"B9",X"F3",X"21",X"F3",X"90",X"F2",X"04",X"F2",X"7C",X"F1",X"F9",X"F0",X"7B",X"F0",X"03",X"F0",
		X"8D",X"EF",X"1E",X"EF",X"B3",X"EE",X"4C",X"EE",X"E9",X"ED",X"89",X"ED",X"2E",X"ED",X"D6",X"EC",
		X"81",X"EC",X"32",X"EC",X"E4",X"EB",X"9A",X"EB",X"54",X"EB",X"11",X"EB",X"CF",X"EA",X"92",X"EA",
		X"56",X"EA",X"1F",X"EA",X"E9",X"E9",X"B6",X"E9",X"86",X"E9",X"57",X"E9",X"2B",X"E9",X"01",X"E9",
		X"DA",X"E8",X"B4",X"E8",X"8F",X"E8",X"71",X"E8",X"4F",X"E8",X"33",X"E8",X"17",X"E8",X"FE",X"E7",
		X"E4",X"E7",X"CE",X"E7",X"BD",X"E7",X"50",X"E8",X"9F",X"E9",X"5A",X"EB",X"63",X"ED",X"91",X"EF",
		X"DD",X"F1",X"2C",X"F4",X"81",X"F6",X"CC",X"F8",X"0E",X"FB",X"45",X"FD",X"6B",X"FF",X"80",X"01",
		X"8A",X"03",X"82",X"05",X"68",X"07",X"40",X"09",X"08",X"0B",X"C1",X"0C",X"6B",X"0E",X"05",X"10",
		X"94",X"11",X"13",X"13",X"85",X"14",X"EA",X"15",X"42",X"17",X"8E",X"18",X"CF",X"19",X"03",X"1B",
		X"2D",X"1C",X"4A",X"1D",X"5F",X"1E",X"69",X"1F",X"69",X"20",X"60",X"21",X"4E",X"22",X"31",X"23",
		X"0D",X"24",X"DF",X"24",X"AB",X"25",X"6E",X"26",X"29",X"27",X"DC",X"27",X"88",X"28",X"2F",X"29",
		X"CE",X"29",X"65",X"2A",X"F7",X"2A",X"82",X"2B",X"07",X"2C",X"86",X"2C",X"01",X"2D",X"75",X"2D",
		X"E4",X"2D",X"4F",X"2E",X"B4",X"2E",X"14",X"2F",X"6F",X"2F",X"C7",X"2F",X"19",X"30",X"68",X"30",
		X"B1",X"30",X"F7",X"30",X"3A",X"31",X"79",X"31",X"B4",X"31",X"EC",X"31",X"1F",X"32",X"51",X"32",
		X"7E",X"32",X"AA",X"32",X"D0",X"32",X"F5",X"32",X"18",X"33",X"37",X"33",X"55",X"33",X"6D",X"33",
		X"85",X"33",X"9B",X"33",X"AD",X"33",X"BE",X"33",X"CD",X"33",X"D9",X"33",X"E4",X"33",X"ED",X"33",
		X"F3",X"33",X"F9",X"33",X"FA",X"33",X"FC",X"33",X"FC",X"33",X"FC",X"33",X"F6",X"33",X"F3",X"33",
		X"EA",X"33",X"E4",X"33",X"DA",X"33",X"CF",X"33",X"C3",X"33",X"B6",X"33",X"A9",X"33",X"99",X"33",
		X"89",X"33",X"78",X"33",X"64",X"33",X"51",X"33",X"3D",X"33",X"28",X"33",X"10",X"33",X"FC",X"32",
		X"CE",X"32",X"E9",X"31",X"62",X"30",X"7D",X"2E",X"55",X"2C",X"0B",X"2A",X"AF",X"27",X"4D",X"25",
		X"EA",X"22",X"90",X"20",X"43",X"1E",X"FE",X"1B",X"CA",X"19",X"A7",X"17",X"92",X"15",X"8D",X"13",
		X"99",X"11",X"B3",X"0F",X"DF",X"0D",X"18",X"0C",X"60",X"0A",X"B6",X"08",X"1C",X"07",X"8D",X"05",
		X"0B",X"04",X"98",X"02",X"32",X"01",X"D6",X"FF",X"86",X"FE",X"41",X"FD",X"07",X"FC",X"D9",X"FA",
		X"B4",X"F9",X"9B",X"F8",X"8A",X"F7",X"83",X"F6",X"83",X"F5",X"8E",X"F4",X"A2",X"F3",X"BD",X"F2",
		X"E0",X"F1",X"0D",X"F1",X"3F",X"F0",X"7A",X"EF",X"BD",X"EE",X"05",X"EE",X"55",X"ED",X"A9",X"EC",
		X"05",X"EC",X"68",X"EB",X"D0",X"EA",X"3F",X"EA",X"B2",X"E9",X"2B",X"E9",X"A9",X"E8",X"2E",X"E8",
		X"B5",X"E7",X"41",X"E7",X"D4",X"E6",X"69",X"E6",X"04",X"E6",X"A3",X"E5",X"46",X"E5",X"EC",X"E4",
		X"97",X"E4",X"45",X"E4",X"F7",X"E3",X"AC",X"E3",X"65",X"E3",X"22",X"E3",X"E0",X"E2",X"A3",X"E2",
		X"68",X"E2",X"2F",X"E2",X"FB",X"E1",X"C9",X"E1",X"9A",X"E1",X"6C",X"E1",X"41",X"E1",X"18",X"E1",
		X"F3",X"E0",X"D0",X"E0",X"AD",X"E0",X"90",X"E0",X"71",X"E0",X"56",X"E0",X"3D",X"E0",X"24",X"E0",
		X"0F",X"E0",X"FB",X"DF",X"E8",X"DF",X"D6",X"DF",X"C8",X"DF",X"BB",X"DF",X"AE",X"DF",X"A4",X"DF",
		X"9A",X"DF",X"92",X"DF",X"8B",X"DF",X"86",X"DF",X"81",X"DF",X"7E",X"DF",X"7C",X"DF",X"79",X"DF",
		X"7B",X"DF",X"7D",X"DF",X"7E",X"DF",X"81",X"DF",X"86",X"DF",X"8A",X"DF",X"90",X"DF",X"97",X"DF",
		X"9E",X"DF",X"A6",X"DF",X"B0",X"DF",X"BA",X"DF",X"C4",X"DF",X"CF",X"DF",X"DB",X"DF",X"E6",X"DF",
		X"F5",X"DF",X"01",X"E0",X"10",X"E0",X"1D",X"E0",X"2C",X"E0",X"3D",X"E0",X"4D",X"E0",X"5D",X"E0",
		X"6E",X"E0",X"7F",X"E0",X"92",X"E0",X"A3",X"E0",X"B8",X"E0",X"CB",X"E0",X"DE",X"E0",X"F2",X"E0",
		X"06",X"E1",X"16",X"E1",X"57",X"E1",X"53",X"E2",X"D6",X"E3",X"B0",X"E5",X"C0",X"E7",X"EE",X"E9",
		X"29",X"EC",X"69",X"EE",X"A7",X"F0",X"DB",X"F2",X"07",X"F5",X"22",X"F7",X"32",X"F9",X"30",X"FB",
		X"22",X"FD",X"01",X"FF",X"D3",X"00",X"95",X"02",X"49",X"04",X"EE",X"05",X"86",X"07",X"0D",X"09",
		X"8C",X"0A",X"F7",X"0B",X"5B",X"0D",X"AF",X"0E",X"FB",X"0F",X"37",X"11",X"6C",X"12",X"93",X"13",
		X"B4",X"14",X"C3",X"15",X"D1",X"16",X"C8",X"17",X"EE",X"18",X"F8",X"19",X"D7",X"1A",X"BC",X"1B",
		X"8D",X"1C",X"5E",X"1D",X"22",X"1E",X"E2",X"1E",X"9A",X"1F",X"48",X"20",X"F1",X"20",X"95",X"21",
		X"30",X"22",X"C7",X"22",X"56",X"23",X"E0",X"23",X"62",X"24",X"E1",X"24",X"5A",X"25",X"CD",X"25",
		X"3F",X"26",X"8D",X"26",X"27",X"26",X"28",X"25",X"CD",X"23",X"35",X"22",X"7B",X"20",X"AB",X"1E",
		X"D3",X"1C",X"FA",X"1A",X"23",X"19",X"55",X"17",X"8F",X"15",X"D5",X"13",X"28",X"12",X"85",X"10",
		X"EE",X"0E",X"67",X"0D",X"E8",X"0B",X"79",X"0A",X"14",X"09",X"BA",X"07",X"6B",X"06",X"29",X"05",
		X"EE",X"03",X"C3",X"02",X"9C",X"01",X"85",X"00",X"6F",X"FF",X"C5",X"FE",X"DB",X"FE",X"68",X"FF",
		X"4B",X"00",X"5E",X"01",X"94",X"02",X"DA",X"03",X"2B",X"05",X"7C",X"06",X"CB",X"07",X"15",X"09",
		X"5A",X"0A",X"95",X"0B",X"C8",X"0C",X"F1",X"0D",X"12",X"0F",X"29",X"10",X"36",X"11",X"38",X"12",
		X"35",X"13",X"27",X"14",X"10",X"15",X"F3",X"15",X"CC",X"16",X"9B",X"17",X"65",X"18",X"28",X"19",
		X"D3",X"19",X"D6",X"19",X"39",X"19",X"3A",X"18",X"F7",X"16",X"90",X"15",X"11",X"14",X"85",X"12",
		X"F5",X"10",X"68",X"0F",X"DE",X"0D",X"5D",X"0C",X"E4",X"0A",X"76",X"09",X"11",X"08",X"B5",X"06",
		X"64",X"05",X"20",X"04",X"E6",X"02",X"B5",X"01",X"8E",X"00",X"73",X"FF",X"60",X"FE",X"56",X"FD",
		X"53",X"FC",X"5D",X"FB",X"6D",X"FA",X"85",X"F9",X"A6",X"F8",X"CF",X"F7",X"FD",X"F6",X"35",X"F6",
		X"74",X"F5",X"B9",X"F4",X"04",X"F4",X"56",X"F3",X"AE",X"F2",X"0E",X"F2",X"72",X"F1",X"DC",X"F0",
		X"4C",X"F0",X"C1",X"EF",X"3B",X"EF",X"BC",X"EE",X"3E",X"EE",X"C7",X"ED",X"55",X"ED",X"E8",X"EC",
		X"7D",X"EC",X"18",X"EC",X"B5",X"EB",X"59",X"EB",X"FF",X"EA",X"AA",X"EA",X"56",X"EA",X"08",X"EA",
		X"BC",X"E9",X"73",X"E9",X"2F",X"E9",X"EE",X"E8",X"AE",X"E8",X"72",X"E8",X"37",X"E8",X"01",X"E8",
		X"CC",X"E7",X"9C",X"E7",X"6B",X"E7",X"3F",X"E7",X"14",X"E7",X"ED",X"E6",X"C6",X"E6",X"A3",X"E6",
		X"81",X"E6",X"61",X"E6",X"42",X"E6",X"27",X"E6",X"0C",X"E6",X"F3",X"E5",X"DB",X"E5",X"C7",X"E5",
		X"B2",X"E5",X"A2",X"E5",X"8B",X"E5",X"AE",X"E5",X"83",X"E6",X"D3",X"E7",X"74",X"E9",X"48",X"EB",
		X"37",X"ED",X"34",X"EF",X"35",X"F1",X"36",X"F3",X"2C",X"F5",X"1B",X"F7",X"FE",X"F8",X"D4",X"FA",
		X"9B",X"FC",X"57",X"FE",X"04",X"00",X"A4",X"01",X"35",X"03",X"B9",X"04",X"32",X"06",X"9E",X"07",
		X"FA",X"08",X"4E",X"0A",X"95",X"0B",X"D1",X"0C",X"01",X"0E",X"28",X"0F",X"45",X"10",X"56",X"11",
		X"5D",X"12",X"5D",X"13",X"51",X"14",X"3D",X"15",X"22",X"16",X"FD",X"16",X"D1",X"17",X"9B",X"18",
		X"60",X"19",X"1D",X"1A",X"D1",X"1A",X"80",X"1B",X"28",X"1C",X"CA",X"1C",X"63",X"1D",X"F9",X"1D",
		X"87",X"1E",X"11",X"1F",X"92",X"1F",X"14",X"20",X"8B",X"20",X"FE",X"20",X"6D",X"21",X"D8",X"21",
		X"3C",X"22",X"A1",X"22",X"DF",X"22",X"6E",X"22",X"77",X"21",X"2B",X"20",X"A9",X"1E",X"06",X"1D",
		X"52",X"1B",X"98",X"19",X"DB",X"17",X"23",X"16",X"72",X"14",X"CB",X"12",X"2D",X"11",X"9B",X"0F",
		X"14",X"0E",X"99",X"0C",X"2B",X"0B",X"C5",X"09",X"6D",X"08",X"1F",X"07",X"DC",X"05",X"A4",X"04",
		X"77",X"03",X"53",X"02",X"39",X"01",X"28",X"00",X"22",X"FF",X"23",X"FE",X"2D",X"FD",X"40",X"FC",
		X"5A",X"FB",X"7C",X"FA",X"A7",X"F9",X"D8",X"F8",X"12",X"F8",X"52",X"F7",X"97",X"F6",X"E4",X"F5",
		X"38",X"F5",X"92",X"F4",X"F1",X"F3",X"57",X"F3",X"C2",X"F2",X"33",X"F2",X"A8",X"F1",X"23",X"F1",
		X"A2",X"F0",X"28",X"F0",X"B2",X"EF",X"40",X"EF",X"D1",X"EE",X"67",X"EE",X"03",X"EE",X"A1",X"ED",
		X"44",X"ED",X"EB",X"EC",X"95",X"EC",X"42",X"EC",X"F1",X"EB",X"A7",X"EB",X"5F",X"EB",X"19",X"EB",
		X"D7",X"EA",X"96",X"EA",X"5B",X"EA",X"21",X"EA",X"EA",X"E9",X"B4",X"E9",X"82",X"E9",X"52",X"E9",
		X"23",X"E9",X"FA",X"E8",X"D2",X"E8",X"AA",X"E8",X"85",X"E8",X"63",X"E8",X"42",X"E8",X"24",X"E8",
		X"05",X"E8",X"EB",X"E7",X"D1",X"E7",X"B9",X"E7",X"A2",X"E7",X"8D",X"E7",X"7A",X"E7",X"69",X"E7",
		X"58",X"E7",X"48",X"E7",X"3B",X"E7",X"2E",X"E7",X"23",X"E7",X"18",X"E7",X"10",X"E7",X"07",X"E7",
		X"01",X"E7",X"FC",X"E6",X"F8",X"E6",X"F4",X"E6",X"F1",X"E6",X"EE",X"E6",X"EE",X"E6",X"ED",X"E6",
		X"EF",X"E6",X"F0",X"E6",X"F2",X"E6",X"F6",X"E6",X"F9",X"E6",X"FE",X"E6",X"02",X"E7",X"0A",X"E7",
		X"0F",X"E7",X"16",X"E7",X"1E",X"E7",X"26",X"E7",X"2E",X"E7",X"39",X"E7",X"42",X"E7",X"4C",X"E7",
		X"58",X"E7",X"64",X"E7",X"6E",X"E7",X"7B",X"E7",X"86",X"E7",X"94",X"E7",X"A0",X"E7",X"AF",X"E7",
		X"BE",X"E7",X"CB",X"E7",X"DB",X"E7",X"E9",X"E7",X"F9",X"E7",X"09",X"E8",X"17",X"E8",X"28",X"E8",
		X"3A",X"E8",X"48",X"E8",X"5A",X"E8",X"6D",X"E8",X"02",X"E9",X"2A",X"EA",X"AA",X"EB",X"65",X"ED",
		X"41",X"EF",X"2F",X"F1",X"23",X"F3",X"17",X"F5",X"05",X"F7",X"EC",X"F8",X"C7",X"FA",X"96",X"FC",
		X"58",X"FE",X"0C",X"00",X"B1",X"01",X"4C",X"03",X"D8",X"04",X"58",X"06",X"CA",X"07",X"32",X"09",
		X"8C",X"0A",X"D9",X"0B",X"1C",X"0D",X"52",X"0E",X"80",X"0F",X"A2",X"10",X"B9",X"11",X"C7",X"12",
		X"CA",X"13",X"C5",X"14",X"B7",X"15",X"A1",X"16",X"81",X"17",X"5B",X"18",X"2A",X"19",X"F2",X"19",
		X"B4",X"1A",X"6D",X"1B",X"1F",X"1C",X"CB",X"1C",X"70",X"1D",X"0E",X"1E",X"A9",X"1E",X"3A",X"1F",
		X"C6",X"1F",X"4D",X"20",X"CF",X"20",X"4A",X"21",X"C2",X"21",X"33",X"22",X"9E",X"22",X"07",X"23",
		X"6B",X"23",X"C9",X"23",X"26",X"24",X"7B",X"24",X"CE",X"24",X"1D",X"25",X"68",X"25",X"B0",X"25",
		X"F2",X"25",X"33",X"26",X"70",X"26",X"AB",X"26",X"E1",X"26",X"15",X"27",X"45",X"27",X"74",X"27",
		X"9E",X"27",X"C7",X"27",X"EC",X"27",X"11",X"28",X"30",X"28",X"51",X"28",X"6A",X"28",X"84",X"28",
		X"9D",X"28",X"B3",X"28",X"C7",X"28",X"DA",X"28",X"E8",X"28",X"FC",X"28",X"EC",X"28",X"47",X"28",
		X"22",X"27",X"B6",X"25",X"12",X"24",X"5A",X"22",X"86",X"20",X"ED",X"1E",X"3A",X"1D",X"60",X"1B",
		X"A0",X"19",X"DE",X"17",X"2F",X"16",X"87",X"14",X"EF",X"12",X"5F",X"11",X"DE",X"0F",X"67",X"0E",
		X"FE",X"0C",X"9F",X"0B",X"4C",X"0A",X"04",X"09",X"C8",X"07",X"94",X"06",X"6C",X"05",X"4D",X"04",
		X"38",X"03",X"2B",X"02",X"28",X"01",X"2E",X"00",X"3B",X"FF",X"53",X"FE",X"70",X"FD",X"98",X"FC",
		X"C4",X"FB",X"F9",X"FA",X"35",X"FA",X"77",X"F9",X"C0",X"F8",X"10",X"F8",X"65",X"F7",X"C2",X"F6",
		X"23",X"F6",X"8A",X"F5",X"F7",X"F4",X"6A",X"F4",X"E1",X"F3",X"5D",X"F3",X"DD",X"F2",X"65",X"F2",
		X"EE",X"F1",X"7D",X"F1",X"10",X"F1",X"A9",X"F0",X"44",X"F0",X"E2",X"EF",X"85",X"EF",X"2D",X"EF",
		X"D7",X"EE",X"85",X"EE",X"35",X"EE",X"EA",X"ED",X"A1",X"ED",X"5C",X"ED",X"1B",X"ED",X"DA",X"EC",
		X"9D",X"EC",X"64",X"EC",X"2B",X"EC",X"F6",X"EB",X"C3",X"EB",X"94",X"EB",X"65",X"EB",X"3A",X"EB",
		X"11",X"EB",X"E9",X"EA",X"C2",X"EA",X"A1",X"EA",X"7E",X"EA",X"60",X"EA",X"40",X"EA",X"27",X"EA",
		X"06",X"EA",X"2C",X"EA",X"F0",X"EA",X"19",X"EC",X"86",X"ED",X"19",X"EF",X"C2",X"F0",X"79",X"F2",
		X"32",X"F4",X"E9",X"F5",X"99",X"F7",X"3E",X"F9",X"DD",X"FA",X"6E",X"FC",X"F7",X"FD",X"71",X"FF",
		X"DF",X"00",X"42",X"02",X"9A",X"03",X"E6",X"04",X"28",X"06",X"5F",X"07",X"8B",X"08",X"AC",X"09",
		X"C4",X"0A",X"D1",X"0B",X"D7",X"0C",X"D1",X"0D",X"BF",X"0E",X"25",X"0F",X"FB",X"0E",X"7A",X"0E",
		X"BD",X"0D",X"DB",X"0C",X"E0",X"0B",X"D7",X"0A",X"CC",X"09",X"BD",X"08",X"B0",X"07",X"A9",X"06",
		X"A5",X"05",X"A9",X"04",X"B2",X"03",X"C5",X"02",X"DC",X"01",X"FD",X"00",X"24",X"00",X"52",X"FF",
		X"87",X"FE",X"C2",X"FD",X"06",X"FD",X"4D",X"FC",X"9E",X"FB",X"F2",X"FA",X"4F",X"FA",X"AC",X"F9",
		X"40",X"F9",X"71",X"F9",X"0F",X"FA",X"F7",X"FA",X"0A",X"FC",X"3C",X"FD",X"7D",X"FE",X"C2",X"FF",
		X"0A",X"01",X"4F",X"02",X"90",X"03",X"CA",X"04",X"FB",X"05",X"25",X"07",X"45",X"08",X"5B",X"09",
		X"6A",X"0A",X"6F",X"0B",X"6B",X"0C",X"5F",X"0D",X"4A",X"0E",X"2E",X"0F",X"08",X"10",X"DA",X"10",
		X"A7",X"11",X"6A",X"12",X"26",X"13",X"DC",X"13",X"8D",X"14",X"34",X"15",X"D8",X"15",X"73",X"16",
		X"09",X"17",X"9B",X"17",X"25",X"18",X"A9",X"18",X"2B",X"19",X"A4",X"19",X"1B",X"1A",X"8D",X"1A",
		X"FB",X"1A",X"63",X"1B",X"C7",X"1B",X"26",X"1C",X"82",X"1C",X"D8",X"1C",X"2D",X"1D",X"7C",X"1D",
		X"CA",X"1D",X"11",X"1E",X"58",X"1E",X"99",X"1E",X"D9",X"1E",X"12",X"1F",X"50",X"1F",X"67",X"1F",
		X"EA",X"1E",X"00",X"1E",X"CC",X"1C",X"69",X"1B",X"EF",X"19",X"63",X"18",X"D5",X"16",X"45",X"15",
		X"BB",X"13",X"36",X"12",X"BA",X"10",X"47",X"0F",X"DE",X"0D",X"82",X"0C",X"2D",X"0B",X"E5",X"09",
		X"A5",X"08",X"71",X"07",X"47",X"06",X"27",X"05",X"0E",X"04",X"00",X"03",X"F9",X"01",X"FF",X"00",
		X"0A",X"00",X"22",X"FF",X"3A",X"FE",X"B5",X"FD",X"C4",X"FD",X"31",X"FE",X"E0",X"FE",X"B3",X"FF",
		X"A1",X"00",X"99",X"01",X"9E",X"02",X"A0",X"03",X"A4",X"04",X"A2",X"05",X"9B",X"06",X"8D",X"07",
		X"79",X"08",X"5F",X"09",X"3D",X"0A",X"14",X"0B",X"E2",X"0B",X"AB",X"0C",X"6C",X"0D",X"26",X"0E",
		X"DA",X"0E",X"88",X"0F",X"2E",X"10",X"CF",X"10",X"6B",X"11",X"00",X"12",X"8F",X"12",X"1A",X"13",
		X"9E",X"13",X"1D",X"14",X"97",X"14",X"0E",X"15",X"7E",X"15",X"EC",X"15",X"55",X"16",X"B9",X"16",
		X"19",X"17",X"75",X"17",X"CE",X"17",X"21",X"18",X"73",X"18",X"C0",X"18",X"09",X"19",X"52",X"19",
		X"94",X"19",X"D5",X"19",X"12",X"1A",X"4D",X"1A",X"83",X"1A",X"B9",X"1A",X"EB",X"1A",X"1C",X"1B",
		X"45",X"1B",X"76",X"1B",X"5C",X"1B",X"B1",X"1A",X"AB",X"19",X"67",X"18",X"00",X"17",X"82",X"15",
		X"FD",X"13",X"71",X"12",X"E8",X"10",X"65",X"0F",X"EB",X"0D",X"76",X"0C",X"0E",X"0B",X"AF",X"09",
		X"5A",X"08",X"10",X"07",X"D0",X"05",X"99",X"04",X"6E",X"03",X"4C",X"02",X"33",X"01",X"24",X"00",
		X"20",X"FF",X"22",X"FE",X"2F",X"FD",X"43",X"FC",X"5F",X"FB",X"81",X"FA",X"AD",X"F9",X"DD",X"F8",
		X"19",X"F8",X"5A",X"F7",X"A0",X"F6",X"EF",X"F5",X"43",X"F5",X"9E",X"F4",X"FD",X"F3",X"63",X"F3",
		X"CE",X"F2",X"3F",X"F2",X"B7",X"F1",X"31",X"F1",X"B2",X"F0",X"37",X"F0",X"C2",X"EF",X"4E",X"EF",
		X"DF",X"EE",X"79",X"EE",X"12",X"EE",X"B2",X"ED",X"54",X"ED",X"FA",X"EC",X"A4",X"EC",X"53",X"EC",
		X"08",X"EC",X"2B",X"EC",X"D5",X"EC",X"C7",X"ED",X"EF",X"EE",X"35",X"F0",X"8E",X"F1",X"ED",X"F2",
		X"51",X"F4",X"B1",X"F5",X"0B",X"F7",X"5F",X"F8",X"AA",X"F9",X"EE",X"FA",X"27",X"FC",X"57",X"FD",
		X"7E",X"FE",X"9A",X"FF",X"AE",X"00",X"BA",X"01",X"BB",X"02",X"B3",X"03",X"A4",X"04",X"8C",X"05",
		X"6D",X"06",X"47",X"07",X"16",X"08",X"E5",X"08",X"82",X"09",X"90",X"09",X"35",X"09",X"96",X"08",
		X"CA",X"07",X"E3",X"06",X"EC",X"05",X"ED",X"04",X"EB",X"03",X"EA",X"02",X"EC",X"01",X"F2",X"00",
		X"FF",X"FF",X"11",X"FF",X"2D",X"FE",X"4D",X"FD",X"75",X"FC",X"A2",X"FB",X"DA",X"FA",X"15",X"FA",
		X"59",X"F9",X"A0",X"F8",X"F1",X"F7",X"47",X"F7",X"A4",X"F6",X"03",X"F6",X"6D",X"F5",X"D9",X"F4",
		X"A7",X"F4",X"FE",X"F4",X"A4",X"F5",X"83",X"F6",X"82",X"F7",X"96",X"F8",X"B5",X"F9",X"D9",X"FA",
		X"FD",X"FB",X"1D",X"FD",X"37",X"FE",X"4E",X"FF",X"5A",X"00",X"5D",X"01",X"5C",X"02",X"54",X"03",
		X"41",X"04",X"28",X"05",X"07",X"06",X"DE",X"06",X"AD",X"07",X"76",X"08",X"37",X"09",X"F2",X"09",
		X"A6",X"0A",X"53",X"0B",X"FD",X"0B",X"88",X"0C",X"89",X"0C",X"1E",X"0C",X"6E",X"0B",X"93",X"0A",
		X"9A",X"09",X"92",X"08",X"81",X"07",X"70",X"06",X"5D",X"05",X"4F",X"04",X"46",X"03",X"44",X"02",
		X"48",X"01",X"53",X"00",X"66",X"FF",X"7F",X"FE",X"A2",X"FD",X"CB",X"FC",X"FA",X"FB",X"30",X"FB",
		X"6F",X"FA",X"B2",X"F9",X"FD",X"F8",X"4F",X"F8",X"A6",X"F7",X"04",X"F7",X"66",X"F6",X"D0",X"F5",
		X"3D",X"F5",X"B0",X"F4",X"29",X"F4",X"A6",X"F3",X"26",X"F3",X"B1",X"F2",X"21",X"F2",X"A1",X"F1",
		X"39",X"F1",X"CD",X"F0",X"6B",X"F0",X"09",X"F0",X"AD",X"EF",X"51",X"EF",X"FC",X"EE",X"A9",X"EE",
		X"5A",X"EE",X"0D",X"EE",X"C5",X"ED",X"7E",X"ED",X"3C",X"ED",X"FC",X"EC",X"BF",X"EC",X"83",X"EC",
		X"4C",X"EC",X"16",X"EC",X"E4",X"EB",X"B2",X"EB",X"85",X"EB",X"59",X"EB",X"2E",X"EB",X"06",X"EB",
		X"E0",X"EA",X"BC",X"EA",X"9B",X"EA",X"7A",X"EA",X"5C",X"EA",X"40",X"EA",X"25",X"EA",X"0A",X"EA",
		X"F3",X"E9",X"DB",X"E9",X"C8",X"E9",X"B3",X"E9",X"A2",X"E9",X"91",X"E9",X"83",X"E9",X"75",X"E9",
		X"67",X"E9",X"5B",X"E9",X"52",X"E9",X"47",X"E9",X"40",X"E9",X"34",X"E9",X"65",X"E9",X"1C",X"EA",
		X"27",X"EB",X"6A",X"EC",X"CC",X"ED",X"41",X"EF",X"C1",X"F0",X"42",X"F2",X"C1",X"F3",X"3A",X"F5",
		X"AB",X"F6",X"14",X"F8",X"73",X"F9",X"C8",X"FA",X"13",X"FC",X"53",X"FD",X"8A",X"FE",X"B6",X"FF",
		X"D8",X"00",X"EF",X"01",X"FF",X"02",X"06",X"04",X"02",X"05",X"F7",X"05",X"E2",X"06",X"C6",X"07",
		X"A3",X"08",X"72",X"09",X"CC",X"09",X"AD",X"09",X"47",X"09",X"AE",X"08",X"F4",X"07",X"25",X"07",
		X"4F",X"06",X"72",X"05",X"92",X"04",X"B7",X"03",X"DE",X"02",X"09",X"02",X"39",X"01",X"6F",X"00",
		X"AC",X"FF",X"EC",X"FE",X"37",X"FE",X"85",X"FD",X"D8",X"FC",X"31",X"FC",X"90",X"FB",X"F7",X"FA",
		X"5F",X"FA",X"CF",X"F9",X"44",X"F9",X"BD",X"F8",X"3B",X"F8",X"BE",X"F7",X"46",X"F7",X"D2",X"F6",
		X"61",X"F6",X"F6",X"F5",X"8E",X"F5",X"2B",X"F5",X"C9",X"F4",X"6F",X"F4",X"14",X"F4",X"BD",X"F3",
		X"6C",X"F3",X"1E",X"F3",X"D1",X"F2",X"88",X"F2",X"42",X"F2",X"FF",X"F1",X"BE",X"F1",X"81",X"F1",
		X"45",X"F1",X"0C",X"F1",X"D5",X"F0",X"A3",X"F0",X"70",X"F0",X"42",X"F0",X"13",X"F0",X"E9",X"EF",
		X"BF",X"EF",X"F8",X"EF",X"A5",X"F0",X"98",X"F1",X"BC",X"F2",X"FB",X"F3",X"4C",X"F5",X"A2",X"F6",
		X"F9",X"F7",X"4D",X"F9",X"9D",X"FA",X"E5",X"FB",X"25",X"FD",X"5C",X"FE",X"8B",X"FF",X"AF",X"00",
		X"CB",X"01",X"DF",X"02",X"E8",X"03",X"E9",X"04",X"E1",X"05",X"D2",X"06",X"B7",X"07",X"9A",X"08",
		X"70",X"09",X"40",X"0A",X"08",X"0B",X"CC",X"0B",X"6D",X"0C",X"8A",X"0C",X"47",X"0C",X"C4",X"0B",
		X"16",X"0B",X"50",X"0A",X"79",X"09",X"9C",X"08",X"B9",X"07",X"D8",X"06",X"F6",X"05",X"1D",X"05",
		X"47",X"04",X"76",X"03",X"AB",X"02",X"E6",X"01",X"28",X"01",X"6D",X"00",X"BD",X"FF",X"10",X"FF",
		X"68",X"FE",X"C6",X"FD",X"2C",X"FD",X"93",X"FC",X"03",X"FC",X"76",X"FB",X"F0",X"FA",X"6B",X"FA",
		X"38",X"FA",X"82",X"FA",X"16",X"FB",X"DE",X"FB",X"C5",X"FC",X"C0",X"FD",X"C3",X"FE",X"CB",X"FF",
		X"D2",X"00",X"D7",X"01",X"D9",X"02",X"D2",X"03",X"C8",X"04",X"B4",X"05",X"9B",X"06",X"7A",X"07",
		X"51",X"08",X"21",X"09",X"EA",X"09",X"AC",X"0A",X"68",X"0B",X"1D",X"0C",X"CA",X"0C",X"73",X"0D",
		X"15",X"0E",X"B2",X"0E",X"48",X"0F",X"DA",X"0F",X"64",X"10",X"EB",X"10",X"6C",X"11",X"E9",X"11",
		X"60",X"12",X"D4",X"12",X"41",X"13",X"AC",X"13",X"12",X"14",X"74",X"14",X"D3",X"14",X"2D",X"15",
		X"83",X"15",X"D6",X"15",X"25",X"16",X"71",X"16",X"BA",X"16",X"00",X"17",X"43",X"17",X"82",X"17",
		X"BF",X"17",X"F7",X"17",X"31",X"18",X"64",X"18",X"97",X"18",X"C4",X"18",X"F6",X"18",X"E5",X"18",
		X"5D",X"18",X"88",X"17",X"7F",X"16",X"58",X"15",X"1F",X"14",X"DF",X"12",X"9A",X"11",X"58",X"10",
		X"19",X"0F",X"E1",X"0D",X"AF",X"0C",X"88",X"0B",X"66",X"0A",X"4D",X"09",X"3C",X"08",X"36",X"07",
		X"35",X"06",X"40",X"05",X"50",X"04",X"69",X"03",X"8A",X"02",X"B1",X"01",X"E0",X"00",X"18",X"00",
		X"55",X"FF",X"99",X"FE",X"EA",X"FD",X"AC",X"FD",X"D6",X"FD",X"41",X"FE",X"DA",X"FE",X"8E",X"FF",
		X"53",X"00",X"20",X"01",X"F3",X"01",X"C5",X"02",X"96",X"03",X"60",X"04",X"2A",X"05",X"EC",X"05",
		X"AA",X"06",X"62",X"07",X"12",X"08",X"BF",X"08",X"64",X"09",X"06",X"0A",X"A1",X"0A",X"36",X"0B",
		X"C6",X"0B",X"50",X"0C",X"D7",X"0C",X"57",X"0D",X"D4",X"0D",X"49",X"0E",X"BD",X"0E",X"2B",X"0F",
		X"96",X"0F",X"FB",X"0F",X"5F",X"10",X"BD",X"10",X"17",X"11",X"6E",X"11",X"C2",X"11",X"13",X"12",
		X"5F",X"12",X"A7",X"12",X"F0",X"12",X"31",X"13",X"74",X"13",X"B1",X"13",X"ED",X"13",X"24",X"14",
		X"5B",X"14",X"8D",X"14",X"BF",X"14",X"EE",X"14",X"1B",X"15",X"44",X"15",X"6F",X"15",X"92",X"15",
		X"BA",X"15",X"BC",X"15",X"48",X"15",X"82",X"14",X"86",X"13",X"69",X"12",X"39",X"11",X"01",X"10",
		X"C3",X"0E",X"8A",X"0D",X"51",X"0C",X"1E",X"0B",X"F1",X"09",X"CC",X"08",X"B1",X"07",X"9E",X"06",
		X"93",X"05",X"90",X"04",X"96",X"03",X"A2",X"02",X"B7",X"01",X"D4",X"00",X"FB",X"FF",X"28",X"FF",
		X"59",X"FE",X"95",X"FD",X"D5",X"FC",X"1E",X"FC",X"6A",X"FB",X"0F",X"FB",X"24",X"FB",X"7C",X"FB",
		X"07",X"FC",X"AC",X"FC",X"67",X"FD",X"2B",X"FE",X"F3",X"FE",X"BB",X"FF",X"84",X"00",X"48",X"01",
		X"0A",X"02",X"C6",X"02",X"7C",X"03",X"2D",X"04",X"D9",X"04",X"7D",X"05",X"21",X"06",X"BC",X"06",
		X"51",X"07",X"E2",X"07",X"6E",X"08",X"F4",X"08",X"78",X"09",X"F3",X"09",X"6D",X"0A",X"E2",X"0A",
		X"51",X"0B",X"BD",X"0B",X"23",X"0C",X"88",X"0C",X"E7",X"0C",X"44",X"0D",X"9E",X"0D",X"F3",X"0D",
		X"43",X"0E",X"93",X"0E",X"DE",X"0E",X"27",X"0F",X"6B",X"0F",X"AF",X"0F",X"EF",X"0F",X"2C",X"10",
		X"66",X"10",X"9F",X"10",X"D4",X"10",X"06",X"11",X"38",X"11",X"66",X"11",X"93",X"11",X"BF",X"11",
		X"E7",X"11",X"0C",X"12",X"30",X"12",X"53",X"12",X"76",X"12",X"93",X"12",X"B1",X"12",X"CD",X"12",
		X"E7",X"12",X"00",X"13",X"17",X"13",X"2C",X"13",X"41",X"13",X"54",X"13",X"67",X"13",X"77",X"13",
		X"86",X"13",X"96",X"13",X"A1",X"13",X"AD",X"13",X"B8",X"13",X"C2",X"13",X"CA",X"13",X"D2",X"13",
		X"DA",X"13",X"E1",X"13",X"E6",X"13",X"E8",X"13",X"ED",X"13",X"EE",X"13",X"F3",X"13",X"E8",X"13",
		X"76",X"13",X"AC",X"12",X"AC",X"11",X"8B",X"10",X"52",X"0F",X"12",X"0E",X"CB",X"0C",X"9D",X"0B",
		X"68",X"0A",X"24",X"09",X"F1",X"07",X"C0",X"06",X"9C",X"05",X"7E",X"04",X"69",X"03",X"5D",X"02",
		X"5C",X"01",X"60",X"00",X"6F",X"FF",X"84",X"FE",X"A3",X"FD",X"C6",X"FC",X"F3",X"FB",X"27",X"FB",
		X"61",X"FA",X"A3",X"F9",X"E9",X"F8",X"68",X"F8",X"5B",X"F8",X"98",X"F8",X"08",X"F9",X"97",X"F9",
		X"3B",X"FA",X"EA",X"FA",X"A2",X"FB",X"58",X"FC",X"12",X"FD",X"C7",X"FD",X"7A",X"FE",X"28",X"FF",
		X"D2",X"FF",X"74",X"00",X"15",X"01",X"AD",X"01",X"44",X"02",X"D4",X"02",X"61",X"03",X"E7",X"03",
		X"6A",X"04",X"E8",X"04",X"61",X"05",X"D8",X"05",X"48",X"06",X"B4",X"06",X"17",X"07",X"1B",X"07",
		X"BF",X"06",X"29",X"06",X"6A",X"05",X"94",X"04",X"B0",X"03",X"C5",X"02",X"D8",X"01",X"EB",X"00",
		X"03",X"00",X"1F",X"FF",X"3F",X"FE",X"67",X"FD",X"94",X"FC",X"C7",X"FB",X"00",X"FB",X"41",X"FA",
		X"88",X"F9",X"D5",X"F8",X"29",X"F8",X"83",X"F7",X"E2",X"F6",X"45",X"F6",X"B0",X"F5",X"1F",X"F5",
		X"96",X"F4",X"0B",X"F4",X"AD",X"F3",X"C0",X"F3",X"1C",X"F4",X"AC",X"F4",X"5C",X"F5",X"20",X"F6",
		X"EF",X"F6",X"C3",X"F7",X"98",X"F8",X"6D",X"F9",X"3D",X"FA",X"0C",X"FB",X"D4",X"FB",X"96",X"FC",
		X"53",X"FD",X"0C",X"FE",X"BE",X"FE",X"6A",X"FF",X"10",X"00",X"B1",X"00",X"4C",X"01",X"E2",X"01",
		X"74",X"02",X"00",X"03",X"87",X"03",X"0C",X"04",X"86",X"04",X"FF",X"04",X"24",X"05",X"E5",X"04",
		X"6C",X"04",X"C7",X"03",X"0A",X"03",X"3C",X"02",X"69",X"01",X"91",X"00",X"BA",X"FF",X"E4",X"FE",
		X"14",X"FE",X"48",X"FD",X"81",X"FC",X"C0",X"FB",X"04",X"FB",X"4F",X"FA",X"9E",X"F9",X"F5",X"F8",
		X"50",X"F8",X"B3",X"F7",X"19",X"F7",X"86",X"F6",X"F8",X"F5",X"70",X"F5",X"EB",X"F4",X"6C",X"F4",
		X"EF",X"F3",X"90",X"F3",X"9C",X"F3",X"F8",X"F3",X"85",X"F4",X"34",X"F5",X"F6",X"F5",X"C4",X"F6",
		X"99",X"F7",X"70",X"F8",X"45",X"F9",X"16",X"FA",X"E4",X"FA",X"AC",X"FB",X"6F",X"FC",X"2D",X"FD",
		X"E4",X"FD",X"98",X"FE",X"44",X"FF",X"EB",X"FF",X"8C",X"00",X"28",X"01",X"C0",X"01",X"51",X"02",
		X"DD",X"02",X"64",X"03",X"E8",X"03",X"66",X"04",X"E1",X"04",X"57",X"05",X"C7",X"05",X"35",X"06",
		X"9E",X"06",X"05",X"07",X"67",X"07",X"C5",X"07",X"1F",X"08",X"77",X"08",X"CC",X"08",X"1D",X"09",
		X"69",X"09",X"B5",X"09",X"FC",X"09",X"42",X"0A",X"85",X"0A",X"C5",X"0A",X"01",X"0B",X"3D",X"0B",
		X"76",X"0B",X"AE",X"0B",X"E1",X"0B",X"13",X"0C",X"42",X"0C",X"70",X"0C",X"9A",X"0C",X"C4",X"0C",
		X"EE",X"0C",X"15",X"0D",X"36",X"0D",X"59",X"0D",X"79",X"0D",X"9A",X"0D",X"B6",X"0D",X"D4",X"0D",
		X"EF",X"0D",X"07",X"0E",X"20",X"0E",X"38",X"0E",X"4D",X"0E",X"62",X"0E",X"74",X"0E",X"87",X"0E",
		X"96",X"0E",X"A6",X"0E",X"B4",X"0E",X"C2",X"0E",X"CF",X"0E",X"DA",X"0E",X"E5",X"0E",X"EE",X"0E",
		X"F8",X"0E",X"01",X"0F",X"08",X"0F",X"0E",X"0F",X"14",X"0F",X"19",X"0F",X"1E",X"0F",X"21",X"0F",
		X"25",X"0F",X"27",X"0F",X"27",X"0F",X"29",X"0F",X"2B",X"0F",X"2A",X"0F",X"29",X"0F",X"28",X"0F",
		X"26",X"0F",X"24",X"0F",X"22",X"0F",X"1E",X"0F",X"1A",X"0F",X"16",X"0F",X"13",X"0F",X"0E",X"0F",
		X"08",X"0F",X"03",X"0F",X"FE",X"0E",X"F7",X"0E",X"F2",X"0E",X"EA",X"0E",X"E3",X"0E",X"D4",X"0E",
		X"6E",X"0E",X"B6",X"0D",X"CF",X"0C",X"C8",X"0B",X"AD",X"0A",X"8A",X"09",X"64",X"08",X"3F",X"07",
		X"1C",X"06",X"FF",X"04",X"E9",X"03",X"DA",X"02",X"D3",X"01",X"D2",X"00",X"DD",X"FF",X"ED",X"FE",
		X"03",X"FE",X"23",X"FD",X"4B",X"FC",X"78",X"FB",X"AF",X"FA",X"EB",X"F9",X"2F",X"F9",X"78",X"F8",
		X"C7",X"F7",X"1E",X"F7",X"7B",X"F6",X"DC",X"F5",X"45",X"F5",X"B0",X"F4",X"24",X"F4",X"9B",X"F3",
		X"17",X"F3",X"98",X"F2",X"1E",X"F2",X"A9",X"F1",X"38",X"F1",X"CB",X"F0",X"61",X"F0",X"FD",X"EF",
		X"9B",X"EF",X"3F",X"EF",X"E6",X"EE",X"8F",X"EE",X"3E",X"EE",X"EE",X"ED",X"A2",X"ED",X"5B",X"ED",
		X"14",X"ED",X"D2",X"EC",X"91",X"EC",X"54",X"EC",X"1A",X"EC",X"E2",X"EB",X"AD",X"EB",X"CB",X"EB",
		X"3D",X"EC",X"E2",X"EC",X"AC",X"ED",X"87",X"EE",X"70",X"EF",X"5F",X"F0",X"50",X"F1",X"3D",X"F2",
		X"29",X"F3",X"0F",X"F4",X"F0",X"F4",X"CA",X"F5",X"A0",X"F6",X"6F",X"F7",X"39",X"F8",X"FA",X"F8",
		X"B6",X"F9",X"6C",X"FA",X"1D",X"FB",X"C7",X"FB",X"6B",X"FC",X"0A",X"FD",X"A5",X"FD",X"3A",X"FE",
		X"CA",X"FE",X"53",X"FF",X"DA",X"FF",X"5A",X"00",X"D8",X"00",X"50",X"01",X"C4",X"01",X"35",X"02",
		X"A3",X"02",X"0B",X"03",X"70",X"03",X"D2",X"03",X"30",X"04",X"8A",X"04",X"E3",X"04",X"35",X"05",
		X"87",X"05",X"D6",X"05",X"21",X"06",X"69",X"06",X"AF",X"06",X"F2",X"06",X"33",X"07",X"70",X"07",
		X"AD",X"07",X"E6",X"07",X"1D",X"08",X"52",X"08",X"86",X"08",X"A6",X"08",X"68",X"08",X"E6",X"07",
		X"35",X"07",X"6A",X"06",X"8D",X"05",X"A9",X"04",X"C2",X"03",X"D7",X"02",X"F2",X"01",X"11",X"01",
		X"36",X"00",X"5E",X"FF",X"8C",X"FE",X"C2",X"FD",X"FD",X"FC",X"3F",X"FC",X"86",X"FB",X"D6",X"FA",
		X"29",X"FA",X"83",X"F9",X"E3",X"F8",X"48",X"F8",X"B4",X"F7",X"23",X"F7",X"98",X"F6",X"12",X"F6",
		X"92",X"F5",X"15",X"F5",X"9E",X"F4",X"29",X"F4",X"BB",X"F3",X"50",X"F3",X"E8",X"F2",X"85",X"F2",
		X"25",X"F2",X"C9",X"F1",X"71",X"F1",X"1D",X"F1",X"CB",X"F0",X"7D",X"F0",X"32",X"F0",X"E8",X"EF",
		X"A2",X"EF",X"61",X"EF",X"23",X"EF",X"E4",X"EE",X"AB",X"EE",X"74",X"EE",X"3F",X"EE",X"0B",X"EE",
		X"DA",X"ED",X"AC",X"ED",X"7F",X"ED",X"55",X"ED",X"2E",X"ED",X"07",X"ED",X"E2",X"EC",X"BF",X"EC",
		X"9F",X"EC",X"80",X"EC",X"63",X"EC",X"47",X"EC",X"2B",X"EC",X"13",X"EC",X"FD",X"EB",X"E6",X"EB",
		X"D2",X"EB",X"BF",X"EB",X"AD",X"EB",X"9C",X"EB",X"8C",X"EB",X"7F",X"EB",X"73",X"EB",X"66",X"EB",
		X"5B",X"EB",X"52",X"EB",X"48",X"EB",X"41",X"EB",X"3A",X"EB",X"34",X"EB",X"2E",X"EB",X"29",X"EB",
		X"4D",X"EB",X"CA",X"EB",X"7E",X"EC",X"58",X"ED",X"44",X"EE",X"40",X"EF",X"3E",X"F0",X"44",X"F1",
		X"29",X"F2",X"18",X"F3",X"16",X"F4",X"07",X"F5",X"F7",X"F5",X"DB",X"F6",X"BD",X"F7",X"95",X"F8",
		X"68",X"F9",X"33",X"FA",X"F7",X"FA",X"B6",X"FB",X"70",X"FC",X"20",X"FD",X"CC",X"FD",X"73",X"FE",
		X"14",X"FF",X"AE",X"FF",X"45",X"00",X"CF",X"00",X"0C",X"01",X"F9",X"00",X"B7",X"00",X"50",X"00",
		X"D8",X"FF",X"52",X"FF",X"C5",X"FE",X"35",X"FE",X"A5",X"FD",X"15",X"FD",X"86",X"FC",X"FC",X"FB",
		X"75",X"FB",X"F2",X"FA",X"74",X"FA",X"F8",X"F9",X"82",X"F9",X"0E",X"F9",X"9F",X"F8",X"34",X"F8",
		X"CE",X"F7",X"69",X"F7",X"0A",X"F7",X"AF",X"F6",X"55",X"F6",X"00",X"F6",X"AC",X"F5",X"5D",X"F5",
		X"12",X"F5",X"C9",X"F4",X"83",X"F4",X"3E",X"F4",X"FD",X"F3",X"C0",X"F3",X"84",X"F3",X"4A",X"F3",
		X"14",X"F3",X"DF",X"F2",X"AD",X"F2",X"7C",X"F2",X"4C",X"F2",X"22",X"F2",X"F7",X"F1",X"CF",X"F1",
		X"A8",X"F1",X"83",X"F1",X"61",X"F1",X"3F",X"F1",X"1E",X"F1",X"00",X"F1",X"E4",X"F0",X"C9",X"F0",
		X"AE",X"F0",X"98",X"F0",X"83",X"F0",X"AF",X"F0",X"29",X"F1",X"D1",X"F1",X"98",X"F2",X"71",X"F3",
		X"53",X"F4",X"3B",X"F5",X"23",X"F6",X"09",X"F7",X"EB",X"F7",X"C9",X"F8",X"A2",X"F9",X"76",X"FA",
		X"42",X"FB",X"07",X"FC",X"C6",X"FC",X"81",X"FD",X"34",X"FE",X"E3",X"FE",X"8D",X"FF",X"2D",X"00",
		X"CA",X"00",X"63",X"01",X"F5",X"01",X"84",X"02",X"0C",X"03",X"92",X"03",X"FE",X"03",X"12",X"04",
		X"E6",X"03",X"92",X"03",X"21",X"03",X"A2",X"02",X"19",X"02",X"8A",X"01",X"F9",X"00",X"67",X"00",
		X"D8",X"FF",X"4D",X"FF",X"C3",X"FE",X"3D",X"FE",X"BA",X"FD",X"3C",X"FD",X"C5",X"FC",X"4E",X"FC",
		X"DC",X"FB",X"6E",X"FB",X"03",X"FB",X"9C",X"FA",X"39",X"FA",X"DA",X"F9",X"7F",X"F9",X"24",X"F9",
		X"CF",X"F8",X"7E",X"F8",X"2E",X"F8",X"E2",X"F7",X"99",X"F7",X"51",X"F7",X"0F",X"F7",X"CC",X"F6",
		X"8E",X"F6",X"52",X"F6",X"19",X"F6",X"E1",X"F5",X"AD",X"F5",X"79",X"F5",X"48",X"F5",X"18",X"F5",
		X"EA",X"F4",X"C1",X"F4",X"97",X"F4",X"70",X"F4",X"4A",X"F4",X"25",X"F4",X"04",X"F4",X"E3",X"F3",
		X"C4",X"F3",X"A6",X"F3",X"8A",X"F3",X"6F",X"F3",X"55",X"F3",X"3D",X"F3",X"25",X"F3",X"10",X"F3",
		X"FB",X"F2",X"E8",X"F2",X"D5",X"F2",X"C3",X"F2",X"B2",X"F2",X"A3",X"F2",X"97",X"F2",X"89",X"F2",
		X"7D",X"F2",X"72",X"F2",X"67",X"F2",X"5C",X"F2",X"54",X"F2",X"4C",X"F2",X"45",X"F2",X"3E",X"F2",
		X"38",X"F2",X"33",X"F2",X"2E",X"F2",X"2B",X"F2",X"28",X"F2",X"24",X"F2",X"22",X"F2",X"20",X"F2",
		X"20",X"F2",X"20",X"F2",X"1F",X"F2",X"20",X"F2",X"21",X"F2",X"22",X"F2",X"24",X"F2",X"27",X"F2",
		X"2A",X"F2",X"2D",X"F2",X"31",X"F2",X"35",X"F2",X"38",X"F2",X"3D",X"F2",X"43",X"F2",X"48",X"F2",
		X"4D",X"F2",X"53",X"F2",X"5B",X"F2",X"60",X"F2",X"67",X"F2",X"6E",X"F2",X"74",X"F2",X"7D",X"F2",
		X"85",X"F2",X"8D",X"F2",X"95",X"F2",X"9E",X"F2",X"AD",X"F2",X"02",X"F3",X"96",X"F3",X"51",X"F4",
		X"28",X"F5",X"09",X"F6",X"F3",X"F6",X"DF",X"F7",X"CA",X"F8",X"B3",X"F9",X"97",X"FA",X"77",X"FB",
		X"4F",X"FC",X"23",X"FD",X"F1",X"FD",X"B6",X"FE",X"74",X"FF",X"30",X"00",X"E3",X"00",X"91",X"01",
		X"39",X"02",X"DC",X"02",X"78",X"03",X"11",X"04",X"A2",X"04",X"31",X"05",X"B7",X"05",X"3F",X"06",
		X"9D",X"06",X"AB",X"06",X"88",X"06",X"3E",X"06",X"DC",X"05",X"6E",X"05",X"F6",X"04",X"7A",X"04",
		X"FD",X"03",X"7F",X"03",X"03",X"03",X"88",X"02",X"12",X"02",X"9E",X"01",X"2D",X"01",X"C1",X"00",
		X"57",X"00",X"F1",X"FF",X"8E",X"FF",X"2D",X"FF",X"CF",X"FE",X"77",X"FE",X"20",X"FE",X"CD",X"FD",
		X"7C",X"FD",X"2F",X"FD",X"E5",X"FC",X"9F",X"FC",X"9A",X"FC",X"D9",X"FC",X"40",X"FD",X"C5",X"FD",
		X"58",X"FE",X"F6",X"FE",X"99",X"FF",X"3F",X"00",X"E1",X"00",X"83",X"01",X"21",X"02",X"BC",X"02",
		X"53",X"03",X"E5",X"03",X"72",X"04",X"FB",X"04",X"7F",X"05",X"00",X"06",X"7A",X"06",X"F4",X"06",
		X"67",X"07",X"D4",X"07",X"40",X"08",X"A8",X"08",X"0B",X"09",X"6B",X"09",X"C7",X"09",X"21",X"0A",
		X"76",X"0A",X"CA",X"0A",X"19",X"0B",X"65",X"0B",X"AE",X"0B",X"F4",X"0B",X"38",X"0C",X"7A",X"0C",
		X"B7",X"0C",X"F4",X"0C",X"2E",X"0D",X"64",X"0D",X"9A",X"0D",X"CB",X"0D",X"FE",X"0D",X"2B",X"0E",
		X"59",X"0E",X"82",X"0E",X"AB",X"0E",X"D1",X"0E",X"F6",X"0E",X"1A",X"0F",X"3C",X"0F",X"5B",X"0F",
		X"7B",X"0F",X"95",X"0F",X"B2",X"0F",X"98",X"0F",X"37",X"0F",X"B4",X"0E",X"0F",X"0E",X"5E",X"0D",
		X"A1",X"0C",X"E3",X"0B",X"21",X"0B",X"62",X"0A",X"A5",X"09",X"EC",X"08",X"35",X"08",X"87",X"07",
		X"DA",X"06",X"35",X"06",X"94",X"05",X"F8",X"04",X"61",X"04",X"D0",X"03",X"43",X"03",X"B9",X"02",
		X"37",X"02",X"B6",X"01",X"3C",X"01",X"C2",X"00",X"51",X"00",X"E2",X"FF",X"A3",X"FF",X"AB",X"FF",
		X"DD",X"FF",X"2F",X"00",X"94",X"00",X"05",X"01",X"7E",X"01",X"F8",X"01",X"75",X"02",X"EF",X"02",
		X"69",X"03",X"E1",X"03",X"52",X"04",X"C3",X"04",X"31",X"05",X"9B",X"05",X"FF",X"05",X"62",X"06",
		X"C1",X"06",X"1E",X"07",X"75",X"07",X"CC",X"07",X"1D",X"08",X"6C",X"08",X"BA",X"08",X"01",X"09",
		X"48",X"09",X"8C",X"09",X"CE",X"09",X"0D",X"0A",X"49",X"0A",X"83",X"0A",X"BA",X"0A",X"F0",X"0A",
		X"24",X"0B",X"55",X"0B",X"85",X"0B",X"B2",X"0B",X"DD",X"0B",X"06",X"0C",X"2E",X"0C",X"52",X"0C",
		X"78",X"0C",X"99",X"0C",X"BB",X"0C",X"DB",X"0C",X"F8",X"0C",X"16",X"0D",X"30",X"0D",X"4A",X"0D",
		X"63",X"0D",X"78",X"0D",X"90",X"0D",X"A5",X"0D",X"BA",X"0D",X"AB",X"0D",X"57",X"0D",X"DA",X"0C",
		X"40",X"0C",X"94",X"0B",X"DE",X"0A",X"24",X"0A",X"69",X"09",X"AF",X"08",X"F7",X"07",X"42",X"07",
		X"92",X"06",X"E8",X"05",X"40",X"05",X"9F",X"04",X"03",X"04",X"6A",X"03",X"D8",X"02",X"4A",X"02",
		X"C1",X"01",X"3B",X"01",X"BB",X"00",X"40",X"00",X"CA",X"FF",X"55",X"FF",X"E4",X"FE",X"79",X"FE",
		X"11",X"FE",X"AC",X"FD",X"4B",X"FD",X"EE",X"FC",X"93",X"FC",X"3B",X"FC",X"E9",X"FB",X"99",X"FB",
		X"4A",X"FB",X"F6",X"FA",X"A6",X"FA",X"62",X"FA",X"1F",X"FA",X"DC",X"F9",X"9E",X"F9",X"61",X"F9",
		X"28",X"F9",X"F0",X"F8",X"B9",X"F8",X"86",X"F8",X"54",X"F8",X"24",X"F8",X"F6",X"F7",X"CB",X"F7",
		X"A0",X"F7",X"78",X"F7",X"51",X"F7",X"2C",X"F7",X"07",X"F7",X"E7",X"F6",X"C5",X"F6",X"A7",X"F6",
		X"88",X"F6",X"6C",X"F6",X"50",X"F6",X"37",X"F6",X"21",X"F6",X"08",X"F6",X"F2",X"F5",X"DD",X"F5",
		X"CA",X"F5",X"B7",X"F5",X"A4",X"F5",X"93",X"F5",X"83",X"F5",X"74",X"F5",X"67",X"F5",X"59",X"F5",
		X"4D",X"F5",X"41",X"F5",X"37",X"F5",X"2D",X"F5",X"24",X"F5",X"1C",X"F5",X"14",X"F5",X"0C",X"F5",
		X"06",X"F5",X"00",X"F5",X"FA",X"F4",X"F6",X"F4",X"F1",X"F4",X"EE",X"F4",X"EB",X"F4",X"E9",X"F4",
		X"E6",X"F4",X"E4",X"F4",X"E3",X"F4",X"E4",X"F4",X"E3",X"F4",X"E2",X"F4",X"E2",X"F4",X"E5",X"F4",
		X"E7",X"F4",X"E7",X"F4",X"EA",X"F4",X"EC",X"F4",X"EF",X"F4",X"F2",X"F4",X"F6",X"F4",X"F9",X"F4",
		X"FE",X"F4",X"02",X"F5",X"07",X"F5",X"0C",X"F5",X"10",X"F5",X"17",X"F5",X"1C",X"F5",X"21",X"F5",
		X"27",X"F5",X"2F",X"F5",X"34",X"F5",X"39",X"F5",X"42",X"F5",X"48",X"F5",X"51",X"F5",X"57",X"F5",
		X"5E",X"F5",X"66",X"F5",X"6F",X"F5",X"77",X"F5",X"80",X"F5",X"88",X"F5",X"8E",X"F5",X"97",X"F5",
		X"9F",X"F5",X"A7",X"F5",X"B1",X"F5",X"BB",X"F5",X"C3",X"F5",X"CB",X"F5",X"D6",X"F5",X"DF",X"F5",
		X"EA",X"F5",X"F2",X"F5",X"FC",X"F5",X"05",X"F6",X"0F",X"F6",X"18",X"F6",X"24",X"F6",X"2C",X"F6",
		X"36",X"F6",X"40",X"F6",X"4A",X"F6",X"54",X"F6",X"5E",X"F6",X"68",X"F6",X"72",X"F6",X"7D",X"F6",
		X"86",X"F6",X"92",X"F6",X"9B",X"F6",X"A6",X"F6",X"B0",X"F6",X"BB",X"F6",X"C5",X"F6",X"D0",X"F6",
		X"DA",X"F6",X"E5",X"F6",X"FA",X"F6",X"4A",X"F7",X"C8",X"F7",X"63",X"F8",X"0F",X"F9",X"C5",X"F9",
		X"82",X"FA",X"3F",X"FB",X"FB",X"FB",X"B5",X"FC",X"6B",X"FD",X"1B",X"FE",X"CA",X"FE",X"72",X"FF",
		X"13",X"00",X"B1",X"00",X"49",X"01",X"DD",X"01",X"6C",X"02",X"F6",X"02",X"7B",X"03",X"FB",X"03",
		X"78",X"04",X"F0",X"04",X"65",X"05",X"D3",X"05",X"3F",X"06",X"A7",X"06",X"0C",X"07",X"6C",X"07",
		X"CA",X"07",X"23",X"08",X"7A",X"08",X"CD",X"08",X"1E",X"09",X"6B",X"09",X"B6",X"09",X"FD",X"09",
		X"42",X"0A",X"84",X"0A",X"C3",X"0A",X"01",X"0B",X"3B",X"0B",X"74",X"0B",X"AA",X"0B",X"DE",X"0B",
		X"0F",X"0C",X"3F",X"0C",X"6C",X"0C",X"9A",X"0C",X"C4",X"0C",X"EA",X"0C",X"12",X"0D",X"36",X"0D",
		X"59",X"0D",X"7B",X"0D",X"9A",X"0D",X"B9",X"0D",X"D6",X"0D",X"F2",X"0D",X"0B",X"0E",X"24",X"0E",
		X"3B",X"0E",X"52",X"0E",X"67",X"0E",X"7B",X"0E",X"8E",X"0E",X"9F",X"0E",X"B0",X"0E",X"BF",X"0E",
		X"CD",X"0E",X"DB",X"0E",X"E8",X"0E",X"F5",X"0E",X"00",X"0F",X"09",X"0F",X"13",X"0F",X"1B",X"0F",
		X"22",X"0F",X"2A",X"0F",X"31",X"0F",X"35",X"0F",X"39",X"0F",X"3F",X"0F",X"41",X"0F",X"45",X"0F",
		X"47",X"0F",X"49",X"0F",X"4A",X"0F",X"4C",X"0F",X"4C",X"0F",X"4B",X"0F",X"4A",X"0F",X"4A",X"0F",
		X"47",X"0F",X"46",X"0F",X"43",X"0F",X"41",X"0F",X"3C",X"0F",X"39",X"0F",X"37",X"0F",X"30",X"0F",
		X"2B",X"0F",X"27",X"0F",X"22",X"0F",X"1B",X"0F",X"15",X"0F",X"10",X"0F",X"09",X"0F",X"02",X"0F",
		X"F9",X"0E",X"BF",X"0E",X"55",X"0E",X"CF",X"0D",X"36",X"0D",X"91",X"0C",X"E6",X"0B",X"3A",X"0B",
		X"8D",X"0A",X"E3",X"09",X"3D",X"09",X"99",X"08",X"FA",X"07",X"5E",X"07",X"C7",X"06",X"35",X"06",
		X"A8",X"05",X"1F",X"05",X"9A",X"04",X"19",X"04",X"9D",X"03",X"26",X"03",X"B1",X"02",X"41",X"02",
		X"D4",X"01",X"6B",X"01",X"07",X"01",X"A3",X"00",X"47",X"00",X"EC",X"FF",X"94",X"FF",X"3E",X"FF",
		X"EC",X"FE",X"9D",X"FE",X"50",X"FE",X"06",X"FE",X"BF",X"FD",X"7A",X"FD",X"3A",X"FD",X"F9",X"FC",
		X"BA",X"FC",X"82",X"FC",X"49",X"FC",X"10",X"FC",X"DB",X"FB",X"A8",X"FB",X"79",X"FB",X"49",X"FB",
		X"1D",X"FB",X"EF",X"FA",X"C7",X"FA",X"9D",X"FA",X"76",X"FA",X"51",X"FA",X"2D",X"FA",X"0C",X"FA",
		X"13",X"FA",X"4C",X"FA",X"A7",X"FA",X"13",X"FB",X"8C",X"FB",X"0C",X"FC",X"90",X"FC",X"14",X"FD",
		X"96",X"FD",X"17",X"FE",X"96",X"FE",X"13",X"FF",X"8C",X"FF",X"00",X"00",X"72",X"00",X"DE",X"00",
		X"4A",X"01",X"AF",X"01",X"13",X"02",X"75",X"02",X"D1",X"02",X"2B",X"03",X"80",X"03",X"D4",X"03",
		X"24",X"04",X"73",X"04",X"BC",X"04",X"04",X"05",X"4B",X"05",X"8D",X"05",X"CF",X"05",X"0D",X"06",
		X"47",X"06",X"82",X"06",X"B8",X"06",X"F0",X"06",X"22",X"07",X"55",X"07",X"82",X"07",X"B0",X"07",
		X"DD",X"07",X"07",X"08",X"2E",X"08",X"56",X"08",X"79",X"08",X"9E",X"08",X"BF",X"08",X"E1",X"08",
		X"FF",X"08",X"1F",X"09",X"38",X"09",X"55",X"09",X"6F",X"09",X"8A",X"09",X"9A",X"09",X"77",X"09",
		X"2E",X"09",X"C9",X"08",X"55",X"08",X"D9",X"07",X"55",X"07",X"CF",X"06",X"4A",X"06",X"C6",X"05",
		X"45",X"05",X"C5",X"04",X"4A",X"04",X"D2",X"03",X"5D",X"03",X"EC",X"02",X"7D",X"02",X"14",X"02",
		X"AD",X"01",X"4A",X"01",X"E9",X"00",X"8D",X"00",X"34",X"00",X"DE",X"FF",X"8B",X"FF",X"3A",X"FF",
		X"EC",X"FE",X"A1",X"FE",X"58",X"FE",X"13",X"FE",X"CF",X"FD",X"8E",X"FD",X"50",X"FD",X"12",X"FD",
		X"D8",X"FC",X"A1",X"FC",X"6A",X"FC",X"37",X"FC",X"04",X"FC",X"D3",X"FB",X"A6",X"FB",X"78",X"FB",
		X"4D",X"FB",X"25",X"FB",X"FC",X"FA",X"D8",X"FA",X"B2",X"FA",X"8F",X"FA",X"6C",X"FA",X"4D",X"FA",
		X"2E",X"FA",X"11",X"FA",X"F4",X"F9",X"D9",X"F9",X"BF",X"F9",X"A5",X"F9",X"8E",X"F9",X"77",X"F9",
		X"61",X"F9",X"4C",X"F9",X"39",X"F9",X"26",X"F9",X"14",X"F9",X"04",X"F9",X"F4",X"F8",X"E4",X"F8",
		X"D5",X"F8",X"C7",X"F8",X"BB",X"F8",X"AE",X"F8",X"A4",X"F8",X"99",X"F8",X"8E",X"F8",X"85",X"F8",
		X"7C",X"F8",X"74",X"F8",X"6C",X"F8",X"66",X"F8",X"5F",X"F8",X"58",X"F8",X"54",X"F8",X"4E",X"F8",
		X"49",X"F8",X"45",X"F8",X"41",X"F8",X"3F",X"F8",X"3B",X"F8",X"39",X"F8",X"38",X"F8",X"36",X"F8",
		X"34",X"F8",X"36",X"F8",X"26",X"F8",X"1D",X"F8",X"21",X"F8",X"20",X"F8",X"22",X"F8",X"21",X"F8",
		X"23",X"F8",X"25",X"F8",X"27",X"F8",X"29",X"F8",X"2C",X"F8",X"2E",X"F8",X"31",X"F8",X"34",X"F8",
		X"38",X"F8",X"3C",X"F8",X"40",X"F8",X"42",X"F8",X"46",X"F8",X"4A",X"F8",X"50",X"F8",X"55",X"F8",
		X"59",X"F8",X"5E",X"F8",X"63",X"F8",X"68",X"F8",X"6E",X"F8",X"73",X"F8",X"79",X"F8",X"7F",X"F8",
		X"84",X"F8",X"8B",X"F8",X"90",X"F8",X"97",X"F8",X"9D",X"F8",X"A4",X"F8",X"AB",X"F8",X"B1",X"F8",
		X"B7",X"F8",X"BF",X"F8",X"C6",X"F8",X"CD",X"F8",X"D3",X"F8",X"DA",X"F8",X"E3",X"F8",X"E8",X"F8",
		X"FB",X"F8",X"3F",X"F9",X"A0",X"F9",X"18",X"FA",X"98",X"FA",X"20",X"FB",X"AD",X"FB",X"3A",X"FC",
		X"C6",X"FC",X"51",X"FD",X"D8",X"FD",X"5C",X"FE",X"DB",X"FE",X"58",X"FF",X"D2",X"FF",X"45",X"00",
		X"B6",X"00",X"24",X"01",X"8E",X"01",X"F5",X"01",X"57",X"02",X"B8",X"02",X"13",X"03",X"6D",X"03",
		X"C3",X"03",X"15",X"04",X"66",X"04",X"B2",X"04",X"FC",X"04",X"44",X"05",X"89",X"05",X"CB",X"05",
		X"0C",X"06",X"49",X"06",X"85",X"06",X"BF",X"06",X"F5",X"06",X"2C",X"07",X"5E",X"07",X"90",X"07",
		X"BD",X"07",X"EB",X"07",X"18",X"08",X"41",X"08",X"68",X"08",X"8E",X"08",X"B4",X"08",X"D7",X"08",
		X"F8",X"08",X"1A",X"09",X"39",X"09",X"57",X"09",X"72",X"09",X"8E",X"09",X"A7",X"09",X"C0",X"09",
		X"D6",X"09",X"EE",X"09",X"02",X"0A",X"17",X"0A",X"2B",X"0A",X"3D",X"0A",X"4F",X"0A",X"5F",X"0A",
		X"6E",X"0A",X"7D",X"0A",X"8B",X"0A",X"99",X"0A",X"A3",X"0A",X"B0",X"0A",X"BC",X"0A",X"C6",X"0A",
		X"CE",X"0A",X"D7",X"0A",X"DF",X"0A",X"E5",X"0A",X"EB",X"0A",X"F3",X"0A",X"F8",X"0A",X"FC",X"0A",
		X"00",X"0B",X"05",X"0B",X"09",X"0B",X"0D",X"0B",X"0E",X"0B",X"11",X"0B",X"13",X"0B",X"14",X"0B",
		X"15",X"0B",X"15",X"0B",X"13",X"0B",X"15",X"0B",X"15",X"0B",X"14",X"0B",X"12",X"0B",X"11",X"0B",
		X"0D",X"0B",X"0C",X"0B",X"09",X"0B",X"06",X"0B",X"03",X"0B",X"01",X"0B",X"FC",X"0A",X"F8",X"0A",
		X"F5",X"0A",X"F0",X"0A",X"EB",X"0A",X"E6",X"0A",X"E2",X"0A",X"DD",X"0A",X"D1",X"0A",X"A1",X"0A",
		X"52",X"0A",X"EC",X"09",X"7B",X"09",X"01",X"09",X"85",X"08",X"06",X"08",X"8A",X"07",X"0D",X"07",
		X"94",X"06",X"1D",X"06",X"A7",X"05",X"38",X"05",X"CA",X"04",X"60",X"04",X"F8",X"03",X"95",X"03",
		X"35",X"03",X"D7",X"02",X"7F",X"02",X"27",X"02",X"D3",X"01",X"81",X"01",X"32",X"01",X"E6",X"00",
		X"9F",X"00",X"55",X"00",X"23",X"00",X"1C",X"00",X"2D",X"00",X"53",X"00",X"84",X"00",X"BD",X"00",
		X"F9",X"00",X"37",X"01",X"78",X"01",X"B8",X"01",X"F6",X"01",X"34",X"02",X"70",X"02",X"AA",X"02",
		X"E2",X"02",X"18",X"03",X"4D",X"03",X"81",X"03",X"B3",X"03",X"E4",X"03",X"12",X"04",X"3E",X"04",
		X"69",X"04",X"91",X"04",X"B8",X"04",X"E0",X"04",X"04",X"05",X"28",X"05",X"48",X"05",X"69",X"05",
		X"88",X"05",X"A6",X"05",X"C3",X"05",X"DE",X"05",X"F8",X"05",X"12",X"06",X"29",X"06",X"41",X"06",
		X"57",X"06",X"6D",X"06",X"81",X"06",X"94",X"06",X"A7",X"06",X"B7",X"06",X"C9",X"06",X"DA",X"06",
		X"E7",X"06",X"F6",X"06",X"03",X"07",X"10",X"07",X"1B",X"07",X"29",X"07",X"32",X"07",X"3D",X"07",
		X"47",X"07",X"4F",X"07",X"5A",X"07",X"60",X"07",X"66",X"07",X"6E",X"07",X"75",X"07",X"7A",X"07",
		X"80",X"07",X"84",X"07",X"89",X"07",X"8D",X"07",X"91",X"07",X"95",X"07",X"97",X"07",X"9B",X"07",
		X"9E",X"07",X"9E",X"07",X"A1",X"07",X"A1",X"07",X"A2",X"07",X"A2",X"07",X"A3",X"07",X"A3",X"07",
		X"A2",X"07",X"A2",X"07",X"A3",X"07",X"A1",X"07",X"9F",X"07",X"82",X"07",X"42",X"07",X"F0",X"06",
		X"8F",X"06",X"28",X"06",X"BD",X"05",X"51",X"05",X"E5",X"04",X"79",X"04",X"10",X"04",X"A7",X"03",
		X"42",X"03",X"E0",X"02",X"81",X"02",X"25",X"02",X"CC",X"01",X"76",X"01",X"22",X"01",X"D2",X"00",
		X"83",X"00",X"37",X"00",X"F0",X"FF",X"A9",X"FF",X"66",X"FF",X"24",X"FF",X"E5",X"FE",X"A7",X"FE",
		X"74",X"FE",X"67",X"FE",X"73",X"FE",X"94",X"FE",X"C0",X"FE",X"F1",X"FE",X"29",X"FF",X"62",X"FF",
		X"9D",X"FF",X"D6",X"FF",X"0F",X"00",X"48",X"00",X"80",X"00",X"B5",X"00",X"EA",X"00",X"1D",X"01",
		X"4D",X"01",X"7C",X"01",X"AB",X"01",X"D7",X"01",X"02",X"02",X"2C",X"02",X"53",X"02",X"7A",X"02",
		X"9E",X"02",X"C2",X"02",X"E4",X"02",X"06",X"03",X"23",X"03",X"42",X"03",X"60",X"03",X"7E",X"03",
		X"98",X"03",X"B1",X"03",X"CC",X"03",X"E1",X"03",X"FA",X"03",X"0F",X"04",X"25",X"04",X"39",X"04",
		X"4D",X"04",X"5F",X"04",X"6F",X"04",X"81",X"04",X"92",X"04",X"A3",X"04",X"B1",X"04",X"BE",X"04",
		X"CD",X"04",X"DA",X"04",X"E5",X"04",X"F1",X"04",X"FB",X"04",X"06",X"05",X"10",X"05",X"1A",X"05",
		X"21",X"05",X"29",X"05",X"32",X"05",X"38",X"05",X"41",X"05",X"46",X"05",X"4C",X"05",X"52",X"05",
		X"57",X"05",X"5C",X"05",X"60",X"05",X"65",X"05",X"68",X"05",X"6B",X"05",X"70",X"05",X"71",X"05",
		X"74",X"05",X"77",X"05",X"78",X"05",X"7B",X"05",X"7A",X"05",X"7B",X"05",X"7D",X"05",X"7F",X"05",
		X"7F",X"05",X"7E",X"05",X"7C",X"05",X"5A",X"05",X"21",X"05",X"D5",X"04",X"83",X"04",X"27",X"04",
		X"CB",X"03",X"6C",X"03",X"0D",X"03",X"B2",X"02",X"55",X"02",X"FC",X"01",X"A5",X"01",X"50",X"01",
		X"00",X"01",X"B0",X"00",X"64",X"00",X"19",X"00",X"D3",X"FF",X"8E",X"FF",X"4C",X"FF",X"0A",X"FF",
		X"CB",X"FE",X"90",X"FE",X"56",X"FE",X"1E",X"FE",X"E7",X"FD",X"B4",X"FD",X"8E",X"FD",X"89",X"FD",
		X"99",X"FD",X"B9",X"FD",X"E0",X"FD",X"10",X"FE",X"40",X"FE",X"73",X"FE",X"A8",X"FE",X"DC",X"FE",
		X"0E",X"FF",X"41",X"FF",X"72",X"FF",X"A2",X"FF",X"D0",X"FF",X"FC",X"FF",X"27",X"00",X"50",X"00",
		X"7A",X"00",X"A1",X"00",X"C5",X"00",X"EB",X"00",X"0E",X"01",X"30",X"01",X"50",X"01",X"70",X"01",
		X"90",X"01",X"AC",X"01",X"AF",X"01",X"95",X"01",X"6C",X"01",X"39",X"01",X"FF",X"00",X"C1",X"00",
		X"81",X"00",X"3F",X"00",X"FF",X"FF",X"C1",X"FF",X"82",X"FF",X"45",X"FF",X"08",X"FF",X"CE",X"FE",
		X"97",X"FE",X"60",X"FE",X"2E",X"FE",X"F9",X"FD",X"C9",X"FD",X"9B",X"FD",X"6D",X"FD",X"41",X"FD",
		X"18",X"FD",X"EE",X"FC",X"C8",X"FC",X"A2",X"FC",X"7F",X"FC",X"5C",X"FC",X"39",X"FC",X"1A",X"FC",
		X"FC",X"FB",X"DE",X"FB",X"C2",X"FB",X"A8",X"FB",X"8D",X"FB",X"74",X"FB",X"5D",X"FB",X"45",X"FB",
		X"2E",X"FB",X"1B",X"FB",X"05",X"FB",X"F4",X"FA",X"E1",X"FA",X"D0",X"FA",X"C0",X"FA",X"AF",X"FA",
		X"A0",X"FA",X"92",X"FA",X"85",X"FA",X"76",X"FA",X"6A",X"FA",X"5F",X"FA",X"54",X"FA",X"49",X"FA",
		X"40",X"FA",X"36",X"FA",X"2D",X"FA",X"27",X"FA",X"1F",X"FA",X"17",X"FA",X"11",X"FA",X"0B",X"FA",
		X"05",X"FA",X"00",X"FA",X"FB",X"F9",X"F7",X"F9",X"F3",X"F9",X"F0",X"F9",X"ED",X"F9",X"E9",X"F9",
		X"E7",X"F9",X"E6",X"F9",X"E3",X"F9",X"E1",X"F9",X"E0",X"F9",X"DF",X"F9",X"DF",X"F9",X"E0",X"F9",
		X"DF",X"F9",X"DF",X"F9",X"E1",X"F9",X"E0",X"F9",X"E2",X"F9",X"E3",X"F9",X"E4",X"F9",X"E6",X"F9",
		X"E6",X"F9",X"EA",X"F9",X"EB",X"F9",X"EF",X"F9",X"F1",X"F9",X"F2",X"F9",X"F5",X"F9",X"FA",X"F9",
		X"FD",X"F9",X"01",X"FA",X"04",X"FA",X"08",X"FA",X"0B",X"FA",X"10",X"FA",X"14",X"FA",X"19",X"FA",
		X"1E",X"FA",X"20",X"FA",X"25",X"FA",X"2A",X"FA",X"2E",X"FA",X"33",X"FA",X"39",X"FA",X"3D",X"FA",
		X"50",X"FA",X"7E",X"FA",X"B9",X"FA",X"00",X"FB",X"4C",X"FB",X"99",X"FB",X"E9",X"FB",X"39",X"FC",
		X"89",X"FC",X"D6",X"FC",X"23",X"FD",X"6D",X"FD",X"B5",X"FD",X"FB",X"FD",X"40",X"FE",X"80",X"FE",
		X"C2",X"FE",X"FE",X"FE",X"3A",X"FF",X"73",X"FF",X"AB",X"FF",X"E0",X"FF",X"14",X"00",X"46",X"00",
		X"77",X"00",X"A6",X"00",X"D4",X"00",X"FB",X"00",X"0C",X"01",X"06",X"01",X"F4",X"00",X"DA",X"00",
		X"BA",X"00",X"96",X"00",X"72",X"00",X"4B",X"00",X"24",X"00",X"FE",X"FF",X"DA",X"FF",X"B6",X"FF",
		X"91",X"FF",X"6F",X"FF",X"4E",X"FF",X"2D",X"FF",X"0E",X"FF",X"EF",X"FE",X"D3",X"FE",X"B7",X"FE",
		X"9C",X"FE",X"80",X"FE",X"68",X"FE",X"51",X"FE",X"3B",X"FE",X"23",X"FE",X"0F",X"FE",X"F9",X"FD",
		X"E6",X"FD",X"D5",X"FD",X"C2",X"FD",X"B1",X"FD",X"A0",X"FD",X"90",X"FD",X"81",X"FD",X"72",X"FD",
		X"66",X"FD",X"57",X"FD",X"4B",X"FD",X"3F",X"FD",X"33",X"FD",X"28",X"FD",X"1F",X"FD",X"15",X"FD",
		X"0B",X"FD",X"03",X"FD",X"FA",X"FC",X"F2",X"FC",X"EB",X"FC",X"E4",X"FC",X"DF",X"FC",X"D7",X"FC",
		X"D1",X"FC",X"CC",X"FC",X"C6",X"FC",X"D8",X"FC",X"FB",X"FC",X"2B",X"FD",X"60",X"FD",X"9C",X"FD",
		X"D8",X"FD",X"16",X"FE",X"55",X"FE",X"91",X"FE",X"CD",X"FE",X"09",X"FF",X"43",X"FF",X"7B",X"FF",
		X"B0",X"FF",X"E6",X"FF",X"17",X"00",X"4A",X"00",X"79",X"00",X"A6",X"00",X"D2",X"00",X"FE",X"00",
		X"28",X"01",X"4E",X"01",X"76",X"01",X"9A",X"01",X"BE",X"01",X"E1",X"01",X"FA",X"01",X"FE",X"01",
		X"F2",X"01",X"DB",X"01",X"BE",X"01",X"9E",X"01",X"79",X"01",X"56",X"01",X"32",X"01",X"0E",X"01",
		X"E9",X"00",X"C7",X"00",X"A3",X"00",X"82",X"00",X"60",X"00",X"42",X"00",X"23",X"00",X"07",X"00",
		X"EA",X"FF",X"D0",X"FF",X"B4",X"FF",X"9B",X"FF",X"83",X"FF",X"6C",X"FF",X"55",X"FF",X"3F",X"FF",
		X"29",X"FF",X"15",X"FF",X"12",X"FF",X"22",X"FF",X"3D",X"FF",X"61",X"FF",X"87",X"FF",X"B0",X"FF",
		X"DD",X"FF",X"09",X"00",X"34",X"00",X"5F",X"00",X"8A",X"00",X"B3",X"00",X"DC",X"00",X"03",X"01",
		X"29",X"01",X"4E",X"01",X"71",X"01",X"93",X"01",X"B2",X"01",X"D3",X"01",X"F2",X"01",X"0F",X"02",
		X"2B",X"02",X"47",X"02",X"61",X"02",X"7A",X"02",X"93",X"02",X"A6",X"02",X"A7",X"02",X"95",X"02",
		X"7D",X"02",X"5E",X"02",X"3B",X"02",X"15",X"02",X"EF",X"01",X"CB",X"01",X"A3",X"01",X"7E",X"01",
		X"5A",X"01",X"37",X"01",X"14",X"01",X"F2",X"00",X"D1",X"00",X"B3",X"00",X"93",X"00",X"77",X"00",
		X"5A",X"00",X"3F",X"00",X"24",X"00",X"0A",X"00",X"F3",X"FF",X"DC",X"FF",X"C5",X"FF",X"AF",X"FF",
		X"9A",X"FF",X"92",X"FF",X"9C",X"FF",X"AF",X"FF",X"CB",X"FF",X"EB",X"FF",X"0E",X"00",X"32",X"00",
		X"58",X"00",X"7D",X"00",X"A1",X"00",X"C6",X"00",X"E9",X"00",X"0B",X"01",X"2C",X"01",X"4D",X"01",
		X"6D",X"01",X"8C",X"01",X"A8",X"01",X"C4",X"01",X"DD",X"01",X"F8",X"01",X"11",X"02",X"2B",X"02",
		X"40",X"02",X"55",X"02",X"6D",X"02",X"81",X"02",X"94",X"02",X"A8",X"02",X"BA",X"02",X"CB",X"02",
		X"DC",X"02",X"ED",X"02",X"FC",X"02",X"0B",X"03",X"1A",X"03",X"25",X"03",X"34",X"03",X"40",X"03",
		X"4B",X"03",X"57",X"03",X"63",X"03",X"6C",X"03",X"77",X"03",X"81",X"03",X"88",X"03",X"92",X"03",
		X"99",X"03",X"A2",X"03",X"A8",X"03",X"B0",X"03",X"B6",X"03",X"BB",X"03",X"C1",X"03",X"C7",X"03",
		X"C3",X"03",X"B0",X"03",X"93",X"03",X"6E",X"03",X"48",X"03",X"1D",X"03",X"F1",X"02",X"C5",X"02",
		X"9B",X"02",X"71",X"02",X"47",X"02",X"1F",X"02",X"F7",X"01",X"D1",X"01",X"AC",X"01",X"87",X"01",
		X"65",X"01",X"43",X"01",X"23",X"01",X"04",X"01",X"E6",X"00",X"C8",X"00",X"AD",X"00",X"92",X"00",
		X"78",X"00",X"5D",X"00",X"46",X"00",X"31",X"00",X"28",X"00",X"2F",X"00",X"3D",X"00",X"4E",X"00",
		X"66",X"00",X"7D",X"00",X"97",X"00",X"B1",X"00",X"CB",X"00",X"E6",X"00",X"FE",X"00",X"18",X"01",
		X"30",X"01",X"47",X"01",X"5C",X"01",X"73",X"01",X"88",X"01",X"9B",X"01",X"B0",X"01",X"C2",X"01",
		X"D3",X"01",X"E4",X"01",X"F6",X"01",X"06",X"02",X"15",X"02",X"23",X"02",X"32",X"02",X"40",X"02",
		X"4D",X"02",X"5A",X"02",X"64",X"02",X"71",X"02",X"7B",X"02",X"86",X"02",X"90",X"02",X"99",X"02",
		X"A2",X"02",X"AA",X"02",X"B3",X"02",X"BC",X"02",X"C3",X"02",X"CA",X"02",X"D1",X"02",X"D6",X"02",
		X"DD",X"02",X"E2",X"02",X"E8",X"02",X"EE",X"02",X"F2",X"02",X"F6",X"02",X"FB",X"02",X"FF",X"02",
		X"02",X"03",X"04",X"03",X"09",X"03",X"0D",X"03",X"10",X"03",X"11",X"03",X"15",X"03",X"18",X"03",
		X"19",X"03",X"1A",X"03",X"1C",X"03",X"1B",X"03",X"23",X"03",X"26",X"03",X"26",X"03",X"28",X"03",
		X"28",X"03",X"29",X"03",X"29",X"03",X"2A",X"03",X"29",X"03",X"29",X"03",X"27",X"03",X"28",X"03",
		X"28",X"03",X"27",X"03",X"26",X"03",X"25",X"03",X"23",X"03",X"22",X"03",X"17",X"03",X"03",X"03",
		X"E6",X"02",X"C7",X"02",X"A3",X"02",X"7F",X"02",X"5A",X"02",X"36",X"02",X"12",X"02",X"F0",X"01",
		X"CC",X"01",X"AB",X"01",X"89",X"01",X"6A",X"01",X"4C",X"01",X"2E",X"01",X"11",X"01",X"F5",X"00",
		X"DA",X"00",X"C1",X"00",X"A8",X"00",X"90",X"00",X"7A",X"00",X"63",X"00",X"4F",X"00",X"38",X"00",
		X"24",X"00",X"14",X"00",X"0E",X"00",X"13",X"00",X"1C",X"00",X"2A",X"00",X"37",X"00",X"48",X"00",
		X"59",X"00",X"6B",X"00",X"7E",X"00",X"8F",X"00",X"9F",X"00",X"B2",X"00",X"BF",X"00",X"D0",X"00",
		X"DE",X"00",X"EC",X"00",X"FC",X"00",X"09",X"01",X"18",X"01",X"22",X"01",X"2F",X"01",X"3B",X"01",
		X"47",X"01",X"52",X"01",X"5C",X"01",X"64",X"01",X"6E",X"01",X"71",X"01",X"6B",X"01",X"5D",X"01",
		X"4C",X"01",X"36",X"01",X"23",X"01",X"0D",X"01",X"F5",X"00",X"E0",X"00",X"CA",X"00",X"B5",X"00",
		X"A0",X"00",X"8C",X"00",X"77",X"00",X"65",X"00",X"52",X"00",X"42",X"00",X"2F",X"00",X"1F",X"00",
		X"0F",X"00",X"01",X"00",X"F3",X"FF",X"E4",X"FF",X"D7",X"FF",X"CA",X"FF",X"BE",X"FF",X"B2",X"FF",
		X"A6",X"FF",X"9C",X"FF",X"92",X"FF",X"87",X"FF",X"7F",X"FF",X"75",X"FF",X"6C",X"FF",X"64",X"FF",
		X"5C",X"FF",X"56",X"FF",X"4E",X"FF",X"47",X"FF",X"40",X"FF",X"39",X"FF",X"33",X"FF",X"2D",X"FF",
		X"29",X"FF",X"24",X"FF",X"1F",X"FF",X"1A",X"FF",X"15",X"FF",X"11",X"FF",X"0F",X"FF",X"0C",X"FF",
		X"08",X"FF",X"05",X"FF",X"02",X"FF",X"FF",X"FE",X"01",X"FF",X"0A",X"FF",X"1A",X"FF",X"2C",X"FF",
		X"3F",X"FF",X"53",X"FF",X"6B",X"FF",X"80",X"FF",X"96",X"FF",X"AC",X"FF",X"C1",X"FF",X"D4",X"FF",
		X"E8",X"FF",X"FB",X"FF",X"0D",X"00",X"1F",X"00",X"30",X"00",X"41",X"00",X"52",X"00",X"60",X"00",
		X"6F",X"00",X"7E",X"00",X"8D",X"00",X"98",X"00",X"A6",X"00",X"B3",X"00",X"BF",X"00",X"CB",X"00",
		X"D6",X"00",X"E0",X"00",X"E9",X"00",X"F3",X"00",X"FC",X"00",X"05",X"01",X"0F",X"01",X"15",X"01",
		X"1D",X"01",X"26",X"01",X"2D",X"01",X"33",X"01",X"3A",X"01",X"40",X"01",X"47",X"01",X"4C",X"01",
		X"52",X"01",X"56",X"01",X"5C",X"01",X"60",X"01",X"65",X"01",X"6A",X"01",X"6C",X"01",X"70",X"01",
		X"74",X"01",X"77",X"01",X"7C",X"01",X"7B",X"01",X"77",X"01",X"6C",X"01",X"61",X"01",X"52",X"01",
		X"43",X"01",X"34",X"01",X"24",X"01",X"16",X"01",X"07",X"01",X"F9",X"00",X"EA",X"00",X"DD",X"00",
		X"CF",X"00",X"C2",X"00",X"B5",X"00",X"AA",X"00",X"9C",X"00",X"94",X"00",X"88",X"00",X"7C",X"00",
		X"74",X"00",X"6B",X"00",X"61",X"00",X"58",X"00",X"50",X"00",X"47",X"00",X"3F",X"00",X"39",X"00",
		X"33",X"00",X"2B",X"00",X"27",X"00",X"20",X"00",X"19",X"00",X"15",X"00",X"10",X"00",X"0A",X"00",
		X"05",X"00",X"01",X"00",X"FE",X"FF",X"F9",X"FF",X"F5",X"FF",X"F1",X"FF",X"EE",X"FF",X"EC",X"FF",
		X"E8",X"FF",X"E5",X"FF",X"E4",X"FF",X"E1",X"FF",X"E0",X"FF",X"DD",X"FF",X"DB",X"FF",X"D9",X"FF",
		X"D7",X"FF",X"D6",X"FF",X"D5",X"FF",X"DA",X"FF",X"E0",X"FF",X"E9",X"FF",X"F3",X"FF",X"FD",X"FF",
		X"08",X"00",X"13",X"00",X"1C",X"00",X"27",X"00",X"32",X"00",X"3D",X"00",X"47",X"00",X"51",X"00",
		X"5A",X"00",X"63",X"00",X"6B",X"00",X"72",X"00",X"7A",X"00",X"84",X"00",X"89",X"00",X"90",X"00",
		X"97",X"00",X"9E",X"00",X"A5",X"00",X"AA",X"00",X"AF",X"00",X"B4",X"00",X"B9",X"00",X"BF",X"00",
		X"C4",X"00",X"C9",X"00",X"CC",X"00",X"D1",X"00",X"D5",X"00",X"DA",X"00",X"DC",X"00",X"E0",X"00",
		X"E2",X"00",X"E6",X"00",X"E8",X"00",X"EC",X"00",X"EC",X"00",X"EF",X"00",X"F0",X"00",X"F3",X"00",
		X"F4",X"00",X"F6",X"00",X"F9",X"00",X"FA",X"00",X"FC",X"00",X"FD",X"00",X"FE",X"00",X"00",X"01",
		X"00",X"01",X"00",X"01",X"FF",X"00",X"FB",X"00",X"F6",X"00",X"F2",X"00",X"ED",X"00",X"E7",X"00",
		X"E2",X"00",X"DC",X"00",X"D7",X"00",X"D1",X"00",X"CD",X"00",X"C8",X"00",X"C4",X"00",X"BE",X"00",
		X"BC",X"00",X"B6",X"00",X"B2",X"00",X"B0",X"00",X"AC",X"00",X"A9",X"00",X"A7",X"00",X"A2",X"00",
		X"A0",X"00",X"9D",X"00",X"9B",X"00",X"98",X"00",X"97",X"00",X"95",X"00",X"93",X"00",X"91",X"00",
		X"91",X"00",X"8D",X"00",X"8D",X"00",X"8A",X"00",X"8B",X"00",X"8A",X"00",X"88",X"00",X"88",X"00",
		X"87",X"00",X"86",X"00",X"86",X"00",X"85",X"00",X"86",X"00",X"85",X"00",X"85",X"00",X"86",X"00",
		X"85",X"00",X"85",X"00",X"85",X"00",X"84",X"00",X"85",X"00",X"86",X"00",X"86",X"00",X"86",X"00",
		X"86",X"00",X"87",X"00",X"87",X"00",X"88",X"00",X"8A",X"00",X"8B",X"00",X"8B",X"00",X"8B",X"00",
		X"8D",X"00",X"8E",X"00",X"8F",X"00",X"90",X"00",X"90",X"00",X"91",X"00",X"93",X"00",X"95",X"00",
		X"95",X"00",X"96",X"00",X"98",X"00",X"99",X"00",X"9A",X"00",X"9C",X"00",X"9E",X"00",X"9E",X"00",
		X"A0",X"00",X"A0",X"00",X"A2",X"00",X"A3",X"00",X"A6",X"00",X"A8",X"00",X"A9",X"00",X"AB",X"00",
		X"AC",X"00",X"AF",X"00",X"AF",X"00",X"B1",X"00",X"B2",X"00",X"B3",X"00",X"B5",X"00",X"B7",X"00",
		X"BA",X"00",X"BC",X"00",X"BE",X"00",X"BF",X"00",X"C0",X"00",X"C2",X"00",X"C4",X"00",X"C5",X"00",
		X"C7",X"00",X"C9",X"00",X"CA",X"00",X"CD",X"00",X"CE",X"00",X"D1",X"00",X"D2",X"00",X"D2",X"00",
		X"D5",X"00",X"D7",X"00",X"D7",X"00",X"DC",X"00",X"DB",X"00",X"DD",X"00",X"E0",X"00",X"E2",X"00",
		X"E5",X"00",X"E5",X"00",X"E6",X"00",X"EA",X"00",X"EB",X"00",X"EC",X"00",X"EF",X"00",X"F2",X"00",
		X"F3",X"00",X"F4",X"00",X"F4",X"00",X"F8",X"00",X"FA",X"00",X"FB",X"00",X"FE",X"00",X"FF",X"00",
		X"01",X"01",X"04",X"01",X"04",X"01",X"06",X"01",X"08",X"01",X"09",X"01",X"0C",X"01",X"0E",X"01",
		X"0F",X"01",X"12",X"01",X"12",X"01",X"16",X"01",X"16",X"01",X"1B",X"01",X"1D",X"01",X"1E",X"01",
		X"1F",X"01",X"22",X"01",X"24",X"01",X"26",X"01",X"28",X"01",X"2A",X"01",X"2B",X"01",X"2D",X"01",
		X"2D",X"01",X"31",X"01",X"32",X"01",X"34",X"01",X"35",X"01",X"38",X"01",X"38",X"01",X"3B",X"01",
		X"3D",X"01",X"3F",X"01",X"40",X"01",X"42",X"01",X"44",X"01",X"45",X"01",X"46",X"01",X"49",X"01",
		X"48",X"01",X"4A",X"01",X"4D",X"01",X"4F",X"01",X"4F",X"01",X"52",X"01",X"53",X"01",X"57",X"01",
		X"56",X"01",X"59",X"01",X"58",X"01",X"5D",X"01",X"5C",X"01",X"60",X"01",X"5F",X"01",X"62",X"01",
		X"63",X"01",X"67",X"01",X"65",X"01",X"69",X"01",X"6A",X"01",X"6C",X"01",X"6C",X"01",X"70",X"01",
		X"70",X"01",X"72",X"01",X"72",X"01",X"75",X"01",X"75",X"01",X"78",X"01",X"7A",X"01",X"7B",X"01",
		X"7D",X"01",X"7F",X"01",X"80",X"01",X"81",X"01",X"83",X"01",X"85",X"01",X"87",X"01",X"87",X"01",
		X"8B",X"01",X"88",X"01",X"8B",X"01",X"88",X"01",X"90",X"01",X"8E",X"01",X"98",X"01",X"94",X"01",
		X"9E",X"01",X"8D",X"01",X"98",X"01",X"76",X"01",X"98",X"01",X"B0",X"B0",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"01",X"00",X"FE",X"FF",X"00",X"00",
		X"FE",X"FF",X"00",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"FE",X"FF",X"01",X"00",X"FE",X"FF",X"00",X"00",X"FE",X"FF",X"02",X"00",X"FD",X"FF",
		X"04",X"00",X"FD",X"FF",X"05",X"00",X"FC",X"FF",X"05",X"00",X"FB",X"FF",X"06",X"00",X"FA",X"FF",
		X"08",X"00",X"F9",X"FF",X"08",X"00",X"F8",X"FF",X"09",X"00",X"F6",X"FF",X"0B",X"00",X"F4",X"FF",
		X"0C",X"00",X"F3",X"FF",X"0D",X"00",X"F1",X"FF",X"0E",X"00",X"F1",X"FF",X"0F",X"00",X"F0",X"FF",
		X"11",X"00",X"EE",X"FF",X"12",X"00",X"ED",X"FF",X"15",X"00",X"EC",X"FF",X"15",X"00",X"EA",X"FF",
		X"17",X"00",X"E8",X"FF",X"18",X"00",X"E7",X"FF",X"1A",X"00",X"E5",X"FF",X"1A",X"00",X"E4",X"FF",
		X"1D",X"00",X"E4",X"FF",X"1D",X"00",X"E2",X"FF",X"1E",X"00",X"E2",X"FF",X"1F",X"00",X"E0",X"FF",
		X"22",X"00",X"DF",X"FF",X"21",X"00",X"DE",X"FF",X"24",X"00",X"DC",X"FF",X"25",X"00",X"D9",X"FF",
		X"29",X"00",X"D2",X"FF",X"39",X"00",X"A5",X"FF",X"3A",X"01",X"EA",X"14",X"1E",X"12",X"46",X"0C",
		X"F0",X"07",X"19",X"02",X"8C",X"01",X"C3",X"0B",X"35",X"16",X"F7",X"20",X"F8",X"21",X"DE",X"1B",
		X"7E",X"17",X"F1",X"11",X"62",X"0D",X"08",X"08",X"46",X"03",X"E9",X"FF",X"17",X"09",X"15",X"13",
		X"6E",X"1E",X"85",X"22",X"38",X"1D",X"8C",X"18",X"6E",X"13",X"B0",X"0E",X"9E",X"09",X"04",X"05",
		X"D4",X"FF",X"66",X"03",X"65",X"0E",X"2A",X"18",X"E8",X"21",X"C6",X"1F",X"AC",X"1A",X"DB",X"15",
		X"09",X"11",X"2F",X"0C",X"6E",X"07",X"7A",X"02",X"08",X"FF",X"EF",X"06",X"53",X"11",X"C9",X"1B",
		X"1C",X"22",X"2F",X"1D",X"A7",X"18",X"65",X"13",X"DD",X"0E",X"95",X"09",X"31",X"05",X"8E",X"FF",
		X"DE",X"00",X"C8",X"0B",X"AD",X"15",X"20",X"20",X"BE",X"1F",X"19",X"1A",X"79",X"15",X"49",X"10",
		X"7E",X"0B",X"72",X"06",X"70",X"01",X"44",X"FE",X"40",X"07",X"89",X"11",X"A0",X"1C",X"D5",X"20",
		X"51",X"1B",X"D0",X"16",X"77",X"11",X"E6",X"0C",X"99",X"07",X"27",X"03",X"D4",X"FD",X"59",X"02",
		X"32",X"0D",X"50",X"17",X"6B",X"20",X"A3",X"1D",X"85",X"18",X"B7",X"13",X"D6",X"0E",X"FD",X"09",
		X"3A",X"05",X"34",X"00",X"81",X"FD",X"5F",X"06",X"59",X"10",X"FD",X"1A",X"41",X"20",X"3E",X"1B",
		X"BD",X"16",X"A5",X"11",X"1F",X"0D",X"07",X"08",X"A0",X"03",X"31",X"FE",X"8D",X"FE",X"20",X"09",
		X"B2",X"12",X"AB",X"1D",X"E1",X"1E",X"1C",X"19",X"BE",X"14",X"74",X"0F",X"ED",X"0A",X"B1",X"05",
		X"30",X"01",X"55",X"FC",X"8D",X"02",X"39",X"0D",X"C4",X"17",X"A7",X"1F",X"52",X"1B",X"82",X"16",
		X"57",X"11",X"9E",X"0C",X"65",X"07",X"D8",X"02",X"3B",X"FD",X"2B",X"FE",X"3C",X"09",X"21",X"13",
		X"DD",X"1D",X"21",X"1D",X"76",X"17",X"BD",X"12",X"92",X"0D",X"A8",X"08",X"AD",X"03",X"78",X"FE",
		X"23",X"FC",X"EF",X"05",X"24",X"10",X"68",X"1B",X"E9",X"1D",X"23",X"18",X"8C",X"13",X"28",X"0E",
		X"6A",X"09",X"22",X"04",X"4E",X"FF",X"11",X"FB",X"6A",X"03",X"1E",X"0E",X"36",X"19",X"25",X"1E",
		X"93",X"18",X"FF",X"13",X"8C",X"0E",X"E9",X"09",X"88",X"04",X"F9",X"FF",X"DB",X"FA",X"C4",X"00",
		X"97",X"0B",X"33",X"16",X"33",X"1E",X"D2",X"19",X"05",X"15",X"E3",X"0F",X"31",X"0B",X"0A",X"06",
		X"85",X"01",X"0B",X"FC",X"33",X"FC",X"C5",X"06",X"6D",X"10",X"65",X"1B",X"96",X"1C",X"DE",X"16",
		X"87",X"12",X"49",X"0D",X"D4",X"08",X"AA",X"03",X"4A",X"FF",X"2C",X"FA",X"20",X"FF",X"C9",X"09",
		X"AD",X"13",X"BE",X"1C",X"81",X"1A",X"52",X"15",X"BC",X"10",X"D0",X"0B",X"33",X"07",X"55",X"02",
		X"B4",X"FD",X"BB",X"F9",X"E7",X"00",X"1D",X"0B",X"47",X"15",X"DE",X"1C",X"38",X"19",X"6A",X"14",
		X"AB",X"0F",X"F8",X"0A",X"40",X"06",X"96",X"01",X"CE",X"FC",X"7C",X"F9",X"64",X"01",X"67",X"0B",
		X"AB",X"15",X"9C",X"1C",X"76",X"18",X"CC",X"13",X"E7",X"0E",X"44",X"0A",X"5D",X"05",X"CA",X"00",
		X"AD",X"FB",X"7C",X"F9",X"05",X"03",X"DD",X"0C",X"C4",X"17",X"3D",X"1C",X"92",X"16",X"43",X"12",
		X"EE",X"0C",X"7F",X"08",X"31",X"03",X"DD",X"FE",X"4D",X"F9",X"46",X"FC",X"41",X"07",X"2C",X"11",
		X"6A",X"1B",X"73",X"19",X"FA",X"13",X"4C",X"0F",X"3B",X"0A",X"6F",X"05",X"84",X"00",X"88",X"FB",
		X"B5",X"F8",X"E7",X"01",X"DA",X"0B",X"EA",X"16",X"A5",X"1B",X"0D",X"16",X"B8",X"11",X"71",X"0C",
		X"03",X"08",X"CA",X"02",X"81",X"FE",X"F9",X"F8",X"D8",X"FA",X"79",X"05",X"1E",X"0F",X"71",X"19",
		X"D6",X"19",X"53",X"14",X"FB",X"0F",X"D7",X"0A",X"70",X"06",X"52",X"01",X"09",X"FD",X"E3",X"F7",
		X"7B",X"FC",X"22",X"07",X"D3",X"10",X"5A",X"1A",X"9C",X"18",X"5E",X"13",X"ED",X"0E",X"F2",X"09",
		X"7D",X"05",X"84",X"00",X"2C",X"FC",X"62",X"F7",X"0F",X"FD",X"94",X"07",X"49",X"11",X"58",X"1A",
		X"F8",X"17",X"E6",X"12",X"66",X"0E",X"8A",X"09",X"0B",X"05",X"2C",X"00",X"C4",X"FB",X"29",X"F7",
		X"D7",X"FC",X"47",X"07",X"F5",X"10",X"F0",X"19",X"AD",X"17",X"98",X"12",X"0C",X"0E",X"2A",X"09",
		X"95",X"04",X"B1",X"FF",X"20",X"FB",X"CC",X"F6",X"AA",X"FD",X"1F",X"08",X"5E",X"12",X"5A",X"1A",
		X"2D",X"16",X"70",X"11",X"6E",X"0C",X"C3",X"07",X"BA",X"02",X"29",X"FE",X"D3",X"F8",X"AB",X"F7",
		X"B2",X"01",X"91",X"0B",X"99",X"16",X"1E",X"19",X"72",X"13",X"05",X"0F",X"B3",X"09",X"23",X"05",
		X"DF",X"FF",X"57",X"FB",X"62",X"F6",X"78",X"FC",X"45",X"07",X"E5",X"11",X"D7",X"19",X"41",X"15",
		X"81",X"10",X"3B",X"0B",X"90",X"06",X"3D",X"01",X"C5",X"FC",X"09",X"F7",X"E8",X"F8",X"31",X"04",
		X"49",X"0E",X"71",X"18",X"BC",X"16",X"4B",X"11",X"66",X"0C",X"5A",X"07",X"4B",X"02",X"75",X"FD",
		X"08",X"F8",X"1B",X"F7",X"B3",X"01",X"A7",X"0B",X"08",X"17",X"E7",X"17",X"F8",X"11",X"82",X"0D",
		X"2F",X"08",X"8C",X"03",X"60",X"FE",X"AF",X"F9",X"77",X"F5",X"6B",X"FD",X"E3",X"07",X"98",X"12",
		X"00",X"19",X"FB",X"13",X"6C",X"0F",X"40",X"0A",X"B4",X"05",X"8B",X"00",X"29",X"FC",X"AA",X"F6",
		X"65",X"F7",X"0E",X"02",X"9B",X"0B",X"77",X"16",X"87",X"17",X"DB",X"11",X"90",X"0D",X"60",X"08",
		X"F7",X"03",X"D7",X"FE",X"88",X"FA",X"5C",X"F5",X"8A",X"F9",X"41",X"04",X"E7",X"0D",X"90",X"17",
		X"20",X"16",X"C6",X"10",X"5B",X"0C",X"5D",X"07",X"E4",X"02",X"F0",X"FD",X"87",X"F9",X"E1",X"F4",
		X"9D",X"FA",X"12",X"05",X"D5",X"0E",X"B2",X"17",X"5B",X"15",X"3C",X"10",X"BF",X"0B",X"E2",X"06",
		X"59",X"02",X"81",X"FD",X"FA",X"F8",X"A0",X"F4",X"07",X"FB",X"74",X"05",X"7A",X"0F",X"B5",X"17",
		X"7C",X"14",X"84",X"0F",X"C2",X"0A",X"F3",X"05",X"23",X"01",X"67",X"FC",X"66",X"F7",X"C0",X"F4",
		X"07",X"FE",X"F8",X"07",X"08",X"13",X"BF",X"17",X"0A",X"12",X"B4",X"0D",X"59",X"08",X"E2",X"03",
		X"93",X"FE",X"36",X"FA",X"AC",X"F4",X"25",X"F8",X"42",X"03",X"48",X"0D",X"29",X"17",X"93",X"14",
		X"45",X"0F",X"69",X"0A",X"72",X"05",X"70",X"00",X"AA",X"FB",X"4F",X"F6",X"08",X"F5",X"6F",X"FF",
		X"87",X"09",X"90",X"14",X"1D",X"16",X"5F",X"10",X"CA",X"0B",X"7B",X"06",X"BB",X"01",X"8D",X"FC",
		X"AB",X"F7",X"EC",X"F3",X"8E",X"FC",X"F7",X"06",X"58",X"12",X"0B",X"17",X"1F",X"11",X"A9",X"0C",
		X"2A",X"07",X"8A",X"02",X"24",X"FD",X"81",X"F8",X"9B",X"F3",X"70",X"FA",X"51",X"05",X"63",X"10",
		X"ED",X"16",X"C1",X"11",X"17",X"0D",X"A4",X"07",X"F9",X"02",X"86",X"FD",X"F5",X"F8",X"90",X"F3",
		X"F7",X"F8",X"31",X"04",X"FF",X"0E",X"AE",X"16",X"1E",X"12",X"4D",X"0D",X"E3",X"07",X"2D",X"03",
		X"B7",X"FD",X"2B",X"F9",X"87",X"F3",X"02",X"F8",X"6D",X"03",X"13",X"0E",X"6F",X"16",X"44",X"12",
		X"5B",X"0D",X"F8",X"07",X"3A",X"03",X"C0",X"FD",X"36",X"F9",X"76",X"F3",X"69",X"F7",X"E8",X"02",
		X"84",X"0D",X"34",X"16",X"46",X"12",X"4B",X"0D",X"EF",X"07",X"27",X"03",X"B0",X"FD",X"21",X"F9",
		X"5D",X"F3",X"18",X"F7",X"99",X"02",X"36",X"0D",X"03",X"16",X"28",X"12",X"2B",X"0D",X"D4",X"07",
		X"0F",X"03",X"A4",X"FD",X"21",X"F9",X"59",X"F3",X"45",X"F6",X"B5",X"01",X"E5",X"0B",X"86",X"15",
		X"E4",X"12",X"AF",X"0D",X"B6",X"08",X"D5",X"03",X"C5",X"FE",X"1B",X"FA",X"B1",X"F4",X"B9",X"F3",
		X"F8",X"FD",X"E0",X"07",X"D1",X"12",X"F3",X"14",X"5B",X"0F",X"F1",X"0A",X"B4",X"05",X"34",X"01",
		X"0A",X"FC",X"A1",X"F7",X"88",X"F2",X"77",X"F7",X"40",X"02",X"35",X"0C",X"3D",X"15",X"BB",X"12",
		X"92",X"0D",X"F0",X"08",X"0C",X"04",X"61",X"FF",X"91",X"FA",X"D2",X"F5",X"50",X"F2",X"46",X"FA",
		X"5B",X"04",X"CC",X"0E",X"88",X"15",X"3F",X"11",X"9E",X"0C",X"BE",X"07",X"25",X"03",X"51",X"FE",
		X"C8",X"F9",X"CA",X"F4",X"6D",X"F2",X"87",X"FB",X"43",X"05",X"DF",X"0F",X"68",X"15",X"72",X"10",
		X"0C",X"0C",X"FD",X"06",X"85",X"02",X"7C",X"FD",X"18",X"F9",X"C0",X"F3",X"33",X"F3",X"66",X"FD",
		X"1E",X"07",X"F4",X"11",X"92",X"14",X"DA",X"0E",X"8E",X"0A",X"40",X"05",X"D3",X"00",X"8B",X"FB",
		X"34",X"F7",X"DA",X"F1",X"AF",X"F6",X"B5",X"01",X"D9",X"0B",X"F5",X"14",X"A2",X"11",X"8E",X"0C",
		X"9B",X"07",X"C2",X"02",X"B5",X"FD",X"09",X"F9",X"9D",X"F3",X"E4",X"F2",X"83",X"FD",X"83",X"07",
		X"77",X"12",X"99",X"13",X"E2",X"0D",X"4C",X"09",X"07",X"04",X"4B",X"FF",X"26",X"FA",X"41",X"F5",
		X"98",X"F1",X"42",X"FA",X"A6",X"04",X"FF",X"0F",X"A3",X"14",X"DC",X"0E",X"64",X"0A",X"EC",X"04",
		X"51",X"00",X"EB",X"FA",X"54",X"F6",X"54",X"F1",X"C8",X"F7",X"C3",X"02",X"8E",X"0D",X"95",X"14",
		X"E6",X"0F",X"30",X"0B",X"EA",X"05",X"48",X"01",X"FF",X"FB",X"8D",X"F7",X"F9",X"F1",X"77",X"F4",
		X"74",X"FF",X"66",X"09",X"99",X"13",X"28",X"12",X"C6",X"0C",X"22",X"08",X"1F",X"03",X"67",X"FE",
		X"82",X"F9",X"AB",X"F4",X"2F",X"F1",X"57",X"F9",X"87",X"03",X"26",X"0E",X"4E",X"14",X"A5",X"0F",
		X"11",X"0B",X"00",X"06",X"71",X"01",X"5C",X"FC",X"EC",X"F7",X"7D",X"F2",X"A8",X"F2",X"43",X"FD",
		X"06",X"07",X"D2",X"11",X"10",X"13",X"5D",X"0D",X"EF",X"08",X"AE",X"03",X"1C",X"FF",X"EF",X"F9",
		X"55",X"F5",X"C4",X"F0",X"B9",X"F7",X"79",X"02",X"1F",X"0D",X"17",X"14",X"73",X"0F",X"BA",X"0A",
		X"7E",X"05",X"D7",X"00",X"8E",X"FB",X"16",X"F7",X"74",X"F1",X"EE",X"F3",X"04",X"FF",X"08",X"09",
		X"22",X"13",X"79",X"11",X"27",X"0C",X"67",X"07",X"6F",X"02",X"9C",X"FD",X"CA",X"F8",X"C9",X"F3",
		X"DD",X"F0",X"AC",X"F9",X"C7",X"03",X"95",X"0E",X"B8",X"13",X"A0",X"0E",X"2D",X"0A",X"05",X"05",
		X"8E",X"00",X"6D",X"FB",X"1A",X"F7",X"A9",X"F1",X"8A",X"F2",X"2D",X"FD",X"AD",X"06",X"6B",X"11",
		X"CD",X"12",X"17",X"0D",X"E4",X"08",X"B3",X"03",X"62",X"FF",X"3F",X"FA",X"09",X"F6",X"B3",X"F0",
		X"1A",X"F4",X"BE",X"FE",X"4B",X"08",X"42",X"12",X"E1",X"11",X"70",X"0C",X"25",X"08",X"1B",X"03",
		X"BF",X"FE",X"BC",X"F9",X"7A",X"F5",X"68",X"F0",X"A3",X"F4",X"35",X"FF",X"B7",X"08",X"6E",X"12",
		X"92",X"11",X"35",X"0C",X"EA",X"07",X"EE",X"02",X"93",X"FE",X"99",X"F9",X"58",X"F5",X"4F",X"F0",
		X"76",X"F4",X"0E",X"FF",X"7F",X"08",X"61",X"12",X"8A",X"11",X"1E",X"0C",X"DD",X"07",X"D9",X"02",
		X"83",X"FE",X"85",X"F9",X"4B",X"F5",X"39",X"F0",X"38",X"F4",X"DF",X"FE",X"42",X"08",X"66",X"12",
		X"83",X"11",X"06",X"0C",X"D3",X"07",X"C2",X"02",X"7A",X"FE",X"6C",X"F9",X"45",X"F5",X"10",X"F0",
		X"FC",X"F3",X"AC",X"FE",X"14",X"08",X"1E",X"12",X"62",X"11",X"FE",X"0B",X"BE",X"07",X"B7",X"02",
		X"68",X"FE",X"60",X"F9",X"33",X"F5",X"01",X"F0",X"D4",X"F3",X"77",X"FE",X"E6",X"07",X"D7",X"11",
		X"48",X"11",X"F5",X"0B",X"AA",X"07",X"AB",X"02",X"54",X"FE",X"54",X"F9",X"1D",X"F5",X"FD",X"EF",
		X"B1",X"F3",X"43",X"FE",X"B6",X"07",X"9B",X"11",X"3A",X"11",X"E6",X"0B",X"9A",X"07",X"9D",X"02",
		X"3E",X"FE",X"3C",X"F9",X"F7",X"F4",X"D9",X"EF",X"F1",X"F3",X"9D",X"FE",X"56",X"08",X"03",X"12",
		X"87",X"10",X"40",X"0B",X"B5",X"06",X"B8",X"01",X"16",X"FD",X"25",X"F8",X"74",X"F3",X"7E",X"EF",
		X"1A",X"F7",X"90",X"01",X"23",X"0C",X"CF",X"12",X"22",X"0E",X"7A",X"09",X"56",X"04",X"B8",X"FF",
		X"89",X"FA",X"11",X"F6",X"84",X"F0",X"EA",X"F1",X"EE",X"FC",X"DF",X"06",X"51",X"11",X"A4",X"10",
		X"21",X"0B",X"6C",X"06",X"53",X"01",X"77",X"FC",X"88",X"F7",X"6A",X"F2",X"BB",X"EF",X"39",X"F9",
		X"6E",X"03",X"C3",X"0E",X"1F",X"12",X"51",X"0C",X"DC",X"07",X"6E",X"02",X"D5",X"FD",X"7B",X"F8",
		X"DE",X"F3",X"17",X"EF",X"5F",X"F6",X"48",X"01",X"36",X"0C",X"76",X"12",X"5A",X"0D",X"AD",X"08",
		X"4C",X"03",X"A0",X"FE",X"3E",X"F9",X"AD",X"F4",X"4F",X"EF",X"91",X"F4",X"C2",X"FF",X"71",X"0A",
		X"91",X"12",X"0C",X"0E",X"30",X"09",X"DB",X"03",X"20",X"FF",X"B9",X"F9",X"2D",X"F5",X"87",X"EF",
		X"68",X"F3",X"B7",X"FE",X"48",X"09",X"81",X"12",X"87",X"0E",X"7E",X"09",X"4B",X"04",X"7D",X"FF",
		X"34",X"FA",X"A3",X"F5",X"FB",X"EF",X"E6",X"F1",X"06",X"FD",X"1D",X"07",X"56",X"11",X"D7",X"0F",
		X"7A",X"0A",X"B3",X"05",X"B7",X"00",X"DA",X"FB",X"06",X"F7",X"F4",X"F1",X"56",X"EF",X"80",X"F8",
		X"90",X"02",X"87",X"0D",X"00",X"12",X"A4",X"0C",X"42",X"08",X"09",X"03",X"99",X"FE",X"68",X"F9",
		X"1C",X"F5",X"A3",X"EF",X"C6",X"F1",X"85",X"FC",X"2A",X"06",X"79",X"10",X"94",X"10",X"0B",X"0B",
		X"B6",X"06",X"9B",X"01",X"31",X"FD",X"21",X"F8",X"CD",X"F3",X"DD",X"EE",X"E6",X"F3",X"78",X"FE",
		X"49",X"08",X"73",X"11",X"75",X"0F",X"4F",X"0A",X"D2",X"05",X"ED",X"00",X"6C",X"FC",X"8A",X"F7",
		X"17",X"F3",X"A8",X"EE",X"D5",X"F4",X"3D",X"FF",X"28",X"09",X"B8",X"11",X"E0",X"0E",X"E6",X"09",
		X"3F",X"05",X"6D",X"00",X"C0",X"FB",X"F4",X"F6",X"33",X"F2",X"9C",X"EE",X"CE",X"F6",X"10",X"01",
		X"AE",X"0B",X"29",X"12",X"24",X"0D",X"A1",X"08",X"79",X"03",X"EF",X"FE",X"C1",X"F9",X"59",X"F5",
		X"CF",X"EF",X"C5",X"F0",X"AC",X"FB",X"6A",X"05",X"69",X"10",X"4C",X"10",X"85",X"0A",X"0C",X"06",
		X"CE",X"00",X"25",X"FC",X"08",X"F7",X"3B",X"F2",X"6F",X"EE",X"23",X"F7",X"99",X"01",X"9E",X"0C",
		X"A6",X"11",X"2C",X"0C",X"A6",X"07",X"46",X"02",X"AF",X"FD",X"57",X"F8",X"D2",X"F3",X"84",X"EE",
		X"F3",X"F3",X"FF",X"FE",X"AB",X"09",X"CF",X"11",X"78",X"0D",X"A8",X"08",X"5E",X"03",X"AA",X"FE",
		X"4E",X"F9",X"CB",X"F4",X"18",X"EF",X"B9",X"F1",X"17",X"FD",X"44",X"07",X"0C",X"11",X"BC",X"0E",
		X"7E",X"09",X"91",X"04",X"AC",X"FF",X"A7",X"FA",X"F7",X"F5",X"9C",X"F0",X"44",X"EF",X"5D",X"F9",
		X"4A",X"03",X"4B",X"0E",X"DE",X"10",X"4E",X"0B",X"E8",X"06",X"AE",X"01",X"34",X"FD",X"07",X"F8",
		X"A7",X"F3",X"76",X"EE",X"EF",X"F2",X"C4",X"FD",X"AA",X"07",X"F9",X"10",X"D0",X"0E",X"9A",X"09",
		X"F6",X"04",X"07",X"00",X"50",X"FB",X"75",X"F6",X"99",X"F1",X"3C",X"EE",X"00",X"F7",X"39",X"01",
		X"18",X"0C",X"98",X"11",X"2B",X"0C",X"C0",X"07",X"71",X"02",X"F4",X"FD",X"A3",X"F8",X"49",X"F4",
		X"A5",X"EE",X"B3",X"F1",X"FA",X"FC",X"FC",X"06",X"DA",X"10",X"A5",X"0E",X"56",X"09",X"78",X"04",
		X"85",X"FF",X"86",X"FA",X"C7",X"F5",X"73",X"F0",X"0C",X"EF",X"2A",X"F9",X"2D",X"03",X"2A",X"0E",
		X"92",X"10",X"F6",X"0A",X"88",X"06",X"4C",X"01",X"C7",X"FC",X"9A",X"F7",X"2B",X"F3",X"20",X"EE",
		X"5C",X"F3",X"27",X"FE",X"3C",X"08",X"02",X"11",X"29",X"0E",X"17",X"09",X"60",X"04",X"8C",X"FF",
		X"CE",X"FA",X"0F",X"F6",X"32",X"F1",X"26",X"EE",X"D3",X"F6",X"D1",X"00",X"89",X"0B",X"70",X"11",
		X"5A",X"0C",X"F1",X"07",X"C7",X"02",X"4F",X"FE",X"26",X"F9",X"CC",X"F4",X"42",X"EF",X"FE",X"EF",
		X"A1",X"FA",X"73",X"04",X"25",X"0F",X"D3",X"0F",X"3A",X"0A",X"BE",X"05",X"89",X"00",X"EC",X"FB",
		X"CC",X"F6",X"1C",X"F2",X"DC",X"ED",X"75",X"F5",X"FD",X"FF",X"E9",X"0A",X"3A",X"11",X"36",X"0C",
		X"A0",X"07",X"5A",X"02",X"C4",X"FD",X"80",X"F8",X"16",X"F4",X"8C",X"EE",X"34",X"F1",X"3B",X"FC",
		X"1A",X"06",X"6B",X"10",X"DB",X"0E",X"72",X"09",X"D9",X"04",X"D5",X"FF",X"27",X"FB",X"3F",X"F6",
		X"78",X"F1",X"E5",X"ED",X"E8",X"F5",X"1A",X"00",X"B4",X"0A",X"15",X"11",X"8E",X"0C",X"F7",X"07",
		X"FC",X"02",X"6B",X"FE",X"78",X"F9",X"01",X"F5",X"CC",X"EF",X"AA",X"EE",X"BF",X"F8",X"41",X"02",
		X"3C",X"0D",X"F2",X"10",X"50",X"0B",X"22",X"07",X"FD",X"01",X"A7",X"FD",X"96",X"F8",X"5A",X"F4",
		X"02",X"EF",X"92",X"EF",X"F2",X"F9",X"4C",X"03",X"13",X"0E",X"86",X"10",X"DF",X"0A",X"BF",X"06",
		X"A0",X"01",X"59",X"FD",X"4D",X"F8",X"1F",X"F4",X"CD",X"EE",X"B2",X"EF",X"22",X"FA",X"65",X"03",
		X"30",X"0E",X"76",X"10",X"CF",X"0A",X"B8",X"06",X"96",X"01",X"5A",X"FD",X"46",X"F8",X"27",X"F4",
		X"BF",X"EE",X"83",X"EF",X"00",X"FA",X"4A",X"03",X"FA",X"0D",X"53",X"10",X"DB",X"0A",X"B2",X"06",
		X"9C",X"01",X"57",X"FD",X"4C",X"F8",X"22",X"F4",X"C7",X"EE",X"84",X"EF",X"D7",X"F9",X"31",X"03",
		X"C6",X"0D",X"41",X"10",X"E2",X"0A",X"AE",X"06",X"A1",X"01",X"54",X"FD",X"4E",X"F8",X"20",X"F4",
		X"C6",X"EE",X"8E",X"EF",X"E0",X"F9",X"5F",X"03",X"01",X"0E",X"06",X"10",X"86",X"0A",X"40",X"06",
		X"12",X"01",X"B1",X"FC",X"85",X"F7",X"3F",X"F3",X"DD",X"ED",X"73",X"F1",X"73",X"FC",X"43",X"06",
		X"23",X"10",X"58",X"0E",X"F6",X"08",X"55",X"04",X"51",X"FF",X"92",X"FA",X"A9",X"F5",X"C4",X"F0",
		X"95",X"ED",X"9F",X"F6",X"BB",X"00",X"AC",X"0B",X"DA",X"10",X"69",X"0B",X"09",X"07",X"D2",X"01",
		X"61",X"FD",X"35",X"F8",X"E8",X"F3",X"6F",X"EE",X"03",X"F0",X"AC",X"FA",X"4C",X"04",X"D3",X"0E",
		X"5E",X"0F",X"E0",X"09",X"8A",X"05",X"70",X"00",X"08",X"FC",X"F5",X"F6",X"AC",X"F2",X"89",X"ED",
		X"EC",X"F1",X"C6",X"FC",X"5B",X"06",X"50",X"10",X"57",X"0E",X"08",X"09",X"87",X"04",X"91",X"FF",
		X"F7",X"FA",X"0C",X"F6",X"62",X"F1",X"5A",X"ED",X"C9",X"F4",X"33",X"FF",X"BC",X"09",X"A6",X"10",
		X"42",X"0C",X"91",X"07",X"7E",X"02",X"DD",X"FD",X"BB",X"F8",X"42",X"F4",X"BD",X"EE",X"63",X"EF",
		X"2A",X"FA",X"12",X"04",X"C7",X"0E",X"01",X"0F",X"71",X"09",X"D8",X"04",X"B4",X"FF",X"FC",X"FA",
		X"F7",X"F5",X"25",X"F1",X"5F",X"ED",X"6D",X"F5",X"CD",X"FF",X"97",X"0A",X"99",X"10",X"AF",X"0B",
		X"2B",X"07",X"FF",X"01",X"7F",X"FD",X"57",X"F8",X"FF",X"F3",X"81",X"EE",X"71",X"EF",X"05",X"FA",
		X"B2",X"03",X"44",X"0E",X"74",X"0F",X"DA",X"09",X"91",X"05",X"68",X"00",X"08",X"FC",X"E8",X"F6",
		X"A6",X"F2",X"76",X"ED",X"B5",X"F1",X"5F",X"FC",X"1A",X"06",X"B4",X"0F",X"4C",X"0E",X"07",X"09",
		X"9F",X"04",X"A5",X"FF",X"35",X"FB",X"3F",X"F6",X"E6",X"F1",X"27",X"ED",X"DB",X"F2",X"60",X"FD",
		X"27",X"07",X"25",X"10",X"C5",X"0D",X"BA",X"08",X"3B",X"04",X"65",X"FF",X"E7",X"FA",X"12",X"F6",
		X"A7",X"F1",X"29",X"ED",X"11",X"F3",X"7D",X"FD",X"3C",X"07",X"15",X"10",X"B3",X"0D",X"AC",X"08",
		X"21",X"04",X"4C",X"FF",X"BA",X"FA",X"E0",X"F5",X"4E",X"F1",X"17",X"ED",X"11",X"F4",X"82",X"FE",
		X"CC",X"08",X"AA",X"10",X"85",X"0C",X"D0",X"07",X"D4",X"02",X"31",X"FE",X"2C",X"F9",X"A6",X"F4",
		X"51",X"EF",X"34",X"EE",X"3F",X"F8",X"25",X"02",X"26",X"0D",X"B7",X"0F",X"18",X"0A",X"AD",X"05",
		X"64",X"00",X"DB",X"FB",X"9D",X"F6",X"19",X"F2",X"26",X"ED",X"31",X"F3",X"07",X"FE",X"A8",X"08",
		X"97",X"10",X"2A",X"0C",X"6A",X"07",X"2F",X"02",X"87",X"FD",X"3B",X"F8",X"C5",X"F3",X"0B",X"EE",
		X"D3",X"EF",X"28",X"FB",X"38",X"05",X"80",X"0F",X"E3",X"0D",X"70",X"08",X"93",X"03",X"8C",X"FE",
		X"83",X"F9",X"B2",X"F4",X"46",X"EF",X"4B",X"EE",X"E3",X"F8",X"E6",X"02",X"41",X"0E",X"28",X"0F",
		X"4D",X"09",X"CF",X"04",X"87",X"FF",X"E2",X"FA",X"BD",X"F5",X"05",X"F1",X"F4",X"EC",X"18",X"F5",
		X"8E",X"FF",X"5A",X"0A",X"7F",X"10",X"60",X"0B",X"DC",X"06",X"AD",X"01",X"2A",X"FD",X"FE",X"F7",
		X"A4",X"F3",X"25",X"EE",X"5A",X"EF",X"2A",X"FA",X"BB",X"03",X"91",X"0E",X"13",X"0F",X"6A",X"09",
		X"1E",X"05",X"F4",X"FF",X"8F",X"FB",X"74",X"F6",X"22",X"F2",X"19",X"ED",X"05",X"F2",X"AD",X"FC",
		X"7D",X"06",X"BB",X"0F",X"BF",X"0D",X"86",X"08",X"0D",X"04",X"21",X"FF",X"9F",X"FA",X"BC",X"F5",
		X"3E",X"F1",X"F7",X"EC",X"7C",X"F3",X"CE",X"FD",X"CA",X"07",X"0A",X"10",X"20",X"0D",X"26",X"08",
		X"99",X"03",X"CF",X"FE",X"42",X"FA",X"7F",X"F5",X"F2",X"F0",X"F5",X"EC",X"D4",X"F3",X"0B",X"FE",
		X"FC",X"07",X"1A",X"10",X"0D",X"0D",X"1C",X"08",X"92",X"03",X"CC",X"FE",X"43",X"FA",X"80",X"F5",
		X"F9",X"F0",X"EA",X"EC",X"B2",X"F3",X"F2",X"FD",X"DB",X"07",X"2C",X"10",X"19",X"0D",X"1F",X"08",
		X"9C",X"03",X"D1",X"FE",X"4E",X"FA",X"82",X"F5",X"07",X"F1",X"E4",X"EC",X"8F",X"F3",X"D7",X"FD",
		X"BC",X"07",X"4E",X"10",X"1D",X"0D",X"26",X"08",X"A2",X"03",X"D5",X"FE",X"58",X"FA",X"86",X"F5",
		X"14",X"F1",X"CD",X"EC",X"69",X"F3",X"C0",X"FD",X"9F",X"07",X"32",X"10",X"1D",X"0D",X"30",X"08",
		X"A7",X"03",X"DE",X"FE",X"5C",X"FA",X"8F",X"F5",X"1A",X"F1",X"C6",X"EC",X"4C",X"F3",X"A7",X"FD",
		X"81",X"07",X"03",X"10",X"24",X"0D",X"3B",X"08",X"AA",X"03",X"E9",X"FE",X"5F",X"FA",X"98",X"F5",
		X"16",X"F1",X"D9",X"EC",X"61",X"F3",X"C7",X"FD",X"D0",X"07",X"17",X"10",X"C3",X"0C",X"E8",X"07",
		X"21",X"03",X"62",X"FE",X"94",X"F9",X"E3",X"F4",X"E8",X"EF",X"35",X"ED",X"2B",X"F6",X"48",X"00",
		X"11",X"0B",X"18",X"10",X"CB",X"0A",X"5B",X"06",X"1D",X"01",X"9E",X"FC",X"5E",X"F7",X"01",X"F3",
		X"74",X"ED",X"4F",X"F0",X"81",X"FB",X"76",X"05",X"6B",X"0F",X"90",X"0D",X"38",X"08",X"6A",X"03",
		X"72",X"FE",X"81",X"F9",X"B1",X"F4",X"6C",X"EF",X"A5",X"ED",X"A8",X"F7",X"CC",X"01",X"F9",X"0C",
		X"46",X"0F",X"90",X"09",X"0B",X"05",X"B3",X"FF",X"09",X"FB",X"CC",X"F5",X"0D",X"F1",X"C9",X"EC",
		X"C4",X"F4",X"67",X"FF",X"71",X"0A",X"2C",X"10",X"C7",X"0A",X"40",X"06",X"E8",X"00",X"5D",X"FC",
		X"0D",X"F7",X"A6",X"F2",X"34",X"ED",X"07",X"F1",X"14",X"FC",X"25",X"06",X"92",X"0F",X"44",X"0D",
		X"0F",X"08",X"52",X"03",X"6B",X"FE",X"A3",X"F9",X"DA",X"F4",X"E7",X"EF",X"0E",X"ED",X"0C",X"F6",
		X"17",X"00",X"D8",X"0A",X"33",X"10",X"F0",X"0A",X"8D",X"06",X"67",X"01",X"F6",X"FC",X"CF",X"F7",
		X"7A",X"F3",X"FD",X"ED",X"14",X"EF",X"C7",X"F9",X"82",X"03",X"4A",X"0E",X"AC",X"0E",X"09",X"09",
		X"99",X"04",X"66",X"FF",X"D1",X"FA",X"AF",X"F5",X"0D",X"F1",X"C5",X"EC",X"3D",X"F4",X"C0",X"FE",
		X"A5",X"09",X"46",X"10",X"37",X"0B",X"A6",X"06",X"5C",X"01",X"C7",X"FC",X"74",X"F7",X"0A",X"F3",
		X"5F",X"ED",X"47",X"F0",X"9B",X"FB",X"B9",X"05",X"92",X"0F",X"26",X"0D",X"DC",X"07",X"E9",X"02",
		X"FB",X"FD",X"E1",X"F8",X"2A",X"F4",X"A0",X"EE",X"4F",X"EE",X"25",X"F9",X"37",X"03",X"5D",X"0E",
		X"67",X"0E",X"B1",X"08",X"FF",X"03",X"C8",X"FE",X"E3",X"F9",X"DD",X"F4",X"AE",X"EF",X"56",X"ED",
		X"53",X"F7",X"A9",X"01",X"F0",X"0C",X"16",X"0F",X"57",X"09",X"BF",X"04",X"6C",X"FF",X"B4",X"FA",
		X"85",X"F5",X"B7",X"F0",X"C3",X"EC",X"05",X"F5",X"7F",X"FF",X"83",X"0A",X"2F",X"10",X"B7",X"0A",
		X"47",X"06",X"F4",X"00",X"79",X"FC",X"31",X"F7",X"E0",X"F2",X"49",X"ED",X"1A",X"F0",X"3A",X"FB",
		X"F7",X"04",X"40",X"0F",X"E4",X"0D",X"6E",X"08",X"EE",X"03",X"E7",X"FE",X"4C",X"FA",X"5A",X"F5",
		X"AE",X"F0",X"C1",X"EC",X"61",X"F4",X"B8",X"FE",X"62",X"09",X"25",X"10",X"77",X"0B",X"DF",X"06",
		X"B9",X"01",X"25",X"FD",X"F9",X"F7",X"88",X"F3",X"FD",X"ED",X"01",X"EF",X"D7",X"F9",X"BA",X"03",
		X"84",X"0E",X"4C",X"0E",X"AE",X"08",X"19",X"04",X"EE",X"FE",X"2F",X"FA",X"23",X"F5",X"3A",X"F0",
		X"DD",X"EC",X"DE",X"F5",X"32",X"00",X"64",X"0B",X"DB",X"0F",X"23",X"0A",X"AA",X"05",X"42",X"00",
		X"AA",X"FB",X"54",X"F6",X"C2",X"F1",X"BA",X"EC",X"F6",X"F2",X"EC",X"FD",X"C7",X"08",X"13",X"10",
		X"56",X"0B",X"A2",X"06",X"45",X"01",X"9E",X"FC",X"35",X"F7",X"BC",X"F2",X"10",X"ED",X"FA",X"F0",
		X"69",X"FC",X"DD",X"06",X"CF",X"0F",X"3F",X"0C",X"37",X"07",X"FE",X"01",X"33",X"FD",X"DB",X"F7",
		X"49",X"F3",X"8E",X"ED",X"EB",X"EF",X"56",X"FB",X"AA",X"05",X"85",X"0F",X"DA",X"0C",X"92",X"07",
		X"7A",X"02",X"8D",X"FD",X"49",X"F8",X"9C",X"F3",X"E9",X"ED",X"52",X"EF",X"AA",X"FA",X"F1",X"04",
		X"4B",X"0F",X"39",X"0D",X"C7",X"07",X"C2",X"02",X"C0",X"FD",X"89",X"F8",X"C9",X"F3",X"1D",X"EE",
		X"00",X"EF",X"47",X"FA",X"80",X"04",X"19",X"0F",X"82",X"0D",X"FF",X"07",X"1B",X"03",X"13",X"FE",
		X"06",X"F9",X"40",X"F4",X"D1",X"EE",X"E3",X"ED",X"60",X"F8",X"5B",X"02",X"7F",X"0D",X"DB",X"0E",
		X"2D",X"09",X"B4",X"04",X"78",X"FF",X"E1",X"FA",X"C0",X"F5",X"2B",X"F1",X"A9",X"EC",X"73",X"F3",
		X"03",X"FE",X"83",X"08",X"11",X"10",X"DA",X"0B",X"28",X"07",X"24",X"02",X"85",X"FD",X"79",X"F8",
		X"FC",X"F3",X"93",X"EE",X"F6",X"ED",X"40",X"F8",X"1C",X"02",X"09",X"0D",X"10",X"0F",X"74",X"09",
		X"02",X"05",X"C2",X"FF",X"31",X"FB",X"FD",X"F5",X"6E",X"F1",X"A3",X"EC",X"24",X"F3",X"E6",X"FD",
		X"9C",X"08",X"0E",X"10",X"8A",X"0B",X"D2",X"06",X"95",X"01",X"EE",X"FC",X"A4",X"F7",X"2C",X"F3",
		X"82",X"ED",X"BC",X"EF",X"02",X"FB",X"1A",X"05",X"4D",X"0F",X"4E",X"0D",X"E4",X"07",X"02",X"03",
		X"03",X"FE",X"F3",X"F8",X"2C",X"F4",X"B0",X"EE",X"06",X"EE",X"C9",X"F8",X"DE",X"02",X"1C",X"0E",
		X"68",X"0E",X"A9",X"08",X"FA",X"03",X"BE",X"FE",X"DB",X"F9",X"CF",X"F4",X"A1",X"EF",X"36",X"ED",
		X"26",X"F7",X"81",X"01",X"D3",X"0C",X"FD",X"0E",X"3A",X"09",X"95",X"04",X"3E",X"FF",X"6E",X"FA",
		X"3D",X"F5",X"3E",X"F0",X"C7",X"EC",X"12",X"F6",X"A8",X"00",X"F6",X"0B",X"56",X"0F",X"94",X"09",
		X"F8",X"04",X"8C",X"FF",X"CB",X"FA",X"7C",X"F5",X"9F",X"F0",X"97",X"EC",X"70",X"F5",X"26",X"00",
		X"75",X"0B",X"7F",X"0F",X"CB",X"09",X"2A",X"05",X"B9",X"FF",X"F9",X"FA",X"A6",X"F5",X"CD",X"F0",
		X"90",X"EC",X"01",X"F5",X"C5",X"FF",X"EE",X"0A",X"B3",X"0F",X"22",X"0A",X"99",X"05",X"31",X"00",
		X"9B",X"FB",X"46",X"F6",X"C0",X"F1",X"AF",X"EC",X"9B",X"F2",X"71",X"FD",X"07",X"08",X"15",X"10",
		X"E3",X"0B",X"19",X"07",X"06",X"02",X"5C",X"FD",X"47",X"F8",X"C5",X"F3",X"5E",X"EE",X"39",X"EE",
		X"A9",X"F8",X"5E",X"02",X"51",X"0D",X"05",X"0F",X"67",X"09",X"0B",X"05",X"D6",X"FF",X"59",X"FB",
		X"2B",X"F6",X"BA",X"F1",X"B0",X"EC",X"35",X"F2",X"09",X"FD",X"61",X"07",X"D0",X"0F",X"45",X"0C",
		X"57",X"07",X"54",X"02",X"93",X"FD",X"7B",X"F8",X"E2",X"F3",X"69",X"EE",X"42",X"EE",X"F3",X"F8",
		X"DD",X"02",X"05",X"0E",X"95",X"0E",X"CD",X"08",X"46",X"04",X"00",X"FF",X"4C",X"FA",X"2B",X"F5",
		X"55",X"F0",X"9B",X"EC",X"61",X"F5",X"CB",X"FF",X"C4",X"0A",X"DE",X"0F",X"77",X"0A",X"00",X"06",
		X"B7",X"00",X"3A",X"FC",X"F9",X"F6",X"A3",X"F2",X"24",X"ED",X"3D",X"F0",X"50",X"FB",X"18",X"05",
		X"20",X"0F",X"AF",X"0D",X"49",X"08",X"C3",X"03",X"C0",X"FE",X"28",X"FA",X"38",X"F5",X"98",X"F0",
		X"A1",X"EC",X"14",X"F4",X"56",X"FE",X"C3",X"08",X"FA",X"0F",X"E8",X"0B",X"32",X"07",X"5E",X"02",
		X"B7",X"FD",X"EA",X"F8",X"55",X"F4",X"62",X"EF",X"F7",X"EC",X"30",X"F6",X"E9",X"FF",X"A2",X"0A",
		X"24",X"10",X"08",X"0B",X"AD",X"06",X"B2",X"01",X"41",X"FD",X"5A",X"F8",X"F6",X"F3",X"DC",X"EE",
		X"5A",X"ED",X"F7",X"F6",X"80",X"00",X"34",X"0B",X"0C",X"10",X"CB",X"0A",X"8A",X"06",X"7F",X"01",
		X"1E",X"FD",X"23",X"F8",X"CC",X"F3",X"88",X"EE",X"BE",X"ED",X"D1",X"F7",X"70",X"01",X"58",X"0C",
		X"AA",X"0F",X"EE",X"09",X"BA",X"05",X"72",X"00",X"17",X"FC",X"D7",X"F6",X"92",X"F2",X"1C",X"ED",
		X"75",X"F0",X"58",X"FB",X"51",X"05",X"43",X"0F",X"71",X"0D",X"19",X"08",X"6A",X"03",X"68",X"FE",
		X"9B",X"F9",X"BA",X"F4",X"B7",X"EF",X"08",X"ED",X"43",X"F6",X"4C",X"00",X"64",X"0B",X"CC",X"0F",
		X"4D",X"0A",X"F3",X"05",X"B1",X"00",X"44",X"FC",X"0D",X"F7",X"C6",X"F2",X"46",X"ED",X"EC",X"EF",
		X"B1",X"FA",X"72",X"04",X"8C",X"0E",X"1C",X"0E",X"AA",X"08",X"47",X"04",X"32",X"FF",X"C2",X"FA",
		X"B4",X"F5",X"59",X"F1",X"88",X"EC",X"71",X"F2",X"04",X"FD",X"F6",X"06",X"D2",X"0F",X"E7",X"0C",
		X"E4",X"07",X"51",X"03",X"7C",X"FE",X"EC",X"F9",X"18",X"F5",X"8E",X"F0",X"8B",X"EC",X"C2",X"F3",
		X"01",X"FE",X"1E",X"08",X"26",X"10",X"65",X"0C",X"9A",X"07",X"F4",X"02",X"3F",X"FE",X"A7",X"F9",
		X"F1",X"F4",X"5A",X"F0",X"87",X"EC",X"00",X"F4",X"28",X"FE",X"3C",X"08",X"09",X"10",X"5E",X"0C",
		X"A0",X"07",X"F6",X"02",X"4A",X"FE",X"AD",X"F9",X"FD",X"F4",X"61",X"F0",X"99",X"EC",X"EB",X"F3",
		X"14",X"FE",X"20",X"08",X"E5",X"0F",X"6E",X"0C",X"A9",X"07",X"02",X"03",X"54",X"FE",X"B8",X"F9",
		X"0A",X"F5",X"6C",X"F0",X"AA",X"EC",X"D6",X"F3",X"FE",X"FD",X"06",X"08",X"D0",X"0F",X"83",X"0C",
		X"B1",X"07",X"12",X"03",X"60",X"FE",X"C6",X"F9",X"14",X"F5",X"77",X"F0",X"AD",X"EC",X"BC",X"F3",
		X"EB",X"FD",X"E6",X"07",X"CC",X"0F",X"95",X"0C",X"B7",X"07",X"21",X"03",X"67",X"FE",X"D4",X"F9",
		X"1C",X"F5",X"86",X"F0",X"A0",X"EC",X"A3",X"F3",X"D5",X"FD",X"CA",X"07",X"D9",X"0F",X"A9",X"0C",
		X"BD",X"07",X"31",X"03",X"6F",X"FE",X"E3",X"F9",X"22",X"F5",X"97",X"F0",X"9E",X"EC",X"86",X"F3",
		X"BF",X"FD",X"B2",X"07",X"F5",X"0F",X"B6",X"0C",X"C8",X"07",X"41",X"03",X"77",X"FE",X"F3",X"F9",
		X"2B",X"F5",X"AC",X"F0",X"95",X"EC",X"69",X"F3",X"AB",X"FD",X"9A",X"07",X"1A",X"10",X"C0",X"0C",
		X"D3",X"07",X"4C",X"03",X"82",X"FE",X"01",X"FA",X"32",X"F5",X"BE",X"F0",X"7C",X"EC",X"47",X"F3",
		X"97",X"FD",X"81",X"07",X"E8",X"0F",X"C8",X"0C",X"E2",X"07",X"54",X"03",X"90",X"FE",X"07",X"FA",
		X"41",X"F5",X"C7",X"F0",X"91",X"EC",X"37",X"F3",X"81",X"FD",X"68",X"07",X"C2",X"0F",X"D6",X"0C",
		X"EE",X"07",X"61",X"03",X"9C",X"FE",X"14",X"FA",X"4E",X"F5",X"CF",X"F0",X"A3",X"EC",X"23",X"F3",
		X"6B",X"FD",X"4D",X"07",X"AB",X"0F",X"E9",X"0C",X"F5",X"07",X"6E",X"03",X"A8",X"FE",X"22",X"FA",
		X"58",X"F5",X"DC",X"F0",X"A9",X"EC",X"0A",X"F3",X"56",X"FD",X"31",X"07",X"A4",X"0F",X"FE",X"0C",
		X"FC",X"07",X"7D",X"03",X"AF",X"FE",X"30",X"FA",X"63",X"F5",X"EB",X"F0",X"9E",X"EC",X"EF",X"F2",
		X"42",X"FD",X"15",X"07",X"B0",X"0F",X"12",X"0D",X"03",X"08",X"8E",X"03",X"B8",X"FE",X"3F",X"FA",
		X"6C",X"F5",X"FB",X"F0",X"A1",X"EC",X"D2",X"F2",X"2F",X"FD",X"FA",X"06",X"CA",X"0F",X"23",X"0D",
		X"0B",X"08",X"9C",X"03",X"C0",X"FE",X"4F",X"FA",X"72",X"F5",X"10",X"F1",X"9B",X"EC",X"B3",X"F2",
		X"1B",X"FD",X"DF",X"06",X"ED",X"0F",X"2E",X"0D",X"17",X"08",X"AB",X"03",X"CB",X"FE",X"5F",X"FA",
		X"79",X"F5",X"22",X"F1",X"88",X"EC",X"92",X"F2",X"09",X"FD",X"C9",X"06",X"BA",X"0F",X"30",X"0D",
		X"2A",X"08",X"B2",X"03",X"DB",X"FE",X"64",X"FA",X"8A",X"F5",X"24",X"F1",X"97",X"EC",X"AB",X"F2",
		X"31",X"FD",X"1E",X"07",X"DD",X"0F",X"D0",X"0C",X"DE",X"07",X"26",X"03",X"5C",X"FE",X"98",X"F9",
		X"DC",X"F4",X"F1",X"EF",X"EC",X"EC",X"86",X"F5",X"B6",X"FF",X"73",X"0A",X"EC",X"0F",X"D9",X"0A",
		X"55",X"06",X"26",X"01",X"A1",X"FC",X"74",X"F7",X"16",X"F3",X"97",X"ED",X"5F",X"EF",X"5A",X"FA",
		X"FF",X"03",X"84",X"0E",X"5F",X"0E",X"CB",X"08",X"68",X"04",X"4F",X"FF",X"D2",X"FA",X"C8",X"F5",
		X"58",X"F1",X"AF",X"EC",X"B1",X"F2",X"34",X"FD",X"4B",X"07",X"C1",X"0F",X"C4",X"0C",X"CE",X"07",
		X"26",X"03",X"5C",X"FE",X"B7",X"F9",X"F6",X"F4",X"48",X"F0",X"A3",X"EC",X"87",X"F4",X"A4",X"FE",
		X"F5",X"08",X"24",X"10",X"FC",X"0B",X"5C",X"07",X"91",X"02",X"F7",X"FD",X"3C",X"F9",X"A6",X"F4",
		X"D7",X"EF",X"C4",X"EC",X"2F",X"F5",X"19",X"FF",X"6F",X"09",X"20",X"10",X"D3",X"0B",X"48",X"07",
		X"7B",X"02",X"F0",X"FD",X"31",X"F9",X"A8",X"F4",X"D4",X"EF",X"E0",X"EC",X"20",X"F5",X"0A",X"FF",
		X"50",X"09",X"08",X"10",X"E8",X"0B",X"51",X"07",X"89",X"02",X"FA",X"FD",X"3E",X"F9",X"B5",X"F4",
		X"E0",X"EF",X"EC",X"EC",X"06",X"F5",X"F8",X"FE",X"32",X"09",X"00",X"10",X"FA",X"0B",X"5A",X"07",
		X"99",X"02",X"04",X"FE",X"4D",X"F9",X"BF",X"F4",X"EF",X"EF",X"E7",X"EC",X"EB",X"F4",X"E6",X"FE",
		X"14",X"09",X"0A",X"10",X"0B",X"0C",X"64",X"07",X"A6",X"02",X"11",X"FE",X"59",X"F9",X"CB",X"F4",
		X"F9",X"EF",X"DA",X"EC",X"E4",X"F4",X"F3",X"FE",X"3B",X"09",X"19",X"10",X"CE",X"0B",X"2C",X"07",
		X"43",X"02",X"AD",X"FD",X"BC",X"F8",X"3B",X"F4",X"05",X"EF",X"9A",X"ED",X"60",X"F7",X"32",X"01",
		X"31",X"0C",X"A2",X"0F",X"0E",X"0A",X"BA",X"05",X"70",X"00",X"FE",X"FB",X"B9",X"F6",X"5F",X"F2",
		X"FE",X"EC",X"4A",X"F1",X"3D",X"FC",X"76",X"06",X"BC",X"0F",X"D6",X"0C",X"B9",X"07",X"CF",X"02",
		X"F0",X"FD",X"EA",X"F8",X"34",X"F4",X"D3",X"EE",X"F2",X"ED",X"81",X"F8",X"70",X"02",X"BA",X"0D",
		X"F1",X"0E",X"09",X"09",X"8C",X"04",X"3A",X"FF",X"89",X"FA",X"5D",X"F5",X"7F",X"F0",X"D9",X"EC",
		X"87",X"F5",X"09",X"00",X"42",X"0B",X"B8",X"0F",X"2F",X"0A",X"9F",X"05",X"39",X"00",X"94",X"FB",
		X"37",X"F6",X"9C",X"F1",X"A0",X"EC",X"72",X"F3",X"7D",X"FE",X"63",X"09",X"10",X"10",X"00",X"0B",
		X"51",X"06",X"E9",X"00",X"3F",X"FC",X"D5",X"F6",X"47",X"F2",X"E2",X"EC",X"37",X"F2",X"6D",X"FD",
		X"31",X"08",X"2C",X"10",X"94",X"0B",X"BA",X"06",X"60",X"01",X"A6",X"FC",X"3E",X"F7",X"AB",X"F2",
		X"1A",X"ED",X"76",X"F1",X"CA",X"FC",X"72",X"07",X"31",X"10",X"EC",X"0B",X"F8",X"06",X"A7",X"01",
		X"E1",X"FC",X"79",X"F7",X"E2",X"F2",X"3C",X"ED",X"12",X"F1",X"72",X"FC",X"10",X"07",X"27",X"10",
		X"1E",X"0C",X"15",X"07",X"CB",X"01",X"FA",X"FC",X"95",X"F7",X"F9",X"F2",X"4D",X"ED",X"E9",X"F0",
		X"55",X"FC",X"E9",X"06",X"18",X"10",X"3A",X"0C",X"2F",X"07",X"F4",X"01",X"2D",X"FD",X"DC",X"F7",
		X"50",X"F3",X"A0",X"ED",X"DD",X"EF",X"0A",X"FB",X"2D",X"05",X"60",X"0F",X"77",X"0D",X"21",X"08",
		X"57",X"03",X"60",X"FE",X"7D",X"F9",X"AF",X"F4",X"91",X"EF",X"4D",X"ED",X"DD",X"F6",X"CF",X"00",
		X"F3",X"0B",X"E3",X"0F",X"38",X"0A",X"F0",X"05",X"A6",X"00",X"44",X"FC",X"06",X"F7",X"C8",X"F2",
		X"4E",X"ED",X"47",X"F0",X"06",X"FB",X"CC",X"04",X"CB",X"0E",X"26",X"0E",X"BC",X"08",X"58",X"04",
		X"46",X"FF",X"D7",X"FA",X"CD",X"F5",X"71",X"F1",X"A7",X"EC",X"A0",X"F2",X"2E",X"FD",X"21",X"07",
		X"F4",X"0F",X"08",X"0D",X"07",X"08",X"76",X"03",X"A2",X"FE",X"13",X"FA",X"41",X"F5",X"BA",X"F0",
		X"A8",X"EC",X"D3",X"F3",X"15",X"FE",X"28",X"08",X"3C",X"10",X"96",X"0C",X"C9",X"07",X"27",X"03",
		X"70",X"FE",X"DA",X"F9",X"20",X"F5",X"91",X"F0",X"A3",X"EC",X"FD",X"F3",X"2F",X"FE",X"38",X"08",
		X"1D",X"10",X"95",X"0C",X"D2",X"07",X"2E",X"03",X"7E",X"FE",X"E2",X"F9",X"32",X"F5",X"98",X"F0",
		X"C1",X"EC",X"EC",X"F3",X"1B",X"FE",X"20",X"08",X"FD",X"0F",X"A9",X"0C",X"DD",X"07",X"3C",X"03",
		X"89",X"FE",X"EF",X"F9",X"3E",X"F5",X"A5",X"F0",X"D0",X"EC",X"D6",X"F3",X"07",X"FE",X"04",X"08",
		X"EE",X"0F",X"BE",X"0C",X"E3",X"07",X"4A",X"03",X"93",X"FE",X"FE",X"F9",X"48",X"F5",X"B2",X"F0",
		X"D0",X"EC",X"BF",X"F3",X"F4",X"FD",X"E8",X"07",X"EE",X"0F",X"D4",X"0C",X"EA",X"07",X"5B",X"03",
		X"9E",X"FE",X"0E",X"FA",X"51",X"F5",X"C3",X"F0",X"C2",X"EC",X"A3",X"F3",X"DF",X"FD",X"CD",X"07",
		X"FF",X"0F",X"E5",X"0C",X"F2",X"07",X"6B",X"03",X"A4",X"FE",X"1F",X"FA",X"5B",X"F5",X"D5",X"F0",
		X"C7",X"EC",X"87",X"F3",X"CC",X"FD",X"B3",X"07",X"22",X"10",X"F2",X"0C",X"00",X"08",X"79",X"03",
		X"B1",X"FE",X"2C",X"FA",X"63",X"F5",X"E9",X"F0",X"BC",X"EC",X"67",X"F3",X"BA",X"FD",X"99",X"07",
		X"34",X"10",X"F5",X"0C",X"0F",X"08",X"77",X"03",X"B0",X"FE",X"14",X"FA",X"4C",X"F5",X"A6",X"F0",
		X"CB",X"EC",X"46",X"F4",X"A1",X"FE",X"F7",X"08",X"54",X"10",X"F0",X"0B",X"44",X"07",X"47",X"02",
		X"A7",X"FD",X"A4",X"F8",X"1F",X"F4",X"C9",X"EE",X"17",X"EE",X"6E",X"F8",X"2E",X"02",X"61",X"0D",
		X"5F",X"0F",X"8D",X"09",X"35",X"05",X"E3",X"FF",X"5F",X"FB",X"21",X"F6",X"9E",X"F1",X"C6",X"EC",
		X"4E",X"F3",X"1C",X"FE",X"C5",X"08",X"66",X"10",X"AD",X"0B",X"F7",X"06",X"BB",X"01",X"15",X"FD",
		X"CB",X"F7",X"4F",X"F3",X"AE",X"ED",X"FF",X"EF",X"36",X"FB",X"69",X"05",X"61",X"0F",X"61",X"0D",
		X"0D",X"08",X"20",X"03",X"28",X"FE",X"12",X"F9",X"51",X"F4",X"D4",X"EE",X"44",X"EE",X"15",X"F9",
		X"2C",X"03",X"49",X"0E",X"92",X"0E",X"C5",X"08",X"1A",X"04",X"DB",X"FE",X"FA",X"F9",X"EE",X"F4",
		X"BD",X"EF",X"77",X"ED",X"96",X"F7",X"C0",X"01",X"68",X"0D",X"52",X"0F",X"43",X"09",X"BE",X"04",
		X"52",X"FF",X"8F",X"FA",X"56",X"F5",X"52",X"F0",X"1C",X"ED",X"91",X"F6",X"F2",X"00",X"8D",X"0C",
		X"91",X"0F",X"A4",X"09",X"15",X"05",X"A4",X"FF",X"E0",X"FA",X"9A",X"F5",X"A9",X"F0",X"00",X"ED",
		X"F6",X"F5",X"84",X"00",X"0F",X"0C",X"B9",X"0F",X"D5",X"09",X"49",X"05",X"CC",X"FF",X"12",X"FB",
		X"BB",X"F5",X"D9",X"F0",X"EF",X"EC",X"B5",X"F5",X"4D",X"00",X"E0",X"0B",X"CC",X"0F",X"EC",X"09",
		X"58",X"05",X"E1",X"FF",X"22",X"FB",X"D1",X"F5",X"F9",X"F0",X"E8",X"EC",X"39",X"F5",X"D5",X"FF",
		X"15",X"0B",X"FE",X"0F",X"7B",X"0A",X"FB",X"05",X"9A",X"00",X"0C",X"FC",X"B7",X"F6",X"47",X"F2",
		X"FB",X"EC",X"0E",X"F2",X"0F",X"FD",X"53",X"07",X"47",X"10",X"A8",X"0C",X"AA",X"07",X"C4",X"02",
		X"FE",X"FD",X"0C",X"F9",X"6B",X"F4",X"36",X"EF",X"B9",X"ED",X"A7",X"F7",X"65",X"01",X"74",X"0C",
		X"DC",X"0F",X"41",X"0A",X"FE",X"05",X"C6",X"00",X"68",X"FC",X"3E",X"F7",X"00",X"F3",X"90",X"ED",
		X"F8",X"EF",X"AC",X"FA",X"44",X"04",X"88",X"0E",X"B0",X"0E",X"2E",X"09",X"E2",X"04",X"CE",X"FF",
		X"6E",X"FB",X"62",X"F6",X"1D",X"F2",X"11",X"ED",X"83",X"F1",X"1A",X"FC",X"C5",X"05",X"45",X"0F",
		X"03",X"0E",X"BE",X"08",X"5F",X"04",X"6D",X"FF",X"04",X"FB",X"15",X"F6",X"C3",X"F1",X"FA",X"EC",
		X"09",X"F2",X"87",X"FC",X"28",X"06",X"71",X"0F",X"E6",X"0D",X"AF",X"08",X"50",X"04",X"68",X"FF",
		X"01",X"FB",X"18",X"F6",X"C8",X"F1",X"F5",X"EC",X"F1",X"F1",X"77",X"FC",X"0B",X"06",X"77",X"0F",
		X"FA",X"0D",X"B6",X"08",X"61",X"04",X"72",X"FF",X"0F",X"FB",X"23",X"F6",X"D7",X"F1",X"FF",X"EC",
		X"D5",X"F1",X"66",X"FC",X"EE",X"05",X"90",X"0F",X"11",X"0E",X"BC",X"08",X"72",X"04",X"79",X"FF",
		X"20",X"FB",X"29",X"F6",X"EB",X"F1",X"FD",X"EC",X"B4",X"F1",X"53",X"FC",X"D3",X"05",X"A8",X"0F",
		X"20",X"0E",X"C7",X"08",X"82",X"04",X"83",X"FF",X"30",X"FB",X"30",X"F6",X"00",X"F2",X"EF",X"EC",
		X"94",X"F1",X"40",X"FC",X"BF",X"05",X"77",X"0F",X"1D",X"0E",X"DC",X"08",X"83",X"04",X"89",X"FF",
		X"21",X"FB",X"21",X"F6",X"D0",X"F1",X"DA",X"EC",X"45",X"F2",X"0F",X"FD",X"EF",X"06",X"40",X"10",
		X"35",X"0D",X"1E",X"08",X"6B",X"03",X"8F",X"FE",X"C6",X"F9",X"00",X"F5",X"05",X"F0",X"4A",X"ED",
		X"55",X"F6",X"69",X"00",X"6D",X"0B",X"13",X"10",X"B6",X"0A",X"4C",X"06",X"0C",X"01",X"95",X"FC",
		X"5B",X"F7",X"0B",X"F3",X"8B",X"ED",X"53",X"F0",X"2C",X"FB",X"F8",X"04",X"06",X"0F",X"3A",X"0E",
		X"D5",X"08",X"5E",X"04",X"53",X"FF",X"D0",X"FA",X"CE",X"F5",X"5A",X"F1",X"CA",X"EC",X"62",X"F3",
		X"EC",X"FD",X"03",X"08",X"7C",X"10",X"BF",X"0C",X"E8",X"07",X"2E",X"03",X"75",X"FE",X"C2",X"F9",
		X"14",X"F5",X"4C",X"F0",X"14",X"ED",X"2F",X"F5",X"37",X"FF",X"8E",X"09",X"71",X"10",X"17",X"0C",
		X"76",X"07",X"AE",X"02",X"15",X"FE",X"5A",X"F9",X"C9",X"F4",X"EF",X"EF",X"38",X"ED",X"C3",X"F5",
		X"94",X"FF",X"F9",X"09",X"83",X"10",X"F4",X"0B",X"6A",X"07",X"A1",X"02",X"10",X"FE",X"59",X"F9",
		X"CA",X"F4",X"FB",X"EF",X"23",X"ED",X"AD",X"F5",X"80",X"FF",X"E8",X"09",X"8D",X"10",X"FC",X"0B",
		X"7C",X"07",X"AB",X"02",X"1F",X"FE",X"64",X"F9",X"D9",X"F4",X"08",X"F0",X"0E",X"ED",X"91",X"F5",
		X"71",X"FF",X"C9",X"09",X"66",X"10",X"0E",X"0C",X"87",X"07",X"B7",X"02",X"2D",X"FE",X"6E",X"F9",
		X"E7",X"F4",X"0F",X"F0",X"28",X"ED",X"78",X"F5",X"61",X"FF",X"A9",X"09",X"50",X"10",X"22",X"0C",
		X"91",X"07",X"C6",X"02",X"39",X"FE",X"74",X"F9",X"ED",X"F4",X"05",X"F0",X"45",X"ED",X"CF",X"F5",
		X"C9",X"FF",X"58",X"0A",X"53",X"10",X"8B",X"0B",X"13",X"07",X"FD",X"01",X"7E",X"FD",X"67",X"F8",
		X"04",X"F4",X"95",X"EE",X"9F",X"EE",X"18",X"F9",X"E7",X"02",X"AF",X"0D",X"44",X"0F",X"94",X"09",
		X"32",X"05",X"F1",X"FF",X"70",X"FB",X"41",X"F6",X"CC",X"F1",X"F1",X"EC",X"08",X"F3",X"CF",X"FD",
		X"0D",X"08",X"49",X"10",X"9F",X"0C",X"B8",X"07",X"DF",X"02",X"24",X"FE",X"46",X"F9",X"AA",X"F4",
		X"92",X"EF",X"9C",X"ED",X"10",X"F7",X"D6",X"00",X"B1",X"0B",X"29",X"10",X"EE",X"0A",X"96",X"06",
		X"7E",X"01",X"14",X"FD",X"0B",X"F8",X"BF",X"F3",X"65",X"EE",X"B6",X"EE",X"3D",X"F9",X"B2",X"02",
		X"9D",X"0D",X"AB",X"0F",X"E5",X"09",X"B0",X"05",X"71",X"00",X"15",X"FC",X"DC",X"F6",X"94",X"F2",
		X"44",X"ED",X"83",X"F1",X"57",X"FC",X"68",X"06",X"D1",X"0F",X"6D",X"0D",X"3B",X"08",X"76",X"03",
		X"88",X"FE",X"A9",X"F9",X"DC",X"F4",X"BA",X"EF",X"9F",X"ED",X"56",X"F7",X"5C",X"01",X"9C",X"0C",
		X"C1",X"0F",X"08",X"0A",X"9A",X"05",X"3F",X"00",X"AC",X"FB",X"62",X"F6",X"D3",X"F1",X"E6",X"EC",
		X"5F",X"F3",X"4C",X"FE",X"03",X"09",X"5E",X"10",X"9E",X"0B",X"E1",X"06",X"97",X"01",X"ED",X"FC",
		X"95",X"F7",X"14",X"F3",X"76",X"ED",X"E0",X"F0",X"19",X"FC",X"81",X"06",X"06",X"10",X"CC",X"0C",
		X"AF",X"07",X"8E",X"02",X"B4",X"FD",X"74",X"F8",X"D2",X"F3",X"27",X"EE",X"53",X"EF",X"94",X"FA",
		X"D4",X"04",X"35",X"0F",X"99",X"0D",X"2F",X"08",X"34",X"03",X"31",X"FE",X"08",X"F9",X"44",X"F4",
		X"AD",X"EE",X"77",X"EE",X"8F",X"F9",X"C8",X"03",X"9F",X"0E",X"15",X"0E",X"7B",X"08",X"9B",X"03",
		X"78",X"FE",X"64",X"F9",X"80",X"F4",X"07",X"EF",X"1E",X"EE",X"EA",X"F8",X"33",X"03",X"3C",X"0E",
		X"58",X"0E",X"A3",X"08",X"CF",X"03",X"9D",X"FE",X"91",X"F9",X"9C",X"F4",X"31",X"EF",X"F0",X"ED",
		X"95",X"F8",X"E8",X"02",X"08",X"0E",X"6E",X"0E",X"AF",X"08",X"E1",X"03",X"A6",X"FE",X"9F",X"F9",
		X"9F",X"F4",X"39",X"EF",X"D8",X"ED",X"80",X"F8",X"D6",X"02",X"FE",X"0D",X"64",X"0E",X"AC",X"08",
		X"D3",X"03",X"9E",X"FE",X"8E",X"F9",X"9A",X"F4",X"2F",X"EF",X"C6",X"ED",X"57",X"F8",X"9C",X"02",
		X"B2",X"0D",X"A5",X"0E",X"E8",X"08",X"48",X"04",X"08",X"FF",X"43",X"FA",X"2C",X"F5",X"46",X"F0",
		X"17",X"ED",X"BF",X"F5",X"FE",X"FF",X"2B",X"0B",X"F8",X"0F",X"6C",X"0A",X"04",X"06",X"BB",X"00",
		X"3D",X"FC",X"03",X"F7",X"9D",X"F2",X"5A",X"ED",X"8F",X"F0",X"4F",X"FB",X"40",X"05",X"33",X"0F",
		X"A5",X"0D",X"48",X"08",X"AF",X"03",X"A7",X"FE",X"F3",X"F9",X"01",X"F5",X"27",X"F0",X"13",X"ED",
		X"8A",X"F5",X"C9",X"FF",X"D1",X"0A",X"DD",X"0F",X"86",X"0A",X"08",X"06",X"BD",X"00",X"2B",X"FC",
		X"E8",X"F6",X"65",X"F2",X"2C",X"ED",X"3A",X"F1",X"34",X"FC",X"8C",X"06",X"F1",X"0F",X"8F",X"0C",
		X"69",X"07",X"69",X"02",X"8B",X"FD",X"69",X"F8",X"BF",X"F3",X"34",X"EE",X"93",X"EE",X"93",X"F9",
		X"AF",X"03",X"69",X"0E",X"EC",X"0D",X"60",X"08",X"94",X"03",X"76",X"FE",X"7F",X"F9",X"8F",X"F4",
		X"4D",X"EF",X"9B",X"ED",X"97",X"F7",X"DF",X"01",X"14",X"0D",X"DC",X"0E",X"F9",X"08",X"65",X"04",
		X"06",X"FF",X"41",X"FA",X"0D",X"F5",X"11",X"F0",X"2A",X"ED",X"43",X"F6",X"A4",X"00",X"18",X"0C",
		X"76",X"0F",X"83",X"09",X"0D",X"05",X"A4",X"FF",X"09",X"FB",X"C0",X"F5",X"20",X"F1",X"AE",X"EC",
		X"93",X"F3",X"4C",X"FE",X"04",X"09",X"D9",X"0F",X"43",X"0B",X"97",X"06",X"71",X"01",X"D5",X"FC",
		X"B3",X"F7",X"3A",X"F3",X"EA",X"ED",X"F8",X"EE",X"7E",X"F9",X"58",X"03",X"D1",X"0D",X"77",X"0E",
		X"E3",X"08",X"86",X"04",X"5F",X"FF",X"EA",X"FA",X"D3",X"F5",X"6B",X"F1",X"B2",X"EC",X"29",X"F2",
		X"AA",X"FC",X"B3",X"06",X"C8",X"0F",X"DC",X"0C",X"BB",X"07",X"30",X"03",X"49",X"FE",X"BB",X"F9",
		X"DE",X"F4",X"4D",X"F0",X"BA",X"EC",X"10",X"F4",X"43",X"FE",X"7B",X"08",X"E9",X"0F",X"FA",X"0B",
		X"35",X"07",X"82",X"02",X"D1",X"FD",X"29",X"F9",X"7A",X"F4",X"C4",X"EF",X"F7",X"EC",X"F7",X"F4",
		X"07",X"FF",X"70",X"09",X"E2",X"0F",X"56",X"0B",X"BB",X"06",X"CB",X"01",X"2D",X"FD",X"3F",X"F8",
		X"AE",X"F3",X"92",X"EE",X"10",X"EE",X"D6",X"F7",X"AA",X"01",X"AB",X"0C",X"20",X"0F",X"6A",X"09",
		X"19",X"05",X"CE",X"FF",X"50",X"FB",X"1B",X"F6",X"98",X"F1",X"EB",X"EC",X"24",X"F2",X"CE",X"FC",
		X"56",X"07",X"C5",X"0F",X"0C",X"0C",X"16",X"07",X"28",X"02",X"5A",X"FD",X"69",X"F8",X"B8",X"F3",
		X"9F",X"EE",X"10",X"EE",X"D3",X"F7",X"B3",X"01",X"A0",X"0C",X"10",X"0F",X"74",X"09",X"26",X"05",
		X"F1",X"FF",X"84",X"FB",X"64",X"F6",X"08",X"F2",X"14",X"ED",X"8B",X"F0",X"3F",X"FB",X"01",X"05",
		X"C7",X"0E",X"9D",X"0D",X"39",X"08",X"CF",X"03",X"CD",X"FE",X"49",X"FA",X"57",X"F5",X"C6",X"F0",
		X"D9",X"EC",X"12",X"F3",X"6E",X"FD",X"D6",X"07",X"AB",X"0F",X"EC",X"0B",X"0D",X"07",X"2B",X"02",
		X"65",X"FD",X"7E",X"F8",X"C6",X"F3",X"BE",X"EE",X"E1",X"ED",X"A0",X"F7",X"AF",X"01",X"9A",X"0C",
		X"DF",X"0E",X"34",X"09",X"C6",X"04",X"7A",X"FF",X"E8",X"FA",X"B0",X"F5",X"11",X"F1",X"DD",X"EC",
		X"28",X"F3",X"C8",X"FD",X"AC",X"08",X"DF",X"0F",X"13",X"0B",X"60",X"06",X"22",X"01",X"71",X"FC",
		X"2F",X"F7",X"9A",X"F2",X"4A",X"ED",X"3D",X"F0",X"29",X"FB",X"8D",X"05",X"1D",X"0F",X"A7",X"0C",
		X"50",X"07",X"67",X"02",X"61",X"FD",X"57",X"F8",X"78",X"F3",X"47",X"EE",X"BB",X"EE",X"3B",X"F9",
		X"80",X"03",X"6A",X"0E",X"BF",X"0D",X"EB",X"07",X"45",X"03",X"FC",X"FD",X"21",X"F9",X"06",X"F4",
		X"FF",X"EE",X"D5",X"ED",X"E7",X"F7",X"3B",X"02",X"8F",X"0D",X"4E",X"0E",X"5F",X"08",X"C6",X"03",
		X"68",X"FE",X"99",X"F9",X"66",X"F4",X"70",X"EF",X"5D",X"ED",X"0C",X"F7",X"7F",X"01",X"E2",X"0C",
		X"96",X"0E",X"A9",X"08",X"12",X"04",X"A6",X"FE",X"DC",X"F9",X"9A",X"F4",X"B2",X"EF",X"20",X"ED",
		X"6E",X"F6",X"EB",X"00",X"35",X"0C",X"E0",X"0E",X"18",X"09",X"94",X"04",X"3A",X"FF",X"92",X"FA",
		X"5D",X"F5",X"9F",X"F0",X"D3",X"EC",X"E2",X"F3",X"4B",X"FE",X"37",X"09",X"CC",X"0F",X"DE",X"0A",
		X"34",X"06",X"1B",X"01",X"71",X"FC",X"64",X"F7",X"CE",X"F2",X"C6",X"ED",X"33",X"EF",X"7B",X"F9",
		X"45",X"03",X"0A",X"0E",X"4E",X"0E",X"82",X"08",X"41",X"04",X"0A",X"FF",X"A2",X"FA",X"89",X"F5",
		X"17",X"F1",X"EC",X"EC",X"26",X"F2",X"80",X"FC",X"AD",X"06",X"31",X"0F",X"9B",X"0C",X"76",X"07",
		X"F1",X"02",X"08",X"FE",X"7C",X"F9",X"A1",X"F4",X"07",X"F0",X"F9",X"EC",X"0D",X"F4",X"02",X"FE",
		X"6D",X"08",X"8F",X"0F",X"C6",X"0B",X"F7",X"06",X"52",X"02",X"92",X"FD",X"FA",X"F8",X"40",X"F4",
		X"9C",X"EF",X"29",X"ED",X"B2",X"F4",X"8C",X"FE",X"F1",X"08",X"93",X"0F",X"8D",X"0B",X"DB",X"06",
		X"30",X"02",X"83",X"FD",X"E5",X"F8",X"3D",X"F4",X"8E",X"EF",X"2B",X"ED",X"A0",X"F4",X"82",X"FE",
		X"D0",X"08",X"89",X"0F",X"9A",X"0B",X"E3",X"06",X"39",X"02",X"8A",X"FD",X"EF",X"F8",X"42",X"F4",
		X"9F",X"EF",X"2A",X"ED",X"75",X"F4",X"75",X"FE",X"AE",X"08",X"91",X"0F",X"94",X"0B",X"D9",X"06",
		X"19",X"02",X"68",X"FD",X"AE",X"F8",X"FA",X"F3",X"28",X"EF",X"7E",X"ED",X"E3",X"F5",X"E2",X"FF",
		X"AE",X"0A",X"70",X"0F",X"39",X"0A",X"CB",X"05",X"A2",X"00",X"18",X"FC",X"00",X"F7",X"75",X"F2",
		X"9B",X"ED",X"AB",X"EF",X"28",X"FA",X"4F",X"04",X"56",X"0E",X"74",X"0D",X"E9",X"07",X"59",X"03",
		X"2D",X"FE",X"81",X"F9",X"69",X"F4",X"A8",X"EF",X"50",X"ED",X"BB",X"F5",X"12",X"00",X"43",X"0B",
		X"42",X"0F",X"96",X"09",X"21",X"05",X"C4",X"FF",X"29",X"FB",X"E3",X"F5",X"3B",X"F1",X"17",X"ED",
		X"AF",X"F2",X"53",X"FD",X"39",X"08",X"8D",X"0F",X"14",X"0B",X"2B",X"06",X"02",X"01",X"2D",X"FC",
		X"05",X"F7",X"3F",X"F2",X"7D",X"ED",X"75",X"F0",X"25",X"FB",X"9B",X"05",X"28",X"0F",X"94",X"0C",
		X"48",X"07",X"84",X"02",X"80",X"FD",X"B3",X"F8",X"C7",X"F3",X"F9",X"EE",X"ED",X"ED",X"F0",X"F6",
		X"F8",X"00",X"0E",X"0C",X"2D",X"0F",X"61",X"09",X"20",X"05",X"DA",X"FF",X"6F",X"FB",X"4C",X"F6",
		X"D5",X"F1",X"4D",X"ED",X"A8",X"F0",X"E7",X"FA",X"00",X"05",X"81",X"0E",X"5F",X"0D",X"EB",X"07",
		X"92",X"03",X"7A",X"FE",X"0E",X"FA",X"08",X"F5",X"9A",X"F0",X"2F",X"ED",X"F3",X"F2",X"02",X"FD",
		X"4F",X"07",X"79",X"0F",X"3F",X"0C",X"39",X"07",X"B4",X"02",X"D2",X"FD",X"52",X"F9",X"72",X"F4",
		X"FE",X"EF",X"4F",X"ED",X"FD",X"F3",X"ED",X"FD",X"44",X"08",X"B4",X"0F",X"C7",X"0B",X"FB",X"06",
		X"59",X"02",X"94",X"FD",X"FE",X"F8",X"2C",X"F4",X"A4",X"EF",X"7C",X"ED",X"EE",X"F4",X"F4",X"FE",
		X"9A",X"09",X"B9",X"0F",X"C9",X"0A",X"37",X"06",X"3B",X"01",X"90",X"FC",X"A6",X"F7",X"F0",X"F2",
		X"47",X"EE",X"E7",X"EE",X"91",X"F8",X"A9",X"02",X"64",X"0D",X"56",X"0E",X"87",X"08",X"32",X"04",
		X"DE",X"FE",X"5C",X"FA",X"25",X"F5",X"91",X"F0",X"3F",X"ED",X"C3",X"F3",X"25",X"FE",X"35",X"09",
		X"D5",X"0F",X"9E",X"0A",X"FC",X"05",X"C2",X"00",X"0E",X"FC",X"E3",X"F6",X"29",X"F2",X"AB",X"ED",
		X"B4",X"F0",X"23",X"FB",X"BF",X"05",X"F6",X"0E",X"6E",X"0C",X"09",X"07",X"37",X"02",X"1D",X"FD",
		X"35",X"F8",X"2C",X"F3",X"77",X"EE",X"F6",X"EE",X"FF",X"F8",X"69",X"03",X"36",X"0E",X"A7",X"0D",
		X"C2",X"07",X"32",X"03",X"D6",X"FD",X"17",X"F9",X"DA",X"F3",X"1E",X"EF",X"FA",X"ED",X"7E",X"F7",
		X"F8",X"01",X"32",X"0D",X"48",X"0E",X"4E",X"08",X"C7",X"03",X"58",X"FE",X"A1",X"F9",X"50",X"F4",
		X"95",X"EF",X"C8",X"ED",X"89",X"F6",X"19",X"01",X"68",X"0C",X"98",X"0E",X"AC",X"08",X"21",X"04",
		X"A9",X"FE",X"F2",X"F9",X"9A",X"F4",X"DC",X"EF",X"B1",X"ED",X"FD",X"F5",X"99",X"00",X"F6",X"0B",
		X"C3",X"0E",X"DF",X"08",X"50",X"04",X"D4",X"FE",X"1B",X"FA",X"BC",X"F4",X"FE",X"EF",X"A7",X"ED",
		X"BE",X"F5",X"63",X"00",X"CC",X"0B",X"D5",X"0E",X"F0",X"08",X"5F",X"04",X"E0",X"FE",X"27",X"FA",
		X"C3",X"F4",X"06",X"F0",X"A0",X"ED",X"B5",X"F5",X"5F",X"00",X"D2",X"0B",X"DC",X"0E",X"E5",X"08",
		X"5D",X"04",X"D4",X"FE",X"1F",X"FA",X"B6",X"F4",X"FC",X"EF",X"9C",X"ED",X"D6",X"F5",X"7D",X"00",
		X"03",X"0C",X"DE",X"0E",X"C9",X"08",X"4C",X"04",X"BA",X"FE",X"0B",X"FA",X"98",X"F4",X"E2",X"EF",
		X"94",X"ED",X"14",X"F6",X"B9",X"00",X"56",X"0C",X"E0",X"0E",X"A0",X"08",X"2E",X"04",X"92",X"FE",
		X"EA",X"F9",X"70",X"F4",X"D0",X"EF",X"C6",X"ED",X"64",X"F6",X"14",X"01",X"87",X"0C",X"AD",X"0E",
		X"7A",X"08",X"FE",X"03",X"6C",X"FE",X"B9",X"F9",X"48",X"F4",X"AC",X"EF",X"0D",X"EE",X"C8",X"F6",
		X"81",X"01",X"C0",X"0C",X"6B",X"0E",X"56",X"08",X"C4",X"03",X"42",X"FE",X"7E",X"F9",X"1B",X"F4",
		X"7D",X"EF",X"56",X"EE",X"35",X"F7",X"FA",X"01",X"03",X"0D",X"2D",X"0E",X"2F",X"08",X"A1",X"03",
		X"2D",X"FE",X"7B",X"F9",X"22",X"F4",X"A1",X"EF",X"27",X"EE",X"83",X"F6",X"FC",X"00",X"1F",X"0C",
		X"EE",X"0E",X"F4",X"08",X"9B",X"04",X"36",X"FF",X"AE",X"FA",X"70",X"F5",X"DA",X"F0",X"A2",X"ED",
		X"17",X"F3",X"54",X"FD",X"17",X"08",X"65",X"0F",X"7B",X"0B",X"7A",X"06",X"B7",X"01",X"C9",X"FC",
		X"16",X"F8",X"1A",X"F3",X"D6",X"EE",X"EF",X"EE",X"DA",X"F7",X"05",X"02",X"C2",X"0C",X"A4",X"0E",
		X"CA",X"08",X"75",X"04",X"25",X"FF",X"9E",X"FA",X"6C",X"F5",X"CF",X"F0",X"BD",X"ED",X"3A",X"F3",
		X"94",X"FD",X"75",X"08",X"70",X"0F",X"0D",X"0B",X"25",X"06",X"1A",X"01",X"3F",X"FC",X"38",X"F7",
		X"59",X"F2",X"2D",X"EE",X"43",X"F0",X"83",X"FA",X"1F",X"05",X"E5",X"0E",X"C3",X"0C",X"40",X"07",
		X"86",X"02",X"53",X"FD",X"86",X"F8",X"57",X"F3",X"F5",X"EE",X"1C",X"EF",X"48",X"F8",X"E7",X"02",
		X"83",X"0D",X"E3",X"0D",X"04",X"08",X"7A",X"03",X"13",X"FE",X"65",X"F9",X"0C",X"F4",X"A2",X"EF",
		X"6D",X"EE",X"C8",X"F6",X"75",X"01",X"83",X"0C",X"9B",X"0E",X"87",X"08",X"19",X"04",X"8E",X"FE",
		X"F6",X"F9",X"7C",X"F4",X"17",X"F0",X"0D",X"EE",X"D7",X"F5",X"8C",X"00",X"DA",X"0B",X"FF",X"0E",
		X"E1",X"08",X"75",X"04",X"DF",X"FE",X"47",X"FA",X"C7",X"F4",X"58",X"F0",X"E9",X"ED",X"47",X"F5",
		X"0F",X"00",X"6B",X"0B",X"34",X"0F",X"0E",X"09",X"A8",X"04",X"07",X"FF",X"75",X"FA",X"E6",X"F4",
		X"7D",X"F0",X"E2",X"ED",X"05",X"F5",X"C7",X"FF",X"27",X"0B",X"51",X"0F",X"4F",X"09",X"E5",X"04",
		X"66",X"FF",X"D1",X"FA",X"78",X"F5",X"EA",X"F0",X"E7",X"ED",X"6F",X"F3",X"CD",X"FD",X"CB",X"08",
		X"71",X"0F",X"EC",X"0A",X"1A",X"06",X"19",X"01",X"47",X"FC",X"64",X"F7",X"81",X"F2",X"A0",X"EE",
		X"CE",X"EF",X"51",X"F9",X"95",X"03",X"C4",X"0D",X"F3",X"0D",X"46",X"08",X"F5",X"03",X"B7",X"FE",
		X"44",X"FA",X"16",X"F5",X"B4",X"F0",X"06",X"EE",X"7E",X"F3",X"B7",X"FD",X"7E",X"08",X"6A",X"0F",
		X"34",X"0B",X"4C",X"06",X"5F",X"01",X"7C",X"FC",X"9D",X"F7",X"A6",X"F2",X"BA",X"EE",X"E2",X"EF",
		X"5F",X"F9",X"E2",X"03",X"16",X"0E",X"96",X"0D",X"D4",X"07",X"5C",X"03",X"00",X"FE",X"71",X"F9",
		X"14",X"F4",X"E3",X"EF",X"7A",X"EE",X"1D",X"F6",X"98",X"00",X"AD",X"0B",X"3D",X"0F",X"48",X"09",
		X"FE",X"04",X"9D",X"FF",X"1F",X"FB",X"ED",X"F5",X"55",X"F1",X"2B",X"EE",X"25",X"F2",X"14",X"FC",
		X"BA",X"06",X"48",X"0F",X"69",X"0C",X"03",X"07",X"98",X"02",X"67",X"FD",X"06",X"F9",X"C3",X"F3",
		X"E1",X"EF",X"64",X"EE",X"98",X"F5",X"C2",X"FF",X"76",X"0A",X"6E",X"0F",X"57",X"0A",X"D9",X"05",
		X"DA",X"00",X"2F",X"FC",X"58",X"F7",X"83",X"F2",X"D0",X"EE",X"05",X"F0",X"10",X"F9",X"6B",X"03",
		X"93",X"0D",X"12",X"0E",X"45",X"08",X"F6",X"03",X"A0",X"FE",X"2C",X"FA",X"E5",X"F4",X"92",X"F0",
		X"55",X"EE",X"36",X"F4",X"84",X"FE",X"7D",X"09",X"6B",X"0F",X"8C",X"0A",X"D1",X"05",X"AD",X"00",
		X"E7",X"FB",X"D4",X"F6",X"03",X"F2",X"8A",X"EE",X"1D",X"F1",X"38",X"FB",X"FD",X"05",X"45",X"0F",
		X"62",X"0C",X"F7",X"06",X"38",X"02",X"09",X"FD",X"43",X"F8",X"06",X"F3",X"1D",X"EF",X"D0",X"EF",
		X"D7",X"F8",X"9D",X"03",X"E6",X"0D",X"9F",X"0D",X"C6",X"07",X"40",X"03",X"D3",X"FD",X"34",X"F9",
		X"C3",X"F3",X"B1",X"EF",X"0A",X"EF",X"3B",X"F7",X"0D",X"02",X"E2",X"0C",X"6E",X"0E",X"4F",X"08",
		X"EF",X"03",X"56",X"FE",X"D4",X"F9",X"3C",X"F4",X"2C",X"F0",X"97",X"EE",X"3A",X"F6",X"0B",X"01",
		X"35",X"0C",X"E0",X"0E",X"B1",X"08",X"52",X"04",X"B3",X"FE",X"29",X"FA",X"92",X"F4",X"69",X"F0",
		X"86",X"EE",X"A9",X"F5",X"7A",X"00",X"C4",X"0B",X"1E",X"0F",X"E4",X"08",X"8B",X"04",X"E0",X"FE",
		X"61",X"FA",X"C6",X"F4",X"9C",X"F0",X"7D",X"EE",X"19",X"F5",X"A1",X"FF",X"FE",X"0A",X"7A",X"0F",
		X"97",X"09",X"33",X"05",X"CD",X"FF",X"3B",X"FB",X"FC",X"F5",X"64",X"F1",X"91",X"EE",X"6D",X"F2",
		X"69",X"FC",X"37",X"07",X"52",X"0F",X"0F",X"0C",X"C4",X"06",X"33",X"02",X"0E",X"FD",X"93",X"F8",
		X"4F",X"F3",X"B0",X"EF",X"31",X"EF",X"E6",X"F6",X"13",X"01",X"EA",X"0B",X"53",X"0F",X"81",X"09",
		X"4C",X"05",X"1D",X"00",X"A2",X"FB",X"B1",X"F6",X"0A",X"F2",X"F1",X"EE",X"B9",X"F0",X"C2",X"F9",
		X"FA",X"03",X"C3",X"0D",X"1A",X"0E",X"70",X"08",X"47",X"04",X"1B",X"FF",X"C7",X"FA",X"C2",X"F5",
		X"59",X"F1",X"AF",X"EE",X"A4",X"F1",X"35",X"FB",X"60",X"05",X"84",X"0E",X"78",X"0D",X"F8",X"07",
		X"C8",X"03",X"A0",X"FE",X"55",X"FA",X"34",X"F5",X"03",X"F1",X"A9",X"EE",X"BA",X"F2",X"A8",X"FC",
		X"31",X"07",X"70",X"0F",X"41",X"0C",X"07",X"07",X"86",X"02",X"63",X"FD",X"F0",X"F8",X"A6",X"F3",
		X"01",X"F0",X"2A",X"EF",X"61",X"F6",X"B7",X"00",X"92",X"0B",X"25",X"0F",X"83",X"09",X"23",X"05",
		X"D3",X"FF",X"47",X"FB",X"13",X"F6",X"82",X"F1",X"CC",X"EE",X"52",X"F2",X"62",X"FC",X"49",X"07",
		X"8F",X"0F",X"CD",X"0B",X"A6",X"06",X"CC",X"01",X"BB",X"FC",X"EF",X"F7",X"BF",X"F2",X"65",X"EF",
		X"5B",X"F0",X"49",X"F9",X"26",X"04",X"1E",X"0E",X"8D",X"0D",X"A1",X"07",X"37",X"03",X"B7",X"FD",
		X"39",X"F9",X"A9",X"F3",X"08",X"F0",X"5B",X"EF",X"49",X"F7",X"F1",X"01",X"12",X"0D",X"A7",X"0E",
		X"5F",X"08",X"1B",X"04",X"75",X"FE",X"03",X"FA",X"63",X"F4",X"82",X"F0",X"22",X"EF",X"FA",X"F5",
		X"96",X"00",X"E9",X"0B",X"03",X"0F",X"01",X"09",X"95",X"04",X"06",X"FF",X"73",X"FA",X"E9",X"F4",
		X"C7",X"F0",X"14",X"EF",X"22",X"F5",X"C8",X"FF",X"1B",X"0B",X"36",X"0F",X"62",X"09",X"E3",X"04",
		X"56",X"FF",X"BD",X"FA",X"3A",X"F5",X"FC",X"F0",X"0C",X"EF",X"6D",X"F4",X"EB",X"FE",X"1B",X"0A",
		X"63",X"0F",X"24",X"0A",X"7F",X"05",X"43",X"00",X"8D",X"FB",X"6E",X"F6",X"B1",X"F1",X"16",X"EF",
		X"F9",X"F1",X"B9",X"FB",X"7E",X"06",X"49",X"0F",X"7A",X"0C",X"19",X"07",X"96",X"02",X"64",X"FD",
		X"F5",X"F8",X"9E",X"F3",X"21",X"F0",X"72",X"EF",X"3D",X"F6",X"81",X"00",X"31",X"0B",X"4F",X"0F",
		X"F6",X"09",X"90",X"05",X"85",X"00",X"EA",X"FB",X"1B",X"F7",X"4B",X"F2",X"93",X"EF",X"A0",X"F0",
		X"1D",X"F9",X"54",X"03",X"87",X"0D",X"96",X"0E",X"B0",X"08",X"A6",X"04",X"68",X"FF",X"1C",X"FB",
		X"16",X"F6",X"AC",X"F1",X"55",X"EF",X"9D",X"F1",X"92",X"FA",X"C9",X"04",X"41",X"0E",X"EE",X"0D",
		X"3D",X"08",X"2B",X"04",X"FE",X"FE",X"BE",X"FA",X"BA",X"F5",X"73",X"F1",X"58",X"EF",X"EB",X"F1",
		X"03",X"FB",X"20",X"05",X"7C",X"0E",X"D1",X"0D",X"2C",X"08",X"1D",X"04",X"FA",X"FE",X"BC",X"FA",
		X"BC",X"F5",X"7E",X"F1",X"6D",X"EF",X"D5",X"F1",X"EF",X"FA",X"04",X"05",X"98",X"0E",X"E8",X"0D",
		X"31",X"08",X"31",X"04",X"FF",X"FE",X"CF",X"FA",X"C0",X"F5",X"96",X"F1",X"6F",X"EF",X"BF",X"F1",
		X"D5",X"FA",X"12",X"05",X"90",X"0E",X"D4",X"0D",X"07",X"08",X"09",X"04",X"AA",X"FE",X"86",X"FA",
		X"2C",X"F5",X"45",X"F1",X"57",X"EF",X"2E",X"F3",X"C8",X"FC",X"8F",X"07",X"44",X"0F",X"34",X"0C",
		X"D1",X"06",X"68",X"02",X"1F",X"FD",X"C9",X"F8",X"51",X"F3",X"5E",X"F0",X"D6",X"EF",X"1C",X"F7",
		X"99",X"01",X"52",X"0C",X"F2",X"0E",X"15",X"09",X"C0",X"04",X"60",X"FF",X"DD",X"FA",X"8D",X"F5",
		X"51",X"F1",X"7F",X"EF",X"79",X"F3",X"9F",X"FD",X"A4",X"08",X"7F",X"0F",X"16",X"0B",X"2C",X"06",
		X"1F",X"01",X"36",X"FC",X"3C",X"F7",X"40",X"F2",X"AE",X"EF",X"76",X"F1",X"DA",X"FA",X"D2",X"05",
		X"2E",X"0F",X"AF",X"0C",X"06",X"07",X"6E",X"02",X"15",X"FD",X"7F",X"F8",X"0D",X"F3",X"2E",X"F0",
		X"73",X"F0",X"5F",X"F8",X"22",X"03",X"72",X"0D",X"3D",X"0E",X"55",X"08",X"12",X"04",X"A2",X"FE",
		X"48",X"FA",X"DA",X"F4",X"FE",X"F0",X"99",X"EF",X"38",X"F4",X"37",X"FE",X"0E",X"09",X"81",X"0F",
		X"3C",X"0B",X"59",X"06",X"9C",X"01",X"AB",X"FC",X"21",X"F8",X"F1",X"F2",X"48",X"F0",X"4E",X"F0",
		X"9A",X"F7",X"14",X"02",X"78",X"0C",X"09",X"0F",X"14",X"09",X"F6",X"04",X"8C",X"FF",X"35",X"FB",
		X"E5",X"F5",X"BA",X"F1",X"A7",X"EF",X"76",X"F2",X"46",X"FC",X"1C",X"07",X"6E",X"0F",X"39",X"0C",
		X"D4",X"06",X"44",X"02",X"01",X"FD",X"7D",X"F8",X"11",X"F3",X"63",X"F0",X"6E",X"F0",X"2F",X"F8",
		X"FD",X"02",X"56",X"0D",X"50",X"0E",X"57",X"08",X"0E",X"04",X"94",X"FE",X"37",X"FA",X"B7",X"F4",
		X"FD",X"F0",X"D3",X"EF",X"A5",X"F4",X"D5",X"FE",X"B6",X"09",X"88",X"0F",X"C1",X"0A",X"0F",X"06",
		X"1E",X"01",X"51",X"FC",X"96",X"F7",X"8D",X"F2",X"30",X"F0",X"E8",X"F0",X"BB",X"F8",X"45",X"03",
		X"47",X"0D",X"9B",X"0E",X"AC",X"08",X"A5",X"04",X"47",X"FF",X"0F",X"FB",X"D1",X"F5",X"C7",X"F1",
		X"E1",X"EF",X"52",X"F2",X"54",X"FB",X"D5",X"05",X"B5",X"0E",X"67",X"0D",X"CE",X"07",X"B6",X"03",
		X"6B",X"FE",X"4D",X"FA",X"FC",X"F4",X"6B",X"F1",X"DB",X"EF",X"19",X"F3",X"98",X"FC",X"F9",X"06",
		X"3D",X"0F",X"D0",X"0C",X"82",X"07",X"4B",X"03",X"28",X"FE",X"01",X"FA",X"C2",X"F4",X"4F",X"F1",
		X"EE",X"EF",X"5F",X"F3",X"E8",X"FC",X"47",X"07",X"4C",X"0F",X"99",X"0C",X"54",X"07",X"09",X"03",
		X"D7",X"FD",X"A7",X"F9",X"38",X"F4",X"1C",X"F1",X"F2",X"EF",X"AA",X"F4",X"E0",X"FE",X"90",X"09",
		X"D2",X"0F",X"EF",X"0A",X"3F",X"06",X"57",X"01",X"7D",X"FC",X"C3",X"F7",X"B6",X"F2",X"7A",X"F0",
		X"EE",X"F0",X"FA",X"F8",X"95",X"03",X"01",X"0E",X"52",X"0E",X"28",X"08",X"17",X"04",X"86",X"FE",
		X"56",X"FA",X"BB",X"F4",X"66",X"F1",X"FC",X"EF",X"56",X"F4",X"4D",X"FE",X"38",X"09",X"DC",X"0F",
		X"2F",X"0B",X"67",X"06",X"9D",X"01",X"B7",X"FC",X"27",X"F8",X"03",X"F3",X"A8",X"F0",X"B9",X"F0",
		X"8A",X"F7",X"E2",X"01",X"37",X"0C",X"1B",X"0F",X"83",X"09",X"49",X"05",X"29",X"00",X"B6",X"FB",
		X"CB",X"F6",X"42",X"F2",X"68",X"F0",X"79",X"F1",X"C5",X"F9",X"40",X"04",X"23",X"0E",X"2B",X"0E",
		X"3A",X"08",X"2F",X"04",X"B4",X"FE",X"86",X"FA",X"08",X"F5",X"84",X"F1",X"2D",X"F0",X"FF",X"F3",
		X"C2",X"FD",X"C4",X"08",X"8C",X"0F",X"61",X"0B",X"62",X"06",X"91",X"01",X"8D",X"FC",X"D8",X"F7",
		X"B7",X"F2",X"A4",X"F0",X"4A",X"F1",X"5B",X"F9",X"25",X"04",X"4F",X"0E",X"D8",X"0D",X"DF",X"07",
		X"99",X"03",X"0A",X"FE",X"B6",X"F9",X"01",X"F4",X"31",X"F1",X"50",X"F0",X"39",X"F6",X"1B",X"01",
		X"E2",X"0B",X"25",X"0F",X"1E",X"09",X"D6",X"04",X"3B",X"FF",X"D4",X"FA",X"30",X"F5",X"98",X"F1",
		X"49",X"F0",X"9F",X"F4",X"D8",X"FE",X"43",X"0A",X"D7",X"0F",X"17",X"0A",X"93",X"05",X"1E",X"00",
		X"7E",X"FB",X"10",X"F6",X"CF",X"F1",X"62",X"F0",X"87",X"F3",X"79",X"FD",X"E3",X"08",X"AF",X"0F",
		X"DD",X"0A",X"FE",X"05",X"C0",X"00",X"E3",X"FB",X"A8",X"F6",X"00",X"F2",X"80",X"F0",X"DF",X"F2",
		X"A0",X"FC",X"06",X"08",X"8D",X"0F",X"53",X"0B",X"41",X"06",X"1D",X"01",X"21",X"FC",X"FD",X"F6",
		X"2A",X"F2",X"95",X"F0",X"8C",X"F2",X"26",X"FC",X"8F",X"07",X"78",X"0F",X"94",X"0B",X"60",X"06",
		X"4F",X"01",X"3F",X"FC",X"29",X"F7",X"39",X"F2",X"A6",X"F0",X"70",X"F2",X"F3",X"FB",X"63",X"07",
		X"74",X"0F",X"A8",X"0B",X"6C",X"06",X"5D",X"01",X"47",X"FC",X"33",X"F7",X"3B",X"F2",X"AE",X"F0",
		X"81",X"F2",X"F1",X"FB",X"6C",X"07",X"81",X"0F",X"A3",X"0B",X"66",X"06",X"57",X"01",X"42",X"FC",
		X"35",X"F7",X"46",X"F2",X"C0",X"F0",X"5B",X"F2",X"89",X"FB",X"D0",X"06",X"43",X"0F",X"45",X"0C",
		X"D9",X"06",X"2A",X"02",X"EF",X"FC",X"51",X"F8",X"00",X"F3",X"1C",X"F1",X"3C",X"F1",X"9B",X"F8",
		X"3A",X"03",X"CA",X"0D",X"8E",X"0E",X"66",X"08",X"57",X"04",X"CF",X"FE",X"9D",X"FA",X"14",X"F5",
		X"C9",X"F1",X"A8",X"F0",X"F5",X"F3",X"8D",X"FD",X"76",X"08",X"B8",X"0F",X"A5",X"0B",X"A4",X"06",
		X"E8",X"01",X"DF",X"FC",X"43",X"F8",X"10",X"F3",X"2E",X"F1",X"4B",X"F1",X"5A",X"F8",X"0D",X"03",
		X"8C",X"0D",X"8E",X"0E",X"68",X"08",X"4E",X"04",X"A9",X"FE",X"71",X"FA",X"B5",X"F4",X"B2",X"F1",
		X"B1",X"F0",X"FD",X"F4",X"53",X"FF",X"64",X"0A",X"A0",X"0F",X"2E",X"0A",X"9C",X"05",X"55",X"00",
		X"AB",X"FB",X"79",X"F6",X"2D",X"F2",X"EF",X"F0",X"AF",X"F2",X"D2",X"FB",X"C6",X"06",X"2B",X"0F",
		X"97",X"0C",X"24",X"07",X"AD",X"02",X"6C",X"FD",X"0F",X"F9",X"A0",X"F3",X"7A",X"F1",X"F6",X"F0",
		X"67",X"F6",X"E9",X"00",X"62",X"0B",X"79",X"0F",X"ED",X"09",X"A4",X"05",X"7C",X"00",X"FC",X"FB",
		X"0C",X"F7",X"7E",X"F2",X"23",X"F1",X"DB",X"F1",X"5B",X"F9",X"D8",X"03",X"B8",X"0D",X"88",X"0E",
		X"A5",X"08",X"AD",X"04",X"56",X"FF",X"2C",X"FB",X"F2",X"F5",X"27",X"F2",X"0A",X"F1",X"74",X"F2",
		X"E8",X"FA",X"52",X"05",X"B8",X"0E",X"F1",X"0D",X"21",X"08",X"35",X"04",X"DF",X"FE",X"D1",X"FA",
		X"87",X"F5",X"12",X"F2",X"0B",X"F1",X"C3",X"F2",X"62",X"FB",X"BB",X"05",X"D8",X"0E",X"C2",X"0D",
		X"14",X"08",X"20",X"04",X"D7",X"FE",X"C8",X"FA",X"88",X"F5",X"0F",X"F2",X"19",X"F1",X"D8",X"F2",
		X"4A",X"FB",X"AB",X"05",X"A8",X"0E",X"C6",X"0D",X"24",X"08",X"29",X"04",X"E6",X"FE",X"D3",X"FA",
		X"95",X"F5",X"06",X"F2",X"2C",X"F1",X"D9",X"F2",X"2E",X"FB",X"95",X"05",X"87",X"0E",X"D4",X"0D",
		X"31",X"08",X"34",X"04",X"F3",X"FE",X"DC",X"FA",X"A4",X"F5",X"18",X"F2",X"41",X"F1",X"CB",X"F2",
		X"17",X"FB",X"7A",X"05",X"74",X"0E",X"E3",X"0D",X"3C",X"08",X"3F",X"04",X"03",X"FF",X"E3",X"FA",
		X"B2",X"F5",X"2A",X"F2",X"53",X"F1",X"B2",X"F2",X"02",X"FB",X"5C",X"05",X"71",X"0E",X"F8",X"0D",
		X"44",X"08",X"4B",X"04",X"0E",X"FF",X"EF",X"FA",X"C0",X"F5",X"3A",X"F2",X"5E",X"F1",X"93",X"F2",
		X"E9",X"FA",X"47",X"05",X"79",X"0E",X"0C",X"0E",X"2D",X"08",X"46",X"04",X"D9",X"FE",X"D1",X"FA",
		X"57",X"F5",X"36",X"F2",X"43",X"F1",X"74",X"F3",X"61",X"FC",X"42",X"07",X"2F",X"0F",X"AB",X"0C",
		X"22",X"07",X"DF",X"02",X"79",X"FD",X"48",X"F9",X"B0",X"F3",X"F5",X"F1",X"2F",X"F1",X"71",X"F6",
		X"FE",X"00",X"AF",X"0B",X"52",X"0F",X"A1",X"09",X"44",X"05",X"ED",X"FF",X"6B",X"FB",X"14",X"F6",
		X"50",X"F2",X"70",X"F1",X"41",X"F3",X"A3",X"FC",X"C2",X"07",X"7B",X"0F",X"DD",X"0B",X"AC",X"06",
		X"D8",X"01",X"C0",X"FC",X"F6",X"F7",X"E3",X"F2",X"B2",X"F1",X"1A",X"F2",X"B5",X"F9",X"BF",X"04",
		X"A6",X"0E",X"97",X"0D",X"92",X"07",X"43",X"03",X"AF",X"FD",X"57",X"F9",X"B4",X"F3",X"03",X"F2",
		X"67",X"F1",X"01",X"F7",X"D0",X"01",X"5F",X"0C",X"0C",X"0F",X"26",X"09",X"F2",X"04",X"7C",X"FF",
		X"2B",X"FB",X"B7",X"F5",X"59",X"F2",X"87",X"F1",X"60",X"F3",X"83",X"FC",X"65",X"07",X"4E",X"0F",
		X"7E",X"0C",X"1D",X"07",X"C0",X"02",X"7F",X"FD",X"40",X"F9",X"D5",X"F3",X"14",X"F2",X"77",X"F1",
		X"14",X"F6",X"30",X"00",X"F4",X"0A",X"CA",X"0F",X"3D",X"0A",X"DD",X"05",X"B2",X"00",X"1A",X"FC",
		X"14",X"F7",X"A5",X"F2",X"C6",X"F1",X"80",X"F2",X"51",X"FA",X"2B",X"05",X"E8",X"0E",X"9D",X"0D",
		X"AA",X"07",X"77",X"03",X"E9",X"FD",X"A7",X"F9",X"FD",X"F3",X"27",X"F2",X"8E",X"F1",X"80",X"F6",
		X"08",X"01",X"E0",X"0B",X"4C",X"0F",X"59",X"09",X"0D",X"05",X"83",X"FF",X"1D",X"FB",X"7F",X"F5",
		X"61",X"F2",X"A3",X"F1",X"47",X"F4",X"20",X"FE",X"74",X"09",X"C5",X"0F",X"C0",X"0A",X"04",X"06",
		X"C0",X"00",X"FE",X"FB",X"B6",X"F6",X"9D",X"F2",X"CB",X"F1",X"20",X"F3",X"3E",X"FC",X"8C",X"07",
		X"72",X"0F",X"D4",X"0B",X"93",X"06",X"A2",X"01",X"89",X"FC",X"8C",X"F7",X"C9",X"F2",X"F3",X"F1",
		X"B3",X"F2",X"04",X"FB",X"50",X"06",X"2D",X"0F",X"88",X"0C",X"ED",X"06",X"32",X"02",X"E0",X"FC",
		X"13",X"F8",X"E9",X"F2",X"0F",X"F2",X"74",X"F2",X"48",X"FA",X"8B",X"05",X"F8",X"0E",X"EE",X"0C",
		X"27",X"07",X"80",X"02",X"19",X"FD",X"5A",X"F8",X"10",X"F3",X"1F",X"F2",X"5E",X"F2",X"E0",X"F9",
		X"2A",X"05",X"CC",X"0E",X"34",X"0D",X"4E",X"07",X"CC",X"02",X"51",X"FD",X"C7",X"F8",X"56",X"F3",
		X"47",X"F2",X"08",X"F2",X"70",X"F8",X"4E",X"03",X"CB",X"0D",X"70",X"0E",X"53",X"08",X"32",X"04",
		X"9A",X"FE",X"65",X"FA",X"BB",X"F4",X"6F",X"F2",X"D3",X"F1",X"0C",X"F5",X"AE",X"FE",X"C2",X"09",
		X"F5",X"0F",X"FF",X"0A",X"50",X"06",X"6B",X"01",X"97",X"FC",X"E6",X"F7",X"0A",X"F3",X"4A",X"F2",
		X"28",X"F2",X"46",X"F8",X"D2",X"02",X"F3",X"0C",X"EC",X"0E",X"25",X"09",X"0B",X"05",X"C5",X"FF",
		X"79",X"FB",X"4F",X"F6",X"B8",X"F2",X"2C",X"F2",X"E1",X"F2",X"8D",X"FA",X"00",X"05",X"91",X"0E",
		X"11",X"0E",X"4D",X"08",X"4A",X"04",X"FD",X"FE",X"DD",X"FA",X"91",X"F5",X"9D",X"F2",X"20",X"F2",
		X"58",X"F3",X"A0",X"FB",X"1E",X"06",X"37",X"0F",X"7F",X"0D",X"C7",X"07",X"BB",X"03",X"52",X"FE",
		X"40",X"FA",X"A6",X"F4",X"8D",X"F2",X"FF",X"F1",X"8F",X"F4",X"35",X"FE",X"11",X"09",X"9D",X"0F",
		X"78",X"0B",X"7E",X"06",X"C0",X"01",X"BF",X"FC",X"16",X"F8",X"2E",X"F3",X"85",X"F2",X"2B",X"F2",
		X"AE",X"F8",X"91",X"03",X"9E",X"0D",X"60",X"0E",X"61",X"08",X"30",X"04",X"9D",X"FE",X"5A",X"FA",
		X"A1",X"F4",X"94",X"F2",X"15",X"F2",X"69",X"F5",X"9A",X"FF",X"C6",X"0A",X"B4",X"0F",X"0C",X"0A",
		X"A1",X"05",X"2C",X"00",X"A9",X"FB",X"2C",X"F6",X"D1",X"F2",X"3C",X"F2",X"D8",X"F3",X"EF",X"FC",
		X"38",X"08",X"94",X"0F",X"89",X"0B",X"65",X"06",X"6C",X"01",X"66",X"FC",X"5E",X"F7",X"E8",X"F2",
		X"7A",X"F2",X"0A",X"F3",X"2B",X"FB",X"73",X"06",X"6A",X"0F",X"84",X"0C",X"F0",X"06",X"36",X"02",
		X"ED",X"FC",X"1E",X"F8",X"1D",X"F3",X"9E",X"F2",X"9D",X"F2",X"03",X"FA",X"52",X"05",X"24",X"0F",
		X"27",X"0D",X"46",X"07",X"B9",X"02",X"3E",X"FD",X"99",X"F8",X"51",X"F3",X"B9",X"F2",X"66",X"F2",
		X"55",X"F9",X"A7",X"04",X"BE",X"0E",X"79",X"0D",X"7D",X"07",X"FC",X"02",X"71",X"FD",X"D4",X"F8",
		X"72",X"F3",X"C6",X"F2",X"58",X"F2",X"FE",X"F8",X"53",X"04",X"92",X"0E",X"A7",X"0D",X"92",X"07",
		X"20",X"03",X"82",X"FD",X"F2",X"F8",X"78",X"F3",X"D5",X"F2",X"5C",X"F2",X"ED",X"F8",X"36",X"04",
		X"9B",X"0E",X"B2",X"0D",X"95",X"07",X"21",X"03",X"84",X"FD",X"EE",X"F8",X"76",X"F3",X"D7",X"F2",
		X"6A",X"F2",X"CF",X"F8",X"F9",X"03",X"5D",X"0E",X"F8",X"0D",X"DC",X"07",X"93",X"03",X"FB",X"FD",
		X"9E",X"F9",X"11",X"F4",X"E8",X"F2",X"4F",X"F2",X"C9",X"F6",X"2D",X"01",X"F4",X"0B",X"49",X"0F",
		X"7F",X"09",X"37",X"05",X"D5",X"FF",X"73",X"FB",X"0F",X"F6",X"EE",X"F2",X"A1",X"F2",X"95",X"F3",
		X"E3",X"FB",X"BB",X"06",X"32",X"0F",X"F2",X"0C",X"63",X"07",X"21",X"03",X"D1",X"FD",X"9C",X"F9",
		X"3C",X"F4",X"FC",X"F2",X"66",X"F2",X"AD",X"F5",X"2C",X"FF",X"0E",X"0A",X"BB",X"0F",X"27",X"0B",
		X"65",X"06",X"BE",X"01",X"D8",X"FC",X"64",X"F8",X"7B",X"F3",X"06",X"F3",X"6F",X"F2",X"29",X"F7",
		X"ED",X"00",X"AE",X"0B",X"C3",X"0F",X"42",X"0A",X"F2",X"05",X"0E",X"01",X"71",X"FC",X"CE",X"F7",
		X"43",X"F3",X"09",X"F3",X"8B",X"F2",X"BA",X"F7",X"93",X"01",X"27",X"0C",X"A8",X"0F",X"06",X"0A",
		X"DB",X"05",X"E4",X"00",X"66",X"FC",X"B0",X"F7",X"54",X"F3",X"0A",X"F3",X"A0",X"F2",X"AB",X"F7",
		X"92",X"01",X"00",X"0C",X"8C",X"0F",X"19",X"0A",X"E2",X"05",X"F3",X"00",X"71",X"FC",X"BB",X"F7",
		X"6B",X"F3",X"14",X"F3",X"A9",X"F2",X"8B",X"F7",X"80",X"01",X"D9",X"0B",X"79",X"0F",X"2F",X"0A",
		X"E7",X"05",X"02",X"01",X"77",X"FC",X"CE",X"F7",X"76",X"F3",X"22",X"F3",X"A7",X"F2",X"67",X"F7",
		X"70",X"01",X"B5",X"0B",X"77",X"0F",X"42",X"0A",X"EC",X"05",X"15",X"01",X"7D",X"FC",X"DE",X"F7",
		X"7A",X"F3",X"33",X"F3",X"96",X"F2",X"43",X"F7",X"5B",X"01",X"98",X"0B",X"84",X"0F",X"4F",X"0A",
		X"F7",X"05",X"21",X"01",X"87",X"FC",X"ED",X"F7",X"83",X"F3",X"3E",X"F3",X"A2",X"F2",X"42",X"F7",
		X"3C",X"01",X"8A",X"0B",X"98",X"0F",X"5A",X"0A",X"FF",X"05",X"2D",X"01",X"8F",X"FC",X"FA",X"F7",
		X"86",X"F3",X"45",X"F3",X"B3",X"F2",X"47",X"F7",X"15",X"01",X"8A",X"0B",X"B2",X"0F",X"63",X"0A",
		X"0C",X"06",X"3A",X"01",X"9A",X"FC",X"06",X"F8",X"85",X"F3",X"4E",X"F3",X"BF",X"F2",X"42",X"F7",
		X"EE",X"00",X"91",X"0B",X"D3",X"0F",X"65",X"0A",X"1A",X"06",X"42",X"01",X"A8",X"FC",X"0E",X"F8",
		X"85",X"F3",X"54",X"F3",X"D1",X"F2",X"27",X"F7",X"DB",X"00",X"6B",X"0B",X"AE",X"0F",X"7C",X"0A",
		X"1F",X"06",X"50",X"01",X"B0",X"FC",X"1A",X"F8",X"9B",X"F3",X"62",X"F3",X"D6",X"F2",X"07",X"F7",
		X"C9",X"00",X"46",X"0B",X"98",X"0F",X"94",X"0A",X"23",X"06",X"60",X"01",X"B8",X"FC",X"29",X"F8",
		X"AB",X"F3",X"71",X"F3",X"D4",X"F2",X"E2",X"F6",X"BA",X"00",X"20",X"0B",X"94",X"0F",X"A4",X"0A",
		X"2F",X"06",X"6E",X"01",X"C2",X"FC",X"34",X"F8",X"BB",X"F3",X"7B",X"F3",X"D2",X"F2",X"B6",X"F6",
		X"AF",X"00",X"FB",X"0A",X"A6",X"0F",X"A7",X"0A",X"3F",X"06",X"6F",X"01",X"D1",X"FC",X"2A",X"F8",
		X"C6",X"F3",X"7B",X"F3",X"E5",X"F2",X"20",X"F7",X"66",X"01",X"BD",X"0B",X"70",X"0F",X"E3",X"09",
		X"A7",X"05",X"6E",X"00",X"04",X"FC",X"CE",X"F6",X"5D",X"F3",X"6A",X"F3",X"77",X"F3",X"4E",X"FA",
		X"1C",X"05",X"9A",X"0E",X"C8",X"0D",X"E0",X"07",X"BA",X"03",X"45",X"FE",X"0C",X"FA",X"9D",X"F4",
		X"85",X"F3",X"0F",X"F3",X"85",X"F5",X"B9",X"FE",X"CB",X"09",X"F7",X"0F",X"28",X"0B",X"71",X"06",
		X"A6",X"01",X"D4",X"FC",X"2B",X"F8",X"C0",X"F3",X"9F",X"F3",X"00",X"F3",X"9C",X"F7",X"B8",X"01",
		X"1D",X"0C",X"53",X"0F",X"D4",X"09",X"8D",X"05",X"84",X"00",X"09",X"FC",X"20",X"F7",X"7E",X"F3",
		X"AC",X"F3",X"14",X"F3",X"CD",X"F8",X"35",X"03",X"21",X"0D",X"E4",X"0E",X"44",X"09",X"25",X"05",
		X"0D",X"00",X"B5",X"FB",X"B9",X"F6",X"76",X"F3",X"B0",X"F3",X"2F",X"F3",X"3A",X"F9",X"92",X"03",
		X"58",X"0D",X"D1",X"0E",X"2E",X"09",X"17",X"05",X"03",X"00",X"B2",X"FB",X"BB",X"F6",X"88",X"F3",
		X"B2",X"F3",X"49",X"F3",X"3C",X"F9",X"6F",X"03",X"4E",X"0D",X"E3",X"0E",X"36",X"09",X"23",X"05",
		X"0F",X"00",X"BD",X"FB",X"C7",X"F6",X"93",X"F3",X"B9",X"F3",X"5C",X"F3",X"33",X"F9",X"4C",X"03",
		X"51",X"0D",X"FA",X"0E",X"3E",X"09",X"32",X"05",X"19",X"00",X"C8",X"FB",X"D2",X"F6",X"9A",X"F3",
		X"C0",X"F3",X"6A",X"F3",X"1F",X"F9",X"2C",X"03",X"62",X"0D",X"1B",X"0F",X"3B",X"09",X"48",X"05",
		X"19",X"00",X"DE",X"FB",X"CF",X"F6",X"A7",X"F3",X"BD",X"F3",X"84",X"F3",X"50",X"F9",X"AC",X"03",
		X"C1",X"0D",X"C8",X"0E",X"B7",X"08",X"C7",X"04",X"53",X"FF",X"29",X"FB",X"BF",X"F5",X"B7",X"F3",
		X"93",X"F3",X"31",X"F4",X"24",X"FC",X"42",X"07",X"4B",X"0F",X"94",X"0C",X"22",X"07",X"AF",X"02",
		X"72",X"FD",X"F3",X"F8",X"1C",X"F4",X"F2",X"F3",X"3C",X"F3",X"33",X"F7",X"4A",X"01",X"00",X"0C",
		X"43",X"0F",X"B8",X"09",X"63",X"05",X"32",X"00",X"BE",X"FB",X"9A",X"F6",X"AA",X"F3",X"D7",X"F3",
		X"CB",X"F3",X"67",X"FA",X"FB",X"04",X"85",X"0E",X"0A",X"0E",X"2F",X"08",X"27",X"04",X"CF",X"FE",
		X"A7",X"FA",X"5C",X"F5",X"D1",X"F3",X"A5",X"F3",X"77",X"F4",X"4C",X"FC",X"09",X"07",X"24",X"0F",
		X"0C",X"0D",X"91",X"07",X"6D",X"03",X"36",X"FE",X"0C",X"FA",X"E4",X"F4",X"E3",X"F3",X"98",X"F3",
		X"D9",X"F4",X"20",X"FD",X"C7",X"07",X"5B",X"0F",X"AF",X"0C",X"64",X"07",X"31",X"03",X"16",X"FE",
		X"E4",X"F9",X"DA",X"F4",X"EB",X"F3",X"A2",X"F3",X"F4",X"F4",X"2A",X"FD",X"BE",X"07",X"6D",X"0F",
		X"B7",X"0C",X"6B",X"07",X"3B",X"03",X"20",X"FE",X"ED",X"F9",X"EA",X"F4",X"F4",X"F3",X"AE",X"F3",
		X"F9",X"F4",X"0C",X"FD",X"A7",X"07",X"84",X"0F",X"C7",X"0C",X"75",X"07",X"47",X"03",X"2B",X"FE",
		X"F9",X"F9",X"F7",X"F4",X"F8",X"F3",X"BA",X"F3",X"F5",X"F4",X"ED",X"FC",X"95",X"07",X"A8",X"0F",
		X"D0",X"0C",X"7F",X"07",X"52",X"03",X"34",X"FE",X"03",X"FA",X"02",X"F5",X"FD",X"F3",X"CB",X"F3",
		X"E1",X"F4",X"CF",X"FC",X"80",X"07",X"72",X"0F",X"DA",X"0C",X"8B",X"07",X"5B",X"03",X"41",X"FE",
		X"0D",X"FA",X"0A",X"F5",X"FE",X"F3",X"DC",X"F3",X"BF",X"F4",X"B6",X"FC",X"68",X"07",X"4A",X"0F",
		X"E6",X"0C",X"96",X"07",X"66",X"03",X"4B",X"FE",X"19",X"FA",X"0D",X"F5",X"02",X"F4",X"E8",X"F3",
		X"A4",X"F4",X"A4",X"FC",X"4A",X"07",X"32",X"0F",X"F8",X"0C",X"99",X"07",X"6C",X"03",X"3F",X"FE",
		X"08",X"FA",X"E9",X"F4",X"1B",X"F4",X"D6",X"F3",X"0D",X"F5",X"A3",X"FD",X"AD",X"08",X"9D",X"0F",
		X"E1",X"0B",X"CB",X"06",X"35",X"02",X"2D",X"FD",X"90",X"F8",X"30",X"F4",X"5B",X"F4",X"A0",X"F3",
		X"C2",X"F7",X"D3",X"01",X"90",X"0C",X"F7",X"0E",X"48",X"09",X"E5",X"04",X"97",X"FF",X"14",X"FB",
		X"D3",X"F5",X"11",X"F4",X"0C",X"F4",X"DA",X"F4",X"33",X"FD",X"7C",X"08",X"A6",X"0F",X"7F",X"0B",
		X"83",X"06",X"84",X"01",X"A3",X"FC",X"88",X"F7",X"F0",X"F3",X"65",X"F4",X"E4",X"F3",X"1E",X"FA",
		X"46",X"05",X"CF",X"0E",X"51",X"0D",X"75",X"07",X"FC",X"02",X"93",X"FD",X"EA",X"F8",X"4A",X"F4",
		X"7B",X"F4",X"AF",X"F3",X"61",X"F8",X"FD",X"02",X"CC",X"0D",X"4A",X"0E",X"41",X"08",X"D6",X"03",
		X"55",X"FE",X"BA",X"F9",X"AD",X"F4",X"67",X"F4",X"D2",X"F3",X"51",X"F7",X"92",X"01",X"B2",X"0C",
		X"C7",X"0E",X"D3",X"08",X"5D",X"04",X"D4",X"FE",X"3A",X"FA",X"F6",X"F4",X"5B",X"F4",X"EB",X"F3",
		X"B4",X"F6",X"B0",X"00",X"04",X"0C",X"09",X"0F",X"2E",X"09",X"A9",X"04",X"21",X"FF",X"81",X"FA",
		X"28",X"F5",X"58",X"F4",X"00",X"F4",X"63",X"F6",X"38",X"00",X"A5",X"0B",X"29",X"0F",X"5A",X"09",
		X"CE",X"04",X"46",X"FF",X"A1",X"FA",X"43",X"F5",X"5D",X"F4",X"0A",X"F4",X"4B",X"F6",X"09",X"00",
		X"88",X"0B",X"30",X"0F",X"6A",X"09",X"D5",X"04",X"50",X"FF",X"A3",X"FA",X"4C",X"F5",X"66",X"F4",
		X"14",X"F4",X"56",X"F6",X"11",X"00",X"99",X"0B",X"2D",X"0F",X"5C",X"09",X"CB",X"04",X"3E",X"FF",
		X"94",X"FA",X"44",X"F5",X"74",X"F4",X"12",X"F4",X"7D",X"F6",X"3E",X"00",X"D3",X"0B",X"23",X"0F",
		X"3B",X"09",X"B2",X"04",X"1F",X"FF",X"76",X"FA",X"2F",X"F5",X"88",X"F4",X"0C",X"F4",X"AF",X"F6",
		X"86",X"00",X"1D",X"0C",X"1F",X"0F",X"22",X"09",X"AD",X"04",X"26",X"FF",X"8D",X"FA",X"55",X"F5",
		X"81",X"F4",X"2F",X"F4",X"0B",X"F6",X"2B",X"FF",X"8E",X"0A",X"76",X"0F",X"50",X"0A",X"A7",X"05",
		X"7B",X"00",X"D0",X"FB",X"9E",X"F6",X"43",X"F4",X"9D",X"F4",X"6F",X"F4",X"23",X"FB",X"18",X"06",
		X"F5",X"0E",X"15",X"0D",X"8E",X"07",X"28",X"03",X"FA",X"FD",X"7B",X"F9",X"CC",X"F4",X"AE",X"F4",
		X"28",X"F4",X"59",X"F6",X"33",X"FF",X"3B",X"0A",X"93",X"0F",X"F6",X"0A",X"2D",X"06",X"76",X"01",
		X"A2",X"FC",X"F7",X"F7",X"51",X"F4",X"DF",X"F4",X"FE",X"F3",X"ED",X"F7",X"AE",X"01",X"4A",X"0C",
		X"29",X"0F",X"D5",X"09",X"71",X"05",X"8C",X"00",X"F5",X"FB",X"31",X"F7",X"49",X"F4",X"E8",X"F4",
		X"05",X"F4",X"C0",X"F8",X"D6",X"02",X"14",X"0D",X"E6",X"0E",X"66",X"09",X"2B",X"05",X"34",X"00",
		X"C0",X"FB",X"EE",X"F6",X"59",X"F4",X"E2",X"F4",X"21",X"F4",X"F5",X"F8",X"04",X"03",X"15",X"0D",
		X"E0",X"0E",X"60",X"09",X"31",X"05",X"31",X"00",X"CC",X"FB",X"EE",X"F6",X"66",X"F4",X"E1",X"F4",
		X"3A",X"F4",X"EE",X"F8",X"EC",X"02",X"F3",X"0C",X"F0",X"0E",X"65",X"09",X"3D",X"05",X"2A",X"00",
		X"CC",X"FB",X"D3",X"F6",X"72",X"F4",X"E0",X"F4",X"57",X"F4",X"91",X"F9",X"02",X"04",X"D6",X"0D",
		X"4D",X"0E",X"8A",X"08",X"5C",X"04",X"0F",X"FF",X"AE",X"FA",X"9D",X"F5",X"B1",X"F4",X"9B",X"F4",
		X"55",X"F5",X"01",X"FD",X"3F",X"08",X"71",X"0F",X"E3",X"0B",X"AA",X"06",X"FE",X"01",X"F4",X"FC",
		X"2F",X"F8",X"83",X"F4",X"0B",X"F5",X"45",X"F4",X"65",X"F8",X"6D",X"02",X"05",X"0D",X"C3",X"0E",
		X"16",X"09",X"BC",X"04",X"97",X"FF",X"10",X"FB",X"28",X"F6",X"96",X"F4",X"E5",X"F4",X"A2",X"F4",
		X"71",X"FB",X"55",X"06",X"2F",X"0F",X"2B",X"0D",X"AB",X"07",X"66",X"03",X"45",X"FE",X"DC",X"F9",
		X"26",X"F5",X"DE",X"F4",X"9D",X"F4",X"B2",X"F5",X"98",X"FD",X"9E",X"08",X"8D",X"0F",X"E6",X"0B",
		X"C1",X"06",X"3B",X"02",X"30",X"FD",X"98",X"F8",X"A8",X"F4",X"2B",X"F5",X"46",X"F4",X"93",X"F7",
		X"51",X"01",X"76",X"0C",X"3C",X"0F",X"63",X"09",X"0E",X"05",X"C9",X"FF",X"36",X"FB",X"2A",X"F6",
		X"B7",X"F4",X"EB",X"F4",X"F5",X"F4",X"70",X"FC",X"D1",X"07",X"AA",X"0F",X"E8",X"0B",X"AE",X"06",
		X"E2",X"01",X"DA",X"FC",X"E8",X"F7",X"A3",X"F4",X"2B",X"F5",X"7F",X"F4",X"76",X"F9",X"4B",X"04",
		X"3F",X"0E",X"A5",X"0D",X"D3",X"07",X"54",X"03",X"F7",X"FD",X"42",X"F9",X"D5",X"F4",X"36",X"F5",
		X"68",X"F4",X"AB",X"F7",X"DA",X"01",X"FD",X"0C",X"C1",X"0E",X"A8",X"08",X"41",X"04",X"C5",X"FE",
		X"1F",X"FA",X"2A",X"F5",X"1E",X"F5",X"99",X"F4",X"BD",X"F6",X"E3",X"FF",X"6E",X"0B",X"55",X"0F",
		X"C2",X"09",X"3C",X"05",X"FB",X"FF",X"55",X"FB",X"4B",X"F6",X"D5",X"F4",X"0C",X"F5",X"03",X"F5",
		X"06",X"FC",X"44",X"07",X"9B",X"0F",X"68",X"0C",X"06",X"07",X"8A",X"02",X"6B",X"FD",X"D4",X"F8",
		X"D8",X"F4",X"51",X"F5",X"86",X"F4",X"4B",X"F7",X"70",X"00",X"87",X"0B",X"4E",X"0F",X"29",X"0A",
		X"99",X"05",X"B6",X"00",X"07",X"FC",X"33",X"F7",X"A6",X"F4",X"66",X"F5",X"87",X"F4",X"1F",X"F9",
		X"1F",X"03",X"8D",X"0D",X"BA",X"0E",X"FE",X"08",X"CB",X"04",X"BB",X"FF",X"49",X"FB",X"74",X"F6",
		X"CE",X"F4",X"4B",X"F5",X"CB",X"F4",X"30",X"FA",X"70",X"04",X"26",X"0E",X"3B",X"0E",X"8D",X"08",
		X"6D",X"04",X"52",X"FF",X"F4",X"FA",X"1E",X"F6",X"F4",X"F4",X"31",X"F5",X"13",X"F5",X"21",X"FB",
		X"E1",X"05",X"BA",X"0E",X"5A",X"0D",X"BA",X"07",X"73",X"03",X"3F",X"FE",X"BD",X"F9",X"45",X"F5",
		X"4F",X"F5",X"D9",X"F4",X"22",X"F6",X"B1",X"FE",X"1D",X"0A",X"A8",X"0F",X"BF",X"0A",X"EF",X"05",
		X"01",X"01",X"24",X"FC",X"3C",X"F7",X"D5",X"F4",X"7A",X"F5",X"B3",X"F4",X"15",X"FA",X"F1",X"04",
		X"90",X"0E",X"96",X"0D",X"D0",X"07",X"80",X"03",X"40",X"FE",X"B6",X"F9",X"4B",X"F5",X"62",X"F5",
		X"E6",X"F4",X"38",X"F6",X"83",X"FE",X"DC",X"09",X"C6",X"0F",X"12",X"0B",X"48",X"06",X"88",X"01",
		X"B9",X"FC",X"FE",X"F7",X"E8",X"F4",X"8A",X"F5",X"C2",X"F4",X"0D",X"F8",X"6E",X"01",X"2B",X"0C",
		X"17",X"0F",X"D1",X"09",X"58",X"05",X"7D",X"00",X"D9",X"FB",X"26",X"F7",X"EE",X"F4",X"8F",X"F5",
		X"CD",X"F4",X"20",X"F9",X"E3",X"02",X"27",X"0D",X"AA",X"0E",X"46",X"09",X"EC",X"04",X"0D",X"00",
		X"7D",X"FB",X"D7",X"F6",X"FC",X"F4",X"91",X"F5",X"DF",X"F4",X"73",X"F9",X"43",X"03",X"56",X"0D",
		X"97",X"0E",X"2F",X"09",X"E0",X"04",X"03",X"00",X"79",X"FB",X"DA",X"F6",X"04",X"F5",X"99",X"F5",
		X"E8",X"F4",X"5B",X"F9",X"25",X"03",X"4C",X"0D",X"AC",X"0E",X"35",X"09",X"EE",X"04",X"0D",X"00",
		X"83",X"FB",X"E4",X"F6",X"06",X"F5",X"A6",X"F5",X"E6",X"F4",X"41",X"F9",X"07",X"03",X"4F",X"0D",
		X"C8",X"0E",X"39",X"09",X"FB",X"04",X"14",X"00",X"8F",X"FB",X"EB",X"F6",X"07",X"F5",X"B4",X"F5",
		X"DB",X"F4",X"1D",X"F9",X"E8",X"02",X"5F",X"0D",X"E7",X"0E",X"37",X"09",X"0F",X"05",X"15",X"00",
		X"A0",X"FB",X"E5",X"F6",X"10",X"F5",X"BB",X"F5",X"E2",X"F4",X"00",X"F9",X"DC",X"02",X"2E",X"0D",
		X"D9",X"0E",X"45",X"09",X"19",X"05",X"1D",X"00",X"B0",X"FB",X"E0",X"F6",X"1B",X"F5",X"BD",X"F5",
		X"F8",X"F4",X"03",X"F9",X"C3",X"02",X"04",X"0D",X"CF",X"0E",X"57",X"09",X"1F",X"05",X"29",X"00",
		X"B7",X"FB",X"E8",X"F6",X"2D",X"F5",X"BC",X"F5",X"0A",X"F5",X"5B",X"F9",X"6E",X"03",X"A0",X"0D",
		X"66",X"0E",X"B7",X"08",X"76",X"04",X"4F",X"FF",X"C5",X"FA",X"1E",X"F6",X"69",X"F5",X"89",X"F5",
		X"9D",X"F5",X"27",X"FC",X"5D",X"07",X"2D",X"0F",X"45",X"0C",X"EC",X"06",X"57",X"02",X"4B",X"FD",
		X"8D",X"F8",X"2F",X"F5",X"D8",X"F5",X"16",X"F5",X"A9",X"F7",X"FD",X"00",X"FB",X"0B",X"19",X"0F",
		X"B0",X"09",X"34",X"05",X"37",X"00",X"8E",X"FB",X"CC",X"F6",X"49",X"F5",X"CD",X"F5",X"2E",X"F5",
		X"1B",X"FA",X"6B",X"04",X"3A",X"0E",X"ED",X"0D",X"5B",X"08",X"11",X"04",X"0B",X"FF",X"7E",X"FA",
		X"16",X"F6",X"78",X"F5",X"B7",X"F5",X"62",X"F5",X"7E",X"FB",X"39",X"06",X"2A",X"0F",X"3B",X"0D",
		X"C1",X"07",X"80",X"03",X"84",X"FE",X"03",X"FA",X"DC",X"F5",X"98",X"F5",X"A7",X"F5",X"95",X"F5",
		X"0C",X"FC",X"D5",X"06",X"4C",X"0F",X"FC",X"0C",X"9D",X"07",X"61",X"03",X"6B",X"FE",X"F3",X"F9",
		X"D0",X"F5",X"AC",X"F5",X"A3",X"F5",X"B6",X"F5",X"08",X"FC",X"CA",X"06",X"17",X"0F",X"FC",X"0C",
		X"99",X"07",X"5B",X"03",X"4C",X"FE",X"D4",X"F9",X"B1",X"F5",X"C9",X"F5",X"8B",X"F5",X"03",X"F6",
		X"25",X"FD",X"74",X"08",X"89",X"0F",X"DD",X"0B",X"A0",X"06",X"20",X"02",X"0D",X"FD",X"68",X"F8",
		X"4E",X"F5",X"17",X"F6",X"2E",X"F5",X"2F",X"F8",X"6C",X"01",X"BC",X"0C",X"D5",X"0E",X"28",X"09",
		X"A5",X"04",X"85",X"FF",X"BB",X"FA",X"35",X"F6",X"AE",X"F5",X"BC",X"F5",X"EF",X"F5",X"03",X"FD",
		X"82",X"08",X"9D",X"0F",X"51",X"0B",X"3F",X"06",X"55",X"01",X"5C",X"FC",X"72",X"F7",X"68",X"F5",
		X"0C",X"F6",X"5E",X"F5",X"39",X"FA",X"4F",X"05",X"A8",X"0E",X"ED",X"0C",X"4A",X"07",X"A4",X"02",
		X"68",X"FD",X"87",X"F8",X"6A",X"F5",X"24",X"F6",X"45",X"F5",X"B3",X"F8",X"C5",X"02",X"97",X"0D",
		X"2F",X"0E",X"4C",X"08",X"D7",X"03",X"96",X"FE",X"DA",X"F9",X"C4",X"F5",X"F8",X"F5",X"9C",X"F5",
		X"8E",X"F6",X"95",X"FE",X"19",X"0A",X"4F",X"0F",X"B8",X"0A",X"CB",X"05",X"0A",X"01",X"1A",X"FC",
		X"78",X"F7",X"6D",X"F5",X"3B",X"F6",X"47",X"F5",X"44",X"F9",X"43",X"03",X"BA",X"0D",X"54",X"0E",
		X"A0",X"08",X"4C",X"04",X"47",X"FF",X"9F",X"FA",X"53",X"F6",X"C8",X"F5",X"F9",X"F5",X"C5",X"F5",
		X"65",X"FB",X"1B",X"06",X"C2",X"0E",X"17",X"0D",X"B4",X"07",X"56",X"03",X"6B",X"FE",X"C5",X"F9",
		X"DC",X"F5",X"F9",X"F5",X"D9",X"F5",X"25",X"F6",X"8E",X"FC",X"68",X"07",X"1E",X"0F",X"86",X"0C",
		X"52",X"07",X"F0",X"02",X"0F",X"FE",X"70",X"F9",X"C0",X"F5",X"16",X"F6",X"C4",X"F5",X"73",X"F6",
		X"56",X"FD",X"87",X"08",X"53",X"0F",X"CB",X"0B",X"AB",X"06",X"22",X"02",X"23",X"FD",X"80",X"F8",
		X"98",X"F5",X"49",X"F6",X"88",X"F5",X"B2",X"F7",X"D1",X"00",X"FC",X"0B",X"E8",X"0E",X"8D",X"09",
		X"E6",X"04",X"EC",X"FF",X"0A",X"FB",X"A4",X"F6",X"D0",X"F5",X"27",X"F6",X"CA",X"F5",X"DE",X"FB",
		X"48",X"07",X"21",X"0F",X"07",X"0C",X"AD",X"06",X"F7",X"01",X"DD",X"FC",X"0D",X"F8",X"AA",X"F5",
		X"54",X"F6",X"93",X"F5",X"43",X"F9",X"7C",X"03",X"20",X"0E",X"BC",X"0D",X"EA",X"07",X"60",X"03",
		X"18",X"FE",X"40",X"F9",X"B6",X"F5",X"56",X"F6",X"A6",X"F5",X"8D",X"F7",X"03",X"01",X"68",X"0C",
		X"8F",X"0E",X"EA",X"08",X"38",X"04",X"03",X"FF",X"07",X"FA",X"00",X"F6",X"3A",X"F6",X"D6",X"F5",
		X"04",X"F7",X"69",X"FF",X"2D",X"0B",X"15",X"0F",X"8D",X"09",X"CB",X"04",X"90",X"FF",X"95",X"FA",
		X"45",X"F6",X"2B",X"F6",X"F5",X"F5",X"B9",X"F6",X"6D",X"FE",X"62",X"0A",X"57",X"0F",X"F6",X"09",
		X"1C",X"05",X"EA",X"FF",X"E5",X"FA",X"74",X"F6",X"22",X"F6",X"0C",X"F6",X"8F",X"F6",X"E6",X"FD",
		X"E9",X"09",X"71",X"0F",X"2D",X"0A",X"46",X"05",X"15",X"00",X"09",X"FB",X"8D",X"F6",X"22",X"F6",
		X"1A",X"F6",X"81",X"F6",X"B3",X"FD",X"B3",X"09",X"6E",X"0F",X"43",X"0A",X"50",X"05",X"24",X"00",
		X"0F",X"FB",X"91",X"F6",X"27",X"F6",X"22",X"F6",X"81",X"F6",X"B8",X"FD",X"B6",X"09",X"5A",X"0F",
		X"40",X"0A",X"43",X"05",X"1A",X"00",X"FD",X"FA",X"89",X"F6",X"30",X"F6",X"28",X"F6",X"8B",X"F6",
		X"E6",X"FD",X"DF",X"09",X"42",X"0F",X"23",X"0A",X"27",X"05",X"FA",X"FF",X"DE",X"FA",X"6E",X"F6",
		X"3E",X"F6",X"29",X"F6",X"98",X"F6",X"2D",X"FE",X"2E",X"0A",X"22",X"0F",X"FA",X"09",X"FD",X"04",
		X"D2",X"FF",X"B3",X"FA",X"5D",X"F6",X"49",X"F6",X"2C",X"F6",X"A5",X"F6",X"8A",X"FE",X"96",X"0A",
		X"09",X"0F",X"C0",X"09",X"D2",X"04",X"9C",X"FF",X"83",X"FA",X"5A",X"F6",X"58",X"F6",X"2A",X"F6",
		X"C6",X"F6",X"EF",X"FE",X"12",X"0B",X"F4",X"0E",X"7F",X"09",X"9F",X"04",X"5F",X"FF",X"4D",X"FA",
		X"4D",X"F6",X"6E",X"F6",X"1F",X"F6",X"1F",X"F7",X"6E",X"FF",X"97",X"0B",X"E9",X"0E",X"31",X"09",
		X"6E",X"04",X"25",X"FF",X"22",X"FA",X"47",X"F6",X"7A",X"F6",X"25",X"F6",X"15",X"F7",X"0D",X"FF",
		X"04",X"0B",X"0B",X"0F",X"C8",X"09",X"FD",X"04",X"F1",X"FF",X"FC",X"FA",X"AE",X"F6",X"46",X"F6",
		X"6F",X"F6",X"49",X"F6",X"0F",X"FC",X"56",X"07",X"5F",X"0F",X"FE",X"0B",X"AC",X"06",X"18",X"02",
		X"07",X"FD",X"63",X"F8",X"F5",X"F5",X"BA",X"F6",X"F2",X"F5",X"34",X"F8",X"C9",X"00",X"2C",X"0C",
		X"EB",X"0E",X"8E",X"09",X"FC",X"04",X"26",X"00",X"4C",X"FB",X"0D",X"F7",X"2A",X"F6",X"B0",X"F6",
		X"F2",X"F5",X"DA",X"F9",X"19",X"04",X"E5",X"0D",X"DB",X"0D",X"56",X"08",X"F6",X"03",X"14",X"FF",
		X"5A",X"FA",X"91",X"F6",X"5F",X"F6",X"8F",X"F6",X"3A",X"F6",X"25",X"FB",X"B3",X"05",X"8B",X"0E",
		X"2D",X"0D",X"D6",X"07",X"74",X"03",X"A3",X"FE",X"EE",X"F9",X"78",X"F6",X"71",X"F6",X"8E",X"F6",
		X"51",X"F6",X"8D",X"FB",X"24",X"06",X"AE",X"0E",X"08",X"0D",X"BF",X"07",X"60",X"03",X"97",X"FE",
		X"E0",X"F9",X"77",X"F6",X"77",X"F6",X"9A",X"F6",X"41",X"F6",X"6E",X"FB",X"0D",X"06",X"AC",X"0E",
		X"1D",X"0D",X"C2",X"07",X"6E",X"03",X"9F",X"FE",X"E8",X"F9",X"70",X"F6",X"82",X"F6",X"9F",X"F6",
		X"40",X"F6",X"5B",X"FB",X"F1",X"05",X"BC",X"0E",X"33",X"0D",X"C2",X"07",X"7D",X"03",X"A1",X"FE",
		X"FA",X"F9",X"7E",X"F6",X"90",X"F6",X"9F",X"F6",X"58",X"F6",X"55",X"FB",X"CF",X"05",X"E0",X"0E",
		X"42",X"0D",X"C7",X"07",X"8C",X"03",X"A4",X"FE",X"0C",X"FA",X"89",X"F6",X"9D",X"F6",X"9B",X"F6",
		X"71",X"F6",X"3E",X"FB",X"C1",X"05",X"AA",X"0E",X"40",X"0D",X"C0",X"07",X"83",X"03",X"81",X"FE",
		X"E5",X"F9",X"72",X"F6",X"BB",X"F6",X"87",X"F6",X"AA",X"F6",X"60",X"FC",X"A7",X"07",X"27",X"0F",
		X"11",X"0C",X"A7",X"06",X"41",X"02",X"14",X"FD",X"97",X"F8",X"30",X"F6",X"FE",X"F6",X"32",X"F6",
		X"41",X"F8",X"9F",X"00",X"52",X"0C",X"DE",X"0E",X"36",X"09",X"9D",X"04",X"97",X"FF",X"A5",X"FA",
		X"CD",X"F6",X"A2",X"F6",X"B2",X"F6",X"A0",X"F6",X"81",X"FC",X"01",X"08",X"38",X"0F",X"67",X"0B",
		X"20",X"06",X"61",X"01",X"35",X"FC",X"B0",X"F7",X"62",X"F6",X"F6",X"F6",X"41",X"F6",X"F5",X"F9",
		X"D0",X"04",X"7C",X"0E",X"DB",X"0C",X"39",X"07",X"90",X"02",X"54",X"FD",X"8F",X"F8",X"54",X"F6",
		X"03",X"F7",X"49",X"F6",X"D3",X"F8",X"90",X"02",X"6C",X"0D",X"C4",X"0D",X"FF",X"07",X"52",X"03",
		X"16",X"FE",X"23",X"F9",X"59",X"F6",X"05",X"F7",X"62",X"F6",X"3B",X"F8",X"19",X"01",X"AD",X"0C",
		X"4F",X"0E",X"7F",X"08",X"CC",X"03",X"90",X"FE",X"82",X"F9",X"62",X"F6",X"08",X"F7",X"73",X"F6",
		X"EA",X"F7",X"2E",X"00",X"20",X"0C",X"A9",X"0E",X"EE",X"08",X"36",X"04",X"1A",X"FF",X"08",X"FA",
		X"A4",X"F6",X"E0",X"F6",X"B7",X"F6",X"F2",X"F6",X"CE",X"FD",X"B0",X"09",X"14",X"0F",X"98",X"0A",
		X"92",X"05",X"CE",X"00",X"C0",X"FB",X"73",X"F7",X"8D",X"F6",X"0F",X"F7",X"68",X"F6",X"C2",X"F9",
		X"0B",X"04",X"F0",X"0D",X"85",X"0D",X"FD",X"07",X"86",X"03",X"8B",X"FE",X"BD",X"F9",X"9B",X"F6",
		X"F6",X"F6",X"C4",X"F6",X"E7",X"F6",X"AF",X"FC",X"E7",X"07",X"2C",X"0F",X"E5",X"0B",X"A2",X"06",
		X"3B",X"02",X"39",X"FD",X"BC",X"F8",X"7D",X"F6",X"1C",X"F7",X"A1",X"F6",X"61",X"F7",X"7A",X"FE",
		X"DE",X"09",X"11",X"0F",X"FD",X"0A",X"FC",X"05",X"8E",X"01",X"99",X"FC",X"4F",X"F8",X"86",X"F6",
		X"2A",X"F7",X"98",X"F6",X"BF",X"F7",X"4D",X"FF",X"89",X"0A",X"07",X"0F",X"AB",X"0A",X"CD",X"05",
		X"58",X"01",X"73",X"FC",X"34",X"F8",X"8F",X"F6",X"2F",X"F7",X"9F",X"F6",X"B3",X"F7",X"53",X"FF",
		X"7F",X"0A",X"15",X"0F",X"AC",X"0A",X"D5",X"05",X"61",X"01",X"7E",X"FC",X"39",X"F8",X"91",X"F6",
		X"3A",X"F7",X"A1",X"F6",X"CF",X"F7",X"39",X"FF",X"6E",X"0A",X"35",X"0F",X"B1",X"0A",X"E4",X"05",
		X"66",X"01",X"8A",X"FC",X"38",X"F8",X"97",X"F6",X"43",X"F7",X"A6",X"F6",X"E2",X"F7",X"1A",X"FF",
		X"66",X"0A",X"5D",X"0F",X"AE",X"0A",X"F5",X"05",X"68",X"01",X"9D",X"FC",X"2C",X"F8",X"A1",X"F6",
		X"43",X"F7",X"B3",X"F6",X"E0",X"F7",X"00",X"FF",X"48",X"0A",X"3C",X"0F",X"BD",X"0A",X"FC",X"05",
		X"73",X"01",X"A4",X"FC",X"3E",X"F8",X"B0",X"F6",X"45",X"F7",X"BF",X"F6",X"EB",X"F7",X"23",X"FF",
		X"94",X"0A",X"1B",X"0F",X"6F",X"0A",X"9B",X"05",X"FD",X"00",X"02",X"FC",X"CE",X"F7",X"BC",X"F6",
		X"57",X"F7",X"A0",X"F6",X"01",X"F9",X"43",X"02",X"05",X"0D",X"14",X"0E",X"9B",X"08",X"F9",X"03",
		X"13",X"FF",X"0F",X"FA",X"EA",X"F6",X"1F",X"F7",X"13",X"F7",X"06",X"F7",X"8B",X"FC",X"D8",X"07",
		X"0E",X"0F",X"A0",X"0B",X"60",X"06",X"D9",X"01",X"C8",X"FC",X"5F",X"F8",X"C3",X"F6",X"5E",X"F7",
		X"C6",X"F6",X"4C",X"F8",X"1E",X"00",X"9F",X"0B",X"E3",X"0E",X"BE",X"09",X"16",X"05",X"64",X"00",
		X"74",X"FB",X"92",X"F7",X"E2",X"F6",X"63",X"F7",X"B5",X"F6",X"5A",X"F9",X"74",X"02",X"19",X"0D",
		X"45",X"0E",X"D8",X"08",X"61",X"04",X"A5",X"FF",X"C8",X"FA",X"57",X"F7",X"FD",X"F6",X"5F",X"F7",
		X"BD",X"F6",X"E5",X"F9",X"77",X"03",X"94",X"0D",X"F1",X"0D",X"86",X"08",X"21",X"04",X"66",X"FF",
		X"99",X"FA",X"4A",X"F7",X"0E",X"F7",X"60",X"F7",X"C9",X"F6",X"04",X"FA",X"7F",X"03",X"B4",X"0D",
		X"FC",X"0D",X"82",X"08",X"2A",X"04",X"6B",X"FF",X"A4",X"FA",X"45",X"F7",X"17",X"F7",X"61",X"F7",
		X"D9",X"F6",X"FA",X"F9",X"5E",X"03",X"B6",X"0D",X"02",X"0E",X"8B",X"08",X"33",X"04",X"74",X"FF",
		X"AA",X"FA",X"3F",X"F7",X"23",X"F7",X"63",X"F7",X"E8",X"F6",X"DF",X"F9",X"4A",X"03",X"83",X"0D",
		X"F3",X"0D",X"9E",X"08",X"35",X"04",X"83",X"FF",X"AC",X"FA",X"49",X"F7",X"29",X"F7",X"6A",X"F7",
		X"EF",X"F6",X"C0",X"F9",X"33",X"03",X"5A",X"0D",X"F3",X"0D",X"AE",X"08",X"3B",X"04",X"8E",X"FF",
		X"B5",X"FA",X"60",X"F7",X"29",X"F7",X"74",X"F7",X"EE",X"F6",X"98",X"F9",X"1D",X"03",X"38",X"0D",
		X"FF",X"0D",X"B6",X"08",X"48",X"04",X"96",X"FF",X"C1",X"FA",X"6D",X"F7",X"30",X"F7",X"7C",X"F7",
		X"F1",X"F6",X"80",X"F9",X"06",X"03",X"1E",X"0D",X"17",X"0E",X"B5",X"08",X"57",X"04",X"8D",X"FF",
		X"C7",X"FA",X"68",X"F7",X"42",X"F7",X"79",X"F7",X"FC",X"F6",X"EB",X"F9",X"1F",X"04",X"C4",X"0D",
		X"71",X"0D",X"E5",X"07",X"79",X"03",X"7D",X"FE",X"AD",X"F9",X"07",X"F7",X"81",X"F7",X"45",X"F7",
		X"74",X"F7",X"FB",X"FC",X"7E",X"08",X"07",X"0F",X"1D",X"0B",X"E4",X"05",X"46",X"01",X"17",X"FC",
		X"E8",X"F7",X"24",X"F7",X"9A",X"F7",X"06",X"F7",X"91",X"F9",X"4D",X"03",X"A9",X"0D",X"5E",X"0D",
		X"B3",X"07",X"1E",X"03",X"F1",X"FD",X"30",X"F9",X"12",X"F7",X"9C",X"F7",X"32",X"F7",X"F5",X"F7",
		X"A3",X"FF",X"B4",X"0B",X"8F",X"0E",X"1A",X"09",X"48",X"04",X"47",X"FF",X"1C",X"FA",X"36",X"F7",
		X"84",X"F7",X"5F",X"F7",X"89",X"F7",X"9C",X"FD",X"8E",X"09",X"DC",X"0E",X"25",X"0A",X"0C",X"05",
		X"22",X"00",X"E1",X"FA",X"78",X"F7",X"6F",X"F7",X"7E",X"F7",X"5A",X"F7",X"57",X"FC",X"1D",X"08",
		X"F8",X"0E",X"D6",X"0A",X"86",X"05",X"B3",X"00",X"59",X"FB",X"AC",X"F7",X"5F",X"F7",X"98",X"F7",
		X"41",X"F7",X"9C",X"FB",X"31",X"07",X"FF",X"0E",X"3B",X"0B",X"D0",X"05",X"FF",X"00",X"A2",X"FB",
		X"CA",X"F7",X"5C",X"F7",X"A3",X"F7",X"3B",X"F7",X"3C",X"FB",X"B7",X"06",X"F3",X"0E",X"73",X"0B",
		X"EF",X"05",X"26",X"01",X"BE",X"FB",X"DC",X"F7",X"5E",X"F7",X"AD",X"F7",X"3E",X"F7",X"21",X"FB",
		X"89",X"06",X"E6",X"0E",X"7D",X"0B",X"F8",X"05",X"2A",X"01",X"C2",X"FB",X"DF",X"F7",X"68",X"F7",
		X"AF",X"F7",X"48",X"F7",X"2E",X"FB",X"9B",X"06",X"D8",X"0E",X"6D",X"0B",X"E8",X"05",X"19",X"01",
		X"AC",X"FB",X"D9",X"F7",X"73",X"F7",X"B2",X"F7",X"54",X"F7",X"5D",X"FB",X"D9",X"06",X"CF",X"0E",
		X"46",X"0B",X"CB",X"05",X"F6",X"00",X"8A",X"FB",X"C8",X"F7",X"81",X"F7",X"B0",X"F7",X"60",X"F7",
		X"9F",X"FB",X"3E",X"07",X"D0",X"0E",X"11",X"0B",X"A2",X"05",X"C8",X"00",X"58",X"FB",X"AF",X"F7",
		X"90",X"F7",X"B0",X"F7",X"6B",X"F7",X"EB",X"FB",X"BD",X"07",X"DA",X"0E",X"CF",X"0A",X"73",X"05",
		X"90",X"00",X"21",X"FB",X"94",X"F7",X"9E",X"F7",X"B2",X"F7",X"72",X"F7",X"3C",X"FC",X"50",X"08",
		X"F4",X"0E",X"83",X"0A",X"3F",X"05",X"4C",X"00",X"EE",X"FA",X"97",X"F7",X"A6",X"F7",X"B6",X"F7",
		X"76",X"F7",X"92",X"FC",X"EF",X"08",X"1B",X"0F",X"30",X"0A",X"08",X"05",X"04",X"00",X"B1",X"FA",
		X"95",X"F7",X"B1",X"F7",X"B3",X"F7",X"93",X"F7",X"14",X"FD",X"75",X"09",X"FB",X"0E",X"E6",X"09",
		X"C7",X"04",X"BE",X"FF",X"72",X"FA",X"8F",X"F7",X"C0",X"F7",X"AF",X"F7",X"C2",X"F7",X"B1",X"FD",
		X"F3",X"09",X"C0",X"0E",X"99",X"09",X"83",X"04",X"75",X"FF",X"2C",X"FA",X"85",X"F7",X"D1",X"F7",
		X"A6",X"F7",X"ED",X"F7",X"4E",X"FE",X"81",X"0A",X"8A",X"0E",X"4A",X"09",X"3E",X"04",X"29",X"FF",
		X"E2",X"F9",X"77",X"F7",X"E1",X"F7",X"A1",X"F7",X"13",X"F8",X"E9",X"FE",X"17",X"0B",X"61",X"0E",
		X"F2",X"08",X"00",X"04",X"D4",X"FE",X"AF",X"F9",X"72",X"F7",X"F0",X"F7",X"9B",X"F7",X"2C",X"F8",
		X"3F",X"FF",X"5F",X"0B",X"5B",X"0E",X"FA",X"08",X"16",X"04",X"17",X"FF",X"E7",X"F9",X"81",X"F7",
		X"E5",X"F7",X"BD",X"F7",X"D9",X"F7",X"39",X"FD",X"FB",X"08",X"E6",X"0E",X"84",X"0A",X"67",X"05",
		X"B7",X"00",X"85",X"FB",X"00",X"F8",X"AF",X"F7",X"F7",X"F7",X"88",X"F7",X"DB",X"F9",X"58",X"03",
		X"9A",X"0D",X"62",X"0D",X"CA",X"07",X"56",X"03",X"57",X"FE",X"9C",X"F9",X"87",X"F7",X"F4",X"F7",
		X"CC",X"F7",X"C1",X"F7",X"2A",X"FC",X"8B",X"07",X"D3",X"0E",X"AF",X"0B",X"62",X"06",X"0D",X"02",
		X"EB",X"FC",X"D5",X"F8",X"8E",X"F7",X"0F",X"F8",X"AD",X"F7",X"38",X"F8",X"11",X"FE",X"90",X"09",
		X"FE",X"0E",X"B8",X"0A",X"B9",X"05",X"56",X"01",X"41",X"FC",X"79",X"F8",X"A2",X"F7",X"13",X"F8",
		X"AC",X"F7",X"72",X"F8",X"E7",X"FE",X"48",X"0A",X"EA",X"0E",X"5B",X"0A",X"85",X"05",X"17",X"01",
		X"16",X"FC",X"68",X"F8",X"AE",X"F7",X"14",X"F8",X"B5",X"F7",X"79",X"F8",X"E6",X"FE",X"5B",X"0A",
		X"0D",X"0F",X"51",X"0A",X"92",X"05",X"15",X"01",X"27",X"FC",X"6A",X"F8",X"BD",X"F7",X"13",X"F8",
		X"C7",X"F7",X"60",X"F8",X"CF",X"FE",X"36",X"0A",X"E1",X"0E",X"61",X"0A",X"9B",X"05",X"1F",X"01",
		X"33",X"FC",X"6F",X"F8",X"C3",X"F7",X"12",X"F8",X"D6",X"F7",X"40",X"F8",X"B4",X"FE",X"13",X"0A",
		X"C4",X"0E",X"75",X"0A",X"9E",X"05",X"2B",X"01",X"3B",X"FC",X"71",X"F8",X"C9",X"F7",X"17",X"F8",
		X"DF",X"F7",X"34",X"F8",X"A1",X"FE",X"EF",X"09",X"B8",X"0E",X"86",X"0A",X"A1",X"05",X"38",X"01",
		X"3C",X"FC",X"73",X"F8",X"CA",X"F7",X"27",X"F8",X"D8",X"F7",X"63",X"F8",X"3C",X"FF",X"C3",X"0A",
		X"8A",X"0E",X"D8",X"09",X"F3",X"04",X"5F",X"00",X"39",X"FB",X"24",X"F8",X"E6",X"F7",X"2E",X"F8",
		X"BD",X"F7",X"E6",X"F9",X"35",X"03",X"8B",X"0D",X"32",X"0D",X"A8",X"07",X"14",X"03",X"08",X"FE",
		X"5F",X"F9",X"D0",X"F7",X"25",X"F8",X"FD",X"F7",X"31",X"F8",X"1C",X"FE",X"DC",X"09",X"A1",X"0E",
		X"DB",X"09",X"DD",X"04",X"0D",X"00",X"D4",X"FA",X"F9",X"F7",X"0F",X"F8",X"25",X"F8",X"CF",X"F7",
		X"27",X"FB",X"75",X"06",X"C1",X"0E",X"87",X"0B",X"0D",X"06",X"6B",X"01",X"09",X"FC",X"5C",X"F8",
		X"F0",X"F7",X"3D",X"F8",X"D7",X"F7",X"F7",X"F9",X"CB",X"03",X"E2",X"0D",X"95",X"0C",X"EE",X"06",
		X"41",X"02",X"EE",X"FC",X"96",X"F8",X"ED",X"F7",X"3F",X"F8",X"ED",X"F7",X"31",X"F9",X"18",X"02",
		X"31",X"0D",X"46",X"0D",X"7A",X"07",X"D1",X"02",X"78",X"FD",X"F5",X"F8",X"E8",X"F7",X"46",X"F8",
		X"FB",X"F7",X"CA",X"F8",X"09",X"01",X"BC",X"0C",X"A6",X"0D",X"D3",X"07",X"1F",X"03",X"D1",X"FD",
		X"27",X"F9",X"EB",X"F7",X"49",X"F8",X"07",X"F8",X"97",X"F8",X"7B",X"00",X"6E",X"0C",X"D4",X"0D",
		X"01",X"08",X"47",X"03",X"F8",X"FD",X"3D",X"F9",X"F2",X"F7",X"4C",X"F8",X"10",X"F8",X"8F",X"F8",
		X"46",X"00",X"48",X"0C",X"DC",X"0D",X"10",X"08",X"4B",X"03",X"01",X"FE",X"3A",X"F9",X"F7",X"F7",
		X"51",X"F8",X"17",X"F8",X"A0",X"F8",X"56",X"00",X"47",X"0C",X"C8",X"0D",X"07",X"08",X"3B",X"03",
		X"F3",X"FD",X"26",X"F9",X"FC",X"F7",X"57",X"F8",X"1A",X"F8",X"BF",X"F8",X"93",X"00",X"61",X"0C",
		X"A4",X"0D",X"EA",X"07",X"1B",X"03",X"CF",X"FD",X"15",X"F9",X"03",X"F8",X"5D",X"F8",X"1B",X"F8",
		X"E6",X"F8",X"F1",X"00",X"95",X"0C",X"78",X"0D",X"BE",X"07",X"F3",X"02",X"9D",X"FD",X"0C",X"F9",
		X"0B",X"F8",X"63",X"F8",X"1C",X"F8",X"12",X"F9",X"69",X"01",X"DE",X"0C",X"46",X"0D",X"87",X"07",
		X"C1",X"02",X"60",X"FD",X"FA",X"F8",X"16",X"F8",X"6A",X"F8",X"1B",X"F8",X"3F",X"F9",X"F0",X"01",
		X"3C",X"0D",X"15",X"0D",X"45",X"07",X"8E",X"02",X"19",X"FD",X"E5",X"F8",X"1E",X"F8",X"72",X"F8",
		X"19",X"F8",X"6A",X"F9",X"7E",X"02",X"AB",X"0D",X"E0",X"0C",X"FE",X"06",X"55",X"02",X"CD",X"FC",
		X"C7",X"F8",X"28",X"F8",X"78",X"F8",X"19",X"F8",X"8B",X"F9",X"1C",X"03",X"F3",X"0D",X"9F",X"0C",
		X"B6",X"06",X"16",X"02",X"82",X"FC",X"9F",X"F8",X"37",X"F8",X"78",X"F8",X"21",X"F8",X"B3",X"F9",
		X"CD",X"03",X"02",X"0E",X"46",X"0C",X"77",X"06",X"C8",X"01",X"3E",X"FC",X"7E",X"F8",X"46",X"F8",
		X"76",X"F8",X"2B",X"F8",X"22",X"FA",X"7F",X"04",X"21",X"0E",X"EC",X"0B",X"38",X"06",X"79",X"01",
		X"FB",X"FB",X"79",X"F8",X"50",X"F8",X"78",X"F8",X"31",X"F8",X"89",X"FA",X"36",X"05",X"4E",X"0E",
		X"8C",X"0B",X"F7",X"05",X"2A",X"01",X"B3",X"FB",X"70",X"F8",X"5D",X"F8",X"7A",X"F8",X"36",X"F8",
		X"EB",X"FA",X"F0",X"05",X"89",X"0E",X"32",X"0B",X"B2",X"05",X"DE",X"00",X"67",X"FB",X"63",X"F8",
		X"68",X"F8",X"7E",X"F8",X"36",X"F8",X"45",X"FB",X"AD",X"06",X"D0",X"0E",X"D8",X"0A",X"6B",X"05",
		X"92",X"00",X"17",X"FB",X"56",X"F8",X"73",X"F8",X"83",X"F8",X"35",X"F8",X"9C",X"FB",X"63",X"07",
		X"C4",X"0E",X"89",X"0A",X"1D",X"05",X"4B",X"00",X"C3",X"FA",X"44",X"F8",X"7C",X"F8",X"89",X"F8",
		X"3B",X"F8",X"04",X"FC",X"11",X"08",X"98",X"0E",X"31",X"0A",X"D9",X"04",X"F4",X"FF",X"91",X"FA",
		X"4E",X"F8",X"84",X"F8",X"88",X"F8",X"58",X"F8",X"A2",X"FC",X"B3",X"08",X"7F",X"0E",X"D1",X"09",
		X"9D",X"04",X"9A",X"FF",X"5F",X"FA",X"51",X"F8",X"90",X"F8",X"84",X"F8",X"74",X"F8",X"37",X"FD",
		X"60",X"09",X"70",X"0E",X"71",X"09",X"5C",X"04",X"41",X"FF",X"28",X"FA",X"52",X"F8",X"9A",X"F8",
		X"80",X"F8",X"88",X"F8",X"C4",X"FD",X"12",X"0A",X"6F",X"0E",X"0B",X"09",X"1D",X"04",X"E5",X"FE",
		X"EC",X"F9",X"52",X"F8",X"A6",X"F8",X"7D",X"F8",X"9B",X"F8",X"47",X"FE",X"C9",X"0A",X"71",X"0E",
		X"AA",X"08",X"D8",X"03",X"93",X"FE",X"A7",X"F9",X"55",X"F8",X"AA",X"F8",X"86",X"F8",X"98",X"F8",
		X"E2",X"FE",X"3B",X"0B",X"10",X"0E",X"68",X"08",X"87",X"03",X"49",X"FE",X"7A",X"F9",X"66",X"F8",
		X"A7",X"F8",X"92",X"F8",X"B2",X"F8",X"8B",X"FF",X"AC",X"0B",X"C1",X"0D",X"19",X"08",X"3F",X"03",
		X"F3",X"FD",X"5E",X"F9",X"71",X"F8",X"AD",X"F8",X"8F",X"F8",X"F3",X"F8",X"44",X"00",X"21",X"0C",
		X"7A",X"0D",X"C6",X"07",X"FB",X"02",X"99",X"FD",X"40",X"F9",X"7A",X"F8",X"B6",X"F8",X"8B",X"F8",
		X"2D",X"F9",X"F8",X"00",X"A2",X"0C",X"3A",X"0D",X"70",X"07",X"B5",X"02",X"3F",X"FD",X"1A",X"F9",
		X"83",X"F8",X"BD",X"F8",X"87",X"F8",X"5D",X"F9",X"A7",X"01",X"2F",X"0D",X"05",X"0D",X"18",X"07",
		X"77",X"02",X"E9",X"FC",X"F8",X"F8",X"88",X"F8",X"C7",X"F8",X"85",X"F8",X"69",X"F9",X"94",X"01",
		X"0B",X"0D",X"31",X"0D",X"71",X"07",X"D7",X"02",X"8C",X"FD",X"4F",X"F9",X"89",X"F8",X"BF",X"F8",
		X"AB",X"F8",X"C2",X"F8",X"86",X"FE",X"5E",X"0A",X"4D",X"0E",X"48",X"09",X"6B",X"04",X"A2",X"FF",
		X"90",X"FA",X"87",X"F8",X"BC",X"F8",X"C0",X"F8",X"8D",X"F8",X"75",X"FA",X"4B",X"04",X"E1",X"0D",
		X"85",X"0C",X"EE",X"06",X"99",X"02",X"6B",X"FD",X"6B",X"F9",X"88",X"F8",X"D1",X"F8",X"B5",X"F8",
		X"A7",X"F8",X"AD",X"FC",X"EB",X"07",X"74",X"0E",X"F7",X"0A",X"C5",X"05",X"70",X"01",X"3B",X"FC",
		X"E4",X"F8",X"A4",X"F8",X"D1",X"F8",X"B9",X"F8",X"BD",X"F8",X"0D",X"FE",X"AD",X"09",X"8C",X"0E",
		X"28",X"0A",X"3D",X"05",X"D5",X"00",X"BB",X"FB",X"C1",X"F8",X"B6",X"F8",X"D3",X"F8",X"BE",X"F8",
		X"D5",X"F8",X"A4",X"FE",X"2B",X"0A",X"78",X"0E",X"EC",X"09",X"1D",X"05",X"B4",X"00",X"A3",X"FB",
		X"BC",X"F8",X"C1",X"F8",X"D4",X"F8",X"C3",X"F8",X"E6",X"F8",X"AF",X"FE",X"02",X"0A",X"65",X"0E",
		X"F9",X"09",X"27",X"05",X"BB",X"00",X"B1",X"FB",X"CF",X"F8",X"C5",X"F8",X"DB",X"F8",X"C8",X"F8",
		X"F3",X"F8",X"A3",X"FE",X"D8",X"09",X"5F",X"0E",X"03",X"0A",X"30",X"05",X"C2",X"00",X"BD",X"FB",
		X"DB",X"F8",X"CA",X"F8",X"E0",X"F8",X"CF",X"F8",X"FC",X"F8",X"8C",X"FE",X"B5",X"09",X"68",X"0E",
		X"0D",X"0A",X"3B",X"05",X"C7",X"00",X"CB",X"FB",X"E4",X"F8",X"CF",X"F8",X"E2",X"F8",X"D7",X"F8",
		X"FB",X"F8",X"6B",X"FE",X"9C",X"09",X"79",X"0E",X"12",X"0A",X"3A",X"05",X"BE",X"00",X"B5",X"FB",
		X"E4",X"F8",X"D6",X"F8",X"ED",X"F8",X"D2",X"F8",X"36",X"F9",X"A6",X"FF",X"08",X"0B",X"03",X"0E",
		X"FD",X"08",X"39",X"04",X"7E",X"FF",X"7A",X"FA",X"B2",X"F8",X"EE",X"F8",X"EF",X"F8",X"C1",X"F8",
		X"89",X"FA",X"5A",X"04",X"D5",X"0D",X"2E",X"0C",X"A7",X"06",X"32",X"02",X"F8",X"FC",X"24",X"F9",
		X"D8",X"F8",X"EF",X"F8",X"F7",X"F8",X"CF",X"F8",X"D9",X"FD",X"96",X"09",X"84",X"0E",X"C9",X"09",
		X"E7",X"04",X"4B",X"00",X"3C",X"FB",X"DB",X"F8",X"EC",X"F8",X"FD",X"F8",X"DA",X"F8",X"91",X"F9",
		X"F0",X"00",X"F1",X"0B",X"AB",X"0D",X"7C",X"08",X"E6",X"03",X"2F",X"FF",X"59",X"FA",X"C6",X"F8",
		X"FB",X"F8",X"03",X"F9",X"D2",X"F8",X"11",X"FA",X"94",X"02",X"EF",X"0C",X"2E",X"0D",X"DF",X"07",
		X"73",X"03",X"A8",X"FE",X"0B",X"FA",X"C9",X"F8",X"04",X"F9",X"06",X"F9",X"D4",X"F8",X"4B",X"FA",
		X"15",X"03",X"1A",X"0D",X"0B",X"0D",X"BE",X"07",X"60",X"03",X"93",X"FE",X"0B",X"FA",X"CF",X"F8",
		X"0C",X"F9",X"09",X"F9",X"E0",X"F8",X"4F",X"FA",X"F9",X"02",X"FC",X"0C",X"17",X"0D",X"C6",X"07",
		X"68",X"03",X"98",X"FE",X"1D",X"FA",X"DA",X"F8",X"0E",X"F9",X"0F",X"F9",X"E7",X"F8",X"47",X"FA",
		X"D3",X"02",X"EE",X"0C",X"24",X"0D",X"CE",X"07",X"73",X"03",X"A2",X"FE",X"2B",X"FA",X"E2",X"F8",
		X"10",X"F9",X"16",X"F9",X"ED",X"F8",X"34",X"FA",X"AA",X"02",X"F1",X"0C",X"36",X"0D",X"D7",X"07",
		X"7B",X"03",X"AB",X"FE",X"36",X"FA",X"E8",X"F8",X"15",X"F9",X"1C",X"F9",X"F0",X"F8",X"18",X"FA",
		X"82",X"02",X"02",X"0D",X"49",X"0D",X"D8",X"07",X"87",X"03",X"B1",X"FE",X"3F",X"FA",X"E9",X"F8",
		X"1B",X"F9",X"21",X"F9",X"F7",X"F8",X"F6",X"F9",X"6A",X"02",X"FF",X"0C",X"54",X"0D",X"DD",X"07",
		X"94",X"03",X"B5",X"FE",X"48",X"FA",X"E7",X"F8",X"29",X"F9",X"1E",X"F9",X"04",X"F9",X"05",X"FA",
		X"7B",X"02",X"EE",X"0C",X"31",X"0D",X"AF",X"07",X"5C",X"03",X"55",X"FE",X"0E",X"FA",X"EE",X"F8",
		X"30",X"F9",X"22",X"F9",X"01",X"F9",X"11",X"FB",X"53",X"05",X"FB",X"0D",X"B6",X"0B",X"3A",X"06",
		X"D4",X"01",X"83",X"FC",X"30",X"F9",X"1C",X"F9",X"27",X"F9",X"32",X"F9",X"0E",X"F9",X"B6",X"FE",
		X"88",X"0A",X"1C",X"0E",X"01",X"09",X"3E",X"04",X"79",X"FF",X"88",X"FA",X"FC",X"F8",X"33",X"F9",
		X"33",X"F9",X"0D",X"F9",X"45",X"FA",X"07",X"03",X"47",X"0D",X"BF",X"0C",X"46",X"07",X"E9",X"02",
		X"D9",X"FD",X"CD",X"F9",X"0C",X"F9",X"37",X"F9",X"3B",X"F9",X"01",X"F9",X"41",X"FB",X"8F",X"05",
		X"25",X"0E",X"CE",X"0B",X"69",X"06",X"27",X"02",X"05",X"FD",X"82",X"F9",X"1C",X"F9",X"3C",X"F9",
		X"40",X"F9",X"0C",X"F9",X"FF",X"FB",X"9F",X"06",X"48",X"0E",X"5A",X"0B",X"1E",X"06",X"D8",X"01",
		X"C3",X"FC",X"6F",X"F9",X"27",X"F9",X"3B",X"F9",X"4A",X"F9",X"07",X"F9",X"06",X"FC",X"BE",X"06",
		X"68",X"0E",X"53",X"0B",X"1E",X"06",X"DB",X"01",X"C9",X"FC",X"77",X"F9",X"29",X"F9",X"43",X"F9",
		X"4D",X"F9",X"0E",X"F9",X"00",X"FC",X"A4",X"06",X"5D",X"0E",X"56",X"0B",X"2A",X"06",X"E3",X"01",
		X"D3",X"FC",X"7A",X"F9",X"2C",X"F9",X"4A",X"F9",X"4E",X"F9",X"1B",X"F9",X"05",X"FC",X"81",X"06",
		X"32",X"0E",X"60",X"0B",X"33",X"06",X"E9",X"01",X"DE",X"FC",X"7A",X"F9",X"34",X"F9",X"4F",X"F9",
		X"52",X"F9",X"27",X"F9",X"01",X"FC",X"5C",X"06",X"13",X"0E",X"6B",X"0B",X"3B",X"06",X"F2",X"01",
		X"E5",X"FC",X"76",X"F9",X"3D",X"F9",X"51",X"F9",X"58",X"F9",X"2B",X"F9",X"F2",X"FB",X"35",X"06",
		X"06",X"0E",X"76",X"0B",X"42",X"06",X"FC",X"01",X"EA",X"FC",X"6F",X"F9",X"47",X"F9",X"54",X"F9",
		X"62",X"F9",X"2E",X"F9",X"D8",X"FB",X"13",X"06",X"08",X"0E",X"86",X"0B",X"48",X"06",X"07",X"02",
		X"EF",X"FC",X"84",X"F9",X"45",X"F9",X"5D",X"F9",X"61",X"F9",X"39",X"F9",X"2C",X"FC",X"EE",X"06",
		X"20",X"0E",X"E4",X"0A",X"A7",X"05",X"3E",X"01",X"04",X"FC",X"51",X"F9",X"59",X"F9",X"62",X"F9",
		X"61",X"F9",X"61",X"F9",X"18",X"FF",X"DA",X"0A",X"F2",X"0D",X"8E",X"08",X"E7",X"03",X"F5",X"FE",
		X"48",X"FA",X"37",X"F9",X"6D",X"F9",X"6C",X"F9",X"42",X"F9",X"E2",X"FA",X"75",X"04",X"F8",X"0D",
		X"E2",X"0B",X"6A",X"06",X"0E",X"02",X"D2",X"FC",X"88",X"F9",X"5C",X"F9",X"6B",X"F9",X"73",X"F9",
		X"4C",X"F9",X"E1",X"FC",X"FB",X"07",X"2B",X"0E",X"58",X"0A",X"48",X"05",X"DA",X"00",X"BD",X"FB",
		X"4F",X"F9",X"6E",X"F9",X"6D",X"F9",X"72",X"F9",X"71",X"F9",X"61",X"FE",X"A6",X"09",X"14",X"0E",
		X"89",X"09",X"C6",X"04",X"38",X"00",X"52",X"FB",X"4A",X"F9",X"7A",X"F9",X"6F",X"F9",X"79",X"F9",
		X"86",X"F9",X"F5",X"FE",X"20",X"0A",X"00",X"0E",X"4C",X"09",X"A6",X"04",X"10",X"00",X"41",X"FB",
		X"45",X"F9",X"85",X"F9",X"6C",X"F9",X"85",X"F9",X"83",X"F9",X"EB",X"FE",X"09",X"0A",X"02",X"0E",
		X"47",X"09",X"97",X"04",X"F2",X"FF",X"1C",X"FB",X"47",X"F9",X"8A",X"F9",X"75",X"F9",X"7F",X"F9",
		X"C6",X"F9",X"7C",X"00",X"B8",X"0B",X"74",X"0D",X"FF",X"07",X"8A",X"03",X"72",X"FE",X"30",X"FA",
		X"5C",X"F9",X"8D",X"F9",X"82",X"F9",X"6B",X"F9",X"4F",X"FB",X"93",X"05",X"F2",X"0D",X"11",X"0B",
		X"B8",X"05",X"26",X"01",X"DC",X"FB",X"69",X"F9",X"89",X"F9",X"84",X"F9",X"87",X"F9",X"D1",X"F9",
		X"AC",X"00",X"34",X"0C",X"16",X"0D",X"63",X"07",X"DA",X"02",X"84",X"FD",X"B7",X"F9",X"7F",X"F9",
		X"85",X"F9",X"A0",X"F9",X"51",X"F9",X"BF",X"FD",X"A1",X"09",X"E5",X"0D",X"C0",X"08",X"E2",X"03",
		X"C2",X"FE",X"3C",X"FA",X"72",X"F9",X"94",X"F9",X"98",X"F9",X"6E",X"F9",X"33",X"FC",X"61",X"07",
		X"77",X"0E",X"E8",X"09",X"E5",X"04",X"06",X"00",X"0A",X"FB",X"60",X"F9",X"A1",X"F9",X"8F",X"F9",
		X"8A",X"F9",X"38",X"FA",X"B2",X"02",X"21",X"0D",X"6C",X"0C",X"C2",X"06",X"63",X"02",X"1C",X"FD",
		X"BC",X"F9",X"89",X"F9",X"9C",X"F9",X"A1",X"F9",X"78",X"F9",X"B4",X"FC",X"C3",X"07",X"59",X"0E",
		X"1A",X"0A",X"26",X"05",X"80",X"00",X"6D",X"FB",X"66",X"F9",X"B0",X"F9",X"8F",X"F9",X"AA",X"F9",
		X"CF",X"F9",X"7A",X"00",X"C7",X"0B",X"32",X"0D",X"A8",X"07",X"2B",X"03",X"EB",X"FD",X"F5",X"F9",
		X"89",X"F9",X"A8",X"F9",X"A5",X"F9",X"88",X"F9",X"61",X"FC",X"96",X"07",X"42",X"0E",X"D2",X"09",
		X"CC",X"04",X"EC",X"FF",X"F2",X"FA",X"76",X"F9",X"B2",X"F9",X"A6",X"F9",X"98",X"F9",X"79",X"FA",
		X"5A",X"03",X"6D",X"0D",X"F6",X"0B",X"5A",X"06",X"EB",X"01",X"9C",X"FC",X"AD",X"F9",X"A6",X"F9",
		X"AA",X"F9",X"B9",X"F9",X"8B",X"F9",X"C0",X"FD",X"44",X"09",X"32",X"0E",X"39",X"09",X"7F",X"04",
		X"B4",X"FF",X"EC",X"FA",X"7B",X"F9",X"C1",X"F9",X"A5",X"F9",X"B6",X"F9",X"00",X"FA",X"F5",X"00",
		X"E5",X"0B",X"20",X"0D",X"CC",X"07",X"5F",X"03",X"64",X"FE",X"4C",X"FA",X"96",X"F9",X"B8",X"F9",
		X"B9",X"F9",X"A2",X"F9",X"97",X"FA",X"DB",X"02",X"06",X"0D",X"7B",X"0C",X"1A",X"07",X"CC",X"02",
		X"C3",X"FD",X"11",X"FA",X"A3",X"F9",X"B9",X"F9",X"C2",X"F9",X"9F",X"F9",X"DE",X"FA",X"91",X"03",
		X"48",X"0D",X"3C",X"0C",X"EA",X"06",X"A3",X"02",X"A0",X"FD",X"0B",X"FA",X"A9",X"F9",X"C2",X"F9",
		X"C5",X"F9",X"AB",X"F9",X"DD",X"FA",X"84",X"03",X"27",X"0D",X"40",X"0C",X"F3",X"06",X"AB",X"02",
		X"A9",X"FD",X"12",X"FA",X"AC",X"F9",X"C7",X"F9",X"C7",X"F9",X"B4",X"F9",X"C8",X"FA",X"62",X"03",
		X"0B",X"0D",X"4C",X"0C",X"F9",X"06",X"B5",X"02",X"B0",X"FD",X"18",X"FA",X"AD",X"F9",X"D0",X"F9",
		X"C7",X"F9",X"BE",X"F9",X"AD",X"FA",X"63",X"03",X"10",X"0D",X"39",X"0C",X"CB",X"06",X"81",X"02",
		X"58",X"FD",X"FC",X"F9",X"B9",X"F9",X"D3",X"F9",X"CF",X"F9",X"B4",X"F9",X"D7",X"FB",X"31",X"06",
		X"13",X"0E",X"A1",X"0A",X"73",X"05",X"E2",X"00",X"B6",X"FB",X"9D",X"F9",X"E0",X"F9",X"C4",X"F9",
		X"E1",X"F9",X"DF",X"F9",X"BB",X"FF",X"41",X"0B",X"51",X"0D",X"DA",X"07",X"5D",X"03",X"34",X"FE",
		X"29",X"FA",X"BA",X"F9",X"DE",X"F9",X"D6",X"F9",X"C6",X"F9",X"0E",X"FB",X"B3",X"04",X"8E",X"0D",
		X"65",X"0B",X"0A",X"06",X"AA",X"01",X"76",X"FC",X"D5",X"F9",X"D6",X"F9",X"DC",X"F9",X"E4",X"F9",
		X"BD",X"F9",X"D2",X"FC",X"BA",X"07",X"31",X"0E",X"0A",X"0A",X"1F",X"05",X"9E",X"00",X"98",X"FB",
		X"B1",X"F9",X"EA",X"F9",X"D7",X"F9",X"F0",X"F9",X"BD",X"F9",X"DA",X"FD",X"16",X"09",X"2D",X"0E",
		X"69",X"09",X"BB",X"04",X"24",X"00",X"46",X"FB",X"AD",X"F9",X"F3",X"F9",X"D9",X"F9",X"F6",X"F9",
		X"C9",X"F9",X"2C",X"FE",X"62",X"09",X"27",X"0E",X"46",X"09",X"B4",X"04",X"0D",X"00",X"51",X"FB",
		X"B5",X"F9",X"FA",X"F9",X"DC",X"F9",X"FC",X"F9",X"D3",X"F9",X"58",X"FE",X"A3",X"09",X"07",X"0E",
		X"EF",X"08",X"64",X"04",X"87",X"FF",X"EB",X"FA",X"B4",X"F9",X"07",X"FA",X"D9",X"F9",X"08",X"FA",
		X"F6",X"F9",X"07",X"01",X"0A",X"0C",X"BB",X"0C",X"42",X"07",X"C4",X"02",X"8E",X"FD",X"09",X"FA",
		X"F3",X"F9",X"E4",X"F9",X"0D",X"FA",X"B9",X"F9",X"2B",X"FC",X"30",X"07",X"E6",X"0D",X"C3",X"09",
		X"BC",X"04",X"DE",X"FF",X"F6",X"FA",X"C4",X"F9",X"0A",X"FA",X"E8",X"F9",X"00",X"FA",X"7F",X"FA",
		X"F4",X"02",X"4B",X"0D",X"9D",X"0B",X"12",X"06",X"71",X"01",X"23",X"FC",X"D7",X"F9",X"06",X"FA",
		X"EE",X"F9",X"11",X"FA",X"F0",X"F9",X"3B",X"00",X"B4",X"0B",X"BF",X"0C",X"0B",X"07",X"75",X"02",
		X"06",X"FD",X"E5",X"F9",X"07",X"FA",X"F5",X"F9",X"11",X"FA",X"E2",X"F9",X"E2",X"FD",X"99",X"09",
		X"DA",X"0D",X"6A",X"08",X"DD",X"03",X"A9",X"FE",X"90",X"FA",X"E1",X"F9",X"10",X"FA",X"FE",X"F9",
		X"FC",X"F9",X"05",X"FB",X"08",X"04",X"AB",X"0D",X"67",X"0B",X"01",X"06",X"8F",X"01",X"60",X"FC",
		X"EA",X"F9",X"11",X"FA",X"FC",X"F9",X"20",X"FA",X"DB",X"F9",X"2E",X"FD",X"6F",X"08",X"D1",X"0D",
		X"45",X"09",X"73",X"04",X"98",X"FF",X"E1",X"FA",X"DD",X"F9",X"20",X"FA",X"FC",X"F9",X"21",X"FA",
		X"2A",X"FA",X"F8",X"01",X"A1",X"0C",X"17",X"0C",X"8F",X"06",X"09",X"02",X"B5",X"FC",X"EA",X"F9",
		X"1E",X"FA",X"02",X"FA",X"29",X"FA",X"EA",X"F9",X"F9",X"FD",X"BD",X"09",X"A6",X"0D",X"3B",X"08",
		X"A3",X"03",X"61",X"FE",X"77",X"FA",X"FC",X"F9",X"1D",X"FA",X"15",X"FA",X"05",X"FA",X"72",X"FB",
		X"29",X"05",X"05",X"0E",X"B5",X"0A",X"77",X"05",X"E0",X"00",X"D2",X"FB",X"F4",X"F9",X"24",X"FA",
		X"11",X"FA",X"2B",X"FA",X"05",X"FA",X"80",X"FE",X"F5",X"09",X"95",X"0D",X"7B",X"08",X"EB",X"03",
		X"FC",X"FE",X"AC",X"FA",X"FD",X"F9",X"29",X"FA",X"1A",X"FA",X"25",X"FA",X"56",X"FA",X"25",X"01",
		X"0A",X"0C",X"D7",X"0C",X"50",X"07",X"07",X"03",X"ED",X"FD",X"66",X"FA",X"0D",X"FA",X"28",X"FA",
		X"22",X"FA",X"22",X"FA",X"96",X"FA",X"91",X"02",X"B2",X"0C",X"43",X"0C",X"DB",X"06",X"97",X"02",
		X"85",X"FD",X"48",X"FA",X"1B",X"FA",X"27",X"FA",X"2D",X"FA",X"1C",X"FA",X"C7",X"FA",X"E8",X"02",
		X"E0",X"0C",X"2C",X"0C",X"C6",X"06",X"8B",X"02",X"7C",X"FD",X"46",X"FA",X"21",X"FA",X"2B",X"FA",
		X"33",X"FA",X"20",X"FA",X"D9",X"FA",X"C7",X"02",X"F4",X"0C",X"41",X"0C",X"C6",X"06",X"98",X"02",
		X"7F",X"FD",X"4A",X"FA",X"21",X"FA",X"34",X"FA",X"32",X"FA",X"2A",X"FA",X"D8",X"FA",X"AD",X"02",
		X"E2",X"0C",X"42",X"0C",X"CE",X"06",X"A4",X"02",X"7F",X"FD",X"46",X"FA",X"25",X"FA",X"3A",X"FA",
		X"32",X"FA",X"37",X"FA",X"CD",X"FA",X"94",X"02",X"AF",X"0C",X"3C",X"0C",X"DC",X"06",X"AB",X"02",
		X"87",X"FD",X"4B",X"FA",X"2B",X"FA",X"40",X"FA",X"35",X"FA",X"3E",X"FA",X"BA",X"FA",X"71",X"02",
		X"8C",X"0C",X"3F",X"0C",X"E8",X"06",X"AE",X"02",X"94",X"FD",X"5C",X"FA",X"2E",X"FA",X"45",X"FA",
		X"37",X"FA",X"48",X"FA",X"9F",X"FA",X"6B",X"02",X"8B",X"0C",X"26",X"0C",X"C2",X"06",X"76",X"02",
		X"43",X"FD",X"43",X"FA",X"3C",X"FA",X"41",X"FA",X"49",X"FA",X"32",X"FA",X"97",X"FB",X"25",X"05",
		X"E8",X"0D",X"9B",X"0A",X"6E",X"05",X"CF",X"00",X"CF",X"FB",X"20",X"FA",X"51",X"FA",X"3D",X"FA",
		X"59",X"FA",X"35",X"FA",X"F2",X"FE",X"B0",X"0A",X"47",X"0D",X"9D",X"07",X"2A",X"03",X"CF",X"FD",
		X"6D",X"FA",X"40",X"FA",X"4A",X"FA",X"56",X"FA",X"30",X"FA",X"1C",X"FC",X"8D",X"06",X"DE",X"0D",
		X"86",X"09",X"8B",X"04",X"83",X"FF",X"E9",X"FA",X"2A",X"FA",X"5F",X"FA",X"43",X"FA",X"5E",X"FA",
		X"B0",X"FA",X"87",X"03",X"64",X"0D",X"DA",X"0A",X"84",X"05",X"B3",X"00",X"AF",X"FB",X"28",X"FA",
		X"64",X"FA",X"45",X"FA",X"68",X"FA",X"56",X"FA",X"45",X"00",X"9C",X"0B",X"B3",X"0C",X"F3",X"06",
		X"97",X"02",X"30",X"FD",X"4D",X"FA",X"56",X"FA",X"54",X"FA",X"64",X"FA",X"3D",X"FA",X"1A",X"FC",
		X"37",X"06",X"EF",X"0D",X"FE",X"09",X"08",X"05",X"4E",X"00",X"90",X"FB",X"30",X"FA",X"6C",X"FA",
		X"4A",X"FA",X"79",X"FA",X"32",X"FA",X"AC",X"FE",X"2E",X"0A",X"44",X"0D",X"F5",X"07",X"73",X"03",
		X"43",X"FE",X"9F",X"FA",X"4B",X"FA",X"68",X"FA",X"5C",X"FA",X"62",X"FA",X"06",X"FB",X"44",X"04",
		X"73",X"0D",X"A9",X"0A",X"6D",X"05",X"A9",X"00",X"B6",X"FB",X"3B",X"FA",X"71",X"FA",X"58",X"FA",
		X"78",X"FA",X"62",X"FA",X"07",X"00",X"B7",X"0B",X"A7",X"0C",X"C3",X"06",X"56",X"02",X"D0",X"FC",
		X"40",X"FA",X"74",X"FA",X"58",X"FA",X"84",X"FA",X"2C",X"FA",X"B0",X"FD",X"5A",X"09",X"49",X"0D",
		X"F3",X"07",X"40",X"03",X"E4",X"FD",X"7C",X"FA",X"6B",X"FA",X"63",X"FA",X"7D",X"FA",X"47",X"FA",
		X"9E",X"FC",X"8A",X"07",X"A8",X"0D",X"B3",X"08",X"E0",X"03",X"8E",X"FE",X"B2",X"FA",X"5E",X"FA",
		X"76",X"FA",X"70",X"FA",X"69",X"FA",X"AF",X"FB",X"AC",X"05",X"F3",X"0D",X"C2",X"09",X"C1",X"04",
		X"C8",X"FF",X"23",X"FB",X"4E",X"FA",X"83",X"FA",X"68",X"FA",X"88",X"FA",X"8D",X"FA",X"18",X"01",
		X"06",X"0C",X"46",X"0C",X"9C",X"06",X"47",X"02",X"E9",X"FC",X"59",X"FA",X"7D",X"FA",X"73",X"FA",
		X"83",X"FA",X"64",X"FA",X"0C",X"FC",X"0F",X"06",X"FA",X"0D",X"DD",X"09",X"F3",X"04",X"1E",X"00",
		X"76",X"FB",X"54",X"FA",X"8D",X"FA",X"6E",X"FA",X"96",X"FA",X"6C",X"FA",X"B1",X"FF",X"54",X"0B",
		X"C6",X"0C",X"06",X"07",X"A3",X"02",X"33",X"FD",X"74",X"FA",X"82",X"FA",X"7C",X"FA",X"8D",X"FA",
		X"64",X"FA",X"9A",X"FC",X"56",X"07",X"BA",X"0D",X"E0",X"08",X"14",X"04",X"E1",X"FE",X"D7",X"FA",
		X"6D",X"FA",X"8E",X"FA",X"7E",X"FA",X"8C",X"FA",X"04",X"FB",X"55",X"04",X"7C",X"0D",X"37",X"0A",
		X"0B",X"05",X"0B",X"00",X"52",X"FB",X"63",X"FA",X"99",X"FA",X"7C",X"FA",X"9D",X"FA",X"B9",X"FA",
		X"52",X"02",X"BB",X"0C",X"27",X"0B",X"A2",X"05",X"D3",X"00",X"C1",X"FB",X"68",X"FA",X"99",X"FA",
		X"82",X"FA",X"A1",X"FA",X"97",X"FA",X"E1",X"00",X"16",X"0C",X"EB",X"0B",X"3C",X"06",X"A0",X"01",
		X"60",X"FC",X"65",X"FA",X"A2",X"FA",X"7D",X"FA",X"B3",X"FA",X"50",X"FA",X"DF",X"FD",X"58",X"09",
		X"3A",X"0D",X"06",X"08",X"75",X"03",X"40",X"FE",X"C1",X"FA",X"87",X"FA",X"9B",X"FA",X"91",X"FA",
		X"9C",X"FA",X"F0",X"FA",X"FC",X"02",X"CF",X"0C",X"45",X"0B",X"EF",X"05",X"6D",X"01",X"58",X"FC",
		X"6D",X"FA",X"A8",X"FA",X"8A",X"FA",X"B1",X"FA",X"6D",X"FA",X"31",X"FD",X"0E",X"08",X"8A",X"0D",
		X"9A",X"08",X"ED",X"03",X"C4",X"FE",X"E3",X"FA",X"89",X"FA",X"A5",X"FA",X"97",X"FA",X"A7",X"FA",
		X"FD",X"FA",X"2B",X"03",X"FA",X"0C",X"D4",X"0A",X"80",X"05",X"B4",X"00",X"CC",X"FB",X"77",X"FA",
		X"B4",X"FA",X"8F",X"FA",X"C4",X"FA",X"73",X"FA",X"70",X"FF",X"26",X"0B",X"A3",X"0C",X"F6",X"06",
		X"8F",X"02",X"2D",X"FD",X"92",X"FA",X"A7",X"FA",X"A2",X"FA",X"AD",X"FA",X"98",X"FA",X"D1",X"FB",
		X"A8",X"05",X"A6",X"0D",X"D6",X"09",X"F5",X"04",X"1F",X"00",X"98",X"FB",X"7E",X"FA",X"BD",X"FA",
		X"95",X"FA",X"CE",X"FA",X"6F",X"FA",X"3E",X"FE",X"42",X"09",X"48",X"0D",X"30",X"08",X"C0",X"03",
		X"AE",X"FE",X"EB",X"FA",X"93",X"FA",X"BF",X"FA",X"9A",X"FA",X"D3",X"FA",X"7B",X"FA",X"DA",X"FF",
		X"F5",X"0A",X"AD",X"0C",X"67",X"07",X"14",X"03",X"00",X"FE",X"C9",X"FA",X"A3",X"FA",X"BB",X"FA",
		X"A5",X"FA",X"CF",X"FA",X"A0",X"FA",X"A6",X"00",X"7D",X"0B",X"6A",X"0C",X"23",X"07",X"D7",X"02",
		X"C4",X"FD",X"BB",X"FA",X"AE",X"FA",X"BC",X"FA",X"AE",X"FA",X"C9",X"FA",X"D6",X"FA",X"BD",X"01",
		X"61",X"0C",X"C1",X"0B",X"5E",X"06",X"F1",X"01",X"CE",X"FC",X"9B",X"FA",X"C3",X"FA",X"B1",X"FA",
		X"CA",X"FA",X"9D",X"FA",X"25",X"FC",X"33",X"06",X"75",X"0D",X"68",X"09",X"8A",X"04",X"86",X"FF",
		X"4C",X"FB",X"9E",X"FA",X"CE",X"FA",X"AA",X"FA",X"E0",X"FA",X"9D",X"FA",X"F1",X"00",X"FD",X"0B",
		X"C0",X"0B",X"37",X"06",X"9D",X"01",X"60",X"FC",X"9B",X"FA",X"D0",X"FA",X"B8",X"FA",X"D8",X"FA",
		X"9E",X"FA",X"E9",X"FD",X"7E",X"09",X"32",X"0D",X"73",X"07",X"F5",X"02",X"7E",X"FD",X"BB",X"FA",
		X"C5",X"FA",X"C3",X"FA",X"D2",X"FA",X"AA",X"FA",X"61",X"FC",X"44",X"07",X"79",X"0D",X"7E",X"08",
		X"CD",X"03",X"6A",X"FE",X"D3",X"FA",X"C3",X"FA",X"CD",X"FA",X"C8",X"FA",X"D0",X"FA",X"5E",X"FB",
		X"D0",X"03",X"43",X"0D",X"67",X"0A",X"2B",X"05",X"6C",X"00",X"AE",X"FB",X"AB",X"FA",X"DA",X"FA",
		X"C5",X"FA",X"E3",X"FA",X"AE",X"FA",X"6A",X"FE",X"B7",X"09",X"32",X"0D",X"A4",X"07",X"52",X"03",
		X"07",X"FE",X"D5",X"FA",X"C7",X"FA",X"D9",X"FA",X"C6",X"FA",X"EB",X"FA",X"DC",X"FA",X"2D",X"02",
		X"A8",X"0C",X"3B",X"0B",X"E7",X"05",X"4D",X"01",X"41",X"FC",X"A9",X"FA",X"E9",X"FA",X"C3",X"FA",
		X"F5",X"FA",X"9D",X"FA",X"31",X"FD",X"94",X"08",X"54",X"0D",X"FA",X"07",X"7D",X"03",X"10",X"FE",
		X"D1",X"FA",X"D5",X"FA",X"DB",X"FA",X"D8",X"FA",X"DE",X"FA",X"88",X"FB",X"73",X"04",X"68",X"0D",
		X"D1",X"09",X"B9",X"04",X"AB",X"FF",X"60",X"FB",X"C3",X"FA",X"EB",X"FA",X"CF",X"FA",X"FC",X"FA",
		X"CC",X"FA",X"BC",X"01",X"96",X"0C",X"05",X"0B",X"94",X"05",X"BC",X"00",X"CD",X"FB",X"B7",X"FA",
		X"F4",X"FA",X"CE",X"FA",X"02",X"FB",X"BD",X"FA",X"2C",X"00",X"77",X"0B",X"CA",X"0B",X"1F",X"06",
		X"70",X"01",X"21",X"FC",X"B9",X"FA",X"F6",X"FA",X"D6",X"FA",X"01",X"FB",X"BE",X"FA",X"3A",X"FF",
		X"BF",X"0A",X"36",X"0C",X"78",X"06",X"D0",X"01",X"6B",X"FC",X"C0",X"FA",X"F8",X"FA",X"DC",X"FA",
		X"03",X"FB",X"C1",X"FA",X"BE",X"FE",X"51",X"0A",X"6B",X"0C",X"A5",X"06",X"FF",X"01",X"8D",X"FC",
		X"C4",X"FA",X"F9",X"FA",X"E0",X"FA",X"04",X"FB",X"C3",X"FA",X"90",X"FE",X"23",X"0A",X"78",X"0C",
		X"B0",X"06",X"0B",X"02",X"8F",X"FC",X"C5",X"FA",X"01",X"FB",X"E4",X"FA",X"0B",X"FB",X"C6",X"FA",
		X"98",X"FE",X"2A",X"0A",X"6A",X"0C",X"A5",X"06",X"FE",X"01",X"7D",X"FC",X"C3",X"FA",X"05",X"FB",
		X"E4",X"FA",X"11",X"FB",X"C6",X"FA",X"C5",X"FE",X"5E",X"0A",X"49",X"0C",X"87",X"06",X"D6",X"01",
		X"70",X"FC",X"CC",X"FA",X"07",X"FB",X"EA",X"FA",X"14",X"FB",X"C6",X"FA",X"06",X"FF",X"B5",X"0A",
		X"1F",X"0C",X"5E",X"06",X"A3",X"01",X"56",X"FC",X"D4",X"FA",X"09",X"FB",X"ED",X"FA",X"1A",X"FB",
		X"C6",X"FA",X"52",X"FF",X"2A",X"0B",X"EF",X"0B",X"27",X"06",X"65",X"01",X"33",X"FC",X"DD",X"FA",
		X"0B",X"FB",X"F3",X"FA",X"1E",X"FB",X"C3",X"FA",X"A2",X"FF",X"B9",X"0B",X"C3",X"0B",X"E9",X"05",
		X"21",X"01",X"06",X"FC",X"E5",X"FA",X"0D",X"FB",X"F5",X"FA",X"22",X"FB",X"D0",X"FA",X"2D",X"00",
		X"EB",X"0B",X"6A",X"0B",X"B2",X"05",X"CE",X"00",X"D7",X"FB",X"EB",X"FA",X"12",X"FB",X"F9",X"FA",
		X"25",X"FB",X"ED",X"FA",X"DE",X"00",X"1A",X"0C",X"0D",X"0B",X"75",X"05",X"7E",X"00",X"A0",X"FB",
		X"EF",X"FA",X"17",X"FB",X"FE",X"FA",X"25",X"FB",X"05",X"FB",X"90",X"01",X"59",X"0C",X"AD",X"0A",
		X"35",X"05",X"27",X"00",X"88",X"FB",X"F4",X"FA",X"19",X"FB",X"01",X"FB",X"26",X"FB",X"19",X"FB",
		X"40",X"02",X"AE",X"0C",X"4A",X"0A",X"F7",X"04",X"CA",X"FF",X"78",X"FB",X"F9",X"FA",X"1F",X"FB",
		X"03",X"FB",X"2D",X"FB",X"24",X"FB",X"DF",X"02",X"FF",X"0C",X"09",X"0A",X"D4",X"04",X"B0",X"FF",
		X"79",X"FB",X"00",X"FB",X"20",X"FB",X"08",X"FB",X"30",X"FB",X"0E",X"FB",X"4D",X"01",X"08",X"0C",
		X"23",X"0B",X"B2",X"05",X"00",X"01",X"0B",X"FC",X"F4",X"FA",X"25",X"FB",X"0C",X"FB",X"31",X"FB",
		X"E8",X"FA",X"7F",X"FD",X"6B",X"08",X"05",X"0D",X"DA",X"07",X"69",X"03",X"18",X"FE",X"17",X"FB",
		X"18",X"FB",X"20",X"FB",X"15",X"FB",X"32",X"FB",X"30",X"FB",X"26",X"02",X"5F",X"0C",X"D2",X"0A",
		X"80",X"05",X"C5",X"00",X"ED",X"FB",X"FE",X"FA",X"2C",X"FB",X"14",X"FB",X"3C",X"FB",X"EC",X"FA",
		X"0B",X"FE",X"91",X"09",X"B4",X"0C",X"13",X"07",X"96",X"02",X"32",X"FD",X"07",X"FB",X"26",X"FB",
		X"24",X"FB",X"2A",X"FB",X"1C",X"FB",X"60",X"FC",X"6D",X"06",X"3E",X"0D",X"61",X"08",X"AF",X"03",
		X"3E",X"FE",X"20",X"FB",X"25",X"FB",X"2D",X"FB",X"21",X"FB",X"3B",X"FB",X"63",X"FB",X"48",X"04",
		X"7A",X"0D",X"47",X"09",X"5D",X"04",X"07",X"FF",X"5E",X"FB",X"1B",X"FB",X"36",X"FB",X"1D",X"FB",
		X"48",X"FB",X"3A",X"FB",X"FC",X"02",X"02",X"0D",X"EB",X"09",X"BF",X"04",X"9B",X"FF",X"83",X"FB",
		X"1F",X"FB",X"38",X"FB",X"24",X"FB",X"4A",X"FB",X"1F",X"FB",X"08",X"01",X"D8",X"0B",X"29",X"0B",
		X"B5",X"05",X"06",X"01",X"10",X"FC",X"0E",X"FB",X"3D",X"FB",X"29",X"FB",X"47",X"FB",X"0B",X"FB",
		X"4C",X"FD",X"F8",X"07",X"02",X"0D",X"EF",X"07",X"7D",X"03",X"32",X"FE",X"30",X"FB",X"33",X"FB",
		X"3A",X"FB",X"2F",X"FB",X"4D",X"FB",X"2F",X"FB",X"F5",X"00",X"AC",X"0B",X"69",X"0B",X"F4",X"05",
		X"68",X"01",X"66",X"FC",X"1C",X"FB",X"3F",X"FB",X"37",X"FB",X"46",X"FB",X"26",X"FB",X"D4",X"FC",
		X"15",X"07",X"1A",X"0D",X"22",X"08",X"8E",X"03",X"2A",X"FE",X"31",X"FB",X"3C",X"FB",X"43",X"FB",
		X"36",X"FB",X"54",X"FB",X"61",X"FB",X"1B",X"03",X"DE",X"0C",X"ED",X"09",X"D4",X"04",X"C0",X"FF",
		X"9E",X"FB",X"2D",X"FB",X"4C",X"FB",X"34",X"FB",X"60",X"FB",X"22",X"FB",X"7B",X"00",X"9B",X"0B",
		X"36",X"0B",X"A3",X"05",X"DA",X"00",X"ED",X"FB",X"28",X"FB",X"4F",X"FB",X"39",X"FB",X"63",X"FB",
		X"08",X"FB",X"CE",X"FE",X"A7",X"0A",X"04",X"0C",X"30",X"06",X"8A",X"01",X"52",X"FC",X"2F",X"FB",
		X"4C",X"FB",X"44",X"FB",X"5A",X"FB",X"1F",X"FB",X"CD",X"FD",X"46",X"09",X"A9",X"0C",X"F6",X"06",
		X"81",X"02",X"25",X"FD",X"38",X"FB",X"49",X"FB",X"53",X"FB",X"46",X"FB",X"57",X"FB",X"D8",X"FB",
		X"DD",X"04",X"4A",X"0D",X"37",X"09",X"69",X"04",X"5B",X"FF",X"97",X"FB",X"3D",X"FB",X"58",X"FB",
		X"43",X"FB",X"6F",X"FB",X"14",X"FB",X"74",X"FE",X"E9",X"09",X"86",X"0C",X"F2",X"06",X"9B",X"02",
		X"53",X"FD",X"3B",X"FB",X"4F",X"FB",X"5B",X"FB",X"4A",X"FB",X"68",X"FB",X"84",X"FB",X"8E",X"03",
		X"EE",X"0C",X"C4",X"09",X"C4",X"04",X"C1",X"FF",X"B0",X"FB",X"43",X"FB",X"60",X"FB",X"4A",X"FB",
		X"76",X"FB",X"18",X"FB",X"21",X"FF",X"DB",X"0A",X"EE",X"0B",X"2B",X"06",X"9F",X"01",X"79",X"FC",
		X"44",X"FB",X"5A",X"FB",X"5C",X"FB",X"5F",X"FB",X"4E",X"FB",X"DB",X"FC",X"13",X"07",X"FF",X"0C",
		X"08",X"08",X"80",X"03",X"2D",X"FE",X"4F",X"FB",X"5E",X"FB",X"61",X"FB",X"57",X"FB",X"77",X"FB",
		X"4B",X"FB",X"CB",X"00",X"97",X"0B",X"5C",X"0B",X"E8",X"05",X"74",X"01",X"87",X"FC",X"4B",X"FB",
		X"5E",X"FB",X"68",X"FB",X"5F",X"FB",X"6D",X"FB",X"C6",X"FB",X"31",X"04",X"E1",X"0C",X"C3",X"09",
		X"E1",X"04",X"22",X"00",X"CC",X"FB",X"51",X"FB",X"67",X"FB",X"67",X"FB",X"6A",X"FB",X"60",X"FB",
		X"54",X"FC",X"FD",X"05",X"46",X"0D",X"F1",X"08",X"65",X"04",X"7A",X"FF",X"AA",X"FB",X"58",X"FB",
		X"6E",X"FB",X"67",X"FB",X"75",X"FB",X"57",X"FB",X"9F",X"FC",X"9A",X"06",X"3E",X"0D",X"A4",X"08",
		X"31",X"04",X"2B",X"FF",X"98",X"FB",X"5D",X"FB",X"74",X"FB",X"64",X"FB",X"82",X"FB",X"4A",X"FB",
		X"CA",X"FD",X"83",X"08",X"D3",X"0C",X"68",X"07",X"16",X"03",X"C3",X"FD",X"6A",X"FB",X"67",X"FB",
		X"7D",X"FB",X"60",X"FB",X"97",X"FB",X"43",X"FB",X"A7",X"01",X"6B",X"0C",X"97",X"0A",X"3D",X"05",
		X"78",X"00",X"FB",X"FB",X"65",X"FB",X"73",X"FB",X"75",X"FB",X"80",X"FB",X"59",X"FB",X"46",X"FD",
		X"3C",X"08",X"F0",X"0C",X"76",X"07",X"1C",X"03",X"CD",X"FD",X"70",X"FB",X"70",X"FB",X"82",X"FB",
		X"68",X"FB",X"9A",X"FB",X"4B",X"FB",X"CF",X"00",X"85",X"0B",X"42",X"0B",X"E5",X"05",X"7A",X"01",
		X"8B",X"FC",X"5C",X"FB",X"7D",X"FB",X"7F",X"FB",X"76",X"FB",X"90",X"FB",X"B5",X"FB",X"5D",X"03",
		X"D5",X"0C",X"EB",X"09",X"E9",X"04",X"1B",X"00",X"ED",X"FB",X"71",X"FB",X"80",X"FB",X"7E",X"FB",
		X"8B",X"FB",X"63",X"FB",X"3E",X"FD",X"02",X"08",X"DC",X"0C",X"77",X"07",X"0E",X"03",X"B6",X"FD",
		X"75",X"FB",X"7A",X"FB",X"8E",X"FB",X"71",X"FB",X"A4",X"FB",X"70",X"FB",X"A7",X"02",X"E1",X"0C",
		X"DD",X"09",X"C0",X"04",X"BE",X"FF",X"C4",X"FB",X"7D",X"FB",X"87",X"FB",X"82",X"FB",X"9C",X"FB",
		X"58",X"FB",X"2D",X"FE",X"88",X"09",X"6A",X"0C",X"BF",X"06",X"6C",X"02",X"2B",X"FD",X"77",X"FB",
		X"82",X"FB",X"95",X"FB",X"7A",X"FB",X"AA",X"FB",X"7E",X"FB",X"3B",X"02",X"42",X"0C",X"6F",X"0A",
		X"46",X"05",X"AD",X"00",X"26",X"FC",X"7B",X"FB",X"88",X"FB",X"95",X"FB",X"87",X"FB",X"9A",X"FB",
		X"16",X"FC",X"C4",X"04",X"0B",X"0D",X"41",X"09",X"82",X"04",X"AC",X"FF",X"D8",X"FB",X"87",X"FB",
		X"8E",X"FB",X"95",X"FB",X"92",X"FB",X"8D",X"FB",X"9E",X"FC",X"F7",X"05",X"05",X"0D",X"BD",X"08",
		X"30",X"04",X"48",X"FF",X"C2",X"FB",X"8D",X"FB",X"91",X"FB",X"97",X"FB",X"98",X"FB",X"8D",X"FB",
		X"B4",X"FC",X"46",X"06",X"15",X"0D",X"82",X"08",X"05",X"04",X"F8",X"FE",X"B4",X"FB",X"8F",X"FB",
		X"9B",X"FB",X"93",X"FB",X"AA",X"FB",X"76",X"FB",X"01",X"FE",X"A6",X"08",X"6E",X"0C",X"19",X"07",
		X"B9",X"02",X"71",X"FD",X"7A",X"FB",X"9A",X"FB",X"9F",X"FB",X"91",X"FB",X"B7",X"FB",X"9E",X"FB",
		X"4A",X"02",X"40",X"0C",X"FD",X"09",X"DF",X"04",X"F0",X"FF",X"DA",X"FB",X"93",X"FB",X"9F",X"FB",
		X"9D",X"FB",X"AD",X"FB",X"83",X"FB",X"B2",X"FD",X"44",X"08",X"89",X"0C",X"2F",X"07",X"DB",X"02",
		X"84",X"FD",X"7F",X"FB",X"A0",X"FB",X"A9",X"FB",X"94",X"FB",X"C6",X"FB",X"66",X"FB",X"7B",X"00",
		X"96",X"0B",X"3B",X"0B",X"C6",X"05",X"60",X"01",X"90",X"FC",X"97",X"FB",X"9C",X"FB",X"B2",X"FB",
		X"97",X"FB",X"C4",X"FB",X"BB",X"FB",X"A7",X"02",X"51",X"0C",X"38",X"0A",X"1F",X"05",X"8D",X"00",
		X"2B",X"FC",X"A1",X"FB",X"9F",X"FB",X"B5",X"FB",X"9D",X"FB",X"C0",X"FB",X"F2",X"FB",X"8F",X"03",
		X"8A",X"0C",X"D5",X"09",X"E3",X"04",X"46",X"00",X"16",X"FC",X"A7",X"FB",X"A1",X"FB",X"BB",X"FB",
		X"9F",X"FB",X"C6",X"FB",X"EA",X"FB",X"90",X"03",X"A8",X"0C",X"D7",X"09",X"E5",X"04",X"4D",X"00",
		X"1E",X"FC",X"AA",X"FB",X"A4",X"FB",X"C0",X"FB",X"A1",X"FB",X"D0",X"FB",X"C7",X"FB",X"6C",X"03",
		X"CE",X"0C",X"DB",X"09",X"EF",X"04",X"54",X"00",X"25",X"FC",X"AA",X"FB",X"AB",X"FB",X"C1",X"FB",
		X"A6",X"FB",X"D0",X"FB",X"CB",X"FB",X"5C",X"03",X"91",X"0C",X"DE",X"09",X"F8",X"04",X"5B",X"00",
		X"25",X"FC",X"AA",X"FB",X"B0",X"FB",X"C2",X"FB",X"AC",X"FB",X"CF",X"FB",X"DE",X"FB",X"46",X"03",
		X"63",X"0C",X"E7",X"09",X"FE",X"04",X"65",X"00",X"23",X"FC",X"AE",X"FB",X"B4",X"FB",X"C4",X"FB",
		X"B1",X"FB",X"D1",X"FB",X"EB",X"FB",X"25",X"03",X"45",X"0C",X"F5",X"09",X"06",X"05",X"6D",X"00",
		X"19",X"FC",X"B3",X"FB",X"B6",X"FB",X"C8",X"FB",X"B4",X"FB",X"D5",X"FB",X"EC",X"FB",X"FF",X"02",
		X"39",X"0C",X"04",X"0A",X"09",X"05",X"74",X"00",X"27",X"FC",X"BA",X"FB",X"B7",X"FB",X"CE",X"FB",
		X"B4",X"FB",X"DE",X"FB",X"E2",X"FB",X"D6",X"02",X"40",X"0C",X"12",X"0A",X"0D",X"05",X"80",X"00",
		X"36",X"FC",X"C1",X"FB",X"B7",X"FB",X"D5",X"FB",X"B3",X"FB",X"E7",X"FB",X"CC",X"FB",X"AE",X"02",
		X"56",X"0C",X"1F",X"0A",X"12",X"05",X"8B",X"00",X"40",X"FC",X"C5",X"FB",X"BA",X"FB",X"DB",X"FB",
		X"B4",X"FB",X"F1",X"FB",X"AA",X"FB",X"86",X"02",X"7C",X"0C",X"25",X"0A",X"19",X"05",X"92",X"00",
		X"47",X"FC",X"C6",X"FB",X"C0",X"FB",X"DD",X"FB",X"BA",X"FB",X"EF",X"FB",X"BE",X"FB",X"81",X"02",
		X"3A",X"0C",X"28",X"0A",X"22",X"05",X"9A",X"00",X"4C",X"FC",X"C5",X"FB",X"C4",X"FB",X"DC",X"FB",
		X"C0",X"FB",X"EF",X"FB",X"CC",X"FB",X"6E",X"02",X"08",X"0C",X"2F",X"0A",X"2A",X"05",X"A3",X"00",
		X"4C",X"FC",X"C7",X"FB",X"CA",X"FB",X"E0",X"FB",X"C6",X"FB",X"F0",X"FB",X"D7",X"FB",X"4F",X"02",
		X"E9",X"0B",X"3B",X"0A",X"30",X"05",X"AB",X"00",X"46",X"FC",X"CC",X"FB",X"CD",X"FB",X"E3",X"FB",
		X"C8",X"FB",X"F4",X"FB",X"DB",X"FB",X"3A",X"02",X"E8",X"0B",X"27",X"0A",X"13",X"05",X"74",X"00",
		X"28",X"FC",X"D6",X"FB",X"CD",X"FB",X"E7",X"FB",X"CC",X"FB",X"EF",X"FB",X"39",X"FC",X"CD",X"04",
		X"C7",X"0C",X"85",X"08",X"E6",X"03",X"B5",X"FE",X"D4",X"FB",X"E1",X"FB",X"DB",X"FB",X"DE",X"FB",
		X"ED",X"FB",X"B9",X"FB",X"CB",X"FE",X"B7",X"09",X"A8",X"0B",X"2B",X"06",X"BD",X"01",X"CD",X"FC",
		X"D4",X"FB",X"D4",X"FB",X"F0",X"FB",X"CD",X"FB",X"07",X"FC",X"D2",X"FB",X"59",X"02",X"12",X"0C",
		X"D6",X"09",X"CD",X"04",X"0B",X"00",X"0A",X"FC",X"E5",X"FB",X"D8",X"FB",X"F3",X"FB",X"DA",X"FB",
		X"F4",X"FB",X"63",X"FC",X"DA",X"04",X"91",X"0C",X"A6",X"08",X"07",X"04",X"03",X"FF",X"E9",X"FB",
		X"E8",X"FB",X"E2",X"FB",X"E9",X"FB",X"F1",X"FB",X"CE",X"FB",X"60",X"FD",X"0F",X"08",X"5F",X"0C",
		X"DE",X"06",X"84",X"02",X"3E",X"FD",X"CF",X"FB",X"E5",X"FB",X"F7",X"FB",X"D8",X"FB",X"15",X"FC",
		X"B0",X"FB",X"FD",X"01",X"31",X"0C",X"9B",X"09",X"7E",X"04",X"75",X"FF",X"ED",X"FB",X"F3",X"FB",
		X"E6",X"FB",X"EF",X"FB",X"FC",X"FB",X"CC",X"FB",X"8D",X"FE",X"A9",X"09",X"66",X"0B",X"D2",X"05",
		X"22",X"01",X"6C",X"FC",X"F3",X"FB",X"DF",X"FB",X"04",X"FC",X"E5",X"FB",X"FB",X"FB",X"F5",X"FC",
		X"5E",X"07",X"7E",X"0C",X"C3",X"06",X"42",X"02",X"FD",X"FC",X"E9",X"FB",X"E6",X"FB",X"09",X"FC",
		X"DF",X"FB",X"13",X"FC",X"5C",X"FC",X"60",X"05",X"9F",X"0C",X"A7",X"07",X"1A",X"03",X"A1",X"FD",
		X"D5",X"FB",X"F4",X"FB",X"01",X"FC",X"E6",X"FB",X"1F",X"FC",X"BC",X"FB",X"94",X"01",X"03",X"0C",
		X"D2",X"09",X"A2",X"04",X"BF",X"FF",X"FD",X"FB",X"07",X"FC",X"E7",X"FB",X"0C",X"FC",X"F2",X"FB",
		X"FE",X"FB",X"12",X"FD",X"43",X"07",X"A5",X"0C",X"2F",X"07",X"EA",X"02",X"9F",X"FD",X"E4",X"FB",
		X"FA",X"FB",X"03",X"FC",X"F4",X"FB",X"1A",X"FC",X"D1",X"FB",X"3B",X"FF",X"E8",X"09",X"6A",X"0B",
		X"04",X"06",X"A8",X"01",X"D6",X"FC",X"F1",X"FB",X"F7",X"FB",X"0F",X"FC",X"F0",X"FB",X"26",X"FC",
		X"D4",X"FB",X"B5",X"00",X"08",X"0B",X"B3",X"0A",X"76",X"05",X"04",X"01",X"8F",X"FC",X"00",X"FC",
		X"F6",X"FB",X"16",X"FC",X"F0",X"FB",X"2B",X"FC",X"E0",X"FB",X"3D",X"01",X"4D",X"0B",X"79",X"0A",
		X"52",X"05",X"DE",X"00",X"7E",X"FC",X"02",X"FC",X"F9",X"FB",X"19",X"FC",X"F3",X"FB",X"2F",X"FC",
		X"E3",X"FB",X"24",X"01",X"39",X"0B",X"85",X"0A",X"57",X"05",X"EA",X"00",X"7C",X"FC",X"08",X"FC",
		X"FB",X"FB",X"1E",X"FC",X"F7",X"FB",X"34",X"FC",X"DD",X"FB",X"F8",X"00",X"31",X"0B",X"94",X"0A",
		X"5B",X"05",X"F3",X"00",X"74",X"FC",X"0C",X"FC",X"FF",X"FB",X"21",X"FC",X"F8",X"FB",X"3B",X"FC",
		X"CE",X"FB",X"C6",X"00",X"3D",X"0B",X"A3",X"0A",X"60",X"05",X"FA",X"00",X"75",X"FC",X"10",X"FC",
		X"01",X"FC",X"25",X"FC",X"FB",X"FB",X"3C",X"FC",X"CD",X"FB",X"AA",X"00",X"54",X"0B",X"B6",X"0A",
		X"63",X"05",X"05",X"01",X"85",X"FC",X"17",X"FC",X"04",X"FC",X"29",X"FC",X"00",X"FC",X"3E",X"FC",
		X"DB",X"FB",X"A9",X"00",X"30",X"0B",X"B7",X"0A",X"6A",X"05",X"0C",X"01",X"93",X"FC",X"1A",X"FC",
		X"05",X"FC",X"2C",X"FC",X"02",X"FC",X"40",X"FC",X"E3",X"FB",X"A0",X"00",X"F6",X"0A",X"B4",X"0A",
		X"76",X"05",X"13",X"01",X"9D",X"FC",X"1B",X"FC",X"08",X"FC",X"2F",X"FC",X"06",X"FC",X"43",X"FC",
		X"EA",X"FB",X"8A",X"00",X"CB",X"0A",X"BB",X"0A",X"7D",X"05",X"1C",X"01",X"A5",X"FC",X"1C",X"FC",
		X"0E",X"FC",X"31",X"FC",X"09",X"FC",X"45",X"FC",X"ED",X"FB",X"67",X"00",X"B2",X"0A",X"C6",X"0A",
		X"83",X"05",X"24",X"01",X"A5",X"FC",X"1E",X"FC",X"12",X"FC",X"35",X"FC",X"0D",X"FC",X"4B",X"FC",
		X"E8",X"FB",X"39",X"00",X"A7",X"0A",X"D4",X"0A",X"89",X"05",X"2B",X"01",X"9F",X"FC",X"22",X"FC",
		X"13",X"FC",X"39",X"FC",X"0C",X"FC",X"52",X"FC",X"EF",X"FB",X"34",X"01",X"59",X"0B",X"01",X"0A",
		X"D6",X"04",X"19",X"00",X"40",X"FC",X"37",X"FC",X"10",X"FC",X"40",X"FC",X"12",X"FC",X"46",X"FC",
		X"7C",X"FC",X"9D",X"05",X"68",X"0C",X"82",X"07",X"F5",X"02",X"C3",X"FD",X"15",X"FC",X"24",X"FC",
		X"37",X"FC",X"16",X"FC",X"5A",X"FC",X"D3",X"FB",X"8B",X"00",X"48",X"0B",X"DC",X"09",X"9F",X"04",
		X"99",X"FF",X"22",X"FC",X"42",X"FC",X"1B",X"FC",X"3F",X"FC",X"28",X"FC",X"28",X"FC",X"1D",X"FE",
		X"19",X"09",X"6F",X"0B",X"AB",X"05",X"0D",X"01",X"6C",X"FC",X"42",X"FC",X"14",X"FC",X"4E",X"FC",
		X"18",X"FC",X"4F",X"FC",X"C6",X"FC",X"E8",X"06",X"FA",X"0B",X"8C",X"06",X"E6",X"01",X"C3",X"FC",
		X"32",X"FC",X"21",X"FC",X"4D",X"FC",X"1B",X"FC",X"5A",X"FC",X"66",X"FC",X"77",X"05",X"41",X"0C",
		X"1C",X"07",X"6B",X"02",X"27",X"FD",X"30",X"FC",X"28",X"FC",X"4E",X"FC",X"1D",X"FC",X"63",X"FC",
		X"43",X"FC",X"A0",X"04",X"59",X"0C",X"72",X"07",X"B2",X"02",X"5F",X"FD",X"2E",X"FC",X"2E",X"FC",
		X"4F",X"FC",X"21",X"FC",X"66",X"FC",X"35",X"FC",X"33",X"04",X"57",X"0C",X"99",X"07",X"CD",X"02",
		X"75",X"FD",X"2D",X"FC",X"32",X"FC",X"51",X"FC",X"25",X"FC",X"6A",X"FC",X"30",X"FC",X"16",X"04",
		X"4B",X"0C",X"99",X"07",X"CA",X"02",X"6B",X"FD",X"2D",X"FC",X"35",X"FC",X"54",X"FC",X"28",X"FC",
		X"6F",X"FC",X"2B",X"FC",X"36",X"04",X"3D",X"0C",X"7E",X"07",X"B8",X"02",X"4B",X"FD",X"30",X"FC",
		X"37",X"FC",X"58",X"FC",X"28",X"FC",X"77",X"FC",X"27",X"FC",X"81",X"04",X"33",X"0C",X"4D",X"07",
		X"90",X"02",X"34",X"FD",X"3C",X"FC",X"32",X"FC",X"62",X"FC",X"24",X"FC",X"80",X"FC",X"31",X"FC",
		X"EF",X"04",X"2A",X"0C",X"1D",X"07",X"6E",X"02",X"2D",X"FD",X"43",X"FC",X"36",X"FC",X"63",X"FC",
		X"29",X"FC",X"80",X"FC",X"15",X"FC",X"93",X"03",X"26",X"0C",X"0E",X"08",X"47",X"03",X"09",X"FE",
		X"2C",X"FC",X"52",X"FC",X"4F",X"FC",X"46",X"FC",X"6A",X"FC",X"16",X"FC",X"7A",X"FF",X"48",X"0A",
		X"7F",X"0A",X"20",X"05",X"6E",X"00",X"59",X"FC",X"6A",X"FC",X"2E",X"FC",X"73",X"FC",X"2B",X"FC",
		X"87",X"FC",X"2E",X"FC",X"E4",X"03",X"29",X"0C",X"4F",X"08",X"94",X"03",X"9F",X"FE",X"2B",X"FC",
		X"68",X"FC",X"3D",X"FC",X"69",X"FC",X"42",X"FC",X"65",X"FC",X"34",X"FD",X"B9",X"06",X"05",X"0C",
		X"10",X"07",X"B0",X"02",X"B1",X"FD",X"38",X"FC",X"5D",X"FC",X"4E",X"FC",X"5D",X"FC",X"59",X"FC",
		X"4B",X"FC",X"F5",X"FD",X"2F",X"08",X"C1",X"0B",X"51",X"06",X"0B",X"02",X"07",X"FD",X"4F",X"FC",
		X"49",X"FC",X"6C",X"FC",X"41",X"FC",X"89",X"FC",X"02",X"FC",X"01",X"00",X"B6",X"0A",X"24",X"0A",
		X"D6",X"04",X"0E",X"00",X"55",X"FC",X"75",X"FC",X"3E",X"FC",X"7B",X"FC",X"41",X"FC",X"81",X"FC",
		X"A0",X"FC",X"E7",X"05",X"0B",X"0C",X"F2",X"06",X"68",X"02",X"4A",X"FD",X"56",X"FC",X"50",X"FC",
		X"74",X"FC",X"41",X"FC",X"96",X"FC",X"02",X"FC",X"94",X"00",X"0A",X"0B",X"C2",X"09",X"92",X"04",
		X"BF",X"FF",X"48",X"FC",X"80",X"FC",X"40",X"FC",X"84",X"FC",X"43",X"FC",X"90",X"FC",X"8A",X"FC",
		X"DF",X"04",X"57",X"0C",X"BE",X"07",X"33",X"03",X"34",X"FE",X"3B",X"FC",X"74",X"FC",X"56",X"FC",
		X"74",X"FC",X"60",X"FC",X"67",X"FC",X"8E",X"FD",X"AF",X"07",X"A4",X"0B",X"52",X"06",X"DF",X"01",
		X"02",X"FD",X"67",X"FC",X"54",X"FC",X"7F",X"FC",X"4D",X"FC",X"9D",X"FC",X"0F",X"FC",X"14",X"01",
		X"50",X"0B",X"59",X"09",X"37",X"04",X"30",X"FF",X"3D",X"FC",X"86",X"FC",X"53",X"FC",X"80",X"FC",
		X"60",X"FC",X"6E",X"FC",X"9E",X"FD",X"2A",X"08",X"59",X"0B",X"D3",X"05",X"42",X"01",X"A1",X"FC",
		X"80",X"FC",X"4D",X"FC",X"91",X"FC",X"48",X"FC",X"AC",X"FC",X"35",X"FC",X"E2",X"02",X"D6",X"0B",
		X"73",X"08",X"AD",X"03",X"96",X"FE",X"34",X"FC",X"8F",X"FC",X"58",X"FC",X"89",X"FC",X"62",X"FC",
		X"7F",X"FC",X"3C",X"FD",X"08",X"07",X"DD",X"0B",X"A1",X"06",X"38",X"02",X"5F",X"FD",X"64",X"FC",
		X"6E",X"FC",X"7C",X"FC",X"6B",X"FC",X"8D",X"FC",X"4A",X"FC",X"6A",X"FF",X"1A",X"0A",X"7D",X"0A",
		X"FE",X"04",X"65",X"00",X"69",X"FC",X"9A",X"FC",X"4D",X"FC",X"A2",X"FC",X"4D",X"FC",X"B3",X"FC",
		X"88",X"FC",X"DF",X"04",X"18",X"0C",X"42",X"07",X"A7",X"02",X"93",X"FD",X"66",X"FC",X"72",X"FC",
		X"87",X"FC",X"6A",X"FC",X"9F",X"FC",X"3F",X"FC",X"B0",X"00",X"39",X"0B",X"8D",X"09",X"2E",X"04",
		X"5F",X"FF",X"49",X"FC",X"A4",X"FC",X"55",X"FC",X"A3",X"FC",X"5B",X"FC",X"A4",X"FC",X"11",X"FD",
		X"9E",X"06",X"13",X"0C",X"9F",X"06",X"3D",X"02",X"59",X"FD",X"74",X"FC",X"77",X"FC",X"89",X"FC",
		X"75",X"FC",X"9B",X"FC",X"51",X"FC",X"16",X"FF",X"A2",X"09",X"A2",X"0A",X"45",X"05",X"B7",X"00",
		X"82",X"FC",X"9E",X"FC",X"5E",X"FC",X"A7",X"FC",X"5B",X"FC",X"BE",X"FC",X"3C",X"FC",X"88",X"02",
		X"BB",X"0B",X"88",X"08",X"92",X"03",X"91",X"FE",X"51",X"FC",X"9E",X"FC",X"70",X"FC",X"98",X"FC",
		X"7F",X"FC",X"79",X"FC",X"1E",X"FE",X"BE",X"08",X"F4",X"0A",X"61",X"05",X"AD",X"00",X"73",X"FC",
		X"AA",X"FC",X"5F",X"FC",X"B1",X"FC",X"5C",X"FC",X"C8",X"FC",X"65",X"FC",X"8F",X"04",X"E9",X"0B",
		X"4D",X"07",X"BA",X"02",X"A4",X"FD",X"70",X"FC",X"89",X"FC",X"90",X"FC",X"81",X"FC",X"A6",X"FC",
		X"55",X"FC",X"D0",X"FE",X"7F",X"09",X"99",X"0A",X"37",X"05",X"9E",X"00",X"8C",X"FC",X"AA",X"FC",
		X"6B",X"FC",X"B1",X"FC",X"6A",X"FC",X"C4",X"FC",X"51",X"FC",X"D1",X"01",X"99",X"0B",X"04",X"09",
		X"F3",X"03",X"29",X"FF",X"58",X"FC",X"B6",X"FC",X"6B",X"FC",X"B8",X"FC",X"6E",X"FC",X"BE",X"FC",
		X"F4",X"FC",X"4D",X"06",X"B9",X"0B",X"7E",X"06",X"FA",X"01",X"26",X"FD",X"95",X"FC",X"7C",X"FC",
		X"AC",X"FC",X"76",X"FC",X"C7",X"FC",X"4D",X"FC",X"65",X"01",X"7A",X"0B",X"CD",X"08",X"AD",X"03",
		X"B4",X"FE",X"61",X"FC",X"B2",X"FC",X"7C",X"FC",X"AF",X"FC",X"87",X"FC",X"9E",X"FC",X"04",X"FE",
		X"85",X"08",X"3F",X"0B",X"75",X"05",X"08",X"01",X"AF",X"FC",X"BB",X"FC",X"6E",X"FC",X"C3",X"FC",
		X"6D",X"FC",X"D8",X"FC",X"4F",X"FC",X"CE",X"01",X"69",X"0B",X"E8",X"08",X"E1",X"03",X"1C",X"FF",
		X"5D",X"FC",X"C6",X"FC",X"73",X"FC",X"C6",X"FC",X"74",X"FC",X"D5",X"FC",X"99",X"FC",X"A2",X"04",
		X"E5",X"0B",X"90",X"07",X"F2",X"02",X"22",X"FE",X"6F",X"FC",X"B7",X"FC",X"85",X"FC",X"BA",X"FC",
		X"85",X"FC",X"C0",X"FC",X"EF",X"FC",X"05",X"06",X"BF",X"0B",X"F3",X"06",X"81",X"02",X"BA",X"FD",
		X"80",X"FC",X"AC",X"FC",X"93",X"FC",X"B3",X"FC",X"95",X"FC",X"B5",X"FC",X"29",X"FD",X"6B",X"06",
		X"B6",X"0B",X"B5",X"06",X"50",X"02",X"88",X"FD",X"91",X"FC",X"A3",X"FC",X"A3",X"FC",X"A6",X"FC",
		X"AC",X"FC",X"96",X"FC",X"1C",X"FE",X"6B",X"08",X"F9",X"0A",X"81",X"05",X"06",X"01",X"B7",X"FC",
		X"C5",X"FC",X"7E",X"FC",X"D2",X"FC",X"79",X"FC",X"F0",X"FC",X"39",X"FC",X"12",X"02",X"6D",X"0B",
		X"59",X"08",X"67",X"03",X"67",X"FE",X"74",X"FC",X"C0",X"FC",X"96",X"FC",X"BA",X"FC",X"A5",X"FC",
		X"A6",X"FC",X"C2",X"FD",X"1D",X"08",X"00",X"0B",X"94",X"05",X"0B",X"01",X"BE",X"FC",X"C4",X"FC",
		X"8C",X"FC",X"CD",X"FC",X"8D",X"FC",X"E1",X"FC",X"62",X"FC",X"FB",X"00",X"FC",X"0A",X"57",X"09",
		X"17",X"04",X"74",X"FF",X"70",X"FC",X"E2",X"FC",X"7E",X"FC",X"E4",X"FC",X"7A",X"FC",X"00",X"FD",
		X"58",X"FC",X"78",X"03",X"A3",X"0B",X"D1",X"07",X"18",X"03",X"2C",X"FE",X"7C",X"FC",X"CB",X"FC",
		X"9C",X"FC",X"C9",X"FC",X"A6",X"FC",X"B9",X"FC",X"D5",X"FD",X"F9",X"07",X"09",X"0B",X"81",X"05",
		X"E6",X"00",X"A8",X"FC",X"D7",X"FC",X"8C",X"FC",X"E0",X"FC",X"89",X"FC",X"FD",X"FC",X"5C",X"FC",
		X"30",X"03",X"99",X"0B",X"98",X"07",X"CD",X"02",X"D5",X"FD",X"9A",X"FC",X"BA",X"FC",X"BB",X"FC",
		X"B4",X"FC",X"D0",X"FC",X"88",X"FC",X"B4",X"FE",X"54",X"09",X"4B",X"0A",X"DD",X"04",X"3F",X"00",
		X"94",X"FC",X"E4",X"FC",X"90",X"FC",X"E6",X"FC",X"8E",X"FC",X"FD",X"FC",X"70",X"FC",X"82",X"02",
		X"7B",X"0B",X"59",X"08",X"6C",X"03",X"9E",X"FE",X"7C",X"FC",X"E5",X"FC",X"96",X"FC",X"E6",X"FC",
		X"96",X"FC",X"F7",X"FC",X"E5",X"FC",X"BC",X"05",X"9C",X"0B",X"89",X"06",X"0A",X"02",X"50",X"FD",
		X"C2",X"FC",X"AC",X"FC",X"D7",X"FC",X"A8",X"FC",X"F1",X"FC",X"6E",X"FC",X"BB",X"FF",X"48",X"0A",
		X"7F",X"09",X"22",X"04",X"57",X"FF",X"81",X"FC",X"F2",X"FC",X"96",X"FC",X"F1",X"FC",X"98",X"FC",
		X"F8",X"FC",X"36",X"FD",X"F9",X"06",X"6B",X"0B",X"BD",X"05",X"3C",X"01",X"D6",X"FC",X"EA",X"FC",
		X"9B",X"FC",X"F0",X"FC",X"9C",X"FC",X"07",X"FD",X"74",X"FC",X"86",X"01",X"4E",X"0B",X"AA",X"08",
		X"8E",X"03",X"CF",X"FE",X"83",X"FC",X"F4",X"FC",X"9C",X"FC",X"F6",X"FC",X"9B",X"FC",X"08",X"FD",
		X"B9",X"FC",X"5D",X"05",X"84",X"0B",X"CA",X"06",X"3D",X"02",X"8F",X"FD",X"AC",X"FC",X"D9",X"FC",
		X"BC",X"FC",X"DF",X"FC",X"BC",X"FC",X"DE",X"FC",X"BF",X"FD",X"8C",X"07",X"2F",X"0B",X"DA",X"05",
		X"7C",X"01",X"21",X"FD",X"D1",X"FC",X"C3",X"FC",X"D3",X"FC",X"CE",X"FC",X"D5",X"FC",X"C5",X"FC",
		X"4E",X"FE",X"5D",X"08",X"F0",X"0A",X"81",X"05",X"33",X"01",X"FD",X"FC",X"DE",X"FC",X"BC",X"FC",
		X"DF",X"FC",X"C8",X"FC",X"E1",X"FC",X"BF",X"FC",X"5A",X"FE",X"52",X"08",X"DD",X"0A",X"83",X"05",
		X"34",X"01",X"FC",X"FC",X"E2",X"FC",X"BE",X"FC",X"E3",X"FC",X"C9",X"FC",X"E5",X"FC",X"BD",X"FC",
		X"33",X"FE",X"2B",X"08",X"D8",X"0A",X"8F",X"05",X"38",X"01",X"F8",X"FC",X"E3",X"FC",X"C2",X"FC",
		X"E5",X"FC",X"CD",X"FC",X"E8",X"FC",X"BC",X"FC",X"19",X"FE",X"11",X"08",X"DE",X"0A",X"9C",X"05",
		X"38",X"01",X"F3",X"FC",X"E6",X"FC",X"CA",X"FC",X"E4",X"FC",X"D4",X"FC",X"E5",X"FC",X"C7",X"FC",
		X"21",X"FE",X"FC",X"07",X"EF",X"0A",X"A2",X"05",X"3E",X"01",X"09",X"FD",X"E4",X"FC",X"CF",X"FC",
		X"E2",X"FC",X"DC",X"FC",X"E1",X"FC",X"D6",X"FC",X"1D",X"FE",X"F0",X"07",X"0A",X"0B",X"A3",X"05",
		X"4B",X"01",X"17",X"FD",X"E7",X"FC",X"D4",X"FC",X"E2",X"FC",X"E3",X"FC",X"DD",X"FC",X"E3",X"FC",
		X"0B",X"FE",X"F1",X"07",X"2E",X"0B",X"9C",X"05",X"5B",X"01",X"1A",X"FD",X"EB",X"FC",X"D2",X"FC",
		X"E9",X"FC",X"E3",X"FC",X"E1",X"FC",X"E6",X"FC",X"00",X"FE",X"C3",X"07",X"16",X"0B",X"AA",X"05",
		X"60",X"01",X"20",X"FD",X"EE",X"FC",X"D5",X"FC",X"ED",X"FC",X"E3",X"FC",X"E7",X"FC",X"E6",X"FC",
		X"E6",X"FD",X"91",X"07",X"02",X"0B",X"B7",X"05",X"67",X"01",X"25",X"FD",X"ED",X"FC",X"D8",X"FC",
		X"EE",X"FC",X"E5",X"FC",X"EB",X"FC",X"E8",X"FC",X"C1",X"FD",X"6B",X"07",X"FC",X"0A",X"C4",X"05",
		X"6C",X"01",X"23",X"FD",X"F1",X"FC",X"DB",X"FC",X"F2",X"FC",X"E7",X"FC",X"F1",X"FC",X"E3",X"FC",
		X"BE",X"FD",X"48",X"07",X"06",X"0B",X"C8",X"05",X"70",X"01",X"16",X"FD",X"FB",X"FC",X"D6",X"FC",
		X"FF",X"FC",X"DD",X"FC",X"05",X"FD",X"C9",X"FC",X"58",X"FE",X"92",X"08",X"62",X"0A",X"E2",X"04",
		X"68",X"00",X"BF",X"FC",X"25",X"FD",X"B8",X"FC",X"27",X"FD",X"B5",X"FC",X"3E",X"FD",X"81",X"FC",
		X"1C",X"02",X"09",X"0B",X"03",X"08",X"F0",X"02",X"49",X"FE",X"B4",X"FC",X"16",X"FD",X"D1",X"FC",
		X"16",X"FD",X"D1",X"FC",X"1A",X"FD",X"7A",X"FD",X"CF",X"06",X"25",X"0B",X"B8",X"05",X"3C",X"01",
		X"FA",X"FC",X"0C",X"FD",X"D8",X"FC",X"0E",X"FD",X"DD",X"FC",X"1A",X"FD",X"B9",X"FC",X"E8",X"FE",
		X"34",X"09",X"FC",X"09",X"A2",X"04",X"25",X"00",X"C2",X"FC",X"24",X"FD",X"C8",X"FC",X"23",X"FD",
		X"CB",X"FC",X"35",X"FD",X"A5",X"FC",X"F6",X"00",X"E7",X"0A",X"C0",X"08",X"77",X"03",X"D1",X"FE",
		X"9D",X"FC",X"36",X"FD",X"BE",X"FC",X"35",X"FD",X"BB",X"FC",X"49",X"FD",X"E5",X"FC",X"D4",X"05",
		X"42",X"0B",X"E8",X"05",X"4F",X"01",X"FE",X"FC",X"1D",X"FD",X"D4",X"FC",X"23",X"FD",X"D4",X"FC",
		X"39",X"FD",X"A5",X"FC",X"2D",X"01",X"1C",X"0B",X"4C",X"08",X"15",X"03",X"5C",X"FE",X"B3",X"FC",
		X"2B",X"FD",X"D2",X"FC",X"2B",X"FD",X"D2",X"FC",X"37",X"FD",X"5B",X"FD",X"DC",X"06",X"23",X"0B",
		X"89",X"05",X"19",X"01",X"EF",X"FC",X"26",X"FD",X"D9",X"FC",X"24",X"FD",X"E1",X"FC",X"30",X"FD",
		X"B9",X"FC",X"74",X"FF",X"7A",X"09",X"A6",X"09",X"3E",X"04",X"BA",X"FF",X"B6",X"FC",X"3C",X"FD",
		X"CA",X"FC",X"3B",X"FD",X"CA",X"FC",X"54",X"FD",X"A5",X"FC",X"8B",X"02",X"56",X"0B",X"9E",X"07",
		X"A2",X"02",X"F9",X"FD",X"D1",X"FC",X"24",X"FD",X"EA",X"FC",X"23",X"FD",X"EE",X"FC",X"1A",X"FD",
		X"25",X"FE",X"62",X"08",X"54",X"0A",X"85",X"04",X"F0",X"FF",X"B3",X"FC",X"43",X"FD",X"CF",X"FC",
		X"41",X"FD",X"D1",X"FC",X"53",X"FD",X"D0",X"FC",X"48",X"04",X"38",X"0B",X"8B",X"06",X"CB",X"01",
		X"67",X"FD",X"0E",X"FD",X"FC",X"FC",X"1A",X"FD",X"FF",X"FC",X"23",X"FD",X"E5",X"FC",X"0C",X"FF",
		X"10",X"09",X"E7",X"09",X"3F",X"04",X"D6",X"FF",X"AA",X"FC",X"55",X"FD",X"C6",X"FC",X"55",X"FD",
		X"C5",X"FC",X"71",X"FD",X"83",X"FC",X"9F",X"01",X"CC",X"0A",X"3C",X"08",X"28",X"03",X"AB",X"FE",
		X"BF",X"FC",X"49",X"FD",X"D4",X"FC",X"50",X"FD",X"CC",X"FC",X"6D",X"FD",X"B3",X"FC",X"6D",X"03",
		X"5A",X"0B",X"63",X"07",X"98",X"02",X"21",X"FE",X"D2",X"FC",X"3E",X"FD",X"E0",X"FC",X"4A",X"FD",
		X"D4",X"FC",X"68",X"FD",X"CD",X"FC",X"0E",X"04",X"60",X"0B",X"1B",X"07",X"6D",X"02",X"02",X"FE",
		X"E1",X"FC",X"3B",X"FD",X"E7",X"FC",X"4A",X"FD",X"DB",X"FC",X"6D",X"FD",X"C2",X"FC",X"F1",X"03",
		X"3B",X"0B",X"21",X"07",X"74",X"02",X"0E",X"FE",X"E4",X"FC",X"3C",X"FD",X"EC",X"FC",X"4B",X"FD",
		X"DC",X"FC",X"72",X"FD",X"A6",X"FC",X"C3",X"03",X"24",X"0B",X"2B",X"07",X"7D",X"02",X"16",X"FE",
		X"E6",X"FC",X"3E",X"FD",X"F1",X"FC",X"4C",X"FD",X"E3",X"FC",X"6E",X"FD",X"BA",X"FC",X"AD",X"03",
		X"11",X"0B",X"3B",X"07",X"7F",X"02",X"1D",X"FE",X"E2",X"FC",X"43",X"FD",X"F2",X"FC",X"50",X"FD",
		X"E5",X"FC",X"6C",X"FD",X"CB",X"FC",X"99",X"03",X"0E",X"0B",X"4D",X"07",X"81",X"02",X"21",X"FE",
		X"DE",X"FC",X"4C",X"FD",X"EF",X"FC",X"55",X"FD",X"E5",X"FC",X"72",X"FD",X"D2",X"FC",X"80",X"03",
		X"1D",X"0B",X"5A",X"07",X"84",X"02",X"22",X"FE",X"DA",X"FC",X"54",X"FD",X"EC",X"FC",X"5C",X"FD",
		X"E3",X"FC",X"7A",X"FD",X"CD",X"FC",X"65",X"03",X"3C",X"0B",X"5F",X"07",X"8B",X"02",X"21",X"FE",
		X"DD",X"FC",X"5A",X"FD",X"ED",X"FC",X"63",X"FD",X"E1",X"FC",X"83",X"FD",X"C2",X"FC",X"47",X"03",
		X"38",X"0B",X"63",X"07",X"94",X"02",X"31",X"FE",X"E4",X"FC",X"58",X"FD",X"F0",X"FC",X"64",X"FD",
		X"E5",X"FC",X"89",X"FD",X"B1",X"FC",X"1C",X"03",X"0D",X"0B",X"69",X"07",X"9D",X"02",X"3C",X"FE",
		X"EB",X"FC",X"55",X"FD",X"F7",X"FC",X"61",X"FD",X"EA",X"FC",X"8A",X"FD",X"A1",X"FC",X"EE",X"02",
		X"F6",X"0A",X"70",X"07",X"A9",X"02",X"42",X"FE",X"F3",X"FC",X"54",X"FD",X"01",X"FD",X"5E",X"FD",
		X"F4",X"FC",X"7F",X"FD",X"BB",X"FC",X"EC",X"02",X"E2",X"0A",X"68",X"07",X"89",X"02",X"28",X"FE",
		X"F9",X"FC",X"55",X"FD",X"04",X"FD",X"60",X"FD",X"F7",X"FC",X"81",X"FD",X"F8",X"FC",X"44",X"05",
		X"21",X"0B",X"D8",X"05",X"4F",X"01",X"24",X"FD",X"4F",X"FD",X"11",X"FD",X"4F",X"FD",X"15",X"FD",
		X"5D",X"FD",X"E7",X"FC",X"69",X"FF",X"BD",X"09",X"EA",X"08",X"6E",X"03",X"D3",X"FE",X"D8",X"FC",
		X"6C",X"FD",X"FD",X"FC",X"6D",X"FD",X"FB",X"FC",X"7E",X"FD",X"41",X"FD",X"5C",X"06",X"CD",X"0A",
		X"EF",X"04",X"68",X"00",X"E7",X"FC",X"7A",X"FD",X"F3",X"FC",X"78",X"FD",X"F0",X"FC",X"97",X"FD",
		X"BC",X"FC",X"9B",X"03",X"E7",X"0A",X"49",X"06",X"5A",X"01",X"31",X"FD",X"56",X"FD",X"14",X"FD",
		X"60",X"FD",X"0F",X"FD",X"7B",X"FD",X"D5",X"FC",X"C7",X"01",X"B1",X"0A",X"31",X"07",X"F8",X"01",
		X"8B",X"FD",X"3B",X"FD",X"2B",X"FD",X"4F",X"FD",X"21",X"FD",X"6A",X"FD",X"E9",X"FC",X"B1",X"00",
		X"78",X"0A",X"C0",X"07",X"53",X"02",X"D6",X"FD",X"2A",X"FD",X"3D",X"FD",X"42",X"FD",X"31",X"FD",
		X"5D",X"FD",X"FB",X"FC",X"1F",X"00",X"47",X"0A",X"0A",X"08",X"81",X"02",X"FB",X"FD",X"22",X"FD",
		X"46",X"FD",X"3F",X"FD",X"38",X"FD",X"59",X"FD",X"06",X"FD",X"EF",X"FF",X"24",X"0A",X"1F",X"08",
		X"8A",X"02",X"02",X"FE",X"21",X"FD",X"49",X"FD",X"3F",X"FD",X"3D",X"FD",X"5B",X"FD",X"0A",X"FD",
		X"01",X"00",X"16",X"0A",X"11",X"08",X"7D",X"02",X"EE",X"FD",X"28",X"FD",X"4A",X"FD",X"45",X"FD",
		X"3C",X"FD",X"62",X"FD",X"05",X"FD",X"41",X"00",X"1D",X"0A",X"E0",X"07",X"60",X"02",X"C6",X"FD",
		X"30",X"FD",X"44",X"FD",X"4D",X"FD",X"38",X"FD",X"6C",X"FD",X"FB",X"FC",X"9F",X"00",X"39",X"0A",
		X"9E",X"07",X"34",X"02",X"B4",X"FD",X"3F",X"FD",X"3E",X"FD",X"58",X"FD",X"30",X"FD",X"79",X"FD",
		X"F1",X"FC",X"D0",X"00",X"43",X"0A",X"9E",X"07",X"49",X"02",X"D1",X"FD",X"34",X"FD",X"52",X"FD",
		X"45",X"FD",X"50",X"FD",X"51",X"FD",X"3A",X"FD",X"DD",X"FE",X"18",X"09",X"42",X"09",X"6E",X"03",
		X"14",X"FF",X"EC",X"FC",X"91",X"FD",X"0C",X"FD",X"91",X"FD",X"05",X"FD",X"AD",X"FD",X"F1",X"FC",
		X"4C",X"04",X"01",X"0B",X"07",X"06",X"51",X"01",X"61",X"FD",X"5F",X"FD",X"3A",X"FD",X"60",X"FD",
		X"43",X"FD",X"67",X"FD",X"2B",X"FD",X"29",X"FF",X"4F",X"09",X"0E",X"09",X"45",X"03",X"EC",X"FE",
		X"F7",X"FC",X"8F",X"FD",X"17",X"FD",X"8C",X"FD",X"16",X"FD",X"9C",X"FD",X"54",X"FD",X"EE",X"05",
		X"6A",X"0A",X"EE",X"04",X"2F",X"00",X"F0",X"FC",X"99",X"FD",X"11",X"FD",X"98",X"FD",X"0A",X"FD",
		X"BC",X"FD",X"B7",X"FC",X"C6",X"02",X"E7",X"0A",X"90",X"06",X"AE",X"01",X"89",X"FD",X"59",X"FD",
		X"4C",X"FD",X"5C",X"FD",X"54",X"FD",X"5E",X"FD",X"48",X"FD",X"5E",X"FE",X"77",X"08",X"96",X"09",
		X"E6",X"03",X"86",X"FF",X"EC",X"FC",X"9F",X"FD",X"16",X"FD",X"98",X"FD",X"18",X"FD",X"AE",X"FD",
		X"E2",X"FC",X"98",X"01",X"4A",X"0A",X"A5",X"07",X"6B",X"02",X"2B",X"FE",X"21",X"FD",X"81",X"FD",
		X"32",X"FD",X"89",X"FD",X"2A",X"FD",X"9C",X"FD",X"68",X"FD",X"F4",X"05",X"7A",X"0A",X"F9",X"04",
		X"5E",X"00",X"12",X"FD",X"98",X"FD",X"26",X"FD",X"93",X"FD",X"26",X"FD",X"AA",X"FD",X"EB",X"FC",
		X"A3",X"01",X"5B",X"0A",X"38",X"07",X"F9",X"01",X"B5",X"FD",X"4C",X"FD",X"65",X"FD",X"5B",X"FD",
		X"67",X"FD",X"61",X"FD",X"56",X"FD",X"7B",X"FE",X"51",X"08",X"6C",X"09",X"C1",X"03",X"54",X"FF",
		X"F6",X"FC",X"AD",X"FD",X"1C",X"FD",X"A8",X"FD",X"18",X"FD",X"C6",X"FD",X"DB",X"FC",X"93",X"02",
		X"7A",X"0A",X"03",X"07",X"EA",X"01",X"DA",X"FD",X"3A",X"FD",X"86",X"FD",X"39",X"FD",X"9A",X"FD",
		X"29",X"FD",X"BD",X"FD",X"28",X"FD",X"89",X"05",X"D8",X"0A",X"71",X"05",X"F7",X"00",X"55",X"FD",
		X"77",X"FD",X"5A",X"FD",X"66",X"FD",X"73",X"FD",X"54",X"FD",X"88",X"FD",X"DE",X"FD",X"E0",X"06",
		X"4B",X"0A",X"D4",X"04",X"6E",X"00",X"37",X"FD",X"88",X"FD",X"52",X"FD",X"72",X"FD",X"6C",X"FD",
		X"62",X"FD",X"7B",X"FD",X"1B",X"FE",X"55",X"07",X"26",X"0A",X"A4",X"04",X"4D",X"00",X"30",X"FD",
		X"8E",X"FD",X"52",X"FD",X"76",X"FD",X"6E",X"FD",X"63",X"FD",X"84",X"FD",X"F8",X"FD",X"5D",X"07",
		X"49",X"0A",X"9C",X"04",X"5D",X"00",X"22",X"FD",X"9A",X"FD",X"4B",X"FD",X"81",X"FD",X"66",X"FD",
		X"6E",X"FD",X"7C",X"FD",X"DD",X"FD",X"25",X"07",X"2F",X"0A",X"A9",X"04",X"61",X"00",X"18",X"FD",
		X"A4",X"FD",X"45",X"FD",X"8E",X"FD",X"5F",X"FD",X"7F",X"FD",X"6B",X"FD",X"04",X"FE",X"67",X"07",
		X"FE",X"09",X"47",X"04",X"0B",X"00",X"02",X"FD",X"C0",X"FD",X"2D",X"FD",X"B0",X"FD",X"38",X"FD",
		X"BB",X"FD",X"10",X"FD",X"49",X"00",X"82",X"09",X"41",X"08",X"A6",X"02",X"75",X"FE",X"1E",X"FD",
		X"B2",X"FD",X"37",X"FD",X"B3",X"FD",X"32",X"FD",X"CC",X"FD",X"44",X"FD",X"41",X"05",X"62",X"0A",
		X"38",X"05",X"7C",X"00",X"39",X"FD",X"A0",X"FD",X"53",X"FD",X"93",X"FD",X"61",X"FD",X"93",X"FD",
		X"4E",X"FD",X"18",X"FF",X"0C",X"09",X"0A",X"09",X"4C",X"03",X"27",X"FF",X"13",X"FD",X"C1",X"FD",
		X"37",X"FD",X"BB",X"FD",X"36",X"FD",X"D1",X"FD",X"01",X"FD",X"5D",X"01",X"FD",X"09",X"AA",X"07",
		X"58",X"02",X"4A",X"FE",X"35",X"FD",X"B1",X"FD",X"3F",X"FD",X"BE",X"FD",X"2E",X"FD",X"EA",X"FD",
		X"E9",X"FC",X"70",X"04",X"D2",X"0A",X"7A",X"05",X"E1",X"00",X"55",X"FD",X"A3",X"FD",X"58",X"FD",
		X"9C",X"FD",X"62",X"FD",X"A5",X"FD",X"3D",X"FD",X"52",X"FF",X"88",X"09",X"6C",X"08",X"A9",X"02",
		X"82",X"FE",X"38",X"FD",X"B0",X"FD",X"51",X"FD",X"B0",X"FD",X"4F",X"FD",X"BE",X"FD",X"A2",X"FD",
		X"69",X"06",X"EB",X"09",X"24",X"04",X"9D",X"FF",X"0D",X"FD",X"D2",X"FD",X"35",X"FD",X"D1",X"FD",
		X"2D",X"FD",X"F6",X"FD",X"E1",X"FC",X"35",X"04",X"BF",X"0A",X"2B",X"05",X"75",X"00",X"2A",X"FD",
		X"C9",X"FD",X"42",X"FD",X"C6",X"FD",X"3C",X"FD",X"E6",X"FD",X"F6",X"FC",X"B0",X"02",X"72",X"0A",
		X"FF",X"05",X"F3",X"00",X"64",X"FD",X"AF",X"FD",X"59",X"FD",X"B4",X"FD",X"53",X"FD",X"D3",X"FD",
		X"0F",X"FD",X"C8",X"01",X"3B",X"0A",X"76",X"06",X"3E",X"01",X"85",X"FD",X"A2",X"FD",X"67",X"FD",
		X"AC",X"FD",X"5E",X"FD",X"C8",X"FD",X"1D",X"FD",X"57",X"01",X"1B",X"0A",X"AE",X"06",X"60",X"01",
		X"93",X"FD",X"A0",X"FD",X"6A",X"FD",X"AB",X"FD",X"63",X"FD",X"C9",X"FD",X"21",X"FD",X"39",X"01",
		X"13",X"0A",X"B8",X"06",X"5E",X"01",X"97",X"FD",X"A2",X"FD",X"6E",X"FD",X"AD",X"FD",X"66",X"FD",
		X"CE",X"FD",X"1E",X"FD",X"4F",X"01",X"27",X"0A",X"9B",X"06",X"4D",X"01",X"89",X"FD",X"AC",X"FD",
		X"68",X"FD",X"B7",X"FD",X"5D",X"FD",X"DA",X"FD",X"12",X"FD",X"7F",X"01",X"40",X"0A",X"8C",X"06",
		X"47",X"01",X"90",X"FD",X"A7",X"FD",X"74",X"FD",X"AB",X"FD",X"75",X"FD",X"BC",X"FD",X"4A",X"FD",
		X"FD",X"FF",X"52",X"09",X"E2",X"07",X"44",X"02",X"3F",X"FE",X"58",X"FD",X"BC",X"FD",X"69",X"FD",
		X"C2",X"FD",X"61",X"FD",X"D6",X"FD",X"8B",X"FD",X"D3",X"05",X"FD",X"09",X"97",X"04",X"0E",X"00",
		X"39",X"FD",X"D0",X"FD",X"60",X"FD",X"C5",X"FD",X"66",X"FD",X"D4",X"FD",X"38",X"FD",X"6C",X"00",
		X"80",X"09",X"AE",X"07",X"27",X"02",X"2E",X"FE",X"63",X"FD",X"BA",X"FD",X"73",X"FD",X"C0",X"FD",
		X"6E",X"FD",X"CA",X"FD",X"CD",X"FD",X"BD",X"06",X"9E",X"09",X"CE",X"03",X"6E",X"FF",X"33",X"FD",
		X"E0",X"FD",X"54",X"FD",X"DF",X"FD",X"4C",X"FD",X"05",X"FE",X"08",X"FD",X"E0",X"03",X"67",X"0A",
		X"1B",X"05",X"58",X"00",X"35",X"FD",X"E1",X"FD",X"59",X"FD",X"DE",X"FD",X"54",X"FD",X"FF",X"FD",
		X"00",X"FD",X"34",X"02",X"74",X"0A",X"0E",X"06",X"EF",X"00",X"6B",X"FD",X"C8",X"FD",X"71",X"FD",
		X"C9",X"FD",X"6E",X"FD",X"E4",X"FD",X"29",X"FD",X"2A",X"01",X"01",X"0A",X"AD",X"06",X"4E",X"01",
		X"A2",X"FD",X"B2",X"FD",X"85",X"FD",X"BB",X"FD",X"80",X"FD",X"D5",X"FD",X"44",X"FD",X"9B",X"00",
		X"BE",X"09",X"FF",X"06",X"7F",X"01",X"BD",X"FD",X"A9",X"FD",X"91",X"FD",X"B4",X"FD",X"8A",X"FD",
		X"CD",X"FD",X"51",X"FD",X"62",X"00",X"A3",X"09",X"1A",X"07",X"8D",X"01",X"C4",X"FD",X"AA",X"FD",
		X"92",X"FD",X"B7",X"FD",X"8B",X"FD",X"CF",X"FD",X"55",X"FD",X"32",X"00",X"77",X"09",X"61",X"07",
		X"C5",X"01",X"FC",X"FD",X"8E",X"FD",X"B3",X"FD",X"95",X"FD",X"B9",X"FD",X"95",X"FD",X"BA",X"FD",
		X"3A",X"FE",X"C2",X"07",X"1A",X"09",X"21",X"03",X"EF",X"FE",X"39",X"FD",X"F4",X"FD",X"5C",X"FD",
		X"F4",X"FD",X"55",X"FD",X"19",X"FE",X"06",X"FD",X"B1",X"02",X"5D",X"0A",X"19",X"06",X"19",X"01",
		X"A4",X"FD",X"AE",X"FD",X"A8",X"FD",X"A1",X"FD",X"BF",X"FD",X"8F",X"FD",X"D7",X"FD",X"BE",X"FD",
		X"21",X"06",X"D1",X"09",X"5D",X"04",X"FF",X"FF",X"56",X"FD",X"DF",X"FD",X"84",X"FD",X"C9",X"FD",
		X"9A",X"FD",X"BD",X"FD",X"A1",X"FD",X"67",X"FE",X"E4",X"07",X"4A",X"09",X"7D",X"03",X"74",X"FF",
		X"48",X"FD",X"F0",X"FD",X"76",X"FD",X"DB",X"FD",X"8A",X"FD",X"D7",X"FD",X"82",X"FD",X"D8",X"FE",
		X"7E",X"08",X"F5",X"08",X"34",X"03",X"43",X"FF",X"4B",X"FD",X"F3",X"FD",X"76",X"FD",X"E1",X"FD",
		X"86",X"FD",X"DF",X"FD",X"79",X"FD",X"04",X"FF",X"5D",X"08",X"DF",X"08",X"3C",X"03",X"44",X"FF",
		X"4C",X"FD",X"F6",X"FD",X"75",X"FD",X"E6",X"FD",X"84",X"FD",X"E7",X"FD",X"75",X"FD",X"20",X"FF",
		X"2E",X"08",X"D6",X"08",X"23",X"03",X"35",X"FF",X"43",X"FD",X"06",X"FE",X"68",X"FD",X"FE",X"FD",
		X"6A",X"FD",X"13",X"FE",X"31",X"FD",X"64",X"00",X"9E",X"09",X"8C",X"07",X"E4",X"01",X"41",X"FE",
		X"75",X"FD",X"EE",X"FD",X"7A",X"FD",X"FC",X"FD",X"6A",X"FD",X"23",X"FE",X"3A",X"FD",X"3B",X"05",
		X"27",X"0A",X"6E",X"04",X"F4",X"FF",X"53",X"FD",X"FA",X"FD",X"80",X"FD",X"EB",X"FD",X"87",X"FD",
		X"F7",X"FD",X"5F",X"FD",X"E7",X"FF",X"2E",X"09",X"DF",X"07",X"3B",X"02",X"7B",X"FE",X"72",X"FD",
		X"F2",X"FD",X"80",X"FD",X"FA",X"FD",X"74",X"FD",X"1E",X"FE",X"36",X"FD",X"BB",X"02",X"00",X"0A",
		X"21",X"06",X"1A",X"01",X"C2",X"FD",X"B5",X"FD",X"C9",X"FD",X"A6",X"FD",X"E0",X"FD",X"92",X"FD",
		X"04",X"FE",X"7B",X"FD",X"33",X"05",X"F5",X"09",X"81",X"04",X"17",X"00",X"65",X"FD",X"FA",X"FD",
		X"8C",X"FD",X"ED",X"FD",X"95",X"FD",X"F4",X"FD",X"74",X"FD",X"C8",X"FF",X"D2",X"08",X"D6",X"07",
		X"14",X"02",X"61",X"FE",X"83",X"FD",X"F2",X"FD",X"8F",X"FD",X"F8",X"FD",X"84",X"FD",X"13",X"FE",
		X"84",X"FD",X"E1",X"05",X"B8",X"09",X"CD",X"03",X"6D",X"FF",X"51",X"FD",X"11",X"FE",X"7C",X"FD",
		X"0C",X"FE",X"75",X"FD",X"2C",X"FE",X"2F",X"FD",X"F5",X"02",X"FF",X"09",X"3B",X"05",X"54",X"00",
		X"7C",X"FD",X"F8",X"FD",X"93",X"FD",X"F8",X"FD",X"8D",X"FD",X"17",X"FE",X"3D",X"FD",X"3A",X"01",
		X"01",X"0A",X"37",X"06",X"E7",X"00",X"A6",X"FD",X"E0",X"FD",X"AB",X"FD",X"DD",X"FD",X"AF",X"FD",
		X"EC",X"FD",X"8A",X"FD",X"BA",X"FF",X"E6",X"08",X"A2",X"07",X"E8",X"01",X"3C",X"FE",X"9C",X"FD",
		X"EA",X"FD",X"A4",X"FD",X"F5",X"FD",X"96",X"FD",X"15",X"FE",X"85",X"FD",X"4F",X"05",X"D2",X"09",
		X"38",X"04",X"DF",X"FF",X"66",X"FD",X"0F",X"FE",X"90",X"FD",X"FE",X"FD",X"9C",X"FD",X"00",X"FE",
		X"8A",X"FD",X"70",X"FF",X"43",X"08",X"4D",X"08",X"7B",X"02",X"CE",X"FE",X"66",X"FD",X"1B",X"FE",
		X"7F",X"FD",X"1E",X"FE",X"79",X"FD",X"38",X"FE",X"37",X"FD",X"31",X"01",X"85",X"09",X"17",X"07",
		X"A7",X"01",X"4D",X"FE",X"8F",X"FD",X"08",X"FE",X"8E",X"FD",X"19",X"FE",X"7C",X"FD",X"41",X"FE",
		X"28",X"FD",X"14",X"02",X"EE",X"09",X"7F",X"06",X"5B",X"01",X"15",X"FE",X"A9",X"FD",X"F6",X"FD",
		X"9F",X"FD",X"0C",X"FE",X"8D",X"FD",X"37",X"FE",X"3A",X"FD",X"3E",X"02",X"DD",X"09",X"63",X"06",
		X"5E",X"01",X"0D",X"FE",X"B5",X"FD",X"EF",X"FD",X"AB",X"FD",X"04",X"FE",X"97",X"FD",X"2A",X"FE",
		X"4F",X"FD",X"22",X"02",X"BC",X"09",X"6F",X"06",X"66",X"01",X"0E",X"FE",X"B7",X"FD",X"F2",X"FD",
		X"AF",X"FD",X"05",X"FE",X"9A",X"FD",X"2E",X"FE",X"51",X"FD",X"70",X"02",X"C5",X"09",X"10",X"06",
		X"06",X"01",X"E6",X"FD",X"CD",X"FD",X"E6",X"FD",X"BC",X"FD",X"FE",X"FD",X"A4",X"FD",X"2A",X"FE",
		X"74",X"FD",X"5D",X"05",X"B6",X"09",X"EE",X"03",X"AB",X"FF",X"6D",X"FD",X"20",X"FE",X"9A",X"FD",
		X"14",X"FE",X"9E",X"FD",X"28",X"FE",X"61",X"FD",X"7C",X"00",X"71",X"09",X"BE",X"06",X"40",X"01",
		X"F8",X"FD",X"D1",X"FD",X"E1",X"FD",X"D1",X"FD",X"EA",X"FD",X"CF",X"FD",X"EA",X"FD",X"74",X"FE",
		X"49",X"07",X"93",X"08",X"81",X"02",X"AF",X"FE",X"8C",X"FD",X"1C",X"FE",X"A0",X"FD",X"1F",X"FE",
		X"95",X"FD",X"42",X"FE",X"62",X"FD",X"52",X"05",X"8B",X"09",X"87",X"03",X"59",X"FF",X"78",X"FD",
		X"28",X"FE",X"9B",X"FD",X"23",X"FE",X"94",X"FD",X"44",X"FE",X"50",X"FD",X"A7",X"02",X"C1",X"09",
		X"6E",X"05",X"70",X"00",X"AC",X"FD",X"00",X"FE",X"C9",X"FD",X"F1",X"FD",X"D9",X"FD",X"EB",X"FD",
		X"DA",X"FD",X"AC",X"FE",X"60",X"07",X"9B",X"08",X"BB",X"02",X"F3",X"FE",X"86",X"FD",X"27",X"FE",
		X"A2",X"FD",X"28",X"FE",X"9C",X"FD",X"43",X"FE",X"56",X"FD",X"35",X"01",X"82",X"09",X"6B",X"06",
		X"0B",X"01",X"FA",X"FD",X"D5",X"FD",X"F8",X"FD",X"CC",X"FD",X"07",X"FE",X"BE",X"FD",X"21",X"FE",
		X"D3",X"FD",X"52",X"06",X"18",X"09",X"0E",X"03",X"1C",X"FF",X"87",X"FD",X"2C",X"FE",X"A5",X"FD",
		X"2B",X"FE",X"9E",X"FD",X"4C",X"FE",X"5A",X"FD",X"12",X"03",X"B6",X"09",X"F5",X"04",X"1D",X"00",
		X"96",X"FD",X"1C",X"FE",X"BD",X"FD",X"11",X"FE",X"C7",X"FD",X"16",X"FE",X"AD",X"FD",X"81",X"FF",
		X"67",X"08",X"C9",X"07",X"EA",X"01",X"70",X"FE",X"A8",X"FD",X"21",X"FE",X"AF",X"FD",X"2D",X"FE",
		X"A1",X"FD",X"52",X"FE",X"5D",X"FD",X"D1",X"02",X"A5",X"09",X"7C",X"05",X"8A",X"00",X"D3",X"FD",
		X"F4",X"FD",X"EE",X"FD",X"E2",X"FD",X"05",X"FE",X"CE",X"FD",X"25",X"FE",X"CF",X"FD",X"2C",X"06",
		X"52",X"09",X"3B",X"03",X"4E",X"FF",X"7D",X"FD",X"3E",X"FE",X"A6",X"FD",X"38",X"FE",X"A5",X"FD",
		X"52",X"FE",X"5A",X"FD",X"52",X"01",X"A1",X"09",X"0A",X"06",X"BC",X"00",X"DE",X"FD",X"F7",X"FD",
		X"E9",X"FD",X"F3",X"FD",X"F2",X"FD",X"F4",X"FD",X"EB",X"FD",X"D1",X"FE",X"BC",X"07",X"F9",X"07",
		X"EC",X"01",X"6B",X"FE",X"BD",X"FD",X"1E",X"FE",X"C5",X"FD",X"24",X"FE",X"BC",X"FD",X"3E",X"FE",
		X"BE",X"FD",X"1A",X"06",X"23",X"09",X"D8",X"02",X"02",X"FF",X"94",X"FD",X"3C",X"FE",X"AF",X"FD",
		X"3B",X"FE",X"A7",X"FD",X"5E",X"FE",X"79",X"FD",X"D0",X"04",X"86",X"09",X"89",X"03",X"55",X"FF",
		X"8E",X"FD",X"40",X"FE",X"B1",X"FD",X"3E",X"FE",X"A9",X"FD",X"60",X"FE",X"68",X"FD",X"E5",X"03",
		X"94",X"09",X"FD",X"03",X"81",X"FF",X"8F",X"FD",X"41",X"FE",X"B4",X"FD",X"3F",X"FE",X"AD",X"FD",
		X"62",X"FE",X"64",X"FD",X"76",X"03",X"99",X"09",X"30",X"04",X"98",X"FF",X"91",X"FD",X"3F",X"FE",
		X"B8",X"FD",X"3D",X"FE",X"B1",X"FD",X"61",X"FE",X"66",X"FD",X"0C",X"03",X"97",X"09",X"8C",X"04",
		X"CB",X"FF",X"96",X"FD",X"3C",X"FE",X"C2",X"FD",X"35",X"FE",X"C3",X"FD",X"4B",X"FE",X"84",X"FD",
		X"8A",X"00",X"36",X"09",X"86",X"06",X"F1",X"00",X"14",X"FE",X"E7",X"FD",X"15",X"FE",X"DF",X"FD",
		X"28",X"FE",X"CB",X"FD",X"4C",X"FE",X"AA",X"FD",X"8A",X"05",X"5C",X"09",X"68",X"03",X"6B",X"FF",
		X"97",X"FD",X"45",X"FE",X"C1",X"FD",X"3B",X"FE",X"C5",X"FD",X"4C",X"FE",X"90",X"FD",X"77",X"00",
		X"39",X"09",X"A0",X"06",X"FE",X"00",X"1B",X"FE",X"EC",X"FD",X"15",X"FE",X"E8",X"FD",X"23",X"FE",
		X"DF",X"FD",X"38",X"FE",X"F2",X"FD",X"77",X"06",X"A7",X"08",X"75",X"02",X"D0",X"FE",X"B2",X"FD",
		X"42",X"FE",X"C4",X"FD",X"46",X"FE",X"B9",X"FD",X"6B",X"FE",X"7C",X"FD",X"5F",X"04",X"88",X"09",
		X"AF",X"03",X"74",X"FF",X"9E",X"FD",X"4E",X"FE",X"C1",X"FD",X"4A",X"FE",X"BA",X"FD",X"6C",X"FE",
		X"6C",X"FD",X"9C",X"02",X"76",X"09",X"A5",X"04",X"C8",X"FF",X"A7",X"FD",X"45",X"FE",X"CF",X"FD",
		X"40",X"FE",X"C6",X"FD",X"62",X"FE",X"75",X"FD",X"80",X"01",X"5F",X"09",X"48",X"05",X"1F",X"00",
		X"BE",X"FD",X"36",X"FE",X"E2",X"FD",X"2D",X"FE",X"E8",X"FD",X"37",X"FE",X"C3",X"FD",X"CC",X"FF",
		X"D3",X"08",X"14",X"07",X"30",X"01",X"47",X"FE",X"DE",X"FD",X"34",X"FE",X"DA",X"FD",X"45",X"FE",
		X"C6",X"FD",X"6E",X"FE",X"8C",X"FD",X"DF",X"04",X"8E",X"09",X"B9",X"03",X"95",X"FF",X"A8",X"FD",
		X"49",X"FE",X"D9",X"FD",X"39",X"FE",X"E5",X"FD",X"3B",X"FE",X"D3",X"FD",X"83",X"FF",X"2A",X"08",
		X"74",X"07",X"81",X"01",X"5C",X"FE",X"D8",X"FD",X"3F",X"FE",X"D8",X"FD",X"4B",X"FE",X"C8",X"FD",
		X"71",X"FE",X"8F",X"FD",X"AA",X"04",X"6F",X"09",X"88",X"03",X"6B",X"FF",X"AC",X"FD",X"55",X"FE",
		X"CF",X"FD",X"51",X"FE",X"CA",X"FD",X"70",X"FE",X"78",X"FD",X"5C",X"01",X"50",X"09",X"83",X"05",
		X"52",X"00",X"E7",X"FD",X"27",X"FE",X"02",X"FE",X"1A",X"FE",X"11",X"FE",X"11",X"FE",X"1D",X"FE",
		X"6E",X"FE",X"D3",X"06",X"55",X"08",X"39",X"02",X"D5",X"FE",X"BC",X"FD",X"5A",X"FE",X"CE",X"FD",
		X"5B",X"FE",X"C8",X"FD",X"7B",X"FE",X"80",X"FD",X"22",X"01",X"3D",X"09",X"36",X"06",X"C5",X"00",
		X"2F",X"FE",X"F2",X"FD",X"3C",X"FE",X"E4",X"FD",X"55",X"FE",X"CB",X"FD",X"84",X"FE",X"78",X"FD",
		X"24",X"03",X"55",X"09",X"EA",X"04",X"18",X"00",X"F8",X"FD",X"17",X"FE",X"24",X"FE",X"FC",X"FD",
		X"44",X"FE",X"DF",X"FD",X"74",X"FE",X"A4",X"FD",X"2B",X"04",X"41",X"09",X"5A",X"04",X"D3",X"FF",
		X"E7",X"FD",X"27",X"FE",X"1A",X"FE",X"09",X"FE",X"3C",X"FE",X"E9",X"FD",X"6E",X"FE",X"AC",X"FD",
		X"49",X"04",X"43",X"09",X"40",X"04",X"D5",X"FF",X"E2",X"FD",X"2B",X"FE",X"18",X"FE",X"0D",X"FE",
		X"3C",X"FE",X"ED",X"FD",X"72",X"FE",X"98",X"FD",X"1B",X"04",X"5F",X"09",X"3C",X"04",X"E8",X"FF",
		X"DC",X"FD",X"38",X"FE",X"11",X"FE",X"19",X"FE",X"36",X"FE",X"F5",X"FD",X"6D",X"FE",X"98",X"FD",
		X"09",X"04",X"81",X"09",X"2F",X"04",X"F1",X"FF",X"CB",X"FD",X"4B",X"FE",X"02",X"FE",X"2D",X"FE",
		X"21",X"FE",X"10",X"FE",X"4B",X"FE",X"F3",X"FD",X"5C",X"05",X"F5",X"08",X"FC",X"02",X"42",X"FF",
		X"BE",X"FD",X"68",X"FE",X"E1",X"FD",X"5E",X"FE",X"E8",X"FD",X"6B",X"FE",X"BB",X"FD",X"22",X"00",
		X"A3",X"08",X"90",X"06",X"CE",X"00",X"3B",X"FE",X"0A",X"FE",X"3C",X"FE",X"05",X"FE",X"4A",X"FE",
		X"F6",X"FD",X"69",X"FE",X"DA",X"FD",X"AB",X"05",X"A4",X"08",X"73",X"02",X"D2",X"FE",X"D0",X"FD",
		X"68",X"FE",X"E1",X"FD",X"6C",X"FE",X"D7",X"FD",X"94",X"FE",X"86",X"FD",X"6A",X"03",X"74",X"09",
		X"DB",X"03",X"87",X"FF",X"CF",X"FD",X"63",X"FE",X"EF",X"FD",X"5D",X"FE",X"EB",X"FD",X"7B",X"FE",
		X"A2",X"FD",X"33",X"01",X"06",X"09",X"5C",X"05",X"23",X"00",X"EB",X"FD",X"45",X"FE",X"14",X"FE",
		X"34",X"FE",X"23",X"FE",X"2C",X"FE",X"2D",X"FE",X"AB",X"FE",X"ED",X"06",X"04",X"08",X"E9",X"01",
		X"B1",X"FE",X"DE",X"FD",X"69",X"FE",X"EC",X"FD",X"6D",X"FE",X"E2",X"FD",X"8C",X"FE",X"98",X"FD",
		X"55",X"01",X"F9",X"08",X"A5",X"05",X"5B",X"00",X"13",X"FE",X"2C",X"FE",X"33",X"FE",X"19",X"FE",
		X"4A",X"FE",X"05",X"FE",X"70",X"FE",X"DC",X"FD",X"54",X"05",X"D3",X"08",X"B3",X"02",X"13",X"FF",
		X"D4",X"FD",X"72",X"FE",X"EB",X"FD",X"71",X"FE",X"E5",X"FD",X"92",X"FE",X"92",X"FD",X"71",X"01",
		X"09",X"09",X"1E",X"05",X"F6",X"FF",X"EF",X"FD",X"4E",X"FE",X"18",X"FE",X"41",X"FE",X"24",X"FE",
		X"40",X"FE",X"1B",X"FE",X"20",X"FF",X"A4",X"07",X"62",X"07",X"58",X"01",X"80",X"FE",X"FA",X"FD",
		X"64",X"FE",X"FC",X"FD",X"70",X"FE",X"E9",X"FD",X"99",X"FE",X"9A",X"FD",X"06",X"03",X"25",X"09",
		X"6E",X"04",X"C0",X"FF",X"F1",X"FD",X"50",X"FE",X"24",X"FE",X"34",X"FE",X"41",X"FE",X"1E",X"FE",
		X"64",X"FE",X"0D",X"FE",X"C1",X"05",X"B4",X"08",X"BA",X"02",X"27",X"FF",X"E3",X"FD",X"6A",X"FE",
		X"09",X"FE",X"57",X"FE",X"1D",X"FE",X"4E",X"FE",X"27",X"FE",X"C4",X"FE",X"F2",X"06",X"F3",X"07",
		X"02",X"02",X"D0",X"FE",X"F0",X"FD",X"6B",X"FE",X"09",X"FE",X"62",X"FE",X"12",X"FE",X"5F",X"FE",
		X"0C",X"FE",X"25",X"FF",X"5C",X"07",X"A4",X"07",X"B8",X"01",X"B9",X"FE",X"F2",X"FD",X"73",X"FE",
		X"FE",X"FD",X"74",X"FE",X"FD",X"FD",X"85",X"FE",X"D3",X"FD",X"50",X"00",X"56",X"08",X"7C",X"06",
		X"C3",X"00",X"4F",X"FE",X"17",X"FE",X"61",X"FE",X"0A",X"FE",X"75",X"FE",X"F5",X"FD",X"A4",X"FE",
		X"9C",X"FD",X"D0",X"03",X"FB",X"08",X"77",X"03",X"49",X"FF",X"E7",X"FD",X"73",X"FE",X"0C",X"FE",
		X"6B",X"FE",X"10",X"FE",X"74",X"FE",X"ED",X"FD",X"E4",X"FF",X"25",X"08",X"88",X"06",X"BF",X"00",
		X"4C",X"FE",X"21",X"FE",X"60",X"FE",X"12",X"FE",X"75",X"FE",X"FB",X"FD",X"A8",X"FE",X"97",X"FD",
		X"44",X"03",X"1E",X"09",X"0F",X"04",X"A3",X"FF",X"02",X"FE",X"5E",X"FE",X"2F",X"FE",X"46",X"FE",
		X"48",X"FE",X"2F",X"FE",X"6B",X"FE",X"31",X"FE",X"92",X"05",X"89",X"08",X"92",X"02",X"0F",X"FF",
		X"E8",X"FD",X"82",X"FE",X"05",X"FE",X"7C",X"FE",X"0A",X"FE",X"88",X"FE",X"E5",X"FD",X"DF",X"FF",
		X"23",X"08",X"78",X"06",X"96",X"00",X"44",X"FE",X"2D",X"FE",X"60",X"FE",X"1E",X"FE",X"73",X"FE",
		X"0A",X"FE",X"9C",X"FE",X"C8",X"FD",X"E5",X"04",X"96",X"08",X"85",X"02",X"F7",X"FE",X"F6",X"FD",
		X"83",X"FE",X"0A",X"FE",X"85",X"FE",X"FF",X"FD",X"A8",X"FE",X"AE",X"FD",X"5C",X"02",X"48",X"09",
		X"26",X"04",X"9A",X"FF",X"FE",X"FD",X"75",X"FE",X"1C",X"FE",X"71",X"FE",X"1B",X"FE",X"87",X"FE",
		X"E4",X"FD",X"6C",X"00",X"93",X"08",X"6A",X"05",X"15",X"00",X"1F",X"FE",X"5D",X"FE",X"37",X"FE",
		X"5A",X"FE",X"3B",X"FE",X"63",X"FE",X"1D",X"FE",X"73",X"FF",X"E1",X"07",X"83",X"06",X"90",X"00",
		X"44",X"FE",X"3A",X"FE",X"5D",X"FE",X"30",X"FE",X"6E",X"FE",X"20",X"FE",X"90",X"FE",X"04",X"FE",
		X"4F",X"05",X"68",X"08",X"55",X"02",X"FA",X"FE",X"FD",X"FD",X"88",X"FE",X"13",X"FE",X"85",X"FE",
		X"13",X"FE",X"99",X"FE",X"E0",X"FD",X"43",X"00",X"4E",X"08",X"10",X"06",X"74",X"00",X"44",X"FE",
		X"3E",X"FE",X"66",X"FE",X"2D",X"FE",X"7C",X"FE",X"16",X"FE",X"A7",X"FE",X"C4",X"FD",X"24",X"04",
		X"CD",X"08",X"FC",X"02",X"17",X"FF",X"FE",X"FD",X"8A",X"FE",X"1A",X"FE",X"84",X"FE",X"18",X"FE",
		X"9B",X"FE",X"DC",X"FD",X"74",X"00",X"7C",X"08",X"75",X"05",X"17",X"00",X"2F",X"FE",X"59",X"FE",
		X"4E",X"FE",X"4E",X"FE",X"5A",X"FE",X"4B",X"FE",X"5B",X"FE",X"DF",X"FE",X"60",X"07",X"3A",X"07",
		X"D9",X"00",X"7B",X"FE",X"2D",X"FE",X"77",X"FE",X"2C",X"FE",X"81",X"FE",X"20",X"FE",X"9D",X"FE",
		X"14",X"FE",X"BF",X"05",X"01",X"08",X"A0",X"01",X"BC",X"FE",X"19",X"FE",X"88",X"FE",X"20",X"FE",
		X"92",X"FE",X"11",X"FE",X"B8",X"FE",X"BE",X"FD",X"AA",X"04",X"66",X"08",X"22",X"02",X"E2",X"FE",
		X"10",X"FE",X"8F",X"FE",X"1D",X"FE",X"96",X"FE",X"10",X"FE",X"BD",X"FE",X"B9",X"FD",X"22",X"04",
		X"8E",X"08",X"6A",X"02",X"F5",X"FE",X"10",X"FE",X"92",X"FE",X"1D",X"FE",X"99",X"FE",X"10",X"FE",
		X"C2",X"FE",X"B4",X"FD",X"E7",X"03",X"97",X"08",X"84",X"02",X"FA",X"FE",X"11",X"FE",X"92",X"FE",
		X"20",X"FE",X"97",X"FE",X"14",X"FE",X"BF",X"FE",X"B8",X"FD",X"69",X"03",X"BD",X"08",X"02",X"03",
		X"28",X"FF",X"0D",X"FE",X"95",X"FE",X"25",X"FE",X"93",X"FE",X"21",X"FE",X"A8",X"FE",X"E6",X"FD",
		X"E4",X"00",X"95",X"08",X"43",X"05",X"04",X"00",X"47",X"FE",X"5A",X"FE",X"68",X"FE",X"4A",X"FE",
		X"7C",X"FE",X"34",X"FE",X"A2",X"FE",X"10",X"FE",X"18",X"05",X"57",X"08",X"46",X"02",X"04",X"FF",
		X"10",X"FE",X"99",X"FE",X"26",X"FE",X"97",X"FE",X"23",X"FE",X"AD",X"FE",X"EB",X"FD",X"B7",X"00",
		X"72",X"08",X"46",X"05",X"FC",X"FF",X"48",X"FE",X"60",X"FE",X"65",X"FE",X"56",X"FE",X"73",X"FE",
		X"4C",X"FE",X"81",X"FE",X"9E",X"FE",X"D0",X"06",X"77",X"07",X"FF",X"00",X"8F",X"FE",X"34",X"FE",
		X"8C",X"FE",X"32",X"FE",X"99",X"FE",X"20",X"FE",X"C4",X"FE",X"C7",X"FD",X"CD",X"03",X"A0",X"08",
		X"E2",X"02",X"23",X"FF",X"19",X"FE",X"96",X"FE",X"36",X"FE",X"8D",X"FE",X"3B",X"FE",X"95",X"FE",
		X"23",X"FE",X"9D",X"FF",X"A0",X"07",X"8A",X"06",X"95",X"00",X"74",X"FE",X"41",X"FE",X"8D",X"FE",
		X"35",X"FE",X"9D",X"FE",X"22",X"FE",X"C7",X"FE",X"D1",X"FD",X"43",X"02",X"ED",X"08",X"3C",X"04",
		X"AA",X"FF",X"37",X"FE",X"79",X"FE",X"5D",X"FE",X"66",X"FE",X"72",X"FE",X"56",X"FE",X"88",X"FE",
		X"7B",X"FE",X"34",X"06",X"A7",X"07",X"58",X"01",X"C2",X"FE",X"2A",X"FE",X"9F",X"FE",X"2F",X"FE",
		X"A6",X"FE",X"21",X"FE",X"CC",X"FE",X"CF",X"FD",X"ED",X"02",X"EE",X"08",X"51",X"03",X"34",X"FF",
		X"23",X"FE",X"9B",X"FE",X"3B",X"FE",X"99",X"FE",X"39",X"FE",X"AE",X"FE",X"FB",X"FD",X"7B",X"00",
		X"56",X"08",X"F4",X"04",X"CC",X"FF",X"46",X"FE",X"7B",X"FE",X"5F",X"FE",X"75",X"FE",X"61",X"FE",
		X"7D",X"FE",X"4B",X"FE",X"7F",X"FF",X"A9",X"07",X"0D",X"06",X"31",X"00",X"60",X"FE",X"66",X"FE",
		X"75",X"FE",X"62",X"FE",X"7C",X"FE",X"60",X"FE",X"79",X"FE",X"F1",X"FE",X"2A",X"07",X"B6",X"06",
		X"6F",X"00",X"76",X"FE",X"57",X"FE",X"85",X"FE",X"56",X"FE",X"8C",X"FE",X"4F",X"FE",X"94",X"FE",
		X"A9",X"FE",X"D7",X"06",X"06",X"07",X"94",X"00",X"81",X"FE",X"52",X"FE",X"8B",X"FE",X"52",X"FE",
		X"91",X"FE",X"4C",X"FE",X"9E",X"FE",X"92",X"FE",X"A8",X"06",X"1C",X"07",X"A2",X"00",X"85",X"FE",
		X"50",X"FE",X"8F",X"FE",X"52",X"FE",X"93",X"FE",X"4D",X"FE",X"9D",X"FE",X"9A",X"FE",X"9D",X"06",
		X"05",X"07",X"9C",X"00",X"87",X"FE",X"56",X"FE",X"8D",X"FE",X"56",X"FE",X"92",X"FE",X"55",X"FE",
		X"95",X"FE",X"B1",X"FE",X"B2",X"06",X"D1",X"06",X"89",X"00",X"82",X"FE",X"5C",X"FE",X"88",X"FE",
		X"5F",X"FE",X"8A",X"FE",X"60",X"FE",X"89",X"FE",X"D3",X"FE",X"DF",X"06",X"88",X"06",X"64",X"00",
		X"7C",X"FE",X"65",X"FE",X"83",X"FE",X"66",X"FE",X"86",X"FE",X"6A",X"FE",X"7C",X"FE",X"F7",X"FE",
		X"25",X"07",X"33",X"06",X"36",X"00",X"70",X"FE",X"71",X"FE",X"7C",X"FE",X"72",X"FE",X"7D",X"FE",
		X"79",X"FE",X"6D",X"FE",X"1E",X"FF",X"7A",X"07",X"DF",X"05",X"FF",X"FF",X"67",X"FE",X"77",X"FE",
		X"7A",X"FE",X"73",X"FE",X"81",X"FE",X"72",X"FE",X"7F",X"FE",X"D7",X"FE",X"DA",X"06",X"9C",X"06",
		X"84",X"00",X"96",X"FE",X"57",X"FE",X"9D",X"FE",X"4F",X"FE",X"AE",X"FE",X"3C",X"FE",X"DA",X"FE",
		X"EE",X"FD",X"0D",X"04",X"6B",X"08",X"6A",X"02",X"13",X"FF",X"3B",X"FE",X"AA",X"FE",X"50",X"FE",
		X"A3",X"FE",X"56",X"FE",X"AA",X"FE",X"3F",X"FE",X"B6",X"FF",X"A2",X"07",X"ED",X"05",X"28",X"00",
		X"89",X"FE",X"60",X"FE",X"9E",X"FE",X"55",X"FE",X"B0",X"FE",X"3F",X"FE",X"D7",X"FE",X"09",X"FE",
		X"E9",X"04",X"31",X"08",X"AE",X"01",X"D1",X"FE",X"41",X"FE",X"B1",X"FE",X"4C",X"FE",X"B6",X"FE",
		X"40",X"FE",X"DB",X"FE",X"E6",X"FD",X"35",X"02",X"77",X"08",X"6A",X"03",X"4A",X"FF",X"49",X"FE",
		X"A2",X"FE",X"61",X"FE",X"9B",X"FE",X"69",X"FE",X"A0",X"FE",X"58",X"FE",X"55",X"FF",X"4B",X"07",
		X"2D",X"06",X"4F",X"00",X"9A",X"FE",X"5B",X"FE",X"AA",X"FE",X"52",X"FE",X"BB",X"FE",X"3E",X"FE",
		X"E7",X"FE",X"DD",X"FD",X"A2",X"02",X"70",X"08",X"82",X"03",X"57",X"FF",X"55",X"FE",X"96",X"FE",
		X"7A",X"FE",X"82",X"FE",X"8F",X"FE",X"70",X"FE",X"AC",X"FE",X"77",X"FE",X"D5",X"05",X"B0",X"07",
		X"32",X"01",X"C4",X"FE",X"49",X"FE",X"BA",X"FE",X"4D",X"FE",X"C0",X"FE",X"44",X"FE",X"DD",X"FE",
		X"FC",X"FD",X"AA",X"01",X"86",X"08",X"F7",X"03",X"5D",X"FF",X"5B",X"FE",X"9B",X"FE",X"77",X"FE",
		X"92",X"FE",X"7D",X"FE",X"94",X"FE",X"70",X"FE",X"44",X"FF",X"29",X"07",X"08",X"06",X"27",X"00",
		X"8D",X"FE",X"71",X"FE",X"A0",X"FE",X"6B",X"FE",X"AC",X"FE",X"5E",X"FE",X"C3",X"FE",X"66",X"FE",
		X"DC",X"05",X"5D",X"07",X"D2",X"00",X"BB",X"FE",X"56",X"FE",X"B9",X"FE",X"55",X"FE",X"C2",X"FE",
		X"45",X"FE",X"EB",X"FE",X"FE",X"FD",X"AC",X"04",X"F2",X"07",X"5D",X"01",X"C9",X"FE",X"50",X"FE",
		X"BE",X"FE",X"52",X"FE",X"C8",X"FE",X"42",X"FE",X"F6",X"FE",X"DA",X"FD",X"CD",X"03",X"26",X"08",
		X"BD",X"01",X"D3",X"FE",X"52",X"FE",X"C1",X"FE",X"55",X"FE",X"CA",X"FE",X"42",X"FE",X"F9",X"FE",
		X"D4",X"FD",X"65",X"03",X"3B",X"08",X"EC",X"01",X"DC",X"FE",X"52",X"FE",X"C2",X"FE",X"54",X"FE",
		X"CC",X"FE",X"43",X"FE",X"FB",X"FE",X"D8",X"FD",X"56",X"03",X"40",X"08",X"F1",X"01",X"DF",X"FE",
		X"55",X"FE",X"C4",X"FE",X"57",X"FE",X"CD",X"FE",X"48",X"FE",X"FA",X"FE",X"E3",X"FD",X"85",X"03",
		X"41",X"08",X"D4",X"01",X"E8",X"FE",X"50",X"FE",X"C9",X"FE",X"55",X"FE",X"D3",X"FE",X"43",X"FE",
		X"FF",X"FE",X"E9",X"FD",X"E7",X"03",X"42",X"08",X"A7",X"01",X"EB",X"FE",X"51",X"FE",X"CB",X"FE",
		X"59",X"FE",X"D1",X"FE",X"48",X"FE",X"FB",X"FE",X"E8",X"FD",X"15",X"03",X"59",X"08",X"5B",X"02",
		X"F7",X"FE",X"59",X"FE",X"BF",X"FE",X"69",X"FE",X"BC",X"FE",X"67",X"FE",X"CD",X"FE",X"3F",X"FE",
		X"61",X"00",X"EE",X"07",X"11",X"05",X"AE",X"FF",X"8D",X"FE",X"82",X"FE",X"AE",X"FE",X"71",X"FE",
		X"C2",X"FE",X"5B",X"FE",X"EC",X"FE",X"14",X"FE",X"5D",X"04",X"2B",X"08",X"D4",X"01",X"F1",X"FE",
		X"5B",X"FE",X"C5",X"FE",X"69",X"FE",X"C3",X"FE",X"68",X"FE",X"D4",X"FE",X"3B",X"FE",X"9A",X"00",
		X"08",X"08",X"A0",X"04",X"87",X"FF",X"84",X"FE",X"96",X"FE",X"9C",X"FE",X"90",X"FE",X"A5",X"FE",
		X"8A",X"FE",X"AD",X"FE",X"C0",X"FE",X"5B",X"06",X"7E",X"06",X"53",X"00",X"AF",X"FE",X"75",X"FE",
		X"BE",X"FE",X"6B",X"FE",X"CF",X"FE",X"57",X"FE",X"FB",X"FE",X"FB",X"FD",X"89",X"03",X"38",X"08",
		X"35",X"02",X"F9",X"FE",X"66",X"FE",X"BF",X"FE",X"79",X"FE",X"B6",X"FE",X"84",X"FE",X"B4",X"FE",
		X"82",X"FE",X"23",X"FF",X"D5",X"06",X"38",X"06",X"4D",X"00",X"B8",X"FE",X"73",X"FE",X"C6",X"FE",
		X"6F",X"FE",X"D2",X"FE",X"61",X"FE",X"F2",X"FE",X"17",X"FE",X"94",X"01",X"27",X"08",X"E0",X"03",
		X"60",X"FF",X"84",X"FE",X"A1",X"FE",X"9F",X"FE",X"93",X"FE",X"B1",X"FE",X"87",X"FE",X"C5",X"FE",
		X"9C",X"FE",X"CB",X"05",X"FD",X"06",X"B4",X"00",X"CB",X"FE",X"70",X"FE",X"CB",X"FE",X"6E",X"FE",
		X"D6",X"FE",X"5D",X"FE",X"FF",X"FE",X"FB",X"FD",X"CB",X"02",X"1C",X"08",X"7C",X"02",X"0E",X"FF",
		X"70",X"FE",X"C2",X"FE",X"81",X"FE",X"BE",X"FE",X"85",X"FE",X"C2",X"FE",X"74",X"FE",X"6E",X"FF",
		X"15",X"07",X"C2",X"05",X"FA",X"FF",X"B6",X"FE",X"7C",X"FE",X"CB",X"FE",X"72",X"FE",X"DC",X"FE",
		X"5F",X"FE",X"04",X"FF",X"08",X"FE",X"39",X"02",X"1E",X"08",X"7A",X"03",X"40",X"FF",X"91",X"FE",
		X"9E",X"FE",X"B5",X"FE",X"86",X"FE",X"CF",X"FE",X"69",X"FE",X"03",X"FF",X"01",X"FE",X"D9",X"03",
		X"E6",X"07",X"38",X"02",X"0D",X"FF",X"82",X"FE",X"B3",X"FE",X"A1",X"FE",X"9E",X"FE",X"BB",X"FE",
		X"82",X"FE",X"EB",X"FE",X"39",X"FE",X"A8",X"04",X"AB",X"07",X"B7",X"01",X"FF",X"FE",X"7B",X"FE",
		X"C2",X"FE",X"93",X"FE",X"AF",X"FE",X"AA",X"FE",X"97",X"FE",X"D3",X"FE",X"66",X"FE",X"1F",X"05",
		X"6A",X"07",X"2E",X"01",X"F1",X"FE",X"6E",X"FE",X"D7",X"FE",X"7A",X"FE",X"D2",X"FE",X"80",X"FE",
		X"D8",X"FE",X"6D",X"FE",X"D1",X"FF",X"2E",X"07",X"81",X"05",X"D4",X"FF",X"BB",X"FE",X"86",X"FE",
		X"D0",X"FE",X"7D",X"FE",X"DD",X"FE",X"6D",X"FE",X"02",X"FF",X"22",X"FE",X"C1",X"03",X"D0",X"07",
		X"D9",X"01",X"FB",X"FE",X"7E",X"FE",X"CB",X"FE",X"8C",X"FE",X"C9",X"FE",X"8F",X"FE",X"CF",X"FE",
		X"7B",X"FE",X"C2",X"FF",X"34",X"07",X"8E",X"05",X"DF",X"FF",X"BF",X"FE",X"85",X"FE",X"D7",X"FE",
		X"7A",X"FE",X"E6",X"FE",X"67",X"FE",X"10",X"FF",X"0C",X"FE",X"B9",X"01",X"0F",X"08",X"88",X"03",
		X"4A",X"FF",X"98",X"FE",X"AC",X"FE",X"B7",X"FE",X"9A",X"FE",X"CE",X"FE",X"83",X"FE",X"F8",X"FE",
		X"3E",X"FE",X"1E",X"04",X"C3",X"07",X"A7",X"01",X"FD",X"FE",X"7D",X"FE",X"D3",X"FE",X"8F",X"FE",
		X"CD",X"FE",X"91",X"FE",X"D6",X"FE",X"77",X"FE",X"FE",X"FF",X"7F",X"07",X"F0",X"04",X"98",X"FF",
		X"B1",X"FE",X"9E",X"FE",X"C5",X"FE",X"96",X"FE",X"D1",X"FE",X"88",X"FE",X"EF",X"FE",X"67",X"FE",
		X"EA",X"04",X"2F",X"07",X"E8",X"00",X"E4",X"FE",X"82",X"FE",X"DE",X"FE",X"83",X"FE",X"E1",X"FE",
		X"7E",X"FE",X"F9",X"FE",X"45",X"FE",X"D7",X"00",X"B4",X"07",X"4A",X"04",X"6D",X"FF",X"B5",X"FE",
		X"9D",X"FE",X"D0",X"FE",X"8D",X"FE",X"E6",X"FE",X"74",X"FE",X"17",X"FF",X"13",X"FE",X"4C",X"03",
		X"FF",X"07",X"2F",X"02",X"03",X"FF",X"8B",X"FE",X"CE",X"FE",X"A1",X"FE",X"C1",X"FE",X"AE",X"FE",
		X"B7",X"FE",X"BD",X"FE",X"E7",X"FE",X"09",X"06",X"57",X"06",X"37",X"00",X"D3",X"FE",X"8A",X"FE",
		X"E1",X"FE",X"86",X"FE",X"EF",X"FE",X"76",X"FE",X"16",X"FF",X"13",X"FE",X"79",X"02",X"E5",X"07",
		X"57",X"02",X"F2",X"FE",X"96",X"FE",X"D1",X"FE",X"9F",X"FE",X"D0",X"FE",X"9E",X"FE",X"DE",X"FE",
		X"7C",X"FE",X"2A",X"00",X"B9",X"07",X"55",X"04",X"61",X"FF",X"B2",X"FE",X"B0",X"FE",X"C2",X"FE",
		X"AC",X"FE",X"C7",X"FE",X"AC",X"FE",X"C8",X"FE",X"FE",X"FE",X"8D",X"06",X"9A",X"05",X"C1",X"FF",
		X"BA",X"FE",X"A6",X"FE",X"CE",X"FE",X"A2",X"FE",X"D7",X"FE",X"9B",X"FE",X"E8",X"FE",X"A7",X"FE",
		X"A0",X"05",X"5B",X"06",X"0B",X"00",X"C5",X"FE",X"9E",X"FE",X"DA",X"FE",X"98",X"FE",X"E5",X"FE",
		X"8E",X"FE",X"FE",X"FE",X"75",X"FE",X"14",X"05",X"BA",X"06",X"4C",X"00",X"D1",X"FE",X"9A",X"FE",
		X"E0",X"FE",X"97",X"FE",X"E9",X"FE",X"8A",X"FE",X"05",X"FF",X"63",X"FE",X"CE",X"04",X"DD",X"06",
		X"65",X"00",X"D1",X"FE",X"9B",X"FE",X"E0",X"FE",X"98",X"FE",X"EB",X"FE",X"8C",X"FE",X"07",X"FF",
		X"62",X"FE",X"BD",X"04",X"DC",X"06",X"60",X"00",X"CE",X"FE",X"9E",X"FE",X"E1",X"FE",X"9A",X"FE",
		X"EA",X"FE",X"8D",X"FE",X"06",X"FF",X"66",X"FE",X"DD",X"04",X"BE",X"06",X"53",X"00",X"D0",X"FE",
		X"A0",X"FE",X"E3",X"FE",X"9B",X"FE",X"EC",X"FE",X"8F",X"FE",X"08",X"FF",X"68",X"FE",X"0C",X"05",
		X"A0",X"06",X"4B",X"00",X"D5",X"FE",X"9E",X"FE",X"E7",X"FE",X"99",X"FE",X"F2",X"FE",X"8A",X"FE",
		X"17",X"FF",X"41",X"FE",X"B7",X"03",X"78",X"07",X"46",X"01",X"F3",X"FE",X"9B",X"FE",X"E6",X"FE",
		X"A1",X"FE",X"E9",X"FE",X"9D",X"FE",X"FA",X"FE",X"6F",X"FE",X"79",X"00",X"63",X"07",X"3F",X"04",
		X"5B",X"FF",X"C8",X"FE",X"B1",X"FE",X"DC",X"FE",X"A8",X"FE",X"EB",X"FE",X"96",X"FE",X"10",X"FF",
		X"56",X"FE",X"1F",X"04",X"4A",X"07",X"15",X"01",X"F3",X"FE",X"9C",X"FE",X"EC",X"FE",X"9F",X"FE",
		X"EF",X"FE",X"97",X"FE",X"0B",X"FF",X"58",X"FE",X"04",X"01",X"97",X"07",X"5B",X"03",X"12",X"FF",
		X"BA",X"FE",X"C8",X"FE",X"C7",X"FE",X"C5",X"FE",X"CC",X"FE",X"C4",X"FE",X"CB",X"FE",X"45",X"FF",
		X"E5",X"06",X"27",X"05",X"83",X"FF",X"DE",X"FE",X"A8",X"FE",X"E8",X"FE",X"A6",X"FE",X"F2",X"FE",
		X"9C",X"FE",X"07",X"FF",X"8A",X"FE",X"B5",X"05",X"1B",X"06",X"F9",X"FF",X"DF",X"FE",X"A7",X"FE",
		X"EE",X"FE",X"A3",X"FE",X"F6",X"FE",X"98",X"FE",X"15",X"FF",X"69",X"FE",X"D8",X"04",X"9F",X"06",
		X"4E",X"00",X"E0",X"FE",X"A5",X"FE",X"F2",X"FE",X"A1",X"FE",X"FB",X"FE",X"90",X"FE",X"21",X"FF",
		X"45",X"FE",X"73",X"03",X"71",X"07",X"46",X"01",X"F7",X"FE",X"A8",X"FE",X"EE",X"FE",X"AB",X"FE",
		X"EE",X"FE",X"A8",X"FE",X"FE",X"FE",X"80",X"FE",X"58",X"00",X"39",X"07",X"41",X"04",X"4D",X"FF",
		X"D9",X"FE",X"B4",X"FE",X"EC",X"FE",X"A8",X"FE",X"FD",X"FE",X"95",X"FE",X"25",X"FF",X"45",X"FE",
		X"7C",X"03",X"83",X"07",X"76",X"01",X"04",X"FF",X"AB",X"FE",X"EA",X"FE",X"B5",X"FE",X"E7",X"FE",
		X"B9",X"FE",X"EE",X"FE",X"A2",X"FE",X"EE",X"FF",X"15",X"07",X"7C",X"04",X"55",X"FF",X"DF",X"FE",
		X"B5",X"FE",X"EB",X"FE",X"B2",X"FE",X"F5",X"FE",X"A5",X"FE",X"10",X"FF",X"8B",X"FE",X"23",X"05",
		X"60",X"06",X"2F",X"00",X"E6",X"FE",X"AD",X"FE",X"F7",X"FE",X"A7",X"FE",X"02",X"FF",X"97",X"FE",
		X"28",X"FF",X"47",X"FE",X"65",X"03",X"60",X"07",X"03",X"01",X"FB",X"FE",X"A8",X"FE",X"FF",X"FE",
		X"A4",X"FE",X"09",X"FF",X"92",X"FE",X"34",X"FF",X"2D",X"FE",X"3F",X"02",X"E3",X"07",X"AB",X"01",
		X"17",X"FF",X"A4",X"FE",X"FF",X"FE",X"A6",X"FE",X"06",X"FF",X"99",X"FE",X"2A",X"FF",X"41",X"FE",
		X"91",X"01",X"C0",X"07",X"2E",X"02",X"13",X"FF",X"B3",X"FE",X"F3",X"FE",X"B6",X"FE",X"FA",X"FE",
		X"A9",X"FE",X"1A",X"FF",X"59",X"FE",X"3F",X"01",X"B7",X"07",X"63",X"02",X"1A",X"FF",X"B4",X"FE",
		X"F6",X"FE",X"B5",X"FE",X"FE",X"FE",X"A9",X"FE",X"1D",X"FF",X"5B",X"FE",X"26",X"01",X"B6",X"07",
		X"7B",X"02",X"16",X"FF",X"BC",X"FE",X"ED",X"FE",X"C1",X"FE",X"EF",X"FE",X"BC",X"FE",X"00",X"FF",
		X"93",X"FE",X"43",X"00",X"22",X"07",X"DC",X"03",X"2D",X"FF",X"DD",X"FE",X"C7",X"FE",X"EE",X"FE",
		X"BF",X"FE",X"FB",X"FE",X"AE",X"FE",X"1F",X"FF",X"6F",X"FE",X"D0",X"04",X"9B",X"06",X"70",X"00",
		X"F8",X"FE",X"B1",X"FE",X"00",X"FF",X"B2",X"FE",X"04",X"FF",X"AF",X"FE",X"16",X"FF",X"7F",X"FE",
		X"8D",X"00",X"31",X"07",X"B5",X"03",X"24",X"FF",X"E2",X"FE",X"C8",X"FE",X"F2",X"FE",X"C2",X"FE",
		X"FF",X"FE",X"B2",X"FE",X"20",X"FF",X"7F",X"FE",X"17",X"05",X"4B",X"06",X"21",X"00",X"FC",X"FE",
		X"B1",X"FE",X"07",X"FF",X"B0",X"FE",X"12",X"FF",X"A1",X"FE",X"37",X"FF",X"4D",X"FE",X"BE",X"02",
		X"6C",X"07",X"50",X"01",X"FB",X"FE",X"BE",X"FE",X"FC",X"FE",X"BB",X"FE",X"07",X"FF",X"AE",X"FE",
		X"28",X"FF",X"5F",X"FE",X"3C",X"01",X"A2",X"07",X"60",X"02",X"19",X"FF",X"C6",X"FE",X"F5",X"FE",
		X"C9",X"FE",X"F9",X"FE",X"C2",X"FE",X"0D",X"FF",X"90",X"FE",X"82",X"00",X"40",X"07",X"2C",X"03",
		X"1C",X"FF",X"DB",X"FE",X"E1",X"FE",X"DE",X"FE",X"E1",X"FE",X"DE",X"FE",X"EB",X"FE",X"CC",X"FE",
		X"B1",X"FF",X"A6",X"06",X"6A",X"04",X"38",X"FF",X"F2",X"FE",X"C5",X"FE",X"FF",X"FE",X"C0",X"FE",
		X"0C",X"FF",X"AE",X"FE",X"31",X"FF",X"68",X"FE",X"2F",X"04",X"BF",X"06",X"AC",X"00",X"F5",X"FE",
		X"C6",X"FE",X"FD",X"FE",X"C8",X"FE",X"FC",X"FE",X"CC",X"FE",X"03",X"FF",X"B3",X"FE",X"F2",X"FF",
		X"C2",X"06",X"60",X"04",X"3E",X"FF",X"F6",X"FE",X"C4",X"FE",X"04",X"FF",X"C0",X"FE",X"11",X"FF",
		X"AF",X"FE",X"34",X"FF",X"67",X"FE",X"86",X"03",X"02",X"07",X"D9",X"00",X"F2",X"FE",X"C8",X"FE",
		X"02",X"FF",X"C6",X"FE",X"0A",X"FF",X"BB",X"FE",X"24",X"FF",X"7C",X"FE",X"EB",X"00",X"50",X"07",
		X"D3",X"02",X"19",X"FF",X"E0",X"FE",X"E8",X"FE",X"E7",X"FE",X"E7",X"FE",X"E9",X"FE",X"E9",X"FE",
		X"E1",X"FE",X"86",X"FF",X"89",X"06",X"66",X"04",X"23",X"FF",X"01",X"FF",X"C7",X"FE",X"06",X"FF",
		X"C6",X"FE",X"0F",X"FF",X"BD",X"FE",X"26",X"FF",X"AF",X"FE",X"EF",X"05",X"63",X"05",X"66",X"FF",
		X"13",X"FF",X"B9",X"FE",X"18",X"FF",X"B9",X"FE",X"1F",X"FF",X"AD",X"FE",X"41",X"FF",X"72",X"FE",
		X"60",X"05",X"D8",X"05",X"A7",X"FF",X"13",X"FF",X"B9",X"FE",X"19",X"FF",X"BB",X"FE",X"21",X"FF",
		X"AB",X"FE",X"46",X"FF",X"65",X"FE",X"FF",X"04",X"0E",X"06",X"C4",X"FF",X"16",X"FF",X"B9",X"FE",
		X"1C",X"FF",X"B8",X"FE",X"26",X"FF",X"A7",X"FE",X"4D",X"FF",X"5B",X"FE",X"E5",X"04",X"22",X"06",
		X"C4",X"FF",X"1A",X"FF",X"B7",X"FE",X"20",X"FF",X"B7",X"FE",X"2B",X"FF",X"A5",X"FE",X"53",X"FF",
		X"4D",X"FE",X"FE",X"04",X"23",X"06",X"A7",X"FF",X"1F",X"FF",X"B6",X"FE",X"23",X"FF",X"B8",X"FE",
		X"2C",X"FF",X"A7",X"FE",X"50",X"FF",X"62",X"FE",X"02",X"05",X"F2",X"05",X"88",X"FF",X"16",X"FF",
		X"BD",X"FE",X"1E",X"FF",X"BF",X"FE",X"25",X"FF",X"B2",X"FE",X"44",X"FF",X"7E",X"FE",X"FA",X"04",
		X"F5",X"05",X"9E",X"FF",X"13",X"FF",X"C1",X"FE",X"1E",X"FF",X"BF",X"FE",X"29",X"FF",X"AF",X"FE",
		X"51",X"FF",X"54",X"FE",X"38",X"03",X"E6",X"06",X"F9",X"00",X"07",X"FF",X"D6",X"FE",X"08",X"FF",
		X"DB",X"FE",X"08",X"FF",X"DD",X"FE",X"0E",X"FF",X"C8",X"FE",X"D2",X"FF",X"9F",X"06",X"2D",X"04",
		X"4F",X"FF",X"06",X"FF",X"D2",X"FE",X"14",X"FF",X"CC",X"FE",X"20",X"FF",X"BB",X"FE",X"48",X"FF",
		X"62",X"FE",X"60",X"03",X"D2",X"06",X"CF",X"00",X"12",X"FF",X"CF",X"FE",X"15",X"FF",X"D0",X"FE",
		X"19",X"FF",X"CC",X"FE",X"2F",X"FF",X"93",X"FE",X"8F",X"00",X"6B",X"07",X"BB",X"02",X"0D",X"FF",
		X"F8",X"FE",X"ED",X"FE",X"FD",X"FE",X"EC",X"FE",X"02",X"FF",X"E8",X"FE",X"07",X"FF",X"37",X"FF",
		X"E3",X"05",X"E7",X"04",X"63",X"FF",X"14",X"FF",X"CF",X"FE",X"1F",X"FF",X"CA",X"FE",X"29",X"FF",
		X"BB",X"FE",X"4C",X"FF",X"6C",X"FE",X"7C",X"02",X"09",X"07",X"8D",X"01",X"F0",X"FE",X"F8",X"FE",
		X"F0",X"FE",X"00",X"FF",X"E7",X"FE",X"11",X"FF",X"D3",X"FE",X"38",X"FF",X"9A",X"FE",X"32",X"05",
		X"0A",X"06",X"D6",X"FF",X"2C",X"FF",X"BF",X"FE",X"2F",X"FF",X"C4",X"FE",X"2F",X"FF",X"BE",X"FE",
		X"45",X"FF",X"88",X"FE",X"BC",X"00",X"18",X"07",X"EB",X"02",X"0F",X"FF",X"0E",X"FF",X"DE",X"FE",
		X"16",X"FF",X"D8",X"FE",X"25",X"FF",X"C6",X"FE",X"48",X"FF",X"8D",X"FE",X"63",X"05",X"9A",X"05",
		X"81",X"FF",X"27",X"FF",X"C8",X"FE",X"2B",X"FF",X"C8",X"FE",X"32",X"FF",X"BD",X"FE",X"55",X"FF",
		X"6F",X"FE",X"3F",X"03",X"9C",X"06",X"9E",X"00",X"0F",X"FF",X"DC",X"FE",X"1D",X"FF",X"D9",X"FE",
		X"24",X"FF",X"CC",X"FE",X"45",X"FF",X"7E",X"FE",X"BB",X"01",X"25",X"07",X"67",X"01",X"02",X"FF",
		X"E9",X"FE",X"12",X"FF",X"E4",X"FE",X"1B",X"FF",X"D7",X"FE",X"39",X"FF",X"95",X"FE",X"E2",X"00",
		X"5C",X"07",X"F5",X"01",X"FB",X"FE",X"F5",X"FE",X"08",X"FF",X"EE",X"FE",X"11",X"FF",X"E6",X"FE",
		X"2A",X"FF",X"B0",X"FE",X"8D",X"00",X"4E",X"07",X"52",X"02",X"FE",X"FE",X"FD",X"FE",X"03",X"FF",
		X"F6",X"FE",X"0C",X"FF",X"ED",X"FE",X"21",X"FF",X"BB",X"FE",X"5D",X"00",X"40",X"07",X"76",X"02",
		X"FA",X"FE",X"02",X"FF",X"FF",X"FE",X"FC",X"FE",X"0A",X"FF",X"F2",X"FE",X"1F",X"FF",X"C2",X"FE",
		X"4A",X"00",X"38",X"07",X"70",X"02",X"F5",X"FE",X"07",X"FF",X"03",X"FF",X"FB",X"FE",X"0C",X"FF",
		X"F2",X"FE",X"22",X"FF",X"C3",X"FE",X"4F",X"00",X"17",X"07",X"56",X"02",X"FA",X"FE",X"05",X"FF",
		X"04",X"FF",X"FA",X"FE",X"0F",X"FF",X"F3",X"FE",X"22",X"FF",X"C3",X"FE",X"7C",X"00",X"FF",X"06",
		X"58",X"02",X"FD",X"FE",X"07",X"FF",X"00",X"FF",X"03",X"FF",X"06",X"FF",X"03",X"FF",X"0B",X"FF",
		X"F7",X"FE",X"92",X"FF",X"62",X"06",X"F4",X"03",X"2C",X"FF",X"29",X"FF",X"DB",X"FE",X"2F",X"FF",
		X"D6",X"FE",X"3C",X"FF",X"C2",X"FE",X"69",X"FF",X"5C",X"FE",X"63",X"03",X"AD",X"06",X"99",X"00",
		X"25",X"FF",X"E4",X"FE",X"23",X"FF",X"E9",X"FE",X"20",X"FF",X"EE",X"FE",X"25",X"FF",X"DF",X"FE",
		X"C6",X"FF",X"72",X"06",X"CA",X"03",X"20",X"FF",X"31",X"FF",X"D8",X"FE",X"36",X"FF",X"D3",X"FE",
		X"44",X"FF",X"BF",X"FE",X"72",X"FF",X"58",X"FE",X"3A",X"04",X"24",X"06",X"BB",X"FF",X"2D",X"FF",
		X"D8",X"FE",X"35",X"FF",X"DA",X"FE",X"3B",X"FF",X"CF",X"FE",X"5A",X"FF",X"84",X"FE",X"17",X"02",
		X"C3",X"06",X"57",X"01",X"0D",X"FF",X"01",X"FF",X"0F",X"FF",X"04",X"FF",X"0D",X"FF",X"08",X"FF",
		X"0C",X"FF",X"0A",X"FF",X"66",X"FF",X"D7",X"05",X"78",X"04",X"55",X"FF",X"2F",X"FF",X"DE",X"FE",
		X"34",X"FF",X"DE",X"FE",X"3B",X"FF",X"D4",X"FE",X"56",X"FF",X"96",X"FE",X"4D",X"01",X"F5",X"06",
		X"26",X"02",X"F0",X"FE",X"23",X"FF",X"F0",X"FE",X"28",X"FF",X"E9",X"FE",X"3B",X"FF",X"D2",X"FE",
		X"67",X"FF",X"74",X"FE",X"7B",X"04",X"0B",X"06",X"C7",X"FF",X"3B",X"FF",X"D9",X"FE",X"3B",X"FF",
		X"DE",X"FE",X"3E",X"FF",X"D8",X"FE",X"56",X"FF",X"9A",X"FE",X"06",X"01",X"00",X"07",X"E6",X"01",
		X"FA",X"FE",X"16",X"FF",X"07",X"FF",X"14",X"FF",X"0A",X"FF",X"15",X"FF",X"0B",X"FF",X"0B",X"FF",
		X"95",X"FF",X"19",X"06",X"B9",X"03",X"1F",X"FF",X"30",X"FF",X"EA",X"FE",X"31",X"FF",X"EB",X"FE",
		X"3A",X"FF",X"DF",X"FE",X"55",X"FF",X"C0",X"FE",X"10",X"05",X"00",X"05",X"4A",X"FF",X"43",X"FF",
		X"D9",X"FE",X"46",X"FF",X"D9",X"FE",X"4F",X"FF",X"C8",X"FE",X"79",X"FF",X"69",X"FE",X"73",X"04",
		X"B7",X"05",X"7B",X"FF",X"46",X"FF",X"D5",X"FE",X"49",X"FF",X"D7",X"FE",X"53",X"FF",X"C5",X"FE",
		X"7F",X"FF",X"5F",X"FE",X"16",X"04",X"0C",X"06",X"A1",X"FF",X"41",X"FF",X"D9",X"FE",X"48",X"FF",
		X"D8",X"FE",X"54",X"FF",X"C8",X"FE",X"7E",X"FF",X"5F",X"FE",X"D6",X"03",X"29",X"06",X"B4",X"FF",
		X"42",X"FF",X"DA",X"FE",X"4B",X"FF",X"DA",X"FE",X"55",X"FF",X"C6",X"FE",X"82",X"FF",X"5C",X"FE",
		X"BE",X"03",X"27",X"06",X"B9",X"FF",X"43",X"FF",X"DA",X"FE",X"4B",X"FF",X"DC",X"FE",X"56",X"FF",
		X"C8",X"FE",X"82",X"FF",X"5D",X"FE",X"B1",X"03",X"03",X"06",X"B0",X"FF",X"48",X"FF",X"DA",X"FE",
		X"4C",X"FF",X"DC",X"FE",X"56",X"FF",X"CA",X"FE",X"80",X"FF",X"69",X"FE",X"BF",X"03",X"DB",X"05",
		X"B1",X"FF",X"44",X"FF",X"E0",X"FE",X"4A",X"FF",X"E1",X"FE",X"53",X"FF",X"D1",X"FE",X"7A",X"FF",
		X"6D",X"FE",X"BB",X"02",X"9A",X"06",X"82",X"00",X"23",X"FF",X"00",X"FF",X"2C",X"FF",X"02",X"FF",
		X"2D",X"FF",X"07",X"FF",X"2E",X"FF",X"F8",X"FE",X"B3",X"FF",X"87",X"06",X"7B",X"03",X"F9",X"FE",
		X"4C",X"FF",X"E5",X"FE",X"4A",X"FF",X"E1",X"FE",X"58",X"FF",X"CF",X"FE",X"84",X"FF",X"66",X"FE",
		X"2C",X"03",X"7A",X"06",X"44",X"00",X"29",X"FF",X"FD",X"FE",X"34",X"FF",X"00",X"FF",X"33",X"FF",
		X"FF",X"FE",X"3F",X"FF",X"DE",X"FE",X"37",X"00",X"96",X"06",X"80",X"02",X"FC",X"FE",X"35",X"FF",
		X"01",X"FF",X"32",X"FF",X"05",X"FF",X"33",X"FF",X"01",X"FF",X"3B",X"FF",X"36",X"FF",X"A9",X"05",
		X"09",X"04",X"1E",X"FF",X"4A",X"FF",X"EF",X"FE",X"44",X"FF",X"F1",X"FE",X"4B",X"FF",X"E6",X"FE",
		X"67",X"FF",X"BC",X"FE",X"82",X"04",X"12",X"05",X"66",X"FF",X"50",X"FF",X"E5",X"FE",X"51",X"FF",
		X"E6",X"FE",X"5A",X"FF",X"D6",X"FE",X"81",X"FF",X"80",X"FE",X"C6",X"03",X"A4",X"05",X"A1",X"FF",
		X"4E",X"FF",X"E7",X"FE",X"53",X"FF",X"E8",X"FE",X"5A",X"FF",X"D6",X"FE",X"83",X"FF",X"75",X"FE",
		X"B0",X"02",X"87",X"06",X"65",X"00",X"25",X"FF",X"07",X"FF",X"33",X"FF",X"0B",X"FF",X"30",X"FF",
		X"0F",X"FF",X"33",X"FF",X"05",X"FF",X"AB",X"FF",X"61",X"06",X"66",X"03",X"F7",X"FE",X"54",X"FF",
		X"EC",X"FE",X"51",X"FF",X"EC",X"FE",X"5A",X"FF",X"DC",X"FE",X"81",X"FF",X"7F",X"FE",X"8F",X"02",
		X"6F",X"06",X"B4",X"00",X"22",X"FF",X"15",X"FF",X"29",X"FF",X"19",X"FF",X"27",X"FF",X"1E",X"FF",
		X"25",X"FF",X"1A",X"FF",X"8C",X"FF",X"18",X"06",X"82",X"03",X"F9",X"FE",X"55",X"FF",X"F0",X"FE",
		X"51",X"FF",X"F1",X"FE",X"5B",X"FF",X"DF",X"FE",X"83",X"FF",X"8C",X"FE",X"F9",X"03",X"7A",X"05",
		X"91",X"FF",X"56",X"FF",X"EC",X"FE",X"59",X"FF",X"ED",X"FE",X"60",X"FF",X"DE",X"FE",X"85",X"FF",
		X"81",X"FE",X"B6",X"02",X"4C",X"06",X"38",X"00",X"32",X"FF",X"06",X"FF",X"43",X"FF",X"03",X"FF",
		X"4A",X"FF",X"F8",X"FE",X"67",X"FF",X"B1",X"FE",X"A0",X"01",X"62",X"06",X"EB",X"00",X"1C",X"FF",
		X"1A",X"FF",X"31",X"FF",X"14",X"FF",X"3C",X"FF",X"0A",X"FF",X"53",X"FF",X"D2",X"FE",X"02",X"01",
		X"62",X"06",X"5B",X"01",X"14",X"FF",X"27",X"FF",X"29",X"FF",X"1C",X"FF",X"36",X"FF",X"15",X"FF",
		X"49",X"FF",X"E3",X"FE",X"BB",X"00",X"5A",X"06",X"8E",X"01",X"10",X"FF",X"2D",X"FF",X"28",X"FF",
		X"21",X"FF",X"31",X"FF",X"18",X"FF",X"46",X"FF",X"E6",X"FE",X"AE",X"00",X"55",X"06",X"92",X"01",
		X"0C",X"FF",X"31",X"FF",X"27",X"FF",X"24",X"FF",X"32",X"FF",X"19",X"FF",X"4A",X"FF",X"E6",X"FE",
		X"C7",X"00",X"5B",X"06",X"6E",X"01",X"0C",X"FF",X"2C",X"FF",X"2D",X"FF",X"1F",X"FF",X"39",X"FF",
		X"13",X"FF",X"54",X"FF",X"D6",X"FE",X"FF",X"00",X"6A",X"06",X"39",X"01",X"0D",X"FF",X"29",X"FF",
		X"31",X"FF",X"1E",X"FF",X"3D",X"FF",X"11",X"FF",X"56",X"FF",X"D8",X"FE",X"E8",X"00",X"6A",X"06",
		X"78",X"01",X"03",X"FF",X"3A",X"FF",X"20",X"FF",X"33",X"FF",X"21",X"FF",X"37",X"FF",X"1E",X"FF",
		X"40",X"FF",X"36",X"FF",X"A9",X"05",X"AB",X"03",X"05",X"FF",X"6B",X"FF",X"EF",X"FE",X"67",X"FF",
		X"F0",X"FE",X"6F",X"FF",X"DE",X"FE",X"98",X"FF",X"7D",X"FE",X"57",X"02",X"53",X"06",X"87",X"00",
		X"30",X"FF",X"21",X"FF",X"35",X"FF",X"28",X"FF",X"2F",X"FF",X"32",X"FF",X"29",X"FF",X"3B",X"FF",
		X"51",X"FF",X"C5",X"05",X"75",X"03",X"02",X"FF",X"6A",X"FF",X"F8",X"FE",X"60",X"FF",X"FC",X"FE",
		X"67",X"FF",X"F0",X"FE",X"87",X"FF",X"AE",X"FE",X"CA",X"03",X"3D",X"05",X"8F",X"FF",X"5D",X"FF",
		X"FF",X"FE",X"5E",X"FF",X"00",X"FF",X"66",X"FF",X"F2",X"FE",X"86",X"FF",X"A0",X"FE",X"C8",X"01",
		X"73",X"06",X"E7",X"00",X"1D",X"FF",X"32",X"FF",X"2C",X"FF",X"36",X"FF",X"27",X"FF",X"41",X"FF",
		X"1A",X"FF",X"59",X"FF",X"10",X"FF",X"25",X"05",X"62",X"04",X"2D",X"FF",X"67",X"FF",X"FE",X"FE",
		X"5E",X"FF",X"07",X"FF",X"5C",X"FF",X"07",X"FF",X"68",X"FF",X"E6",X"FE",X"84",X"00",X"1A",X"06",
		X"4E",X"02",X"01",X"FF",X"62",X"FF",X"06",X"FF",X"61",X"FF",X"00",X"FF",X"6C",X"FF",X"EE",X"FE",
		X"97",X"FF",X"95",X"FE",X"71",X"03",X"7E",X"05",X"BE",X"FF",X"59",X"FF",X"09",X"FF",X"59",X"FF",
		X"10",X"FF",X"59",X"FF",X"0E",X"FF",X"6A",X"FF",X"DB",X"FE",X"F3",X"00",X"28",X"06",X"76",X"01",
		X"0E",X"FF",X"49",X"FF",X"24",X"FF",X"44",X"FF",X"23",X"FF",X"4A",X"FF",X"1C",X"FF",X"5B",X"FF",
		X"23",X"FF",X"17",X"05",X"21",X"04",X"1C",X"FF",X"72",X"FF",X"FC",X"FE",X"6B",X"FF",X"02",X"FF",
		X"6E",X"FF",X"FC",X"FE",X"83",X"FF",X"C5",X"FE",X"1F",X"01",X"1A",X"06",X"B9",X"01",X"02",X"FF",
		X"65",X"FF",X"08",X"FF",X"67",X"FF",X"01",X"FF",X"78",X"FF",X"EA",X"FE",X"A5",X"FF",X"86",X"FE",
		X"EE",X"02",X"FE",X"05",X"58",X"00",X"25",X"FF",X"41",X"FF",X"27",X"FF",X"51",X"FF",X"15",X"FF",
		X"68",X"FF",X"F7",X"FE",X"9C",X"FF",X"8B",X"FE",X"BE",X"03",X"AD",X"05",X"E0",X"FF",X"48",X"FF",
		X"26",X"FF",X"3F",X"FF",X"3C",X"FF",X"2C",X"FF",X"56",X"FF",X"0C",X"FF",X"88",X"FF",X"A8",X"FE",
		X"0A",X"04",X"81",X"05",X"A0",X"FF",X"64",X"FF",X"11",X"FF",X"59",X"FF",X"22",X"FF",X"4A",X"FF",
		X"34",X"FF",X"3B",X"FF",X"49",X"FF",X"45",X"FF",X"07",X"05",X"F2",X"03",X"16",X"FF",X"83",X"FF",
		X"F7",X"FE",X"7A",X"FF",X"FF",X"FE",X"7B",X"FF",X"F4",X"FE",X"96",X"FF",X"AD",X"FE",X"98",X"01",
		X"0C",X"06",X"CA",X"00",X"29",X"FF",X"41",X"FF",X"35",X"FF",X"45",X"FF",X"2F",X"FF",X"4F",X"FF",
		X"22",X"FF",X"66",X"FF",X"18",X"FF",X"01",X"05",X"F2",X"03",X"1C",X"FF",X"81",X"FF",X"FE",X"FE",
		X"76",X"FF",X"07",X"FF",X"78",X"FF",X"FF",X"FE",X"8B",X"FF",X"C9",X"FE",X"F5",X"00",X"4C",X"06",
		X"BC",X"01",X"03",X"FF",X"66",X"FF",X"15",X"FF",X"68",X"FF",X"10",X"FF",X"75",X"FF",X"FC",X"FE",
		X"9C",X"FF",X"A5",X"FE",X"51",X"02",X"DD",X"05",X"68",X"00",X"3F",X"FF",X"38",X"FF",X"3F",X"FF",
		X"43",X"FF",X"36",X"FF",X"50",X"FF",X"27",X"FF",X"68",X"FF",X"16",X"FF",X"31",X"05",X"C5",X"03",
		X"10",X"FF",X"84",X"FF",X"00",X"FF",X"7A",X"FF",X"07",X"FF",X"7F",X"FF",X"F9",X"FE",X"A2",X"FF",
		X"A2",X"FE",X"77",X"02",X"A5",X"05",X"F6",X"FF",X"5C",X"FF",X"1C",X"FF",X"62",X"FF",X"1E",X"FF",
		X"66",X"FF",X"18",X"FF",X"7B",X"FF",X"E0",X"FE",X"F9",X"00",X"20",X"06",X"34",X"01",X"1E",X"FF",
		X"4E",X"FF",X"38",X"FF",X"49",X"FF",X"3D",X"FF",X"49",X"FF",X"41",X"FF",X"3C",X"FF",X"D5",X"FF",
		X"AE",X"05",X"35",X"02",X"EF",X"FE",X"73",X"FF",X"1B",X"FF",X"65",X"FF",X"24",X"FF",X"69",X"FF",
		X"1D",X"FF",X"7C",X"FF",X"07",X"FF",X"14",X"05",X"A0",X"03",X"09",X"FF",X"8C",X"FF",X"02",X"FF",
		X"7F",X"FF",X"07",X"FF",X"86",X"FF",X"F8",X"FE",X"AA",X"FF",X"A0",X"FE",X"49",X"02",X"B1",X"05",
		X"3A",X"00",X"48",X"FF",X"3B",X"FF",X"47",X"FF",X"44",X"FF",X"3E",X"FF",X"54",X"FF",X"2F",X"FF",
		X"6C",X"FF",X"18",X"FF",X"1F",X"05",X"E6",X"03",X"13",X"FF",X"8F",X"FF",X"02",X"FF",X"84",X"FF",
		X"08",X"FF",X"88",X"FF",X"FC",X"FE",X"A9",X"FF",X"AA",X"FE",X"C7",X"01",X"1E",X"06",X"A1",X"00",
		X"3C",X"FF",X"45",X"FF",X"46",X"FF",X"48",X"FF",X"42",X"FF",X"50",X"FF",X"3B",X"FF",X"57",X"FF",
		X"64",X"FF",X"6A",X"05",X"BB",X"02",X"F7",X"FE",X"86",X"FF",X"11",X"FF",X"79",X"FF",X"17",X"FF",
		X"7C",X"FF",X"0D",X"FF",X"97",X"FF",X"E0",X"FE",X"99",X"04",X"1C",X"04",X"24",X"FF",X"88",X"FF",
		X"0F",X"FF",X"7E",X"FF",X"12",X"FF",X"84",X"FF",X"07",X"FF",X"A4",X"FF",X"B9",X"FE",X"59",X"03",
		X"D9",X"04",X"5A",X"FF",X"7E",X"FF",X"14",X"FF",X"7B",X"FF",X"17",X"FF",X"81",X"FF",X"08",X"FF",
		X"A7",X"FF",X"B0",X"FE",X"94",X"02",X"42",X"05",X"89",X"FF",X"74",X"FF",X"1A",X"FF",X"7A",X"FF",
		X"1B",X"FF",X"82",X"FF",X"0B",X"FF",X"A5",X"FF",X"B2",X"FE",X"2F",X"02",X"6E",X"05",X"B2",X"FF",
		X"6F",X"FF",X"20",X"FF",X"77",X"FF",X"1E",X"FF",X"7F",X"FF",X"0F",X"FF",X"A2",X"FF",X"BA",X"FE",
		X"12",X"02",X"73",X"05",X"BA",X"FF",X"6B",X"FF",X"23",X"FF",X"74",X"FF",X"23",X"FF",X"7D",X"FF",
		X"15",X"FF",X"A1",X"FF",X"C1",X"FE",X"28",X"02",X"62",X"05",X"BA",X"FF",X"6E",X"FF",X"24",X"FF",
		X"77",X"FF",X"1F",X"FF",X"80",X"FF",X"13",X"FF",X"A4",X"FF",X"BF",X"FE",X"68",X"02",X"42",X"05",
		X"B0",X"FF",X"72",X"FF",X"22",X"FF",X"79",X"FF",X"22",X"FF",X"81",X"FF",X"14",X"FF",X"A4",X"FF",
		X"C2",X"FE",X"88",X"02",X"44",X"05",X"B8",X"FF",X"74",X"FF",X"24",X"FF",X"79",X"FF",X"26",X"FF",
		X"7C",X"FF",X"1D",X"FF",X"95",X"FF",X"E2",X"FE",X"FA",X"00",X"D6",X"05",X"E8",X"00",X"2E",X"FF",
		X"64",X"FF",X"3E",X"FF",X"66",X"FF",X"38",X"FF",X"72",X"FF",X"25",X"FF",X"95",X"FF",X"E4",X"FE",
		X"6F",X"04",X"FC",X"03",X"1B",X"FF",X"9E",X"FF",X"0D",X"FF",X"8E",X"FF",X"16",X"FF",X"8E",X"FF",
		X"11",X"FF",X"A5",X"FF",X"D3",X"FE",X"2E",X"01",X"C8",X"05",X"C8",X"00",X"35",X"FF",X"61",X"FF",
		X"43",X"FF",X"62",X"FF",X"41",X"FF",X"69",X"FF",X"3A",X"FF",X"73",X"FF",X"5D",X"FF",X"0F",X"05",
		X"CB",X"02",X"EE",X"FE",X"99",X"FF",X"19",X"FF",X"87",X"FF",X"1F",X"FF",X"8C",X"FF",X"0F",X"FF",
		X"B0",X"FF",X"BD",X"FE",X"EE",X"03",X"A5",X"04",X"4C",X"FF",X"98",X"FF",X"14",X"FF",X"8C",X"FF",
		X"20",X"FF",X"8A",X"FF",X"1D",X"FF",X"9B",X"FF",X"EE",X"FE",X"CD",X"00",X"F6",X"05",X"6D",X"01",
		X"1C",X"FF",X"7C",X"FF",X"2D",X"FF",X"7C",X"FF",X"28",X"FF",X"8A",X"FF",X"16",X"FF",X"B0",X"FF",
		X"C5",X"FE",X"D5",X"02",X"1D",X"05",X"C1",X"FF",X"63",X"FF",X"44",X"FF",X"61",X"FF",X"4F",X"FF",
		X"57",X"FF",X"5C",X"FF",X"4A",X"FF",X"6D",X"FF",X"56",X"FF",X"FC",X"04",X"E2",X"02",X"EE",X"FE",
		X"A6",X"FF",X"12",X"FF",X"94",X"FF",X"1A",X"FF",X"99",X"FF",X"0E",X"FF",X"BB",X"FF",X"BE",X"FE",
		X"CC",X"02",X"EE",X"04",X"93",X"FF",X"7A",X"FF",X"33",X"FF",X"77",X"FF",X"38",X"FF",X"79",X"FF",
		X"35",X"FF",X"89",X"FF",X"09",X"FF",X"B0",X"00",X"B9",X"05",X"53",X"01",X"25",X"FF",X"77",X"FF",
		X"3C",X"FF",X"75",X"FF",X"38",X"FF",X"82",X"FF",X"25",X"FF",X"A9",X"FF",X"D9",X"FE",X"69",X"03",
		X"AE",X"04",X"74",X"FF",X"82",X"FF",X"35",X"FF",X"75",X"FF",X"45",X"FF",X"68",X"FF",X"54",X"FF",
		X"57",X"FF",X"6E",X"FF",X"4E",X"FF",X"F8",X"04",X"59",X"03",X"0D",X"FF",X"A6",X"FF",X"1B",X"FF",
		X"8F",X"FF",X"2D",X"FF",X"85",X"FF",X"37",X"FF",X"7E",X"FF",X"37",X"FF",X"C7",X"FF",X"3E",X"05",
		X"85",X"02",X"FE",X"FE",X"A7",X"FF",X"1A",X"FF",X"94",X"FF",X"27",X"FF",X"8D",X"FF",X"30",X"FF",
		X"8C",X"FF",X"24",X"FF",X"FD",X"FF",X"61",X"05",X"46",X"02",X"02",X"FF",X"A4",X"FF",X"1E",X"FF",
		X"93",X"FF",X"2A",X"FF",X"8E",X"FF",X"2D",X"FF",X"90",X"FF",X"20",X"FF",X"13",X"00",X"80",X"05",
		X"4A",X"02",X"08",X"FF",X"A2",X"FF",X"20",X"FF",X"94",X"FF",X"2A",X"FF",X"91",X"FF",X"2E",X"FF",
		X"93",X"FF",X"1E",X"FF",X"27",X"00",X"A6",X"05",X"4F",X"02",X"09",X"FF",X"A2",X"FF",X"1F",X"FF",
		X"95",X"FF",X"28",X"FF",X"95",X"FF",X"29",X"FF",X"9C",X"FF",X"10",X"FF",X"56",X"00",X"A0",X"05",
		X"05",X"02",X"06",X"FF",X"A5",X"FF",X"1D",X"FF",X"9E",X"FF",X"1D",X"FF",X"A4",X"FF",X"12",X"FF",
		X"C4",X"FF",X"CA",X"FE",X"C5",X"01",X"3E",X"05",X"38",X"00",X"43",X"FF",X"70",X"FF",X"4D",X"FF",
		X"74",X"FF",X"49",X"FF",X"7D",X"FF",X"3E",X"FF",X"90",X"FF",X"3F",X"FF",X"BB",X"04",X"CB",X"02",
		X"FA",X"FE",X"A5",X"FF",X"26",X"FF",X"94",X"FF",X"2D",X"FF",X"9A",X"FF",X"1F",X"FF",X"BF",X"FF",
		X"C9",X"FE",X"41",X"03",X"9B",X"04",X"5D",X"FF",X"A2",X"FF",X"26",X"FF",X"98",X"FF",X"2D",X"FF",
		X"99",X"FF",X"24",X"FF",X"B4",X"FF",X"DD",X"FE",X"6F",X"01",X"37",X"05",X"08",X"00",X"67",X"FF",
		X"52",X"FF",X"75",X"FF",X"4E",X"FF",X"7B",X"FF",X"46",X"FF",X"90",X"FF",X"15",X"FF",X"BF",X"00",
		X"84",X"05",X"8E",X"00",X"48",X"FF",X"67",X"FF",X"64",X"FF",X"5E",X"FF",X"6D",X"FF",X"59",X"FF",
		X"7B",X"FF",X"35",X"FF",X"5C",X"00",X"9B",X"05",X"F8",X"00",X"3C",X"FF",X"6F",X"FF",X"5E",X"FF",
		X"64",X"FF",X"67",X"FF",X"5E",X"FF",X"71",X"FF",X"49",X"FF",X"11",X"00",X"95",X"05",X"8B",X"01",
		X"20",X"FF",X"91",X"FF",X"3F",X"FF",X"8A",X"FF",X"3D",X"FF",X"92",X"FF",X"2D",X"FF",X"B6",X"FF",
		X"E3",X"FE",X"03",X"04",X"90",X"03",X"F8",X"FE",X"BA",X"FF",X"1E",X"FF",X"A3",X"FF",X"2B",X"FF",
		X"A0",X"FF",X"29",X"FF",X"B2",X"FF",X"F7",X"FE",X"E1",X"00",X"64",X"05",X"DD",X"00",X"2A",X"FF",
		X"91",X"FF",X"3D",X"FF",X"92",X"FF",X"37",X"FF",X"A1",X"FF",X"20",X"FF",X"CA",X"FF",X"C9",X"FE",
		X"E9",X"02",X"BC",X"04",X"C1",X"FF",X"71",X"FF",X"60",X"FF",X"63",X"FF",X"74",X"FF",X"50",X"FF",
		X"8C",X"FF",X"34",X"FF",X"BC",X"FF",X"DE",X"FE",X"09",X"04",X"34",X"04",X"57",X"FF",X"98",X"FF",
		X"44",X"FF",X"7D",X"FF",X"61",X"FF",X"64",X"FF",X"7A",X"FF",X"49",X"FF",X"A6",X"FF",X"02",X"FF",
		X"50",X"04",X"EE",X"03",X"3D",X"FF",X"A3",X"FF",X"3C",X"FF",X"86",X"FF",X"56",X"FF",X"70",X"FF",
		X"70",X"FF",X"54",X"FF",X"97",X"FF",X"18",X"FF",X"1A",X"04",X"E6",X"03",X"3E",X"FF",X"A6",X"FF",
		X"39",X"FF",X"8C",X"FF",X"52",X"FF",X"77",X"FF",X"69",X"FF",X"5E",X"FF",X"8F",X"FF",X"28",X"FF",
		X"EE",X"03",X"D9",X"03",X"29",X"FF",X"B5",X"FF",X"2A",X"FF",X"9E",X"FF",X"3F",X"FF",X"8F",X"FF",
		X"4D",X"FF",X"84",X"FF",X"55",X"FF",X"B3",X"FF",X"FF",X"04",X"60",X"02",X"F3",X"FE",X"C7",X"FF",
		X"19",X"FF",X"B7",X"FF",X"20",X"FF",X"BA",X"FF",X"12",X"FF",X"DE",X"FF",X"BA",X"FE",X"6C",X"02",
		X"FB",X"04",X"B8",X"FF",X"86",X"FF",X"52",X"FF",X"7E",X"FF",X"5D",X"FF",X"7B",X"FF",X"5F",X"FF",
		X"7C",X"FF",X"52",X"FF",X"F9",X"FF",X"20",X"05",X"54",X"01",X"19",X"FF",X"9C",X"FF",X"46",X"FF",
		X"8E",X"FF",X"4C",X"FF",X"92",X"FF",X"45",X"FF",X"A2",X"FF",X"40",X"FF",X"AB",X"04",X"AE",X"02",
		X"05",X"FF",X"B8",X"FF",X"2D",X"FF",X"A7",X"FF",X"34",X"FF",X"AE",X"FF",X"25",X"FF",X"D3",X"FF",
		X"C4",X"FE",X"16",X"03",X"07",X"04",X"2D",X"FF",X"B6",X"FF",X"30",X"FF",X"A4",X"FF",X"3D",X"FF",
		X"A0",X"FF",X"3D",X"FF",X"AD",X"FF",X"17",X"FF",X"A6",X"00",X"0F",X"05",X"F4",X"00",X"29",X"FF",
		X"A0",X"FF",X"41",X"FF",X"A0",X"FF",X"3A",X"FF",X"AF",X"FF",X"22",X"FF",X"DB",X"FF",X"C1",X"FE",
		X"F0",X"02",X"73",X"04",X"74",X"FF",X"93",X"FF",X"56",X"FF",X"7D",X"FF",X"6D",X"FF",X"6B",X"FF",
		X"83",X"FF",X"51",X"FF",X"A9",X"FF",X"17",X"FF",X"EE",X"03",X"70",X"03",X"1F",X"FF",X"B2",X"FF",
		X"3F",X"FF",X"96",X"FF",X"58",X"FF",X"82",X"FF",X"6B",X"FF",X"70",X"FF",X"83",X"FF",X"6A",X"FF",
		X"60",X"04",X"F1",X"02",X"0B",X"FF",X"C0",X"FF",X"32",X"FF",X"A6",X"FF",X"43",X"FF",X"9D",X"FF",
		X"4A",X"FF",X"9C",X"FF",X"43",X"FF",X"17",X"00",X"18",X"05",X"D0",X"01",X"12",X"FF",X"B8",X"FF",
		X"34",X"FF",X"AD",X"FF",X"38",X"FF",X"B4",X"FF",X"28",X"FF",X"D5",X"FF",X"DA",X"FE",X"42",X"02",
		X"97",X"04",X"B6",X"FF",X"8E",X"FF",X"5B",X"FF",X"89",X"FF",X"61",X"FF",X"85",X"FF",X"63",X"FF",
		X"8A",X"FF",X"52",X"FF",X"1E",X"00",X"2C",X"05",X"54",X"01",X"2B",X"FF",X"A0",X"FF",X"4E",X"FF",
		X"98",X"FF",X"4F",X"FF",X"9F",X"FF",X"41",X"FF",X"BD",X"FF",X"09",X"FF",X"02",X"04",X"E7",X"02",
		X"FA",X"FE",X"CA",X"FF",X"2C",X"FF",X"B6",X"FF",X"35",X"FF",X"BB",X"FF",X"25",X"FF",X"DF",X"FF",
		X"D0",X"FE",X"78",X"03",X"D7",X"03",X"0C",X"FF",X"CB",X"FF",X"2F",X"FF",X"B2",X"FF",X"3D",X"FF",
		X"B1",X"FF",X"36",X"FF",X"CA",X"FF",X"F4",X"FE",X"45",X"01",X"D0",X"04",X"13",X"00",X"6E",X"FF",
		X"77",X"FF",X"73",X"FF",X"7D",X"FF",X"6B",X"FF",X"8B",X"FF",X"5A",X"FF",X"AA",X"FF",X"24",X"FF",
		X"06",X"04",X"F6",X"02",X"F8",X"FE",X"D1",X"FF",X"2C",X"FF",X"B8",X"FF",X"3C",X"FF",X"B2",X"FF",
		X"3D",X"FF",X"BB",X"FF",X"20",X"FF",X"8D",X"00",X"2B",X"05",X"41",X"01",X"26",X"FF",X"B5",X"FF",
		X"3E",X"FF",X"B0",X"FF",X"3F",X"FF",X"B9",X"FF",X"30",X"FF",X"D3",X"FF",X"F2",X"FE",X"4B",X"01",
		X"0D",X"05",X"71",X"00",X"4C",X"FF",X"9A",X"FF",X"55",X"FF",X"A2",X"FF",X"4B",X"FF",X"B0",X"FF",
		X"37",X"FF",X"D3",X"FF",X"E6",X"FE",X"B8",X"01",X"DB",X"04",X"F7",X"FF",X"6F",X"FF",X"80",X"FF",
		X"6C",X"FF",X"8F",X"FF",X"5D",X"FF",X"A1",X"FF",X"46",X"FF",X"C9",X"FF",X"FB",X"FE",X"72",X"03",
		X"A0",X"03",X"34",X"FF",X"BE",X"FF",X"44",X"FF",X"A9",X"FF",X"4F",X"FF",X"A4",X"FF",X"51",X"FF",
		X"B0",X"FF",X"2D",X"FF",X"A7",X"00",X"EB",X"04",X"B4",X"00",X"50",X"FF",X"94",X"FF",X"63",X"FF",
		X"93",X"FF",X"5F",X"FF",X"9F",X"FF",X"4E",X"FF",X"C2",X"FF",X"0B",X"FF",X"8C",X"03",X"79",X"03",
		X"25",X"FF",X"CA",X"FF",X"3C",X"FF",X"B2",X"FF",X"4E",X"FF",X"A6",X"FF",X"57",X"FF",X"A1",X"FF",
		X"57",X"FF",X"E4",X"FF",X"A4",X"04",X"BE",X"01",X"00",X"FF",X"D4",X"FF",X"30",X"FF",X"C4",X"FF",
		X"39",X"FF",X"C4",X"FF",X"33",X"FF",X"D4",X"FF",X"09",X"FF",X"EC",X"00",X"C0",X"04",X"D7",X"00",
		X"30",X"FF",X"B8",X"FF",X"44",X"FF",X"BA",X"FF",X"40",X"FF",X"C4",X"FF",X"31",X"FF",X"DF",X"FF",
		X"F4",X"FE",X"68",X"01",X"BA",X"04",X"7B",X"00",X"4B",X"FF",X"A9",X"FF",X"52",X"FF",X"AF",X"FF",
		X"49",X"FF",X"BB",X"FF",X"39",X"FF",X"DA",X"FF",X"FA",X"FE",X"4F",X"01",X"B2",X"04",X"75",X"00",
		X"4B",X"FF",X"A8",X"FF",X"54",X"FF",X"AE",X"FF",X"4B",X"FF",X"BD",X"FF",X"3A",X"FF",X"DA",X"FF",
		X"FB",X"FE",X"1E",X"01",X"B9",X"04",X"75",X"00",X"48",X"FF",X"AD",X"FF",X"52",X"FF",X"B3",X"FF",
		X"4A",X"FF",X"BF",X"FF",X"3B",X"FF",X"DD",X"FF",X"FB",X"FE",X"32",X"01",X"C9",X"04",X"6E",X"00",
		X"46",X"FF",X"AF",X"FF",X"51",X"FF",X"B3",X"FF",X"48",X"FF",X"C1",X"FF",X"39",X"FF",X"DF",X"FF",
		X"FB",X"FE",X"43",X"01",X"DE",X"04",X"6F",X"00",X"4C",X"FF",X"AD",X"FF",X"53",X"FF",X"B4",X"FF",
		X"4B",X"FF",X"C1",X"FF",X"3A",X"FF",X"DF",X"FF",X"F9",X"FE",X"53",X"01",X"FF",X"04",X"76",X"00",
		X"57",X"FF",X"A6",X"FF",X"5C",X"FF",X"AE",X"FF",X"55",X"FF",X"BA",X"FF",X"43",X"FF",X"D9",X"FF",
		X"00",X"FF",X"57",X"01",X"E0",X"04",X"5E",X"00",X"5F",X"FF",X"A0",X"FF",X"63",X"FF",X"AA",X"FF",
		X"56",X"FF",X"BC",X"FF",X"3E",X"FF",X"E6",X"FF",X"E0",X"FE",X"75",X"02",X"0C",X"04",X"6D",X"FF",
		X"AE",X"FF",X"62",X"FF",X"9B",X"FF",X"73",X"FF",X"92",X"FF",X"7C",X"FF",X"8C",X"FF",X"7D",X"FF",
		X"CC",X"FF",X"90",X"04",X"6E",X"01",X"26",X"FF",X"C0",X"FF",X"52",X"FF",X"B3",X"FF",X"56",X"FF",
		X"BB",X"FF",X"46",X"FF",X"DE",X"FF",X"F1",X"FE",X"1A",X"03",X"40",X"03",X"16",X"FF",X"DE",X"FF",
		X"3C",X"FF",X"C7",X"FF",X"47",X"FF",X"CA",X"FF",X"3C",X"FF",X"E8",X"FF",X"ED",X"FE",X"1A",X"02",
		X"3F",X"04",X"6F",X"FF",X"BA",X"FF",X"57",X"FF",X"B0",X"FF",X"5D",X"FF",X"B3",X"FF",X"54",X"FF",
		X"CD",X"FF",X"15",X"FF",X"4C",X"01",X"AE",X"04",X"B9",X"FF",X"9E",X"FF",X"6A",X"FF",X"A2",X"FF",
		X"6C",X"FF",X"A4",X"FF",X"67",X"FF",X"B4",X"FF",X"3D",X"FF",X"AF",X"00",X"9D",X"04",X"27",X"00",
		X"7F",X"FF",X"83",X"FF",X"90",X"FF",X"80",X"FF",X"95",X"FF",X"78",X"FF",X"A3",X"FF",X"56",X"FF",
		X"62",X"00",X"95",X"04",X"57",X"00",X"72",X"FF",X"8B",X"FF",X"8A",X"FF",X"84",X"FF",X"91",X"FF",
		X"7D",X"FF",X"9D",X"FF",X"60",X"FF",X"51",X"00",X"9A",X"04",X"5B",X"00",X"71",X"FF",X"8C",X"FF",
		X"8C",X"FF",X"83",X"FF",X"95",X"FF",X"7B",X"FF",X"A4",X"FF",X"58",X"FF",X"6E",X"00",X"A8",X"04",
		X"48",X"00",X"72",X"FF",X"8F",X"FF",X"87",X"FF",X"8A",X"FF",X"8A",X"FF",X"8B",X"FF",X"8C",X"FF",
		X"85",X"FF",X"C5",X"FF",X"58",X"04",X"2B",X"01",X"37",X"FF",X"C1",X"FF",X"5A",X"FF",X"B9",X"FF",
		X"5B",X"FF",X"C2",X"FF",X"4A",X"FF",X"E6",X"FF",X"FC",X"FE",X"48",X"03",X"3E",X"03",X"20",X"FF",
		X"D8",X"FF",X"50",X"FF",X"BD",X"FF",X"61",X"FF",X"B4",X"FF",X"67",X"FF",X"B6",X"FF",X"53",X"FF",
		X"41",X"00",X"74",X"04",X"DE",X"00",X"45",X"FF",X"BC",X"FF",X"60",X"FF",X"B8",X"FF",X"5E",X"FF",
		X"C1",X"FF",X"4D",X"FF",X"E4",X"FF",X"05",X"FF",X"77",X"03",X"F4",X"02",X"07",X"FF",X"E8",X"FF",
		X"44",X"FF",X"CD",X"FF",X"50",X"FF",X"CC",X"FF",X"47",X"FF",X"E9",X"FF",X"FE",X"FE",X"C4",X"01",
		X"24",X"04",X"97",X"FF",X"B0",X"FF",X"6F",X"FF",X"A6",X"FF",X"7A",X"FF",X"9F",X"FF",X"7F",X"FF",
		X"9D",X"FF",X"7E",X"FF",X"D0",X"FF",X"3F",X"04",X"51",X"01",X"2B",X"FF",X"D2",X"FF",X"53",X"FF",
		X"C8",X"FF",X"54",X"FF",X"D0",X"FF",X"44",X"FF",X"F4",X"FF",X"F0",X"FE",X"FF",X"01",X"16",X"04",
		X"A6",X"FF",X"9E",X"FF",X"87",X"FF",X"8C",X"FF",X"9B",X"FF",X"79",X"FF",X"B2",X"FF",X"5E",X"FF",
		X"DC",X"FF",X"0E",X"FF",X"33",X"03",X"1C",X"03",X"37",X"FF",X"D0",X"FF",X"64",X"FF",X"AD",X"FF",
		X"7D",X"FF",X"99",X"FF",X"94",X"FF",X"80",X"FF",X"B5",X"FF",X"57",X"FF",X"E3",X"03",X"88",X"02",
		X"1C",X"FF",X"DE",X"FF",X"56",X"FF",X"BD",X"FF",X"6E",X"FF",X"AB",X"FF",X"80",X"FF",X"9A",X"FF",
		X"99",X"FF",X"8F",X"FF",X"1A",X"04",X"26",X"02",X"0A",X"FF",X"EF",X"FF",X"44",X"FF",X"D5",X"FF",
		X"52",X"FF",X"CE",X"FF",X"56",X"FF",X"D6",X"FF",X"3A",X"FF",X"87",X"00",X"53",X"04",X"A7",X"00",
		X"50",X"FF",X"C2",X"FF",X"65",X"FF",X"C1",X"FF",X"62",X"FF",X"CA",X"FF",X"51",X"FF",X"ED",X"FF",
		X"04",X"FF",X"1F",X"03",X"F5",X"02",X"27",X"FF",X"DF",X"FF",X"54",X"FF",X"C5",X"FF",X"63",X"FF",
		X"C2",X"FF",X"62",X"FF",X"CD",X"FF",X"41",X"FF",X"93",X"00",X"58",X"04",X"93",X"00",X"56",X"FF",
		X"C0",X"FF",X"67",X"FF",X"C2",X"FF",X"60",X"FF",X"D3",X"FF",X"46",X"FF",X"FD",X"FF",X"ED",X"FE",
		X"78",X"02",X"D1",X"03",X"67",X"FF",X"B8",X"FF",X"7E",X"FF",X"98",X"FF",X"9A",X"FF",X"82",X"FF",
		X"B4",X"FF",X"64",X"FF",X"E1",X"FF",X"10",X"FF",X"43",X"03",X"1D",X"03",X"2E",X"FF",X"D4",X"FF",
		X"6A",X"FF",X"AE",X"FF",X"88",X"FF",X"96",X"FF",X"A1",X"FF",X"79",X"FF",X"CB",X"FF",X"32",X"FF",
		X"87",X"03",X"CA",X"02",X"1E",X"FF",X"DF",X"FF",X"61",X"FF",X"B9",X"FF",X"7D",X"FF",X"A3",X"FF",
		X"96",X"FF",X"88",X"FF",X"BB",X"FF",X"4B",X"FF",X"A1",X"03",X"AC",X"02",X"0A",X"FF",X"F6",X"FF",
		X"4B",X"FF",X"D2",X"FF",X"63",X"FF",X"C2",X"FF",X"71",X"FF",X"B9",X"FF",X"77",X"FF",X"DB",X"FF",
		X"01",X"04",X"49",X"01",X"2A",X"FF",X"E4",X"FF",X"52",X"FF",X"D6",X"FF",X"56",X"FF",X"DC",X"FF",
		X"48",X"FF",X"FE",X"FF",X"F6",X"FE",X"25",X"02",X"88",X"03",X"62",X"FF",X"CE",X"FF",X"6F",X"FF",
		X"B7",X"FF",X"7D",X"FF",X"AD",X"FF",X"85",X"FF",X"AA",X"FF",X"88",X"FF",X"CF",X"FF",X"01",X"04",
		X"5D",X"01",X"2A",X"FF",X"E7",X"FF",X"55",X"FF",X"D9",X"FF",X"57",X"FF",X"E2",X"FF",X"47",X"FF",
		X"FF",X"FF",X"05",X"FF",X"7F",X"01",X"4C",X"04",X"EB",X"FF",X"86",X"FF",X"AE",X"FF",X"7C",X"FF",
		X"BE",X"FF",X"6A",X"FF",X"D2",X"FF",X"50",X"FF",X"FD",X"FF",X"FA",X"FE",X"3B",X"02",X"B0",X"03",
		X"8C",X"FF",X"AD",X"FF",X"92",X"FF",X"94",X"FF",X"AB",X"FF",X"7E",X"FF",X"C4",X"FF",X"60",X"FF",
		X"F3",X"FF",X"03",X"FF",X"89",X"02",X"75",X"03",X"65",X"FF",X"C4",X"FF",X"82",X"FF",X"A3",X"FF",
		X"9C",X"FF",X"8D",X"FF",X"B6",X"FF",X"6E",X"FF",X"E5",X"FF",X"12",X"FF",X"A2",X"02",X"6C",X"03",
		X"47",X"FF",X"DA",X"FF",X"6E",X"FF",X"B8",X"FF",X"88",X"FF",X"A4",X"FF",X"9E",X"FF",X"8C",X"FF",
		X"C3",X"FF",X"46",X"FF",X"5E",X"03",X"33",X"02",X"10",X"FF",X"FC",X"FF",X"4C",X"FF",X"E1",X"FF",
		X"5D",X"FF",X"DC",X"FF",X"58",X"FF",X"EE",X"FF",X"26",X"FF",X"04",X"01",X"EE",X"03",X"E9",X"FF",
		X"9B",X"FF",X"9D",X"FF",X"99",X"FF",X"A1",X"FF",X"94",X"FF",X"AA",X"FF",X"8C",X"FF",X"B6",X"FF",
		X"93",X"FF",X"F9",X"03",X"4D",X"01",X"31",X"FF",X"E0",X"FF",X"65",X"FF",X"CE",X"FF",X"6B",X"FF",
		X"D3",X"FF",X"60",X"FF",X"F0",X"FF",X"1D",X"FF",X"13",X"03",X"7B",X"02",X"20",X"FF",X"F3",X"FF",
		X"58",X"FF",X"DA",X"FF",X"60",X"FF",X"DF",X"FF",X"53",X"FF",X"03",X"00",X"FE",X"FE",X"67",X"02",
		X"82",X"03",X"38",X"FF",X"E9",X"FF",X"61",X"FF",X"D0",X"FF",X"71",X"FF",X"C9",X"FF",X"76",X"FF",
		X"CD",X"FF",X"60",X"FF",X"5C",X"00",X"21",X"04",X"A3",X"00",X"5A",X"FF",X"D0",X"FF",X"70",X"FF",
		X"D0",X"FF",X"6B",X"FF",X"DC",X"FF",X"54",X"FF",X"05",X"00",X"FC",X"FE",X"71",X"02",X"7F",X"03",
		X"4E",X"FF",X"D3",X"FF",X"7E",X"FF",X"B3",X"FF",X"97",X"FF",X"9D",X"FF",X"AE",X"FF",X"83",X"FF",
		X"D5",X"FF",X"40",X"FF",X"3F",X"03",X"7A",X"02",X"2A",X"FF",X"EA",X"FF",X"6B",X"FF",X"C7",X"FF",
		X"84",X"FF",X"B3",X"FF",X"99",X"FF",X"9D",X"FF",X"B6",X"FF",X"77",X"FF",X"8D",X"03",X"EF",X"01",
		X"2B",X"FF",X"EC",X"FF",X"69",X"FF",X"CB",X"FF",X"80",X"FF",X"B9",X"FF",X"92",X"FF",X"A7",X"FF",
		X"AA",X"FF",X"91",X"FF",X"A8",X"03",X"D1",X"01",X"2E",X"FF",X"EB",X"FF",X"69",X"FF",X"CC",X"FF",
		X"80",X"FF",X"BC",X"FF",X"91",X"FF",X"AA",X"FF",X"A9",X"FF",X"96",X"FF",X"B4",X"03",X"DF",X"01",
		X"28",X"FF",X"F1",X"FF",X"63",X"FF",X"D3",X"FF",X"7A",X"FF",X"C3",X"FF",X"8C",X"FF",X"B1",X"FF",
		X"A1",X"FF",X"A6",X"FF",X"C1",X"03",X"D3",X"01",X"18",X"FF",X"02",X"00",X"54",X"FF",X"E6",X"FF",
		X"64",X"FF",X"DE",X"FF",X"68",X"FF",X"E4",X"FF",X"54",X"FF",X"5C",X"00",X"D4",X"03",X"88",X"00",
		X"5D",X"FF",X"DA",X"FF",X"71",X"FF",X"D7",X"FF",X"6E",X"FF",X"E0",X"FF",X"5D",X"FF",X"05",X"00",
		X"0A",X"FF",X"9D",X"02",X"B6",X"02",X"34",X"FF",X"EE",X"FF",X"69",X"FF",X"D5",X"FF",X"76",X"FF",
		X"D2",X"FF",X"72",X"FF",X"E5",X"FF",X"41",X"FF",X"E5",X"00",X"DA",X"03",X"C2",X"FF",X"B4",X"FF",
		X"94",X"FF",X"B1",X"FF",X"9A",X"FF",X"AE",X"FF",X"9D",X"FF",X"AF",X"FF",X"95",X"FF",X"FA",X"FF",
		X"D4",X"03",X"AA",X"00",X"6A",X"FF",X"C9",X"FF",X"89",X"FF",X"BF",X"FF",X"8B",X"FF",X"C1",X"FF",
		X"86",X"FF",X"CF",X"FF",X"82",X"FF",X"C2",X"03",X"5C",X"01",X"3F",X"FF",X"E6",X"FF",X"72",X"FF",
		X"D5",X"FF",X"7A",X"FF",X"D6",X"FF",X"6F",X"FF",X"EE",X"FF",X"41",X"FF",X"9D",X"03",X"C4",X"01",
		X"2C",X"FF",X"F3",X"FF",X"68",X"FF",X"DB",X"FF",X"73",X"FF",X"DD",X"FF",X"68",X"FF",X"FB",X"FF",
		X"28",X"FF",X"46",X"03",X"0B",X"02",X"22",X"FF",X"FE",X"FF",X"61",X"FF",X"E4",X"FF",X"6B",X"FF",
		X"E6",X"FF",X"60",X"FF",X"05",X"00",X"10",X"FF",X"22",X"02",X"00",X"03",X"4A",X"FF",X"E8",X"FF",
		X"76",X"FF",X"CE",X"FF",X"87",X"FF",X"C5",X"FF",X"8C",X"FF",X"C4",X"FF",X"89",X"FF",X"05",X"00",
		X"BA",X"03",X"C7",X"00",X"59",X"FF",X"DF",X"FF",X"76",X"FF",X"D9",X"FF",X"76",X"FF",X"E2",X"FF",
		X"66",X"FF",X"02",X"00",X"19",X"FF",X"08",X"02",X"29",X"03",X"5C",X"FF",X"E3",X"FF",X"7C",X"FF",
		X"CB",X"FF",X"8C",X"FF",X"C3",X"FF",X"91",X"FF",X"C7",X"FF",X"83",X"FF",X"29",X"00",X"B9",X"03",
		X"60",X"00",X"7B",X"FF",X"C7",X"FF",X"90",X"FF",X"C1",X"FF",X"90",X"FF",X"C9",X"FF",X"83",X"FF",
		X"E3",X"FF",X"53",X"FF",X"73",X"03",X"D4",X"01",X"23",X"FF",X"03",X"00",X"5F",X"FF",X"ED",X"FF",
		X"68",X"FF",X"EF",X"FF",X"5D",X"FF",X"0B",X"00",X"19",X"FF",X"91",X"01",X"AA",X"03",X"9F",X"FF",
		X"C0",X"FF",X"A0",X"FF",X"AA",X"FF",X"B5",X"FF",X"9A",X"FF",X"C7",X"FF",X"80",X"FF",X"F1",X"FF",
		X"2B",X"FF",X"DA",X"02",X"35",X"02",X"1A",X"FF",X"05",X"00",X"66",X"FF",X"E4",X"FF",X"78",X"FF",
		X"D8",X"FF",X"7F",X"FF",X"DB",X"FF",X"73",X"FF",X"47",X"00",X"AB",X"03",X"80",X"00",X"70",X"FF",
		X"D7",X"FF",X"83",X"FF",X"D4",X"FF",X"82",X"FF",X"DD",X"FF",X"72",X"FF",X"FD",X"FF",X"26",X"FF",
		X"B3",X"02",X"3E",X"02",X"23",X"FF",X"04",X"00",X"67",X"FF",X"E9",X"FF",X"73",X"FF",X"E8",X"FF",
		X"6C",X"FF",X"FE",X"FF",X"33",X"FF",X"1C",X"01",X"83",X"03",X"A9",X"FF",X"C0",X"FF",X"A2",X"FF",
		X"B1",X"FF",X"B0",X"FF",X"A3",X"FF",X"C2",X"FF",X"8D",X"FF",X"E4",X"FF",X"4A",X"FF",X"16",X"03",
		X"CD",X"01",X"25",X"FF",X"05",X"00",X"68",X"FF",X"E7",X"FF",X"7A",X"FF",X"DE",X"FF",X"80",X"FF",
		X"E1",X"FF",X"6E",X"FF",X"5A",X"00",X"AE",X"03",X"89",X"00",X"6D",X"FF",X"E0",X"FF",X"7E",X"FF",
		X"DF",X"FF",X"7B",X"FF",X"EA",X"FF",X"67",X"FF",X"0F",X"00",X"14",X"FF",X"38",X"02",X"15",X"03",
		X"49",X"FF",X"F5",X"FF",X"7B",X"FF",X"D9",X"FF",X"8B",X"FF",X"CD",X"FF",X"91",X"FF",X"D1",X"FF",
		X"82",X"FF",X"47",X"00",X"AF",X"03",X"5C",X"00",X"85",X"FF",X"CA",X"FF",X"95",X"FF",X"C8",X"FF",
		X"96",X"FF",X"CE",X"FF",X"8B",X"FF",X"E6",X"FF",X"5A",X"FF",X"28",X"03",X"71",X"01",X"39",X"FF",
		X"FB",X"FF",X"73",X"FF",X"E7",X"FF",X"7B",X"FF",X"EA",X"FF",X"6F",X"FF",X"05",X"00",X"2D",X"FF",
		X"A0",X"02",X"2B",X"02",X"2F",X"FF",X"04",X"00",X"6F",X"FF",X"EC",X"FF",X"7A",X"FF",X"EC",X"FF",
		X"6D",X"FF",X"0B",X"00",X"22",X"FF",X"33",X"02",X"B5",X"02",X"35",X"FF",X"07",X"00",X"6C",X"FF",
		X"EE",X"FF",X"76",X"FF",X"F0",X"FF",X"6B",X"FF",X"0E",X"00",X"20",X"FF",X"F5",X"01",X"F5",X"02",
		X"40",X"FF",X"02",X"00",X"6F",X"FF",X"EC",X"FF",X"7A",X"FF",X"EC",X"FF",X"6F",X"FF",X"0B",X"00",
		X"26",X"FF",X"CF",X"01",X"06",X"03",X"46",X"FF",X"00",X"00",X"73",X"FF",X"EB",X"FF",X"7C",X"FF",
		X"E9",X"FF",X"75",X"FF",X"03",X"00",X"37",X"FF",X"38",X"01",X"5B",X"03",X"86",X"FF",X"DE",X"FF",
		X"8F",X"FF",X"CE",X"FF",X"9D",X"FF",X"C5",X"FF",X"A4",X"FF",X"C1",X"FF",X"A7",X"FF",X"E2",X"FF",
		X"87",X"03",X"E8",X"00",X"56",X"FF",X"F5",X"FF",X"79",X"FF",X"EC",X"FF",X"77",X"FF",X"F4",X"FF",
		X"68",X"FF",X"14",X"00",X"20",X"FF",X"95",X"01",X"44",X"03",X"8C",X"FF",X"D0",X"FF",X"A5",X"FF",
		X"B4",X"FF",X"BC",X"FF",X"A2",X"FF",X"D1",X"FF",X"87",X"FF",X"F9",X"FF",X"39",X"FF",X"8F",X"02",
		X"56",X"02",X"44",X"FF",X"F7",X"FF",X"85",X"FF",X"D4",X"FF",X"A1",X"FF",X"BE",X"FF",X"B7",X"FF",
		X"A7",X"FF",X"D8",X"FF",X"6B",X"FF",X"E7",X"02",X"CA",X"01",X"30",X"FF",X"0B",X"00",X"71",X"FF",
		X"ED",X"FF",X"84",X"FF",X"E0",X"FF",X"90",X"FF",X"DB",X"FF",X"91",X"FF",X"00",X"00",X"84",X"03",
		X"C4",X"00",X"5C",X"FF",X"F8",X"FF",X"79",X"FF",X"EF",X"FF",X"7A",X"FF",X"F8",X"FF",X"6A",X"FF",
		X"19",X"00",X"1B",X"FF",X"DC",X"01",X"CA",X"02",X"50",X"FF",X"F8",X"FF",X"84",X"FF",X"DD",X"FF",
		X"95",X"FF",X"D4",X"FF",X"9B",X"FF",X"D6",X"FF",X"8F",X"FF",X"22",X"00",X"9F",X"03",X"7A",X"00",
		X"7B",X"FF",X"E3",X"FF",X"8D",X"FF",X"E2",X"FF",X"88",X"FF",X"EF",X"FF",X"75",X"FF",X"12",X"00",
		X"25",X"FF",X"B3",X"01",X"D8",X"02",X"6A",X"FF",X"E1",X"FF",X"9E",X"FF",X"C2",X"FF",X"B8",X"FF",
		X"AD",X"FF",X"CF",X"FF",X"92",X"FF",X"F7",X"FF",X"45",X"FF",X"D7",X"02",X"23",X"02",X"3D",X"FF",
		X"01",X"00",X"85",X"FF",X"DB",X"FF",X"A0",X"FF",X"C6",X"FF",X"B4",X"FF",X"B0",X"FF",X"D4",X"FF",
		X"83",X"FF",X"15",X"03",X"A1",X"01",X"43",X"FF",X"01",X"00",X"82",X"FF",X"E2",X"FF",X"99",X"FF",
		X"CF",X"FF",X"AC",X"FF",X"BD",X"FF",X"C7",X"FF",X"9A",X"FF",X"27",X"03",X"8A",X"01",X"3E",X"FF",
		X"0C",X"00",X"75",X"FF",X"F0",X"FF",X"88",X"FF",X"E6",X"FF",X"91",X"FF",X"E1",X"FF",X"92",X"FF",
		X"0D",X"00",X"3B",X"03",X"AC",X"00",X"61",X"FF",X"FB",X"FF",X"80",X"FF",X"F2",X"FF",X"80",X"FF",
		X"F8",X"FF",X"72",X"FF",X"13",X"00",X"30",X"FF",X"B3",X"01",X"D0",X"02",X"69",X"FF",X"EF",X"FF",
		X"94",X"FF",X"D5",X"FF",X"A5",X"FF",X"CA",X"FF",X"AC",X"FF",X"C6",X"FF",X"B0",X"FF",X"E3",X"FF",
		X"41",X"03",X"C3",X"00",X"64",X"FF",X"F6",X"FF",X"84",X"FF",X"EE",X"FF",X"84",X"FF",X"F7",X"FF",
		X"76",X"FF",X"14",X"00",X"37",X"FF",X"4A",X"01",X"35",X"03",X"A1",X"FF",X"D0",X"FF",X"B1",X"FF",
		X"B9",X"FF",X"C5",X"FF",X"A8",X"FF",X"D8",X"FF",X"8F",X"FF",X"00",X"00",X"43",X"FF",X"32",X"02",
		X"54",X"02",X"41",X"FF",X"06",X"00",X"86",X"FF",X"E5",X"FF",X"9A",X"FF",X"D7",X"FF",X"A8",X"FF",
		X"CC",X"FF",X"B1",X"FF",X"DB",X"FF",X"58",X"03",X"C8",X"00",X"68",X"FF",X"F6",X"FF",X"89",X"FF",
		X"EE",X"FF",X"8A",X"FF",X"F1",X"FF",X"7C",X"FF",X"10",X"00",X"35",X"FF",X"16",X"02",X"5A",X"02",
		X"41",X"FF",X"0A",X"00",X"7F",X"FF",X"EE",X"FF",X"8E",X"FF",X"E9",X"FF",X"90",X"FF",X"EF",X"FF",
		X"7B",X"FF",X"6F",X"00",X"2C",X"03",X"1F",X"00",X"96",X"FF",X"DD",X"FF",X"99",X"FF",X"E3",X"FF",
		X"91",X"FF",X"F1",X"FF",X"7B",X"FF",X"19",X"00",X"2C",X"FF",X"0D",X"02",X"9E",X"02",X"56",X"FF",
		X"FA",X"FF",X"94",X"FF",X"D7",X"FF",X"AC",X"FF",X"C7",X"FF",X"BE",X"FF",X"B2",X"FF",X"DA",X"FF",
		X"83",X"FF",X"C7",X"02",X"65",X"01",X"42",X"FF",X"10",X"00",X"7C",X"FF",X"F9",X"FF",X"86",X"FF",
		X"F6",X"FF",X"83",X"FF",X"06",X"00",X"58",X"FF",X"EA",X"00",X"F7",X"02",X"B3",X"FF",X"CB",X"FF",
		X"B7",X"FF",X"C0",X"FF",X"C1",X"FF",X"BA",X"FF",X"C9",X"FF",X"B1",X"FF",X"D6",X"FF",X"9E",X"FF",
		X"02",X"03",X"E2",X"00",X"6A",X"FF",X"F7",X"FF",X"91",X"FF",X"E9",X"FF",X"95",X"FF",X"EF",X"FF",
		X"89",X"FF",X"0A",X"00",X"4A",X"FF",X"6A",X"02",X"BE",X"01",X"39",X"FF",X"15",X"00",X"7C",X"FF",
		X"FD",X"FF",X"84",X"FF",X"FE",X"FF",X"77",X"FF",X"20",X"00",X"28",X"FF",X"E5",X"01",X"80",X"02",
		X"3B",X"FF",X"15",X"00",X"7B",X"FF",X"FB",X"FF",X"86",X"FF",X"FC",X"FF",X"7E",X"FF",X"15",X"00",
		X"3C",X"FF",X"68",X"01",X"A9",X"02",X"5F",X"FF",X"05",X"00",X"89",X"FF",X"F1",X"FF",X"93",X"FF",
		X"F1",X"FF",X"8A",X"FF",X"08",X"00",X"4D",X"FF",X"2F",X"01",X"C1",X"02",X"6F",X"FF",X"FF",X"FF",
		X"8E",X"FF",X"EF",X"FF",X"94",X"FF",X"F1",X"FF",X"8D",X"FF",X"06",X"00",X"52",X"FF",X"1F",X"01",
		X"C8",X"02",X"73",X"FF",X"FE",X"FF",X"8E",X"FF",X"EE",X"FF",X"95",X"FF",X"F0",X"FF",X"8B",X"FF",
		X"09",X"00",X"51",X"FF",X"1E",X"01",X"CC",X"02",X"68",X"FF",X"05",X"00",X"8B",X"FF",X"F4",X"FF",
		X"91",X"FF",X"F6",X"FF",X"87",X"FF",X"12",X"00",X"45",X"FF",X"46",X"01",X"CF",X"02",X"56",X"FF",
		X"0E",X"00",X"85",X"FF",X"F9",X"FF",X"90",X"FF",X"F9",X"FF",X"84",X"FF",X"13",X"00",X"47",X"FF",
		X"6C",X"01",X"8C",X"02",X"4B",X"FF",X"0F",X"00",X"86",X"FF",X"F8",X"FF",X"8F",X"FF",X"F9",X"FF",
		X"88",X"FF",X"12",X"00",X"49",X"FF",X"95",X"01",X"50",X"02",X"4A",X"FF",X"10",X"00",X"87",X"FF",
		X"F8",X"FF",X"93",X"FF",X"F9",X"FF",X"89",X"FF",X"11",X"00",X"4B",X"FF",X"C5",X"01",X"1E",X"02",
		X"50",X"FF",X"0F",X"00",X"8B",X"FF",X"F8",X"FF",X"93",X"FF",X"F9",X"FF",X"89",X"FF",X"12",X"00",
		X"47",X"FF",X"FC",X"01",X"ED",X"01",X"51",X"FF",X"0F",X"00",X"89",X"FF",X"F9",X"FF",X"92",X"FF",
		X"FC",X"FF",X"86",X"FF",X"19",X"00",X"3E",X"FF",X"37",X"02",X"BC",X"01",X"4A",X"FF",X"14",X"00",
		X"86",X"FF",X"FE",X"FF",X"8D",X"FF",X"00",X"00",X"84",X"FF",X"1F",X"00",X"37",X"FF",X"81",X"02",
		X"82",X"01",X"49",X"FF",X"15",X"00",X"87",X"FF",X"FA",X"FF",X"93",X"FF",X"F9",X"FF",X"8E",X"FF",
		X"0E",X"00",X"5E",X"FF",X"93",X"02",X"1E",X"01",X"5E",X"FF",X"06",X"00",X"96",X"FF",X"EF",X"FF",
		X"A1",X"FF",X"EE",X"FF",X"9E",X"FF",X"F9",X"FF",X"87",X"FF",X"A9",X"02",X"E3",X"00",X"77",X"FF",
		X"F5",X"FF",X"A4",X"FF",X"E3",X"FF",X"AD",X"FF",X"DF",X"FF",X"AC",X"FF",X"E5",X"FF",X"A9",X"FF",
		X"C6",X"02",X"A3",X"00",X"8B",X"FF",X"E8",X"FF",X"AF",X"FF",X"DB",X"FF",X"B5",X"FF",X"D8",X"FF",
		X"B8",X"FF",X"D8",X"FF",X"C4",X"FF",X"EF",X"02",X"60",X"00",X"A4",X"FF",X"D9",X"FF",X"B9",X"FF",
		X"D1",X"FF",X"C0",X"FF",X"CF",X"FF",X"C1",X"FF",X"D2",X"FF",X"C9",X"FF",X"F9",X"02",X"67",X"00",
		X"9A",X"FF",X"E7",X"FF",X"AE",X"FF",X"E0",X"FF",X"AF",X"FF",X"E6",X"FF",X"A4",X"FF",X"FD",X"FF",
		X"74",X"FF",X"65",X"02",X"5D",X"01",X"55",X"FF",X"15",X"00",X"8C",X"FF",X"FE",X"FF",X"95",X"FF",
		X"FD",X"FF",X"91",X"FF",X"0C",X"00",X"6C",X"FF",X"CB",X"00",X"B3",X"02",X"CD",X"FF",X"C4",X"FF",
		X"D4",X"FF",X"B7",X"FF",X"E4",X"FF",X"A8",X"FF",X"F5",X"FF",X"8E",X"FF",X"1E",X"00",X"39",X"FF",
		X"F4",X"01",X"27",X"02",X"57",X"FF",X"0B",X"00",X"9D",X"FF",X"E4",X"FF",X"B8",X"FF",X"D1",X"FF",
		X"CD",X"FF",X"BA",X"FF",X"EE",X"FF",X"7D",X"FF",X"72",X"02",X"73",X"01",X"4B",X"FF",X"1A",X"00",
		X"8E",X"FF",X"FC",X"FF",X"A0",X"FF",X"EE",X"FF",X"AC",X"FF",X"E5",X"FF",X"B7",X"FF",X"E8",X"FF",
		X"AE",X"02",X"BC",X"00",X"70",X"FF",X"0C",X"00",X"91",X"FF",X"01",X"00",X"94",X"FF",X"04",X"00",
		X"8A",X"FF",X"1A",X"00",X"57",X"FF",X"40",X"01",X"63",X"02",X"87",X"FF",X"F1",X"FF",X"B3",X"FF",
		X"DB",X"FF",X"BF",X"FF",X"D3",X"FF",X"C6",X"FF",X"D0",X"FF",X"CA",X"FF",X"E1",X"FF",X"B9",X"02",
		X"88",X"00",X"8D",X"FF",X"F7",X"FF",X"A5",X"FF",X"F0",X"FF",X"A4",X"FF",X"F8",X"FF",X"96",X"FF",
		X"12",X"00",X"5C",X"FF",X"5A",X"01",X"58",X"02",X"7A",X"FF",X"F6",X"FF",X"B3",X"FF",X"D9",X"FF",
		X"CA",X"FF",X"C6",X"FF",X"DD",X"FF",X"AE",X"FF",X"03",X"00",X"5F",X"FF",X"40",X"02",X"9D",X"01",
		X"56",X"FF",X"17",X"00",X"98",X"FF",X"F4",X"FF",X"B0",X"FF",X"E1",X"FF",X"C3",X"FF",X"CC",X"FF",
		X"E0",X"FF",X"99",X"FF",X"AF",X"02",X"1C",X"01",X"5F",X"FF",X"14",X"00",X"95",X"FF",X"F9",X"FF",
		X"A9",X"FF",X"E8",X"FF",X"BA",X"FF",X"D8",X"FF",X"D2",X"FF",X"B6",X"FF",X"C9",X"02",X"EF",X"00",
		X"69",X"FF",X"10",X"00",X"99",X"FF",X"F7",X"FF",X"AA",X"FF",X"E9",X"FF",X"B9",X"FF",X"D8",X"FF",
		X"D2",X"FF",X"AC",X"FF",X"A8",X"02",X"F9",X"00",X"68",X"FF",X"13",X"00",X"97",X"FF",X"FB",X"FF",
		X"A8",X"FF",X"EE",X"FF",X"B7",X"FF",X"DF",X"FF",X"CD",X"FF",X"BC",X"FF",X"93",X"02",X"FC",X"00",
		X"6A",X"FF",X"14",X"00",X"96",X"FF",X"FC",X"FF",X"A6",X"FF",X"F1",X"FF",X"B3",X"FF",X"E3",X"FF",
		X"C5",X"FF",X"CC",X"FF",X"7F",X"02",X"FA",X"00",X"63",X"FF",X"1C",X"00",X"8D",X"FF",X"0A",X"00",
		X"97",X"FF",X"04",X"00",X"9B",X"FF",X"08",X"00",X"91",X"FF",X"40",X"00",X"CF",X"02",X"25",X"00",
		X"A4",X"FF",X"F7",X"FF",X"A5",X"FF",X"FC",X"FF",X"9F",X"FF",X"07",X"00",X"8D",X"FF",X"29",X"00",
		X"3F",X"FF",X"E5",X"01",X"D3",X"01",X"5B",X"FF",X"16",X"00",X"9C",X"FF",X"FB",X"FF",X"AA",X"FF",
		X"F5",X"FF",X"A9",X"FF",X"FD",X"FF",X"90",X"FF",X"8A",X"00",X"96",X"02",X"B8",X"FF",X"E4",X"FF",
		X"C2",X"FF",X"D9",X"FF",X"C8",X"FF",X"D5",X"FF",X"CC",X"FF",X"D5",X"FF",X"CC",X"FF",X"E7",X"FF",
		X"9F",X"02",X"56",X"00",X"A9",X"FF",X"E9",X"FF",X"BB",X"FF",X"E5",X"FF",X"BC",X"FF",X"E8",X"FF",
		X"B6",X"FF",X"F5",X"FF",X"9D",X"FF",X"59",X"02",X"D4",X"00",X"81",X"FF",X"04",X"00",X"A7",X"FF",
		X"F5",X"FF",X"AD",X"FF",X"F9",X"FF",X"A5",X"FF",X"0B",X"00",X"79",X"FF",X"24",X"02",X"21",X"01",
		X"6E",X"FF",X"11",X"00",X"A0",X"FF",X"FE",X"FF",X"A8",X"FF",X"FF",X"FF",X"9F",X"FF",X"15",X"00",
		X"67",X"FF",X"00",X"02",X"55",X"01",X"62",X"FF",X"1A",X"00",X"99",X"FF",X"04",X"00",X"A2",X"FF",
		X"06",X"00",X"98",X"FF",X"1F",X"00",X"58",X"FF",X"6A",X"01",X"11",X"02",X"6D",X"FF",X"11",X"00",
		X"A2",X"FF",X"F7",X"FF",X"B3",X"FF",X"EF",X"FF",X"BB",X"FF",X"EA",X"FF",X"BF",X"FF",X"F1",X"FF",
		X"96",X"02",X"76",X"00",X"93",X"FF",X"04",X"00",X"A6",X"FF",X"FF",X"FF",X"A4",X"FF",X"05",X"00",
		X"9A",X"FF",X"1B",X"00",X"6D",X"FF",X"F6",X"00",X"4A",X"02",X"BC",X"FF",X"DB",X"FF",X"D8",X"FF",
		X"C6",X"FF",X"E8",X"FF",X"B7",X"FF",X"FB",X"FF",X"A1",X"FF",X"1D",X"00",X"5A",X"FF",X"96",X"01",
		X"F0",X"01",X"80",X"FF",X"01",X"00",X"B9",X"FF",X"E0",X"FF",X"D2",X"FF",X"CB",X"FF",X"E7",X"FF",
		X"B3",X"FF",X"0D",X"00",X"64",X"FF",X"EC",X"01",X"A3",X"01",X"5D",X"FF",X"1F",X"00",X"9D",X"FF",
		X"00",X"00",X"B0",X"FF",X"F1",X"FF",X"BD",X"FF",X"E8",X"FF",X"C1",X"FF",X"F6",X"FF",X"65",X"02",
		X"81",X"00",X"94",X"FF",X"03",X"00",X"AA",X"FF",X"FC",X"FF",X"AD",X"FF",X"00",X"00",X"A1",X"FF",
		X"19",X"00",X"6B",X"FF",X"85",X"01",X"C7",X"01",X"73",X"FF",X"13",X"00",X"A7",X"FF",X"FE",X"FF",
		X"AE",X"FF",X"FC",X"FF",X"AC",X"FF",X"09",X"00",X"8A",X"FF",X"89",X"00",X"8B",X"02",X"A5",X"FF",
		X"F3",X"FF",X"BF",X"FF",X"E5",X"FF",X"CB",X"FF",X"E0",X"FF",X"CC",X"FF",X"E0",X"FF",X"C9",X"FF",
		X"04",X"00",X"66",X"02",X"39",X"00",X"B9",X"FF",X"E7",X"FF",X"C8",X"FF",X"E2",X"FF",X"C8",X"FF",
		X"E6",X"FF",X"C3",X"FF",X"EF",X"FF",X"B7",X"FF",X"40",X"02",X"9B",X"00",X"94",X"FF",X"01",X"00",
		X"B3",X"FF",X"F6",X"FF",X"B8",X"FF",X"F8",X"FF",X"B1",X"FF",X"08",X"00",X"8B",X"FF",X"29",X"02",
		X"CD",X"00",X"85",X"FF",X"09",X"00",X"B0",X"FF",X"FA",X"FF",X"B6",X"FF",X"FB",X"FF",X"AE",X"FF",
		X"0F",X"00",X"81",X"FF",X"12",X"02",X"F1",X"00",X"7A",X"FF",X"14",X"00",X"A5",X"FF",X"03",X"00",
		X"AB",X"FF",X"07",X"00",X"A0",X"FF",X"22",X"00",X"5C",X"FF",X"C6",X"01",X"88",X"01",X"63",X"FF",
		X"22",X"00",X"9F",X"FF",X"08",X"00",X"AC",X"FF",X"02",X"00",X"AB",X"FF",X"0A",X"00",X"98",X"FF",
		X"59",X"00",X"82",X"02",X"E9",X"FF",X"CB",X"FF",X"E7",X"FF",X"C3",X"FF",X"F1",X"FF",X"B9",X"FF",
		X"FF",X"FF",X"A7",X"FF",X"1C",X"00",X"6B",X"FF",X"73",X"01",X"C6",X"01",X"8B",X"FF",X"00",X"00",
		X"C2",X"FF",X"E2",X"FF",X"D6",X"FF",X"D1",X"FF",X"EA",X"FF",X"BA",X"FF",X"0F",X"00",X"6F",X"FF",
		X"14",X"02",X"43",X"01",X"6E",X"FF",X"18",X"00",X"AC",X"FF",X"F9",X"FF",X"C1",X"FF",X"E7",X"FF",
		X"D2",X"FF",X"D4",X"FF",X"F1",X"FF",X"97",X"FF",X"35",X"02",X"EA",X"00",X"6A",X"FF",X"28",X"00",
		X"99",X"FF",X"10",X"00",X"A5",X"FF",X"0D",X"00",X"A8",X"FF",X"11",X"00",X"95",X"FF",X"6E",X"00",
		X"3F",X"02",X"05",X"00",X"C5",X"FF",X"ED",X"FF",X"C4",X"FF",X"F1",X"FF",X"BF",X"FF",X"FB",X"FF",
		X"B2",X"FF",X"12",X"00",X"7E",X"FF",X"E4",X"01",X"2A",X"01",X"7E",X"FF",X"15",X"00",X"AC",X"FF",
		X"02",X"00",X"B3",X"FF",X"01",X"00",X"B2",X"FF",X"0E",X"00",X"93",X"FF",X"90",X"00",X"3C",X"02",
		X"D8",X"FF",X"E0",X"FF",X"DB",X"FF",X"D3",X"FF",X"E8",X"FF",X"C6",X"FF",X"F7",X"FF",X"B4",X"FF",
		X"14",X"00",X"79",X"FF",X"76",X"01",X"A7",X"01",X"79",X"FF",X"13",X"00",X"B6",X"FF",X"F4",X"FF",
		X"CC",X"FF",X"E2",X"FF",X"DC",X"FF",X"D1",X"FF",X"F7",X"FF",X"9E",X"FF",X"F9",X"01",X"13",X"01",
		X"80",X"FF",X"15",X"00",X"B3",X"FF",X"FC",X"FF",X"C4",X"FF",X"ED",X"FF",X"D1",X"FF",X"DE",X"FF",
		X"E7",X"FF",X"BA",X"FF",X"26",X"02",X"D1",X"00",X"8B",X"FF",X"10",X"00",X"B5",X"FF",X"FB",X"FF",
		X"C3",X"FF",X"EE",X"FF",X"D1",X"FF",X"E1",X"FF",X"E4",X"FF",X"C4",X"FF",X"1D",X"02",X"CF",X"00",
		X"8E",X"FF",X"0F",X"00",X"B5",X"FF",X"FB",X"FF",X"C4",X"FF",X"ED",X"FF",X"D3",X"FF",X"DE",X"FF",
		X"E5",X"FF",X"C0",X"FF",X"0C",X"02",X"DB",X"00",X"87",X"FF",X"13",X"00",X"B4",X"FF",X"FD",X"FF",
		X"C4",X"FF",X"EF",X"FF",X"D3",X"FF",X"DE",X"FF",X"EA",X"FF",X"B8",X"FF",X"02",X"02",X"E9",X"00",
		X"7B",X"FF",X"1E",X"00",X"AA",X"FF",X"08",X"00",X"B9",X"FF",X"FD",X"FF",X"C6",X"FF",X"F2",X"FF",
		X"D3",X"FF",X"E3",X"FF",X"08",X"02",X"AA",X"00",X"87",X"FF",X"1E",X"00",X"A5",X"FF",X"12",X"00",
		X"AA",X"FF",X"14",X"00",X"A4",X"FF",X"22",X"00",X"80",X"FF",X"AB",X"00",X"31",X"02",X"AD",X"FF",
		X"F1",X"FF",X"D6",X"FF",X"DD",X"FF",X"E6",X"FF",X"D2",X"FF",X"F1",X"FF",X"C2",X"FF",X"0F",X"00",
		X"82",X"FF",X"25",X"02",X"F1",X"00",X"77",X"FF",X"22",X"00",X"A7",X"FF",X"0D",X"00",X"B3",X"FF",
		X"08",X"00",X"B4",X"FF",X"0D",X"00",X"A5",X"FF",X"57",X"00",X"1B",X"02",X"17",X"00",X"C3",X"FF",
		X"F9",X"FF",X"C1",X"FF",X"00",X"00",X"BA",X"FF",X"09",X"00",X"AB",X"FF",X"22",X"00",X"79",X"FF",
		X"EB",X"00",X"23",X"02",X"8C",X"FF",X"0A",X"00",X"C7",X"FF",X"EC",X"FF",X"D9",X"FF",X"DD",X"FF",
		X"E7",X"FF",X"CE",X"FF",X"02",X"00",X"9C",X"FF",X"CF",X"01",X"FC",X"00",X"84",X"FF",X"1C",X"00",
		X"AD",X"FF",X"0D",X"00",X"B6",X"FF",X"0C",X"00",X"AF",X"FF",X"1D",X"00",X"86",X"FF",X"CD",X"00",
		X"F3",X"01",X"93",X"FF",X"07",X"00",X"C4",X"FF",X"F4",X"FF",X"D0",X"FF",X"E9",X"FF",X"DC",X"FF",
		X"DE",X"FF",X"F0",X"FF",X"BA",X"FF",X"2F",X"02",X"9A",X"00",X"8D",X"FF",X"1E",X"00",X"AA",X"FF",
		X"12",X"00",X"AF",X"FF",X"14",X"00",X"A9",X"FF",X"24",X"00",X"86",X"FF",X"B4",X"00",X"E8",X"01",
		X"DC",X"FF",X"D9",X"FF",X"F0",X"FF",X"C8",X"FF",X"FF",X"FF",X"BA",X"FF",X"11",X"00",X"A5",X"FF",
		X"33",X"00",X"5F",X"FF",X"53",X"01",X"C4",X"01",X"81",X"FF",X"0D",X"00",X"CA",X"FF",X"E9",X"FF",
		X"E5",X"FF",X"D2",X"FF",X"FA",X"FF",X"BA",X"FF",X"20",X"00",X"74",X"FF",X"63",X"01",X"80",X"01",
		X"7B",X"FF",X"17",X"00",X"BF",X"FF",X"F3",X"FF",X"D9",X"FF",X"DF",X"FF",X"F0",X"FF",X"C7",X"FF",
		X"16",X"00",X"7D",X"FF",X"7B",X"01",X"71",X"01",X"6B",X"FF",X"29",X"00",X"AF",X"FF",X"0A",X"00",
		X"C3",X"FF",X"F9",X"FF",X"D2",X"FF",X"EA",X"FF",X"E5",X"FF",X"D0",X"FF",X"CF",X"01",X"B0",X"00",
		X"94",X"FF",X"18",X"00",X"B3",X"FF",X"0C",X"00",X"BB",X"FF",X"0A",X"00",X"B9",X"FF",X"15",X"00",
		X"99",X"FF",X"B4",X"00",X"C5",X"01",X"B3",X"FF",X"FE",X"FF",X"CF",X"FF",X"F1",X"FF",X"D8",X"FF",
		X"ED",X"FF",X"DA",X"FF",X"EC",X"FF",X"D9",X"FF",X"FA",X"FF",X"F8",X"01",X"30",X"00",X"C2",X"FF",
		X"FB",X"FF",X"CD",X"FF",X"FA",X"FF",X"C9",X"FF",X"01",X"00",X"BF",X"FF",X"18",X"00",X"8B",X"FF",
		X"92",X"01",X"F0",X"00",X"89",X"FF",X"1E",X"00",X"B3",X"FF",X"0D",X"00",X"B9",X"FF",X"12",X"00",
		X"B0",X"FF",X"29",X"00",X"75",X"FF",X"7F",X"01",X"51",X"01",X"7A",X"FF",X"24",X"00",X"B1",X"FF",
		X"0E",X"00",X"C0",X"FF",X"07",X"00",X"BE",X"FF",X"0D",X"00",X"B1",X"FF",X"45",X"00",X"03",X"02",
		X"E5",X"FF",X"DE",X"FF",X"F0",X"FF",X"D4",X"FF",X"F8",X"FF",X"CA",X"FF",X"03",X"00",X"BB",X"FF",
		X"24",X"00",X"79",X"FF",X"9A",X"01",X"3E",X"01",X"7E",X"FF",X"20",X"00",X"BA",X"FF",X"04",X"00",
		X"CC",X"FF",X"F4",X"FF",X"DB",X"FF",X"E6",X"FF",X"EF",X"FF",X"C3",X"FF",X"BA",X"01",X"BA",X"00",
		X"93",X"FF",X"1D",X"00",X"B7",X"FF",X"0B",X"00",X"C5",X"FF",X"02",X"00",X"CB",X"FF",X"FC",X"FF",
		X"CF",X"FF",X"04",X"00",X"DB",X"01",X"64",X"00",X"AF",X"FF",X"0E",X"00",X"C1",X"FF",X"04",X"00",
		X"C8",X"FF",X"00",X"00",X"CE",X"FF",X"FD",X"FF",X"CE",X"FF",X"10",X"00",X"E0",X"01",X"4F",X"00",
		X"B7",X"FF",X"08",X"00",X"C7",X"FF",X"02",X"00",X"CD",X"FF",X"FD",X"FF",X"D2",X"FF",X"F8",X"FF",
		X"D8",X"FF",X"F9",X"FF",X"E1",X"01",X"59",X"00",X"B1",X"FF",X"0D",X"00",X"C5",X"FF",X"04",X"00",
		X"CC",X"FF",X"FF",X"FF",X"D2",X"FF",X"F8",X"FF",X"DB",X"FF",X"E8",X"FF",X"E2",X"01",X"5E",X"00",
		X"AA",X"FF",X"17",X"00",X"BA",X"FF",X"0F",X"00",X"BE",X"FF",X"11",X"00",X"BB",X"FF",X"1A",X"00",
		X"A3",X"FF",X"84",X"00",X"B3",X"01",X"E4",X"FF",X"E4",X"FF",X"EF",X"FF",X"DA",X"FF",X"F7",X"FF",
		X"D3",X"FF",X"00",X"00",X"C5",X"FF",X"14",X"00",X"9D",X"FF",X"69",X"01",X"F3",X"00",X"9A",X"FF",
		X"18",X"00",X"C1",X"FF",X"04",X"00",X"CA",X"FF",X"01",X"00",X"CE",X"FF",X"04",X"00",X"C6",X"FF",
		X"2E",X"00",X"CC",X"01",X"08",X"00",X"D4",X"FF",X"FB",X"FF",X"D0",X"FF",X"02",X"00",X"CB",X"FF",
		X"0E",X"00",X"BA",X"FF",X"26",X"00",X"84",X"FF",X"1E",X"01",X"73",X"01",X"93",X"FF",X"14",X"00",
		X"CE",X"FF",X"F7",X"FF",X"E2",X"FF",X"E6",X"FF",X"F3",X"FF",X"D4",X"FF",X"10",X"00",X"9A",X"FF",
		X"4F",X"01",X"19",X"01",X"83",X"FF",X"2A",X"00",X"B5",X"FF",X"13",X"00",X"C2",X"FF",X"0E",X"00",
		X"C6",X"FF",X"0E",X"00",X"BD",X"FF",X"38",X"00",X"F8",X"01",X"F4",X"FF",X"E0",X"FF",X"F2",X"FF",
		X"DB",X"FF",X"F7",X"FF",X"D8",X"FF",X"FF",X"FF",X"CD",X"FF",X"12",X"00",X"A2",X"FF",X"6B",X"01",
		X"CD",X"00",X"9C",X"FF",X"1D",X"00",X"C0",X"FF",X"0E",X"00",X"C7",X"FF",X"0B",X"00",X"C5",X"FF",
		X"14",X"00",X"B1",X"FF",X"69",X"00",X"A8",X"01",X"D9",X"FF",X"ED",X"FF",X"ED",X"FF",X"DF",X"FF",
		X"F8",X"FF",X"D5",X"FF",X"05",X"00",X"C4",X"FF",X"22",X"00",X"89",X"FF",X"70",X"01",X"28",X"01",
		X"8E",X"FF",X"21",X"00",X"C3",X"FF",X"07",X"00",X"D4",X"FF",X"FC",X"FF",X"DD",X"FF",X"F3",X"FF",
		X"E8",X"FF",X"E8",X"FF",X"96",X"01",X"69",X"00",X"B5",X"FF",X"11",X"00",X"C8",X"FF",X"0A",X"00",
		X"C9",X"FF",X"0B",X"00",X"C3",X"FF",X"1C",X"00",X"9E",X"FF",X"E8",X"00",X"45",X"01",X"A3",X"FF",
		X"15",X"00",X"CA",X"FF",X"05",X"00",X"D2",X"FF",X"02",X"00",X"D3",X"FF",X"07",X"00",X"C4",X"FF",
		X"3C",X"00",X"CA",X"01",X"EF",X"FF",X"E6",X"FF",X"F3",X"FF",X"DF",X"FF",X"FA",X"FF",X"D8",X"FF",
		X"03",X"00",X"CA",X"FF",X"1C",X"00",X"98",X"FF",X"49",X"01",X"02",X"01",X"9A",X"FF",X"19",X"00",
		X"CB",X"FF",X"03",X"00",X"DB",X"FF",X"F6",X"FF",X"E7",X"FF",X"EA",X"FF",X"FB",X"FF",X"C2",X"FF",
		X"81",X"01",X"99",X"00",X"9E",X"FF",X"22",X"00",X"BC",X"FF",X"19",X"00",X"BF",X"FF",X"1A",X"00",
		X"BC",X"FF",X"28",X"00",X"99",X"FF",X"A6",X"00",X"CF",X"01",X"B9",X"FF",X"02",X"00",X"E1",X"FF",
		X"F2",X"FF",X"ED",X"FF",X"E6",X"FF",X"F8",X"FF",X"D9",X"FF",X"0B",X"00",X"AF",X"FF",X"BA",X"01",
		X"91",X"00",X"AB",X"FF",X"19",X"00",X"C9",X"FF",X"0D",X"00",X"CC",X"FF",X"0D",X"00",X"C7",X"FF",
		X"1E",X"00",X"A1",X"FF",X"18",X"01",X"F0",X"00",X"A3",X"FF",X"19",X"00",X"C8",X"FF",X"0A",X"00",
		X"D0",X"FF",X"0C",X"00",X"CC",X"FF",X"18",X"00",X"AB",X"FF",X"92",X"00",X"7C",X"01",X"A5",X"FF",
		X"19",X"00",X"C9",X"FF",X"0C",X"00",X"D0",X"FF",X"0A",X"00",X"CA",X"FF",X"18",X"00",X"AA",X"FF",
		X"95",X"00",X"DC",X"01",X"A5",X"FF",X"19",X"00",X"CC",X"FF",X"0B",X"00",X"D3",X"FF",X"08",X"00",
		X"D0",X"FF",X"11",X"00",X"B8",X"FF",X"72",X"00",X"CF",X"01",X"BB",X"FF",X"0B",X"00",X"D5",X"FF",
		X"02",X"00",X"DA",X"FF",X"02",X"00",X"D7",X"FF",X"0B",X"00",X"C1",X"FF",X"5E",X"00",X"D4",X"01",
		X"C1",X"FF",X"0C",X"00",X"D4",X"FF",X"01",X"00",X"D9",X"FF",X"01",X"00",X"D8",X"FF",X"0D",X"00",
		X"C0",X"FF",X"5D",X"00",X"E5",X"01",X"C1",X"FF",X"0B",X"00",X"D5",X"FF",X"01",X"00",X"D9",X"FF",
		X"02",X"00",X"D8",X"FF",X"0B",X"00",X"C6",X"FF",X"4F",X"00",X"C6",X"01",X"C6",X"FF",X"07",X"00",
		X"D8",X"FF",X"FE",X"FF",X"DD",X"FF",X"01",X"00",X"DC",X"FF",X"06",X"00",X"CC",X"FF",X"3E",X"00",
		X"86",X"01",X"CA",X"FF",X"06",X"00",X"DB",X"FF",X"FE",X"FF",X"E0",X"FF",X"FE",X"FF",X"DC",X"FF",
		X"04",X"00",X"CA",X"FF",X"4C",X"00",X"4F",X"01",X"C1",X"FF",X"0D",X"00",X"D7",X"FF",X"04",X"00",
		X"D9",X"FF",X"05",X"00",X"D6",X"FF",X"12",X"00",X"BA",X"FF",X"8E",X"00",X"2E",X"01",X"B0",X"FF",
		X"14",X"00",X"D3",X"FF",X"09",X"00",X"D8",X"FF",X"06",X"00",X"D4",X"FF",X"11",X"00",X"BD",X"FF",
		X"7A",X"00",X"3E",X"01",X"BA",X"FF",X"0E",X"00",X"DA",X"FF",X"00",X"00",X"E0",X"FF",X"FC",X"FF",
		X"E3",X"FF",X"FC",X"FF",X"E5",X"FF",X"04",X"00",X"C3",X"01",X"25",X"00",X"D6",X"FF",X"04",X"00",
		X"DB",X"FF",X"05",X"00",X"D7",X"FF",X"0D",X"00",X"CC",X"FF",X"22",X"00",X"9D",X"FF",X"09",X"01",
		X"35",X"01",X"9B",X"FF",X"22",X"00",X"C9",X"FF",X"0C",X"00",X"D7",X"FF",X"06",X"00",X"DB",X"FF",
		X"05",X"00",X"D8",X"FF",X"1B",X"00",X"CA",X"01",X"0A",X"00",X"E1",X"FF",X"FB",X"FF",X"E3",X"FF",
		X"FD",X"FF",X"E1",X"FF",X"04",X"00",X"D7",X"FF",X"12",X"00",X"B4",X"FF",X"19",X"01",X"99",X"00",
		X"B1",X"FF",X"1B",X"00",X"CD",X"FF",X"11",X"00",X"CE",X"FF",X"13",X"00",X"C5",X"FF",X"2A",X"00",
		X"8F",X"FF",X"4A",X"01",X"25",X"01",X"92",X"FF",X"2C",X"00",X"C1",X"FF",X"19",X"00",X"C9",X"FF",
		X"19",X"00",X"C4",X"FF",X"28",X"00",X"9E",X"FF",X"F2",X"00",X"26",X"01",X"A8",X"FF",X"1C",X"00",
		X"CF",X"FF",X"0D",X"00",X"D8",X"FF",X"0B",X"00",X"D3",X"FF",X"16",X"00",X"B6",X"FF",X"9F",X"00",
		X"31",X"01",X"B1",X"FF",X"16",X"00",X"D5",X"FF",X"08",X"00",X"DD",X"FF",X"03",X"00",X"DE",X"FF",
		X"03",X"00",X"DC",X"FF",X"12",X"00",X"D4",X"01",X"16",X"00",X"DB",X"FF",X"05",X"00",X"DA",X"FF",
		X"08",X"00",X"D5",X"FF",X"11",X"00",X"C8",X"FF",X"28",X"00",X"98",X"FF",X"15",X"01",X"2A",X"01",
		X"A4",X"FF",X"1B",X"00",X"D6",X"FF",X"03",X"00",X"E5",X"FF",X"F8",X"FF",X"F0",X"FF",X"E9",X"FF",
		X"05",X"00",X"C7",X"FF",X"1D",X"01",X"96",X"00",X"B1",X"FF",X"1D",X"00",X"D0",X"FF",X"0D",X"00",
		X"DA",X"FF",X"07",X"00",X"E0",X"FF",X"01",X"00",X"E6",X"FF",X"FE",X"FF",X"56",X"01",X"3A",X"00",
		X"CB",X"FF",X"11",X"00",X"D7",X"FF",X"0C",X"00",X"DA",X"FF",X"0B",X"00",X"D7",X"FF",X"0E",X"00",
		X"CF",X"FF",X"37",X"00",X"87",X"01",X"01",X"00",X"E8",X"FF",X"FF",X"FF",X"E4",X"FF",X"02",X"00",
		X"DF",X"FF",X"09",X"00",X"D7",X"FF",X"1A",X"00",X"B4",X"FF",X"C2",X"00",X"EA",X"00",X"B4",X"FF",
		X"17",X"00",X"D6",X"FF",X"0A",X"00",X"E1",X"FF",X"03",X"00",X"E2",X"FF",X"06",X"00",X"DD",X"FF",
		X"27",X"00",X"61",X"01",X"FF",X"FF",X"EE",X"FF",X"F9",X"FF",X"EB",X"FF",X"FE",X"FF",X"E6",X"FF",
		X"02",X"00",X"DD",X"FF",X"15",X"00",X"B5",X"FF",X"56",X"01",X"8E",X"00",X"B6",X"FF",X"1D",X"00",
		X"D0",X"FF",X"13",X"00",X"D4",X"FF",X"14",X"00",X"D0",X"FF",X"25",X"00",X"A8",X"FF",X"30",X"01",
		X"C8",X"00",X"B3",X"FF",X"1C",X"00",X"D5",X"FF",X"0E",X"00",X"DB",X"FF",X"0C",X"00",X"D9",X"FF",
		X"16",X"00",X"C4",X"FF",X"6C",X"00",X"04",X"01",X"BE",X"FF",X"11",X"00",X"DF",X"FF",X"03",X"00",
		X"E8",X"FF",X"FE",X"FF",X"EE",X"FF",X"F7",X"FF",X"F5",X"FF",X"E7",X"FF",X"18",X"01",X"47",X"00",
		X"C8",X"FF",X"16",X"00",X"D3",X"FF",X"14",X"00",X"D3",X"FF",X"18",X"00",X"CC",X"FF",X"27",X"00",
		X"B0",X"FF",X"8B",X"00",X"8B",X"01",X"CE",X"FF",X"03",X"00",X"EF",X"FF",X"F2",X"FF",X"FD",X"FF",
		X"E8",X"FF",X"08",X"00",X"DB",X"FF",X"1B",X"00",X"BB",X"FF",X"94",X"00",X"FA",X"00",X"C0",X"FF",
		X"0F",X"00",X"E8",X"FF",X"FA",X"FF",X"F6",X"FF",X"F1",X"FF",X"00",X"00",X"E2",X"FF",X"13",X"00",
		X"BE",X"FF",X"C4",X"00",X"D0",X"00",X"B7",X"FF",X"19",X"00",X"DD",X"FF",X"06",X"00",X"EA",X"FF",
		X"FD",X"FF",X"F2",X"FF",X"F2",X"FF",X"03",X"00",X"D4",X"FF",X"5A",X"01",X"7C",X"00",X"BE",X"FF",
		X"1C",X"00",X"D4",X"FF",X"13",X"00",X"D9",X"FF",X"13",X"00",X"D6",X"FF",X"1D",X"00",X"BE",X"FF",
		X"81",X"00",X"37",X"01",X"CD",X"FF",X"0B",X"00",X"E9",X"FF",X"FD",X"FF",X"F2",X"FF",X"F7",X"FF",
		X"F5",X"FF",X"F2",X"FF",X"FF",X"FF",X"E0",X"FF",X"9B",X"01",X"41",X"00",X"D5",X"FF",X"0D",X"00",
		X"E2",X"FF",X"09",X"00",X"E5",X"FF",X"0A",X"00",X"DE",X"FF",X"15",X"00",X"C4",X"FF",X"F4",X"00",
		X"89",X"00",X"C1",X"FF",X"19",X"00",X"DA",X"FF",X"0F",X"00",X"DD",X"FF",X"11",X"00",X"D6",X"FF",
		X"1E",X"00",X"B8",X"FF",X"A9",X"00",X"DB",X"00",X"B5",X"FF",X"1E",X"00",X"D8",X"FF",X"0F",X"00",
		X"E2",X"FF",X"0C",X"00",X"E2",X"FF",X"0F",X"00",X"D5",X"FF",X"4B",X"00",X"22",X"01",X"E3",X"FF",
		X"00",X"00",X"F4",X"FF",X"F8",X"FF",X"F9",X"FF",X"F0",X"FF",X"00",X"00",X"E8",X"FF",X"0F",X"00",
		X"C9",X"FF",X"C4",X"00",X"A1",X"00",X"B9",X"FF",X"20",X"00",X"D8",X"FF",X"11",X"00",X"E1",X"FF",
		X"0A",X"00",X"E8",X"FF",X"05",X"00",X"F0",X"FF",X"F6",X"FF",X"77",X"01",X"50",X"00",X"CA",X"FF",
		X"1A",X"00",X"D8",X"FF",X"15",X"00",X"DB",X"FF",X"14",X"00",X"DD",X"FF",X"11",X"00",X"DB",X"FF",
		X"1A",X"00",X"68",X"01",X"21",X"00",X"DA",X"FF",X"12",X"00",X"DC",X"FF",X"13",X"00",X"DD",X"FF",
		X"14",X"00",X"DA",X"FF",X"18",X"00",X"D3",X"FF",X"30",X"00",X"6B",X"01",X"0E",X"00",X"E4",X"FF",
		X"0B",X"00",X"E1",X"FF",X"10",X"00",X"DF",X"FF",X"14",X"00",X"DB",X"FF",X"1A",X"00",X"CF",X"FF",
		X"3F",X"00",X"84",X"01",X"02",X"00",X"EB",X"FF",X"06",X"00",X"E6",X"FF",X"0B",X"00",X"E3",X"FF",
		X"0F",X"00",X"DF",X"FF",X"14",X"00",X"D2",X"FF",X"3D",X"00",X"58",X"01",X"04",X"00",X"EC",X"FF",
		X"08",X"00",X"E7",X"FF",X"0D",X"00",X"E1",X"FF",X"12",X"00",X"D8",X"FF",X"20",X"00",X"BF",X"FF",
		X"74",X"00",X"43",X"01",X"D1",X"FF",X"08",X"00",X"F2",X"FF",X"F7",X"FF",X"FD",X"FF",X"EF",X"FF",
		X"06",X"00",X"E2",X"FF",X"1A",X"00",X"BB",X"FF",X"58",X"01",X"94",X"00",X"BE",X"FF",X"1F",X"00",
		X"DA",X"FF",X"12",X"00",X"E0",X"FF",X"11",X"00",X"DE",X"FF",X"1B",X"00",X"C6",X"FF",X"70",X"00",
		X"07",X"01",X"C1",X"FF",X"1A",X"00",X"E0",X"FF",X"0C",X"00",X"E8",X"FF",X"09",X"00",X"E8",X"FF",
		X"0C",X"00",X"E1",X"FF",X"32",X"00",X"29",X"01",X"F3",X"FF",X"FC",X"FF",X"F8",X"FF",X"F8",X"FF",
		X"FC",X"FF",X"F4",X"FF",X"00",X"00",X"F0",X"FF",X"08",X"00",X"D9",X"FF",X"E7",X"00",X"35",X"00",
		X"DB",X"FF",X"10",X"00",X"E5",X"FF",X"0B",X"00",X"E6",X"FF",X"0F",X"00",X"E2",X"FF",X"1A",X"00",
		X"C7",X"FF",X"9C",X"00",X"B6",X"00",X"C8",X"FF",X"15",X"00",X"E6",X"FF",X"08",X"00",X"F0",X"FF",
		X"00",X"00",X"F6",X"FF",X"FB",X"FF",X"00",X"00",X"E3",X"FF",X"FD",X"00",X"42",X"00",X"D2",X"FF",
		X"18",X"00",X"DE",X"FF",X"15",X"00",X"DE",X"FF",X"18",X"00",X"D8",X"FF",X"26",X"00",X"BC",X"FF",
		X"8F",X"00",X"1E",X"01",X"C4",X"FF",X"16",X"00",X"E7",X"FF",X"05",X"00",X"F3",X"FF",X"FF",X"FF",
		X"F9",X"FF",X"F9",X"FF",X"01",X"00",X"E7",X"FF",X"EC",X"00",X"23",X"00",X"E4",X"FF",X"0A",X"00",
		X"EB",X"FF",X"08",X"00",X"ED",X"FF",X"0D",X"00",X"E7",X"FF",X"18",X"00",X"CC",X"FF",X"D6",X"00",
		X"93",X"00",X"C8",X"FF",X"1B",X"00",X"E2",X"FF",X"0F",X"00",X"E7",X"FF",X"0B",X"00",X"EA",X"FF",
		X"0E",X"00",X"E4",X"FF",X"24",X"00",X"F2",X"00",X"08",X"00",X"EF",X"FF",X"08",X"00",X"EB",X"FF",
		X"0D",X"00",X"E8",X"FF",X"11",X"00",X"DE",X"FF",X"22",X"00",X"BE",X"FF",X"A4",X"00",X"02",X"01",
		X"BE",X"FF",X"1E",X"00",X"E4",X"FF",X"0C",X"00",X"F0",X"FF",X"03",X"00",X"F8",X"FF",X"FC",X"FF",
		X"02",X"00",X"E7",X"FF",X"50",X"01",X"51",X"00",X"D4",X"FF",X"19",X"00",X"E1",X"FF",X"15",X"00",
		X"E1",X"FF",X"18",X"00",X"DC",X"FF",X"25",X"00",X"BD",X"FF",X"A7",X"00",X"D4",X"00",X"C0",X"FF",
		X"1E",X"00",X"E1",X"FF",X"10",X"00",X"EB",X"FF",X"09",X"00",X"EF",X"FF",X"06",X"00",X"F2",X"FF",
		X"04",X"00",X"D7",X"00",X"0F",X"00",X"EA",X"FF",X"0E",X"00",X"EA",X"FF",X"0E",X"00",X"E6",X"FF",
		X"15",X"00",X"DD",X"FF",X"25",X"00",X"BB",X"FF",X"B5",X"00",X"D2",X"00",X"C3",X"FF",X"1C",X"00",
		X"E7",X"FF",X"0A",X"00",X"F3",X"FF",X"03",X"00",X"FA",X"FF",X"FB",X"FF",X"05",X"00",X"E7",X"FF",
		X"F5",X"00",X"5A",X"00",X"D7",X"FF",X"17",X"00",X"E6",X"FF",X"0F",X"00",X"EA",X"FF",X"0F",X"00",
		X"EB",X"FF",X"13",X"00",X"DE",X"FF",X"4D",X"00",X"D9",X"00",X"E2",X"FF",X"08",X"00",X"F4",X"FF",
		X"02",X"00",X"F8",X"FF",X"00",X"00",X"FC",X"FF",X"FC",X"FF",X"00",X"00",X"F7",X"FF",X"30",X"01",
		X"2A",X"00",X"EA",X"FF",X"0B",X"00",X"F0",X"FF",X"09",X"00",X"EE",X"FF",X"0C",X"00",X"EA",X"FF",
		X"16",X"00",X"D0",X"FF",X"91",X"00",X"78",X"00",X"CD",X"FF",X"1C",X"00",X"E4",X"FF",X"14",X"00",
		X"E6",X"FF",X"15",X"00",X"E0",X"FF",X"23",X"00",X"BF",X"FF",X"BD",X"00",X"B9",X"00",X"BC",X"FF",
		X"26",X"00",X"DE",X"FF",X"19",X"00",X"E4",X"FF",X"18",X"00",X"E0",X"FF",X"22",X"00",X"C6",X"FF",
		X"96",X"00",X"E6",X"00",X"CD",X"FF",X"1A",X"00",X"E7",X"FF",X"0C",X"00",X"EF",X"FF",X"0A",X"00",
		X"F4",X"FF",X"08",X"00",X"F5",X"FF",X"07",X"00",X"3F",X"01",X"1B",X"00",X"EB",X"FF",X"0D",X"00",
		X"EB",X"FF",X"11",X"00",X"EA",X"FF",X"17",X"00",X"E2",X"FF",X"22",X"00",X"C5",X"FF",X"9C",X"00",
		X"D8",X"00",X"D4",X"FF",X"10",X"00",X"F5",X"FF",X"00",X"00",X"01",X"00",X"F6",X"FF",X"0B",X"00",
		X"EC",X"FF",X"1B",X"00",X"C7",X"FF",X"C2",X"00",X"8C",X"00",X"CD",X"FF",X"1C",X"00",X"E9",X"FF",
		X"0A",X"00",X"F6",X"FF",X"03",X"00",X"FD",X"FF",X"F7",X"FF",X"0F",X"00",X"D9",X"FF",X"AA",X"00",
		X"69",X"00",X"D0",X"FF",X"1D",X"00",X"E6",X"FF",X"11",X"00",X"EF",X"FF",X"0C",X"00",X"F3",X"FF",
		X"08",X"00",X"F9",X"FF",X"03",X"00",X"D5",X"00",X"32",X"00",X"E2",X"FF",X"13",X"00",X"ED",X"FF",
		X"10",X"00",X"EE",X"FF",X"11",X"00",X"ED",X"FF",X"15",X"00",X"E3",X"FF",X"38",X"00",X"A8",X"00",
		X"E4",X"FF",X"0C",X"00",X"F6",X"FF",X"04",X"00",X"FC",X"FF",X"01",X"00",X"FE",X"FF",X"02",X"00",
		X"FD",X"FF",X"07",X"00",X"E0",X"00",X"18",X"00",X"F3",X"FF",X"08",X"00",X"F5",X"FF",X"08",X"00",
		X"F5",X"FF",X"0C",X"00",X"EE",X"FF",X"19",X"00",X"D2",X"FF",X"DB",X"00",X"5F",X"00",X"D4",X"FF",
		X"1C",X"00",X"E6",X"FF",X"14",X"00",X"E9",X"FF",X"18",X"00",X"E5",X"FF",X"24",X"00",X"C7",X"FF",
		X"D8",X"00",X"95",X"00",X"CE",X"FF",X"1D",X"00",X"E7",X"FF",X"15",X"00",X"ED",X"FF",X"12",X"00",
		X"EA",X"FF",X"1C",X"00",X"D5",X"FF",X"8D",X"00",X"9D",X"00",X"D8",X"FF",X"18",X"00",X"EE",X"FF",
		X"0E",X"00",X"F2",X"FF",X"10",X"00",X"EF",X"FF",X"15",X"00",X"DE",X"FF",X"6A",X"00",X"A2",X"00",
		X"DA",X"FF",X"16",X"00",X"EF",X"FF",X"0F",X"00",X"F0",X"FF",X"0F",X"00",X"EF",X"FF",X"15",X"00",
		X"DF",X"FF",X"68",X"00",X"A2",X"00",X"DC",X"FF",X"17",X"00",X"EF",X"FF",X"10",X"00",X"F2",X"FF",
		X"10",X"00",X"EE",X"FF",X"18",X"00",X"DA",X"FF",X"7B",X"00",X"AA",X"00",X"D7",X"FF",X"1A",X"00",
		X"EC",X"FF",X"13",X"00",X"EE",X"FF",X"14",X"00",X"E9",X"FF",X"1E",X"00",X"D0",X"FF",X"9B",X"00",
		X"B5",X"00",X"CD",X"FF",X"21",X"00",X"E4",X"FF",X"18",X"00",X"E8",X"FF",X"1A",X"00",X"E1",X"FF",
		X"28",X"00",X"C0",X"FF",X"C5",X"00",X"C1",X"00",X"C0",X"FF",X"28",X"00",X"E1",X"FF",X"1A",X"00",
		X"E6",X"FF",X"1A",X"00",X"E4",X"FF",X"25",X"00",X"C7",X"FF",X"A6",X"00",X"9C",X"00",X"CA",X"FF",
		X"21",X"00",X"E6",X"FF",X"17",X"00",X"EB",X"FF",X"16",X"00",X"E6",X"FF",X"1F",X"00",X"CD",X"FF",
		X"91",X"00",X"99",X"00",X"CD",X"FF",X"1F",X"00",X"E7",X"FF",X"13",X"00",X"EE",X"FF",X"12",X"00",
		X"ED",X"FF",X"18",X"00",X"DF",X"FF",X"56",X"00",X"B9",X"00",X"E7",X"FF",X"0E",X"00",X"F9",X"FF",
		X"04",X"00",X"FE",X"FF",X"02",X"00",X"02",X"00",X"FB",X"FF",X"09",X"00",X"EE",X"FF",X"C2",X"00",
		X"44",X"00",X"E3",X"FF",X"15",X"00",X"EF",X"FF",X"10",X"00",X"F0",X"FF",X"12",X"00",X"EB",X"FF",
		X"1B",X"00",X"DA",X"FF",X"6F",X"00",X"B7",X"00",X"DC",X"FF",X"15",X"00",X"F1",X"FF",X"0B",X"00",
		X"F6",X"FF",X"07",X"00",X"FA",X"FF",X"07",X"00",X"FC",X"FF",X"08",X"00",X"EC",X"00",X"03",X"00",
		X"FD",X"FF",X"04",X"00",X"FC",X"FF",X"06",X"00",X"FB",X"FF",X"07",X"00",X"F9",X"FF",X"0B",X"00",
		X"EF",X"FF",X"CD",X"00",X"30",X"00",X"EE",X"FF",X"0E",X"00",X"F7",X"FF",X"0A",X"00",X"F7",X"FF",
		X"0C",X"00",X"F5",X"FF",X"13",X"00",X"E6",X"FF",X"6B",X"00",X"56",X"00",X"E1",X"FF",X"15",X"00",
		X"F2",X"FF",X"10",X"00",X"F4",X"FF",X"0E",X"00",X"F1",X"FF",X"16",X"00",X"DF",X"FF",X"63",X"00",
		X"72",X"00",X"DA",X"FF",X"1A",X"00",X"EC",X"FF",X"14",X"00",X"ED",X"FF",X"16",X"00",X"E9",X"FF",
		X"23",X"00",X"D1",X"FF",X"85",X"00",X"C3",X"00",X"D4",X"FF",X"1A",X"00",X"F0",X"FF",X"0E",X"00",
		X"F6",X"FF",X"08",X"00",X"FE",X"FF",X"04",X"00",X"03",X"00",X"F8",X"FF",X"E9",X"00",X"2F",X"00",
		X"EA",X"FF",X"11",X"00",X"F3",X"FF",X"0F",X"00",X"F6",X"FF",X"10",X"00",X"F2",X"FF",X"16",X"00",
		X"E5",X"FF",X"4C",X"00",X"A1",X"00",X"EB",X"FF",X"0F",X"00",X"FB",X"FF",X"07",X"00",X"FE",X"FF",
		X"06",X"00",X"FF",X"FF",X"03",X"00",X"02",X"00",X"FF",X"FF",X"EE",X"00",X"1C",X"00",X"F6",X"FF",
		X"0C",X"00",X"F9",X"FF",X"0B",X"00",X"F7",X"FF",X"0D",X"00",X"F3",X"FF",X"18",X"00",X"E1",X"FF",
		X"6E",X"00",X"6E",X"00",X"DA",X"FF",X"1C",X"00",X"EE",X"FF",X"16",X"00",X"EF",X"FF",X"17",X"00",
		X"E9",X"FF",X"22",X"00",X"CD",X"FF",X"9D",X"00",X"AB",X"00",X"C8",X"FF",X"27",X"00",X"E6",X"FF",
		X"1A",X"00",X"EB",X"FF",X"1A",X"00",X"E8",X"FF",X"22",X"00",X"D3",X"FF",X"7F",X"00",X"A8",X"00",
		X"D6",X"FF",X"1C",X"00",X"EE",X"FF",X"12",X"00",X"F2",X"FF",X"12",X"00",X"F1",X"FF",X"19",X"00",
		X"E1",X"FF",X"5E",X"00",X"A4",X"00",X"DD",X"FF",X"1A",X"00",X"F0",X"FF",X"12",X"00",X"F4",X"FF",
		X"12",X"00",X"F2",X"FF",X"19",X"00",X"E2",X"FF",X"5A",X"00",X"A8",X"00",X"DD",X"FF",X"19",X"00",
		X"F0",X"FF",X"11",X"00",X"F4",X"FF",X"13",X"00",X"F2",X"FF",X"19",X"00",X"E2",X"FF",X"53",X"00",
		X"A6",X"00",X"E4",X"FF",X"13",X"00",X"F9",X"FF",X"0A",X"00",X"FE",X"FF",X"06",X"00",X"01",X"00",
		X"03",X"00",X"06",X"00",X"F8",X"FF",X"AA",X"00",X"1C",X"00",X"F3",X"FF",X"10",X"00",X"F7",X"FF",
		X"0E",X"00",X"F6",X"FF",X"10",X"00",X"F3",X"FF",X"1A",X"00",X"DE",X"FF",X"64",X"00",X"8A",X"00",
		X"DC",X"FF",X"1A",X"00",X"F3",X"FF",X"0F",X"00",X"FA",X"FF",X"09",X"00",X"FF",X"FF",X"05",X"00",
		X"05",X"00",X"F9",X"FF",X"C9",X"00",X"32",X"00",X"ED",X"FF",X"14",X"00",X"F5",X"FF",X"10",X"00",
		X"F8",X"FF",X"0E",X"00",X"F8",X"FF",X"0D",X"00",X"FA",X"FF",X"0A",X"00",X"D9",X"00",X"0F",X"00",
		X"F9",X"FF",X"0E",X"00",X"F9",X"FF",X"0D",X"00",X"F9",X"FF",X"0D",X"00",X"F9",X"FF",X"0E",X"00",
		X"F7",X"FF",X"15",X"00",X"9C",X"00",X"06",X"00",X"FB",X"FF",X"0D",X"00",X"F7",X"FF",X"10",X"00",
		X"F5",X"FF",X"16",X"00",X"EE",X"FF",X"23",X"00",X"D3",X"FF",X"A5",X"00",X"81",X"00",X"D6",X"FF",
		X"1E",X"00",X"EF",X"FF",X"15",X"00",X"F5",X"FF",X"11",X"00",X"F8",X"FF",X"11",X"00",X"F6",X"FF",
		X"19",X"00",X"B9",X"00",X"FE",X"FF",X"05",X"00",X"06",X"00",X"FF",X"FF",X"0A",X"00",X"FC",X"FF",
		X"0F",X"00",X"F4",X"FF",X"1A",X"00",X"D9",X"FF",X"9F",X"00",X"77",X"00",X"D7",X"FF",X"22",X"00",
		X"EC",X"FF",X"17",X"00",X"F4",X"FF",X"12",X"00",X"F7",X"FF",X"0E",X"00",X"FB",X"FF",X"0B",X"00",
		X"7A",X"00",X"2D",X"00",X"ED",X"FF",X"19",X"00",X"F2",X"FF",X"17",X"00",X"F1",X"FF",X"17",X"00",
		X"F0",X"FF",X"1B",X"00",X"E8",X"FF",X"33",X"00",X"C2",X"00",X"00",X"00",X"01",X"00",X"0B",X"00",
		X"FB",X"FF",X"10",X"00",X"F5",X"FF",X"13",X"00",X"F1",X"FF",X"1B",X"00",X"E4",X"FF",X"41",X"00",
		X"C4",X"00",X"F0",X"FF",X"0B",X"00",X"04",X"00",X"00",X"00",X"0B",X"00",X"FC",X"FF",X"0D",X"00",
		X"F8",X"FF",X"14",X"00",X"EF",X"FF",X"33",X"00",X"9E",X"00",X"FC",X"FF",X"07",X"00",X"05",X"00",
		X"02",X"00",X"08",X"00",X"FD",X"FF",X"0C",X"00",X"FE",X"FF",X"0E",X"00",X"FA",X"FF",X"1B",X"00",
		X"79",X"00",X"0B",X"00",X"FF",X"FF",X"0B",X"00",X"FE",X"FF",X"0D",X"00",X"FD",X"FF",X"0C",X"00",
		X"FF",X"FF",X"0B",X"00",X"FF",X"FF",X"07",X"00",X"6B",X"00",X"18",X"00",X"F7",X"FF",X"11",X"00",
		X"F8",X"FF",X"11",X"00",X"F9",X"FF",X"0F",X"00",X"FB",X"FF",X"0F",X"00",X"FB",X"FF",X"0F",X"00",
		X"8D",X"00",X"12",X"00",X"F8",X"FF",X"11",X"00",X"F9",X"FF",X"11",X"00",X"F9",X"FF",X"10",X"00",
		X"F7",X"FF",X"13",X"00",X"F8",X"FF",X"19",X"00",X"B0",X"00",X"09",X"00",X"FE",X"FF",X"0D",X"00",
		X"FC",X"FF",X"10",X"00",X"FA",X"FF",X"10",X"00",X"F8",X"FF",X"15",X"00",X"F5",X"FF",X"21",X"00",
		X"AA",X"00",X"FF",X"FF",X"04",X"00",X"09",X"00",X"00",X"00",X"0D",X"00",X"FD",X"FF",X"12",X"00",
		X"F7",X"FF",X"1B",X"00",X"E3",X"FF",X"82",X"00",X"5A",X"00",X"E6",X"FF",X"19",X"00",X"F7",X"FF",
		X"11",X"00",X"FC",X"FF",X"0F",X"00",X"FD",X"FF",X"0E",X"00",X"FC",X"FF",X"16",X"00",X"83",X"00",
		X"0B",X"00",X"02",X"00",X"0B",X"00",X"01",X"00",X"0D",X"00",X"FF",X"FF",X"0E",X"00",X"FC",X"FF",
		X"11",X"00",X"F5",X"FF",X"26",X"00",X"81",X"00",X"F5",X"FF",X"0C",X"00",X"04",X"00",X"05",X"00",
		X"07",X"00",X"03",X"00",X"0C",X"00",X"FE",X"FF",X"11",X"00",X"F4",X"FF",X"42",X"00",X"4D",X"00",
		X"F6",X"FF",X"0F",X"00",X"02",X"00",X"08",X"00",X"05",X"00",X"04",X"00",X"0A",X"00",X"00",X"00",
		X"10",X"00",X"F2",X"FF",X"5F",X"00",X"44",X"00",X"F4",X"FF",X"11",X"00",X"00",X"00",X"0B",X"00",
		X"03",X"00",X"08",X"00",X"08",X"00",X"05",X"00",X"0E",X"00",X"FA",X"FF",X"3A",X"00",X"47",X"00",
		X"F4",X"FF",X"11",X"00",X"FF",X"FF",X"0C",X"00",X"03",X"00",X"0A",X"00",X"08",X"00",X"05",X"00",
		X"0C",X"00",X"FB",X"FF",X"88",X"00",X"25",X"00",X"F9",X"FF",X"10",X"00",X"FF",X"FF",X"0D",X"00",
		X"00",X"00",X"0C",X"00",X"02",X"00",X"0B",X"00",X"02",X"00",X"0C",X"00",X"47",X"00",X"0D",X"00",
		X"02",X"00",X"0C",X"00",X"02",X"00",X"0C",X"00",X"02",X"00",X"0C",X"00",X"02",X"00",X"10",X"00",
		X"F9",X"FF",X"3C",X"00",X"31",X"00",X"FA",X"FF",X"10",X"00",X"00",X"00",X"0C",X"00",X"04",X"00",
		X"0B",X"00",X"05",X"00",X"0A",X"00",X"05",X"00",X"07",X"00",X"89",X"00",X"13",X"00",X"FF",X"FF",
		X"11",X"00",X"00",X"00",X"11",X"00",X"FF",X"FF",X"12",X"00",X"FC",X"FF",X"15",X"00",X"F5",X"FF",
		X"36",X"00",X"4E",X"00",X"00",X"00",X"0B",X"00",X"09",X"00",X"04",X"00",X"0B",X"00",X"03",X"00",
		X"10",X"00",X"FE",X"FF",X"16",X"00",X"F1",X"FF",X"4D",X"00",X"44",X"00",X"F6",X"FF",X"12",X"00",
		X"02",X"00",X"0E",X"00",X"04",X"00",X"0C",X"00",X"04",X"00",X"0A",X"00",X"06",X"00",X"0B",X"00",
		X"43",X"00",X"05",X"00",X"09",X"00",X"06",X"00",X"0B",X"00",X"06",X"00",X"0A",X"00",X"05",X"00",
		X"0A",X"00",X"04",X"00",X"0F",X"00",X"D3",X"00",X"06",X"00",X"08",X"00",X"08",X"00",X"08",X"00",
		X"0A",X"00",X"06",X"00",X"0A",X"00",X"05",X"00",X"0B",X"00",X"05",X"00",X"3D",X"00",X"17",X"00",
		X"02",X"00",X"0C",X"00",X"05",X"00",X"0C",X"00",X"04",X"00",X"0E",X"00",X"03",X"00",X"13",X"00",
		X"F6",X"FF",X"44",X"00",X"45",X"00",X"F2",X"FF",X"17",X"00",X"FE",X"FF",X"13",X"00",X"00",X"00",
		X"13",X"00",X"FF",X"FF",X"15",X"00",X"F9",X"FF",X"2E",X"00",X"3C",X"00",X"FF",X"FF",X"0E",X"00",
		X"07",X"00",X"09",X"00",X"0A",X"00",X"08",X"00",X"0A",X"00",X"04",X"00",X"10",X"00",X"FD",X"FF",
		X"34",X"00",X"32",X"00",X"F8",X"FF",X"13",X"00",X"01",X"00",X"0F",X"00",X"03",X"00",X"0E",X"00",
		X"03",X"00",X"0E",X"00",X"02",X"00",X"12",X"00",X"68",X"00",X"06",X"00",X"08",X"00",X"0A",X"00",
		X"08",X"00",X"0B",X"00",X"07",X"00",X"0B",X"00",X"06",X"00",X"0E",X"00",X"05",X"00",X"25",X"00",
		X"1B",X"00",X"FF",X"FF",X"11",X"00",X"04",X"00",X"11",X"00",X"01",X"00",X"15",X"00",X"FA",X"FF",
		X"20",X"00",X"E3",X"FF",X"90",X"00",X"80",X"00",X"DC",X"FF",X"25",X"00",X"F4",X"FF",X"1D",X"00",
		X"FA",X"FF",X"18",X"00",X"FC",X"FF",X"19",X"00",X"FA",X"FF",X"1F",X"00",X"B5",X"00",X"07",X"00",
		X"05",X"00",X"0D",X"00",X"04",X"00",X"0E",X"00",X"04",X"00",X"10",X"00",X"03",X"00",X"11",X"00",
		X"02",X"00",X"17",X"00",X"46",X"00",X"08",X"00",X"0A",X"00",X"0E",X"00",X"08",X"00",X"10",X"00",
		X"05",X"00",X"12",X"00",X"01",X"00",X"15",X"00",X"F7",X"FF",X"47",X"00",X"2C",X"00",X"00",X"00",
		X"0F",X"00",X"07",X"00",X"0B",X"00",X"0A",X"00",X"08",X"00",X"0E",X"00",X"05",X"00",X"13",X"00",
		X"F8",X"FF",X"57",X"00",X"2E",X"00",X"FB",X"FF",X"12",X"00",X"05",X"00",X"0F",X"00",X"07",X"00",
		X"0C",X"00",X"09",X"00",X"08",X"00",X"0E",X"00",X"04",X"00",X"2A",X"00",X"27",X"00",X"01",X"00",
		X"0E",X"00",X"06",X"00",X"0A",X"00",X"0A",X"00",X"09",X"00",X"0B",X"00",X"06",X"00",X"0F",X"00",
		X"01",X"00",X"23",X"00",X"37",X"00",X"01",X"00",X"0E",X"00",X"08",X"00",X"0A",X"00",X"0C",X"00",
		X"08",X"00",X"0F",X"00",X"03",X"00",X"16",X"00",X"FA",X"FF",X"39",X"00",X"4D",X"00",X"FA",X"FF",
		X"13",X"00",X"08",X"00",X"0C",X"00",X"0D",X"00",X"08",X"00",X"11",X"00",X"01",X"00",X"1A",X"00",
		X"F1",X"FF",X"54",X"00",X"5E",X"00",X"F2",X"FF",X"16",X"00",X"06",X"00",X"0E",X"00",X"0C",X"00",
		X"09",X"00",X"11",X"00",X"02",X"00",X"1D",X"00",X"EB",X"FF",X"74",X"00",X"6C",X"00",X"ED",X"FF",
		X"1E",X"00",X"00",X"00",X"11",X"00",X"09",X"00",X"0A",X"00",X"10",X"00",X"00",X"00",X"1C",X"00",
		X"EA",X"FF",X"86",X"00",X"6A",X"00",X"E6",X"FF",X"20",X"00",X"FC",X"FF",X"16",X"00",X"04",X"00",
		X"10",X"00",X"09",X"00",X"0B",X"00",X"10",X"00",X"FC",X"FF",X"51",X"00",X"3B",X"00",X"F8",X"FF",
		X"16",X"00",X"02",X"00",X"11",X"00",X"06",X"00",X"0D",X"00",X"0C",X"00",X"08",X"00",X"11",X"00",
		X"FB",X"FF",X"55",X"00",X"32",X"00",X"FA",X"FF",X"15",X"00",X"04",X"00",X"10",X"00",X"07",X"00",
		X"0D",X"00",X"0A",X"00",X"0A",X"00",X"0D",X"00",X"03",X"00",X"41",X"00",X"23",X"00",X"01",X"00",
		X"13",X"00",X"07",X"00",X"0F",X"00",X"07",X"00",X"0E",X"00",X"08",X"00",X"0D",X"00",X"06",X"00",
		X"17",X"00",X"30",X"00",X"02",X"00",X"12",X"00",X"06",X"00",X"11",X"00",X"04",X"00",X"13",X"00",
		X"01",X"00",X"16",X"00",X"F9",X"FF",X"32",X"00",X"89",X"00",X"F5",X"FF",X"16",X"00",X"05",X"00",
		X"11",X"00",X"08",X"00",X"0E",X"00",X"0A",X"00",X"0B",X"00",X"0C",X"00",X"07",X"00",X"20",X"00",
		X"15",X"00",X"06",X"00",X"0F",X"00",X"09",X"00",X"0E",X"00",X"07",X"00",X"0F",X"00",X"06",X"00",
		X"13",X"00",X"FE",X"FF",X"4F",X"00",X"28",X"00",X"FE",X"FF",X"15",X"00",X"03",X"00",X"14",X"00",
		X"04",X"00",X"13",X"00",X"01",X"00",X"19",X"00",X"F7",X"FF",X"63",X"00",X"32",X"00",X"FA",X"FF",
		X"18",X"00",X"00",X"00",X"14",X"00",X"02",X"00",X"17",X"00",X"FF",X"FF",X"1F",X"00",X"EB",X"FF",
		X"8E",X"00",X"4D",X"00",X"EF",X"FF",X"1D",X"00",X"FC",X"FF",X"18",X"00",X"FF",X"FF",X"15",X"00",
		X"FF",X"FF",X"15",X"00",X"FD",X"FF",X"24",X"00",X"5D",X"00",X"04",X"00",X"0D",X"00",X"0B",X"00",
		X"0A",X"00",X"0E",X"00",X"07",X"00",X"11",X"00",X"03",X"00",X"18",X"00",X"F5",X"FF",X"7D",X"00",
		X"3E",X"00",X"F4",X"FF",X"1B",X"00",X"FD",X"FF",X"16",X"00",X"00",X"00",X"16",X"00",X"FF",X"FF",
		X"19",X"00",X"F9",X"FF",X"2F",X"00",X"79",X"00",X"FA",X"FF",X"12",X"00",X"06",X"00",X"0E",X"00",
		X"0B",X"00",X"0B",X"00",X"0C",X"00",X"0A",X"00",X"0D",X"00",X"07",X"00",X"1C",X"00",X"13",X"00",
		X"06",X"00",X"0E",X"00",X"08",X"00",X"0F",X"00",X"08",X"00",X"11",X"00",X"06",X"00",X"14",X"00",
		X"FF",X"FF",X"4F",X"00",X"2A",X"00",X"00",X"00",X"14",X"00",X"05",X"00",X"13",X"00",X"08",X"00",
		X"11",X"00",X"07",X"00",X"0F",X"00",X"07",X"00",X"10",X"00",X"08",X"00",X"0F",X"00",X"08",X"00",
		X"10",X"00",X"07",X"00",X"11",X"00",X"07",X"00",X"12",X"00",X"05",X"00",X"15",X"00",X"FE",X"FF",
		X"2A",X"00",X"51",X"00",X"FF",X"FF",X"13",X"00",X"08",X"00",X"0E",X"00",X"0B",X"00",X"0B",X"00",
		X"0C",X"00",X"08",X"00",X"11",X"00",X"00",X"00",X"5B",X"00",X"22",X"00",X"02",X"00",X"13",X"00",
		X"05",X"00",X"11",X"00",X"08",X"00",X"0F",X"00",X"09",X"00",X"0E",X"00",X"0A",X"00",X"0E",X"00",
		X"0A",X"00",X"0E",X"00",X"0B",X"00",X"0E",X"00",X"0A",X"00",X"0D",X"00",X"0B",X"00",X"0C",X"00",
		X"0A",X"00",X"0E",X"00",X"0B",X"00",X"0C",X"00",X"0A",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",
		X"0D",X"00",X"0B",X"00",X"0F",X"00",X"0C",X"00",X"10",X"00",X"06",X"00",X"23",X"00",X"38",X"00",
		X"FF",X"FF",X"14",X"00",X"07",X"00",X"11",X"00",X"08",X"00",X"10",X"00",X"09",X"00",X"10",X"00",
		X"0B",X"00",X"0D",X"00",X"22",X"00",X"13",X"00",X"09",X"00",X"12",X"00",X"0B",X"00",X"10",X"00",
		X"0A",X"00",X"0F",X"00",X"0C",X"00",X"0E",X"00",X"0E",X"00",X"0A",X"00",X"5D",X"00",X"19",X"00",
		X"05",X"00",X"12",X"00",X"08",X"00",X"12",X"00",X"0A",X"00",X"12",X"00",X"08",X"00",X"11",X"00",
		X"0B",X"00",X"0F",X"00",X"67",X"00",X"13",X"00",X"09",X"00",X"12",X"00",X"09",X"00",X"10",X"00",
		X"0A",X"00",X"11",X"00",X"0A",X"00",X"11",X"00",X"09",X"00",X"11",X"00",X"2F",X"00",X"10",X"00",
		X"0A",X"00",X"10",X"00",X"0B",X"00",X"0F",X"00",X"0B",X"00",X"11",X"00",X"08",X"00",X"12",X"00",
		X"06",X"00",X"21",X"00",X"1D",X"00",X"08",X"00",X"10",X"00",X"0B",X"00",X"0E",X"00",X"0C",X"00",
		X"10",X"00",X"0A",X"00",X"12",X"00",X"05",X"00",X"27",X"00",X"27",X"00",X"04",X"00",X"12",X"00",
		X"09",X"00",X"11",X"00",X"0B",X"00",X"0E",X"00",X"0B",X"00",X"0F",X"00",X"0B",X"00",X"0F",X"00",
		X"2B",X"00",X"0D",X"00",X"0C",X"00",X"0D",X"00",X"0C",X"00",X"0D",X"00",X"0C",X"00",X"0D",X"00",
		X"0D",X"00",X"0D",X"00",X"0E",X"00",X"6A",X"00",X"0B",X"00",X"0E",X"00",X"0C",X"00",X"0D",X"00",
		X"0D",X"00",X"0D",X"00",X"0E",X"00",X"0D",X"00",X"0E",X"00",X"0A",X"00",X"84",X"00",X"10",X"00",
		X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0E",X"00",X"0B",X"00",X"0E",X"00",X"0C",X"00",X"0F",X"00",
		X"07",X"00",X"87",X"00",X"12",X"00",X"0A",X"00",X"10",X"00",X"0A",X"00",X"0F",X"00",X"0B",X"00",
		X"0F",X"00",X"0A",X"00",X"10",X"00",X"05",X"00",X"79",X"00",X"15",X"00",X"08",X"00",X"0F",X"00",
		X"0A",X"00",X"0F",X"00",X"0B",X"00",X"10",X"00",X"09",X"00",X"10",X"00",X"07",X"00",X"5D",X"00",
		X"15",X"00",X"0A",X"00",X"10",X"00",X"0A",X"00",X"11",X"00",X"0C",X"00",X"10",X"00",X"0B",X"00",
		X"11",X"00",X"07",X"00",X"3A",X"00",X"12",X"00",X"0B",X"00",X"0F",X"00",X"0D",X"00",X"0E",X"00",
		X"0D",X"00",X"0F",X"00",X"0B",X"00",X"0F",X"00",X"0C",X"00",X"11",X"00",X"0C",X"00",X"0D",X"00",
		X"0D",X"00",X"0E",X"00",X"0D",X"00",X"0E",X"00",X"0D",X"00",X"0E",X"00",X"0C",X"00",X"0D",X"00",
		X"0B",X"00",X"0C",X"00",X"0E",X"00",X"0E",X"00",X"0D",X"00",X"0E",X"00",X"0E",X"00",X"0D",X"00",
		X"0B",X"00",X"0F",X"00",X"0A",X"00",X"20",X"00",X"12",X"00",X"0C",X"00",X"0E",X"00",X"0D",X"00",
		X"0E",X"00",X"0D",X"00",X"0E",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0F",X"00",X"0D",X"00",
		X"0F",X"00",X"0D",X"00",X"0F",X"00",X"0D",X"00",X"0F",X"00",X"0E",X"00",X"0F",X"00",X"0E",X"00",
		X"0F",X"00",X"09",X"00",X"2E",X"00",X"14",X"00",X"09",X"00",X"10",X"00",X"0C",X"00",X"11",X"00",
		X"0B",X"00",X"10",X"00",X"0D",X"00",X"11",X"00",X"0D",X"00",X"11",X"00",X"0C",X"00",X"12",X"00",
		X"0A",X"00",X"11",X"00",X"0A",X"00",X"13",X"00",X"09",X"00",X"13",X"00",X"07",X"00",X"19",X"00",
		X"FE",X"FF",X"37",X"00",X"44",X"00",X"00",X"00",X"15",X"00",X"09",X"00",X"0F",X"00",X"0D",X"00",
		X"0E",X"00",X"10",X"00",X"0C",X"00",X"12",X"00",X"04",X"00",X"29",X"00",X"2E",X"00",X"03",X"00",
		X"14",X"00",X"0A",X"00",X"12",X"00",X"0B",X"00",X"0F",X"00",X"0D",X"00",X"0F",X"00",X"0D",X"00",
		X"0F",X"00",X"0D",X"00",X"0D",X"00",X"0F",X"00",X"0E",X"00",X"0F",X"00",X"0D",X"00",X"10",X"00",
		X"0C",X"00",X"10",X"00",X"0A",X"00",X"14",X"00",X"04",X"00",X"32",X"00",X"28",X"00",X"05",X"00",
		X"14",X"00",X"0A",X"00",X"11",X"00",X"0C",X"00",X"10",X"00",X"0C",X"00",X"10",X"00",X"0D",X"00",
		X"10",X"00",X"0E",X"00",X"0F",X"00",X"0E",X"00",X"0F",X"00",X"0F",X"00",X"0D",X"00",X"0E",X"00",
		X"0F",X"00",X"0E",X"00",X"0E",X"00",X"0D",X"00",X"12",X"00",X"10",X"00",X"0D",X"00",X"10",X"00",
		X"0D",X"00",X"10",X"00",X"0E",X"00",X"10",X"00",X"0E",X"00",X"10",X"00",X"0C",X"00",X"14",X"00",
		X"39",X"00",X"09",X"00",X"11",X"00",X"0C",X"00",X"11",X"00",X"0C",X"00",X"10",X"00",X"0C",X"00",
		X"11",X"00",X"0A",X"00",X"16",X"00",X"51",X"00",X"09",X"00",X"11",X"00",X"0E",X"00",X"0D",X"00",
		X"0E",X"00",X"0E",X"00",X"0F",X"00",X"0C",X"00",X"11",X"00",X"06",X"00",X"30",X"00",X"25",X"00",
		X"03",X"00",X"15",X"00",X"08",X"00",X"13",X"00",X"0B",X"00",X"12",X"00",X"09",X"00",X"12",X"00",
		X"06",X"00",X"1C",X"00",X"5F",X"00",X"06",X"00",X"13",X"00",X"0B",X"00",X"10",X"00",X"0D",X"00",
		X"10",X"00",X"0D",X"00",X"0E",X"00",X"0E",X"00",X"0A",X"00",X"24",X"00",X"1E",X"00",X"06",X"00",
		X"15",X"00",X"08",X"00",X"13",X"00",X"09",X"00",X"14",X"00",X"07",X"00",X"16",X"00",X"03",X"00",
		X"23",X"00",X"70",X"00",X"02",X"00",X"13",X"00",X"0B",X"00",X"0F",X"00",X"0E",X"00",X"0E",X"00",
		X"0D",X"00",X"0E",X"00",X"0F",X"00",X"0C",X"00",X"17",X"00",X"12",X"00",X"0C",X"00",X"0F",X"00",
		X"0E",X"00",X"0F",X"00",X"0E",X"00",X"0F",X"00",X"0E",X"00",X"0F",X"00",X"0D",X"00",X"10",X"00",
		X"0F",X"00",X"0F",X"00",X"0C",X"00",X"0F",X"00",X"0C",X"00",X"10",X"00",X"0B",X"00",X"12",X"00",
		X"07",X"00",X"18",X"00",X"FC",X"FF",X"63",X"00",X"32",X"00",X"FD",X"FF",X"17",X"00",X"05",X"00",
		X"14",X"00",X"09",X"00",X"12",X"00",X"0B",X"00",X"12",X"00",X"0C",X"00",X"0D",X"00",X"1E",X"00",
		X"16",X"00",X"08",X"00",X"13",X"00",X"0A",X"00",X"11",X"00",X"0B",X"00",X"12",X"00",X"0C",X"00",
		X"11",X"00",X"0C",X"00",X"11",X"00",X"0C",X"00",X"11",X"00",X"0C",X"00",X"11",X"00",X"0C",X"00",
		X"11",X"00",X"0C",X"00",X"10",X"00",X"0C",X"00",X"0F",X"00",X"0D",X"00",X"10",X"00",X"0B",X"00",
		X"11",X"00",X"0C",X"00",X"11",X"00",X"0C",X"00",X"10",X"00",X"0A",X"00",X"11",X"00",X"0A",X"00",
		X"11",X"00",X"06",X"00",X"22",X"00",X"29",X"00",X"06",X"00",X"11",X"00",X"0C",X"00",X"10",X"00",
		X"0D",X"00",X"0F",X"00",X"0C",X"00",X"10",X"00",X"0C",X"00",X"0E",X"00",X"0D",X"00",X"10",X"00",
		X"0D",X"00",X"0F",X"00",X"0D",X"00",X"0F",X"00",X"0E",X"00",X"10",X"00",X"0E",X"00",X"0F",X"00",
		X"0D",X"00",X"10",X"00",X"0F",X"00",X"11",X"00",X"0D",X"00",X"10",X"00",X"0D",X"00",X"11",X"00",
		X"0D",X"00",X"10",X"00",X"0D",X"00",X"11",X"00",X"0D",X"00",X"10",X"00",X"0D",X"00",X"12",X"00",
		X"0B",X"00",X"13",X"00",X"09",X"00",X"14",X"00",X"07",X"00",X"19",X"00",X"FE",X"FF",X"3A",X"00",
		X"57",X"00",X"FC",X"FF",X"19",X"00",X"08",X"00",X"15",X"00",X"0A",X"00",X"12",X"00",X"0D",X"00",
		X"10",X"00",X"10",X"00",X"0A",X"00",X"61",X"00",X"1B",X"00",X"06",X"00",X"14",X"00",X"09",X"00",
		X"12",X"00",X"09",X"00",X"12",X"00",X"0A",X"00",X"10",X"00",X"0A",X"00",X"11",X"00",X"0A",X"00",
		X"12",X"00",X"0C",X"00",X"13",X"00",X"0B",X"00",X"14",X"00",X"0A",X"00",X"13",X"00",X"09",X"00",
		X"16",X"00",X"05",X"00",X"28",X"00",X"27",X"00",X"09",X"00",X"12",X"00",X"0E",X"00",X"0E",X"00",
		X"11",X"00",X"0C",X"00",X"14",X"00",X"09",X"00",X"19",X"00",X"01",X"00",X"3F",X"00",X"3A",X"00",
		X"00",X"00",X"17",X"00",X"08",X"00",X"13",X"00",X"0B",X"00",X"10",X"00",X"0C",X"00",X"10",X"00",
		X"0D",X"00",X"0D",X"00",X"17",X"00",X"18",X"00",X"09",X"00",X"10",X"00",X"0C",X"00",X"10",X"00",
		X"0C",X"00",X"0F",X"00",X"0E",X"00",X"10",X"00",X"0E",X"00",X"11",X"00",X"0F",X"00",X"10",X"00",
		X"0D",X"00",X"0E",X"00",X"0E",X"00",X"11",X"00",X"0F",X"00",X"0F",X"00",X"10",X"00",X"0F",X"00",
		X"10",X"00",X"0E",X"00",X"10",X"00",X"0F",X"00",X"0F",X"00",X"0E",X"00",X"0F",X"00",X"0E",X"00",
		X"0F",X"00",X"0F",X"00",X"10",X"00",X"0E",X"00",X"10",X"00",X"0E",X"00",X"10",X"00",X"0D",X"00",
		X"11",X"00",X"0F",X"00",X"0F",X"00",X"0E",X"00",X"0F",X"00",X"0E",X"00",X"10",X"00",X"0D",X"00",
		X"10",X"00",X"0D",X"00",X"11",X"00",X"0C",X"00",X"11",X"00",X"0D",X"00",X"10",X"00",X"0E",X"00",
		X"12",X"00",X"0C",X"00",X"13",X"00",X"09",X"00",X"1C",X"00",X"33",X"00",X"0A",X"00",X"11",X"00",
		X"0E",X"00",X"10",X"00",X"0E",X"00",X"10",X"00",X"0F",X"00",X"0F",X"00",X"0E",X"00",X"10",X"00",
		X"0F",X"00",X"10",X"00",X"0E",X"00",X"10",X"00",X"0E",X"00",X"10",X"00",X"0D",X"00",X"11",X"00",
		X"0C",X"00",X"15",X"00",X"05",X"00",X"43",X"00",X"24",X"00",X"06",X"00",X"16",X"00",X"0A",X"00",
		X"13",X"00",X"0A",X"00",X"14",X"00",X"0C",X"00",X"13",X"00",X"0B",X"00",X"14",X"00",X"17",X"00",
		X"0F",X"00",X"0D",X"00",X"10",X"00",X"0D",X"00",X"10",X"00",X"0E",X"00",X"11",X"00",X"0F",X"00",
		X"0F",X"00",X"0F",X"00",X"10",X"00",X"0E",X"00",X"0F",X"00",X"0D",X"00",X"10",X"00",X"0E",X"00",
		X"10",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"10",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",
		X"0F",X"00",X"0F",X"00",X"0F",X"00",X"10",X"00",X"0E",X"00",X"0F",X"00",X"0D",X"00",X"13",X"00",
		X"08",X"00",X"39",X"00",X"1C",X"00",X"09",X"00",X"14",X"00",X"0C",X"00",X"11",X"00",X"0D",X"00",
		X"11",X"00",X"0D",X"00",X"10",X"00",X"0E",X"00",X"11",X"00",X"0E",X"00",X"10",X"00",X"0E",X"00",
		X"10",X"00",X"0D",X"00",X"10",X"00",X"0F",X"00",X"10",X"00",X"0E",X"00",X"0F",X"00",X"0E",X"00",
		X"0F",X"00",X"0E",X"00",X"10",X"00",X"0E",X"00",X"10",X"00",X"0E",X"00",X"10",X"00",X"0E",X"00",
		X"11",X"00",X"0C",X"00",X"14",X"00",X"1B",X"00",X"0D",X"00",X"10",X"00",X"0E",X"00",X"10",X"00",
		X"0E",X"00",X"10",X"00",X"0F",X"00",X"10",X"00",X"0F",X"00",X"10",X"00",X"0E",X"00",X"0F",X"00",
		X"0D",X"00",X"0F",X"00",X"0F",X"00",X"11",X"00",X"0E",X"00",X"10",X"00",X"0E",X"00",X"12",X"00",
		X"0C",X"00",X"19",X"00",X"25",X"00",X"09",X"00",X"12",X"00",X"0E",X"00",X"10",X"00",X"0F",X"00",
		X"0F",X"00",X"10",X"00",X"0E",X"00",X"11",X"00",X"0D",X"00",X"20",X"00",X"14",X"00",X"0C",X"00",
		X"11",X"00",X"0D",X"00",X"10",X"00",X"0D",X"00",X"10",X"00",X"0F",X"00",X"0F",X"00",X"0E",X"00",
		X"11",X"00",X"0E",X"00",X"0F",X"00",X"10",X"00",X"10",X"00",X"0F",X"00",X"0F",X"00",X"0E",X"00",
		X"10",X"00",X"0E",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"11",X"00",X"0F",X"00",
		X"0F",X"00",X"10",X"00",X"0F",X"00",X"0E",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"10",X"00",
		X"0F",X"00",X"10",X"00",X"0E",X"00",X"0F",X"00",X"0E",X"00",X"0F",X"00",X"0F",X"00",X"10",X"00",
		X"0C",X"00",X"11",X"00",X"0B",X"00",X"35",X"00",X"16",X"00",X"0D",X"00",X"11",X"00",X"0D",X"00",
		X"10",X"00",X"0E",X"00",X"10",X"00",X"0E",X"00",X"11",X"00",X"0F",X"00",X"11",X"00",X"0E",X"00",
		X"0F",X"00",X"0F",X"00",X"11",X"00",X"0F",X"00",X"0F",X"00",X"0E",X"00",X"11",X"00",X"0F",X"00",
		X"10",X"00",X"0E",X"00",X"0F",X"00",X"0D",X"00",X"0F",X"00",X"0F",X"00",X"10",X"00",X"0D",X"00",
		X"0F",X"00",X"0F",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0F",X"00",X"10",X"00",X"0E",X"00",
		X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0E",X"00",X"10",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",
		X"0E",X"00",X"10",X"00",X"0E",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",
		X"0F",X"00",X"10",X"00",X"0F",X"00",X"11",X"00",X"0D",X"00",X"16",X"00",X"17",X"00",X"0D",X"00",
		X"11",X"00",X"0E",X"00",X"10",X"00",X"0F",X"00",X"0F",X"00",X"10",X"00",X"0E",X"00",X"0E",X"00",
		X"10",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",
		X"10",X"00",X"0F",X"00",X"0E",X"00",X"10",X"00",X"10",X"00",X"10",X"00",X"0F",X"00",X"0E",X"00",
		X"0F",X"00",X"0E",X"00",X"0E",X"00",X"10",X"00",X"0E",X"00",X"0F",X"00",X"0E",X"00",X"0E",X"00",
		X"10",X"00",X"0E",X"00",X"0E",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",
		X"10",X"00",X"0F",X"00",X"10",X"00",X"10",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",
		X"10",X"00",X"0F",X"00",X"10",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"10",X"00",X"0F",X"00",
		X"0F",X"00",X"0E",X"00",X"0E",X"00",X"0F",X"00",X"0F",X"00",X"0E",X"00",X"0F",X"00",X"0F",X"00",
		X"0F",X"00",X"10",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0E",X"00",X"0E",X"00",
		X"0F",X"00",X"0E",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",
		X"0E",X"00",X"0F",X"00",X"0D",X"00",X"0E",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"10",X"00",
		X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0E",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",
		X"0F",X"00",X"0E",X"00",X"0F",X"00",X"0F",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0F",X"00",
		X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0E",X"00",X"0E",X"00",X"0F",X"00",X"10",X"00",
		X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0E",X"00",X"0E",X"00",X"10",X"00",X"0F",X"00",X"0E",X"00",
		X"10",X"00",X"0F",X"00",X"10",X"00",X"0E",X"00",X"10",X"00",X"0E",X"00",X"11",X"00",X"0E",X"00",
		X"10",X"00",X"0D",X"00",X"10",X"00",X"0F",X"00",X"10",X"00",X"0D",X"00",X"11",X"00",X"0E",X"00",
		X"11",X"00",X"0A",X"00",X"1E",X"00",X"1E",X"00",X"0A",X"00",X"13",X"00",X"0B",X"00",X"10",X"00",
		X"0D",X"00",X"11",X"00",X"0D",X"00",X"11",X"00",X"0E",X"00",X"10",X"00",X"0E",X"00",X"10",X"00",
		X"0F",X"00",X"0E",X"00",X"0F",X"00",X"10",X"00",X"0E",X"00",X"0F",X"00",X"10",X"00",X"0F",X"00",
		X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"10",X"00",X"0F",X"00",X"0F",X"00",
		X"0F",X"00",X"0E",X"00",X"0F",X"00",X"10",X"00",X"0D",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",
		X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"10",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",
		X"0F",X"00",X"0E",X"00",X"10",X"00",X"0F",X"00",X"0E",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",
		X"10",X"00",X"0E",X"00",X"0F",X"00",X"0E",X"00",X"0F",X"00",X"0E",X"00",X"0F",X"00",X"0E",X"00",
		X"0F",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"10",X"00",X"0E",X"00",X"10",X"00",X"0F",X"00",
		X"10",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0E",X"00",X"0F",X"00",X"0E",X"00",X"0E",X"00",
		X"0F",X"00",X"10",X"00",X"10",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0E",X"00",X"0F",X"00",
		X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"10",X"00",X"0F",X"00",X"0E",X"00",X"0F",X"00",
		X"0F",X"00",X"0E",X"00",X"10",X"00",X"0F",X"00",X"10",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",
		X"0F",X"00",X"0E",X"00",X"0E",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0E",X"00",
		X"10",X"00",X"0E",X"00",X"10",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"11",X"00",X"0B",X"00",
		X"16",X"00",X"19",X"00",X"0C",X"00",X"10",X"00",X"0E",X"00",X"0F",X"00",X"0F",X"00",X"10",X"00",
		X"10",X"00",X"0F",X"00",X"0E",X"00",X"10",X"00",X"0E",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",
		X"0F",X"00",X"0F",X"00",X"0E",X"00",X"0F",X"00",X"0F",X"00",X"10",X"00",X"0E",X"00",X"10",X"00",
		X"0F",X"00",X"0F",X"00",X"10",X"00",X"10",X"00",X"0F",X"00",X"0E",X"00",X"0F",X"00",X"10",X"00",
		X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0D",X"00",X"10",X"00",X"0F",X"00",X"0F",X"00",X"0E",X"00",
		X"0F",X"00",X"10",X"00",X"0E",X"00",X"10",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",
		X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"10",X"00",
		X"0E",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0E",X"00",X"0F",X"00",X"10",X"00",X"10",X"00",
		X"0F",X"00",X"0F",X"00",X"10",X"00",X"0F",X"00",X"10",X"00",X"0F",X"00",X"0F",X"00",X"10",X"00",
		X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0E",X"00",
		X"0F",X"00",X"0F",X"00",X"0E",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0E",X"00",X"0F",X"00",
		X"0E",X"00",X"0E",X"00",X"10",X"00",X"0F",X"00",X"0E",X"00",X"0F",X"00",X"0F",X"00",X"0E",X"00",
		X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0F",X"00",X"10",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",
		X"0F",X"00",X"0F",X"00",X"0E",X"00",X"0E",X"00",X"0F",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",
		X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0D",X"00",X"0F",X"00",X"0E",X"00",X"0D",X"00",X"0D",X"00",
		X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0F",X"00",X"0E",X"00",
		X"0D",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0F",X"00",X"0E",X"00",X"0E",X"00",X"0D",X"00",
		X"0E",X"00",X"0E",X"00",X"0D",X"00",X"0E",X"00",X"0E",X"00",X"0D",X"00",X"0E",X"00",X"0E",X"00",
		X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0D",X"00",X"0D",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",
		X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0D",X"00",X"0D",X"00",
		X"0F",X"00",X"0D",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0F",X"00",X"0E",X"00",
		X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0F",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0D",X"00",
		X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0F",X"00",X"0E",X"00",X"0E",X"00",X"0F",X"00",
		X"0F",X"00",X"0D",X"00",X"0D",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",
		X"0D",X"00",X"0E",X"00",X"0E",X"00",X"0F",X"00",X"0E",X"00",X"0D",X"00",X"0E",X"00",X"0E",X"00",
		X"0F",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0F",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",
		X"0E",X"00",X"0E",X"00",X"0F",X"00",X"0D",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0F",X"00",
		X"0E",X"00",X"0F",X"00",X"0E",X"00",X"0D",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",
		X"0F",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0F",X"00",X"0E",X"00",X"0E",X"00",
		X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0D",X"00",X"0D",X"00",X"0E",X"00",X"0F",X"00",X"0D",X"00",
		X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0E",X"00",X"0E",X"00",
		X"0E",X"00",X"0E",X"00",X"0F",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",
		X"0F",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",
		X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0D",X"00",X"0E",X"00",X"0E",X"00",X"0D",X"00",
		X"0E",X"00",X"10",X"00",X"0D",X"00",X"0E",X"00",X"0E",X"00",X"0D",X"00",X"0E",X"00",X"0E",X"00",
		X"0E",X"00",X"0F",X"00",X"0D",X"00",X"0E",X"00",X"0D",X"00",X"0E",X"00",X"0F",X"00",X"0F",X"00",
		X"0E",X"00",X"0E",X"00",X"0F",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0D",X"00",
		X"0F",X"00",X"0F",X"00",X"0E",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0F",X"00",X"0E",X"00",
		X"0E",X"00",X"0F",X"00",X"0E",X"00",X"0D",X"00",X"0D",X"00",X"0E",X"00",X"0D",X"00",X"0D",X"00",
		X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0F",X"00",X"0D",X"00",X"0E",X"00",X"0D",X"00",
		X"0E",X"00",X"0F",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",
		X"0E",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0D",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",
		X"0E",X"00",X"0E",X"00",X"0F",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0D",X"00",
		X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0F",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0D",X"00",
		X"0E",X"00",X"0C",X"00",X"0D",X"00",X"0E",X"00",X"0E",X"00",X"0D",X"00",X"0E",X"00",X"0D",X"00",
		X"0E",X"00",X"0E",X"00",X"0F",X"00",X"0F",X"00",X"0D",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",
		X"0E",X"00",X"0E",X"00",X"0D",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0F",X"00",X"0F",X"00",
		X"0E",X"00",X"0D",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0D",X"00",X"0E",X"00",
		X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0D",X"00",X"0F",X"00",X"0C",X"00",X"0D",X"00",
		X"0D",X"00",X"0C",X"00",X"0D",X"00",X"0E",X"00",X"0D",X"00",X"0D",X"00",X"0F",X"00",X"0D",X"00",
		X"0E",X"00",X"0D",X"00",X"0E",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",
		X"0E",X"00",X"0C",X"00",X"0C",X"00",X"0E",X"00",X"0C",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",
		X"0E",X"00",X"0C",X"00",X"0E",X"00",X"0D",X"00",X"0E",X"00",X"0D",X"00",X"0E",X"00",X"0D",X"00",
		X"0D",X"00",X"0D",X"00",X"0C",X"00",X"0E",X"00",X"0D",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",
		X"0E",X"00",X"0D",X"00",X"0D",X"00",X"0B",X"00",X"0E",X"00",X"0D",X"00",X"0C",X"00",X"0E",X"00",
		X"0E",X"00",X"0D",X"00",X"0E",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0E",X"00",
		X"0C",X"00",X"0F",X"00",X"0D",X"00",X"0C",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0E",X"00",
		X"0C",X"00",X"0D",X"00",X"0C",X"00",X"0D",X"00",X"0C",X"00",X"0C",X"00",X"0D",X"00",X"0D",X"00",
		X"0B",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0E",X"00",
		X"0D",X"00",X"0D",X"00",X"0C",X"00",X"0D",X"00",X"0E",X"00",X"0D",X"00",X"0D",X"00",X"0C",X"00",
		X"0E",X"00",X"0D",X"00",X"0D",X"00",X"0C",X"00",X"0E",X"00",X"0C",X"00",X"0D",X"00",X"0E",X"00",
		X"0D",X"00",X"0E",X"00",X"0C",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",
		X"0C",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",
		X"0D",X"00",X"0E",X"00",X"0E",X"00",X"0D",X"00",X"0D",X"00",X"0E",X"00",X"0D",X"00",X"0E",X"00",
		X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0C",X"00",X"0E",X"00",X"0E",X"00",X"0D",X"00",X"0D",X"00",
		X"0D",X"00",X"0C",X"00",X"0D",X"00",X"0D",X"00",X"0E",X"00",X"0C",X"00",X"0B",X"00",X"0D",X"00",
		X"0D",X"00",X"0E",X"00",X"0E",X"00",X"0D",X"00",X"0C",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",
		X"0C",X"00",X"0D",X"00",X"0E",X"00",X"0D",X"00",X"0C",X"00",X"0D",X"00",X"0E",X"00",X"0C",X"00",
		X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0E",X"00",X"0C",X"00",X"0D",X"00",X"0C",X"00",X"0E",X"00",
		X"0C",X"00",X"0D",X"00",X"0E",X"00",X"0E",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0E",X"00",
		X"0D",X"00",X"0C",X"00",X"0C",X"00",X"0D",X"00",X"0C",X"00",X"0D",X"00",X"0F",X"00",X"0D",X"00",
		X"0C",X"00",X"0E",X"00",X"0C",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0C",X"00",
		X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0E",X"00",X"0D",X"00",X"0C",X"00",
		X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0E",X"00",X"0D",X"00",X"0C",X"00",X"0C",X"00",
		X"0E",X"00",X"0D",X"00",X"0E",X"00",X"0D",X"00",X"0C",X"00",X"0D",X"00",X"0D",X"00",X"0E",X"00",
		X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",
		X"0C",X"00",X"0D",X"00",X"0D",X"00",X"0B",X"00",X"0D",X"00",X"0C",X"00",X"0C",X"00",X"0D",X"00",
		X"0D",X"00",X"0C",X"00",X"0D",X"00",X"0E",X"00",X"0D",X"00",X"0D",X"00",X"0C",X"00",X"0D",X"00",
		X"0C",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0C",X"00",X"0C",X"00",X"0E",X"00",X"0B",X"00",
		X"0C",X"00",X"0B",X"00",X"0C",X"00",X"0B",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",
		X"0C",X"00",X"0C",X"00",X"0D",X"00",X"0B",X"00",X"0C",X"00",X"0E",X"00",X"0D",X"00",X"0D",X"00",
		X"0C",X"00",X"0B",X"00",X"0C",X"00",X"0D",X"00",X"0C",X"00",X"0D",X"00",X"0D",X"00",X"0C",X"00",
		X"0C",X"00",X"0E",X"00",X"0C",X"00",X"0D",X"00",X"0C",X"00",X"0C",X"00",X"0D",X"00",X"0A",X"00",
		X"0D",X"00",X"0C",X"00",X"0B",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",
		X"0D",X"00",X"0D",X"00",X"0C",X"00",X"0B",X"00",X"0B",X"00",X"0B",X"00",X"0D",X"00",X"0A",X"00",
		X"0C",X"00",X"0B",X"00",X"0C",X"00",X"0D",X"00",X"0D",X"00",X"0C",X"00",X"0C",X"00",X"0D",X"00",
		X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0B",X"00",X"0C",X"00",
		X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0D",X"00",X"0C",X"00",X"0C",X"00",X"0B",X"00",X"0C",X"00",
		X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",
		X"0C",X"00",X"0C",X"00",X"0E",X"00",X"0C",X"00",X"0C",X"00",X"0B",X"00",X"0C",X"00",X"0C",X"00",
		X"0C",X"00",X"0D",X"00",X"0C",X"00",X"0C",X"00",X"0B",X"00",X"0C",X"00",X"0C",X"00",X"0B",X"00",
		X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0B",X"00",X"0B",X"00",X"0C",X"00",X"0C",X"00",
		X"0C",X"00",X"0C",X"00",X"0E",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",
		X"0C",X"00",X"0C",X"00",X"0D",X"00",X"0B",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0B",X"00",
		X"0D",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0B",X"00",X"0C",X"00",X"0D",X"00",
		X"0D",X"00",X"0B",X"00",X"0C",X"00",X"0C",X"00",X"0B",X"00",X"0B",X"00",X"0C",X"00",X"0D",X"00",
		X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0D",X"00",X"0B",X"00",X"0D",X"00",X"0B",X"00",X"0D",X"00",
		X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0A",X"00",X"0D",X"00",X"0D",X"00",X"0C",X"00",X"0B",X"00",
		X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0D",X"00",X"0C",X"00",X"0B",X"00",X"0C",X"00",X"0C",X"00",
		X"0D",X"00",X"0C",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0C",X"00",X"0C",X"00",X"0D",X"00",
		X"0C",X"00",X"0D",X"00",X"0B",X"00",X"0C",X"00",X"0C",X"00",X"0D",X"00",X"0B",X"00",X"0D",X"00",
		X"0C",X"00",X"0D",X"00",X"0B",X"00",X"0C",X"00",X"0D",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",
		X"0C",X"00",X"0B",X"00",X"0C",X"00",X"0B",X"00",X"0C",X"00",X"0C",X"00",X"0E",X"00",X"0C",X"00",
		X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0B",X"00",X"0D",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",
		X"0C",X"00",X"0E",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0B",X"00",X"0C",X"00",X"0C",X"00",
		X"0B",X"00",X"0D",X"00",X"0C",X"00",X"0D",X"00",X"0B",X"00",X"0C",X"00",X"0D",X"00",X"0C",X"00",
		X"0A",X"00",X"0C",X"00",X"0C",X"00",X"0B",X"00",X"0B",X"00",X"0B",X"00",X"0B",X"00",X"0B",X"00",
		X"0B",X"00",X"0B",X"00",X"0B",X"00",X"0C",X"00",X"0A",X"00",X"0B",X"00",X"0B",X"00",X"0B",X"00",
		X"0B",X"00",X"0A",X"00",X"0C",X"00",X"0A",X"00",X"0B",X"00",X"0A",X"00",X"0B",X"00",X"0B",X"00",
		X"0A",X"00",X"0B",X"00",X"0B",X"00",X"0A",X"00",X"0B",X"00",X"0B",X"00",X"0B",X"00",X"0A",X"00",
		X"0A",X"00",X"0B",X"00",X"0B",X"00",X"0B",X"00",X"0A",X"00",X"0B",X"00",X"0B",X"00",X"0A",X"00",
		X"0B",X"00",X"0B",X"00",X"0C",X"00",X"0B",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0B",X"00",
		X"0B",X"00",X"0A",X"00",X"0B",X"00",X"0A",X"00",X"0B",X"00",X"0B",X"00",X"0A",X"00",X"0C",X"00",
		X"0A",X"00",X"0B",X"00",X"0B",X"00",X"0B",X"00",X"0C",X"00",X"0B",X"00",X"0C",X"00",X"0B",X"00",
		X"0C",X"00",X"0B",X"00",X"0B",X"00",X"0A",X"00",X"0B",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",
		X"0B",X"00",X"0A",X"00",X"0B",X"00",X"0B",X"00",X"0B",X"00",X"0A",X"00",X"0C",X"00",X"0C",X"00",
		X"0D",X"00",X"0B",X"00",X"0B",X"00",X"0A",X"00",X"0C",X"00",X"0B",X"00",X"0B",X"00",X"0B",X"00",
		X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0B",X"00",X"0B",X"00",X"0B",X"00",X"0B",X"00",X"0B",X"00",
		X"0C",X"00",X"0B",X"00",X"0B",X"00",X"0B",X"00",X"0B",X"00",X"0B",X"00",X"0B",X"00",X"0A",X"00",
		X"0B",X"00",X"0B",X"00",X"0C",X"00",X"0B",X"00",X"0B",X"00",X"0B",X"00",X"0A",X"00",X"0A",X"00",
		X"0B",X"00",X"0B",X"00",X"0B",X"00",X"0A",X"00",X"0B",X"00",X"0B",X"00",X"0B",X"00",X"0B",X"00",
		X"0B",X"00",X"0B",X"00",X"0B",X"00",X"0A",X"00",X"0B",X"00",X"0B",X"00",X"0B",X"00",X"0B",X"00",
		X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0B",X"00",X"0C",X"00",X"0B",X"00",X"0B",X"00",X"0B",X"00",
		X"0B",X"00",X"0B",X"00",X"0B",X"00",X"0C",X"00",X"0B",X"00",X"0C",X"00",X"0A",X"00",X"0C",X"00",
		X"0C",X"00",X"0C",X"00",X"0B",X"00",X"0B",X"00",X"0B",X"00",X"0B",X"00",X"0B",X"00",X"0A",X"00",
		X"0A",X"00",X"0B",X"00",X"0C",X"00",X"0B",X"00",X"0C",X"00",X"0B",X"00",X"0B",X"00",X"0C",X"00",
		X"0B",X"00",X"0B",X"00",X"0A",X"00",X"0B",X"00",X"0A",X"00",X"0B",X"00",X"0C",X"00",X"0A",X"00",
		X"0A",X"00",X"0B",X"00",X"0A",X"00",X"0A",X"00",X"0B",X"00",X"0A",X"00",X"0A",X"00",X"0B",X"00",
		X"0B",X"00",X"0B",X"00",X"0C",X"00",X"0B",X"00",X"0B",X"00",X"0C",X"00",X"0B",X"00",X"0B",X"00",
		X"0C",X"00",X"0B",X"00",X"0B",X"00",X"0B",X"00",X"0A",X"00",X"0B",X"00",X"0B",X"00",X"0A",X"00",
		X"0B",X"00",X"0A",X"00",X"0B",X"00",X"0B",X"00",X"0B",X"00",X"0B",X"00",X"0B",X"00",X"0B",X"00",
		X"0B",X"00",X"0B",X"00",X"0C",X"00",X"0B",X"00",X"0B",X"00",X"0B",X"00",X"0B",X"00",X"0B",X"00",
		X"0B",X"00",X"0C",X"00",X"0B",X"00",X"0B",X"00",X"0B",X"00",X"0A",X"00",X"0B",X"00",X"0C",X"00",
		X"0A",X"00",X"0C",X"00",X"0A",X"00",X"0A",X"00",X"0B",X"00",X"0C",X"00",X"0B",X"00",X"0B",X"00",
		X"0C",X"00",X"0B",X"00",X"0B",X"00",X"0A",X"00",X"0B",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",
		X"0A",X"00",X"09",X"00",X"0A",X"00",X"0B",X"00",X"0B",X"00",X"0A",X"00",X"09",X"00",X"0A",X"00",
		X"0A",X"00",X"0A",X"00",X"0B",X"00",X"09",X"00",X"0A",X"00",X"09",X"00",X"0A",X"00",X"0B",X"00",
		X"0B",X"00",X"0A",X"00",X"0A",X"00",X"09",X"00",X"0A",X"00",X"0A",X"00",X"0C",X"00",X"0A",X"00",
		X"0B",X"00",X"0B",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0B",X"00",X"0A",X"00",X"09",X"00",
		X"0A",X"00",X"0B",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"09",X"00",
		X"0A",X"00",X"09",X"00",X"09",X"00",X"09",X"00",X"09",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",
		X"0A",X"00",X"0A",X"00",X"09",X"00",X"0A",X"00",X"0C",X"00",X"0A",X"00",X"0B",X"00",X"0A",X"00",
		X"0B",X"00",X"0B",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0B",X"00",X"0A",X"00",
		X"0A",X"00",X"09",X"00",X"09",X"00",X"0A",X"00",X"0A",X"00",X"09",X"00",X"0A",X"00",X"09",X"00",
		X"0B",X"00",X"0A",X"00",X"09",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0C",X"00",X"0B",X"00",
		X"0B",X"00",X"0B",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0B",X"00",X"0A",X"00",X"0A",X"00",
		X"0A",X"00",X"0B",X"00",X"0A",X"00",X"0B",X"00",X"0B",X"00",X"0A",X"00",X"0B",X"00",X"0B",X"00",
		X"09",X"00",X"09",X"00",X"09",X"00",X"0B",X"00",X"09",X"00",X"09",X"00",X"0A",X"00",X"0B",X"00",
		X"0A",X"00",X"0B",X"00",X"0B",X"00",X"09",X"00",X"09",X"00",X"09",X"00",X"09",X"00",X"0A",X"00",
		X"0A",X"00",X"0A",X"00",X"0A",X"00",X"09",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0B",X"00",
		X"0B",X"00",X"0A",X"00",X"0B",X"00",X"0B",X"00",X"0C",X"00",X"0A",X"00",X"09",X"00",X"0A",X"00",
		X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",
		X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"09",X"00",X"08",X"00",X"0A",X"00",
		X"0A",X"00",X"0B",X"00",X"0A",X"00",X"0A",X"00",X"09",X"00",X"0A",X"00",X"09",X"00",X"0A",X"00",
		X"09",X"00",X"0A",X"00",X"09",X"00",X"09",X"00",X"0B",X"00",X"0A",X"00",X"09",X"00",X"0B",X"00",
		X"09",X"00",X"0B",X"00",X"0A",X"00",X"0B",X"00",X"0A",X"00",X"09",X"00",X"0A",X"00",X"0A",X"00",
		X"0A",X"00",X"09",X"00",X"09",X"00",X"0B",X"00",X"09",X"00",X"09",X"00",X"0A",X"00",X"0B",X"00",
		X"09",X"00",X"0A",X"00",X"0A",X"00",X"0B",X"00",X"0B",X"00",X"09",X"00",X"0B",X"00",X"0A",X"00",
		X"0B",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"09",X"00",X"0A",X"00",X"0A",X"00",
		X"0A",X"00",X"09",X"00",X"0B",X"00",X"0A",X"00",X"0A",X"00",X"09",X"00",X"0A",X"00",X"0A",X"00",
		X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0B",X"00",X"09",X"00",X"0A",X"00",X"0B",X"00",X"0A",X"00",
		X"0A",X"00",X"09",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0B",X"00",X"09",X"00",
		X"09",X"00",X"0A",X"00",X"09",X"00",X"0B",X"00",X"0B",X"00",X"09",X"00",X"0B",X"00",X"0B",X"00",
		X"0B",X"00",X"09",X"00",X"0A",X"00",X"0A",X"00",X"0B",X"00",X"0A",X"00",X"0A",X"00",X"09",X"00",
		X"09",X"00",X"09",X"00",X"09",X"00",X"09",X"00",X"08",X"00",X"08",X"00",X"09",X"00",X"09",X"00",
		X"0A",X"00",X"09",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"09",X"00",X"09",X"00",X"09",X"00",
		X"09",X"00",X"09",X"00",X"09",X"00",X"09",X"00",X"09",X"00",X"09",X"00",X"09",X"00",X"0A",X"00",
		X"09",X"00",X"08",X"00",X"09",X"00",X"09",X"00",X"08",X"00",X"09",X"00",X"09",X"00",X"09",X"00",
		X"09",X"00",X"09",X"00",X"0A",X"00",X"09",X"00",X"09",X"00",X"08",X"00",X"09",X"00",X"09",X"00",
		X"09",X"00",X"09",X"00",X"09",X"00",X"09",X"00",X"0A",X"00",X"08",X"00",X"09",X"00",X"09",X"00",
		X"09",X"00",X"09",X"00",X"09",X"00",X"09",X"00",X"0A",X"00",X"08",X"00",X"09",X"00",X"09",X"00",
		X"09",X"00",X"09",X"00",X"09",X"00",X"09",X"00",X"0A",X"00",X"0A",X"00",X"09",X"00",X"09",X"00",
		X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"09",X"00",X"09",X"00",X"08",X"00",
		X"08",X"00",X"08",X"00",X"09",X"00",X"09",X"00",X"0A",X"00",X"09",X"00",X"09",X"00",X"0A",X"00",
		X"0A",X"00",X"0A",X"00",X"09",X"00",X"09",X"00",X"09",X"00",X"09",X"00",X"09",X"00",X"08",X"00",
		X"09",X"00",X"0A",X"00",X"08",X"00",X"09",X"00",X"08",X"00",X"09",X"00",X"09",X"00",X"09",X"00",
		X"09",X"00",X"09",X"00",X"09",X"00",X"09",X"00",X"09",X"00",X"09",X"00",X"08",X"00",X"09",X"00",
		X"09",X"00",X"08",X"00",X"09",X"00",X"0A",X"00",X"08",X"00",X"0A",X"00",X"08",X"00",X"09",X"00",
		X"09",X"00",X"09",X"00",X"09",X"00",X"09",X"00",X"08",X"00",X"08",X"00",X"0A",X"00",X"09",X"00",
		X"09",X"00",X"09",X"00",X"09",X"00",X"0B",X"00",X"09",X"00",X"09",X"00",X"09",X"00",X"09",X"00",
		X"0A",X"00",X"08",X"00",X"08",X"00",X"0A",X"00",X"09",X"00",X"09",X"00",X"0A",X"00",X"09",X"00",
		X"09",X"00",X"09",X"00",X"09",X"00",X"09",X"00",X"08",X"00",X"09",X"00",X"08",X"00",X"09",X"00",
		X"0A",X"00",X"09",X"00",X"08",X"00",X"08",X"00",X"0A",X"00",X"09",X"00",X"09",X"00",X"08",X"00",
		X"08",X"00",X"0A",X"00",X"0B",X"00",X"08",X"00",X"09",X"00",X"09",X"00",X"09",X"00",X"08",X"00",
		X"09",X"00",X"0A",X"00",X"09",X"00",X"09",X"00",X"09",X"00",X"0A",X"00",X"0A",X"00",X"0B",X"00",
		X"09",X"00",X"09",X"00",X"09",X"00",X"0A",X"00",X"08",X"00",X"09",X"00",X"09",X"00",X"09",X"00",
		X"09",X"00",X"0A",X"00",X"09",X"00",X"09",X"00",X"09",X"00",X"0A",X"00",X"08",X"00",X"09",X"00",
		X"09",X"00",X"09",X"00",X"08",X"00",X"09",X"00",X"09",X"00",X"09",X"00",X"09",X"00",X"09",X"00",
		X"0A",X"00",X"0A",X"00",X"0A",X"00",X"09",X"00",X"09",X"00",X"09",X"00",X"09",X"00",X"09",X"00",
		X"09",X"00",X"09",X"00",X"0A",X"00",X"09",X"00",X"0A",X"00",X"09",X"00",X"09",X"00",X"08",X"00",
		X"09",X"00",X"09",X"00",X"08",X"00",X"08",X"00",X"09",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",
		X"0A",X"00",X"09",X"00",X"09",X"00",X"08",X"00",X"09",X"00",X"09",X"00",X"09",X"00",X"09",X"00",
		X"09",X"00",X"08",X"00",X"0A",X"00",X"09",X"00",X"08",X"00",X"09",X"00",X"08",X"00",X"08",X"00",
		X"09",X"00",X"08",X"00",X"09",X"00",X"09",X"00",X"09",X"00",X"08",X"00",X"09",X"00",X"0A",X"00",
		X"09",X"00",X"0A",X"00",X"09",X"00",X"0A",X"00",X"08",X"00",X"09",X"00",X"09",X"00",X"09",X"00",
		X"09",X"00",X"07",X"00",X"08",X"00",X"07",X"00",X"08",X"00",X"08",X"00",X"09",X"00",X"09",X"00",
		X"08",X"00",X"09",X"00",X"08",X"00",X"09",X"00",X"07",X"00",X"08",X"00",X"09",X"00",X"09",X"00",
		X"09",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"09",X"00",X"08",X"00",X"08",X"00",X"07",X"00",
		X"07",X"00",X"07",X"00",X"07",X"00",X"08",X"00",X"08",X"00",X"07",X"00",X"09",X"00",X"0A",X"00",
		X"08",X"00",X"09",X"00",X"08",X"00",X"08",X"00",X"09",X"00",X"08",X"00",X"08",X"00",X"07",X"00",
		X"08",X"00",X"07",X"00",X"08",X"00",X"07",X"00",X"08",X"00",X"08",X"00",X"09",X"00",X"08",X"00",
		X"08",X"00",X"07",X"00",X"09",X"00",X"09",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"09",X"00",
		X"08",X"00",X"08",X"00",X"09",X"00",X"08",X"00",X"08",X"00",X"09",X"00",X"08",X"00",X"06",X"00",
		X"09",X"00",X"09",X"00",X"08",X"00",X"08",X"00",X"09",X"00",X"08",X"00",X"06",X"00",X"09",X"00",
		X"08",X"00",X"07",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",
		X"07",X"00",X"09",X"00",X"07",X"00",X"07",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",
		X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"09",X"00",X"08",X"00",X"07",X"00",X"08",X"00",
		X"08",X"00",X"08",X"00",X"0A",X"00",X"08",X"00",X"09",X"00",X"08",X"00",X"08",X"00",X"08",X"00",
		X"09",X"00",X"09",X"00",X"08",X"00",X"09",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"09",X"00",
		X"09",X"00",X"09",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"07",X"00",X"08",X"00",X"08",X"00",
		X"09",X"00",X"08",X"00",X"07",X"00",X"07",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"07",X"00",
		X"07",X"00",X"09",X"00",X"09",X"00",X"0A",X"00",X"08",X"00",X"08",X"00",X"07",X"00",X"08",X"00",
		X"08",X"00",X"07",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"07",X"00",X"08",X"00",X"08",X"00",
		X"07",X"00",X"08",X"00",X"09",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"07",X"00",X"08",X"00",
		X"08",X"00",X"08",X"00",X"07",X"00",X"07",X"00",X"08",X"00",X"08",X"00",X"09",X"00",X"08",X"00",
		X"07",X"00",X"08",X"00",X"07",X"00",X"08",X"00",X"0A",X"00",X"09",X"00",X"08",X"00",X"08",X"00",
		X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"07",X"00",X"08",X"00",X"09",X"00",
		X"09",X"00",X"08",X"00",X"08",X"00",X"09",X"00",X"08",X"00",X"07",X"00",X"08",X"00",X"07",X"00",
		X"07",X"00",X"08",X"00",X"09",X"00",X"07",X"00",X"08",X"00",X"08",X"00",X"07",X"00",X"08",X"00",
		X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"09",X"00",X"09",X"00",
		X"08",X"00",X"07",X"00",X"09",X"00",X"07",X"00",X"08",X"00",X"06",X"00",X"08",X"00",X"08",X"00",
		X"09",X"00",X"08",X"00",X"09",X"00",X"09",X"00",X"08",X"00",X"07",X"00",X"08",X"00",X"07",X"00",
		X"06",X"00",X"07",X"00",X"08",X"00",X"07",X"00",X"08",X"00",X"08",X"00",X"09",X"00",X"08",X"00",
		X"08",X"00",X"09",X"00",X"08",X"00",X"08",X"00",X"06",X"00",X"09",X"00",X"08",X"00",X"08",X"00",
		X"09",X"00",X"07",X"00",X"08",X"00",X"09",X"00",X"09",X"00",X"07",X"00",X"09",X"00",X"08",X"00",
		X"08",X"00",X"08",X"00",X"07",X"00",X"08",X"00",X"0A",X"00",X"09",X"00",X"08",X"00",X"08",X"00",
		X"08",X"00",X"07",X"00",X"08",X"00",X"09",X"00",X"06",X"00",X"07",X"00",X"08",X"00",X"08",X"00",
		X"08",X"00",X"08",X"00",X"09",X"00",X"07",X"00",X"07",X"00",X"08",X"00",X"08",X"00",X"07",X"00",
		X"08",X"00",X"09",X"00",X"09",X"00",X"09",X"00",X"08",X"00",X"08",X"00",X"09",X"00",X"08",X"00",
		X"09",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"07",X"00",
		X"07",X"00",X"08",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"06",X"00",X"07",X"00",X"07",X"00",
		X"08",X"00",X"06",X"00",X"07",X"00",X"06",X"00",X"08",X"00",X"07",X"00",X"07",X"00",X"06",X"00",
		X"07",X"00",X"07",X"00",X"07",X"00",X"06",X"00",X"09",X"00",X"07",X"00",X"07",X"00",X"07",X"00",
		X"06",X"00",X"05",X"00",X"06",X"00",X"07",X"00",X"06",X"00",X"06",X"00",X"08",X"00",X"06",X"00",
		X"07",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"06",X"00",X"08",X"00",
		X"06",X"00",X"07",X"00",X"08",X"00",X"07",X"00",X"07",X"00",X"09",X"00",X"07",X"00",X"06",X"00",
		X"06",X"00",X"06",X"00",X"07",X"00",X"07",X"00",X"06",X"00",X"07",X"00",X"08",X"00",X"07",X"00",
		X"07",X"00",X"07",X"00",X"06",X"00",X"06",X"00",X"08",X"00",X"06",X"00",X"07",X"00",X"07",X"00",
		X"08",X"00",X"06",X"00",X"07",X"00",X"07",X"00",X"06",X"00",X"08",X"00",X"08",X"00",X"07",X"00",
		X"07",X"00",X"07",X"00",X"06",X"00",X"06",X"00",X"07",X"00",X"07",X"00",X"08",X"00",X"08",X"00",
		X"07",X"00",X"09",X"00",X"08",X"00",X"07",X"00",X"08",X"00",X"07",X"00",X"07",X"00",X"06",X"00",
		X"07",X"00",X"07",X"00",X"07",X"00",X"06",X"00",X"07",X"00",X"06",X"00",X"08",X"00",X"07",X"00",
		X"08",X"00",X"06",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"06",X"00",X"07",X"00",
		X"06",X"00",X"07",X"00",X"06",X"00",X"07",X"00",X"06",X"00",X"07",X"00",X"07",X"00",X"06",X"00",
		X"07",X"00",X"07",X"00",X"08",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"08",X"00",X"07",X"00",
		X"06",X"00",X"06",X"00",X"05",X"00",X"07",X"00",X"07",X"00",X"08",X"00",X"08",X"00",X"07",X"00",
		X"08",X"00",X"09",X"00",X"08",X"00",X"09",X"00",X"07",X"00",X"06",X"00",X"06",X"00",X"07",X"00",
		X"07",X"00",X"06",X"00",X"07",X"00",X"07",X"00",X"08",X"00",X"08",X"00",X"07",X"00",X"07",X"00",
		X"07",X"00",X"06",X"00",X"06",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"06",X"00",
		X"07",X"00",X"06",X"00",X"07",X"00",X"06",X"00",X"08",X"00",X"07",X"00",X"08",X"00",X"08",X"00",
		X"07",X"00",X"07",X"00",X"08",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"07",X"00",
		X"07",X"00",X"08",X"00",X"08",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"06",X"00",
		X"06",X"00",X"06",X"00",X"08",X"00",X"07",X"00",X"08",X"00",X"07",X"00",X"07",X"00",X"07",X"00",
		X"08",X"00",X"07",X"00",X"08",X"00",X"07",X"00",X"07",X"00",X"06",X"00",X"08",X"00",X"07",X"00",
		X"08",X"00",X"07",X"00",X"06",X"00",X"07",X"00",X"07",X"00",X"06",X"00",X"06",X"00",X"07",X"00",
		X"07",X"00",X"08",X"00",X"06",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"06",X"00",X"07",X"00",
		X"08",X"00",X"07",X"00",X"08",X"00",X"07",X"00",X"07",X"00",X"06",X"00",X"07",X"00",X"07",X"00",
		X"07",X"00",X"08",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"07",X"00",
		X"06",X"00",X"07",X"00",X"08",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"06",X"00",X"06",X"00",
		X"07",X"00",X"07",X"00",X"05",X"00",X"07",X"00",X"08",X"00",X"07",X"00",X"06",X"00",X"07",X"00",
		X"08",X"00",X"06",X"00",X"07",X"00",X"08",X"00",X"07",X"00",X"07",X"00",X"08",X"00",X"07",X"00",
		X"08",X"00",X"08",X"00",X"06",X"00",X"07",X"00",X"08",X"00",X"07",X"00",X"06",X"00",X"06",X"00",
		X"07",X"00",X"07",X"00",X"07",X"00",X"08",X"00",X"07",X"00",X"07",X"00",X"09",X"00",X"06",X"00",
		X"07",X"00",X"07",X"00",X"07",X"00",X"06",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"07",X"00",
		X"06",X"00",X"07",X"00",X"06",X"00",X"07",X"00",X"08",X"00",X"07",X"00",X"06",X"00",X"07",X"00",
		X"07",X"00",X"07",X"00",X"07",X"00",X"08",X"00",X"06",X"00",X"07",X"00",X"08",X"00",X"07",X"00",
		X"06",X"00",X"08",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"07",X"00",
		X"08",X"00",X"06",X"00",X"06",X"00",X"07",X"00",X"07",X"00",X"06",X"00",X"06",X"00",X"07",X"00",
		X"05",X"00",X"06",X"00",X"06",X"00",X"06",X"00",X"06",X"00",X"06",X"00",X"05",X"00",X"07",X"00",
		X"06",X"00",X"06",X"00",X"06",X"00",X"06",X"00",X"06",X"00",X"06",X"00",X"06",X"00",X"06",X"00",
		X"05",X"00",X"05",X"00",X"06",X"00",X"06",X"00",X"06",X"00",X"07",X"00",X"06",X"00",X"06",X"00",
		X"05",X"00",X"06",X"00",X"06",X"00",X"07",X"00",X"05",X"00",X"07",X"00",X"06",X"00",X"06",X"00",
		X"07",X"00",X"06",X"00",X"05",X"00",X"06",X"00",X"06",X"00",X"07",X"00",X"05",X"00",X"07",X"00",
		X"05",X"00",X"07",X"00",X"06",X"00",X"08",X"00",X"06",X"00",X"06",X"00",X"06",X"00",X"06",X"00",
		X"06",X"00",X"06",X"00",X"06",X"00",X"06",X"00",X"05",X"00",X"06",X"00",X"05",X"00",X"06",X"00",
		X"07",X"00",X"07",X"00",X"06",X"00",X"08",X"00",X"06",X"00",X"05",X"00",X"04",X"00",X"05",X"00",
		X"07",X"00",X"06",X"00",X"05",X"00",X"07",X"00",X"06",X"00",X"06",X"00",X"06",X"00",X"05",X"00",
		X"06",X"00",X"06",X"00",X"06",X"00",X"07",X"00",X"06",X"00",X"05",X"00",X"06",X"00",X"06",X"00",
		X"07",X"00",X"06",X"00",X"06",X"00",X"06",X"00",X"05",X"00",X"06",X"00",X"06",X"00",X"07",X"00",
		X"06",X"00",X"06",X"00",X"06",X"00",X"06",X"00",X"06",X"00",X"06",X"00",X"05",X"00",X"08",X"00",
		X"06",X"00",X"06",X"00",X"07",X"00",X"06",X"00",X"06",X"00",X"05",X"00",X"06",X"00",X"07",X"00",
		X"06",X"00",X"06",X"00",X"05",X"00",X"06",X"00",X"06",X"00",X"06",X"00",X"06",X"00",X"07",X"00",
		X"06",X"00",X"06",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"06",X"00",X"06",X"00",
		X"06",X"00",X"06",X"00",X"06",X"00",X"07",X"00",X"06",X"00",X"06",X"00",X"06",X"00",X"06",X"00",
		X"07",X"00",X"06",X"00",X"07",X"00",X"07",X"00",X"06",X"00",X"06",X"00",X"05",X"00",X"06",X"00",
		X"05",X"00",X"05",X"00",X"06",X"00",X"06",X"00",X"06",X"00",X"05",X"00",X"05",X"00",X"06",X"00",
		X"06",X"00",X"06",X"00",X"06",X"00",X"06",X"00",X"05",X"00",X"06",X"00",X"06",X"00",X"06",X"00",
		X"06",X"00",X"06",X"00",X"07",X"00",X"06",X"00",X"06",X"00",X"06",X"00",X"06",X"00",X"05",X"00",
		X"05",X"00",X"07",X"00",X"07",X"00",X"05",X"00",X"06",X"00",X"07",X"00",X"07",X"00",X"07",X"00",
		X"05",X"00",X"05",X"00",X"06",X"00",X"06",X"00",X"07",X"00",X"07",X"00",X"06",X"00",X"06",X"00",
		X"06",X"00",X"06",X"00",X"06",X"00",X"05",X"00",X"06",X"00",X"06",X"00",X"05",X"00",X"06",X"00",
		X"07",X"00",X"06",X"00",X"07",X"00",X"06",X"00",X"06",X"00",X"06",X"00",X"06",X"00",X"06",X"00",
		X"06",X"00",X"05",X"00",X"06",X"00",X"06",X"00",X"06",X"00",X"06",X"00",X"05",X"00",X"06",X"00",
		X"06",X"00",X"06",X"00",X"06",X"00",X"07",X"00",X"06",X"00",X"05",X"00",X"05",X"00",X"05",X"00",
		X"06",X"00",X"06",X"00",X"06",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"06",X"00",X"06",X"00",
		X"06",X"00",X"07",X"00",X"05",X"00",X"05",X"00",X"06",X"00",X"07",X"00",X"06",X"00",X"06",X"00",
		X"05",X"00",X"06",X"00",X"06",X"00",X"07",X"00",X"07",X"00",X"05",X"00",X"06",X"00",X"05",X"00",
		X"06",X"00",X"06",X"00",X"06",X"00",X"06",X"00",X"05",X"00",X"06",X"00",X"07",X"00",X"06",X"00",
		X"06",X"00",X"06",X"00",X"06",X"00",X"05",X"00",X"06",X"00",X"06",X"00",X"06",X"00",X"06",X"00",
		X"06",X"00",X"06",X"00",X"06",X"00",X"07",X"00",X"06",X"00",X"06",X"00",X"06",X"00",X"06",X"00",
		X"06",X"00",X"06",X"00",X"07",X"00",X"06",X"00",X"06",X"00",X"05",X"00",X"06",X"00",X"05",X"00",
		X"05",X"00",X"06",X"00",X"06",X"00",X"05",X"00",X"05",X"00",X"06",X"00",X"06",X"00",X"06",X"00",
		X"06",X"00",X"06",X"00",X"05",X"00",X"07",X"00",X"06",X"00",X"04",X"00",X"06",X"00",X"06",X"00",
		X"06",X"00",X"06",X"00",X"06",X"00",X"06",X"00",X"06",X"00",X"06",X"00",X"07",X"00",X"06",X"00",
		X"06",X"00",X"05",X"00",X"06",X"00",X"06",X"00",X"04",X"00",X"06",X"00",X"07",X"00",X"06",X"00",
		X"06",X"00",X"06",X"00",X"06",X"00",X"05",X"00",X"07",X"00",X"05",X"00",X"06",X"00",X"05",X"00",
		X"06",X"00",X"05",X"00",X"05",X"00",X"06",X"00",X"05",X"00",X"06",X"00",X"06",X"00",X"06",X"00",
		X"06",X"00",X"06",X"00",X"06",X"00",X"08",X"00",X"05",X"00",X"06",X"00",X"07",X"00",X"06",X"00",
		X"06",X"00",X"06",X"00",X"05",X"00",X"06",X"00",X"06",X"00",X"07",X"00",X"05",X"00",X"06",X"00",
		X"06",X"00",X"07",X"00",X"07",X"00",X"06",X"00",X"07",X"00",X"06",X"00",X"07",X"00",X"06",X"00",
		X"06",X"00",X"05",X"00",X"07",X"00",X"06",X"00",X"05",X"00",X"04",X"00",X"05",X"00",X"06",X"00",
		X"05",X"00",X"06",X"00",X"04",X"00",X"05",X"00",X"06",X"00",X"05",X"00",X"05",X"00",X"04",X"00",
		X"05",X"00",X"05",X"00",X"06",X"00",X"04",X"00",X"04",X"00",X"06",X"00",X"05",X"00",X"06",X"00",
		X"06",X"00",X"05",X"00",X"06",X"00",X"05",X"00",X"04",X"00",X"05",X"00",X"05",X"00",X"05",X"00",
		X"06",X"00",X"07",X"00",X"05",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"05",X"00",
		X"05",X"00",X"05",X"00",X"07",X"00",X"06",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",
		X"05",X"00",X"05",X"00",X"05",X"00",X"06",X"00",X"06",X"00",X"04",X"00",X"05",X"00",X"06",X"00",
		X"05",X"00",X"04",X"00",X"06",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",
		X"05",X"00",X"05",X"00",X"04",X"00",X"04",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",
		X"07",X"00",X"05",X"00",X"06",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"04",X"00",X"04",X"00",
		X"05",X"00",X"06",X"00",X"06",X"00",X"04",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",
		X"04",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"04",X"00",X"05",X"00",
		X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"06",X"00",X"05",X"00",X"05",X"00",X"04",X"00",
		X"05",X"00",X"05",X"00",X"04",X"00",X"04",X"00",X"05",X"00",X"07",X"00",X"05",X"00",X"06",X"00",
		X"04",X"00",X"04",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"04",X"00",X"06",X"00",X"06",X"00",
		X"04",X"00",X"05",X"00",X"06",X"00",X"04",X"00",X"05",X"00",X"05",X"00",X"04",X"00",X"03",X"00",
		X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"06",X"00",
		X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"06",X"00",X"06",X"00",X"05",X"00",
		X"04",X"00",X"05",X"00",X"05",X"00",X"04",X"00",X"05",X"00",X"05",X"00",X"06",X"00",X"06",X"00",
		X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"04",X"00",X"05",X"00",
		X"06",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"06",X"00",X"06",X"00",
		X"04",X"00",X"05",X"00",X"04",X"00",X"06",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",
		X"05",X"00",X"06",X"00",X"04",X"00",X"05",X"00",X"05",X"00",X"04",X"00",X"05",X"00",X"05",X"00",
		X"05",X"00",X"05",X"00",X"06",X"00",X"05",X"00",X"04",X"00",X"05",X"00",X"05",X"00",X"05",X"00",
		X"05",X"00",X"07",X"00",X"04",X"00",X"04",X"00",X"05",X"00",X"06",X"00",X"07",X"00",X"05",X"00",
		X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"03",X"00",X"05",X"00",X"04",X"00",
		X"05",X"00",X"04",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"04",X"00",X"05",X"00",
		X"05",X"00",X"04",X"00",X"06",X"00",X"05",X"00",X"06",X"00",X"06",X"00",X"05",X"00",X"06",X"00",
		X"05",X"00",X"06",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"07",X"00",X"05",X"00",X"05",X"00",
		X"04",X"00",X"06",X"00",X"05",X"00",X"05",X"00",X"04",X"00",X"05",X"00",X"04",X"00",X"04",X"00",
		X"05",X"00",X"05",X"00",X"05",X"00",X"04",X"00",X"05",X"00",X"04",X"00",X"04",X"00",X"05",X"00",
		X"04",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"06",X"00",X"07",X"00",X"07",X"00",X"05",X"00",
		X"05",X"00",X"05",X"00",X"06",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",
		X"05",X"00",X"05",X"00",X"05",X"00",X"06",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"04",X"00",
		X"07",X"00",X"05",X"00",X"04",X"00",X"05",X"00",X"05",X"00",X"06",X"00",X"06",X"00",X"05",X"00",
		X"04",X"00",X"05",X"00",X"05",X"00",X"06",X"00",X"05",X"00",X"06",X"00",X"05",X"00",X"05",X"00",
		X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"06",X"00",X"04",X"00",X"04",X"00",X"06",X"00",
		X"05",X"00",X"04",X"00",X"05",X"00",X"06",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",
		X"05",X"00",X"06",X"00",X"05",X"00",X"06",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"06",X"00",
		X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"04",X"00",
		X"04",X"00",X"05",X"00",X"06",X"00",X"04",X"00",X"06",X"00",X"04",X"00",X"05",X"00",X"05",X"00",
		X"04",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"06",X"00",X"06",X"00",X"05",X"00",
		X"06",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"04",X"00",X"05",X"00",X"05",X"00",
		X"05",X"00",X"05",X"00",X"05",X"00",X"06",X"00",X"05",X"00",X"05",X"00",X"06",X"00",X"04",X"00",
		X"04",X"00",X"05",X"00",X"06",X"00",X"04",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"04",X"00",
		X"04",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"04",X"00",X"05",X"00",X"05",X"00",X"07",X"00",
		X"05",X"00",X"07",X"00",X"05",X"00",X"04",X"00",X"05",X"00",X"07",X"00",X"05",X"00",X"05",X"00",
		X"05",X"00",X"05",X"00",X"05",X"00",X"06",X"00",X"05",X"00",X"04",X"00",X"05",X"00",X"05",X"00",
		X"05",X"00",X"05",X"00",X"05",X"00",X"04",X"00",X"05",X"00",X"06",X"00",X"04",X"00",X"06",X"00",
		X"04",X"00",X"05",X"00",X"05",X"00",X"06",X"00",X"05",X"00",X"04",X"00",X"05",X"00",X"05",X"00",
		X"04",X"00",X"05",X"00",X"04",X"00",X"06",X"00",X"04",X"00",X"05",X"00",X"05",X"00",X"06",X"00",
		X"05",X"00",X"05",X"00",X"05",X"00",X"04",X"00",X"04",X"00",X"03",X"00",X"05",X"00",X"05",X"00",
		X"05",X"00",X"03",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",
		X"05",X"00",X"03",X"00",X"04",X"00",X"03",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",
		X"04",X"00",X"05",X"00",X"04",X"00",X"05",X"00",X"04",X"00",X"05",X"00",X"05",X"00",X"03",X"00",
		X"03",X"00",X"04",X"00",X"05",X"00",X"06",X"00",X"04",X"00",X"03",X"00",X"03",X"00",X"04",X"00",
		X"04",X"00",X"04",X"00",X"03",X"00",X"04",X"00",X"04",X"00",X"03",X"00",X"04",X"00",X"03",X"00",
		X"05",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"05",X"00",
		X"03",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"05",X"00",X"03",X"00",X"04",X"00",X"04",X"00",
		X"05",X"00",X"04",X"00",X"04",X"00",X"03",X"00",X"05",X"00",X"04",X"00",X"04",X"00",X"04",X"00",
		X"04",X"00",X"04",X"00",X"05",X"00",X"04",X"00",X"05",X"00",X"05",X"00",X"03",X"00",X"04",X"00",
		X"04",X"00",X"04",X"00",X"05",X"00",X"05",X"00",X"04",X"00",X"05",X"00",X"05",X"00",X"03",X"00",
		X"04",X"00",X"04",X"00",X"03",X"00",X"05",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"05",X"00",
		X"04",X"00",X"04",X"00",X"03",X"00",X"03",X"00",X"04",X"00",X"03",X"00",X"04",X"00",X"04",X"00",
		X"02",X"00",X"04",X"00",X"04",X"00",X"03",X"00",X"04",X"00",X"05",X"00",X"06",X"00",X"04",X"00",
		X"04",X"00",X"04",X"00",X"04",X"00",X"03",X"00",X"06",X"00",X"05",X"00",X"04",X"00",X"04",X"00",
		X"05",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"04",X"00",X"04",X"00",X"05",X"00",
		X"04",X"00",X"04",X"00",X"05",X"00",X"05",X"00",X"04",X"00",X"04",X"00",X"05",X"00",X"03",X"00",
		X"04",X"00",X"05",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"06",X"00",X"03",X"00",
		X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"05",X"00",X"04",X"00",
		X"04",X"00",X"04",X"00",X"03",X"00",X"05",X"00",X"04",X"00",X"03",X"00",X"05",X"00",X"04",X"00",
		X"05",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"03",X"00",X"04",X"00",X"03",X"00",
		X"03",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"03",X"00",X"05",X"00",X"03",X"00",
		X"04",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"06",X"00",X"03",X"00",
		X"05",X"00",X"04",X"00",X"05",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"05",X"00",X"04",X"00",
		X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"03",X"00",X"04",X"00",
		X"05",X"00",X"04",X"00",X"04",X"00",X"03",X"00",X"03",X"00",X"04",X"00",X"04",X"00",X"04",X"00",
		X"05",X"00",X"04",X"00",X"03",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"03",X"00",X"04",X"00",
		X"04",X"00",X"04",X"00",X"05",X"00",X"03",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"03",X"00",
		X"03",X"00",X"04",X"00",X"04",X"00",X"05",X"00",X"04",X"00",X"05",X"00",X"05",X"00",X"04",X"00",
		X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"05",X"00",X"04",X"00",X"04",X"00",X"04",X"00",
		X"05",X"00",X"04",X"00",X"05",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"05",X"00",X"04",X"00",
		X"04",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"03",X"00",X"05",X"00",X"03",X"00",X"04",X"00",
		X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"05",X"00",X"05",X"00",
		X"04",X"00",X"03",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"03",X"00",X"03",X"00",X"04",X"00",
		X"03",X"00",X"04",X"00",X"05",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"03",X"00",
		X"03",X"00",X"04",X"00",X"02",X"00",X"04",X"00",X"05",X"00",X"04",X"00",X"02",X"00",X"05",X"00",
		X"04",X"00",X"05",X"00",X"04",X"00",X"05",X"00",X"03",X"00",X"04",X"00",X"05",X"00",X"03",X"00",
		X"04",X"00",X"05",X"00",X"04",X"00",X"04",X"00",X"05",X"00",X"04",X"00",X"04",X"00",X"06",X"00",
		X"05",X"00",X"04",X"00",X"05",X"00",X"04",X"00",X"04",X"00",X"06",X"00",X"04",X"00",X"04",X"00",
		X"05",X"00",X"04",X"00",X"03",X"00",X"04",X"00",X"05",X"00",X"04",X"00",X"04",X"00",X"04",X"00",
		X"04",X"00",X"05",X"00",X"05",X"00",X"03",X"00",X"04",X"00",X"05",X"00",X"04",X"00",X"04",X"00",
		X"04",X"00",X"04",X"00",X"04",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"04",X"00",X"04",X"00",
		X"04",X"00",X"03",X"00",X"03",X"00",X"04",X"00",X"04",X"00",X"05",X"00",X"04",X"00",X"04",X"00",
		X"05",X"00",X"05",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"03",X"00",X"04",X"00",X"04",X"00",
		X"04",X"00",X"03",X"00",X"04",X"00",X"05",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"05",X"00",
		X"05",X"00",X"05",X"00",X"04",X"00",X"05",X"00",X"03",X"00",X"04",X"00",X"03",X"00",X"03",X"00",
		X"03",X"00",X"04",X"00",X"05",X"00",X"03",X"00",X"03",X"00",X"04",X"00",X"04",X"00",X"03",X"00",
		X"04",X"00",X"04",X"00",X"02",X"00",X"05",X"00",X"04",X"00",X"03",X"00",X"04",X"00",X"04",X"00",
		X"05",X"00",X"03",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"03",X"00",X"04",X"00",X"04",X"00",
		X"04",X"00",X"05",X"00",X"04",X"00",X"05",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",
		X"03",X"00",X"04",X"00",X"04",X"00",X"05",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"03",X"00",
		X"04",X"00",X"04",X"00",X"06",X"00",X"05",X"00",X"06",X"00",X"03",X"00",X"04",X"00",X"02",X"00",
		X"03",X"00",X"04",X"00",X"04",X"00",X"03",X"00",X"04",X"00",X"04",X"00",X"03",X"00",X"04",X"00",
		X"04",X"00",X"03",X"00",X"03",X"00",X"04",X"00",X"03",X"00",X"05",X"00",X"04",X"00",X"04",X"00",
		X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"03",X"00",X"05",X"00",X"03",X"00",X"04",X"00",
		X"03",X"00",X"04",X"00",X"05",X"00",X"04",X"00",X"03",X"00",X"03",X"00",X"06",X"00",X"04",X"00",
		X"05",X"00",X"04",X"00",X"05",X"00",X"05",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"05",X"00",
		X"04",X"00",X"04",X"00",X"03",X"00",X"04",X"00",X"05",X"00",X"04",X"00",X"05",X"00",X"04",X"00",
		X"05",X"00",X"04",X"00",X"05",X"00",X"05",X"00",X"02",X"00",X"03",X"00",X"04",X"00",X"02",X"00",
		X"02",X"00",X"04",X"00",X"05",X"00",X"04",X"00",X"05",X"00",X"03",X"00",X"05",X"00",X"04",X"00",
		X"03",X"00",X"04",X"00",X"04",X"00",X"03",X"00",X"04",X"00",X"03",X"00",X"03",X"00",X"06",X"00",
		X"03",X"00",X"04",X"00",X"04",X"00",X"03",X"00",X"04",X"00",X"05",X"00",X"04",X"00",X"04",X"00",
		X"05",X"00",X"04",X"00",X"03",X"00",X"04",X"00",X"03",X"00",X"04",X"00",X"02",X"00",X"04",X"00",
		X"03",X"00",X"02",X"00",X"03",X"00",X"03",X"00",X"01",X"00",X"03",X"00",X"03",X"00",X"03",X"00",
		X"04",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"02",X"00",X"04",X"00",X"04",X"00",
		X"03",X"00",X"03",X"00",X"02",X"00",X"01",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",
		X"03",X"00",X"04",X"00",X"04",X"00",X"02",X"00",X"03",X"00",X"03",X"00",X"04",X"00",X"04",X"00",
		X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"03",X"00",X"04",X"00",X"02",X"00",X"03",X"00",
		X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"02",X"00",X"04",X"00",X"03",X"00",X"03",X"00",
		X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"02",X"00",X"04",X"00",
		X"03",X"00",X"02",X"00",X"03",X"00",X"02",X"00",X"04",X"00",X"03",X"00",X"04",X"00",X"04",X"00",
		X"03",X"00",X"04",X"00",X"03",X"00",X"03",X"00",X"05",X"00",X"03",X"00",X"03",X"00",X"03",X"00",
		X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"04",X"00",X"04",X"00",X"02",X"00",X"02",X"00",
		X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"04",X"00",X"03",X"00",X"04",X"00",
		X"03",X"00",X"03",X"00",X"03",X"00",X"04",X"00",X"05",X"00",X"03",X"00",X"04",X"00",X"03",X"00",
		X"03",X"00",X"03",X"00",X"02",X"00",X"02",X"00",X"03",X"00",X"04",X"00",X"04",X"00",X"03",X"00",
		X"03",X"00",X"04",X"00",X"03",X"00",X"04",X"00",X"03",X"00",X"04",X"00",X"02",X"00",X"03",X"00",
		X"02",X"00",X"02",X"00",X"04",X"00",X"03",X"00",X"02",X"00",X"04",X"00",X"04",X"00",X"04",X"00",
		X"04",X"00",X"03",X"00",X"03",X"00",X"02",X"00",X"01",X"00",X"04",X"00",X"03",X"00",X"03",X"00",
		X"04",X"00",X"02",X"00",X"03",X"00",X"04",X"00",X"04",X"00",X"03",X"00",X"03",X"00",X"03",X"00",
		X"04",X"00",X"02",X"00",X"03",X"00",X"03",X"00",X"02",X"00",X"04",X"00",X"03",X"00",X"03",X"00",
		X"03",X"00",X"03",X"00",X"02",X"00",X"02",X"00",X"04",X"00",X"03",X"00",X"04",X"00",X"04",X"00",
		X"03",X"00",X"03",X"00",X"02",X"00",X"03",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"03",X"00",
		X"01",X"00",X"01",X"00",X"03",X"00",X"03",X"00",X"02",X"00",X"03",X"00",X"03",X"00",X"03",X"00",
		X"03",X"00",X"02",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"02",X"00",X"03",X"00",X"03",X"00",
		X"04",X"00",X"03",X"00",X"04",X"00",X"02",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",
		X"03",X"00",X"02",X"00",X"03",X"00",X"02",X"00",X"03",X"00",X"03",X"00",X"04",X"00",X"03",X"00",
		X"03",X"00",X"02",X"00",X"03",X"00",X"03",X"00",X"02",X"00",X"04",X"00",X"03",X"00",X"03",X"00",
		X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"02",X"00",X"03",X"00",X"03",X"00",X"04",X"00",
		X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"02",X"00",X"03",X"00",X"03",X"00",X"03",X"00",
		X"03",X"00",X"04",X"00",X"03",X"00",X"02",X"00",X"03",X"00",X"04",X"00",X"02",X"00",X"03",X"00",
		X"02",X"00",X"04",X"00",X"02",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",
		X"04",X"00",X"02",X"00",X"04",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"02",X"00",
		X"03",X"00",X"03",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"03",X"00",X"03",X"00",X"02",X"00",
		X"02",X"00",X"03",X"00",X"03",X"00",X"04",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",
		X"04",X"00",X"04",X"00",X"03",X"00",X"02",X"00",X"04",X"00",X"02",X"00",X"04",X"00",X"03",X"00",
		X"02",X"00",X"03",X"00",X"04",X"00",X"03",X"00",X"02",X"00",X"03",X"00",X"03",X"00",X"03",X"00",
		X"03",X"00",X"03",X"00",X"04",X"00",X"01",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",
		X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"04",X"00",X"04",X"00",X"02",X"00",X"03",X"00",
		X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"04",X"00",X"02",X"00",X"03",X"00",X"03",X"00",
		X"03",X"00",X"02",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"02",X"00",X"02",X"00",X"02",X"00",
		X"02",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"04",X"00",X"03",X"00",X"03",X"00",
		X"02",X"00",X"03",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"03",X"00",X"03",X"00",
		X"03",X"00",X"04",X"00",X"03",X"00",X"03",X"00",X"05",X"00",X"03",X"00",X"03",X"00",X"03",X"00",
		X"02",X"00",X"03",X"00",X"04",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"02",X"00",
		X"03",X"00",X"03",X"00",X"02",X"00",X"03",X"00",X"03",X"00",X"02",X"00",X"03",X"00",X"04",X"00",
		X"03",X"00",X"03",X"00",X"04",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",
		X"04",X"00",X"03",X"00",X"04",X"00",X"02",X"00",X"04",X"00",X"04",X"00",X"03",X"00",X"02",X"00",
		X"03",X"00",X"04",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"04",X"00",X"02",X"00",X"04",X"00",
		X"03",X"00",X"03",X"00",X"03",X"00",X"04",X"00",X"02",X"00",X"03",X"00",X"02",X"00",X"03",X"00",
		X"03",X"00",X"03",X"00",X"04",X"00",X"03",X"00",X"03",X"00",X"02",X"00",X"04",X"00",X"03",X"00",
		X"02",X"00",X"02",X"00",X"04",X"00",X"03",X"00",X"02",X"00",X"03",X"00",X"04",X"00",X"03",X"00",
		X"02",X"00",X"03",X"00",X"02",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"05",X"00",
		X"02",X"00",X"03",X"00",X"04",X"00",X"03",X"00",X"03",X"00",X"01",X"00",X"02",X"00",X"03",X"00",
		X"02",X"00",X"03",X"00",X"03",X"00",X"02",X"00",X"03",X"00",X"04",X"00",X"03",X"00",X"03",X"00",
		X"03",X"00",X"02",X"00",X"04",X"00",X"04",X"00",X"03",X"00",X"02",X"00",X"04",X"00",X"03",X"00",
		X"02",X"00",X"03",X"00",X"04",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",
		X"04",X"00",X"02",X"00",X"02",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"02",X"00",
		X"05",X"00",X"04",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"02",X"00",X"03",X"00",
		X"04",X"00",X"04",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"02",X"00",
		X"03",X"00",X"04",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"02",X"00",X"04",X"00",X"02",X"00",
		X"04",X"00",X"02",X"00",X"03",X"00",X"04",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"02",X"00",
		X"04",X"00",X"04",X"00",X"03",X"00",X"03",X"00",X"02",X"00",X"03",X"00",X"02",X"00",X"03",X"00",
		X"04",X"00",X"02",X"00",X"04",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"02",X"00",X"03",X"00",
		X"01",X"00",X"02",X"00",X"03",X"00",X"02",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",
		X"02",X"00",X"04",X"00",X"03",X"00",X"04",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",
		X"03",X"00",X"04",X"00",X"02",X"00",X"03",X"00",X"02",X"00",X"03",X"00",X"04",X"00",X"03",X"00",
		X"03",X"00",X"03",X"00",X"04",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"02",X"00",X"04",X"00",
		X"02",X"00",X"02",X"00",X"03",X"00",X"02",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"04",X"00",
		X"04",X"00",X"02",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",
		X"03",X"00",X"04",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"04",X"00",X"03",X"00",X"03",X"00",
		X"03",X"00",X"03",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"03",X"00",X"03",X"00",X"03",X"00",
		X"04",X"00",X"03",X"00",X"04",X"00",X"04",X"00",X"02",X"00",X"03",X"00",X"03",X"00",X"03",X"00",
		X"04",X"00",X"04",X"00",X"02",X"00",X"03",X"00",X"01",X"00",X"03",X"00",X"03",X"00",X"04",X"00",
		X"03",X"00",X"04",X"00",X"03",X"00",X"03",X"00",X"02",X"00",X"04",X"00",X"01",X"00",X"03",X"00",
		X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"03",X"00",X"03",X"00",X"04",X"00",X"02",X"00",
		X"03",X"00",X"03",X"00",X"04",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"04",X"00",X"03",X"00",
		X"04",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"03",X"00",X"03",X"00",X"04",X"00",X"04",X"00",
		X"04",X"00",X"03",X"00",X"02",X"00",X"03",X"00",X"03",X"00",X"04",X"00",X"03",X"00",X"03",X"00",
		X"04",X"00",X"04",X"00",X"03",X"00",X"02",X"00",X"04",X"00",X"02",X"00",X"03",X"00",X"03",X"00",
		X"03",X"00",X"02",X"00",X"03",X"00",X"03",X"00",X"04",X"00",X"03",X"00",X"03",X"00",X"03",X"00",
		X"02",X"00",X"04",X"00",X"02",X"00",X"04",X"00",X"03",X"00",X"03",X"00",X"04",X"00",X"02",X"00",
		X"03",X"00",X"03",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",
		X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"03",X"00",X"02",X"00",X"03",X"00",
		X"04",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"03",X"00",X"02",X"00",X"02",X"00",
		X"02",X"00",X"01",X"00",X"03",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"03",X"00",
		X"01",X"00",X"02",X"00",X"02",X"00",X"03",X"00",X"02",X"00",X"02",X"00",X"03",X"00",X"02",X"00",
		X"03",X"00",X"02",X"00",X"02",X"00",X"03",X"00",X"01",X"00",X"03",X"00",X"02",X"00",X"03",X"00",
		X"01",X"00",X"02",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"02",X"00",X"02",X"00",X"02",X"00",
		X"03",X"00",X"02",X"00",X"03",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"03",X"00",X"02",X"00",
		X"01",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"01",X"00",
		X"01",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"03",X"00",X"02",X"00",X"02",X"00",X"03",X"00",
		X"02",X"00",X"02",X"00",X"02",X"00",X"03",X"00",X"02",X"00",X"02",X"00",X"03",X"00",X"02",X"00",
		X"02",X"00",X"04",X"00",X"03",X"00",X"00",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"03",X"00",
		X"02",X"00",X"02",X"00",X"02",X"00",X"04",X"00",X"02",X"00",X"03",X"00",X"02",X"00",X"02",X"00",
		X"02",X"00",X"03",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",
		X"02",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"02",X"00",X"03",X"00",X"02",X"00",X"01",X"00",
		X"01",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"02",X"00",
		X"03",X"00",X"02",X"00",X"02",X"00",X"03",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"02",X"00",
		X"02",X"00",X"01",X"00",X"02",X"00",X"03",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"01",X"00",
		X"02",X"00",X"03",X"00",X"03",X"00",X"02",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"03",X"00",
		X"02",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"03",X"00",
		X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"03",X"00",X"01",X"00",
		X"03",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"02",X"00",
		X"02",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"01",X"00",X"02",X"00",X"03",X"00",X"01",X"00",
		X"02",X"00",X"03",X"00",X"03",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",
		X"02",X"00",X"02",X"00",X"03",X"00",X"04",X"00",X"03",X"00",X"02",X"00",X"01",X"00",X"01",X"00",
		X"03",X"00",X"02",X"00",X"03",X"00",X"03",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"03",X"00",
		X"02",X"00",X"03",X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"00",
		X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"02",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"03",X"00",X"03",X"00",X"02",X"00",X"03",X"00",
		X"03",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"02",X"00",
		X"02",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",
		X"02",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"02",X"00",
		X"02",X"00",X"03",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",
		X"01",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",
		X"02",X"00",X"03",X"00",X"02",X"00",X"01",X"00",X"03",X"00",X"02",X"00",X"01",X"00",X"02",X"00",
		X"02",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"03",X"00",X"02",X"00",X"02",X"00",
		X"01",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"03",X"00",X"03",X"00",X"02",X"00",X"03",X"00",
		X"02",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"03",X"00",
		X"03",X"00",X"02",X"00",X"04",X"00",X"02",X"00",X"02",X"00",X"03",X"00",X"03",X"00",X"02",X"00",
		X"03",X"00",X"02",X"00",X"01",X"00",X"03",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"04",X"00",
		X"01",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"03",X"00",X"02",X"00",X"02",X"00",X"03",X"00",
		X"03",X"00",X"03",X"00",X"03",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"02",X"00",
		X"03",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"03",X"00",X"02",X"00",X"02",X"00",
		X"03",X"00",X"01",X"00",X"03",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"03",X"00",
		X"03",X"00",X"02",X"00",X"01",X"00",X"03",X"00",X"02",X"00",X"02",X"00",X"04",X"00",X"02",X"00",
		X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"04",X"00",X"01",X"00",X"02",X"00",
		X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"02",X"00",
		X"01",X"00",X"03",X"00",X"02",X"00",X"03",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",
		X"01",X"00",X"03",X"00",X"02",X"00",X"02",X"00",X"03",X"00",X"02",X"00",X"02",X"00",X"02",X"00",
		X"03",X"00",X"03",X"00",X"02",X"00",X"03",X"00",X"02",X"00",X"04",X"00",X"03",X"00",X"02",X"00",
		X"02",X"00",X"03",X"00",X"02",X"00",X"03",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"02",X"00",
		X"03",X"00",X"04",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"02",X"00",
		X"00",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"01",X"00",
		X"02",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"03",X"00",X"02",X"00",
		X"01",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"03",X"00",X"02",X"00",X"01",X"00",X"02",X"00",
		X"03",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"01",X"00",X"02",X"00",X"02",X"00",
		X"03",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"03",X"00",X"01",X"00",X"02",X"00",X"02",X"00",
		X"02",X"00",X"01",X"00",X"03",X"00",X"02",X"00",X"02",X"00",X"03",X"00",X"02",X"00",X"03",X"00",
		X"03",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"03",X"00",
		X"03",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"03",X"00",X"00",X"00",X"02",X"00",X"02",X"00",
		X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"03",X"00",X"02",X"00",X"02",X"00",
		X"02",X"00",X"02",X"00",X"03",X"00",X"01",X"00",X"02",X"00",X"03",X"00",X"02",X"00",X"03",X"00",
		X"03",X"00",X"02",X"00",X"01",X"00",X"03",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"02",X"00",
		X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"01",X"00",X"02",X"00",X"03",X"00",X"01",X"00",
		X"02",X"00",X"00",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",
		X"01",X"00",X"02",X"00",X"03",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"02",X"00",
		X"03",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"01",X"00",
		X"03",X"00",X"00",X"00",X"02",X"00",X"03",X"00",X"02",X"00",X"02",X"00",X"03",X"00",X"02",X"00",
		X"01",X"00",X"02",X"00",X"03",X"00",X"01",X"00",X"01",X"00",X"03",X"00",X"02",X"00",X"02",X"00",
		X"03",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",
		X"02",X"00",X"02",X"00",X"03",X"00",X"02",X"00",X"01",X"00",X"03",X"00",X"02",X"00",X"02",X"00",
		X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"01",X"00",
		X"02",X"00",X"02",X"00",X"02",X"00",X"03",X"00",X"01",X"00",X"02",X"00",X"03",X"00",X"02",X"00",
		X"02",X"00",X"03",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",
		X"01",X"00",X"02",X"00",X"03",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"02",X"00",
		X"03",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"01",X"00",
		X"02",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"03",X"00",X"03",X"00",X"02",X"00",
		X"00",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",
		X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"03",X"00",X"02",X"00",X"02",X"00",X"02",X"00",
		X"02",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"00",X"00",X"03",X"00",X"02",X"00",
		X"02",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"02",X"00",
		X"01",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"03",X"00",
		X"03",X"00",X"03",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"02",X"00",
		X"02",X"00",X"02",X"00",X"00",X"00",X"03",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"02",X"00",
		X"01",X"00",X"02",X"00",X"01",X"00",X"03",X"00",X"02",X"00",X"03",X"00",X"02",X"00",X"01",X"00",
		X"01",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",
		X"03",X"00",X"03",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",
		X"01",X"00",X"02",X"00",X"04",X"00",X"02",X"00",X"03",X"00",X"02",X"00",X"02",X"00",X"02",X"00",
		X"04",X"00",X"03",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"00",X"00",
		X"02",X"00",X"02",X"00",X"01",X"00",X"03",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"02",X"00",
		X"02",X"00",X"02",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"01",X"00",X"03",X"00",X"02",X"00",
		X"01",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",
		X"01",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"02",X"00",
		X"03",X"00",X"02",X"00",X"03",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",
		X"02",X"00",X"01",X"00",X"02",X"00",X"04",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"01",X"00",
		X"02",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"03",X"00",X"02",X"00",X"02",X"00",X"02",X"00",
		X"02",X"00",X"02",X"00",X"02",X"00",X"03",X"00",X"02",X"00",X"02",X"00",X"03",X"00",X"02",X"00",
		X"02",X"00",X"03",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"02",X"00",
		X"03",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"03",X"00",X"02",X"00",X"02",X"00",
		X"02",X"00",X"01",X"00",X"03",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"02",X"00",
		X"02",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"01",X"00",
		X"01",X"00",X"03",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",
		X"03",X"00",X"02",X"00",X"03",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"03",X"00",X"02",X"00",
		X"01",X"00",X"03",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"02",X"00",
		X"03",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"02",X"00",
		X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"03",X"00",X"01",X"00",X"02",X"00",X"02",X"00",
		X"02",X"00",X"03",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"02",X"00",
		X"01",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",
		X"02",X"00",X"01",X"00",X"01",X"00",X"03",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"02",X"00",
		X"03",X"00",X"02",X"00",X"04",X"00",X"02",X"00",X"02",X"00",X"03",X"00",X"03",X"00",X"03",X"00",
		X"02",X"00",X"03",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"04",X"00",X"02",X"00",X"03",X"00",
		X"02",X"00",X"03",X"00",X"01",X"00",X"03",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"02",X"00",
		X"01",X"00",X"02",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"02",X"00",X"02",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"02",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"02",X"00",X"01",X"00",
		X"02",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"02",X"00",
		X"00",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"02",X"00",
		X"02",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"02",X"00",X"03",X"00",X"00",X"00",X"FF",X"FF",
		X"02",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"02",X"00",
		X"01",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"01",X"00",X"01",X"00",
		X"02",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"02",X"00",
		X"02",X"00",X"01",X"00",X"01",X"00",X"03",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"02",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"02",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"02",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"02",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"02",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"01",X"00",
		X"02",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"02",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"02",X"00",X"00",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"03",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"01",X"00",
		X"02",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"02",X"00",X"01",X"00",
		X"02",X"00",X"02",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"01",X"00",
		X"00",X"00",X"02",X"00",X"02",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"02",X"00",X"01",X"00",
		X"02",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"02",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"01",X"00",
		X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"02",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"03",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"02",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"FF",X"FF",X"02",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"02",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"01",X"00",X"02",X"00",
		X"02",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"01",X"00",
		X"01",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"02",X"00",
		X"01",X"00",X"02",X"00",X"01",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"02",X"00",
		X"01",X"00",X"03",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"02",X"00",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"02",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"03",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"02",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"02",X"00",
		X"02",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"03",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"03",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"02",X"00",
		X"00",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"02",X"00",
		X"02",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"02",X"00",X"01",X"00",
		X"01",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"00",X"00",X"02",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",
		X"00",X"00",X"02",X"00",X"03",X"00",X"02",X"00",X"01",X"00",X"03",X"00",X"02",X"00",X"01",X"00",
		X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"03",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"00",X"00",
		X"02",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"03",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"02",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"02",X"00",
		X"00",X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"02",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"02",X"00",
		X"02",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"02",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"01",X"00",
		X"01",X"00",X"02",X"00",X"01",X"00",X"03",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"02",X"00",
		X"01",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"02",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"02",X"00",
		X"01",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"03",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"02",X"00",
		X"00",X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"02",X"00",
		X"01",X"00",X"03",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"01",X"00",X"02",X"00",X"02",X"00",
		X"00",X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"00",X"00",
		X"02",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"02",X"00",
		X"02",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"02",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"02",X"00",X"00",X"00",
		X"01",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"03",X"00",X"02",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"03",X"00",X"01",X"00",X"FF",X"FF",X"02",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"02",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"02",X"00",X"02",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"02",X"00",X"02",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"02",X"00",X"01",X"00",
		X"02",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"03",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"03",X"00",X"02",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"02",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"02",X"00",X"02",X"00",
		X"02",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"02",X"00",
		X"02",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"02",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"02",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"03",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"02",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"00",X"00",
		X"00",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"03",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"00",X"00",
		X"02",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"02",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"02",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"03",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"02",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"02",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"03",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"02",X"00",
		X"02",X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"01",X"00",
		X"02",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"02",X"00",
		X"01",X"00",X"03",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FE",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"FE",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FE",X"FF",
		X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",X"02",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FE",X"FF",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"FE",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"FE",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"02",X"00",X"00",X"00",
		X"00",X"00",X"02",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FE",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",
		X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FE",X"FF",
		X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"02",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"02",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"02",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"02",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"02",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FE",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FE",X"FF",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"02",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"FF",X"FF",X"01",X"00",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"02",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"01",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FE",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"02",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"02",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"02",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"FE",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",
		X"01",X"00",X"FE",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"02",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FE",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FE",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",X"FE",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"02",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"02",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FE",X"FF",
		X"00",X"00",X"01",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"FE",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"02",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FE",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FE",X"FF",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"02",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"FE",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FE",X"FF",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"01",X"00",X"FF",X"FF",
		X"01",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FE",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FE",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"FE",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"FE",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"02",X"00",
		X"01",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"01",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"02",X"00",
		X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FE",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"FE",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FE",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"02",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"02",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"FE",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FE",X"FF",X"01",X"00",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FE",X"FF",X"01",X"00",X"FE",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"FE",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FE",X"FF",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",
		X"01",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FE",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"02",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FF",X"FF",X"FF",X"01",X"00",X"02",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"02",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"FE",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FE",X"FF",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FE",X"FF",X"00",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"01",X"00",X"FE",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"02",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FE",X"FF",X"01",X"00",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",
		X"02",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"01",X"00",X"02",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"02",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FE",X"FF",X"01",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"02",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"FE",X"FF",X"00",X"00",
		X"00",X"00",X"FE",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"02",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"02",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"01",X"00",X"02",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"02",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"00",X"00",X"FE",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"FF",X"FF",X"01",X"00",X"02",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"02",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"02",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"FE",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FE",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"02",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FE",X"FF",X"FE",X"FF",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"FE",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"FE",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"02",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"FE",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",
		X"FE",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"FE",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FE",X"FF",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"FE",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"FE",X"FF",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"01",X"00",X"FF",X"FF",X"02",X"00",X"FF",X"FF",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"FE",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"02",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",
		X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FE",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"02",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FE",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FE",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",X"02",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"02",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FE",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"FE",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"FE",X"FF",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FE",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"FE",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",
		X"FE",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"02",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"02",X"00",X"00",X"00",
		X"00",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FE",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FE",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"FE",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"02",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"00",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"02",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"02",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FE",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"FE",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"02",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"00",X"FF",X"FF",X"00",X"00",X"02",X"00",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"FE",X"FF",X"FE",X"FF",X"01",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"FE",X"FF",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"00",X"00",X"02",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",
		X"FE",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FE",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"02",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FE",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"02",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FE",X"FF",X"FF",X"FF",X"FE",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"02",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"02",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FE",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"01",X"00",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FE",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FE",X"FF",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FE",X"FF",X"00",X"00",X"FE",X"FF",X"FF",X"FF",
		X"02",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"FE",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FE",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FE",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FE",X"FF",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"FE",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"02",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FE",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FF",X"FE",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"FF",X"FF",X"01",X"00",X"FE",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FE",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FE",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"02",X"00",
		X"02",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"02",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",
		X"02",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FE",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"02",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"02",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FE",X"FF",
		X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"01",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"02",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"00",
		X"01",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"02",X"00",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"FF",X"FF",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"02",X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"FF",X"FF",
		X"FE",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"FE",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"00",
		X"02",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"02",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"FE",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"FE",X"FF",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"02",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"02",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"02",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FE",X"FF",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",
		X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"02",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FE",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"02",X"00",X"00",X"00",X"FF",X"FF",X"FE",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"FE",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"FE",X"FF",X"FE",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"02",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FE",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"02",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"02",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"FE",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"FE",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"02",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"02",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"02",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"01",X"00",X"FE",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"01",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FE",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FE",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"02",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"02",X"00",X"01",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"02",X"00",
		X"FF",X"FF",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"02",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FE",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FE",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"01",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"02",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"02",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"02",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"02",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"02",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"FE",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FE",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",
		X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"02",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FE",X"FF",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FE",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FE",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FE",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FE",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"02",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"02",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"02",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"FE",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FE",X"FF",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"02",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",X"01",X"00",X"01",X"00",
		X"02",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"02",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"01",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FE",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"01",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"FE",X"FF",X"01",X"00",X"FF",X"FF",X"02",X"00",X"00",X"00",X"02",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"02",X"00",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FE",X"FF",X"01",X"00",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"02",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FE",X"FF",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FE",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FE",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"02",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"02",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FE",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"02",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"02",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FE",X"FF",X"FF",X"FF",
		X"FE",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FE",X"FF",
		X"00",X"00",X"FE",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FE",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"FE",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"FE",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FE",X"FF",X"00",X"00",X"FE",X"FF",X"FF",X"FF",X"01",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",X"FE",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",X"FF",X"FF",
		X"00",X"00",X"02",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"01",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"01",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FE",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FE",X"FF",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"02",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"01",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FE",X"FF",X"01",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FE",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"02",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FE",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",
		X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FE",X"FF",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"FE",X"FF",X"00",X"00",X"FF",X"FF",X"FE",X"FF",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FE",X"FF",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"FE",X"FF",X"FE",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"02",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"01",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"FE",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"00",X"00",
		X"02",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",X"01",X"00",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"02",X"00",X"FF",X"FF",X"00",X"00",X"02",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"FF",X"FF",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"B0",X"FB",X"FF",X"05",X"00",
		X"F6",X"FF",X"0B",X"00",X"F2",X"FF",X"12",X"00",X"E9",X"FF",X"1F",X"00",X"D7",X"FF",X"3C",X"00",
		X"A3",X"FF",X"A7",X"00",X"04",X"F6",X"FC",X"F1",X"E0",X"F2",X"B1",X"F1",X"EB",X"F1",X"16",X"F1",
		X"24",X"F1",X"75",X"F0",X"73",X"F0",X"DD",X"EF",X"D1",X"EF",X"4B",X"EF",X"3B",X"EF",X"C2",X"EE",
		X"B0",X"EE",X"42",X"EE",X"2F",X"EE",X"C9",X"ED",X"B7",X"ED",X"5A",X"ED",X"46",X"ED",X"F1",X"EC",
		X"DE",X"EC",X"90",X"EC",X"7E",X"EC",X"36",X"EC",X"25",X"EC",X"E4",X"EB",X"D1",X"EB",X"97",X"EB",
		X"85",X"EB",X"4F",X"EB",X"4A",X"EB",X"64",X"EB",X"CB",X"EB",X"34",X"EC",X"CA",X"EC",X"54",X"ED",
		X"FA",X"ED",X"91",X"EE",X"3A",X"EF",X"D1",X"EF",X"75",X"F0",X"09",X"F1",X"A6",X"F1",X"35",X"F2",
		X"C9",X"F2",X"52",X"F3",X"DD",X"F3",X"60",X"F4",X"E3",X"F4",X"5F",X"F5",X"DB",X"F5",X"51",X"F6",
		X"C3",X"F6",X"34",X"F7",X"A0",X"F7",X"0B",X"F8",X"6F",X"F8",X"D6",X"F8",X"10",X"F9",X"0C",X"F9",
		X"E4",X"F8",X"A0",X"F8",X"4A",X"F8",X"EB",X"F7",X"83",X"F7",X"1C",X"F7",X"B0",X"F6",X"48",X"F6",
		X"DD",X"F5",X"77",X"F5",X"10",X"F5",X"B2",X"F4",X"4F",X"F4",X"F4",X"F3",X"98",X"F3",X"44",X"F3",
		X"ED",X"F2",X"9C",X"F2",X"4C",X"F2",X"01",X"F2",X"B5",X"F1",X"70",X"F1",X"27",X"F1",X"E8",X"F0",
		X"A3",X"F0",X"6F",X"F0",X"74",X"F0",X"AE",X"F0",X"06",X"F1",X"75",X"F1",X"F0",X"F1",X"74",X"F2",
		X"FB",X"F2",X"86",X"F3",X"0D",X"F4",X"97",X"F4",X"1A",X"F5",X"9E",X"F5",X"1D",X"F6",X"9C",X"F6",
		X"15",X"F7",X"8D",X"F7",X"FF",X"F7",X"71",X"F8",X"DD",X"F8",X"47",X"F9",X"AE",X"F9",X"13",X"FA",
		X"74",X"FA",X"D2",X"FA",X"2E",X"FB",X"86",X"FB",X"DE",X"FB",X"17",X"FC",X"0B",X"FC",X"DB",X"FB",
		X"8C",X"FB",X"2C",X"FB",X"C2",X"FA",X"50",X"FA",X"DB",X"F9",X"68",X"F9",X"F3",X"F8",X"80",X"F8",
		X"0E",X"F8",X"9F",X"F7",X"34",X"F7",X"CB",X"F6",X"64",X"F6",X"01",X"F6",X"A1",X"F5",X"44",X"F5",
		X"EA",X"F4",X"93",X"F4",X"3F",X"F4",X"ED",X"F3",X"9B",X"F3",X"51",X"F3",X"07",X"F3",X"BE",X"F2",
		X"7E",X"F2",X"75",X"F2",X"A3",X"F2",X"F2",X"F2",X"58",X"F3",X"CC",X"F3",X"49",X"F4",X"CC",X"F4",
		X"50",X"F5",X"D3",X"F5",X"58",X"F6",X"D7",X"F6",X"56",X"F7",X"D2",X"F7",X"4A",X"F8",X"C1",X"F8",
		X"35",X"F9",X"A4",X"F9",X"10",X"FA",X"79",X"FA",X"E0",X"FA",X"44",X"FB",X"A4",X"FB",X"02",X"FC",
		X"5E",X"FC",X"B6",X"FC",X"0C",X"FD",X"5E",X"FD",X"7B",X"FD",X"60",X"FD",X"22",X"FD",X"CA",X"FC",
		X"64",X"FC",X"F4",X"FB",X"80",X"FB",X"0A",X"FB",X"93",X"FA",X"1C",X"FA",X"A8",X"F9",X"36",X"F9",
		X"C6",X"F8",X"5A",X"F8",X"F1",X"F7",X"8B",X"F7",X"25",X"F7",X"C4",X"F6",X"68",X"F6",X"0E",X"F6",
		X"B5",X"F5",X"60",X"F5",X"0E",X"F5",X"BF",X"F4",X"72",X"F4",X"26",X"F4",X"DF",X"F3",X"99",X"F3",
		X"55",X"F3",X"13",X"F3",X"D6",X"F2",X"98",X"F2",X"5E",X"F2",X"25",X"F2",X"EE",X"F1",X"B9",X"F1",
		X"86",X"F1",X"55",X"F1",X"26",X"F1",X"F7",X"F0",X"CB",X"F0",X"A0",X"F0",X"78",X"F0",X"50",X"F0",
		X"2B",X"F0",X"06",X"F0",X"E3",X"EF",X"C2",X"EF",X"A0",X"EF",X"81",X"EF",X"63",X"EF",X"46",X"EF",
		X"2B",X"EF",X"10",X"EF",X"F7",X"EE",X"0A",X"EF",X"58",X"EF",X"C7",X"EF",X"54",X"F0",X"EA",X"F0",
		X"8C",X"F1",X"30",X"F2",X"D8",X"F2",X"7E",X"F3",X"23",X"F4",X"C3",X"F4",X"64",X"F5",X"FD",X"F5",
		X"94",X"F6",X"28",X"F7",X"B6",X"F7",X"44",X"F8",X"CB",X"F8",X"4E",X"F9",X"CE",X"F9",X"4B",X"FA",
		X"C3",X"FA",X"39",X"FB",X"AA",X"FB",X"18",X"FC",X"83",X"FC",X"ED",X"FC",X"51",X"FD",X"B3",X"FD",
		X"12",X"FE",X"6F",X"FE",X"C8",X"FE",X"21",X"FF",X"74",X"FF",X"C7",X"FF",X"15",X"00",X"62",X"00",
		X"AD",X"00",X"F5",X"00",X"3B",X"01",X"7F",X"01",X"C2",X"01",X"02",X"02",X"41",X"02",X"7E",X"02",
		X"B8",X"02",X"F1",X"02",X"27",X"03",X"5D",X"03",X"91",X"03",X"C2",X"03",X"F1",X"03",X"23",X"04",
		X"4F",X"04",X"7C",X"04",X"85",X"04",X"4F",X"04",X"F4",X"03",X"7C",X"03",X"F8",X"02",X"67",X"02",
		X"D2",X"01",X"3D",X"01",X"A7",X"00",X"13",X"00",X"81",X"FF",X"F2",X"FE",X"66",X"FE",X"DD",X"FD",
		X"57",X"FD",X"D6",X"FC",X"58",X"FC",X"DE",X"FB",X"6A",X"FB",X"F6",X"FA",X"86",X"FA",X"1A",X"FA",
		X"B4",X"F9",X"4C",X"F9",X"EC",X"F8",X"8D",X"F8",X"30",X"F8",X"DE",X"F7",X"C6",X"F7",X"E5",X"F7",
		X"24",X"F8",X"7B",X"F8",X"DD",X"F8",X"4D",X"F9",X"BC",X"F9",X"2E",X"FA",X"A4",X"FA",X"18",X"FB",
		X"88",X"FB",X"F9",X"FB",X"66",X"FC",X"D0",X"FC",X"38",X"FD",X"9E",X"FD",X"00",X"FE",X"60",X"FE",
		X"BD",X"FE",X"17",X"FF",X"6E",X"FF",X"C3",X"FF",X"14",X"00",X"65",X"00",X"B2",X"00",X"FE",X"00",
		X"48",X"01",X"8E",X"01",X"D3",X"01",X"16",X"02",X"57",X"02",X"96",X"02",X"D2",X"02",X"0E",X"03",
		X"46",X"03",X"7D",X"03",X"B3",X"03",X"E7",X"03",X"1A",X"04",X"4A",X"04",X"7B",X"04",X"A8",X"04",
		X"D5",X"04",X"FF",X"04",X"29",X"05",X"51",X"05",X"79",X"05",X"9E",X"05",X"C4",X"05",X"E6",X"05",
		X"08",X"06",X"2A",X"06",X"4B",X"06",X"68",X"06",X"87",X"06",X"A3",X"06",X"C0",X"06",X"DA",X"06",
		X"F4",X"06",X"0D",X"07",X"27",X"07",X"3E",X"07",X"55",X"07",X"66",X"07",X"63",X"07",X"5E",X"07",
		X"5A",X"07",X"57",X"07",X"53",X"07",X"4F",X"07",X"4B",X"07",X"46",X"07",X"43",X"07",X"40",X"07",
		X"3C",X"07",X"39",X"07",X"33",X"07",X"30",X"07",X"2B",X"07",X"29",X"07",X"25",X"07",X"22",X"07",
		X"1C",X"07",X"1A",X"07",X"14",X"07",X"13",X"07",X"A2",X"06",X"F1",X"05",X"46",X"05",X"94",X"04",
		X"E5",X"03",X"34",X"03",X"8A",X"02",X"E2",X"01",X"3D",X"01",X"9D",X"00",X"02",X"00",X"6B",X"FF",
		X"D8",X"FE",X"49",X"FE",X"BD",X"FD",X"38",X"FD",X"B5",X"FC",X"35",X"FC",X"BB",X"FB",X"43",X"FB",
		X"D2",X"FA",X"60",X"FA",X"F7",X"F9",X"8D",X"F9",X"57",X"F9",X"5C",X"F9",X"86",X"F9",X"CA",X"F9",
		X"1D",X"FA",X"7D",X"FA",X"DF",X"FA",X"47",X"FB",X"AE",X"FB",X"17",X"FC",X"7E",X"FC",X"E3",X"FC",
		X"46",X"FD",X"A9",X"FD",X"06",X"FE",X"63",X"FE",X"BD",X"FE",X"14",X"FF",X"69",X"FF",X"BB",X"FF",
		X"0A",X"00",X"5A",X"00",X"A4",X"00",X"EC",X"00",X"33",X"01",X"78",X"01",X"BA",X"01",X"FD",X"01",
		X"39",X"02",X"77",X"02",X"B3",X"02",X"EB",X"02",X"23",X"03",X"59",X"03",X"8D",X"03",X"BE",X"03",
		X"F0",X"03",X"1F",X"04",X"4B",X"04",X"7A",X"04",X"A5",X"04",X"CE",X"04",X"F5",X"04",X"1E",X"05",
		X"42",X"05",X"68",X"05",X"8B",X"05",X"AE",X"05",X"CF",X"05",X"F1",X"05",X"0E",X"06",X"2C",X"06",
		X"49",X"06",X"65",X"06",X"80",X"06",X"9A",X"06",X"B4",X"06",X"CD",X"06",X"E4",X"06",X"FB",X"06",
		X"0C",X"07",X"0B",X"07",X"06",X"07",X"02",X"07",X"FE",X"06",X"FC",X"06",X"F7",X"06",X"F4",X"06",
		X"EF",X"06",X"EB",X"06",X"E9",X"06",X"E5",X"06",X"E0",X"06",X"DE",X"06",X"DA",X"06",X"D6",X"06",
		X"D0",X"06",X"CF",X"06",X"CA",X"06",X"C8",X"06",X"C3",X"06",X"C1",X"06",X"BB",X"06",X"BA",X"06",
		X"B4",X"06",X"B6",X"06",X"8C",X"06",X"E5",X"05",X"36",X"05",X"84",X"04",X"D3",X"03",X"22",X"03",
		X"76",X"02",X"CB",X"01",X"25",X"01",X"83",X"00",X"E5",X"FF",X"4D",X"FF",X"B8",X"FE",X"27",X"FE",
		X"9B",X"FD",X"12",X"FD",X"8E",X"FC",X"0D",X"FC",X"90",X"FB",X"19",X"FB",X"A3",X"FA",X"33",X"FA",
		X"C4",X"F9",X"5A",X"F9",X"F4",X"F8",X"8F",X"F8",X"2F",X"F8",X"D2",X"F7",X"76",X"F7",X"20",X"F7",
		X"CB",X"F6",X"78",X"F6",X"2A",X"F6",X"DC",X"F5",X"92",X"F5",X"4A",X"F5",X"03",X"F5",X"C0",X"F4",
		X"81",X"F4",X"42",X"F4",X"03",X"F4",X"C9",X"F3",X"8F",X"F3",X"59",X"F3",X"25",X"F3",X"F1",X"F2",
		X"BF",X"F2",X"91",X"F2",X"62",X"F2",X"37",X"F2",X"0B",X"F2",X"E4",X"F1",X"BB",X"F1",X"94",X"F1",
		X"6F",X"F1",X"4D",X"F1",X"2A",X"F1",X"09",X"F1",X"E9",X"F0",X"CB",X"F0",X"AF",X"F0",X"92",X"F0",
		X"77",X"F0",X"5E",X"F0",X"46",X"F0",X"2E",X"F0",X"17",X"F0",X"01",X"F0",X"EE",X"EF",X"D9",X"EF",
		X"C6",X"EF",X"B4",X"EF",X"A2",X"EF",X"93",X"EF",X"82",X"EF",X"76",X"EF",X"66",X"EF",X"5A",X"EF",
		X"4A",X"EF",X"56",X"EF",X"A2",X"EF",X"13",X"F0",X"A3",X"F0",X"42",X"F1",X"ED",X"F1",X"9B",X"F2",
		X"4D",X"F3",X"FE",X"F3",X"AB",X"F4",X"58",X"F5",X"00",X"F6",X"A4",X"F6",X"46",X"F7",X"E2",X"F7",
		X"7A",X"F8",X"0F",X"F9",X"9F",X"F9",X"2B",X"FA",X"B3",X"FA",X"38",X"FB",X"B7",X"FB",X"33",X"FC",
		X"AE",X"FC",X"21",X"FD",X"96",X"FD",X"03",X"FE",X"6E",X"FE",X"A3",X"FE",X"9D",X"FE",X"75",X"FE",
		X"33",X"FE",X"E2",X"FD",X"86",X"FD",X"24",X"FD",X"C0",X"FC",X"5C",X"FC",X"F7",X"FB",X"96",X"FB",
		X"32",X"FB",X"D2",X"FA",X"77",X"FA",X"1A",X"FA",X"C3",X"F9",X"6D",X"F9",X"19",X"F9",X"C8",X"F8",
		X"7C",X"F8",X"30",X"F8",X"E5",X"F7",X"9F",X"F7",X"59",X"F7",X"18",X"F7",X"D6",X"F6",X"99",X"F6",
		X"5F",X"F6",X"22",X"F6",X"EB",X"F5",X"B4",X"F5",X"80",X"F5",X"4D",X"F5",X"1D",X"F5",X"ED",X"F4",
		X"BF",X"F4",X"94",X"F4",X"68",X"F4",X"41",X"F4",X"18",X"F4",X"F3",X"F3",X"CE",X"F3",X"AB",X"F3",
		X"89",X"F3",X"67",X"F3",X"47",X"F3",X"29",X"F3",X"0D",X"F3",X"F1",X"F2",X"D5",X"F2",X"BB",X"F2",
		X"A2",X"F2",X"8A",X"F2",X"73",X"F2",X"5D",X"F2",X"48",X"F2",X"33",X"F2",X"20",X"F2",X"0D",X"F2",
		X"FE",X"F1",X"EB",X"F1",X"DC",X"F1",X"CD",X"F1",X"BE",X"F1",X"B0",X"F1",X"A3",X"F1",X"97",X"F1",
		X"8B",X"F1",X"7F",X"F1",X"76",X"F1",X"6B",X"F1",X"60",X"F1",X"58",X"F1",X"50",X"F1",X"48",X"F1",
		X"41",X"F1",X"3B",X"F1",X"33",X"F1",X"2F",X"F1",X"27",X"F1",X"25",X"F1",X"1E",X"F1",X"40",X"F1",
		X"9C",X"F1",X"1D",X"F2",X"B8",X"F2",X"5F",X"F3",X"13",X"F4",X"C7",X"F4",X"7D",X"F5",X"33",X"F6",
		X"E7",X"F6",X"98",X"F7",X"46",X"F8",X"EE",X"F8",X"94",X"F9",X"34",X"FA",X"D1",X"FA",X"69",X"FB",
		X"FD",X"FB",X"8B",X"FC",X"17",X"FD",X"9D",X"FD",X"20",X"FE",X"A0",X"FE",X"1C",X"FF",X"94",X"FF",
		X"07",X"00",X"78",X"00",X"DE",X"00",X"08",X"01",X"FC",X"00",X"CF",X"00",X"8C",X"00",X"3A",X"00",
		X"E1",X"FF",X"81",X"FF",X"1E",X"FF",X"BC",X"FE",X"59",X"FE",X"F8",X"FD",X"98",X"FD",X"3B",X"FD",
		X"E0",X"FC",X"87",X"FC",X"30",X"FC",X"DB",X"FB",X"89",X"FB",X"3B",X"FB",X"ED",X"FA",X"A3",X"FA",
		X"5B",X"FA",X"16",X"FA",X"D4",X"F9",X"93",X"F9",X"53",X"F9",X"16",X"F9",X"DB",X"F8",X"A1",X"F8",
		X"6A",X"F8",X"35",X"F8",X"01",X"F8",X"CE",X"F7",X"9E",X"F7",X"6D",X"F7",X"41",X"F7",X"17",X"F7",
		X"EC",X"F6",X"C4",X"F6",X"9D",X"F6",X"77",X"F6",X"52",X"F6",X"2F",X"F6",X"0D",X"F6",X"EC",X"F5",
		X"CC",X"F5",X"AF",X"F5",X"92",X"F5",X"75",X"F5",X"59",X"F5",X"3E",X"F5",X"25",X"F5",X"0E",X"F5",
		X"F6",X"F4",X"E4",X"F4",X"07",X"F5",X"61",X"F5",X"D9",X"F5",X"69",X"F6",X"05",X"F7",X"AA",X"F7",
		X"52",X"F8",X"FA",X"F8",X"A0",X"F9",X"46",X"FA",X"EA",X"FA",X"87",X"FB",X"23",X"FC",X"BA",X"FC",
		X"4C",X"FD",X"DC",X"FD",X"67",X"FE",X"EF",X"FE",X"72",X"FF",X"F0",X"FF",X"6C",X"00",X"E4",X"00",
		X"57",X"01",X"C9",X"01",X"36",X"02",X"A0",X"02",X"07",X"03",X"6B",X"03",X"CC",X"03",X"2A",X"04",
		X"84",X"04",X"DE",X"04",X"33",X"05",X"85",X"05",X"D6",X"05",X"25",X"06",X"71",X"06",X"B8",X"06",
		X"01",X"07",X"45",X"07",X"87",X"07",X"C7",X"07",X"05",X"08",X"43",X"08",X"7C",X"08",X"B5",X"08",
		X"EC",X"08",X"20",X"09",X"53",X"09",X"86",X"09",X"B6",X"09",X"E3",X"09",X"11",X"0A",X"3B",X"0A",
		X"65",X"0A",X"5D",X"0A",X"1B",X"0A",X"B8",X"09",X"3B",X"09",X"B1",X"08",X"20",X"08",X"87",X"07",
		X"EF",X"06",X"57",X"06",X"C0",X"05",X"2B",X"05",X"9B",X"04",X"0B",X"04",X"83",X"03",X"FD",X"02",
		X"78",X"02",X"FA",X"01",X"7F",X"01",X"07",X"01",X"91",X"00",X"23",X"00",X"B4",X"FF",X"4C",X"FF",
		X"E4",X"FE",X"80",X"FE",X"20",X"FE",X"C2",X"FD",X"67",X"FD",X"0D",X"FD",X"B8",X"FC",X"67",X"FC",
		X"17",X"FC",X"C8",X"FB",X"7E",X"FB",X"35",X"FB",X"EE",X"FA",X"AA",X"FA",X"67",X"FA",X"28",X"FA",
		X"E9",X"F9",X"AC",X"F9",X"74",X"F9",X"3A",X"F9",X"05",X"F9",X"CF",X"F8",X"9D",X"F8",X"6D",X"F8",
		X"3C",X"F8",X"0F",X"F8",X"E1",X"F7",X"B8",X"F7",X"8F",X"F7",X"66",X"F7",X"3F",X"F7",X"1B",X"F7",
		X"1E",X"F7",X"5F",X"F7",X"C3",X"F7",X"43",X"F8",X"CE",X"F8",X"66",X"F9",X"00",X"FA",X"9B",X"FA",
		X"39",X"FB",X"D4",X"FB",X"6B",X"FC",X"00",X"FD",X"91",X"FD",X"20",X"FE",X"AA",X"FE",X"31",X"FF",
		X"B4",X"FF",X"33",X"00",X"AE",X"00",X"26",X"01",X"9A",X"01",X"0A",X"02",X"79",X"02",X"E2",X"02",
		X"4A",X"03",X"AC",X"03",X"0F",X"04",X"63",X"04",X"7C",X"04",X"5E",X"04",X"20",X"04",X"CF",X"03",
		X"6E",X"03",X"06",X"03",X"99",X"02",X"2B",X"02",X"BC",X"01",X"4D",X"01",X"E1",X"00",X"75",X"00",
		X"0E",X"00",X"A9",X"FF",X"45",X"FF",X"E5",X"FE",X"87",X"FE",X"2B",X"FE",X"D4",X"FD",X"7E",X"FD",
		X"2C",X"FD",X"DA",X"FC",X"8C",X"FC",X"41",X"FC",X"F7",X"FB",X"B0",X"FB",X"6B",X"FB",X"2A",X"FB",
		X"EA",X"FA",X"AC",X"FA",X"6F",X"FA",X"35",X"FA",X"FB",X"F9",X"C6",X"F9",X"91",X"F9",X"5E",X"F9",
		X"2B",X"F9",X"FB",X"F8",X"CD",X"F8",X"A1",X"F8",X"76",X"F8",X"4D",X"F8",X"24",X"F8",X"FB",X"F7",
		X"D8",X"F7",X"B3",X"F7",X"8F",X"F7",X"6E",X"F7",X"4D",X"F7",X"2E",X"F7",X"0F",X"F7",X"F3",X"F6",
		X"D6",X"F6",X"BC",X"F6",X"A1",X"F6",X"88",X"F6",X"71",X"F6",X"58",X"F6",X"41",X"F6",X"2E",X"F6",
		X"17",X"F6",X"04",X"F6",X"F1",X"F5",X"DD",X"F5",X"CD",X"F5",X"BC",X"F5",X"AD",X"F5",X"9E",X"F5",
		X"8E",X"F5",X"81",X"F5",X"74",X"F5",X"66",X"F5",X"5A",X"F5",X"4D",X"F5",X"44",X"F5",X"39",X"F5",
		X"30",X"F5",X"26",X"F5",X"1D",X"F5",X"14",X"F5",X"0C",X"F5",X"05",X"F5",X"FF",X"F4",X"F7",X"F4",
		X"F2",X"F4",X"EC",X"F4",X"E6",X"F4",X"E3",X"F4",X"DE",X"F4",X"D8",X"F4",X"D4",X"F4",X"D1",X"F4",
		X"CF",X"F4",X"CC",X"F4",X"C7",X"F4",X"C6",X"F4",X"C5",X"F4",X"C3",X"F4",X"C2",X"F4",X"C1",X"F4",
		X"BF",X"F4",X"BF",X"F4",X"BF",X"F4",X"BF",X"F4",X"C0",X"F4",X"BF",X"F4",X"C0",X"F4",X"C1",X"F4",
		X"C2",X"F4",X"C5",X"F4",X"FA",X"F4",X"68",X"F5",X"F6",X"F5",X"98",X"F6",X"48",X"F7",X"FF",X"F7",
		X"BA",X"F8",X"75",X"F9",X"2F",X"FA",X"E6",X"FA",X"9A",X"FB",X"48",X"FC",X"F4",X"FC",X"9A",X"FD",
		X"3C",X"FE",X"DA",X"FE",X"73",X"FF",X"08",X"00",X"97",X"00",X"24",X"01",X"AD",X"01",X"30",X"02",
		X"B0",X"02",X"2E",X"03",X"A5",X"03",X"1A",X"04",X"8B",X"04",X"F8",X"04",X"64",X"05",X"CB",X"05",
		X"31",X"06",X"92",X"06",X"EF",X"06",X"4A",X"07",X"A1",X"07",X"F8",X"07",X"4B",X"08",X"9B",X"08",
		X"E7",X"08",X"35",X"09",X"7D",X"09",X"C5",X"09",X"09",X"0A",X"4A",X"0A",X"8A",X"0A",X"C8",X"0A",
		X"03",X"0B",X"3E",X"0B",X"76",X"0B",X"AC",X"0B",X"E1",X"0B",X"15",X"0C",X"44",X"0C",X"75",X"0C",
		X"95",X"0C",X"78",X"0C",X"2B",X"0C",X"BF",X"0B",X"42",X"0B",X"B7",X"0A",X"27",X"0A",X"91",X"09",
		X"FB",X"08",X"67",X"08",X"D5",X"07",X"45",X"07",X"B7",X"06",X"2C",X"06",X"A8",X"05",X"24",X"05",
		X"A5",X"04",X"2A",X"04",X"B2",X"03",X"3D",X"03",X"CD",X"02",X"5E",X"02",X"F3",X"01",X"8D",X"01",
		X"28",X"01",X"C7",X"00",X"68",X"00",X"0E",X"00",X"B5",X"FF",X"5F",X"FF",X"0C",X"FF",X"BC",X"FE",
		X"6C",X"FE",X"22",X"FE",X"D9",X"FD",X"90",X"FD",X"4C",X"FD",X"09",X"FD",X"C8",X"FC",X"8A",X"FC",
		X"4E",X"FC",X"13",X"FC",X"D9",X"FB",X"A2",X"FB",X"6D",X"FB",X"39",X"FB",X"07",X"FB",X"D7",X"FA",
		X"A7",X"FA",X"7B",X"FA",X"4F",X"FA",X"25",X"FA",X"FB",X"F9",X"D2",X"F9",X"AC",X"F9",X"89",X"F9",
		X"64",X"F9",X"43",X"F9",X"21",X"F9",X"01",X"F9",X"E1",X"F8",X"C3",X"F8",X"A7",X"F8",X"8B",X"F8",
		X"71",X"F8",X"56",X"F8",X"3D",X"F8",X"27",X"F8",X"0E",X"F8",X"F8",X"F7",X"E2",X"F7",X"CE",X"F7",
		X"B9",X"F7",X"A7",X"F7",X"95",X"F7",X"85",X"F7",X"73",X"F7",X"63",X"F7",X"53",X"F7",X"44",X"F7",
		X"36",X"F7",X"2A",X"F7",X"1B",X"F7",X"0F",X"F7",X"04",X"F7",X"F9",X"F6",X"ED",X"F6",X"E3",X"F6",
		X"DA",X"F6",X"D0",X"F6",X"C8",X"F6",X"C1",X"F6",X"B8",X"F6",X"B1",X"F6",X"AA",X"F6",X"A3",X"F6",
		X"9C",X"F6",X"97",X"F6",X"92",X"F6",X"8C",X"F6",X"87",X"F6",X"84",X"F6",X"80",X"F6",X"7C",X"F6",
		X"78",X"F6",X"75",X"F6",X"72",X"F6",X"70",X"F6",X"6D",X"F6",X"6B",X"F6",X"6E",X"F6",X"A7",X"F6",
		X"14",X"F7",X"A1",X"F7",X"44",X"F8",X"F3",X"F8",X"A5",X"F9",X"5E",X"FA",X"17",X"FB",X"CC",X"FB",
		X"82",X"FC",X"32",X"FD",X"DF",X"FD",X"87",X"FE",X"2C",X"FF",X"CC",X"FF",X"66",X"00",X"FD",X"00",
		X"90",X"01",X"1D",X"02",X"A7",X"02",X"2D",X"03",X"AE",X"03",X"2E",X"04",X"A7",X"04",X"1D",X"05",
		X"90",X"05",X"00",X"06",X"56",X"06",X"6A",X"06",X"53",X"06",X"1C",X"06",X"D2",X"05",X"7C",X"05",
		X"1F",X"05",X"BD",X"04",X"58",X"04",X"F5",X"03",X"92",X"03",X"30",X"03",X"CF",X"02",X"71",X"02",
		X"16",X"02",X"BD",X"01",X"65",X"01",X"10",X"01",X"BD",X"00",X"6E",X"00",X"23",X"00",X"D8",X"FF",
		X"8F",X"FF",X"48",X"FF",X"03",X"FF",X"C1",X"FE",X"81",X"FE",X"45",X"FE",X"39",X"FE",X"69",X"FE",
		X"B9",X"FE",X"24",X"FF",X"9D",X"FF",X"1D",X"00",X"A4",X"00",X"2B",X"01",X"B4",X"01",X"39",X"02",
		X"BF",X"02",X"42",X"03",X"C1",X"03",X"3C",X"04",X"B4",X"04",X"2A",X"05",X"9B",X"05",X"0B",X"06",
		X"76",X"06",X"DE",X"06",X"42",X"07",X"A5",X"07",X"03",X"08",X"5F",X"08",X"B9",X"08",X"0E",X"09",
		X"61",X"09",X"B3",X"09",X"01",X"0A",X"4E",X"0A",X"96",X"0A",X"DF",X"0A",X"23",X"0B",X"66",X"0B",
		X"A5",X"0B",X"E4",X"0B",X"20",X"0C",X"5A",X"0C",X"94",X"0C",X"C9",X"0C",X"FC",X"0C",X"31",X"0D",
		X"60",X"0D",X"90",X"0D",X"BF",X"0D",X"EA",X"0D",X"15",X"0E",X"3F",X"0E",X"67",X"0E",X"8D",X"0E",
		X"B3",X"0E",X"D5",X"0E",X"F9",X"0E",X"18",X"0F",X"38",X"0F",X"2E",X"0F",X"E8",X"0E",X"7C",X"0E",
		X"F9",X"0D",X"67",X"0D",X"CC",X"0C",X"2C",X"0C",X"8B",X"0B",X"EB",X"0A",X"4D",X"0A",X"B0",X"09",
		X"17",X"09",X"81",X"08",X"EF",X"07",X"61",X"07",X"D6",X"06",X"4D",X"06",X"CD",X"05",X"4E",X"05",
		X"D2",X"04",X"5A",X"04",X"E6",X"03",X"75",X"03",X"07",X"03",X"9F",X"02",X"36",X"02",X"D2",X"01",
		X"7C",X"01",X"62",X"01",X"7F",X"01",X"B7",X"01",X"08",X"02",X"65",X"02",X"CC",X"02",X"35",X"03",
		X"A0",X"03",X"0E",X"04",X"79",X"04",X"E4",X"04",X"4B",X"05",X"B1",X"05",X"14",X"06",X"75",X"06",
		X"D3",X"06",X"2F",X"07",X"87",X"07",X"DE",X"07",X"31",X"08",X"82",X"08",X"CE",X"08",X"1B",X"09",
		X"66",X"09",X"AB",X"09",X"F0",X"09",X"33",X"0A",X"73",X"0A",X"B1",X"0A",X"EE",X"0A",X"28",X"0B",
		X"62",X"0B",X"97",X"0B",X"CC",X"0B",X"00",X"0C",X"30",X"0C",X"60",X"0C",X"8F",X"0C",X"BA",X"0C",
		X"E5",X"0C",X"0E",X"0D",X"38",X"0D",X"5D",X"0D",X"83",X"0D",X"A5",X"0D",X"C8",X"0D",X"EA",X"0D",
		X"0A",X"0E",X"2A",X"0E",X"47",X"0E",X"64",X"0E",X"7F",X"0E",X"9A",X"0E",X"B3",X"0E",X"CD",X"0E",
		X"E4",X"0E",X"FB",X"0E",X"10",X"0F",X"25",X"0F",X"38",X"0F",X"4C",X"0F",X"5E",X"0F",X"6C",X"0F",
		X"67",X"0F",X"5E",X"0F",X"56",X"0F",X"4D",X"0F",X"45",X"0F",X"3C",X"0F",X"35",X"0F",X"2C",X"0F",
		X"23",X"0F",X"1B",X"0F",X"13",X"0F",X"0A",X"0F",X"02",X"0F",X"FA",X"0E",X"F2",X"0E",X"EA",X"0E",
		X"E2",X"0E",X"D8",X"0E",X"D2",X"0E",X"C8",X"0E",X"C0",X"0E",X"B8",X"0E",X"AF",X"0E",X"A8",X"0E",
		X"A0",X"0E",X"97",X"0E",X"90",X"0E",X"87",X"0E",X"7E",X"0E",X"77",X"0E",X"6F",X"0E",X"68",X"0E",
		X"60",X"0E",X"57",X"0E",X"50",X"0E",X"47",X"0E",X"3F",X"0E",X"37",X"0E",X"2F",X"0E",X"29",X"0E",
		X"1F",X"0E",X"18",X"0E",X"10",X"0E",X"09",X"0E",X"00",X"0E",X"F9",X"0D",X"F1",X"0D",X"EA",X"0D",
		X"E1",X"0D",X"DB",X"0D",X"D1",X"0D",X"CA",X"0D",X"51",X"0D",X"8A",X"0C",X"D6",X"0B",X"16",X"0B",
		X"62",X"0A",X"AA",X"09",X"FC",X"08",X"4E",X"08",X"A8",X"07",X"03",X"07",X"64",X"06",X"CA",X"05",
		X"35",X"05",X"A3",X"04",X"17",X"04",X"8A",X"03",X"08",X"03",X"86",X"02",X"09",X"02",X"8E",X"01",
		X"1B",X"01",X"A4",X"00",X"4A",X"00",X"2D",X"00",X"42",X"00",X"73",X"00",X"BA",X"00",X"0B",X"01",
		X"66",X"01",X"C6",X"01",X"27",X"02",X"89",X"02",X"E8",X"02",X"49",X"03",X"A7",X"03",X"03",X"04",
		X"5B",X"04",X"B2",X"04",X"07",X"05",X"5A",X"05",X"AA",X"05",X"F7",X"05",X"43",X"06",X"8A",X"06",
		X"D1",X"06",X"16",X"07",X"58",X"07",X"99",X"07",X"D6",X"07",X"12",X"08",X"1E",X"08",X"F1",X"07",
		X"9D",X"07",X"33",X"07",X"BA",X"06",X"35",X"06",X"AD",X"05",X"23",X"05",X"9A",X"04",X"10",X"04",
		X"89",X"03",X"05",X"03",X"85",X"02",X"05",X"02",X"8A",X"01",X"12",X"01",X"9E",X"00",X"2D",X"00",
		X"C1",X"FF",X"57",X"FF",X"EF",X"FE",X"8C",X"FE",X"2C",X"FE",X"CD",X"FD",X"71",X"FD",X"19",X"FD",
		X"C3",X"FC",X"6F",X"FC",X"21",X"FC",X"D2",X"FB",X"88",X"FB",X"3E",X"FB",X"F7",X"FA",X"B1",X"FA",
		X"71",X"FA",X"30",X"FA",X"F2",X"F9",X"B4",X"F9",X"7C",X"F9",X"42",X"F9",X"0C",X"F9",X"D8",X"F8",
		X"A4",X"F8",X"73",X"F8",X"43",X"F8",X"16",X"F8",X"E9",X"F7",X"BD",X"F7",X"92",X"F7",X"6B",X"F7",
		X"45",X"F7",X"20",X"F7",X"FB",X"F6",X"D6",X"F6",X"BE",X"F6",X"E2",X"F6",X"36",X"F7",X"AA",X"F7",
		X"31",X"F8",X"C5",X"F8",X"61",X"F9",X"FE",X"F9",X"9F",X"FA",X"3A",X"FB",X"D7",X"FB",X"72",X"FC",
		X"07",X"FD",X"9B",X"FD",X"28",X"FE",X"B3",X"FE",X"39",X"FF",X"BD",X"FF",X"3A",X"00",X"B7",X"00",
		X"2E",X"01",X"A2",X"01",X"13",X"02",X"82",X"02",X"EB",X"02",X"53",X"03",X"B7",X"03",X"19",X"04",
		X"57",X"04",X"56",X"04",X"2B",X"04",X"E6",X"03",X"8E",X"03",X"2C",X"03",X"C2",X"02",X"55",X"02",
		X"E5",X"01",X"78",X"01",X"0B",X"01",X"9F",X"00",X"37",X"00",X"D2",X"FF",X"6C",X"FF",X"0C",X"FF",
		X"AC",X"FE",X"52",X"FE",X"F8",X"FD",X"A2",X"FD",X"4E",X"FD",X"FD",X"FC",X"AE",X"FC",X"61",X"FC",
		X"17",X"FC",X"CF",X"FB",X"89",X"FB",X"4C",X"FB",X"45",X"FB",X"77",X"FB",X"C6",X"FB",X"30",X"FC",
		X"A5",X"FC",X"22",X"FD",X"A5",X"FD",X"29",X"FE",X"AE",X"FE",X"2F",X"FF",X"B1",X"FF",X"2F",X"00",
		X"AA",X"00",X"22",X"01",X"97",X"01",X"09",X"02",X"79",X"02",X"E3",X"02",X"4D",X"03",X"B2",X"03",
		X"14",X"04",X"71",X"04",X"CF",X"04",X"2A",X"05",X"80",X"05",X"D3",X"05",X"26",X"06",X"5F",X"06",
		X"55",X"06",X"20",X"06",X"CF",X"05",X"6D",X"05",X"FE",X"04",X"88",X"04",X"0E",X"04",X"94",X"03",
		X"1A",X"03",X"A1",X"02",X"2B",X"02",X"B7",X"01",X"44",X"01",X"D6",X"00",X"6A",X"00",X"02",X"00",
		X"9D",X"FF",X"3A",X"FF",X"DB",X"FE",X"7F",X"FE",X"24",X"FE",X"CB",X"FD",X"77",X"FD",X"25",X"FD",
		X"D7",X"FC",X"88",X"FC",X"3F",X"FC",X"2B",X"FC",X"50",X"FC",X"95",X"FC",X"F4",X"FC",X"62",X"FD",
		X"DA",X"FD",X"56",X"FE",X"D5",X"FE",X"53",X"FF",X"D2",X"FF",X"4D",X"00",X"C6",X"00",X"3D",X"01",
		X"B1",X"01",X"21",X"02",X"91",X"02",X"FC",X"02",X"61",X"03",X"C7",X"03",X"2A",X"04",X"87",X"04",
		X"E3",X"04",X"3C",X"05",X"92",X"05",X"E6",X"05",X"37",X"06",X"86",X"06",X"D2",X"06",X"1A",X"07",
		X"62",X"07",X"A7",X"07",X"EA",X"07",X"2C",X"08",X"6A",X"08",X"A7",X"08",X"E1",X"08",X"1B",X"09",
		X"51",X"09",X"86",X"09",X"BA",X"09",X"EC",X"09",X"1C",X"0A",X"4A",X"0A",X"77",X"0A",X"A4",X"0A",
		X"CC",X"0A",X"F6",X"0A",X"1E",X"0B",X"44",X"0B",X"68",X"0B",X"8B",X"0B",X"AD",X"0B",X"CD",X"0B",
		X"ED",X"0B",X"0C",X"0C",X"29",X"0C",X"46",X"0C",X"61",X"0C",X"7B",X"0C",X"94",X"0C",X"AD",X"0C",
		X"C3",X"0C",X"DB",X"0C",X"F0",X"0C",X"04",X"0D",X"18",X"0D",X"2B",X"0D",X"39",X"0D",X"35",X"0D",
		X"2A",X"0D",X"24",X"0D",X"1E",X"0D",X"14",X"0D",X"0C",X"0D",X"07",X"0D",X"FF",X"0C",X"F8",X"0C",
		X"F0",X"0C",X"E9",X"0C",X"E2",X"0C",X"DB",X"0C",X"D2",X"0C",X"CB",X"0C",X"C5",X"0C",X"BE",X"0C",
		X"AC",X"0C",X"28",X"0C",X"7A",X"0B",X"CC",X"0A",X"19",X"0A",X"67",X"09",X"B6",X"08",X"08",X"08",
		X"5C",X"07",X"B7",X"06",X"13",X"06",X"75",X"05",X"DA",X"04",X"43",X"04",X"B1",X"03",X"23",X"03",
		X"99",X"02",X"13",X"02",X"92",X"01",X"14",X"01",X"9A",X"00",X"25",X"00",X"B3",X"FF",X"44",X"FF",
		X"D7",X"FE",X"6E",X"FE",X"09",X"FE",X"A6",X"FD",X"47",X"FD",X"EB",X"FC",X"90",X"FC",X"3B",X"FC",
		X"E5",X"FB",X"95",X"FB",X"46",X"FB",X"F9",X"FA",X"AF",X"FA",X"67",X"FA",X"21",X"FA",X"DE",X"F9",
		X"9D",X"F9",X"5F",X"F9",X"22",X"F9",X"E6",X"F8",X"AC",X"F8",X"76",X"F8",X"3F",X"F8",X"0D",X"F8",
		X"DC",X"F7",X"AA",X"F7",X"7C",X"F7",X"4E",X"F7",X"22",X"F7",X"F8",X"F6",X"CF",X"F6",X"A8",X"F6",
		X"83",X"F6",X"5F",X"F6",X"3C",X"F6",X"19",X"F6",X"F7",X"F5",X"D9",X"F5",X"BA",X"F5",X"9B",X"F5",
		X"80",X"F5",X"65",X"F5",X"4A",X"F5",X"31",X"F5",X"1A",X"F5",X"02",X"F5",X"EB",X"F4",X"D5",X"F4",
		X"C2",X"F4",X"AD",X"F4",X"99",X"F4",X"87",X"F4",X"76",X"F4",X"65",X"F4",X"56",X"F4",X"45",X"F4",
		X"38",X"F4",X"29",X"F4",X"1A",X"F4",X"0F",X"F4",X"03",X"F4",X"F8",X"F3",X"EE",X"F3",X"E3",X"F3",
		X"D8",X"F3",X"D0",X"F3",X"C7",X"F3",X"BF",X"F3",X"B7",X"F3",X"AE",X"F3",X"A9",X"F3",X"A2",X"F3",
		X"9D",X"F3",X"96",X"F3",X"92",X"F3",X"8D",X"F3",X"88",X"F3",X"83",X"F3",X"80",X"F3",X"7D",X"F3",
		X"7A",X"F3",X"77",X"F3",X"75",X"F3",X"72",X"F3",X"70",X"F3",X"71",X"F3",X"6E",X"F3",X"6E",X"F3",
		X"6D",X"F3",X"6D",X"F3",X"6D",X"F3",X"6E",X"F3",X"6D",X"F3",X"6D",X"F3",X"6E",X"F3",X"71",X"F3",
		X"70",X"F3",X"73",X"F3",X"74",X"F3",X"76",X"F3",X"78",X"F3",X"7B",X"F3",X"7C",X"F3",X"7F",X"F3",
		X"82",X"F3",X"87",X"F3",X"88",X"F3",X"8A",X"F3",X"8F",X"F3",X"93",X"F3",X"95",X"F3",X"AD",X"F3",
		X"03",X"F4",X"84",X"F4",X"1E",X"F5",X"CB",X"F5",X"83",X"F6",X"3C",X"F7",X"FA",X"F7",X"B7",X"F8",
		X"71",X"F9",X"28",X"FA",X"DB",X"FA",X"8A",X"FB",X"35",X"FC",X"DC",X"FC",X"7D",X"FD",X"1A",X"FE",
		X"B3",X"FE",X"47",X"FF",X"D8",X"FF",X"63",X"00",X"EA",X"00",X"6D",X"01",X"EE",X"01",X"69",X"02",
		X"E1",X"02",X"53",X"03",X"C5",X"03",X"04",X"04",X"06",X"04",X"E4",X"03",X"A7",X"03",X"5A",X"03",
		X"05",X"03",X"A6",X"02",X"47",X"02",X"E6",X"01",X"84",X"01",X"24",X"01",X"C4",X"00",X"67",X"00",
		X"0C",X"00",X"B5",X"FF",X"5E",X"FF",X"0A",X"FF",X"B7",X"FE",X"69",X"FE",X"1D",X"FE",X"D3",X"FD",
		X"8A",X"FD",X"43",X"FD",X"00",X"FD",X"BD",X"FC",X"80",X"FC",X"3F",X"FC",X"14",X"FC",X"24",X"FC",
		X"65",X"FC",X"C2",X"FC",X"35",X"FD",X"B5",X"FD",X"38",X"FE",X"C1",X"FE",X"4B",X"FF",X"D6",X"FF",
		X"5B",X"00",X"E1",X"00",X"62",X"01",X"E4",X"01",X"5E",X"02",X"D8",X"02",X"4C",X"03",X"BE",X"03",
		X"2C",X"04",X"9A",X"04",X"01",X"05",X"65",X"05",X"C6",X"05",X"26",X"06",X"82",X"06",X"DA",X"06",
		X"31",X"07",X"86",X"07",X"B0",X"07",X"9C",X"07",X"63",X"07",X"0E",X"07",X"AA",X"06",X"3B",X"06",
		X"C6",X"05",X"4F",X"05",X"D5",X"04",X"5E",X"04",X"E7",X"03",X"73",X"03",X"01",X"03",X"92",X"02",
		X"26",X"02",X"BC",X"01",X"55",X"01",X"F2",X"00",X"91",X"00",X"33",X"00",X"D9",X"FF",X"81",X"FF",
		X"2A",X"FF",X"D7",X"FE",X"87",X"FE",X"38",X"FE",X"EE",X"FD",X"A3",X"FD",X"5C",X"FD",X"17",X"FD",
		X"D4",X"FC",X"95",X"FC",X"55",X"FC",X"18",X"FC",X"DE",X"FB",X"A5",X"FB",X"6F",X"FB",X"3A",X"FB",
		X"06",X"FB",X"D4",X"FA",X"A3",X"FA",X"74",X"FA",X"47",X"FA",X"1C",X"FA",X"F1",X"F9",X"C7",X"F9",
		X"A0",X"F9",X"7A",X"F9",X"54",X"F9",X"31",X"F9",X"0E",X"F9",X"ED",X"F8",X"CC",X"F8",X"AE",X"F8",
		X"90",X"F8",X"73",X"F8",X"57",X"F8",X"3E",X"F8",X"23",X"F8",X"09",X"F8",X"F3",X"F7",X"DA",X"F7",
		X"C6",X"F7",X"AF",X"F7",X"9A",X"F7",X"86",X"F7",X"72",X"F7",X"60",X"F7",X"50",X"F7",X"3E",X"F7",
		X"2E",X"F7",X"1E",X"F7",X"10",X"F7",X"02",X"F7",X"F4",X"F6",X"E7",X"F6",X"DA",X"F6",X"CF",X"F6",
		X"C3",X"F6",X"B9",X"F6",X"AF",X"F6",X"A4",X"F6",X"9B",X"F6",X"91",X"F6",X"8A",X"F6",X"82",X"F6",
		X"7A",X"F6",X"73",X"F6",X"6D",X"F6",X"65",X"F6",X"60",X"F6",X"5A",X"F6",X"55",X"F6",X"50",X"F6",
		X"4C",X"F6",X"47",X"F6",X"43",X"F6",X"40",X"F6",X"3C",X"F6",X"39",X"F6",X"36",X"F6",X"34",X"F6",
		X"32",X"F6",X"31",X"F6",X"30",X"F6",X"2D",X"F6",X"2E",X"F6",X"2C",X"F6",X"2B",X"F6",X"2B",X"F6",
		X"2A",X"F6",X"28",X"F6",X"2C",X"F6",X"2B",X"F6",X"2C",X"F6",X"2C",X"F6",X"2D",X"F6",X"2D",X"F6",
		X"30",X"F6",X"30",X"F6",X"34",X"F6",X"34",X"F6",X"36",X"F6",X"38",X"F6",X"3B",X"F6",X"3C",X"F6",
		X"3E",X"F6",X"42",X"F6",X"44",X"F6",X"48",X"F6",X"4B",X"F6",X"4D",X"F6",X"51",X"F6",X"54",X"F6",
		X"57",X"F6",X"5B",X"F6",X"5E",X"F6",X"61",X"F6",X"65",X"F6",X"6A",X"F6",X"6D",X"F6",X"71",X"F6",
		X"75",X"F6",X"78",X"F6",X"7E",X"F6",X"82",X"F6",X"86",X"F6",X"8B",X"F6",X"90",X"F6",X"93",X"F6",
		X"97",X"F6",X"9E",X"F6",X"A1",X"F6",X"A5",X"F6",X"AC",X"F6",X"B1",X"F6",X"B4",X"F6",X"BA",X"F6",
		X"BE",X"F6",X"C4",X"F6",X"C8",X"F6",X"CE",X"F6",X"D4",X"F6",X"D9",X"F6",X"DD",X"F6",X"0F",X"F7",
		X"7B",X"F7",X"0A",X"F8",X"AD",X"F8",X"60",X"F9",X"18",X"FA",X"D7",X"FA",X"94",X"FB",X"51",X"FC",
		X"0B",X"FD",X"C0",X"FD",X"72",X"FE",X"21",X"FF",X"CB",X"FF",X"6E",X"00",X"0F",X"01",X"AB",X"01",
		X"42",X"02",X"D6",X"02",X"63",X"03",X"EC",X"03",X"72",X"04",X"F5",X"04",X"72",X"05",X"ED",X"05",
		X"62",X"06",X"D5",X"06",X"46",X"07",X"B2",X"07",X"1A",X"08",X"80",X"08",X"E1",X"08",X"40",X"09",
		X"9C",X"09",X"F5",X"09",X"4B",X"0A",X"A0",X"0A",X"F0",X"0A",X"3E",X"0B",X"8A",X"0B",X"D4",X"0B",
		X"1B",X"0C",X"5F",X"0C",X"A1",X"0C",X"E2",X"0C",X"21",X"0D",X"5C",X"0D",X"95",X"0D",X"CD",X"0D",
		X"03",X"0E",X"37",X"0E",X"6A",X"0E",X"9B",X"0E",X"CA",X"0E",X"F8",X"0E",X"24",X"0F",X"4F",X"0F",
		X"76",X"0F",X"9F",X"0F",X"C4",X"0F",X"E9",X"0F",X"0E",X"10",X"2E",X"10",X"50",X"10",X"6E",X"10",
		X"8D",X"10",X"AA",X"10",X"C5",X"10",X"E0",X"10",X"FB",X"10",X"14",X"11",X"29",X"11",X"40",X"11",
		X"56",X"11",X"6A",X"11",X"7F",X"11",X"93",X"11",X"A5",X"11",X"B6",X"11",X"C8",X"11",X"CC",X"11",
		X"C0",X"11",X"B7",X"11",X"AC",X"11",X"56",X"11",X"CD",X"10",X"38",X"10",X"90",X"0F",X"E7",X"0E",
		X"37",X"0E",X"89",X"0D",X"DC",X"0C",X"31",X"0C",X"88",X"0B",X"E5",X"0A",X"44",X"0A",X"A8",X"09",
		X"0D",X"09",X"7B",X"08",X"E9",X"07",X"5E",X"07",X"D5",X"06",X"52",X"06",X"D1",X"05",X"54",X"05",
		X"DC",X"04",X"67",X"04",X"F4",X"03",X"87",X"03",X"1B",X"03",X"B5",X"02",X"4F",X"02",X"EE",X"01",
		X"90",X"01",X"32",X"01",X"DA",X"00",X"83",X"00",X"2E",X"00",X"DF",X"FF",X"8F",X"FF",X"42",X"FF",
		X"F8",X"FE",X"B1",X"FE",X"6A",X"FE",X"25",X"FE",X"E6",X"FD",X"A6",X"FD",X"69",X"FD",X"2E",X"FD",
		X"F5",X"FC",X"BA",X"FC",X"85",X"FC",X"50",X"FC",X"1E",X"FC",X"EC",X"FB",X"BD",X"FB",X"8E",X"FB",
		X"66",X"FB",X"73",X"FB",X"B8",X"FB",X"1C",X"FC",X"9A",X"FC",X"21",X"FD",X"B2",X"FD",X"48",X"FE",
		X"DC",X"FE",X"73",X"FF",X"05",X"00",X"95",X"00",X"25",X"01",X"B0",X"01",X"37",X"02",X"BD",X"02",
		X"3B",X"03",X"B9",X"03",X"2F",X"04",X"A5",X"04",X"16",X"05",X"85",X"05",X"F0",X"05",X"59",X"06",
		X"BC",X"06",X"1C",X"07",X"7D",X"07",X"D8",X"07",X"2F",X"08",X"85",X"08",X"D8",X"08",X"29",X"09",
		X"77",X"09",X"C2",X"09",X"0B",X"0A",X"51",X"0A",X"96",X"0A",X"D9",X"0A",X"1A",X"0B",X"56",X"0B",
		X"92",X"0B",X"CC",X"0B",X"05",X"0C",X"3A",X"0C",X"6E",X"0C",X"A2",X"0C",X"D2",X"0C",X"01",X"0D",
		X"2F",X"0D",X"5B",X"0D",X"85",X"0D",X"AE",X"0D",X"D6",X"0D",X"FA",X"0D",X"1F",X"0E",X"44",X"0E",
		X"66",X"0E",X"87",X"0E",X"A7",X"0E",X"C4",X"0E",X"E2",X"0E",X"FC",X"0E",X"1A",X"0F",X"34",X"0F",
		X"4C",X"0F",X"65",X"0F",X"7D",X"0F",X"91",X"0F",X"A7",X"0F",X"BB",X"0F",X"CE",X"0F",X"E1",X"0F",
		X"F3",X"0F",X"02",X"10",X"FD",X"0F",X"F5",X"0F",X"EC",X"0F",X"E2",X"0F",X"D9",X"0F",X"CF",X"0F",
		X"C6",X"0F",X"BE",X"0F",X"B5",X"0F",X"AA",X"0F",X"A1",X"0F",X"9A",X"0F",X"91",X"0F",X"86",X"0F",
		X"80",X"0F",X"76",X"0F",X"6D",X"0F",X"64",X"0F",X"5D",X"0F",X"53",X"0F",X"4A",X"0F",X"42",X"0F",
		X"39",X"0F",X"30",X"0F",X"26",X"0F",X"1E",X"0F",X"15",X"0F",X"0D",X"0F",X"05",X"0F",X"FC",X"0E",
		X"F3",X"0E",X"EB",X"0E",X"E2",X"0E",X"D9",X"0E",X"D1",X"0E",X"C9",X"0E",X"C0",X"0E",X"B8",X"0E",
		X"AF",X"0E",X"A7",X"0E",X"9F",X"0E",X"8F",X"0E",X"FC",X"0D",X"3C",X"0D",X"86",X"0C",X"C9",X"0B",
		X"14",X"0B",X"5C",X"0A",X"AF",X"09",X"01",X"09",X"5A",X"08",X"B7",X"07",X"19",X"07",X"7D",X"06",
		X"E8",X"05",X"56",X"05",X"C8",X"04",X"3F",X"04",X"BA",X"03",X"38",X"03",X"BA",X"02",X"3F",X"02",
		X"CA",X"01",X"58",X"01",X"E9",X"00",X"7B",X"00",X"14",X"00",X"AE",X"FF",X"4C",X"FF",X"EC",X"FE",
		X"90",X"FE",X"36",X"FE",X"DF",X"FD",X"8B",X"FD",X"38",X"FD",X"E9",X"FC",X"9E",X"FC",X"53",X"FC",
		X"0A",X"FC",X"C4",X"FB",X"81",X"FB",X"3F",X"FB",X"00",X"FB",X"C3",X"FA",X"87",X"FA",X"4C",X"FA",
		X"15",X"FA",X"E0",X"F9",X"AC",X"F9",X"79",X"F9",X"4A",X"F9",X"18",X"F9",X"0B",X"F9",X"3D",X"F9",
		X"95",X"F9",X"06",X"FA",X"89",X"FA",X"17",X"FB",X"A8",X"FB",X"3D",X"FC",X"D1",X"FC",X"65",X"FD",
		X"F7",X"FD",X"84",X"FE",X"0F",X"FF",X"96",X"FF",X"1A",X"00",X"9B",X"00",X"17",X"01",X"8F",X"01",
		X"06",X"02",X"78",X"02",X"E7",X"02",X"53",X"03",X"BB",X"03",X"20",X"04",X"83",X"04",X"E2",X"04",
		X"3E",X"05",X"99",X"05",X"ED",X"05",X"41",X"06",X"92",X"06",X"E2",X"06",X"2F",X"07",X"78",X"07",
		X"C0",X"07",X"05",X"08",X"47",X"08",X"89",X"08",X"C8",X"08",X"05",X"09",X"3F",X"09",X"78",X"09",
		X"AE",X"09",X"E4",X"09",X"18",X"0A",X"4A",X"0A",X"7A",X"0A",X"A8",X"0A",X"D5",X"0A",X"02",X"0B",
		X"2B",X"0B",X"54",X"0B",X"7A",X"0B",X"9F",X"0B",X"C5",X"0B",X"E8",X"0B",X"0A",X"0C",X"2A",X"0C",
		X"4A",X"0C",X"68",X"0C",X"85",X"0C",X"A0",X"0C",X"BD",X"0C",X"D6",X"0C",X"F0",X"0C",X"08",X"0D",
		X"1F",X"0D",X"35",X"0D",X"4B",X"0D",X"5E",X"0D",X"73",X"0D",X"86",X"0D",X"95",X"0D",X"90",X"0D",
		X"89",X"0D",X"80",X"0D",X"79",X"0D",X"71",X"0D",X"6B",X"0D",X"61",X"0D",X"5B",X"0D",X"52",X"0D",
		X"4C",X"0D",X"42",X"0D",X"3E",X"0D",X"D6",X"0C",X"31",X"0C",X"8B",X"0B",X"DA",X"0A",X"2B",X"0A",
		X"7A",X"09",X"CC",X"08",X"1F",X"08",X"79",X"07",X"D2",X"06",X"32",X"06",X"93",X"05",X"FD",X"04",
		X"68",X"04",X"D8",X"03",X"4C",X"03",X"C5",X"02",X"41",X"02",X"C1",X"01",X"46",X"01",X"CE",X"00",
		X"59",X"00",X"E9",X"FF",X"7A",X"FF",X"10",X"FF",X"AA",X"FE",X"46",X"FE",X"E4",X"FD",X"86",X"FD",
		X"2A",X"FD",X"D2",X"FC",X"7C",X"FC",X"29",X"FC",X"DB",X"FB",X"8A",X"FB",X"40",X"FB",X"F6",X"FA",
		X"AF",X"FA",X"6B",X"FA",X"28",X"FA",X"E9",X"F9",X"AB",X"F9",X"6D",X"F9",X"34",X"F9",X"FB",X"F8",
		X"C3",X"F8",X"8F",X"F8",X"5C",X"F8",X"2A",X"F8",X"F9",X"F7",X"CD",X"F7",X"9F",X"F7",X"81",X"F7",
		X"A1",X"F7",X"F1",X"F7",X"5E",X"F8",X"DE",X"F8",X"6B",X"F9",X"FE",X"F9",X"95",X"FA",X"2D",X"FB",
		X"C2",X"FB",X"58",X"FC",X"E7",X"FC",X"78",X"FD",X"03",X"FE",X"8A",X"FE",X"0F",X"FF",X"8F",X"FF",
		X"0A",X"00",X"82",X"00",X"FA",X"00",X"6A",X"01",X"DA",X"01",X"44",X"02",X"AE",X"02",X"12",X"03",
		X"74",X"03",X"D3",X"03",X"30",X"04",X"63",X"04",X"58",X"04",X"27",X"04",X"DA",X"03",X"7D",X"03",
		X"15",X"03",X"A7",X"02",X"37",X"02",X"C5",X"01",X"54",X"01",X"E4",X"00",X"76",X"00",X"0A",X"00",
		X"A1",X"FF",X"3A",X"FF",X"D6",X"FE",X"76",X"FE",X"17",X"FE",X"BC",X"FD",X"63",X"FD",X"0D",X"FD",
		X"B9",X"FC",X"68",X"FC",X"19",X"FC",X"CD",X"FB",X"85",X"FB",X"3C",X"FB",X"F7",X"FA",X"B3",X"FA",
		X"73",X"FA",X"35",X"FA",X"F7",X"F9",X"BC",X"F9",X"84",X"F9",X"4D",X"F9",X"19",X"F9",X"E3",X"F8",
		X"B3",X"F8",X"81",X"F8",X"52",X"F8",X"24",X"F8",X"FA",X"F7",X"D0",X"F7",X"A6",X"F7",X"7F",X"F7",
		X"59",X"F7",X"35",X"F7",X"12",X"F7",X"F0",X"F6",X"CE",X"F6",X"AE",X"F6",X"91",X"F6",X"72",X"F6",
		X"56",X"F6",X"3A",X"F6",X"3D",X"F6",X"80",X"F6",X"E7",X"F6",X"6B",X"F7",X"FF",X"F7",X"9D",X"F8",
		X"3E",X"F9",X"E2",X"F9",X"86",X"FA",X"29",X"FB",X"C7",X"FB",X"65",X"FC",X"FE",X"FC",X"93",X"FD",
		X"25",X"FE",X"B3",X"FE",X"3B",X"FF",X"C1",X"FF",X"41",X"00",X"BE",X"00",X"38",X"01",X"B0",X"01",
		X"22",X"02",X"92",X"02",X"FE",X"02",X"66",X"03",X"CE",X"03",X"2A",X"04",X"50",X"04",X"3D",X"04",
		X"0A",X"04",X"BD",X"03",X"63",X"03",X"FF",X"02",X"95",X"02",X"2C",X"02",X"BE",X"01",X"53",X"01",
		X"E8",X"00",X"7E",X"00",X"19",X"00",X"B7",X"FF",X"55",X"FF",X"F7",X"FE",X"9B",X"FE",X"41",X"FE",
		X"EA",X"FD",X"97",X"FD",X"46",X"FD",X"F6",X"FC",X"AA",X"FC",X"61",X"FC",X"17",X"FC",X"D4",X"FB",
		X"8D",X"FB",X"63",X"FB",X"78",X"FB",X"B8",X"FB",X"16",X"FC",X"86",X"FC",X"00",X"FD",X"81",X"FD",
		X"06",X"FE",X"8B",X"FE",X"10",X"FF",X"93",X"FF",X"12",X"00",X"90",X"00",X"0A",X"01",X"83",X"01",
		X"F6",X"01",X"67",X"02",X"D5",X"02",X"40",X"03",X"A7",X"03",X"0B",X"04",X"6E",X"04",X"CD",X"04",
		X"28",X"05",X"80",X"05",X"D5",X"05",X"28",X"06",X"7A",X"06",X"C8",X"06",X"13",X"07",X"5D",X"07",
		X"A4",X"07",X"E8",X"07",X"2B",X"08",X"6E",X"08",X"AB",X"08",X"E8",X"08",X"21",X"09",X"5B",X"09",
		X"91",X"09",X"C6",X"09",X"F9",X"09",X"2A",X"0A",X"5B",X"0A",X"89",X"0A",X"B6",X"0A",X"E0",X"0A",
		X"0A",X"0B",X"33",X"0B",X"59",X"0B",X"7F",X"0B",X"A2",X"0B",X"C6",X"0B",X"E8",X"0B",X"08",X"0C",
		X"27",X"0C",X"46",X"0C",X"62",X"0C",X"7D",X"0C",X"98",X"0C",X"B3",X"0C",X"CD",X"0C",X"E3",X"0C",
		X"FA",X"0C",X"11",X"0D",X"26",X"0D",X"3C",X"0D",X"4D",X"0D",X"62",X"0D",X"70",X"0D",X"69",X"0D",
		X"62",X"0D",X"59",X"0D",X"51",X"0D",X"48",X"0D",X"41",X"0D",X"38",X"0D",X"31",X"0D",X"28",X"0D",
		X"22",X"0D",X"1A",X"0D",X"14",X"0D",X"0A",X"0D",X"04",X"0D",X"F8",X"0C",X"F8",X"0C",X"97",X"0C",
		X"E9",X"0B",X"40",X"0B",X"8B",X"0A",X"DC",X"09",X"29",X"09",X"7B",X"08",X"CD",X"07",X"26",X"07",
		X"80",X"06",X"E0",X"05",X"43",X"05",X"AC",X"04",X"19",X"04",X"89",X"03",X"FD",X"02",X"76",X"02",
		X"F3",X"01",X"74",X"01",X"F7",X"00",X"80",X"00",X"0B",X"00",X"9D",X"FF",X"2D",X"FF",X"CE",X"FE",
		X"AC",X"FE",X"BE",X"FE",X"F1",X"FE",X"38",X"FF",X"8E",X"FF",X"EB",X"FF",X"4E",X"00",X"B2",X"00",
		X"18",X"01",X"7F",X"01",X"E2",X"01",X"43",X"02",X"A4",X"02",X"02",X"03",X"5D",X"03",X"B5",X"03",
		X"0B",X"04",X"5E",X"04",X"AF",X"04",X"FE",X"04",X"4A",X"05",X"95",X"05",X"DD",X"05",X"22",X"06",
		X"64",X"06",X"A8",X"06",X"E5",X"06",X"22",X"07",X"5E",X"07",X"97",X"07",X"CE",X"07",X"03",X"08",
		X"37",X"08",X"6A",X"08",X"9B",X"08",X"CA",X"08",X"F7",X"08",X"23",X"09",X"4C",X"09",X"75",X"09",
		X"9E",X"09",X"C3",X"09",X"E8",X"09",X"0D",X"0A",X"2E",X"0A",X"50",X"0A",X"71",X"0A",X"91",X"0A",
		X"AD",X"0A",X"CA",X"0A",X"E5",X"0A",X"FF",X"0A",X"1A",X"0B",X"33",X"0B",X"4B",X"0B",X"61",X"0B",
		X"76",X"0B",X"8D",X"0B",X"A0",X"0B",X"B6",X"0B",X"C2",X"0B",X"BC",X"0B",X"B4",X"0B",X"AE",X"0B",
		X"A7",X"0B",X"A0",X"0B",X"9A",X"0B",X"93",X"0B",X"8C",X"0B",X"85",X"0B",X"7D",X"0B",X"77",X"0B",
		X"70",X"0B",X"69",X"0B",X"63",X"0B",X"5C",X"0B",X"56",X"0B",X"4E",X"0B",X"46",X"0B",X"41",X"0B",
		X"3B",X"0B",X"33",X"0B",X"2B",X"0B",X"28",X"0B",X"1C",X"0B",X"1B",X"0B",X"B8",X"0A",X"00",X"0A",
		X"51",X"09",X"9B",X"08",X"E8",X"07",X"35",X"07",X"87",X"06",X"DA",X"05",X"34",X"05",X"8F",X"04",
		X"F0",X"03",X"55",X"03",X"BF",X"02",X"2D",X"02",X"A0",X"01",X"15",X"01",X"8F",X"00",X"0E",X"00",
		X"92",X"FF",X"17",X"FF",X"9F",X"FE",X"2E",X"FE",X"BD",X"FD",X"66",X"FD",X"51",X"FD",X"66",X"FD",
		X"9E",X"FD",X"E5",X"FD",X"3B",X"FE",X"98",X"FE",X"FA",X"FE",X"5D",X"FF",X"C2",X"FF",X"23",X"00",
		X"85",X"00",X"E6",X"00",X"43",X"01",X"A0",X"01",X"FA",X"01",X"4E",X"02",X"A3",X"02",X"F6",X"02",
		X"46",X"03",X"92",X"03",X"DE",X"03",X"26",X"04",X"6D",X"04",X"B0",X"04",X"F3",X"04",X"32",X"05",
		X"6F",X"05",X"7D",X"05",X"4F",X"05",X"FE",X"04",X"93",X"04",X"1B",X"04",X"99",X"03",X"11",X"03",
		X"8A",X"02",X"03",X"02",X"7B",X"01",X"F6",X"00",X"72",X"00",X"F3",X"FF",X"78",X"FF",X"FE",X"FE",
		X"87",X"FE",X"14",X"FE",X"A6",X"FD",X"3A",X"FD",X"D3",X"FC",X"6C",X"FC",X"0A",X"FC",X"AA",X"FB",
		X"4D",X"FB",X"F4",X"FA",X"9E",X"FA",X"47",X"FA",X"05",X"FA",X"01",X"FA",X"2C",X"FA",X"78",X"FA",
		X"D6",X"FA",X"42",X"FB",X"B5",X"FB",X"2D",X"FC",X"A6",X"FC",X"1E",X"FD",X"94",X"FD",X"0B",X"FE",
		X"7F",X"FE",X"F0",X"FE",X"5D",X"FF",X"C8",X"FF",X"30",X"00",X"96",X"00",X"F9",X"00",X"56",X"01",
		X"B4",X"01",X"0E",X"02",X"65",X"02",X"B9",X"02",X"0C",X"03",X"5A",X"03",X"A7",X"03",X"F1",X"03",
		X"3B",X"04",X"81",X"04",X"C5",X"04",X"08",X"05",X"47",X"05",X"84",X"05",X"C0",X"05",X"FA",X"05",
		X"32",X"06",X"69",X"06",X"9C",X"06",X"D0",X"06",X"02",X"07",X"30",X"07",X"5F",X"07",X"8C",X"07",
		X"B6",X"07",X"DF",X"07",X"08",X"08",X"30",X"08",X"54",X"08",X"7A",X"08",X"9D",X"08",X"C0",X"08",
		X"DE",X"08",X"FE",X"08",X"1D",X"09",X"3B",X"09",X"57",X"09",X"73",X"09",X"8D",X"09",X"A5",X"09",
		X"C0",X"09",X"D7",X"09",X"ED",X"09",X"03",X"0A",X"18",X"0A",X"2E",X"0A",X"3D",X"0A",X"39",X"0A",
		X"33",X"0A",X"2E",X"0A",X"28",X"0A",X"20",X"0A",X"19",X"0A",X"13",X"0A",X"0E",X"0A",X"08",X"0A",
		X"01",X"0A",X"FB",X"09",X"F5",X"09",X"F1",X"09",X"EA",X"09",X"E3",X"09",X"DD",X"09",X"D7",X"09",
		X"D1",X"09",X"CB",X"09",X"C6",X"09",X"BE",X"09",X"B9",X"09",X"B2",X"09",X"AD",X"09",X"A7",X"09",
		X"A1",X"09",X"99",X"09",X"94",X"09",X"8F",X"09",X"8A",X"09",X"84",X"09",X"7F",X"09",X"78",X"09",
		X"74",X"09",X"6D",X"09",X"67",X"09",X"61",X"09",X"5C",X"09",X"54",X"09",X"50",X"09",X"4B",X"09",
		X"45",X"09",X"3F",X"09",X"39",X"09",X"33",X"09",X"2E",X"09",X"29",X"09",X"25",X"09",X"10",X"09",
		X"78",X"08",X"B9",X"07",X"02",X"07",X"49",X"06",X"95",X"05",X"E2",X"04",X"36",X"04",X"8C",X"03",
		X"E9",X"02",X"45",X"02",X"A9",X"01",X"13",X"01",X"7F",X"00",X"F0",X"FF",X"67",X"FF",X"E0",X"FE",
		X"5E",X"FE",X"DF",X"FD",X"63",X"FD",X"ED",X"FC",X"79",X"FC",X"09",X"FC",X"9E",X"FB",X"35",X"FB",
		X"CE",X"FA",X"6B",X"FA",X"0C",X"FA",X"AF",X"F9",X"56",X"F9",X"FE",X"F8",X"AA",X"F8",X"58",X"F8",
		X"09",X"F8",X"BD",X"F7",X"72",X"F7",X"2B",X"F7",X"E7",X"F6",X"A2",X"F6",X"63",X"F6",X"22",X"F6",
		X"E6",X"F5",X"AB",X"F5",X"73",X"F5",X"3B",X"F5",X"06",X"F5",X"D2",X"F4",X"A2",X"F4",X"71",X"F4",
		X"44",X"F4",X"19",X"F4",X"20",X"F4",X"61",X"F4",X"C7",X"F4",X"3F",X"F5",X"C7",X"F5",X"59",X"F6",
		X"ED",X"F6",X"84",X"F7",X"1B",X"F8",X"B1",X"F8",X"42",X"F9",X"D3",X"F9",X"5E",X"FA",X"E7",X"FA",
		X"6C",X"FB",X"EE",X"FB",X"6C",X"FC",X"E5",X"FC",X"5D",X"FD",X"D0",X"FD",X"41",X"FE",X"AE",X"FE",
		X"18",X"FF",X"7F",X"FF",X"E2",X"FF",X"41",X"00",X"A1",X"00",X"EA",X"00",X"F1",X"00",X"CD",X"00",
		X"89",X"00",X"33",X"00",X"CE",X"FF",X"63",X"FF",X"F5",X"FE",X"84",X"FE",X"12",X"FE",X"A3",X"FD",
		X"35",X"FD",X"C9",X"FC",X"60",X"FC",X"F9",X"FB",X"95",X"FB",X"34",X"FB",X"D6",X"FA",X"7A",X"FA",
		X"21",X"FA",X"CB",X"F9",X"77",X"F9",X"27",X"F9",X"D9",X"F8",X"8D",X"F8",X"44",X"F8",X"FB",X"F7",
		X"B9",X"F7",X"77",X"F7",X"35",X"F7",X"F6",X"F6",X"BA",X"F6",X"7F",X"F6",X"48",X"F6",X"10",X"F6",
		X"DD",X"F5",X"A8",X"F5",X"78",X"F5",X"47",X"F5",X"1A",X"F5",X"EE",X"F4",X"C3",X"F4",X"99",X"F4",
		X"71",X"F4",X"4B",X"F4",X"26",X"F4",X"02",X"F4",X"E0",X"F3",X"BE",X"F3",X"9C",X"F3",X"7F",X"F3",
		X"61",X"F3",X"44",X"F3",X"29",X"F3",X"0E",X"F3",X"00",X"F3",X"2F",X"F3",X"8E",X"F3",X"0A",X"F4",
		X"9A",X"F4",X"37",X"F5",X"D8",X"F5",X"7E",X"F6",X"23",X"F7",X"C7",X"F7",X"6C",X"F8",X"09",X"F9",
		X"A5",X"F9",X"3C",X"FA",X"D1",X"FA",X"61",X"FB",X"EF",X"FB",X"77",X"FC",X"FA",X"FC",X"7A",X"FD",
		X"F7",X"FD",X"70",X"FE",X"E5",X"FE",X"58",X"FF",X"C6",X"FF",X"31",X"00",X"98",X"00",X"00",X"01",
		X"3D",X"01",X"3F",X"01",X"17",X"01",X"D3",X"00",X"7D",X"00",X"1E",X"00",X"B8",X"FF",X"4F",X"FF",
		X"E3",X"FE",X"79",X"FE",X"10",X"FE",X"A9",X"FD",X"43",X"FD",X"E0",X"FC",X"7F",X"FC",X"22",X"FC",
		X"C5",X"FB",X"6D",X"FB",X"16",X"FB",X"C3",X"FA",X"73",X"FA",X"23",X"FA",X"D9",X"F9",X"8E",X"F9",
		X"46",X"F9",X"03",X"F9",X"C0",X"F8",X"7F",X"F8",X"40",X"F8",X"04",X"F8",X"CA",X"F7",X"91",X"F7",
		X"5A",X"F7",X"24",X"F7",X"F1",X"F6",X"BF",X"F6",X"90",X"F6",X"61",X"F6",X"34",X"F6",X"08",X"F6",
		X"DE",X"F5",X"B7",X"F5",X"90",X"F5",X"6C",X"F5",X"45",X"F5",X"23",X"F5",X"00",X"F5",X"E1",X"F4",
		X"C1",X"F4",X"A5",X"F4",X"85",X"F4",X"6A",X"F4",X"4F",X"F4",X"38",X"F4",X"1B",X"F4",X"1F",X"F4",
		X"61",X"F4",X"CB",X"F4",X"50",X"F5",X"E5",X"F5",X"86",X"F6",X"28",X"F7",X"D0",X"F7",X"76",X"F8",
		X"1A",X"F9",X"BD",X"F9",X"5C",X"FA",X"F8",X"FA",X"8F",X"FB",X"22",X"FC",X"B2",X"FC",X"3D",X"FD",
		X"C5",X"FD",X"47",X"FE",X"C8",X"FE",X"44",X"FF",X"BC",X"FF",X"31",X"00",X"A1",X"00",X"0E",X"01",
		X"78",X"01",X"E2",X"01",X"45",X"02",X"A7",X"02",X"04",X"03",X"60",X"03",X"B9",X"03",X"10",X"04",
		X"62",X"04",X"B3",X"04",X"00",X"05",X"4D",X"05",X"96",X"05",X"DC",X"05",X"22",X"06",X"64",X"06",
		X"A5",X"06",X"E5",X"06",X"1F",X"07",X"5B",X"07",X"94",X"07",X"CA",X"07",X"00",X"08",X"34",X"08",
		X"65",X"08",X"95",X"08",X"C2",X"08",X"F1",X"08",X"1B",X"09",X"46",X"09",X"6F",X"09",X"95",X"09",
		X"BC",X"09",X"E1",X"09",X"02",X"0A",X"25",X"0A",X"47",X"0A",X"66",X"0A",X"84",X"0A",X"A2",X"0A",
		X"BF",X"0A",X"D9",X"0A",X"F4",X"0A",X"0C",X"0B",X"26",X"0B",X"3E",X"0B",X"55",X"0B",X"6A",X"0B",
		X"7E",X"0B",X"92",X"0B",X"A6",X"0B",X"B4",X"0B",X"AD",X"0B",X"A7",X"0B",X"A1",X"0B",X"99",X"0B",
		X"93",X"0B",X"8B",X"0B",X"85",X"0B",X"7E",X"0B",X"76",X"0B",X"6F",X"0B",X"68",X"0B",X"62",X"0B",
		X"5A",X"0B",X"55",X"0B",X"4E",X"0B",X"47",X"0B",X"41",X"0B",X"3A",X"0B",X"33",X"0B",X"2A",X"0B",
		X"27",X"0B",X"1F",X"0B",X"19",X"0B",X"11",X"0B",X"0B",X"0B",X"03",X"0B",X"FD",X"0A",X"F6",X"0A",
		X"F1",X"0A",X"E9",X"0A",X"E3",X"0A",X"DD",X"0A",X"D7",X"0A",X"CE",X"0A",X"C9",X"0A",X"C1",X"0A",
		X"C0",X"0A",X"99",X"0A",X"F2",X"09",X"3A",X"09",X"82",X"08",X"CA",X"07",X"16",X"07",X"63",X"06",
		X"B6",X"05",X"0B",X"05",X"68",X"04",X"C7",X"03",X"2B",X"03",X"92",X"02",X"FE",X"01",X"6F",X"01",
		X"E4",X"00",X"5C",X"00",X"DA",X"FF",X"5C",X"FF",X"E0",X"FE",X"68",X"FE",X"F6",X"FD",X"84",X"FD",
		X"18",X"FD",X"AD",X"FC",X"47",X"FC",X"E4",X"FB",X"83",X"FB",X"27",X"FB",X"CC",X"FA",X"74",X"FA",
		X"1F",X"FA",X"CD",X"F9",X"7E",X"F9",X"33",X"F9",X"E7",X"F8",X"9E",X"F8",X"59",X"F8",X"14",X"F8",
		X"D2",X"F7",X"93",X"F7",X"57",X"F7",X"1A",X"F7",X"DF",X"F6",X"AA",X"F6",X"73",X"F6",X"3F",X"F6",
		X"0D",X"F6",X"DC",X"F5",X"AF",X"F5",X"82",X"F5",X"56",X"F5",X"2A",X"F5",X"03",X"F5",X"DA",X"F4",
		X"B6",X"F4",X"90",X"F4",X"6D",X"F4",X"4A",X"F4",X"2B",X"F4",X"0B",X"F4",X"ED",X"F3",X"CE",X"F3",
		X"B1",X"F3",X"97",X"F3",X"7C",X"F3",X"63",X"F3",X"4C",X"F3",X"34",X"F3",X"1E",X"F3",X"09",X"F3",
		X"F5",X"F2",X"E0",X"F2",X"CF",X"F2",X"BB",X"F2",X"AB",X"F2",X"9A",X"F2",X"89",X"F2",X"7B",X"F2",
		X"6C",X"F2",X"5F",X"F2",X"53",X"F2",X"46",X"F2",X"3B",X"F2",X"2F",X"F2",X"24",X"F2",X"1A",X"F2",
		X"12",X"F2",X"09",X"F2",X"00",X"F2",X"F7",X"F1",X"F0",X"F1",X"EA",X"F1",X"E3",X"F1",X"DD",X"F1",
		X"D6",X"F1",X"D2",X"F1",X"CD",X"F1",X"CA",X"F1",X"C5",X"F1",X"C2",X"F1",X"BE",X"F1",X"BC",X"F1",
		X"BA",X"F1",X"B8",X"F1",X"B4",X"F1",X"B3",X"F1",X"B2",X"F1",X"B1",X"F1",X"B0",X"F1",X"AF",X"F1",
		X"B1",X"F1",X"AF",X"F1",X"B0",X"F1",X"B1",X"F1",X"B2",X"F1",X"B2",X"F1",X"B4",X"F1",X"B5",X"F1",
		X"B8",X"F1",X"B9",X"F1",X"BD",X"F1",X"BF",X"F1",X"C1",X"F1",X"C4",X"F1",X"C6",X"F1",X"CA",X"F1",
		X"CD",X"F1",X"D1",X"F1",X"D3",X"F1",X"D7",X"F1",X"DB",X"F1",X"DF",X"F1",X"E3",X"F1",X"E8",X"F1",
		X"EB",X"F1",X"F1",X"F1",X"F5",X"F1",X"FA",X"F1",X"FE",X"F1",X"04",X"F2",X"09",X"F2",X"0E",X"F2",
		X"13",X"F2",X"19",X"F2",X"1F",X"F2",X"24",X"F2",X"29",X"F2",X"2F",X"F2",X"35",X"F2",X"3B",X"F2",
		X"42",X"F2",X"46",X"F2",X"4C",X"F2",X"53",X"F2",X"5A",X"F2",X"61",X"F2",X"66",X"F2",X"6C",X"F2",
		X"73",X"F2",X"7A",X"F2",X"80",X"F2",X"88",X"F2",X"8D",X"F2",X"96",X"F2",X"9A",X"F2",X"A2",X"F2",
		X"A9",X"F2",X"B0",X"F2",X"B8",X"F2",X"BE",X"F2",X"C5",X"F2",X"CC",X"F2",X"D4",X"F2",X"DB",X"F2",
		X"E2",X"F2",X"E9",X"F2",X"F0",X"F2",X"F8",X"F2",X"FE",X"F2",X"05",X"F3",X"0D",X"F3",X"14",X"F3",
		X"1C",X"F3",X"24",X"F3",X"2B",X"F3",X"32",X"F3",X"39",X"F3",X"42",X"F3",X"75",X"F3",X"E3",X"F3",
		X"72",X"F4",X"19",X"F5",X"CF",X"F5",X"8C",X"F6",X"49",X"F7",X"0A",X"F8",X"C8",X"F8",X"84",X"F9",
		X"3C",X"FA",X"F1",X"FA",X"A0",X"FB",X"4C",X"FC",X"F3",X"FC",X"94",X"FD",X"34",X"FE",X"CB",X"FE",
		X"60",X"FF",X"EF",X"FF",X"7B",X"00",X"02",X"01",X"87",X"01",X"06",X"02",X"82",X"02",X"FC",X"02",
		X"6F",X"03",X"D4",X"03",X"F8",X"03",X"EC",X"03",X"C1",X"03",X"7D",X"03",X"2D",X"03",X"D4",X"02",
		X"77",X"02",X"17",X"02",X"B7",X"01",X"56",X"01",X"F9",X"00",X"9A",X"00",X"3F",X"00",X"E5",X"FF",
		X"90",X"FF",X"3C",X"FF",X"E9",X"FE",X"99",X"FE",X"4C",X"FE",X"01",X"FE",X"B8",X"FD",X"72",X"FD",
		X"2D",X"FD",X"EB",X"FC",X"AA",X"FC",X"6D",X"FC",X"30",X"FC",X"F5",X"FB",X"BF",X"FB",X"85",X"FB",
		X"52",X"FB",X"1D",X"FB",X"EE",X"FA",X"BB",X"FA",X"8D",X"FA",X"60",X"FA",X"33",X"FA",X"0A",X"FA",
		X"E2",X"F9",X"B9",X"F9",X"93",X"F9",X"71",X"F9",X"4C",X"F9",X"29",X"F9",X"08",X"F9",X"E8",X"F8",
		X"CA",X"F8",X"AA",X"F8",X"8E",X"F8",X"72",X"F8",X"58",X"F8",X"3D",X"F8",X"24",X"F8",X"0C",X"F8",
		X"FC",X"F7",X"28",X"F8",X"84",X"F8",X"FF",X"F8",X"90",X"F9",X"2B",X"FA",X"D0",X"FA",X"77",X"FB",
		X"1E",X"FC",X"C4",X"FC",X"67",X"FD",X"09",X"FE",X"A5",X"FE",X"3C",X"FF",X"D3",X"FF",X"64",X"00",
		X"F1",X"00",X"79",X"01",X"FE",X"01",X"80",X"02",X"FE",X"02",X"77",X"03",X"ED",X"03",X"5F",X"04",
		X"CC",X"04",X"3A",X"05",X"A1",X"05",X"08",X"06",X"4C",X"06",X"51",X"06",X"2B",X"06",X"EA",X"05",
		X"96",X"05",X"37",X"05",X"D0",X"04",X"66",X"04",X"FB",X"03",X"90",X"03",X"26",X"03",X"BB",X"02",
		X"55",X"02",X"F0",X"01",X"8E",X"01",X"2F",X"01",X"D2",X"00",X"77",X"00",X"20",X"00",X"CC",X"FF",
		X"78",X"FF",X"2A",X"FF",X"DD",X"FE",X"8F",X"FE",X"47",X"FE",X"01",X"FE",X"BB",X"FD",X"7D",X"FD",
		X"75",X"FD",X"A5",X"FD",X"F5",X"FD",X"5D",X"FE",X"D2",X"FE",X"53",X"FF",X"D5",X"FF",X"59",X"00",
		X"DD",X"00",X"60",X"01",X"E1",X"01",X"61",X"02",X"DB",X"02",X"56",X"03",X"CB",X"03",X"3D",X"04",
		X"AA",X"04",X"17",X"05",X"7F",X"05",X"E4",X"05",X"47",X"06",X"A6",X"06",X"01",X"07",X"5C",X"07",
		X"B2",X"07",X"04",X"08",X"58",X"08",X"A6",X"08",X"F2",X"08",X"3D",X"09",X"83",X"09",X"C7",X"09",
		X"0B",X"0A",X"4B",X"0A",X"8A",X"0A",X"C8",X"0A",X"00",X"0B",X"39",X"0B",X"70",X"0B",X"A5",X"0B",
		X"DA",X"0B",X"0A",X"0C",X"3A",X"0C",X"67",X"0C",X"94",X"0C",X"BE",X"0C",X"E9",X"0C",X"11",X"0D",
		X"38",X"0D",X"5C",X"0D",X"80",X"0D",X"A3",X"0D",X"C4",X"0D",X"E5",X"0D",X"02",X"0E",X"22",X"0E",
		X"3E",X"0E",X"59",X"0E",X"73",X"0E",X"8D",X"0E",X"A6",X"0E",X"BE",X"0E",X"D3",X"0E",X"E8",X"0E",
		X"FD",X"0E",X"11",X"0F",X"25",X"0F",X"37",X"0F",X"4A",X"0F",X"52",X"0F",X"48",X"0F",X"40",X"0F",
		X"38",X"0F",X"2F",X"0F",X"25",X"0F",X"1B",X"0F",X"13",X"0F",X"09",X"0F",X"02",X"0F",X"F9",X"0E",
		X"F1",X"0E",X"E6",X"0E",X"E0",X"0E",X"D6",X"0E",X"CF",X"0E",X"60",X"0E",X"B2",X"0D",X"08",X"0D",
		X"52",X"0C",X"A1",X"0B",X"EE",X"0A",X"3F",X"0A",X"8F",X"09",X"E8",X"08",X"42",X"08",X"A1",X"07",
		X"03",X"07",X"6C",X"06",X"D5",X"05",X"47",X"05",X"B9",X"04",X"31",X"04",X"AD",X"03",X"2E",X"03",
		X"B0",X"02",X"38",X"02",X"C4",X"01",X"52",X"01",X"E1",X"00",X"81",X"00",X"60",X"00",X"71",X"00",
		X"A3",X"00",X"EB",X"00",X"3E",X"01",X"9C",X"01",X"FD",X"01",X"62",X"02",X"C6",X"02",X"2C",X"03",
		X"8C",X"03",X"EE",X"03",X"4D",X"04",X"AA",X"04",X"06",X"05",X"5D",X"05",X"B2",X"05",X"04",X"06",
		X"55",X"06",X"A3",X"06",X"EE",X"06",X"37",X"07",X"7D",X"07",X"C2",X"07",X"05",X"08",X"44",X"08",
		X"84",X"08",X"BF",X"08",X"F9",X"08",X"33",X"09",X"68",X"09",X"9E",X"09",X"D0",X"09",X"02",X"0A",
		X"32",X"0A",X"60",X"0A",X"8B",X"0A",X"B7",X"0A",X"DF",X"0A",X"09",X"0B",X"2F",X"0B",X"54",X"0B",
		X"77",X"0B",X"9C",X"0B",X"BB",X"0B",X"DD",X"0B",X"FC",X"0B",X"1B",X"0C",X"37",X"0C",X"52",X"0C",
		X"6D",X"0C",X"87",X"0C",X"A1",X"0C",X"B9",X"0C",X"CF",X"0C",X"E5",X"0C",X"FA",X"0C",X"0F",X"0D",
		X"22",X"0D",X"35",X"0D",X"44",X"0D",X"42",X"0D",X"39",X"0D",X"33",X"0D",X"28",X"0D",X"21",X"0D",
		X"1A",X"0D",X"12",X"0D",X"0A",X"0D",X"01",X"0D",X"F9",X"0C",X"F3",X"0C",X"EA",X"0C",X"E4",X"0C",
		X"DD",X"0C",X"D3",X"0C",X"CC",X"0C",X"C4",X"0C",X"BD",X"0C",X"B6",X"0C",X"AE",X"0C",X"A6",X"0C",
		X"9F",X"0C",X"97",X"0C",X"90",X"0C",X"89",X"0C",X"81",X"0C",X"79",X"0C",X"72",X"0C",X"6A",X"0C",
		X"63",X"0C",X"5D",X"0C",X"54",X"0C",X"4C",X"0C",X"45",X"0C",X"3E",X"0C",X"36",X"0C",X"2E",X"0C",
		X"27",X"0C",X"1F",X"0C",X"19",X"0C",X"11",X"0C",X"09",X"0C",X"02",X"0C",X"FC",X"0B",X"F5",X"0B",
		X"EE",X"0B",X"E5",X"0B",X"DF",X"0B",X"D6",X"0B",X"D2",X"0B",X"C8",X"0B",X"C5",X"0B",X"B9",X"0B",
		X"B5",X"0B",X"3B",X"0B",X"75",X"0A",X"BF",X"09",X"01",X"09",X"4D",X"08",X"95",X"07",X"E7",X"06",
		X"3A",X"06",X"93",X"05",X"EF",X"04",X"52",X"04",X"B7",X"03",X"22",X"03",X"90",X"02",X"03",X"02",
		X"79",X"01",X"F7",X"00",X"74",X"00",X"F8",X"FF",X"7F",X"FF",X"09",X"FF",X"96",X"FE",X"3B",X"FE",
		X"20",X"FE",X"34",X"FE",X"67",X"FE",X"AE",X"FE",X"00",X"FF",X"5C",X"FF",X"BC",X"FF",X"1C",X"00",
		X"7D",X"00",X"DF",X"00",X"3F",X"01",X"9C",X"01",X"F9",X"01",X"53",X"02",X"AA",X"02",X"FF",X"02",
		X"52",X"03",X"A2",X"03",X"F1",X"03",X"3B",X"04",X"85",X"04",X"CC",X"04",X"11",X"05",X"54",X"05",
		X"94",X"05",X"D2",X"05",X"0E",X"06",X"4A",X"06",X"83",X"06",X"B9",X"06",X"EE",X"06",X"22",X"07",
		X"55",X"07",X"85",X"07",X"B2",X"07",X"E0",X"07",X"0D",X"08",X"36",X"08",X"5E",X"08",X"85",X"08",
		X"AB",X"08",X"D1",X"08",X"F4",X"08",X"16",X"09",X"37",X"09",X"58",X"09",X"76",X"09",X"95",X"09",
		X"B1",X"09",X"CD",X"09",X"E7",X"09",X"00",X"0A",X"18",X"0A",X"31",X"0A",X"49",X"0A",X"5F",X"0A",
		X"73",X"0A",X"87",X"0A",X"9D",X"0A",X"A9",X"0A",X"A3",X"0A",X"9D",X"0A",X"95",X"0A",X"8F",X"0A",
		X"88",X"0A",X"81",X"0A",X"7B",X"0A",X"76",X"0A",X"6F",X"0A",X"67",X"0A",X"62",X"0A",X"5A",X"0A",
		X"55",X"0A",X"4F",X"0A",X"48",X"0A",X"42",X"0A",X"3B",X"0A",X"35",X"0A",X"2E",X"0A",X"28",X"0A",
		X"21",X"0A",X"1C",X"0A",X"14",X"0A",X"11",X"0A",X"08",X"0A",X"02",X"0A",X"88",X"09",X"D0",X"08",
		X"21",X"08",X"69",X"07",X"B8",X"06",X"05",X"06",X"57",X"05",X"AA",X"04",X"05",X"04",X"61",X"03",
		X"C5",X"02",X"29",X"02",X"96",X"01",X"04",X"01",X"77",X"00",X"EE",X"FF",X"6B",X"FF",X"E8",X"FE",
		X"6B",X"FE",X"F3",X"FD",X"7D",X"FD",X"0C",X"FD",X"9C",X"FC",X"32",X"FC",X"CC",X"FB",X"65",X"FB",
		X"06",X"FB",X"A5",X"FA",X"4A",X"FA",X"F3",X"F9",X"9C",X"F9",X"49",X"F9",X"F8",X"F8",X"AB",X"F8",
		X"5F",X"F8",X"15",X"F8",X"CE",X"F7",X"89",X"F7",X"47",X"F7",X"07",X"F7",X"C8",X"F6",X"8C",X"F6",
		X"52",X"F6",X"1A",X"F6",X"E3",X"F5",X"AF",X"F5",X"7B",X"F5",X"4B",X"F5",X"1B",X"F5",X"EE",X"F4",
		X"BF",X"F4",X"B4",X"F4",X"E5",X"F4",X"3E",X"F5",X"B4",X"F5",X"39",X"F6",X"C8",X"F6",X"5E",X"F7",
		X"F5",X"F7",X"8D",X"F8",X"23",X"F9",X"B6",X"F9",X"46",X"FA",X"D4",X"FA",X"5E",X"FB",X"E6",X"FB",
		X"69",X"FC",X"EA",X"FC",X"67",X"FD",X"DE",X"FD",X"53",X"FE",X"C3",X"FE",X"31",X"FF",X"9D",X"FF",
		X"04",X"00",X"69",X"00",X"CA",X"00",X"28",X"01",X"80",X"01",X"9F",X"01",X"86",X"01",X"4D",X"01",
		X"FB",X"00",X"9A",X"00",X"31",X"00",X"C3",X"FF",X"53",X"FF",X"E2",X"FE",X"71",X"FE",X"02",X"FE",
		X"96",X"FD",X"2C",X"FD",X"C3",X"FC",X"5E",X"FC",X"FB",X"FB",X"9E",X"FB",X"42",X"FB",X"E7",X"FA",
		X"90",X"FA",X"3C",X"FA",X"EB",X"F9",X"9B",X"F9",X"4F",X"F9",X"04",X"F9",X"BD",X"F8",X"75",X"F8",
		X"47",X"F8",X"5B",X"F8",X"9B",X"F8",X"F5",X"F8",X"62",X"F9",X"DC",X"F9",X"5C",X"FA",X"DE",X"FA",
		X"62",X"FB",X"E5",X"FB",X"66",X"FC",X"E7",X"FC",X"63",X"FD",X"DC",X"FD",X"54",X"FE",X"C8",X"FE",
		X"37",X"FF",X"A5",X"FF",X"0F",X"00",X"76",X"00",X"D9",X"00",X"3A",X"01",X"98",X"01",X"F4",X"01",
		X"4C",X"02",X"A2",X"02",X"F3",X"02",X"44",X"03",X"93",X"03",X"DE",X"03",X"28",X"04",X"71",X"04",
		X"B4",X"04",X"F7",X"04",X"38",X"05",X"76",X"05",X"B3",X"05",X"ED",X"05",X"25",X"06",X"5D",X"06",
		X"94",X"06",X"C5",X"06",X"F7",X"06",X"29",X"07",X"57",X"07",X"83",X"07",X"B0",X"07",X"DA",X"07",
		X"02",X"08",X"29",X"08",X"50",X"08",X"76",X"08",X"99",X"08",X"BC",X"08",X"DD",X"08",X"FC",X"08",
		X"1D",X"09",X"38",X"09",X"58",X"09",X"73",X"09",X"8D",X"09",X"A7",X"09",X"BF",X"09",X"D8",X"09",
		X"EF",X"09",X"04",X"0A",X"1B",X"0A",X"2E",X"0A",X"43",X"0A",X"50",X"0A",X"49",X"0A",X"44",X"0A",
		X"3D",X"0A",X"37",X"0A",X"2F",X"0A",X"2A",X"0A",X"23",X"0A",X"1E",X"0A",X"18",X"0A",X"12",X"0A",
		X"0A",X"0A",X"05",X"0A",X"FE",X"09",X"FA",X"09",X"F0",X"09",X"F1",X"09",X"8B",X"09",X"DE",X"08",
		X"37",X"08",X"83",X"07",X"D5",X"06",X"22",X"06",X"75",X"05",X"C8",X"04",X"22",X"04",X"7F",X"03",
		X"E1",X"02",X"44",X"02",X"AE",X"01",X"1B",X"01",X"8D",X"00",X"02",X"00",X"7F",X"FF",X"FB",X"FE",
		X"7E",X"FE",X"03",X"FE",X"8D",X"FD",X"19",X"FD",X"AA",X"FC",X"3D",X"FC",X"D4",X"FB",X"6E",X"FB",
		X"0D",X"FB",X"AC",X"FA",X"51",X"FA",X"F7",X"F9",X"A0",X"F9",X"4C",X"F9",X"FC",X"F8",X"AA",X"F8",
		X"5E",X"F8",X"14",X"F8",X"CD",X"F7",X"88",X"F7",X"43",X"F7",X"04",X"F7",X"C5",X"F6",X"87",X"F6",
		X"4D",X"F6",X"13",X"F6",X"DC",X"F5",X"A8",X"F5",X"74",X"F5",X"43",X"F5",X"13",X"F5",X"E5",X"F4",
		X"B7",X"F4",X"8C",X"F4",X"63",X"F4",X"3B",X"F4",X"13",X"F4",X"ED",X"F3",X"CA",X"F3",X"A6",X"F3",
		X"85",X"F3",X"65",X"F3",X"46",X"F3",X"28",X"F3",X"0B",X"F3",X"F0",X"F2",X"D3",X"F2",X"BB",X"F2",
		X"A2",X"F2",X"89",X"F2",X"74",X"F2",X"5E",X"F2",X"49",X"F2",X"35",X"F2",X"21",X"F2",X"10",X"F2",
		X"FD",X"F1",X"EE",X"F1",X"DC",X"F1",X"CD",X"F1",X"BF",X"F1",X"B1",X"F1",X"A4",X"F1",X"96",X"F1",
		X"8A",X"F1",X"80",X"F1",X"73",X"F1",X"6A",X"F1",X"61",X"F1",X"57",X"F1",X"50",X"F1",X"47",X"F1",
		X"3F",X"F1",X"39",X"F1",X"32",X"F1",X"2C",X"F1",X"27",X"F1",X"21",X"F1",X"1C",X"F1",X"19",X"F1",
		X"13",X"F1",X"10",X"F1",X"0D",X"F1",X"0A",X"F1",X"07",X"F1",X"05",X"F1",X"05",X"F1",X"02",X"F1",
		X"00",X"F1",X"00",X"F1",X"FF",X"F0",X"FE",X"F0",X"FE",X"F0",X"FF",X"F0",X"FF",X"F0",X"00",X"F1",
		X"00",X"F1",X"01",X"F1",X"03",X"F1",X"05",X"F1",X"07",X"F1",X"08",X"F1",X"0A",X"F1",X"0F",X"F1",
		X"12",X"F1",X"12",X"F1",X"16",X"F1",X"1A",X"F1",X"1C",X"F1",X"20",X"F1",X"24",X"F1",X"26",X"F1",
		X"2D",X"F1",X"2F",X"F1",X"34",X"F1",X"37",X"F1",X"4E",X"F1",X"A8",X"F1",X"2A",X"F2",X"C8",X"F2",
		X"74",X"F3",X"2B",X"F4",X"E7",X"F4",X"A5",X"F5",X"61",X"F6",X"1C",X"F7",X"D4",X"F7",X"88",X"F8",
		X"3A",X"F9",X"E4",X"F9",X"8B",X"FA",X"2E",X"FB",X"CB",X"FB",X"64",X"FC",X"FA",X"FC",X"8B",X"FD",
		X"16",X"FE",X"A1",X"FE",X"23",X"FF",X"A5",X"FF",X"20",X"00",X"9A",X"00",X"0E",X"01",X"7F",X"01",
		X"BE",X"01",X"C1",X"01",X"9F",X"01",X"63",X"01",X"18",X"01",X"C2",X"00",X"64",X"00",X"05",X"00",
		X"A5",X"FF",X"45",X"FF",X"E6",X"FE",X"88",X"FE",X"2A",X"FE",X"D0",X"FD",X"77",X"FD",X"22",X"FD",
		X"D0",X"FC",X"7F",X"FC",X"30",X"FC",X"E4",X"FB",X"9B",X"FB",X"54",X"FB",X"0E",X"FB",X"CC",X"FA",
		X"8A",X"FA",X"4D",X"FA",X"0E",X"FA",X"E2",X"F9",X"F4",X"F9",X"36",X"FA",X"95",X"FA",X"07",X"FB",
		X"88",X"FB",X"0D",X"FC",X"95",X"FC",X"20",X"FD",X"AB",X"FD",X"33",X"FE",X"BA",X"FE",X"3C",X"FF",
		X"BB",X"FF",X"38",X"00",X"B2",X"00",X"27",X"01",X"9A",X"01",X"09",X"02",X"74",X"02",X"DF",X"02",
		X"44",X"03",X"A7",X"03",X"06",X"04",X"62",X"04",X"BE",X"04",X"15",X"05",X"69",X"05",X"BA",X"05",
		X"08",X"06",X"56",X"06",X"A0",X"06",X"E9",X"06",X"2F",X"07",X"72",X"07",X"B4",X"07",X"F4",X"07",
		X"31",X"08",X"6B",X"08",X"A4",X"08",X"DC",X"08",X"12",X"09",X"46",X"09",X"78",X"09",X"A9",X"09",
		X"D7",X"09",X"06",X"0A",X"32",X"0A",X"5C",X"0A",X"84",X"0A",X"AD",X"0A",X"D2",X"0A",X"F8",X"0A",
		X"1A",X"0B",X"3C",X"0B",X"5C",X"0B",X"7E",X"0B",X"9B",X"0B",X"BA",X"0B",X"D5",X"0B",X"F2",X"0B",
		X"0B",X"0C",X"27",X"0C",X"3E",X"0C",X"55",X"0C",X"6C",X"0C",X"83",X"0C",X"95",X"0C",X"A9",X"0C",
		X"BC",X"0C",X"D1",X"0C",X"DD",X"0C",X"D5",X"0C",X"CE",X"0C",X"C6",X"0C",X"BE",X"0C",X"B6",X"0C",
		X"AF",X"0C",X"A7",X"0C",X"A1",X"0C",X"98",X"0C",X"91",X"0C",X"8A",X"0C",X"81",X"0C",X"7B",X"0C",
		X"72",X"0C",X"6C",X"0C",X"63",X"0C",X"5C",X"0C",X"55",X"0C",X"4E",X"0C",X"44",X"0C",X"3F",X"0C",
		X"37",X"0C",X"31",X"0C",X"29",X"0C",X"21",X"0C",X"19",X"0C",X"11",X"0C",X"0B",X"0C",X"04",X"0C",
		X"FB",X"0B",X"F5",X"0B",X"ED",X"0B",X"E7",X"0B",X"E0",X"0B",X"D8",X"0B",X"D1",X"0B",X"CA",X"0B",
		X"C2",X"0B",X"BD",X"0B",X"B3",X"0B",X"AF",X"0B",X"A4",X"0B",X"A4",X"0B",X"79",X"0B",X"C8",X"0A",
		X"0E",X"0A",X"54",X"09",X"9B",X"08",X"E5",X"07",X"33",X"07",X"85",X"06",X"DC",X"05",X"35",X"05",
		X"93",X"04",X"F8",X"03",X"60",X"03",X"CB",X"02",X"3C",X"02",X"B0",X"01",X"29",X"01",X"A4",X"00",
		X"26",X"00",X"AC",X"FF",X"33",X"FF",X"C0",X"FE",X"4F",X"FE",X"E2",X"FD",X"77",X"FD",X"11",X"FD",
		X"AD",X"FC",X"4E",X"FC",X"F0",X"FB",X"94",X"FB",X"3B",X"FB",X"E7",X"FA",X"94",X"FA",X"44",X"FA",
		X"F5",X"F9",X"AC",X"F9",X"62",X"F9",X"1D",X"F9",X"D9",X"F8",X"96",X"F8",X"57",X"F8",X"19",X"F8",
		X"DD",X"F7",X"A3",X"F7",X"6C",X"F7",X"37",X"F7",X"02",X"F7",X"CE",X"F6",X"9E",X"F6",X"6E",X"F6",
		X"43",X"F6",X"4A",X"F6",X"8B",X"F6",X"EC",X"F6",X"67",X"F7",X"EE",X"F7",X"7E",X"F8",X"11",X"F9",
		X"A7",X"F9",X"3E",X"FA",X"CF",X"FA",X"61",X"FB",X"EF",X"FB",X"7A",X"FC",X"04",X"FD",X"88",X"FD",
		X"08",X"FE",X"87",X"FE",X"FE",X"FE",X"74",X"FF",X"E6",X"FF",X"54",X"00",X"C1",X"00",X"28",X"01",
		X"8F",X"01",X"F0",X"01",X"4F",X"02",X"AD",X"02",X"F6",X"02",X"FE",X"02",X"D8",X"02",X"93",X"02",
		X"39",X"02",X"D5",X"01",X"6A",X"01",X"F8",X"00",X"87",X"00",X"16",X"00",X"A3",X"FF",X"35",X"FF",
		X"C8",X"FE",X"5D",X"FE",X"F5",X"FD",X"8F",X"FD",X"2F",X"FD",X"CE",X"FC",X"71",X"FC",X"19",X"FC",
		X"C1",X"FB",X"6B",X"FB",X"1A",X"FB",X"CC",X"FA",X"7E",X"FA",X"33",X"FA",X"EC",X"F9",X"A7",X"F9",
		X"61",X"F9",X"21",X"F9",X"E1",X"F8",X"A3",X"F8",X"69",X"F8",X"2E",X"F8",X"F8",X"F7",X"C1",X"F7",
		X"8C",X"F7",X"5B",X"F7",X"29",X"F7",X"FB",X"F6",X"CD",X"F6",X"A0",X"F6",X"77",X"F6",X"4E",X"F6",
		X"24",X"F6",X"00",X"F6",X"DA",X"F5",X"B7",X"F5",X"94",X"F5",X"73",X"F5",X"53",X"F5",X"34",X"F5",
		X"17",X"F5",X"FC",X"F4",X"DE",X"F4",X"CF",X"F4",X"FE",X"F4",X"5C",X"F5",X"D7",X"F5",X"67",X"F6",
		X"02",X"F7",X"A2",X"F7",X"48",X"F8",X"EC",X"F8",X"90",X"F9",X"30",X"FA",X"CE",X"FA",X"68",X"FB",
		X"01",X"FC",X"92",X"FC",X"21",X"FD",X"AE",X"FD",X"35",X"FE",X"B6",X"FE",X"38",X"FF",X"B2",X"FF",
		X"2A",X"00",X"9E",X"00",X"0F",X"01",X"7C",X"01",X"E7",X"01",X"4E",X"02",X"B3",X"02",X"F1",X"02",
		X"EF",X"02",X"C6",X"02",X"82",X"02",X"2C",X"02",X"CB",X"01",X"65",X"01",X"F8",X"00",X"8E",X"00",
		X"23",X"00",X"B9",X"FF",X"50",X"FF",X"EB",X"FE",X"85",X"FE",X"23",X"FE",X"C4",X"FD",X"68",X"FD",
		X"0D",X"FD",X"B8",X"FC",X"64",X"FC",X"11",X"FC",X"C2",X"FB",X"74",X"FB",X"2B",X"FB",X"E1",X"FA",
		X"9D",X"FA",X"57",X"FA",X"31",X"FA",X"4D",X"FA",X"90",X"FA",X"F0",X"FA",X"60",X"FB",X"DC",X"FB",
		X"5D",X"FC",X"E2",X"FC",X"67",X"FD",X"EC",X"FD",X"6C",X"FE",X"EB",X"FE",X"69",X"FF",X"E4",X"FF",
		X"5A",X"00",X"CE",X"00",X"3E",X"01",X"AC",X"01",X"15",X"02",X"7F",X"02",X"E1",X"02",X"41",X"03",
		X"A1",X"03",X"FB",X"03",X"54",X"04",X"A9",X"04",X"FC",X"04",X"48",X"05",X"5D",X"05",X"3B",X"05",
		X"F7",X"04",X"9B",X"04",X"31",X"04",X"BE",X"03",X"46",X"03",X"CC",X"02",X"52",X"02",X"DA",X"01",
		X"62",X"01",X"EE",X"00",X"7B",X"00",X"0B",X"00",X"A0",X"FF",X"35",X"FF",X"CE",X"FE",X"6A",X"FE",
		X"08",X"FE",X"AA",X"FD",X"4F",X"FD",X"F6",X"FC",X"A1",X"FC",X"4E",X"FC",X"FD",X"FB",X"AF",X"FB",
		X"64",X"FB",X"18",X"FB",X"D2",X"FA",X"8D",X"FA",X"4B",X"FA",X"0A",X"FA",X"CD",X"F9",X"91",X"F9",
		X"55",X"F9",X"1C",X"F9",X"E4",X"F8",X"B1",X"F8",X"7C",X"F8",X"4C",X"F8",X"1B",X"F8",X"EC",X"F7",
		X"BF",X"F7",X"95",X"F7",X"6B",X"F7",X"41",X"F7",X"1B",X"F7",X"F6",X"F6",X"D1",X"F6",X"AD",X"F6",
		X"8D",X"F6",X"6B",X"F6",X"4B",X"F6",X"2D",X"F6",X"0F",X"F6",X"24",X"F6",X"72",X"F6",X"E2",X"F6",
		X"69",X"F7",X"FE",X"F7",X"9C",X"F8",X"3E",X"F9",X"E0",X"F9",X"81",X"FA",X"21",X"FB",X"BE",X"FB",
		X"59",X"FC",X"ED",X"FC",X"81",X"FD",X"0F",X"FE",X"9A",X"FE",X"22",X"FF",X"A5",X"FF",X"23",X"00",
		X"9D",X"00",X"17",X"01",X"8A",X"01",X"FC",X"01",X"69",X"02",X"D3",X"02",X"39",X"03",X"9C",X"03",
		X"FD",X"03",X"5A",X"04",X"B4",X"04",X"0E",X"05",X"63",X"05",X"B5",X"05",X"04",X"06",X"51",X"06",
		X"9D",X"06",X"E5",X"06",X"2C",X"07",X"71",X"07",X"B3",X"07",X"F3",X"07",X"30",X"08",X"6D",X"08",
		X"A7",X"08",X"E0",X"08",X"15",X"09",X"48",X"09",X"7D",X"09",X"AC",X"09",X"DD",X"09",X"0B",X"0A",
		X"37",X"0A",X"61",X"0A",X"8A",X"0A",X"B3",X"0A",X"D8",X"0A",X"FF",X"0A",X"23",X"0B",X"45",X"0B",
		X"66",X"0B",X"86",X"0B",X"A6",X"0B",X"C3",X"0B",X"E0",X"0B",X"FB",X"0B",X"17",X"0C",X"31",X"0C",
		X"49",X"0C",X"60",X"0C",X"76",X"0C",X"8E",X"0C",X"A1",X"0C",X"B7",X"0C",X"CB",X"0C",X"DD",X"0C",
		X"EE",X"0C",X"ED",X"0C",X"E4",X"0C",X"DD",X"0C",X"D5",X"0C",X"CE",X"0C",X"C7",X"0C",X"BD",X"0C",
		X"B5",X"0C",X"AE",X"0C",X"A7",X"0C",X"A0",X"0C",X"96",X"0C",X"90",X"0C",X"88",X"0C",X"80",X"0C",
		X"78",X"0C",X"71",X"0C",X"69",X"0C",X"62",X"0C",X"5B",X"0C",X"54",X"0C",X"4D",X"0C",X"45",X"0C",
		X"3E",X"0C",X"36",X"0C",X"2E",X"0C",X"27",X"0C",X"20",X"0C",X"18",X"0C",X"11",X"0C",X"0A",X"0C",
		X"03",X"0C",X"FC",X"0B",X"F3",X"0B",X"EB",X"0B",X"E6",X"0B",X"DE",X"0B",X"D7",X"0B",X"CF",X"0B",
		X"C9",X"0B",X"C1",X"0B",X"B9",X"0B",X"B4",X"0B",X"AC",X"0B",X"A4",X"0B",X"9E",X"0B",X"96",X"0B",
		X"8F",X"0B",X"87",X"0B",X"81",X"0B",X"7A",X"0B",X"73",X"0B",X"6D",X"0B",X"65",X"0B",X"5F",X"0B",
		X"58",X"0B",X"50",X"0B",X"48",X"0B",X"42",X"0B",X"39",X"0B",X"36",X"0B",X"2D",X"0B",X"27",X"0B",
		X"1F",X"0B",X"1B",X"0B",X"10",X"0B",X"12",X"0B",X"AF",X"0A",X"E9",X"09",X"31",X"09",X"74",X"08",
		X"BC",X"07",X"05",X"07",X"57",X"06",X"A8",X"05",X"01",X"05",X"5D",X"04",X"BE",X"03",X"21",X"03",
		X"8E",X"02",X"FA",X"01",X"6E",X"01",X"E5",X"00",X"5F",X"00",X"DF",X"FF",X"62",X"FF",X"E7",X"FE",
		X"71",X"FE",X"FE",X"FD",X"90",X"FD",X"24",X"FD",X"BB",X"FC",X"57",X"FC",X"F6",X"FB",X"96",X"FB",
		X"39",X"FB",X"E0",X"FA",X"8B",X"FA",X"37",X"FA",X"E5",X"F9",X"97",X"F9",X"4A",X"F9",X"01",X"F9",
		X"BB",X"F8",X"74",X"F8",X"32",X"F8",X"F1",X"F7",X"B1",X"F7",X"76",X"F7",X"3A",X"F7",X"02",X"F7",
		X"CA",X"F6",X"97",X"F6",X"64",X"F6",X"31",X"F6",X"03",X"F6",X"D7",X"F5",X"DE",X"F5",X"1E",X"F6",
		X"80",X"F6",X"F9",X"F6",X"80",X"F7",X"10",X"F8",X"A3",X"F8",X"3A",X"F9",X"CD",X"F9",X"62",X"FA",
		X"F1",X"FA",X"80",X"FB",X"0A",X"FC",X"92",X"FC",X"17",X"FD",X"96",X"FD",X"13",X"FE",X"8C",X"FE",
		X"01",X"FF",X"73",X"FF",X"E2",X"FF",X"4D",X"00",X"B4",X"00",X"19",X"01",X"7C",X"01",X"DB",X"01",
		X"37",X"02",X"91",X"02",X"E6",X"02",X"3A",X"03",X"8C",X"03",X"DC",X"03",X"28",X"04",X"72",X"04",
		X"B9",X"04",X"01",X"05",X"42",X"05",X"84",X"05",X"C4",X"05",X"00",X"06",X"3D",X"06",X"75",X"06",
		X"AD",X"06",X"E3",X"06",X"16",X"07",X"49",X"07",X"79",X"07",X"A8",X"07",X"D6",X"07",X"02",X"08",
		X"2D",X"08",X"56",X"08",X"7D",X"08",X"A4",X"08",X"C9",X"08",X"C0",X"08",X"7B",X"08",X"14",X"08",
		X"97",X"07",X"09",X"07",X"72",X"06",X"D7",X"05",X"3B",X"05",X"9E",X"04",X"04",X"04",X"6C",X"03",
		X"D8",X"02",X"48",X"02",X"BA",X"01",X"30",X"01",X"A9",X"00",X"28",X"00",X"AB",X"FF",X"2F",X"FF",
		X"B9",X"FE",X"44",X"FE",X"D5",X"FD",X"69",X"FD",X"00",X"FD",X"9A",X"FC",X"35",X"FC",X"D5",X"FB",
		X"79",X"FB",X"1F",X"FB",X"C6",X"FA",X"71",X"FA",X"20",X"FA",X"D0",X"F9",X"84",X"F9",X"39",X"F9",
		X"F0",X"F8",X"AA",X"F8",X"66",X"F8",X"26",X"F8",X"E7",X"F7",X"A9",X"F7",X"6E",X"F7",X"33",X"F7",
		X"FB",X"F6",X"C6",X"F6",X"93",X"F6",X"60",X"F6",X"30",X"F6",X"01",X"F6",X"D3",X"F5",X"A8",X"F5",
		X"7E",X"F5",X"55",X"F5",X"2E",X"F5",X"07",X"F5",X"E3",X"F4",X"BF",X"F4",X"9B",X"F4",X"7C",X"F4",
		X"5D",X"F4",X"3D",X"F4",X"1F",X"F4",X"03",X"F4",X"E7",X"F3",X"CE",X"F3",X"B5",X"F3",X"9E",X"F3",
		X"85",X"F3",X"70",X"F3",X"5B",X"F3",X"44",X"F3",X"32",X"F3",X"1E",X"F3",X"0C",X"F3",X"FC",X"F2",
		X"E9",X"F2",X"D9",X"F2",X"CA",X"F2",X"BC",X"F2",X"AE",X"F2",X"A1",X"F2",X"93",X"F2",X"89",X"F2",
		X"7C",X"F2",X"71",X"F2",X"67",X"F2",X"5D",X"F2",X"55",X"F2",X"4D",X"F2",X"44",X"F2",X"3D",X"F2",
		X"35",X"F2",X"2F",X"F2",X"28",X"F2",X"23",X"F2",X"1D",X"F2",X"18",X"F2",X"14",X"F2",X"0F",X"F2",
		X"0B",X"F2",X"09",X"F2",X"05",X"F2",X"03",X"F2",X"02",X"F2",X"FE",X"F1",X"FC",X"F1",X"FB",X"F1",
		X"FA",X"F1",X"F9",X"F1",X"FC",X"F1",X"36",X"F2",X"A5",X"F2",X"35",X"F3",X"D8",X"F3",X"86",X"F4",
		X"3D",X"F5",X"F7",X"F5",X"B1",X"F6",X"67",X"F7",X"1C",X"F8",X"CE",X"F8",X"7D",X"F9",X"27",X"FA",
		X"CB",X"FA",X"6C",X"FB",X"09",X"FC",X"A1",X"FC",X"34",X"FD",X"C3",X"FD",X"4F",X"FE",X"D7",X"FE",
		X"59",X"FF",X"D9",X"FF",X"53",X"00",X"CB",X"00",X"3F",X"01",X"B1",X"01",X"1C",X"02",X"87",X"02",
		X"EE",X"02",X"51",X"03",X"B3",X"03",X"0F",X"04",X"69",X"04",X"C0",X"04",X"17",X"05",X"6A",X"05",
		X"B9",X"05",X"08",X"06",X"52",X"06",X"9B",X"06",X"E1",X"06",X"26",X"07",X"66",X"07",X"A8",X"07",
		X"E5",X"07",X"21",X"08",X"5A",X"08",X"92",X"08",X"CA",X"08",X"FE",X"08",X"30",X"09",X"63",X"09",
		X"90",X"09",X"BD",X"09",X"B7",X"09",X"78",X"09",X"16",X"09",X"9E",X"08",X"17",X"08",X"87",X"07",
		X"F2",X"06",X"5D",X"06",X"C9",X"05",X"34",X"05",X"A3",X"04",X"15",X"04",X"8B",X"03",X"02",X"03",
		X"7E",X"02",X"FD",X"01",X"80",X"01",X"08",X"01",X"91",X"00",X"21",X"00",X"B1",X"FF",X"46",X"FF",
		X"DD",X"FE",X"79",X"FE",X"17",X"FE",X"B7",X"FD",X"5B",X"FD",X"02",X"FD",X"AA",X"FC",X"57",X"FC",
		X"05",X"FC",X"B7",X"FB",X"6A",X"FB",X"21",X"FB",X"D9",X"FA",X"91",X"FA",X"4F",X"FA",X"0F",X"FA",
		X"CF",X"F9",X"92",X"F9",X"55",X"F9",X"1C",X"F9",X"E6",X"F8",X"B0",X"F8",X"7D",X"F8",X"49",X"F8",
		X"19",X"F8",X"EC",X"F7",X"BD",X"F7",X"92",X"F7",X"66",X"F7",X"3F",X"F7",X"17",X"F7",X"EF",X"F6",
		X"CB",X"F6",X"D2",X"F6",X"15",X"F7",X"7A",X"F7",X"FA",X"F7",X"86",X"F8",X"1D",X"F9",X"B9",X"F9",
		X"54",X"FA",X"F1",X"FA",X"8E",X"FB",X"24",X"FC",X"B8",X"FC",X"4B",X"FD",X"DA",X"FD",X"64",X"FE",
		X"EA",X"FE",X"6D",X"FF",X"EB",X"FF",X"66",X"00",X"DD",X"00",X"52",X"01",X"C3",X"01",X"2F",X"02",
		X"99",X"02",X"00",X"03",X"62",X"03",X"C5",X"03",X"18",X"04",X"2C",X"04",X"0D",X"04",X"D0",X"03",
		X"7C",X"03",X"1C",X"03",X"B4",X"02",X"47",X"02",X"D7",X"01",X"68",X"01",X"F9",X"00",X"8D",X"00",
		X"21",X"00",X"BA",X"FF",X"53",X"FF",X"EF",X"FE",X"8F",X"FE",X"31",X"FE",X"D4",X"FD",X"7C",X"FD",
		X"27",X"FD",X"D4",X"FC",X"84",X"FC",X"36",X"FC",X"EA",X"FB",X"A0",X"FB",X"59",X"FB",X"13",X"FB",
		X"D1",X"FA",X"90",X"FA",X"53",X"FA",X"15",X"FA",X"DA",X"F9",X"A0",X"F9",X"6A",X"F9",X"34",X"F9",
		X"00",X"F9",X"D0",X"F8",X"9E",X"F8",X"70",X"F8",X"43",X"F8",X"17",X"F8",X"EE",X"F7",X"C5",X"F7",
		X"9D",X"F7",X"77",X"F7",X"52",X"F7",X"2E",X"F7",X"0D",X"F7",X"EB",X"F6",X"CB",X"F6",X"AE",X"F6",
		X"8E",X"F6",X"72",X"F6",X"56",X"F6",X"42",X"F6",X"67",X"F6",X"C0",X"F6",X"39",X"F7",X"C7",X"F7",
		X"5F",X"F8",X"00",X"F9",X"A3",X"F9",X"48",X"FA",X"EC",X"FA",X"8D",X"FB",X"2B",X"FC",X"C7",X"FC",
		X"5E",X"FD",X"F0",X"FD",X"81",X"FE",X"0A",X"FF",X"94",X"FF",X"17",X"00",X"95",X"00",X"11",X"01",
		X"8B",X"01",X"FE",X"01",X"70",X"02",X"DE",X"02",X"47",X"03",X"B1",X"03",X"13",X"04",X"75",X"04",
		X"D2",X"04",X"2D",X"05",X"87",X"05",X"DC",X"05",X"2F",X"06",X"80",X"06",X"CC",X"06",X"18",X"07",
		X"5F",X"07",X"A7",X"07",X"EC",X"07",X"2F",X"08",X"6D",X"08",X"AC",X"08",X"EA",X"08",X"22",X"09",
		X"5B",X"09",X"90",X"09",X"C5",X"09",X"F8",X"09",X"28",X"0A",X"5A",X"0A",X"87",X"0A",X"B3",X"0A",
		X"DE",X"0A",X"07",X"0B",X"2E",X"0B",X"54",X"0B",X"79",X"0B",X"9E",X"0B",X"C2",X"0B",X"E3",X"0B",
		X"03",X"0C",X"21",X"0C",X"3F",X"0C",X"5C",X"0C",X"77",X"0C",X"93",X"0C",X"AB",X"0C",X"C7",X"0C",
		X"DC",X"0C",X"F4",X"0C",X"09",X"0D",X"1F",X"0D",X"32",X"0D",X"45",X"0D",X"57",X"0D",X"6B",X"0D",
		X"70",X"0D",X"68",X"0D",X"60",X"0D",X"58",X"0D",X"4F",X"0D",X"4A",X"0D",X"3E",X"0D",X"3B",X"0D",
		X"0A",X"0D",X"7D",X"0C",X"E2",X"0B",X"39",X"0B",X"8C",X"0A",X"DB",X"09",X"2D",X"09",X"7E",X"08",
		X"D4",X"07",X"2E",X"07",X"89",X"06",X"EA",X"05",X"4E",X"05",X"B5",X"04",X"23",X"04",X"94",X"03",
		X"09",X"03",X"82",X"02",X"FF",X"01",X"81",X"01",X"06",X"01",X"8E",X"00",X"1B",X"00",X"AA",X"FF",
		X"3E",X"FF",X"D4",X"FE",X"9B",X"FE",X"9F",X"FE",X"C8",X"FE",X"0B",X"FF",X"5C",X"FF",X"B9",X"FF",
		X"1B",X"00",X"80",X"00",X"E8",X"00",X"4D",X"01",X"B4",X"01",X"19",X"02",X"79",X"02",X"D9",X"02",
		X"36",X"03",X"91",X"03",X"E8",X"03",X"3D",X"04",X"90",X"04",X"E0",X"04",X"2E",X"05",X"7A",X"05",
		X"C3",X"05",X"0A",X"06",X"4E",X"06",X"91",X"06",X"D3",X"06",X"03",X"07",X"F6",X"06",X"B9",X"06",
		X"5C",X"06",X"EB",X"05",X"70",X"05",X"ED",X"04",X"65",X"04",X"DF",X"03",X"56",X"03",X"D1",X"02",
		X"4E",X"02",X"CD",X"01",X"4F",X"01",X"D5",X"00",X"5D",X"00",X"EA",X"FF",X"79",X"FF",X"0C",X"FF",
		X"A1",X"FE",X"39",X"FE",X"D5",X"FD",X"74",X"FD",X"16",X"FD",X"BC",X"FC",X"62",X"FC",X"0E",X"FC",
		X"B9",X"FB",X"90",X"FB",X"A2",X"FB",X"DC",X"FB",X"32",X"FC",X"96",X"FC",X"07",X"FD",X"79",X"FD",
		X"F3",X"FD",X"6C",X"FE",X"E3",X"FE",X"59",X"FF",X"CE",X"FF",X"40",X"00",X"AF",X"00",X"1C",X"01",
		X"85",X"01",X"EB",X"01",X"4F",X"02",X"AF",X"02",X"0E",X"03",X"6A",X"03",X"C1",X"03",X"17",X"04",
		X"6A",X"04",X"BA",X"04",X"09",X"05",X"55",X"05",X"9B",X"05",X"E4",X"05",X"28",X"06",X"6B",X"06",
		X"AA",X"06",X"E9",X"06",X"26",X"07",X"61",X"07",X"98",X"07",X"CF",X"07",X"05",X"08",X"38",X"08",
		X"69",X"08",X"9A",X"08",X"C7",X"08",X"F4",X"08",X"20",X"09",X"4A",X"09",X"72",X"09",X"99",X"09",
		X"BF",X"09",X"E4",X"09",X"05",X"0A",X"29",X"0A",X"49",X"0A",X"69",X"0A",X"86",X"0A",X"A5",X"0A",
		X"A3",X"0A",X"61",X"0A",X"FC",X"09",X"79",X"09",X"E8",X"08",X"4B",X"08",X"AA",X"07",X"07",X"07",
		X"66",X"06",X"C4",X"05",X"25",X"05",X"89",X"04",X"F3",X"03",X"5D",X"03",X"CE",X"02",X"43",X"02",
		X"BB",X"01",X"35",X"01",X"B4",X"00",X"3A",X"00",X"C1",X"FF",X"4A",X"FF",X"D8",X"FE",X"6A",X"FE",
		X"FF",X"FD",X"98",X"FD",X"32",X"FD",X"D6",X"FC",X"B1",X"FC",X"C4",X"FC",X"F8",X"FC",X"46",X"FD",
		X"A2",X"FD",X"05",X"FE",X"70",X"FE",X"DD",X"FE",X"49",X"FF",X"B4",X"FF",X"1F",X"00",X"88",X"00",
		X"EF",X"00",X"54",X"01",X"B5",X"01",X"14",X"02",X"6F",X"02",X"C9",X"02",X"20",X"03",X"74",X"03",
		X"C5",X"03",X"16",X"04",X"62",X"04",X"AC",X"04",X"F5",X"04",X"3C",X"05",X"80",X"05",X"C2",X"05",
		X"00",X"06",X"3F",X"06",X"79",X"06",X"B2",X"06",X"EB",X"06",X"21",X"07",X"56",X"07",X"89",X"07",
		X"B9",X"07",X"E7",X"07",X"15",X"08",X"43",X"08",X"6D",X"08",X"97",X"08",X"BE",X"08",X"E6",X"08",
		X"0A",X"09",X"30",X"09",X"53",X"09",X"73",X"09",X"93",X"09",X"B3",X"09",X"D1",X"09",X"EE",X"09",
		X"0B",X"0A",X"27",X"0A",X"2F",X"0A",X"F8",X"09",X"95",X"09",X"17",X"09",X"85",X"08",X"E9",X"07",
		X"48",X"07",X"A4",X"06",X"FE",X"05",X"5C",X"05",X"BB",X"04",X"1D",X"04",X"82",X"03",X"EC",X"02",
		X"5A",X"02",X"CB",X"01",X"41",X"01",X"BA",X"00",X"38",X"00",X"BB",X"FF",X"3F",X"FF",X"C6",X"FE",
		X"53",X"FE",X"E3",X"FD",X"75",X"FD",X"0B",X"FD",X"A6",X"FC",X"43",X"FC",X"0D",X"FC",X"15",X"FC",
		X"43",X"FC",X"8B",X"FC",X"E3",X"FC",X"44",X"FD",X"AD",X"FD",X"18",X"FE",X"84",X"FE",X"F0",X"FE",
		X"5A",X"FF",X"C3",X"FF",X"28",X"00",X"8D",X"00",X"EF",X"00",X"4E",X"01",X"AC",X"01",X"05",X"02",
		X"5B",X"02",X"B1",X"02",X"03",X"03",X"53",X"03",X"9F",X"03",X"EB",X"03",X"33",X"04",X"79",X"04",
		X"BE",X"04",X"F5",X"04",X"EB",X"04",X"B3",X"04",X"5B",X"04",X"F1",X"03",X"77",X"03",X"F8",X"02",
		X"74",X"02",X"EE",X"01",X"69",X"01",X"E7",X"00",X"67",X"00",X"E9",X"FF",X"6F",X"FF",X"F6",X"FE",
		X"81",X"FE",X"0E",X"FE",X"A0",X"FD",X"35",X"FD",X"CD",X"FC",X"68",X"FC",X"06",X"FC",X"A8",X"FB",
		X"4C",X"FB",X"F2",X"FA",X"9B",X"FA",X"48",X"FA",X"F8",X"F9",X"A8",X"F9",X"5D",X"F9",X"15",X"F9",
		X"CD",X"F8",X"86",X"F8",X"43",X"F8",X"02",X"F8",X"C3",X"F7",X"87",X"F7",X"4B",X"F7",X"13",X"F7",
		X"DD",X"F6",X"A7",X"F6",X"74",X"F6",X"42",X"F6",X"14",X"F6",X"E4",X"F5",X"B8",X"F5",X"8C",X"F5",
		X"63",X"F5",X"3A",X"F5",X"13",X"F5",X"ED",X"F4",X"C9",X"F4",X"A6",X"F4",X"85",X"F4",X"64",X"F4",
		X"4C",X"F4",X"6D",X"F4",X"C2",X"F4",X"35",X"F5",X"C0",X"F5",X"54",X"F6",X"F3",X"F6",X"93",X"F7",
		X"34",X"F8",X"D5",X"F8",X"72",X"F9",X"0D",X"FA",X"A6",X"FA",X"3A",X"FB",X"CA",X"FB",X"56",X"FC",
		X"E0",X"FC",X"64",X"FD",X"E6",X"FD",X"63",X"FE",X"DC",X"FE",X"52",X"FF",X"C5",X"FF",X"35",X"00",
		X"A0",X"00",X"08",X"01",X"6E",X"01",X"D3",X"01",X"15",X"02",X"18",X"02",X"F1",X"01",X"AD",X"01",
		X"5A",X"01",X"F7",X"00",X"8E",X"00",X"23",X"00",X"B8",X"FF",X"4A",X"FF",X"DF",X"FE",X"74",X"FE",
		X"0C",X"FE",X"A7",X"FD",X"44",X"FD",X"E4",X"FC",X"87",X"FC",X"2A",X"FC",X"D2",X"FB",X"7D",X"FB",
		X"29",X"FB",X"D9",X"FA",X"8C",X"FA",X"41",X"FA",X"F8",X"F9",X"B1",X"F9",X"6C",X"F9",X"29",X"F9",
		X"EA",X"F8",X"A9",X"F8",X"6E",X"F8",X"33",X"F8",X"FA",X"F7",X"C3",X"F7",X"8F",X"F7",X"5C",X"F7",
		X"2C",X"F7",X"FC",X"F6",X"CC",X"F6",X"A0",X"F6",X"74",X"F6",X"4C",X"F6",X"23",X"F6",X"FC",X"F5",
		X"D5",X"F5",X"B2",X"F5",X"90",X"F5",X"6E",X"F5",X"4D",X"F5",X"2E",X"F5",X"10",X"F5",X"F3",X"F4",
		X"D5",X"F4",X"BD",X"F4",X"A1",X"F4",X"9B",X"F4",X"D8",X"F4",X"3C",X"F5",X"BE",X"F5",X"51",X"F6",
		X"EF",X"F6",X"92",X"F7",X"36",X"F8",X"DD",X"F8",X"81",X"F9",X"23",X"FA",X"C0",X"FA",X"5C",X"FB",
		X"F3",X"FB",X"87",X"FC",X"15",X"FD",X"A0",X"FD",X"28",X"FE",X"AB",X"FE",X"2A",X"FF",X"A6",X"FF",
		X"1E",X"00",X"92",X"00",X"03",X"01",X"70",X"01",X"DB",X"01",X"41",X"02",X"A6",X"02",X"08",X"03",
		X"65",X"03",X"C0",X"03",X"18",X"04",X"6E",X"04",X"C2",X"04",X"11",X"05",X"5F",X"05",X"AB",X"05",
		X"F5",X"05",X"3A",X"06",X"80",X"06",X"C2",X"06",X"03",X"07",X"41",X"07",X"7D",X"07",X"B7",X"07",
		X"F0",X"07",X"25",X"08",X"5B",X"08",X"8E",X"08",X"C0",X"08",X"EF",X"08",X"1E",X"09",X"49",X"09",
		X"76",X"09",X"9F",X"09",X"C6",X"09",X"EF",X"09",X"15",X"0A",X"39",X"0A",X"5A",X"0A",X"7C",X"0A",
		X"9D",X"0A",X"BC",X"0A",X"DA",X"0A",X"F8",X"0A",X"14",X"0B",X"2F",X"0B",X"4A",X"0B",X"62",X"0B",
		X"7B",X"0B",X"93",X"0B",X"A8",X"0B",X"BD",X"0B",X"D3",X"0B",X"E5",X"0B",X"F8",X"0B",X"0D",X"0C",
		X"12",X"0C",X"0B",X"0C",X"04",X"0C",X"FC",X"0B",X"F4",X"0B",X"EC",X"0B",X"E5",X"0B",X"DE",X"0B",
		X"D5",X"0B",X"D0",X"0B",X"C7",X"0B",X"C0",X"0B",X"B9",X"0B",X"B2",X"0B",X"AB",X"0B",X"A4",X"0B",
		X"9E",X"0B",X"97",X"0B",X"8F",X"0B",X"87",X"0B",X"81",X"0B",X"7A",X"0B",X"72",X"0B",X"6C",X"0B",
		X"65",X"0B",X"5E",X"0B",X"56",X"0B",X"50",X"0B",X"47",X"0B",X"42",X"0B",X"3A",X"0B",X"34",X"0B",
		X"2C",X"0B",X"27",X"0B",X"1D",X"0B",X"18",X"0B",X"0D",X"0B",X"0E",X"0B",X"A5",X"0A",X"E6",X"09",
		X"32",X"09",X"75",X"08",X"C2",X"07",X"0B",X"07",X"5D",X"06",X"AF",X"05",X"09",X"05",X"64",X"04",
		X"C6",X"03",X"2A",X"03",X"93",X"02",X"02",X"02",X"74",X"01",X"E9",X"00",X"64",X"00",X"E2",X"FF",
		X"64",X"FF",X"EA",X"FE",X"74",X"FE",X"01",X"FE",X"92",X"FD",X"27",X"FD",X"BE",X"FC",X"58",X"FC",
		X"F7",X"FB",X"96",X"FB",X"3A",X"FB",X"DF",X"FA",X"89",X"FA",X"35",X"FA",X"E5",X"F9",X"96",X"F9",
		X"49",X"F9",X"FF",X"F8",X"B7",X"F8",X"73",X"F8",X"2F",X"F8",X"ED",X"F7",X"B0",X"F7",X"73",X"F7",
		X"36",X"F7",X"FE",X"F6",X"C8",X"F6",X"93",X"F6",X"5E",X"F6",X"2C",X"F6",X"FB",X"F5",X"CE",X"F5",
		X"A1",X"F5",X"75",X"F5",X"4C",X"F5",X"23",X"F5",X"FB",X"F4",X"D7",X"F4",X"B1",X"F4",X"8E",X"F4",
		X"6D",X"F4",X"4C",X"F4",X"2E",X"F4",X"0D",X"F4",X"F2",X"F3",X"D5",X"F3",X"BA",X"F3",X"9F",X"F3",
		X"87",X"F3",X"6F",X"F3",X"57",X"F3",X"42",X"F3",X"2D",X"F3",X"17",X"F3",X"05",X"F3",X"F2",X"F2",
		X"E0",X"F2",X"CE",X"F2",X"BF",X"F2",X"AC",X"F2",X"B7",X"F2",X"FF",X"F2",X"6F",X"F3",X"FB",X"F3",
		X"98",X"F4",X"3E",X"F5",X"EB",X"F5",X"99",X"F6",X"46",X"F7",X"F2",X"F7",X"9B",X"F8",X"3F",X"F9",
		X"E2",X"F9",X"80",X"FA",X"1A",X"FB",X"B0",X"FB",X"40",X"FC",X"CD",X"FC",X"57",X"FD",X"DD",X"FD",
		X"5D",X"FE",X"DB",X"FE",X"55",X"FF",X"CB",X"FF",X"3D",X"00",X"AD",X"00",X"17",X"01",X"7E",X"01",
		X"B0",X"01",X"A6",X"01",X"7C",X"01",X"36",X"01",X"E3",X"00",X"84",X"00",X"21",X"00",X"BB",X"FF",
		X"53",X"FF",X"EB",X"FE",X"87",X"FE",X"23",X"FE",X"BE",X"FD",X"5F",X"FD",X"02",X"FD",X"A7",X"FC",
		X"4F",X"FC",X"F9",X"FB",X"A7",X"FB",X"54",X"FB",X"08",X"FB",X"BD",X"FA",X"72",X"FA",X"2D",X"FA",
		X"E6",X"F9",X"A3",X"F9",X"63",X"F9",X"52",X"F9",X"7C",X"F9",X"CA",X"F9",X"32",X"FA",X"A7",X"FA",
		X"26",X"FB",X"A9",X"FB",X"31",X"FC",X"B9",X"FC",X"3E",X"FD",X"C2",X"FD",X"42",X"FE",X"C2",X"FE",
		X"3C",X"FF",X"B3",X"FF",X"28",X"00",X"99",X"00",X"09",X"01",X"73",X"01",X"DB",X"01",X"41",X"02",
		X"A3",X"02",X"01",X"03",X"5C",X"03",X"B7",X"03",X"0C",X"04",X"61",X"04",X"A5",X"04",X"AB",X"04",
		X"7F",X"04",X"36",X"04",X"D6",X"03",X"6C",X"03",X"F8",X"02",X"80",X"02",X"07",X"02",X"8F",X"01",
		X"17",X"01",X"A0",X"00",X"2E",X"00",X"BC",X"FF",X"4F",X"FF",X"E5",X"FE",X"7C",X"FE",X"16",X"FE",
		X"B3",X"FD",X"55",X"FD",X"F6",X"FC",X"9F",X"FC",X"47",X"FC",X"F3",X"FB",X"A0",X"FB",X"51",X"FB",
		X"05",X"FB",X"B9",X"FA",X"97",X"FA",X"B3",X"FA",X"F3",X"FA",X"50",X"FB",X"BA",X"FB",X"31",X"FC",
		X"AE",X"FC",X"2E",X"FD",X"AC",X"FD",X"2B",X"FE",X"A9",X"FE",X"23",X"FF",X"9C",X"FF",X"10",X"00",
		X"83",X"00",X"F1",X"00",X"5E",X"01",X"C7",X"01",X"2B",X"02",X"8F",X"02",X"ED",X"02",X"4B",X"03",
		X"A6",X"03",X"FC",X"03",X"51",X"04",X"A4",X"04",X"F5",X"04",X"40",X"05",X"8B",X"05",X"D4",X"05",
		X"19",X"06",X"5D",X"06",X"9F",X"06",X"DF",X"06",X"1D",X"07",X"58",X"07",X"93",X"07",X"CB",X"07",
		X"00",X"08",X"36",X"08",X"67",X"08",X"99",X"08",X"C7",X"08",X"F5",X"08",X"21",X"09",X"4B",X"09",
		X"75",X"09",X"9E",X"09",X"C3",X"09",X"E8",X"09",X"0D",X"0A",X"2F",X"0A",X"50",X"0A",X"6F",X"0A",
		X"93",X"0A",X"91",X"0A",X"54",X"0A",X"EF",X"09",X"6F",X"09",X"DF",X"08",X"45",X"08",X"A5",X"07",
		X"03",X"07",X"63",X"06",X"C5",X"05",X"26",X"05",X"8C",X"04",X"F5",X"03",X"64",X"03",X"D4",X"02",
		X"48",X"02",X"C2",X"01",X"3D",X"01",X"BE",X"00",X"41",X"00",X"CB",X"FF",X"56",X"FF",X"E5",X"FE",
		X"77",X"FE",X"0D",X"FE",X"A5",X"FD",X"42",X"FD",X"E2",X"FC",X"83",X"FC",X"28",X"FC",X"D1",X"FB",
		X"79",X"FB",X"26",X"FB",X"D7",X"FA",X"89",X"FA",X"3E",X"FA",X"F4",X"F9",X"AD",X"F9",X"69",X"F9",
		X"27",X"F9",X"E5",X"F8",X"A7",X"F8",X"6D",X"F8",X"32",X"F8",X"F9",X"F7",X"C2",X"F7",X"8F",X"F7",
		X"5C",X"F7",X"2A",X"F7",X"F9",X"F6",X"CB",X"F6",X"9F",X"F6",X"74",X"F6",X"4A",X"F6",X"23",X"F6",
		X"FB",X"F5",X"D6",X"F5",X"B3",X"F5",X"91",X"F5",X"6E",X"F5",X"4D",X"F5",X"2F",X"F5",X"10",X"F5",
		X"F3",X"F4",X"D7",X"F4",X"BB",X"F4",X"A3",X"F4",X"89",X"F4",X"71",X"F4",X"5A",X"F4",X"43",X"F4",
		X"2F",X"F4",X"1B",X"F4",X"07",X"F4",X"F3",X"F3",X"E3",X"F3",X"D1",X"F3",X"C1",X"F3",X"B0",X"F3",
		X"A2",X"F3",X"93",X"F3",X"85",X"F3",X"79",X"F3",X"9D",X"F3",X"FA",X"F3",X"79",X"F4",X"0E",X"F5",
		X"B4",X"F5",X"5E",X"F6",X"0C",X"F7",X"BC",X"F7",X"6B",X"F8",X"17",X"F9",X"C0",X"F9",X"66",X"FA",
		X"07",X"FB",X"A4",X"FB",X"3F",X"FC",X"D3",X"FC",X"64",X"FD",X"F1",X"FD",X"79",X"FE",X"FF",X"FE",
		X"80",X"FF",X"FC",X"FF",X"75",X"00",X"EA",X"00",X"5D",X"01",X"C9",X"01",X"38",X"02",X"91",X"02",
		X"A7",X"02",X"90",X"02",X"5A",X"02",X"0F",X"02",X"B7",X"01",X"57",X"01",X"F1",X"00",X"8B",X"00",
		X"24",X"00",X"BD",X"FF",X"5A",X"FF",X"F6",X"FE",X"95",X"FE",X"36",X"FE",X"DB",X"FD",X"81",X"FD",
		X"2A",X"FD",X"D7",X"FC",X"85",X"FC",X"33",X"FC",X"E7",X"FB",X"9D",X"FB",X"53",X"FB",X"0E",X"FB",
		X"CA",X"FA",X"88",X"FA",X"48",X"FA",X"33",X"FA",X"5B",X"FA",X"A8",X"FA",X"10",X"FB",X"84",X"FB",
		X"05",X"FC",X"89",X"FC",X"13",X"FD",X"99",X"FD",X"20",X"FE",X"A4",X"FE",X"26",X"FF",X"A5",X"FF",
		X"21",X"00",X"99",X"00",X"0D",X"01",X"81",X"01",X"F1",X"01",X"5C",X"02",X"C3",X"02",X"28",X"03",
		X"8B",X"03",X"EA",X"03",X"46",X"04",X"A1",X"04",X"F8",X"04",X"4A",X"05",X"9D",X"05",X"EC",X"05",
		X"38",X"06",X"81",X"06",X"C9",X"06",X"0D",X"07",X"53",X"07",X"94",X"07",X"D2",X"07",X"0F",X"08",
		X"49",X"08",X"84",X"08",X"BA",X"08",X"F0",X"08",X"25",X"09",X"55",X"09",X"86",X"09",X"B6",X"09",
		X"E1",X"09",X"0D",X"0A",X"38",X"0A",X"60",X"0A",X"87",X"0A",X"AD",X"0A",X"D3",X"0A",X"F6",X"0A",
		X"18",X"0B",X"39",X"0B",X"59",X"0B",X"78",X"0B",X"96",X"0B",X"B1",X"0B",X"CD",X"0B",X"E8",X"0B",
		X"01",X"0C",X"17",X"0C",X"2F",X"0C",X"46",X"0C",X"5C",X"0C",X"72",X"0C",X"84",X"0C",X"98",X"0C",
		X"A9",X"0C",X"BB",X"0C",X"B9",X"0C",X"AF",X"0C",X"A9",X"0C",X"A0",X"0C",X"99",X"0C",X"91",X"0C",
		X"89",X"0C",X"83",X"0C",X"7A",X"0C",X"74",X"0C",X"6D",X"0C",X"63",X"0C",X"5E",X"0C",X"55",X"0C",
		X"4E",X"0C",X"45",X"0C",X"40",X"0C",X"37",X"0C",X"2F",X"0C",X"29",X"0C",X"22",X"0C",X"19",X"0C",
		X"11",X"0C",X"0C",X"0C",X"03",X"0C",X"FB",X"0B",X"F5",X"0B",X"EC",X"0B",X"E5",X"0B",X"DF",X"0B",
		X"D7",X"0B",X"D0",X"0B",X"C8",X"0B",X"C1",X"0B",X"B9",X"0B",X"B4",X"0B",X"AB",X"0B",X"A7",X"0B",
		X"9B",X"0B",X"97",X"0B",X"8D",X"0B",X"89",X"0B",X"7F",X"0B",X"7B",X"0B",X"07",X"0B",X"45",X"0A",
		X"90",X"09",X"D2",X"08",X"1D",X"08",X"67",X"07",X"B8",X"06",X"0A",X"06",X"63",X"05",X"BF",X"04",
		X"21",X"04",X"85",X"03",X"EE",X"02",X"5C",X"02",X"CF",X"01",X"46",X"01",X"BF",X"00",X"3D",X"00",
		X"C1",X"FF",X"48",X"FF",X"D2",X"FE",X"5F",X"FE",X"F3",X"FD",X"BB",X"FD",X"C0",X"FD",X"E5",X"FD",
		X"24",X"FE",X"72",X"FE",X"CB",X"FE",X"2A",X"FF",X"8B",X"FF",X"EE",X"FF",X"50",X"00",X"B2",X"00",
		X"12",X"01",X"6E",X"01",X"C9",X"01",X"24",X"02",X"7B",X"02",X"CF",X"02",X"20",X"03",X"71",X"03",
		X"BF",X"03",X"08",X"04",X"51",X"04",X"98",X"04",X"DB",X"04",X"1F",X"05",X"5C",X"05",X"9E",X"05",
		X"C6",X"05",X"B0",X"05",X"6D",X"05",X"0C",X"05",X"99",X"04",X"1B",X"04",X"95",X"03",X"0B",X"03",
		X"82",X"02",X"FA",X"01",X"72",X"01",X"EE",X"00",X"6C",X"00",X"ED",X"FF",X"73",X"FF",X"F9",X"FE",
		X"84",X"FE",X"14",X"FE",X"A6",X"FD",X"3B",X"FD",X"D3",X"FC",X"6F",X"FC",X"0C",X"FC",X"AF",X"FB",
		X"52",X"FB",X"FA",X"FA",X"A2",X"FA",X"5D",X"FA",X"57",X"FA",X"80",X"FA",X"C9",X"FA",X"27",X"FB",
		X"90",X"FB",X"02",X"FC",X"76",X"FC",X"EE",X"FC",X"66",X"FD",X"DD",X"FD",X"50",X"FE",X"C3",X"FE",
		X"32",X"FF",X"A0",X"FF",X"09",X"00",X"6E",X"00",X"D3",X"00",X"34",X"01",X"94",X"01",X"EF",X"01",
		X"48",X"02",X"9E",X"02",X"F1",X"02",X"41",X"03",X"91",X"03",X"DC",X"03",X"27",X"04",X"46",X"04",
		X"2B",X"04",X"E9",X"03",X"8B",X"03",X"1F",X"03",X"A7",X"02",X"2B",X"02",X"AC",X"01",X"2E",X"01",
		X"AE",X"00",X"30",X"00",X"B6",X"FF",X"3F",X"FF",X"C8",X"FE",X"57",X"FE",X"E7",X"FD",X"7B",X"FD",
		X"11",X"FD",X"AB",X"FC",X"4A",X"FC",X"EB",X"FB",X"8D",X"FB",X"32",X"FB",X"DC",X"FA",X"87",X"FA",
		X"35",X"FA",X"E5",X"F9",X"99",X"F9",X"4E",X"F9",X"05",X"F9",X"BF",X"F8",X"7D",X"F8",X"3B",X"F8",
		X"FC",X"F7",X"BF",X"F7",X"82",X"F7",X"4A",X"F7",X"11",X"F7",X"DB",X"F6",X"A8",X"F6",X"76",X"F6",
		X"45",X"F6",X"15",X"F6",X"EA",X"F5",X"BF",X"F5",X"93",X"F5",X"6A",X"F5",X"43",X"F5",X"1C",X"F5",
		X"F8",X"F4",X"D4",X"F4",X"B2",X"F4",X"92",X"F4",X"71",X"F4",X"53",X"F4",X"36",X"F4",X"1A",X"F4",
		X"FD",X"F3",X"E4",X"F3",X"CB",X"F3",X"B2",X"F3",X"9B",X"F3",X"85",X"F3",X"6F",X"F3",X"59",X"F3",
		X"46",X"F3",X"34",X"F3",X"20",X"F3",X"10",X"F3",X"FF",X"F2",X"EF",X"F2",X"DF",X"F2",X"D1",X"F2",
		X"C3",X"F2",X"B6",X"F2",X"A9",X"F2",X"9D",X"F2",X"91",X"F2",X"87",X"F2",X"7D",X"F2",X"73",X"F2",
		X"6A",X"F2",X"64",X"F2",X"97",X"F2",X"FF",X"F2",X"86",X"F3",X"23",X"F4",X"CB",X"F4",X"7B",X"F5",
		X"2D",X"F6",X"E1",X"F6",X"92",X"F7",X"41",X"F8",X"EE",X"F8",X"97",X"F9",X"39",X"FA",X"DA",X"FA",
		X"75",X"FB",X"0E",X"FC",X"9F",X"FC",X"2F",X"FD",X"BA",X"FD",X"41",X"FE",X"C4",X"FE",X"43",X"FF",
		X"BD",X"FF",X"34",X"00",X"A9",X"00",X"19",X"01",X"85",X"01",X"EF",X"01",X"56",X"02",X"B9",X"02",
		X"19",X"03",X"77",X"03",X"D1",X"03",X"2A",X"04",X"7D",X"04",X"D1",X"04",X"1F",X"05",X"6E",X"05",
		X"B9",X"05",X"01",X"06",X"48",X"06",X"8C",X"06",X"CF",X"06",X"0E",X"07",X"4C",X"07",X"88",X"07",
		X"C2",X"07",X"FA",X"07",X"31",X"08",X"65",X"08",X"96",X"08",X"C9",X"08",X"F7",X"08",X"24",X"09",
		X"50",X"09",X"49",X"09",X"07",X"09",X"A6",X"08",X"2A",X"08",X"A2",X"07",X"11",X"07",X"7D",X"06",
		X"E5",X"05",X"50",X"05",X"BA",X"04",X"29",X"04",X"98",X"03",X"0C",X"03",X"83",X"02",X"FF",X"01",
		X"7F",X"01",X"00",X"01",X"86",X"00",X"12",X"00",X"9E",X"FF",X"2E",X"FF",X"C3",X"FE",X"58",X"FE",
		X"F2",X"FD",X"91",X"FD",X"31",X"FD",X"D3",X"FC",X"7A",X"FC",X"24",X"FC",X"CE",X"FB",X"7C",X"FB",
		X"2C",X"FB",X"DF",X"FA",X"96",X"FA",X"4E",X"FA",X"07",X"FA",X"C5",X"F9",X"83",X"F9",X"44",X"F9",
		X"06",X"F9",X"CB",X"F8",X"92",X"F8",X"59",X"F8",X"22",X"F8",X"F0",X"F7",X"BD",X"F7",X"8C",X"F7",
		X"5C",X"F7",X"2F",X"F7",X"03",X"F7",X"D8",X"F6",X"AF",X"F6",X"87",X"F6",X"61",X"F6",X"3C",X"F6",
		X"43",X"F6",X"86",X"F6",X"EB",X"F6",X"69",X"F7",X"F9",X"F7",X"8D",X"F8",X"2A",X"F9",X"C3",X"F9",
		X"63",X"FA",X"FB",X"FA",X"96",X"FB",X"29",X"FC",X"BD",X"FC",X"48",X"FD",X"D6",X"FD",X"57",X"FE",
		X"DF",X"FE",X"5A",X"FF",X"DA",X"FF",X"4D",X"00",X"C5",X"00",X"30",X"01",X"A3",X"01",X"06",X"02",
		X"74",X"02",X"D0",X"02",X"38",X"03",X"8F",X"03",X"F1",X"03",X"42",X"04",X"9F",X"04",X"E9",X"04",
		X"41",X"05",X"86",X"05",X"DB",X"05",X"1A",X"06",X"6B",X"06",X"A5",X"06",X"F0",X"06",X"27",X"07",
		X"71",X"07",X"A0",X"07",X"E7",X"07",X"13",X"08",X"56",X"08",X"7D",X"08",X"BE",X"08",X"E2",X"08",
		X"1E",X"09",X"3E",X"09",X"7B",X"09",X"95",X"09",X"CF",X"09",X"E5",X"09",X"1F",X"0A",X"10",X"0A",
		X"EA",X"09",X"6F",X"09",X"16",X"09",X"58",X"08",X"52",X"08",X"7A",X"0C",X"A3",X"0C",X"8E",X"0C",
		X"8F",X"0C",X"7F",X"0C",X"80",X"0C",X"6F",X"0C",X"71",X"0C",X"60",X"0C",X"61",X"0C",X"51",X"0C",
		X"53",X"0C",X"41",X"0C",X"43",X"0C",X"32",X"0C",X"35",X"0C",X"23",X"0C",X"25",X"0C",X"16",X"0C",
		X"18",X"0C",X"06",X"0C",X"07",X"0C",X"F9",X"0B",X"F8",X"0B",X"E9",X"0B",X"E9",X"0B",X"D9",X"0B",
		X"DB",X"0B",X"CA",X"0B",X"CD",X"0B",X"BD",X"0B",X"BD",X"0B",X"B0",X"0B",X"AE",X"0B",X"A1",X"0B",
		X"A1",X"0B",X"93",X"0B",X"92",X"0B",X"85",X"0B",X"84",X"0B",X"77",X"0B",X"75",X"0B",X"69",X"0B",
		X"67",X"0B",X"5B",X"0B",X"59",X"0B",X"4D",X"0B",X"4B",X"0B",X"41",X"0B",X"3C",X"0B",X"32",X"0B",
		X"2E",X"0B",X"24",X"0B",X"1F",X"0B",X"17",X"0B",X"12",X"0B",X"09",X"0B",X"03",X"0B",X"FB",X"0A",
		X"F4",X"0A",X"EE",X"0A",X"E8",X"0A",X"E0",X"0A",X"DB",X"0A",X"D2",X"0A",X"CE",X"0A",X"C4",X"0A",
		X"BE",X"0A",X"B8",X"0A",X"B1",X"0A",X"AC",X"0A",X"A4",X"0A",X"9D",X"0A",X"96",X"0A",X"8F",X"0A",
		X"8A",X"0A",X"84",X"0A",X"7C",X"0A",X"75",X"0A",X"6E",X"0A",X"69",X"0A",X"62",X"0A",X"5B",X"0A",
		X"55",X"0A",X"4E",X"0A",X"49",X"0A",X"41",X"0A",X"3B",X"0A",X"35",X"0A",X"2E",X"0A",X"27",X"0A",
		X"21",X"0A",X"1B",X"0A",X"14",X"0A",X"0E",X"0A",X"07",X"0A",X"02",X"0A",X"FB",X"09",X"F6",X"09",
		X"EE",X"09",X"E8",X"09",X"E0",X"09",X"DC",X"09",X"D6",X"09",X"CF",X"09",X"C8",X"09",X"C4",X"09",
		X"BB",X"09",X"B7",X"09",X"B0",X"09",X"A9",X"09",X"A4",X"09",X"9C",X"09",X"97",X"09",X"92",X"09",
		X"8B",X"09",X"85",X"09",X"7F",X"09",X"79",X"09",X"72",X"09",X"6D",X"09",X"67",X"09",X"60",X"09",
		X"5C",X"09",X"53",X"09",X"4F",X"09",X"49",X"09",X"44",X"09",X"3D",X"09",X"37",X"09",X"31",X"09",
		X"2B",X"09",X"25",X"09",X"1F",X"09",X"19",X"09",X"15",X"09",X"0E",X"09",X"08",X"09",X"03",X"09",
		X"FE",X"08",X"F6",X"08",X"F1",X"08",X"EB",X"08",X"E6",X"08",X"DF",X"08",X"DA",X"08",X"D5",X"08",
		X"CE",X"08",X"CA",X"08",X"C4",X"08",X"BD",X"08",X"B7",X"08",X"B2",X"08",X"AC",X"08",X"A8",X"08",
		X"A1",X"08",X"9B",X"08",X"97",X"08",X"90",X"08",X"8A",X"08",X"85",X"08",X"7F",X"08",X"7B",X"08",
		X"75",X"08",X"6E",X"08",X"68",X"08",X"64",X"08",X"5E",X"08",X"5A",X"08",X"54",X"08",X"4F",X"08",
		X"49",X"08",X"43",X"08",X"3E",X"08",X"39",X"08",X"32",X"08",X"2D",X"08",X"29",X"08",X"23",X"08",
		X"1D",X"08",X"18",X"08",X"14",X"08",X"0E",X"08",X"08",X"08",X"03",X"08",X"FE",X"07",X"F9",X"07",
		X"F3",X"07",X"EE",X"07",X"EA",X"07",X"E3",X"07",X"DF",X"07",X"D9",X"07",X"D4",X"07",X"CF",X"07",
		X"C9",X"07",X"C5",X"07",X"BF",X"07",X"BB",X"07",X"B5",X"07",X"B0",X"07",X"AC",X"07",X"A5",X"07",
		X"A0",X"07",X"9D",X"07",X"98",X"07",X"92",X"07",X"8C",X"07",X"88",X"07",X"83",X"07",X"7D",X"07",
		X"79",X"07",X"74",X"07",X"6E",X"07",X"69",X"07",X"66",X"07",X"5F",X"07",X"5B",X"07",X"56",X"07",
		X"52",X"07",X"4C",X"07",X"48",X"07",X"42",X"07",X"3D",X"07",X"39",X"07",X"34",X"07",X"2E",X"07",
		X"2B",X"07",X"25",X"07",X"1F",X"07",X"1C",X"07",X"18",X"07",X"11",X"07",X"0D",X"07",X"09",X"07",
		X"04",X"07",X"00",X"07",X"FA",X"06",X"F6",X"06",X"F1",X"06",X"EB",X"06",X"E8",X"06",X"E4",X"06",
		X"DD",X"06",X"D9",X"06",X"D6",X"06",X"CF",X"06",X"CB",X"06",X"C7",X"06",X"C2",X"06",X"BE",X"06",
		X"B8",X"06",X"B5",X"06",X"AF",X"06",X"AB",X"06",X"A7",X"06",X"A2",X"06",X"9E",X"06",X"98",X"06",
		X"94",X"06",X"90",X"06",X"8C",X"06",X"88",X"06",X"83",X"06",X"7E",X"06",X"79",X"06",X"74",X"06",
		X"70",X"06",X"6B",X"06",X"67",X"06",X"63",X"06",X"5E",X"06",X"5B",X"06",X"56",X"06",X"52",X"06",
		X"4C",X"06",X"4A",X"06",X"45",X"06",X"41",X"06",X"3C",X"06",X"37",X"06",X"33",X"06",X"2F",X"06",
		X"2B",X"06",X"25",X"06",X"22",X"06",X"1D",X"06",X"18",X"06",X"15",X"06",X"10",X"06",X"0C",X"06",
		X"09",X"06",X"04",X"06",X"01",X"06",X"FD",X"05",X"F7",X"05",X"F2",X"05",X"EF",X"05",X"EB",X"05",
		X"E7",X"05",X"E4",X"05",X"DE",X"05",X"DA",X"05",X"D7",X"05",X"D2",X"05",X"CF",X"05",X"CA",X"05",
		X"C5",X"05",X"C2",X"05",X"BC",X"05",X"BA",X"05",X"B6",X"05",X"B2",X"05",X"AD",X"05",X"AA",X"05",
		X"A5",X"05",X"A0",X"05",X"9D",X"05",X"9A",X"05",X"95",X"05",X"91",X"05",X"8B",X"05",X"8A",X"05",
		X"86",X"05",X"81",X"05",X"7D",X"05",X"78",X"05",X"75",X"05",X"71",X"05",X"6D",X"05",X"69",X"05",
		X"65",X"05",X"61",X"05",X"5E",X"05",X"59",X"05",X"55",X"05",X"53",X"05",X"4E",X"05",X"4B",X"05",
		X"48",X"05",X"42",X"05",X"3F",X"05",X"3B",X"05",X"38",X"05",X"33",X"05",X"31",X"05",X"2D",X"05",
		X"28",X"05",X"25",X"05",X"21",X"05",X"1C",X"05",X"19",X"05",X"17",X"05",X"12",X"05",X"10",X"05",
		X"0B",X"05",X"08",X"05",X"04",X"05",X"00",X"05",X"FC",X"04",X"F9",X"04",X"F5",X"04",X"F2",X"04",
		X"ED",X"04",X"E9",X"04",X"E6",X"04",X"E3",X"04",X"E0",X"04",X"DC",X"04",X"D8",X"04",X"D5",X"04",
		X"D0",X"04",X"CD",X"04",X"C8",X"04",X"C6",X"04",X"C2",X"04",X"BF",X"04",X"BB",X"04",X"B8",X"04",
		X"B4",X"04",X"B1",X"04",X"AD",X"04",X"AA",X"04",X"A6",X"04",X"A4",X"04",X"9F",X"04",X"9C",X"04",
		X"98",X"04",X"95",X"04",X"93",X"04",X"8E",X"04",X"8B",X"04",X"88",X"04",X"85",X"04",X"81",X"04",
		X"7D",X"04",X"7A",X"04",X"77",X"04",X"74",X"04",X"6F",X"04",X"6C",X"04",X"69",X"04",X"66",X"04",
		X"63",X"04",X"5E",X"04",X"5B",X"04",X"58",X"04",X"55",X"04",X"51",X"04",X"50",X"04",X"4B",X"04",
		X"48",X"04",X"44",X"04",X"42",X"04",X"3E",X"04",X"3B",X"04",X"37",X"04",X"33",X"04",X"30",X"04",
		X"2C",X"04",X"2A",X"04",X"27",X"04",X"24",X"04",X"21",X"04",X"1D",X"04",X"1A",X"04",X"17",X"04",
		X"13",X"04",X"12",X"04",X"0D",X"04",X"0B",X"04",X"08",X"04",X"04",X"04",X"01",X"04",X"FD",X"03",
		X"FB",X"03",X"F8",X"03",X"F4",X"03",X"F0",X"03",X"EE",X"03",X"EA",X"03",X"E8",X"03",X"E5",X"03",
		X"E2",X"03",X"DF",X"03",X"DB",X"03",X"D8",X"03",X"D6",X"03",X"D2",X"03",X"CF",X"03",X"CD",X"03",
		X"C9",X"03",X"C6",X"03",X"C3",X"03",X"C0",X"03",X"BD",X"03",X"BA",X"03",X"B8",X"03",X"B4",X"03",
		X"B2",X"03",X"AE",X"03",X"AC",X"03",X"AA",X"03",X"A8",X"03",X"A3",X"03",X"A1",X"03",X"9D",X"03",
		X"9B",X"03",X"98",X"03",X"95",X"03",X"91",X"03",X"8E",X"03",X"8C",X"03",X"89",X"03",X"86",X"03",
		X"82",X"03",X"80",X"03",X"7C",X"03",X"7A",X"03",X"78",X"03",X"75",X"03",X"72",X"03",X"70",X"03",
		X"6C",X"03",X"68",X"03",X"67",X"03",X"64",X"03",X"61",X"03",X"5D",X"03",X"5B",X"03",X"58",X"03",
		X"55",X"03",X"53",X"03",X"4F",X"03",X"4E",X"03",X"4A",X"03",X"48",X"03",X"46",X"03",X"42",X"03",
		X"40",X"03",X"3D",X"03",X"3B",X"03",X"38",X"03",X"35",X"03",X"32",X"03",X"2E",X"03",X"2C",X"03",
		X"2A",X"03",X"27",X"03",X"25",X"03",X"22",X"03",X"1E",X"03",X"1D",X"03",X"1B",X"03",X"17",X"03",
		X"15",X"03",X"12",X"03",X"10",X"03",X"0D",X"03",X"0C",X"03",X"08",X"03",X"05",X"03",X"02",X"03",
		X"00",X"03",X"FD",X"02",X"FB",X"02",X"F8",X"02",X"F6",X"02",X"F2",X"02",X"F1",X"02",X"ED",X"02",
		X"EC",X"02",X"E9",X"02",X"E7",X"02",X"E4",X"02",X"E2",X"02",X"DE",X"02",X"DD",X"02",X"DB",X"02",
		X"D7",X"02",X"D5",X"02",X"D2",X"02",X"D0",X"02",X"CF",X"02",X"CB",X"02",X"C8",X"02",X"C5",X"02",
		X"C3",X"02",X"C1",X"02",X"BF",X"02",X"BD",X"02",X"BB",X"02",X"B8",X"02",X"B5",X"02",X"B2",X"02",
		X"AF",X"02",X"AE",X"02",X"AA",X"02",X"A7",X"02",X"A6",X"02",X"A4",X"02",X"A3",X"02",X"9F",X"02",
		X"9E",X"02",X"9B",X"02",X"98",X"02",X"96",X"02",X"93",X"02",X"91",X"02",X"8F",X"02",X"8D",X"02",
		X"8A",X"02",X"87",X"02",X"86",X"02",X"83",X"02",X"80",X"02",X"7F",X"02",X"7C",X"02",X"7A",X"02",
		X"77",X"02",X"75",X"02",X"71",X"02",X"72",X"02",X"6E",X"02",X"6A",X"02",X"6C",X"02",X"66",X"02",
		X"65",X"02",X"64",X"02",X"61",X"02",X"5E",X"02",X"5D",X"02",X"5B",X"02",X"58",X"02",X"56",X"02",
		X"54",X"02",X"51",X"02",X"4E",X"02",X"4D",X"02",X"4B",X"02",X"49",X"02",X"46",X"02",X"44",X"02",
		X"42",X"02",X"40",X"02",X"3D",X"02",X"3B",X"02",X"39",X"02",X"37",X"02",X"35",X"02",X"32",X"02",
		X"2F",X"02",X"2E",X"02",X"2D",X"02",X"2B",X"02",X"29",X"02",X"27",X"02",X"24",X"02",X"22",X"02",
		X"20",X"02",X"1E",X"02",X"1B",X"02",X"1A",X"02",X"17",X"02",X"15",X"02",X"12",X"02",X"12",X"02",
		X"10",X"02",X"0C",X"02",X"0B",X"02",X"08",X"02",X"06",X"02",X"05",X"02",X"02",X"02",X"00",X"02",
		X"FF",X"01",X"FE",X"01",X"FC",X"01",X"F8",X"01",X"F7",X"01",X"F4",X"01",X"F4",X"01",X"F0",X"01",
		X"EE",X"01",X"EC",X"01",X"EB",X"01",X"E9",X"01",X"E7",X"01",X"E5",X"01",X"E3",X"01",X"E0",X"01",
		X"E0",X"01",X"DD",X"01",X"DA",X"01",X"D9",X"01",X"D7",X"01",X"D5",X"01",X"D3",X"01",X"D1",X"01",
		X"CE",X"01",X"CC",X"01",X"CC",X"01",X"C9",X"01",X"C8",X"01",X"C5",X"01",X"C4",X"01",X"C3",X"01",
		X"C0",X"01",X"BF",X"01",X"BD",X"01",X"BB",X"01",X"B9",X"01",X"B6",X"01",X"B5",X"01",X"B3",X"01",
		X"B1",X"01",X"AF",X"01",X"AD",X"01",X"AB",X"01",X"AA",X"01",X"A7",X"01",X"A7",X"01",X"A3",X"01",
		X"A1",X"01",X"9F",X"01",X"9E",X"01",X"9E",X"01",X"9B",X"01",X"99",X"01",X"98",X"01",X"96",X"01",
		X"95",X"01",X"91",X"01",X"90",X"01",X"8F",X"01",X"8C",X"01",X"89",X"01",X"87",X"01",X"88",X"01",
		X"86",X"01",X"83",X"01",X"84",X"01",X"7F",X"01",X"80",X"01",X"7E",X"01",X"7B",X"01",X"79",X"01",
		X"77",X"01",X"76",X"01",X"74",X"01",X"71",X"01",X"70",X"01",X"6F",X"01",X"6D",X"01",X"6A",X"01",
		X"6A",X"01",X"68",X"01",X"68",X"01",X"65",X"01",X"62",X"01",X"61",X"01",X"60",X"01",X"5E",X"01",
		X"5C",X"01",X"5B",X"01",X"59",X"01",X"58",X"01",X"55",X"01",X"53",X"01",X"52",X"01",X"50",X"01",
		X"4E",X"01",X"4E",X"01",X"4C",X"01",X"4C",X"01",X"48",X"01",X"47",X"01",X"44",X"01",X"43",X"01",
		X"42",X"01",X"3E",X"01",X"40",X"01",X"3D",X"01",X"3B",X"01",X"39",X"01",X"39",X"01",X"37",X"01",
		X"37",X"01",X"33",X"01",X"32",X"01",X"31",X"01",X"2F",X"01",X"2E",X"01",X"2A",X"01",X"29",X"01",
		X"29",X"01",X"27",X"01",X"25",X"01",X"24",X"01",X"22",X"01",X"22",X"01",X"1F",X"01",X"1D",X"01",
		X"1D",X"01",X"1B",X"01",X"1A",X"01",X"18",X"01",X"16",X"01",X"15",X"01",X"13",X"01",X"11",X"01",
		X"10",X"01",X"0F",X"01",X"0E",X"01",X"0D",X"01",X"0B",X"01",X"09",X"01",X"08",X"01",X"06",X"01",
		X"06",X"01",X"03",X"01",X"01",X"01",X"00",X"01",X"FF",X"00",X"FD",X"00",X"FB",X"00",X"FB",X"00",
		X"F9",X"00",X"F7",X"00",X"F6",X"00",X"F4",X"00",X"F2",X"00",X"F2",X"00",X"F1",X"00",X"EF",X"00",
		X"ED",X"00",X"EC",X"00",X"EB",X"00",X"E9",X"00",X"E8",X"00",X"E7",X"00",X"E6",X"00",X"E3",X"00",
		X"E2",X"00",X"E2",X"00",X"E0",X"00",X"DD",X"00",X"DD",X"00",X"DB",X"00",X"D9",X"00",X"D9",X"00",
		X"D6",X"00",X"D6",X"00",X"D4",X"00",X"D3",X"00",X"D1",X"00",X"D1",X"00",X"D0",X"00",X"CC",X"00",
		X"CD",X"00",X"CB",X"00",X"C9",X"00",X"C7",X"00",X"C7",X"00",X"C6",X"00",X"C4",X"00",X"C3",X"00",
		X"C2",X"00",X"C0",X"00",X"BE",X"00",X"BE",X"00",X"BE",X"00",X"BB",X"00",X"B9",X"00",X"B8",X"00",
		X"B7",X"00",X"B5",X"00",X"B4",X"00",X"B2",X"00",X"B2",X"00",X"B0",X"00",X"AF",X"00",X"AE",X"00",
		X"AC",X"00",X"AC",X"00",X"AA",X"00",X"A8",X"00",X"A7",X"00",X"A7",X"00",X"A5",X"00",X"A3",X"00",
		X"A4",X"00",X"A2",X"00",X"9F",X"00",X"A0",X"00",X"9E",X"00",X"9D",X"00",X"9C",X"00",X"9A",X"00",
		X"99",X"00",X"97",X"00",X"96",X"00",X"95",X"00",X"93",X"00",X"93",X"00",X"91",X"00",X"8F",X"00",
		X"8E",X"00",X"8D",X"00",X"8E",X"00",X"8C",X"00",X"8A",X"00",X"88",X"00",X"87",X"00",X"86",X"00",
		X"84",X"00",X"85",X"00",X"83",X"00",X"82",X"00",X"81",X"00",X"80",X"00",X"7F",X"00",X"7E",X"00",
		X"7C",X"00",X"7B",X"00",X"79",X"00",X"79",X"00",X"76",X"00",X"76",X"00",X"76",X"00",X"73",X"00",
		X"73",X"00",X"71",X"00",X"71",X"00",X"70",X"00",X"6E",X"00",X"6E",X"00",X"6C",X"00",X"6B",X"00",
		X"69",X"00",X"69",X"00",X"67",X"00",X"66",X"00",X"65",X"00",X"64",X"00",X"63",X"00",X"62",X"00",
		X"60",X"00",X"60",X"00",X"5E",X"00",X"5D",X"00",X"5C",X"00",X"5B",X"00",X"5A",X"00",X"59",X"00",
		X"59",X"00",X"57",X"00",X"55",X"00",X"56",X"00",X"54",X"00",X"53",X"00",X"53",X"00",X"50",X"00",
		X"50",X"00",X"4F",X"00",X"4E",X"00",X"4C",X"00",X"4C",X"00",X"4B",X"00",X"49",X"00",X"48",X"00",
		X"48",X"00",X"45",X"00",X"46",X"00",X"45",X"00",X"44",X"00",X"43",X"00",X"41",X"00",X"40",X"00",
		X"3E",X"00",X"3E",X"00",X"3C",X"00",X"3C",X"00",X"3B",X"00",X"3A",X"00",X"39",X"00",X"38",X"00",
		X"37",X"00",X"37",X"00",X"35",X"00",X"34",X"00",X"32",X"00",X"32",X"00",X"30",X"00",X"30",X"00",
		X"2E",X"00",X"2D",X"00",X"2D",X"00",X"2C",X"00",X"2A",X"00",X"2A",X"00",X"2A",X"00",X"27",X"00",
		X"28",X"00",X"26",X"00",X"25",X"00",X"26",X"00",X"22",X"00",X"22",X"00",X"21",X"00",X"21",X"00",
		X"20",X"00",X"1E",X"00",X"1E",X"00",X"1C",X"00",X"1C",X"00",X"1A",X"00",X"1A",X"00",X"19",X"00",
		X"18",X"00",X"17",X"00",X"17",X"00",X"15",X"00",X"13",X"00",X"14",X"00",X"13",X"00",X"13",X"00",
		X"10",X"00",X"0F",X"00",X"0F",X"00",X"0E",X"00",X"0D",X"00",X"0C",X"00",X"0B",X"00",X"0B",X"00",
		X"09",X"00",X"09",X"00",X"08",X"00",X"06",X"00",X"06",X"00",X"06",X"00",X"04",X"00",X"04",X"00",
		X"03",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FE",X"FF",
		X"FD",X"FF",X"FB",X"FF",X"FA",X"FF",X"FA",X"FF",X"F9",X"FF",X"F8",X"FF",X"F7",X"FF",X"F7",X"FF",
		X"F7",X"FF",X"F5",X"FF",X"F3",X"FF",X"F4",X"FF",X"F3",X"FF",X"F2",X"FF",X"F2",X"FF",X"F0",X"FF",
		X"F1",X"FF",X"EF",X"FF",X"ED",X"FF",X"EC",X"FF",X"EC",X"FF",X"EB",X"FF",X"EB",X"FF",X"E9",X"FF",
		X"E8",X"FF",X"E9",X"FF",X"E7",X"FF",X"E6",X"FF",X"E5",X"FF",X"E4",X"FF",X"E4",X"FF",X"E2",X"FF",
		X"E3",X"FF",X"E2",X"FF",X"E0",X"FF",X"E0",X"FF",X"DF",X"FF",X"DE",X"FF",X"DE",X"FF",X"DC",X"FF",
		X"DD",X"FF",X"DB",X"FF",X"DA",X"FF",X"D9",X"FF",X"DB",X"FF",X"DA",X"FF",X"DA",X"FF",X"D7",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
