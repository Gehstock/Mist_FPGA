library IEEE;
use IEEE.std_logic_1164.all;

package mc_pack is
    constant HW_GALAXIAN : integer := 0;
    constant HW_MOONCR   : integer := 1;
    constant HW_AZURIAN  : integer := 2;
    constant HW_BLKHOLE  : integer := 3;
    constant HW_CATACOMB : integer := 4;
    constant HW_CHEWINGG : integer := 5;
    constant HW_DEVILFSH : integer := 6;
    constant HW_KINGBAL  : integer := 7;
    constant HW_MRDONIGH : integer := 8;
    constant HW_OMEGA    : integer := 9;
    constant HW_ORBITRON : integer := 10;
    constant HW_PISCES   : integer := 11;
    constant HW_UNIWARS  : integer := 12;
    constant HW_VICTORY  : integer := 13;
    constant HW_WAROFBUG : integer := 14;
    constant HW_ZIGZAG   : integer := 15; -- doesn't work yet
    constant HW_TRIPLEDR : integer := 16;
end;