library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_PGM_0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_PGM_0 is
	type rom is array(0 to  12287) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
    x"00",x"AF",x"32",x"01",x"70",x"C3",x"C8",x"00", -- 0x0000
    x"41",x"5A",x"55",x"52",x"49",x"41",x"4E",x"20", -- 0x0008
    x"41",x"54",x"54",x"41",x"43",x"4B",x"20",x"43", -- 0x0010
    x"4F",x"50",x"59",x"52",x"49",x"47",x"48",x"54", -- 0x0018
    x"20",x"52",x"41",x"49",x"54",x"20",x"45",x"4C", -- 0x0020
    x"45",x"43",x"54",x"52",x"4F",x"4E",x"49",x"43", -- 0x0028
    x"53",x"20",x"4C",x"54",x"44",x"20",x"31",x"39", -- 0x0030
    x"38",x"32",x"20",x"41",x"4C",x"4C",x"20",x"52", -- 0x0038
    x"49",x"47",x"48",x"54",x"53",x"20",x"52",x"45", -- 0x0040
    x"53",x"45",x"52",x"56",x"45",x"44",x"00",x"00", -- 0x0048
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0050
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0058
    x"00",x"00",x"00",x"00",x"00",x"00",x"F5",x"C5", -- 0x0060
    x"D5",x"E5",x"DD",x"E5",x"FD",x"E5",x"3A",x"00", -- 0x0068
    x"78",x"AF",x"32",x"01",x"70",x"21",x"B6",x"40", -- 0x0070
    x"35",x"21",x"C0",x"41",x"11",x"00",x"58",x"01", -- 0x0078
    x"80",x"00",x"ED",x"B0",x"3A",x"AF",x"40",x"CB", -- 0x0080
    x"67",x"28",x"14",x"11",x"04",x"00",x"06",x"04", -- 0x0088
    x"21",x"63",x"58",x"3E",x"F3",x"96",x"77",x"19", -- 0x0090
    x"3E",x"5E",x"96",x"77",x"19",x"10",x"F4",x"CD", -- 0x0098
    x"F4",x"0F",x"3A",x"BF",x"40",x"A7",x"C4",x"CD", -- 0x00A0
    x"04",x"DD",x"21",x"AF",x"40",x"DD",x"CB",x"00", -- 0x00A8
    x"4E",x"C2",x"C3",x"18",x"CD",x"66",x"22",x"3E", -- 0x00B0
    x"FF",x"32",x"01",x"70",x"FD",x"E1",x"DD",x"E1", -- 0x00B8
    x"E1",x"D1",x"C1",x"F1",x"ED",x"45",x"00",x"00", -- 0x00C0
    x"31",x"00",x"44",x"CD",x"F4",x"12",x"AF",x"21", -- 0x00C8
    x"00",x"60",x"06",x"04",x"77",x"23",x"10",x"FC", -- 0x00D0
    x"3C",x"06",x"04",x"77",x"23",x"10",x"FC",x"AF", -- 0x00D8
    x"06",x"08",x"21",x"00",x"68",x"77",x"23",x"10", -- 0x00E0
    x"FC",x"06",x"08",x"21",x"01",x"70",x"77",x"23", -- 0x00E8
    x"10",x"FC",x"3D",x"32",x"00",x"78",x"21",x"16", -- 0x00F0
    x"11",x"11",x"00",x"40",x"01",x"00",x"01",x"ED", -- 0x00F8
    x"B0",x"06",x"01",x"3A",x"00",x"70",x"CB",x"47", -- 0x0100
    x"28",x"01",x"04",x"78",x"32",x"B2",x"40",x"32", -- 0x0108
    x"B1",x"40",x"CD",x"42",x"13",x"C3",x"BE",x"01", -- 0x0110
    x"31",x"00",x"44",x"DD",x"CB",x"00",x"DE",x"DD", -- 0x0118
    x"CB",x"00",x"96",x"DD",x"CB",x"00",x"8E",x"AF", -- 0x0120
    x"32",x"BF",x"40",x"32",x"EE",x"40",x"32",x"EF", -- 0x0128
    x"40",x"CD",x"42",x"13",x"CD",x"F4",x"12",x"CD", -- 0x0130
    x"B6",x"12",x"DD",x"36",x"1F",x"05",x"DD",x"36", -- 0x0138
    x"1E",x"04",x"21",x"A7",x"01",x"FD",x"21",x"0F", -- 0x0140
    x"53",x"06",x"11",x"CD",x"3F",x"12",x"DD",x"21", -- 0x0148
    x"AF",x"40",x"3A",x"00",x"68",x"CB",x"47",x"20", -- 0x0150
    x"06",x"CB",x"4F",x"20",x"2A",x"18",x"EF",x"DD", -- 0x0158
    x"CB",x"00",x"FE",x"DD",x"CB",x"00",x"B6",x"21", -- 0x0160
    x"D9",x"40",x"CB",x"DE",x"21",x"B8",x"01",x"FD", -- 0x0168
    x"21",x"01",x"51",x"06",x"06",x"CD",x"3F",x"12", -- 0x0170
    x"3A",x"B0",x"40",x"D6",x"01",x"27",x"32",x"B0", -- 0x0178
    x"40",x"CD",x"9E",x"12",x"C3",x"A9",x"05",x"3A", -- 0x0180
    x"B0",x"40",x"FE",x"02",x"38",x"C0",x"21",x"D9", -- 0x0188
    x"40",x"CB",x"DE",x"DD",x"CB",x"00",x"BE",x"DD", -- 0x0190
    x"CB",x"00",x"F6",x"D6",x"02",x"27",x"32",x"B0", -- 0x0198
    x"40",x"CD",x"9E",x"12",x"C3",x"A9",x"05",x"50", -- 0x01A0
    x"55",x"53",x"48",x"40",x"53",x"54",x"41",x"52", -- 0x01A8
    x"54",x"40",x"42",x"55",x"54",x"54",x"4F",x"4E", -- 0x01B0
    x"40",x"40",x"40",x"40",x"40",x"40",x"DD",x"21", -- 0x01B8
    x"C0",x"41",x"CD",x"F4",x"12",x"3E",x"64",x"CD", -- 0x01C0
    x"38",x"13",x"DD",x"36",x"07",x"01",x"DD",x"36", -- 0x01C8
    x"06",x"04",x"FD",x"21",x"23",x"53",x"3E",x"02", -- 0x01D0
    x"CD",x"38",x"13",x"11",x"E0",x"FF",x"21",x"7D", -- 0x01D8
    x"04",x"06",x"14",x"CD",x"64",x"04",x"3E",x"14", -- 0x01E0
    x"CD",x"38",x"13",x"DD",x"36",x"0F",x"02",x"FD", -- 0x01E8
    x"21",x"67",x"52",x"21",x"91",x"04",x"06",x"08", -- 0x01F0
    x"CD",x"64",x"04",x"3E",x"50",x"CD",x"38",x"13", -- 0x01F8
    x"DD",x"36",x"20",x"FC",x"DD",x"36",x"22",x"FC", -- 0x0200
    x"DD",x"36",x"1C",x"00",x"DD",x"36",x"3E",x"00", -- 0x0208
    x"DD",x"36",x"3F",x"01",x"21",x"B0",x"52",x"11", -- 0x0210
    x"99",x"04",x"06",x"0D",x"1A",x"77",x"13",x"23", -- 0x0218
    x"1A",x"77",x"13",x"23",x"23",x"23",x"1A",x"77", -- 0x0220
    x"13",x"23",x"1A",x"77",x"13",x"D5",x"11",x"DB", -- 0x0228
    x"FF",x"19",x"D1",x"10",x"E7",x"3E",x"24",x"32", -- 0x0230
    x"0E",x"51",x"3E",x"1D",x"32",x"EE",x"50",x"21", -- 0x0238
    x"D5",x"03",x"11",x"E0",x"FF",x"FD",x"21",x"BF", -- 0x0240
    x"52",x"06",x"0E",x"CD",x"73",x"04",x"21",x"DD", -- 0x0248
    x"41",x"22",x"C0",x"40",x"21",x"08",x"03",x"22", -- 0x0250
    x"C2",x"40",x"21",x"BF",x"40",x"CB",x"C6",x"CB", -- 0x0258
    x"CE",x"3E",x"FF",x"CD",x"38",x"13",x"CB",x"86", -- 0x0260
    x"CB",x"8E",x"CD",x"F4",x"12",x"3E",x"32",x"CD", -- 0x0268
    x"38",x"13",x"DD",x"36",x"00",x"FC",x"DD",x"36", -- 0x0270
    x"02",x"FC",x"DD",x"36",x"3E",x"00",x"DD",x"36", -- 0x0278
    x"3F",x"01",x"21",x"A0",x"52",x"11",x"99",x"04", -- 0x0280
    x"06",x"0D",x"1A",x"77",x"13",x"23",x"1A",x"77", -- 0x0288
    x"13",x"13",x"13",x"D5",x"11",x"DF",x"FF",x"19", -- 0x0290
    x"D1",x"10",x"EF",x"21",x"C1",x"41",x"22",x"C0", -- 0x0298
    x"40",x"21",x"03",x"02",x"22",x"C2",x"40",x"21", -- 0x02A0
    x"BF",x"40",x"CB",x"C6",x"DD",x"36",x"09",x"03", -- 0x02A8
    x"21",x"B3",x"03",x"FD",x"21",x"C4",x"52",x"06", -- 0x02B0
    x"0E",x"CD",x"3F",x"12",x"21",x"D5",x"03",x"11", -- 0x02B8
    x"E0",x"FF",x"FD",x"21",x"BF",x"52",x"06",x"0E", -- 0x02C0
    x"CD",x"73",x"04",x"3E",x"32",x"CD",x"38",x"13", -- 0x02C8
    x"11",x"00",x"42",x"21",x"C1",x"03",x"01",x"14", -- 0x02D0
    x"00",x"ED",x"B0",x"21",x"CE",x"41",x"06",x"10", -- 0x02D8
    x"36",x"60",x"23",x"36",x"04",x"23",x"10",x"F8", -- 0x02E0
    x"06",x"06",x"36",x"00",x"23",x"36",x"04",x"23", -- 0x02E8
    x"10",x"F8",x"DD",x"21",x"BF",x"40",x"DD",x"CB", -- 0x02F0
    x"00",x"DE",x"21",x"E3",x"03",x"06",x"05",x"C5", -- 0x02F8
    x"11",x"C4",x"40",x"01",x"0A",x"00",x"ED",x"B0", -- 0x0300
    x"FD",x"2A",x"CC",x"40",x"EB",x"2A",x"CA",x"40", -- 0x0308
    x"EB",x"DD",x"CB",x"00",x"D6",x"1A",x"BE",x"20", -- 0x0310
    x"FC",x"23",x"FD",x"36",x"00",x"01",x"DD",x"CB", -- 0x0318
    x"00",x"56",x"20",x"FA",x"C1",x"10",x"D8",x"3E", -- 0x0320
    x"32",x"CD",x"38",x"13",x"FD",x"21",x"B8",x"52", -- 0x0328
    x"DD",x"21",x"B8",x"51",x"21",x"4C",x"04",x"11", -- 0x0330
    x"E0",x"FF",x"06",x"02",x"FD",x"E5",x"DD",x"E5", -- 0x0338
    x"C5",x"7E",x"FD",x"77",x"00",x"23",x"FD",x"19", -- 0x0340
    x"7E",x"FD",x"77",x"00",x"23",x"3E",x"32",x"CD", -- 0x0348
    x"38",x"13",x"06",x"0A",x"7E",x"DD",x"77",x"00", -- 0x0350
    x"23",x"DD",x"19",x"10",x"F7",x"3E",x"32",x"CD", -- 0x0358
    x"38",x"13",x"C1",x"DD",x"E1",x"FD",x"E1",x"DD", -- 0x0360
    x"23",x"DD",x"23",x"DD",x"23",x"FD",x"23",x"FD", -- 0x0368
    x"23",x"FD",x"23",x"10",x"C7",x"3E",x"FF",x"CD", -- 0x0370
    x"38",x"13",x"AF",x"32",x"BF",x"40",x"CD",x"F4", -- 0x0378
    x"12",x"3E",x"32",x"CD",x"38",x"13",x"CD",x"B6", -- 0x0380
    x"12",x"CD",x"AA",x"12",x"3A",x"BC",x"40",x"3C", -- 0x0388
    x"FE",x"05",x"20",x"02",x"3E",x"01",x"32",x"BC", -- 0x0390
    x"40",x"32",x"1E",x"40",x"21",x"AF",x"40",x"CB", -- 0x0398
    x"D6",x"E5",x"CD",x"93",x"06",x"E1",x"CB",x"8E", -- 0x03A0
    x"3E",x"40",x"CD",x"38",x"13",x"CD",x"AA",x"12", -- 0x03A8
    x"C3",x"BE",x"01",x"46",x"41",x"54",x"41",x"4C", -- 0x03B0
    x"49",x"54",x"59",x"40",x"53",x"43",x"4F",x"52", -- 0x03B8
    x"45",x"00",x"14",x"03",x"3F",x"00",x"18",x"00", -- 0x03C0
    x"5C",x"00",x"13",x"06",x"6F",x"00",x"15",x"06", -- 0x03C8
    x"8B",x"00",x"32",x"04",x"A2",x"13",x"1F",x"20", -- 0x03D0
    x"29",x"22",x"19",x"17",x"18",x"24",x"10",x"01", -- 0x03D8
    x"09",x"08",x"02",x"1A",x"04",x"A9",x"51",x"0A", -- 0x03E0
    x"01",x"D2",x"41",x"00",x"42",x"50",x"24",x"04", -- 0x03E8
    x"AC",x"51",x"0A",x"01",x"D8",x"41",x"04",x"42", -- 0x03F0
    x"4C",x"2E",x"04",x"AF",x"51",x"0A",x"01",x"DE", -- 0x03F8
    x"41",x"08",x"42",x"50",x"38",x"04",x"B2",x"51", -- 0x0400
    x"0A",x"01",x"E4",x"41",x"0C",x"42",x"4C",x"42", -- 0x0408
    x"04",x"B5",x"51",x"0A",x"01",x"EA",x"41",x"10", -- 0x0410
    x"42",x"4C",x"10",x"05",x"03",x"10",x"20",x"1F", -- 0x0418
    x"19",x"1E",x"24",x"23",x"01",x"00",x"00",x"10", -- 0x0420
    x"20",x"1F",x"19",x"1E",x"24",x"23",x"02",x"00", -- 0x0428
    x"00",x"10",x"20",x"1F",x"19",x"1E",x"24",x"23", -- 0x0430
    x"01",x"05",x"00",x"10",x"20",x"1F",x"19",x"1E", -- 0x0438
    x"24",x"23",x"10",x"03",x"00",x"10",x"20",x"1F", -- 0x0440
    x"19",x"1E",x"24",x"23",x"0C",x"10",x"01",x"00", -- 0x0448
    x"00",x"10",x"20",x"1F",x"19",x"1E",x"24",x"23", -- 0x0450
    x"0D",x"10",x"10",x"05",x"00",x"10",x"20",x"1F", -- 0x0458
    x"19",x"1E",x"24",x"23",x"7E",x"FD",x"77",x"00", -- 0x0460
    x"23",x"FD",x"19",x"3E",x"0A",x"CD",x"38",x"13", -- 0x0468
    x"10",x"F2",x"C9",x"7E",x"FD",x"77",x"00",x"23", -- 0x0470
    x"FD",x"19",x"10",x"F7",x"C9",x"22",x"11",x"19", -- 0x0478
    x"24",x"10",x"15",x"1C",x"15",x"13",x"24",x"22", -- 0x0480
    x"1F",x"1E",x"19",x"13",x"23",x"10",x"1C",x"24", -- 0x0488
    x"14",x"20",x"22",x"15",x"23",x"15",x"1E",x"24", -- 0x0490
    x"23",x"68",x"6B",x"68",x"6B",x"69",x"6A",x"69", -- 0x0498
    x"6A",x"6C",x"6F",x"BB",x"B5",x"6D",x"6E",x"BA", -- 0x04A0
    x"B4",x"AC",x"AF",x"BB",x"B5",x"AD",x"AE",x"BA", -- 0x04A8
    x"B4",x"B0",x"B3",x"68",x"6B",x"B1",x"B2",x"69", -- 0x04B0
    x"6A",x"0A",x"0A",x"BD",x"BF",x"68",x"6B",x"BC", -- 0x04B8
    x"BE",x"69",x"6A",x"C1",x"C3",x"B7",x"B9",x"C0", -- 0x04C0
    x"C2",x"B6",x"B8",x"10",x"10",x"0F",x"DC",x"13", -- 0x04C8
    x"05",x"0F",x"DC",x"E0",x"04",x"0F",x"F5",x"DC", -- 0x04D0
    x"2F",x"05",x"F1",x"0F",x"DC",x"63",x"05",x"C9", -- 0x04D8
    x"DD",x"21",x"37",x"40",x"FD",x"21",x"04",x"42", -- 0x04E0
    x"DD",x"CB",x"00",x"56",x"F5",x"C4",x"D6",x"1C", -- 0x04E8
    x"F1",x"C0",x"F5",x"CD",x"67",x"0B",x"E6",x"0F", -- 0x04F0
    x"6F",x"26",x"00",x"29",x"11",x"89",x"05",x"19", -- 0x04F8
    x"7E",x"FD",x"77",x"00",x"23",x"7E",x"FD",x"77", -- 0x0500
    x"03",x"FD",x"36",x"01",x"13",x"DD",x"36",x"00", -- 0x0508
    x"07",x"F1",x"C9",x"21",x"C3",x"40",x"35",x"C0", -- 0x0510
    x"F5",x"36",x"03",x"2B",x"46",x"2A",x"C0",x"40", -- 0x0518
    x"7E",x"3C",x"FE",x"08",x"20",x"02",x"3E",x"01", -- 0x0520
    x"77",x"23",x"23",x"10",x"FB",x"F1",x"C9",x"2A", -- 0x0528
    x"CC",x"40",x"7E",x"A7",x"28",x"01",x"34",x"2A", -- 0x0530
    x"CA",x"40",x"35",x"20",x"05",x"21",x"BF",x"40", -- 0x0538
    x"CB",x"96",x"21",x"C9",x"40",x"35",x"C0",x"36", -- 0x0540
    x"08",x"2B",x"7E",x"A7",x"C8",x"35",x"2A",x"C6", -- 0x0548
    x"40",x"EB",x"2A",x"C4",x"40",x"7E",x"12",x"23", -- 0x0550
    x"22",x"C4",x"40",x"21",x"E0",x"FF",x"19",x"22", -- 0x0558
    x"C6",x"40",x"C9",x"3A",x"92",x"51",x"FE",x"10", -- 0x0560
    x"C8",x"21",x"45",x"40",x"FD",x"21",x"0C",x"42", -- 0x0568
    x"34",x"7E",x"E6",x"18",x"20",x"0A",x"FD",x"36", -- 0x0570
    x"02",x"07",x"3E",x"05",x"32",x"92",x"51",x"C9", -- 0x0578
    x"FD",x"36",x"02",x"06",x"AF",x"32",x"92",x"51", -- 0x0580
    x"C9",x"28",x"94",x"B8",x"94",x"AB",x"76",x"A0", -- 0x0588
    x"A6",x"40",x"A8",x"40",x"78",x"63",x"63",x"85", -- 0x0590
    x"6B",x"73",x"7C",x"59",x"8C",x"79",x"93",x"79", -- 0x0598
    x"99",x"89",x"A4",x"95",x"9C",x"60",x"A0",x"54", -- 0x05A0
    x"A8",x"DD",x"CB",x"00",x"EE",x"CD",x"17",x"13", -- 0x05A8
    x"CD",x"AA",x"12",x"06",x"03",x"3A",x"00",x"68", -- 0x05B0
    x"4F",x"CB",x"7F",x"28",x"02",x"06",x"05",x"78", -- 0x05B8
    x"32",x"1D",x"40",x"06",x"04",x"CB",x"71",x"28", -- 0x05C0
    x"02",x"06",x"02",x"3A",x"00",x"70",x"0F",x"0F", -- 0x05C8
    x"E6",x"01",x"EE",x"01",x"80",x"32",x"F4",x"40", -- 0x05D0
    x"21",x"1D",x"40",x"11",x"00",x"41",x"01",x"1A", -- 0x05D8
    x"00",x"ED",x"B0",x"21",x"A9",x"40",x"06",x"03", -- 0x05E0
    x"AF",x"77",x"23",x"10",x"FC",x"CD",x"4E",x"12", -- 0x05E8
    x"3A",x"AF",x"40",x"CB",x"7F",x"20",x"0D",x"21", -- 0x05F0
    x"AC",x"40",x"06",x"03",x"AF",x"77",x"23",x"10", -- 0x05F8
    x"FC",x"CD",x"57",x"12",x"21",x"BE",x"40",x"06", -- 0x0600
    x"50",x"3A",x"00",x"70",x"CB",x"4F",x"28",x"02", -- 0x0608
    x"06",x"70",x"78",x"F6",x"03",x"77",x"21",x"AF", -- 0x0610
    x"40",x"4E",x"06",x"00",x"CB",x"A6",x"CB",x"69", -- 0x0618
    x"20",x"0B",x"3A",x"00",x"70",x"CB",x"5F",x"28", -- 0x0620
    x"04",x"06",x"01",x"CB",x"E6",x"78",x"32",x"06", -- 0x0628
    x"70",x"32",x"07",x"70",x"11",x"E0",x"FF",x"21", -- 0x0630
    x"9F",x"53",x"06",x"06",x"3E",x"10",x"77",x"19", -- 0x0638
    x"10",x"FC",x"3A",x"1D",x"40",x"32",x"BF",x"53", -- 0x0640
    x"A7",x"28",x"0A",x"47",x"21",x"9F",x"53",x"3E", -- 0x0648
    x"0F",x"77",x"19",x"10",x"FC",x"DD",x"21",x"C0", -- 0x0650
    x"41",x"DD",x"36",x"13",x"02",x"DD",x"36",x"12", -- 0x0658
    x"04",x"DD",x"36",x"17",x"06",x"CD",x"2E",x"08", -- 0x0660
    x"06",x"06",x"C5",x"21",x"02",x"08",x"FD",x"21", -- 0x0668
    x"49",x"52",x"06",x"05",x"CD",x"3F",x"12",x"3E", -- 0x0670
    x"10",x"CD",x"38",x"13",x"21",x"F2",x"07",x"FD", -- 0x0678
    x"21",x"49",x"52",x"06",x"05",x"CD",x"3F",x"12", -- 0x0680
    x"3E",x"0A",x"CD",x"38",x"13",x"C1",x"10",x"DA", -- 0x0688
    x"CD",x"17",x"13",x"21",x"16",x"11",x"11",x"00", -- 0x0690
    x"40",x"01",x"15",x"00",x"ED",x"B0",x"21",x"4D", -- 0x0698
    x"11",x"11",x"37",x"40",x"01",x"70",x"00",x"ED", -- 0x06A0
    x"B0",x"21",x"95",x"0E",x"3A",x"1E",x"40",x"E6", -- 0x06A8
    x"03",x"20",x"03",x"21",x"40",x"10",x"CD",x"07", -- 0x06B0
    x"14",x"CD",x"C4",x"13",x"21",x"AF",x"40",x"CB", -- 0x06B8
    x"CE",x"CD",x"B9",x"07",x"3A",x"01",x"40",x"CB", -- 0x06C0
    x"47",x"C2",x"D2",x"06",x"CD",x"83",x"09",x"C3", -- 0x06C8
    x"C1",x"06",x"DD",x"21",x"37",x"40",x"06",x"07", -- 0x06D0
    x"11",x"10",x"00",x"DD",x"CB",x"00",x"FE",x"DD", -- 0x06D8
    x"19",x"10",x"F8",x"CD",x"B9",x"07",x"3A",x"16", -- 0x06E0
    x"40",x"A7",x"20",x"F7",x"3A",x"01",x"40",x"CB", -- 0x06E8
    x"57",x"28",x"F0",x"21",x"AF",x"40",x"CB",x"56", -- 0x06F0
    x"C0",x"CB",x"8E",x"3E",x"40",x"CD",x"38",x"13", -- 0x06F8
    x"21",x"00",x"68",x"AF",x"06",x"03",x"77",x"23", -- 0x0700
    x"10",x"FC",x"CD",x"17",x"13",x"3A",x"AF",x"40", -- 0x0708
    x"CB",x"77",x"C2",x"45",x"07",x"3A",x"1D",x"40", -- 0x0710
    x"A7",x"C2",x"95",x"07",x"CD",x"46",x"08",x"CD", -- 0x0718
    x"14",x"21",x"3A",x"1D",x"40",x"A7",x"C2",x"95", -- 0x0720
    x"07",x"21",x"06",x"70",x"AF",x"77",x"23",x"77", -- 0x0728
    x"21",x"AF",x"40",x"CB",x"A6",x"CD",x"07",x"08", -- 0x0730
    x"3E",x"64",x"CD",x"38",x"13",x"21",x"AF",x"40", -- 0x0738
    x"CB",x"9E",x"C3",x"BE",x"01",x"3A",x"1D",x"40", -- 0x0740
    x"A7",x"20",x"28",x"CD",x"07",x"08",x"DD",x"36", -- 0x0748
    x"17",x"06",x"3A",x"AF",x"40",x"4F",x"CD",x"2E", -- 0x0750
    x"08",x"3E",x"30",x"CD",x"38",x"13",x"CD",x"46", -- 0x0758
    x"08",x"CD",x"14",x"21",x"3A",x"00",x"41",x"A7", -- 0x0760
    x"20",x"10",x"3A",x"1D",x"40",x"A7",x"20",x"03", -- 0x0768
    x"C3",x"29",x"07",x"3A",x"00",x"41",x"A7",x"CA", -- 0x0770
    x"95",x"07",x"21",x"1D",x"40",x"11",x"00",x"41", -- 0x0778
    x"06",x"1A",x"1A",x"4F",x"7E",x"12",x"71",x"13", -- 0x0780
    x"23",x"10",x"F7",x"21",x"AF",x"40",x"3E",x"20", -- 0x0788
    x"AE",x"77",x"C3",x"95",x"07",x"3A",x"1E",x"40", -- 0x0790
    x"E6",x"03",x"CA",x"16",x"06",x"FD",x"21",x"37", -- 0x0798
    x"40",x"3D",x"20",x"06",x"FD",x"34",x"F7",x"C3", -- 0x07A0
    x"16",x"06",x"3D",x"20",x"06",x"FD",x"34",x"FC", -- 0x07A8
    x"C3",x"16",x"06",x"FD",x"34",x"FA",x"C3",x"16", -- 0x07B0
    x"06",x"3A",x"1E",x"40",x"E6",x"03",x"28",x"1F", -- 0x07B8
    x"CD",x"18",x"0B",x"CD",x"C4",x"08",x"CD",x"F6", -- 0x07C0
    x"25",x"CD",x"96",x"28",x"CD",x"11",x"1F",x"CD", -- 0x07C8
    x"7D",x"20",x"CD",x"08",x"14",x"CD",x"00",x"0C", -- 0x07D0
    x"CD",x"73",x"08",x"CD",x"F2",x"24",x"C9",x"CD", -- 0x07D8
    x"73",x"08",x"CD",x"08",x"14",x"CD",x"30",x"17", -- 0x07E0
    x"CD",x"7F",x"19",x"CD",x"54",x"0E",x"CD",x"4B", -- 0x07E8
    x"25",x"C9",x"40",x"40",x"40",x"40",x"40",x"40", -- 0x07F0
    x"40",x"40",x"40",x"40",x"50",x"4C",x"41",x"59", -- 0x07F8
    x"45",x"52",x"52",x"45",x"41",x"44",x"59",x"DD", -- 0x0800
    x"21",x"C0",x"41",x"DD",x"36",x"13",x"02",x"DD", -- 0x0808
    x"36",x"12",x"04",x"3E",x"01",x"CD",x"38",x"13", -- 0x0810
    x"21",x"25",x"08",x"FD",x"21",x"89",x"52",x"06", -- 0x0818
    x"09",x"CD",x"3F",x"12",x"C9",x"47",x"41",x"4D", -- 0x0820
    x"45",x"40",x"4F",x"56",x"45",x"52",x"21",x"FC", -- 0x0828
    x"07",x"FD",x"21",x"6B",x"52",x"06",x"06",x"CD", -- 0x0830
    x"3F",x"12",x"3E",x"01",x"CB",x"69",x"20",x"02", -- 0x0838
    x"3E",x"02",x"32",x"8B",x"51",x"C9",x"11",x"A9", -- 0x0840
    x"40",x"3A",x"AF",x"40",x"4F",x"CB",x"6F",x"20", -- 0x0848
    x"03",x"11",x"AC",x"40",x"D5",x"21",x"B3",x"40", -- 0x0850
    x"E5",x"06",x"03",x"1A",x"BE",x"38",x"11",x"20", -- 0x0858
    x"04",x"23",x"13",x"10",x"F6",x"D1",x"E1",x"01", -- 0x0860
    x"03",x"00",x"ED",x"B0",x"CD",x"60",x"12",x"C9", -- 0x0868
    x"E1",x"E1",x"C9",x"06",x"01",x"11",x"A9",x"40", -- 0x0870
    x"3A",x"AF",x"40",x"CB",x"6F",x"20",x"05",x"11", -- 0x0878
    x"AC",x"40",x"CB",x"20",x"21",x"BE",x"40",x"78", -- 0x0880
    x"A6",x"C8",x"1A",x"A7",x"20",x"08",x"13",x"7E", -- 0x0888
    x"E6",x"F0",x"4F",x"1A",x"B9",x"D8",x"78",x"AE", -- 0x0890
    x"77",x"21",x"1D",x"40",x"34",x"11",x"E0",x"FF", -- 0x0898
    x"21",x"9F",x"53",x"06",x"06",x"3E",x"10",x"77", -- 0x08A0
    x"19",x"10",x"FC",x"3A",x"1D",x"40",x"32",x"BF", -- 0x08A8
    x"53",x"A7",x"28",x"0A",x"47",x"21",x"9F",x"53", -- 0x08B0
    x"3E",x"0F",x"77",x"19",x"10",x"FC",x"21",x"D9", -- 0x08B8
    x"40",x"CB",x"E6",x"C9",x"3A",x"01",x"40",x"CB", -- 0x08C0
    x"47",x"C0",x"DD",x"21",x"37",x"40",x"FD",x"21", -- 0x08C8
    x"04",x"42",x"3A",x"1E",x"40",x"E6",x"03",x"FE", -- 0x08D0
    x"01",x"CA",x"74",x"25",x"FE",x"02",x"CA",x"4B", -- 0x08D8
    x"27",x"FE",x"03",x"CA",x"58",x"1F",x"C9",x"1E", -- 0x08E0
    x"00",x"3A",x"00",x"42",x"FD",x"96",x"00",x"30", -- 0x08E8
    x"04",x"ED",x"44",x"CB",x"C3",x"47",x"3A",x"03", -- 0x08F0
    x"42",x"FD",x"96",x"03",x"30",x"04",x"ED",x"44", -- 0x08F8
    x"CB",x"CB",x"4F",x"B8",x"38",x"04",x"CB",x"FB", -- 0x0900
    x"48",x"47",x"CB",x"21",x"CB",x"21",x"78",x"B9", -- 0x0908
    x"30",x"0B",x"CB",x"20",x"80",x"30",x"0C",x"0E", -- 0x0910
    x"01",x"06",x"01",x"18",x"0A",x"0E",x"00",x"06", -- 0x0918
    x"02",x"18",x"04",x"0E",x"01",x"06",x"02",x"CB", -- 0x0920
    x"7B",x"28",x"03",x"78",x"41",x"4F",x"CB",x"43", -- 0x0928
    x"28",x"04",x"78",x"ED",x"44",x"47",x"CB",x"4B", -- 0x0930
    x"28",x"04",x"79",x"ED",x"44",x"4F",x"C9",x"DD", -- 0x0938
    x"21",x"37",x"40",x"FD",x"21",x"04",x"42",x"DD", -- 0x0940
    x"7E",x"DF",x"FE",x"07",x"C8",x"06",x"07",x"DD", -- 0x0948
    x"CB",x"00",x"56",x"CA",x"07",x"14",x"CD",x"78", -- 0x0950
    x"09",x"10",x"F4",x"C9",x"DD",x"21",x"37",x"40", -- 0x0958
    x"FD",x"21",x"04",x"42",x"06",x"07",x"FD",x"BE", -- 0x0960
    x"01",x"F5",x"C5",x"E5",x"CC",x"07",x"14",x"E1", -- 0x0968
    x"C1",x"F1",x"CD",x"78",x"09",x"10",x"EF",x"C9", -- 0x0970
    x"11",x"10",x"00",x"DD",x"19",x"11",x"04",x"00", -- 0x0978
    x"FD",x"19",x"C9",x"3A",x"1E",x"40",x"E6",x"03", -- 0x0980
    x"FE",x"01",x"CA",x"98",x"09",x"FE",x"02",x"CA", -- 0x0988
    x"B3",x"09",x"FE",x"03",x"CA",x"CE",x"09",x"C9", -- 0x0990
    x"21",x"2E",x"40",x"7E",x"A7",x"C0",x"3A",x"18", -- 0x0998
    x"40",x"FE",x"01",x"D0",x"21",x"CF",x"40",x"35", -- 0x09A0
    x"C0",x"23",x"35",x"C0",x"36",x"02",x"21",x"1E", -- 0x09A8
    x"40",x"34",x"C9",x"21",x"33",x"40",x"7E",x"A7", -- 0x09B0
    x"C0",x"21",x"16",x"40",x"7E",x"A7",x"C0",x"21", -- 0x09B8
    x"CF",x"40",x"35",x"C0",x"23",x"35",x"C0",x"36", -- 0x09C0
    x"02",x"21",x"1E",x"40",x"34",x"C9",x"21",x"31", -- 0x09C8
    x"40",x"7E",x"A7",x"C0",x"3A",x"19",x"40",x"A7", -- 0x09D0
    x"C0",x"01",x"00",x"01",x"C5",x"CD",x"B9",x"07", -- 0x09D8
    x"3A",x"16",x"40",x"A7",x"20",x"F7",x"C1",x"0B", -- 0x09E0
    x"78",x"B1",x"20",x"F0",x"21",x"AF",x"40",x"CB", -- 0x09E8
    x"8E",x"21",x"00",x"42",x"11",x"01",x"42",x"01", -- 0x09F0
    x"40",x"00",x"36",x"00",x"ED",x"B0",x"3E",x"50", -- 0x09F8
    x"CD",x"38",x"13",x"CD",x"17",x"13",x"3E",x"08", -- 0x0A00
    x"CD",x"38",x"13",x"3A",x"1E",x"40",x"3C",x"32", -- 0x0A08
    x"1E",x"40",x"CD",x"40",x"10",x"3E",x"20",x"CD", -- 0x0A10
    x"38",x"13",x"11",x"00",x"42",x"21",x"29",x"0A", -- 0x0A18
    x"01",x"04",x"00",x"ED",x"B0",x"E1",x"C3",x"BC", -- 0x0A20
    x"06",x"E0",x"11",x"01",x"E0",x"21",x"AF",x"40", -- 0x0A28
    x"CB",x"8E",x"21",x"00",x"68",x"AF",x"77",x"23", -- 0x0A30
    x"77",x"23",x"77",x"31",x"00",x"44",x"21",x"28", -- 0x0A38
    x"40",x"FD",x"21",x"05",x"53",x"AF",x"ED",x"67", -- 0x0A40
    x"FD",x"77",x"00",x"ED",x"67",x"FD",x"77",x"20", -- 0x0A48
    x"ED",x"67",x"2B",x"AF",x"ED",x"67",x"FD",x"77", -- 0x0A50
    x"40",x"ED",x"67",x"FD",x"77",x"60",x"ED",x"67", -- 0x0A58
    x"3E",x"60",x"CD",x"38",x"13",x"21",x"D1",x"41", -- 0x0A60
    x"22",x"C0",x"40",x"21",x"12",x"03",x"22",x"C2", -- 0x0A68
    x"40",x"3E",x"01",x"32",x"BF",x"40",x"06",x"11", -- 0x0A70
    x"FD",x"21",x"05",x"53",x"21",x"EF",x"40",x"E5", -- 0x0A78
    x"CB",x"FE",x"3E",x"01",x"CD",x"38",x"13",x"21", -- 0x0A80
    x"28",x"40",x"7E",x"90",x"27",x"77",x"F5",x"AF", -- 0x0A88
    x"ED",x"67",x"FD",x"77",x"00",x"ED",x"67",x"FD", -- 0x0A90
    x"77",x"20",x"ED",x"67",x"2B",x"F1",x"7E",x"DE", -- 0x0A98
    x"00",x"27",x"77",x"AF",x"ED",x"67",x"FD",x"77", -- 0x0AA0
    x"40",x"ED",x"67",x"FD",x"77",x"60",x"ED",x"67", -- 0x0AA8
    x"16",x"00",x"58",x"E5",x"C5",x"FD",x"E5",x"CD", -- 0x0AB0
    x"72",x"19",x"FD",x"E1",x"C1",x"E1",x"7E",x"A7", -- 0x0AB8
    x"20",x"C0",x"06",x"01",x"23",x"7E",x"A7",x"20", -- 0x0AC0
    x"B9",x"E1",x"CB",x"BE",x"3E",x"60",x"CD",x"38", -- 0x0AC8
    x"13",x"21",x"D1",x"41",x"3E",x"04",x"BE",x"20", -- 0x0AD0
    x"FD",x"AF",x"32",x"BF",x"40",x"21",x"14",x"0B", -- 0x0AD8
    x"FD",x"21",x"65",x"53",x"06",x"04",x"CD",x"3F", -- 0x0AE0
    x"12",x"3E",x"78",x"CD",x"38",x"13",x"CD",x"17", -- 0x0AE8
    x"13",x"21",x"1E",x"40",x"34",x"7E",x"E6",x"C0", -- 0x0AF0
    x"28",x"03",x"3E",x"3D",x"77",x"CD",x"7F",x"26", -- 0x0AF8
    x"21",x"00",x"42",x"36",x"80",x"23",x"36",x"10", -- 0x0B00
    x"23",x"36",x"01",x"23",x"36",x"80",x"CD",x"95", -- 0x0B08
    x"0E",x"C3",x"BC",x"06",x"48",x"4F",x"4D",x"45", -- 0x0B10
    x"DD",x"21",x"37",x"40",x"FD",x"21",x"04",x"42", -- 0x0B18
    x"21",x"16",x"40",x"06",x"07",x"AF",x"77",x"23", -- 0x0B20
    x"10",x"FC",x"06",x"07",x"DD",x"CB",x"00",x"56", -- 0x0B28
    x"28",x"17",x"DD",x"CB",x"00",x"46",x"20",x"11", -- 0x0B30
    x"FD",x"7E",x"01",x"D6",x"13",x"FE",x"07",x"30", -- 0x0B38
    x"08",x"21",x"16",x"40",x"34",x"85",x"6F",x"23", -- 0x0B40
    x"34",x"CD",x"78",x"09",x"10",x"DE",x"C9",x"DD", -- 0x0B48
    x"CB",x"00",x"46",x"C0",x"AF",x"FD",x"77",x"00", -- 0x0B50
    x"FD",x"77",x"01",x"FD",x"77",x"03",x"DD",x"CB", -- 0x0B58
    x"00",x"8E",x"DD",x"CB",x"00",x"96",x"C9",x"E5", -- 0x0B60
    x"21",x"A7",x"40",x"7E",x"0F",x"AE",x"07",x"23", -- 0x0B68
    x"34",x"86",x"EA",x"76",x"0B",x"34",x"2B",x"77", -- 0x0B70
    x"E1",x"C9",x"05",x"20",x"05",x"20",x"05",x"20", -- 0x0B78
    x"05",x"20",x"05",x"20",x"05",x"21",x"05",x"22", -- 0x0B80
    x"05",x"12",x"05",x"02",x"05",x"12",x"05",x"11", -- 0x0B88
    x"05",x"FE",x"05",x"20",x"05",x"2F",x"05",x"1F", -- 0x0B90
    x"05",x"1E",x"05",x"0E",x"05",x"1E",x"05",x"1F", -- 0x0B98
    x"05",x"2F",x"05",x"20",x"05",x"21",x"05",x"11", -- 0x0BA0
    x"05",x"12",x"05",x"02",x"05",x"F2",x"05",x"F1", -- 0x0BA8
    x"05",x"E1",x"05",x"E0",x"05",x"E1",x"05",x"F1", -- 0x0BB0
    x"05",x"F1",x"05",x"F1",x"05",x"F1",x"05",x"F1", -- 0x0BB8
    x"05",x"E1",x"05",x"E0",x"05",x"E1",x"05",x"F1", -- 0x0BC0
    x"05",x"F2",x"05",x"02",x"05",x"12",x"05",x"11", -- 0x0BC8
    x"05",x"21",x"05",x"20",x"05",x"2F",x"05",x"1F", -- 0x0BD0
    x"05",x"1E",x"05",x"0E",x"05",x"FE",x"05",x"FF", -- 0x0BD8
    x"05",x"EF",x"05",x"E0",x"05",x"E0",x"05",x"FF", -- 0x0BE0
    x"05",x"FF",x"05",x"FF",x"05",x"FF",x"05",x"FF", -- 0x0BE8
    x"05",x"FF",x"05",x"FF",x"05",x"FE",x"05",x"0E", -- 0x0BF0
    x"05",x"1E",x"05",x"1F",x"05",x"1E",x"05",x"20", -- 0x0BF8
    x"3A",x"01",x"40",x"CB",x"47",x"C0",x"FD",x"21", -- 0x0C00
    x"00",x"42",x"FD",x"66",x"00",x"FD",x"6E",x"03", -- 0x0C08
    x"DD",x"21",x"37",x"40",x"FD",x"21",x"04",x"42", -- 0x0C10
    x"06",x"07",x"DD",x"CB",x"00",x"56",x"E5",x"C5", -- 0x0C18
    x"C4",x"2B",x"0C",x"C1",x"E1",x"CD",x"78",x"09", -- 0x0C20
    x"10",x"F0",x"C9",x"DD",x"CB",x"00",x"46",x"C0", -- 0x0C28
    x"7C",x"FD",x"96",x"00",x"57",x"30",x"02",x"ED", -- 0x0C30
    x"44",x"FE",x"10",x"D0",x"47",x"3E",x"10",x"90", -- 0x0C38
    x"47",x"7D",x"FD",x"96",x"03",x"4F",x"30",x"02", -- 0x0C40
    x"ED",x"44",x"FE",x"10",x"D0",x"7A",x"F5",x"21", -- 0x0C48
    x"AC",x"14",x"FD",x"7E",x"01",x"D6",x"13",x"FE", -- 0x0C50
    x"06",x"D2",x"C8",x"0C",x"0F",x"0F",x"0F",x"5F", -- 0x0C58
    x"16",x"00",x"19",x"E5",x"21",x"D9",x"0C",x"3A", -- 0x0C60
    x"01",x"42",x"BE",x"28",x"05",x"23",x"23",x"23", -- 0x0C68
    x"18",x"F8",x"23",x"5E",x"23",x"56",x"E1",x"F1", -- 0x0C70
    x"A7",x"FA",x"AF",x"0C",x"CB",x"27",x"85",x"6F", -- 0x0C78
    x"3E",x"00",x"8C",x"67",x"EB",x"1A",x"81",x"C6", -- 0x0C80
    x"20",x"23",x"BE",x"DA",x"BC",x"0C",x"2B",x"13", -- 0x0C88
    x"1A",x"81",x"C6",x"20",x"BE",x"28",x"03",x"D2", -- 0x0C90
    x"C2",x"0C",x"3A",x"1E",x"40",x"E6",x"03",x"CA", -- 0x0C98
    x"79",x"0E",x"CD",x"EB",x"18",x"DD",x"CB",x"00", -- 0x0CA0
    x"C6",x"21",x"01",x"40",x"CB",x"C6",x"C9",x"ED", -- 0x0CA8
    x"44",x"CB",x"27",x"83",x"5F",x"3E",x"00",x"8A", -- 0x0CB0
    x"57",x"C3",x"84",x"0C",x"13",x"13",x"23",x"10", -- 0x0CB8
    x"C4",x"C9",x"23",x"23",x"13",x"10",x"BE",x"C9", -- 0x0CC0
    x"21",x"F1",x"0D",x"FD",x"7E",x"01",x"11",x"20", -- 0x0CC8
    x"00",x"BE",x"23",x"CA",x"63",x"0C",x"19",x"18", -- 0x0CD0
    x"F8",x"10",x"F1",x"0C",x"50",x"11",x"0D",x"11", -- 0x0CD8
    x"31",x"0D",x"91",x"51",x"0D",x"12",x"71",x"0D", -- 0x0CE0
    x"52",x"91",x"0D",x"92",x"B1",x"0D",x"D2",x"D1", -- 0x0CE8
    x"0D",x"25",x"21",x"24",x"21",x"24",x"21",x"29", -- 0x0CF0
    x"23",x"2A",x"23",x"2B",x"23",x"2C",x"23",x"2B", -- 0x0CF8
    x"23",x"2A",x"23",x"29",x"23",x"24",x"21",x"24", -- 0x0D00
    x"21",x"25",x"21",x"50",x"50",x"50",x"50",x"50", -- 0x0D08
    x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"2E", -- 0x0D10
    x"2A",x"2E",x"2B",x"2E",x"2B",x"2C",x"26",x"2C", -- 0x0D18
    x"25",x"2C",x"24",x"2C",x"23",x"2C",x"24",x"2C", -- 0x0D20
    x"25",x"2C",x"26",x"2E",x"2B",x"2E",x"2B",x"2E", -- 0x0D28
    x"2A",x"2C",x"22",x"2C",x"22",x"2C",x"22",x"2C", -- 0x0D30
    x"22",x"2C",x"22",x"2C",x"22",x"29",x"25",x"29", -- 0x0D38
    x"25",x"28",x"26",x"28",x"26",x"28",x"26",x"28", -- 0x0D40
    x"26",x"2A",x"24",x"29",x"25",x"28",x"26",x"27", -- 0x0D48
    x"27",x"28",x"28",x"29",x"27",x"2A",x"26",x"2B", -- 0x0D50
    x"25",x"29",x"27",x"29",x"27",x"29",x"27",x"29", -- 0x0D58
    x"27",x"2A",x"26",x"2A",x"26",x"2D",x"23",x"2D", -- 0x0D60
    x"23",x"2D",x"23",x"2D",x"23",x"2D",x"23",x"2D", -- 0x0D68
    x"23",x"2B",x"2B",x"2B",x"2A",x"2B",x"29",x"2D", -- 0x0D70
    x"2A",x"2B",x"2A",x"2B",x"29",x"2B",x"29",x"2B", -- 0x0D78
    x"26",x"2C",x"25",x"2F",x"24",x"2F",x"24",x"2F", -- 0x0D80
    x"25",x"2F",x"26",x"2F",x"2C",x"2F",x"2C",x"2F", -- 0x0D88
    x"2B",x"24",x"24",x"25",x"22",x"26",x"22",x"25", -- 0x0D90
    x"22",x"25",x"24",x"26",x"24",x"26",x"24",x"29", -- 0x0D98
    x"24",x"2A",x"23",x"2B",x"20",x"2B",x"20",x"2A", -- 0x0DA0
    x"20",x"29",x"20",x"23",x"20",x"23",x"20",x"24", -- 0x0DA8
    x"20",x"2F",x"2B",x"2F",x"2C",x"2F",x"2C",x"2F", -- 0x0DB0
    x"26",x"2F",x"25",x"2F",x"24",x"2F",x"24",x"2C", -- 0x0DB8
    x"25",x"2B",x"26",x"2B",x"29",x"2B",x"29",x"2B", -- 0x0DC0
    x"2A",x"2D",x"2A",x"2B",x"29",x"2B",x"2A",x"2B", -- 0x0DC8
    x"2B",x"24",x"20",x"23",x"20",x"23",x"20",x"29", -- 0x0DD0
    x"20",x"2A",x"20",x"2B",x"20",x"2B",x"20",x"2A", -- 0x0DD8
    x"23",x"29",x"24",x"26",x"24",x"26",x"24",x"25", -- 0x0DE0
    x"24",x"25",x"22",x"26",x"22",x"25",x"22",x"24", -- 0x0DE8
    x"24",x"33",x"0F",x"08",x"0F",x"08",x"0F",x"08", -- 0x0DF0
    x"0F",x"08",x"0F",x"08",x"0F",x"08",x"0F",x"08", -- 0x0DF8
    x"0F",x"08",x"0F",x"08",x"0F",x"06",x"0F",x"04", -- 0x0E00
    x"0F",x"02",x"0F",x"00",x"0F",x"00",x"0F",x"00", -- 0x0E08
    x"0F",x"00",x"B3",x"0F",x"00",x"0F",x"00",x"0F", -- 0x0E10
    x"00",x"0F",x"00",x"0F",x"02",x"0F",x"04",x"0F", -- 0x0E18
    x"06",x"0F",x"08",x"0F",x"08",x"0F",x"08",x"0F", -- 0x0E20
    x"08",x"0F",x"08",x"0F",x"08",x"0F",x"08",x"0F", -- 0x0E28
    x"08",x"0F",x"08",x"97",x"0F",x"06",x"0F",x"05", -- 0x0E30
    x"0F",x"04",x"0F",x"03",x"0F",x"02",x"0F",x"01", -- 0x0E38
    x"0F",x"00",x"0F",x"00",x"0F",x"00",x"0F",x"00", -- 0x0E40
    x"0F",x"00",x"0F",x"00",x"0F",x"00",x"0F",x"00", -- 0x0E48
    x"0F",x"00",x"0F",x"00",x"3A",x"01",x"40",x"CB", -- 0x0E50
    x"47",x"C0",x"FD",x"21",x"00",x"42",x"FD",x"66", -- 0x0E58
    x"00",x"FD",x"6E",x"03",x"FD",x"21",x"04",x"42", -- 0x0E60
    x"06",x"04",x"E5",x"C5",x"CD",x"30",x"0C",x"C1", -- 0x0E68
    x"E1",x"11",x"04",x"00",x"FD",x"19",x"10",x"F2", -- 0x0E70
    x"C9",x"E1",x"E1",x"E1",x"FD",x"7E",x"01",x"FE", -- 0x0E78
    x"33",x"28",x"0A",x"FE",x"B3",x"28",x"06",x"21", -- 0x0E80
    x"01",x"40",x"CB",x"C6",x"C9",x"1A",x"FE",x"08", -- 0x0E88
    x"20",x"F5",x"C3",x"2D",x"0A",x"0E",x"02",x"21", -- 0x0E90
    x"C4",x"41",x"11",x"F0",x"0F",x"1A",x"47",x"13", -- 0x0E98
    x"1A",x"13",x"36",x"00",x"23",x"77",x"23",x"10", -- 0x0EA0
    x"F9",x"0D",x"20",x"F1",x"21",x"11",x"0F",x"46", -- 0x0EA8
    x"23",x"C5",x"5E",x"23",x"56",x"23",x"46",x"23", -- 0x0EB0
    x"4E",x"23",x"D5",x"C5",x"06",x"00",x"ED",x"B0", -- 0x0EB8
    x"C1",x"D1",x"E5",x"21",x"20",x"00",x"19",x"EB", -- 0x0EC0
    x"E1",x"10",x"EF",x"C1",x"10",x"E3",x"3E",x"2C", -- 0x0EC8
    x"06",x"26",x"21",x"A0",x"0F",x"5E",x"23",x"56", -- 0x0ED0
    x"23",x"12",x"10",x"F9",x"C9",x"3A",x"B6",x"40", -- 0x0ED8
    x"A7",x"C0",x"3E",x"0A",x"32",x"B6",x"40",x"3A", -- 0x0EE0
    x"09",x"40",x"CB",x"27",x"21",x"A0",x"0F",x"5F", -- 0x0EE8
    x"16",x"00",x"19",x"5E",x"23",x"56",x"3E",x"2C", -- 0x0EF0
    x"12",x"CD",x"67",x"0B",x"E6",x"1F",x"32",x"09", -- 0x0EF8
    x"40",x"CB",x"27",x"21",x"A0",x"0F",x"5F",x"16", -- 0x0F00
    x"00",x"19",x"5E",x"23",x"56",x"3E",x"10",x"12", -- 0x0F08
    x"C9",x"03",x"42",x"50",x"0C",x"06",x"2D",x"2D", -- 0x0F10
    x"2D",x"92",x"AA",x"10",x"2D",x"2D",x"2D",x"93", -- 0x0F18
    x"A9",x"0B",x"2D",x"2D",x"2D",x"94",x"A8",x"AB", -- 0x0F20
    x"2D",x"2D",x"92",x"95",x"10",x"10",x"2D",x"2D", -- 0x0F28
    x"96",x"A7",x"10",x"10",x"2D",x"98",x"97",x"10", -- 0x0F30
    x"10",x"10",x"2D",x"99",x"A1",x"10",x"10",x"10", -- 0x0F38
    x"98",x"A0",x"A2",x"A6",x"10",x"10",x"9A",x"9F", -- 0x0F40
    x"10",x"A5",x"10",x"10",x"9B",x"9E",x"A3",x"A4", -- 0x0F48
    x"10",x"10",x"9C",x"10",x"10",x"10",x"10",x"10", -- 0x0F50
    x"9D",x"10",x"10",x"10",x"10",x"10",x"59",x"50", -- 0x0F58
    x"08",x"06",x"35",x"2E",x"3D",x"2D",x"2D",x"2D", -- 0x0F60
    x"34",x"2E",x"3C",x"81",x"85",x"88",x"33",x"39", -- 0x0F68
    x"3B",x"2E",x"84",x"87",x"32",x"2D",x"2D",x"80", -- 0x0F70
    x"83",x"2D",x"31",x"2D",x"2D",x"2D",x"2D",x"2D", -- 0x0F78
    x"30",x"38",x"2D",x"2D",x"2D",x"2D",x"2F",x"37", -- 0x0F80
    x"2D",x"3F",x"2D",x"2D",x"10",x"36",x"3A",x"3E", -- 0x0F88
    x"82",x"86",x"90",x"53",x"02",x"05",x"8A",x"8C", -- 0x0F90
    x"8E",x"90",x"10",x"89",x"8B",x"8D",x"8F",x"91", -- 0x0F98
    x"72",x"50",x"D1",x"50",x"EF",x"50",x"0E",x"51", -- 0x0FA0
    x"10",x"51",x"4E",x"51",x"94",x"51",x"F8",x"51", -- 0x0FA8
    x"19",x"52",x"83",x"53",x"5A",x"52",x"78",x"52", -- 0x0FB0
    x"9A",x"52",x"9E",x"52",x"B3",x"52",x"B9",x"52", -- 0x0FB8
    x"BB",x"52",x"DA",x"52",x"DD",x"52",x"FB",x"52", -- 0x0FC0
    x"43",x"53",x"18",x"53",x"1A",x"53",x"1C",x"53", -- 0x0FC8
    x"3D",x"53",x"3E",x"53",x"54",x"53",x"5C",x"53", -- 0x0FD0
    x"77",x"53",x"7D",x"53",x"9A",x"53",x"B8",x"53", -- 0x0FD8
    x"BB",x"53",x"BE",x"53",x"A2",x"53",x"44",x"53", -- 0x0FE0
    x"A7",x"53",x"28",x"53",x"00",x"50",x"00",x"50", -- 0x0FE8
    x"06",x"06",x"17",x"03",x"DD",x"21",x"AF",x"40", -- 0x0FF0
    x"3A",x"00",x"60",x"CB",x"67",x"C2",x"3A",x"10", -- 0x0FF8
    x"DD",x"CB",x"00",x"46",x"28",x"27",x"DD",x"7E", -- 0x1000
    x"01",x"FE",x"99",x"28",x"1C",x"DD",x"35",x"02", -- 0x1008
    x"20",x"17",x"DD",x"7E",x"01",x"C6",x"01",x"27", -- 0x1010
    x"DD",x"77",x"01",x"DD",x"7E",x"03",x"DD",x"77", -- 0x1018
    x"02",x"CD",x"9E",x"12",x"21",x"D9",x"40",x"CB", -- 0x1020
    x"D6",x"DD",x"CB",x"00",x"86",x"DD",x"7E",x"01", -- 0x1028
    x"A7",x"C8",x"DD",x"CB",x"00",x"5E",x"CA",x"18", -- 0x1030
    x"01",x"C9",x"DD",x"CB",x"00",x"C6",x"18",x"ED", -- 0x1038
    x"21",x"CB",x"41",x"36",x"02",x"23",x"23",x"06", -- 0x1040
    x"18",x"3E",x"04",x"77",x"23",x"23",x"10",x"FB", -- 0x1048
    x"21",x"C2",x"10",x"11",x"04",x"42",x"01",x"10", -- 0x1050
    x"00",x"ED",x"B0",x"3A",x"AF",x"40",x"CB",x"67", -- 0x1058
    x"28",x"0A",x"21",x"04",x"42",x"35",x"35",x"21", -- 0x1060
    x"08",x"42",x"35",x"35",x"11",x"E0",x"FF",x"21", -- 0x1068
    x"0E",x"11",x"FD",x"21",x"A5",x"53",x"06",x"08", -- 0x1070
    x"CD",x"73",x"04",x"21",x"BC",x"10",x"11",x"D2", -- 0x1078
    x"41",x"06",x"06",x"7E",x"12",x"13",x"13",x"12", -- 0x1080
    x"13",x"13",x"13",x"13",x"23",x"10",x"F4",x"21", -- 0x1088
    x"A9",x"53",x"DD",x"21",x"D2",x"10",x"06",x"1E", -- 0x1090
    x"E5",x"C5",x"DD",x"5E",x"00",x"DD",x"23",x"DD", -- 0x1098
    x"56",x"00",x"DD",x"23",x"06",x"06",x"73",x"23", -- 0x10A0
    x"72",x"23",x"23",x"10",x"F9",x"C1",x"E1",x"11", -- 0x10A8
    x"E0",x"FF",x"19",x"10",x"E3",x"21",x"99",x"99", -- 0x10B0
    x"22",x"27",x"40",x"C9",x"20",x"90",x"F7",x"63", -- 0x10B8
    x"AA",x"00",x"31",x"33",x"02",x"30",x"21",x"B3", -- 0x10C0
    x"02",x"30",x"10",x"97",x"02",x"30",x"40",x"17", -- 0x10C8
    x"02",x"30",x"10",x"0C",x"CA",x"CB",x"C8",x"C9", -- 0x10D0
    x"0C",x"10",x"10",x"0E",x"0C",x"0D",x"10",x"10", -- 0x10D8
    x"CA",x"CB",x"C8",x"C9",x"10",x"10",x"0D",x"0C", -- 0x10E0
    x"10",x"0E",x"0C",x"10",x"CA",x"CB",x"C8",x"C9", -- 0x10E8
    x"0E",x"10",x"CA",x"CB",x"C8",x"C9",x"0C",x"10", -- 0x10F0
    x"0E",x"0D",x"10",x"0C",x"CA",x"CB",x"C8",x"C9", -- 0x10F8
    x"CA",x"CB",x"C8",x"C9",x"0C",x"0E",x"0C",x"0D", -- 0x1100
    x"0E",x"10",x"0D",x"0C",x"0C",x"10",x"64",x"66", -- 0x1108
    x"18",x"1F",x"1D",x"15",x"67",x"65",x"03",x"00", -- 0x1110
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1118
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1120
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1128
    x"00",x"00",x"00",x"03",x"01",x"0F",x"10",x"0A", -- 0x1130
    x"13",x"08",x"17",x"19",x"20",x"99",x"99",x"01", -- 0x1138
    x"00",x"3C",x"00",x"01",x"15",x"03",x"03",x"23", -- 0x1140
    x"02",x"0A",x"32",x"FF",x"10",x"00",x"00",x"00", -- 0x1148
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1150
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1158
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1160
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1168
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1170
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1178
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1180
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1188
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1190
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1198
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x11A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x11A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x11B0
    x"00",x"00",x"00",x"00",x"00",x"AA",x"02",x"00", -- 0x11B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01", -- 0x11C0
    x"01",x"00",x"50",x"00",x"00",x"00",x"01",x"00", -- 0x11C8
    x"00",x"01",x"00",x"01",x"00",x"00",x"00",x"00", -- 0x11D0
    x"00",x"03",x"00",x"00",x"00",x"00",x"00",x"01", -- 0x11D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"01", -- 0x11E0
    x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00", -- 0x11E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x11F0
    x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x11F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1200
    x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00", -- 0x1208
    x"00",x"00",x"00",x"00",x"00",x"00",x"21",x"23", -- 0x1210
    x"12",x"FD",x"21",x"A0",x"53",x"06",x"1C",x"CD", -- 0x1218
    x"3F",x"12",x"C9",x"53",x"43",x"4F",x"52",x"45", -- 0x1220
    x"5B",x"31",x"40",x"40",x"48",x"49",x"47",x"48", -- 0x1228
    x"40",x"53",x"43",x"4F",x"52",x"45",x"40",x"40", -- 0x1230
    x"53",x"43",x"4F",x"52",x"45",x"5B",x"32",x"11", -- 0x1238
    x"E0",x"FF",x"7E",x"23",x"D6",x"30",x"FD",x"77", -- 0x1240
    x"00",x"FD",x"19",x"10",x"F5",x"C9",x"21",x"A9", -- 0x1248
    x"40",x"FD",x"21",x"81",x"53",x"18",x"12",x"21", -- 0x1250
    x"AC",x"40",x"FD",x"21",x"01",x"51",x"18",x"09", -- 0x1258
    x"21",x"B3",x"40",x"FD",x"21",x"41",x"52",x"18", -- 0x1260
    x"00",x"06",x"03",x"11",x"E0",x"FF",x"0E",x"00", -- 0x1268
    x"7E",x"F5",x"1F",x"1F",x"1F",x"1F",x"CD",x"8A", -- 0x1270
    x"12",x"78",x"FE",x"01",x"CC",x"87",x"12",x"F1", -- 0x1278
    x"CD",x"8A",x"12",x"23",x"10",x"EA",x"C9",x"CB", -- 0x1280
    x"C1",x"C9",x"E6",x"0F",x"20",x"0C",x"CB",x"41", -- 0x1288
    x"20",x"08",x"3E",x"10",x"FD",x"77",x"00",x"FD", -- 0x1290
    x"19",x"C9",x"CB",x"C1",x"18",x"F6",x"FD",x"21", -- 0x1298
    x"7F",x"50",x"21",x"B0",x"40",x"06",x"01",x"C3", -- 0x12A0
    x"6B",x"12",x"21",x"16",x"11",x"11",x"00",x"40", -- 0x12A8
    x"01",x"A9",x"00",x"ED",x"B0",x"C9",x"DD",x"21", -- 0x12B0
    x"C0",x"41",x"DD",x"36",x"00",x"00",x"DD",x"36", -- 0x12B8
    x"01",x"03",x"CD",x"16",x"12",x"DD",x"36",x"02", -- 0x12C0
    x"00",x"DD",x"36",x"03",x"01",x"CD",x"4E",x"12", -- 0x12C8
    x"CD",x"57",x"12",x"CD",x"60",x"12",x"DD",x"36", -- 0x12D0
    x"3E",x"00",x"DD",x"36",x"3F",x"01",x"21",x"EE", -- 0x12D8
    x"12",x"FD",x"21",x"5F",x"51",x"06",x"06",x"CD", -- 0x12E0
    x"3F",x"12",x"CD",x"9E",x"12",x"C9",x"43",x"52", -- 0x12E8
    x"45",x"44",x"49",x"54",x"21",x"00",x"50",x"01", -- 0x12F0
    x"00",x"04",x"36",x"10",x"23",x"0B",x"79",x"B0", -- 0x12F8
    x"20",x"F8",x"21",x"C0",x"41",x"06",x"FF",x"36", -- 0x1300
    x"00",x"23",x"10",x"FB",x"21",x"00",x"42",x"06", -- 0x1308
    x"40",x"36",x"00",x"23",x"10",x"FB",x"C9",x"11", -- 0x1310
    x"03",x"00",x"21",x"02",x"50",x"0E",x"20",x"06", -- 0x1318
    x"1D",x"36",x"10",x"23",x"10",x"FB",x"19",x"0D", -- 0x1320
    x"20",x"F5",x"CD",x"0C",x"13",x"21",x"C4",x"41", -- 0x1328
    x"06",x"1D",x"AF",x"77",x"23",x"10",x"FC",x"C9", -- 0x1330
    x"32",x"B6",x"40",x"3A",x"B6",x"40",x"A7",x"C8", -- 0x1338
    x"18",x"F9",x"3E",x"FF",x"32",x"01",x"70",x"C9", -- 0x1340
    x"3A",x"AF",x"40",x"CB",x"57",x"20",x"23",x"CB", -- 0x1348
    x"6F",x"20",x"1B",x"3A",x"00",x"70",x"CB",x"5F", -- 0x1350
    x"28",x"14",x"3A",x"00",x"68",x"CB",x"3F",x"CB", -- 0x1358
    x"3F",x"47",x"CB",x"A8",x"3A",x"00",x"60",x"CB", -- 0x1360
    x"77",x"78",x"C8",x"CB",x"EF",x"C9",x"3A",x"00", -- 0x1368
    x"60",x"C9",x"21",x"B7",x"40",x"7E",x"23",x"35", -- 0x1370
    x"C0",x"23",x"5E",x"23",x"56",x"13",x"23",x"35", -- 0x1378
    x"20",x"05",x"11",x"96",x"13",x"36",x"14",x"1A", -- 0x1380
    x"47",x"13",x"1A",x"CB",x"EF",x"2B",x"72",x"2B", -- 0x1388
    x"73",x"2B",x"70",x"2B",x"77",x"C9",x"50",x"02", -- 0x1390
    x"5A",x"04",x"3C",x"09",x"46",x"00",x"28",x"02", -- 0x1398
    x"50",x"08",x"5A",x"00",x"5A",x"06",x"50",x"09", -- 0x13A0
    x"4B",x"0A",x"41",x"00",x"05",x"01",x"05",x"02", -- 0x13A8
    x"05",x"04",x"05",x"08",x"5A",x"01",x"50",x"02", -- 0x13B0
    x"46",x"05",x"63",x"01",x"63",x"05",x"3E",x"00", -- 0x13B8
    x"32",x"01",x"70",x"C9",x"11",x"00",x"42",x"21", -- 0x13C0
    x"FF",x"13",x"3A",x"1E",x"40",x"E6",x"03",x"20", -- 0x13C8
    x"03",x"21",x"03",x"14",x"01",x"04",x"00",x"ED", -- 0x13D0
    x"B0",x"21",x"1D",x"40",x"35",x"11",x"E0",x"FF", -- 0x13D8
    x"21",x"9F",x"53",x"06",x"06",x"3E",x"10",x"77", -- 0x13E0
    x"19",x"10",x"FC",x"3A",x"1D",x"40",x"32",x"BF", -- 0x13E8
    x"53",x"A7",x"28",x"0A",x"47",x"21",x"9F",x"53", -- 0x13F0
    x"3E",x"0F",x"77",x"19",x"10",x"FC",x"C9",x"80", -- 0x13F8
    x"10",x"01",x"80",x"E0",x"11",x"01",x"E0",x"E9", -- 0x1400
    x"3A",x"01",x"40",x"CB",x"47",x"C0",x"DD",x"21", -- 0x1408
    x"20",x"42",x"FD",x"21",x"06",x"40",x"06",x"04", -- 0x1410
    x"FD",x"7E",x"00",x"A7",x"28",x"45",x"DD",x"7E", -- 0x1418
    x"03",x"ED",x"44",x"D6",x"14",x"6F",x"DD",x"66", -- 0x1420
    x"01",x"0E",x"00",x"DD",x"E5",x"FD",x"E5",x"C5", -- 0x1428
    x"3A",x"1E",x"40",x"E6",x"03",x"CA",x"6C",x"15", -- 0x1430
    x"FD",x"21",x"04",x"42",x"DD",x"21",x"37",x"40", -- 0x1438
    x"06",x"07",x"DD",x"CB",x"00",x"4E",x"C4",x"70", -- 0x1440
    x"14",x"CD",x"78",x"09",x"10",x"F4",x"79",x"C1", -- 0x1448
    x"FD",x"E1",x"DD",x"E1",x"CB",x"47",x"28",x"0B", -- 0x1450
    x"AF",x"DD",x"77",x"01",x"DD",x"77",x"03",x"FD", -- 0x1458
    x"36",x"00",x"00",x"11",x"08",x"00",x"DD",x"19", -- 0x1460
    x"11",x"04",x"00",x"FD",x"19",x"10",x"A9",x"C9", -- 0x1468
    x"7C",x"FD",x"96",x"00",x"FE",x"10",x"D0",x"57", -- 0x1470
    x"7D",x"FD",x"96",x"03",x"ED",x"44",x"FE",x"10", -- 0x1478
    x"D0",x"5F",x"E5",x"21",x"AC",x"14",x"FD",x"7E", -- 0x1480
    x"01",x"D6",x"13",x"87",x"87",x"87",x"87",x"87", -- 0x1488
    x"CB",x"22",x"82",x"85",x"6F",x"3E",x"00",x"8C", -- 0x1490
    x"67",x"7B",x"BE",x"30",x"0D",x"23",x"BE",x"38", -- 0x1498
    x"09",x"0E",x"FF",x"CD",x"EB",x"18",x"DD",x"CB", -- 0x14A0
    x"00",x"C6",x"E1",x"C9",x"07",x"00",x"07",x"00", -- 0x14A8
    x"07",x"00",x"07",x"00",x"07",x"00",x"07",x"00", -- 0x14B0
    x"07",x"00",x"07",x"00",x"32",x"32",x"32",x"32", -- 0x14B8
    x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"32", -- 0x14C0
    x"32",x"32",x"32",x"32",x"07",x"00",x"07",x"00", -- 0x14C8
    x"07",x"00",x"07",x"00",x"07",x"00",x"07",x"00", -- 0x14D0
    x"07",x"00",x"07",x"00",x"32",x"32",x"32",x"32", -- 0x14D8
    x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"32", -- 0x14E0
    x"32",x"32",x"32",x"32",x"08",x"07",x"09",x"06", -- 0x14E8
    x"0A",x"05",x"0B",x"04",x"0C",x"03",x"0D",x"02", -- 0x14F0
    x"0E",x"01",x"0F",x"00",x"0F",x"00",x"0E",x"01", -- 0x14F8
    x"0D",x"02",x"0C",x"03",x"0B",x"04",x"0A",x"05", -- 0x1500
    x"09",x"06",x"08",x"07",x"00",x"00",x"00",x"00", -- 0x1508
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1510
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1518
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1520
    x"00",x"00",x"00",x"00",x"0F",x"00",x"0F",x"00", -- 0x1528
    x"0F",x"00",x"0F",x"00",x"0F",x"00",x"0F",x"00", -- 0x1530
    x"0F",x"00",x"0F",x"00",x"0F",x"00",x"0F",x"00", -- 0x1538
    x"0F",x"01",x"0F",x"02",x"0F",x"03",x"0F",x"04", -- 0x1540
    x"0F",x"05",x"0F",x"06",x"0C",x"03",x"0C",x"03", -- 0x1548
    x"0C",x"03",x"0C",x"03",x"0D",x"02",x"0E",x"01", -- 0x1550
    x"0F",x"00",x"0F",x"00",x"0F",x"00",x"0F",x"00", -- 0x1558
    x"0E",x"01",x"0D",x"02",x"0C",x"03",x"0C",x"03", -- 0x1560
    x"0C",x"03",x"0C",x"03",x"EB",x"7A",x"2F",x"57", -- 0x1568
    x"1D",x"1D",x"1D",x"CD",x"64",x"16",x"7E",x"FE", -- 0x1570
    x"10",x"28",x"44",x"E5",x"FD",x"E1",x"C5",x"D5", -- 0x1578
    x"21",x"B9",x"16",x"11",x"11",x"00",x"06",x"07", -- 0x1580
    x"BE",x"28",x"07",x"19",x"10",x"FA",x"D1",x"C1", -- 0x1588
    x"18",x"2D",x"23",x"D1",x"C1",x"78",x"CB",x"27", -- 0x1590
    x"85",x"6F",x"3E",x"00",x"8C",x"67",x"79",x"BE", -- 0x1598
    x"28",x"03",x"D2",x"BF",x"15",x"23",x"BE",x"DA", -- 0x15A0
    x"BF",x"15",x"D5",x"FD",x"7E",x"00",x"FE",x"0C", -- 0x15A8
    x"28",x"12",x"FE",x"0E",x"28",x"18",x"FE",x"0D", -- 0x15B0
    x"28",x"2A",x"E6",x"F8",x"20",x"3C",x"D1",x"0E", -- 0x15B8
    x"00",x"C3",x"4E",x"14",x"FD",x"36",x"00",x"10", -- 0x15C0
    x"11",x"00",x"01",x"C3",x"27",x"16",x"FD",x"36", -- 0x15C8
    x"00",x"10",x"11",x"50",x"00",x"FD",x"7E",x"E0", -- 0x15D0
    x"FE",x"0D",x"C2",x"27",x"16",x"FD",x"36",x"E0", -- 0x15D8
    x"10",x"C3",x"27",x"16",x"FD",x"36",x"00",x"10", -- 0x15E0
    x"11",x"50",x"00",x"FD",x"7E",x"20",x"FE",x"0E", -- 0x15E8
    x"C2",x"27",x"16",x"FD",x"36",x"20",x"10",x"C3", -- 0x15F0
    x"27",x"16",x"FD",x"7E",x"00",x"21",x"9B",x"16", -- 0x15F8
    x"06",x"04",x"BE",x"28",x"06",x"23",x"23",x"23", -- 0x1600
    x"10",x"F8",x"C7",x"23",x"5E",x"23",x"56",x"FD", -- 0x1608
    x"19",x"FD",x"36",x"00",x"10",x"FD",x"36",x"01", -- 0x1610
    x"10",x"FD",x"36",x"20",x"10",x"FD",x"36",x"21", -- 0x1618
    x"10",x"11",x"30",x"00",x"C3",x"27",x"16",x"CD", -- 0x1620
    x"72",x"19",x"DD",x"21",x"77",x"40",x"FD",x"21", -- 0x1628
    x"14",x"42",x"06",x"03",x"DD",x"CB",x"00",x"46", -- 0x1630
    x"28",x"0B",x"CD",x"78",x"09",x"10",x"F5",x"0E", -- 0x1638
    x"01",x"D1",x"C3",x"4E",x"14",x"DD",x"36",x"00", -- 0x1640
    x"01",x"FD",x"36",x"01",x"1C",x"FD",x"36",x"02", -- 0x1648
    x"06",x"D1",x"7A",x"2F",x"D6",x"08",x"FD",x"77", -- 0x1650
    x"00",x"3E",x"08",x"83",x"FD",x"77",x"03",x"0E", -- 0x1658
    x"01",x"C3",x"4E",x"14",x"7B",x"E6",x"07",x"4F", -- 0x1660
    x"3E",x"07",x"91",x"4F",x"7B",x"E6",x"F8",x"C6", -- 0x1668
    x"10",x"CB",x"3F",x"CB",x"3F",x"F5",x"21",x"C0", -- 0x1670
    x"41",x"85",x"6F",x"3E",x"00",x"8C",x"67",x"7A", -- 0x1678
    x"86",x"47",x"E6",x"F8",x"6F",x"78",x"E6",x"07", -- 0x1680
    x"47",x"26",x"00",x"29",x"29",x"F1",x"CB",x"3F", -- 0x1688
    x"85",x"6F",x"3E",x"00",x"85",x"6F",x"3E",x"50", -- 0x1690
    x"8C",x"67",x"C9",x"C8",x"00",x"00",x"C9",x"FF", -- 0x1698
    x"FF",x"CA",x"E0",x"FF",x"CB",x"DF",x"FF",x"B9", -- 0x16A0
    x"A9",x"17",x"A1",x"91",x"14",x"89",x"79",x"11", -- 0x16A8
    x"71",x"61",x"0E",x"59",x"49",x"0B",x"41",x"31", -- 0x16B0
    x"08",x"0D",x"04",x"00",x"06",x"00",x"06",x"00", -- 0x16B8
    x"06",x"00",x"06",x"00",x"06",x"00",x"06",x"00", -- 0x16C0
    x"07",x"00",x"0E",x"07",x"00",x"07",x"00",x"07", -- 0x16C8
    x"00",x"07",x"00",x"07",x"00",x"07",x"00",x"05", -- 0x16D0
    x"00",x"05",x"00",x"C8",x"00",x"00",x"00",x"03", -- 0x16D8
    x"00",x"03",x"00",x"04",x"00",x"04",x"00",x"02", -- 0x16E0
    x"00",x"04",x"00",x"05",x"C9",x"07",x"05",x"07", -- 0x16E8
    x"02",x"07",x"00",x"07",x"00",x"07",x"00",x"07", -- 0x16F0
    x"00",x"07",x"00",x"07",x"01",x"CA",x"05",x"00", -- 0x16F8
    x"06",x"00",x"06",x"00",x"05",x"00",x"04",x"00", -- 0x1700
    x"04",x"00",x"03",x"00",x"01",x"00",x"CB",x"07", -- 0x1708
    x"01",x"07",x"02",x"07",x"02",x"07",x"02",x"07", -- 0x1710
    x"02",x"07",x"03",x"07",x"06",x"07",x"06",x"0C", -- 0x1718
    x"32",x"32",x"07",x"01",x"07",x"01",x"07",x"01", -- 0x1720
    x"07",x"01",x"07",x"01",x"07",x"01",x"07",x"01", -- 0x1728
    x"3A",x"01",x"40",x"CB",x"47",x"C0",x"FD",x"21", -- 0x1730
    x"00",x"42",x"21",x"1B",x"18",x"11",x"15",x"00", -- 0x1738
    x"FD",x"7E",x"01",x"BE",x"28",x"03",x"19",x"18", -- 0x1740
    x"FA",x"06",x"0A",x"23",x"FD",x"7E",x"00",x"86", -- 0x1748
    x"ED",x"44",x"57",x"FD",x"7E",x"03",x"23",x"96", -- 0x1750
    x"23",x"5F",x"E5",x"C5",x"CD",x"64",x"16",x"7E", -- 0x1758
    x"FE",x"10",x"CA",x"14",x"18",x"E5",x"DD",x"E1", -- 0x1760
    x"C5",x"D5",x"21",x"B9",x"16",x"11",x"11",x"00", -- 0x1768
    x"06",x"07",x"BE",x"28",x"08",x"19",x"10",x"FA", -- 0x1770
    x"D1",x"C1",x"C3",x"14",x"18",x"23",x"D1",x"C1", -- 0x1778
    x"78",x"CB",x"27",x"85",x"6F",x"3E",x"00",x"8C", -- 0x1780
    x"67",x"79",x"BE",x"D2",x"14",x"18",x"23",x"BE", -- 0x1788
    x"DA",x"14",x"18",x"DD",x"7E",x"00",x"FE",x"0C", -- 0x1790
    x"28",x"0F",x"FE",x"0E",x"28",x"15",x"FE",x"0D", -- 0x1798
    x"28",x"27",x"E6",x"F8",x"20",x"39",x"C3",x"14", -- 0x17A0
    x"18",x"DD",x"36",x"00",x"10",x"11",x"00",x"01", -- 0x17A8
    x"C3",x"09",x"18",x"DD",x"36",x"00",x"10",x"11", -- 0x17B0
    x"50",x"00",x"DD",x"7E",x"E0",x"FE",x"0D",x"C2", -- 0x17B8
    x"09",x"18",x"DD",x"36",x"E0",x"10",x"C3",x"09", -- 0x17C0
    x"18",x"DD",x"36",x"00",x"10",x"11",x"50",x"00", -- 0x17C8
    x"DD",x"7E",x"20",x"FE",x"0E",x"C2",x"09",x"18", -- 0x17D0
    x"DD",x"36",x"20",x"10",x"C3",x"09",x"18",x"DD", -- 0x17D8
    x"7E",x"00",x"21",x"9B",x"16",x"06",x"04",x"BE", -- 0x17E0
    x"28",x"06",x"23",x"23",x"23",x"10",x"F8",x"C7", -- 0x17E8
    x"23",x"5E",x"23",x"56",x"DD",x"19",x"DD",x"36", -- 0x17F0
    x"00",x"10",x"DD",x"36",x"01",x"10",x"DD",x"36", -- 0x17F8
    x"20",x"10",x"DD",x"36",x"21",x"10",x"11",x"30", -- 0x1800
    x"00",x"CD",x"72",x"19",x"21",x"01",x"40",x"CB", -- 0x1808
    x"C6",x"C1",x"E1",x"C9",x"C1",x"E1",x"05",x"C2", -- 0x1810
    x"4C",x"17",x"C9",x"10",x"00",x"01",x"00",x"05", -- 0x1818
    x"02",x"01",x"03",x"09",x"06",x"03",x"06",x"0C", -- 0x1820
    x"0A",x"09",x"0B",x"02",x"0D",x"02",x"0D",x"06", -- 0x1828
    x"50",x"09",x"03",x"06",x"06",x"0C",x"06",x"03", -- 0x1830
    x"0A",x"0F",x"0A",x"09",x"0C",x"03",x"0E",x"05", -- 0x1838
    x"0E",x"0D",x"0E",x"0F",x"0E",x"11",x"00",x"03", -- 0x1840
    x"00",x"05",x"00",x"0B",x"00",x"0D",x"02",x"08", -- 0x1848
    x"05",x"03",x"05",x"0D",x"0C",x"05",x"0C",x"0B", -- 0x1850
    x"0F",x"08",x"D2",x"0F",x"04",x"0D",x"06",x"0C", -- 0x1858
    x"02",x"09",x"06",x"08",x"09",x"06",x"0B",x"03", -- 0x1860
    x"09",x"00",x"04",x"00",x"00",x"06",x"00",x"91", -- 0x1868
    x"0F",x"03",x"0F",x"05",x"0F",x"0B",x"0F",x"0D", -- 0x1870
    x"0D",x"08",x"0A",x"03",x"0A",x"0D",x"03",x"05", -- 0x1878
    x"03",x"0B",x"00",x"08",x"12",x"00",x"0B",x"02", -- 0x1880
    x"09",x"03",x"0D",x"06",x"09",x"07",x"06",x"09", -- 0x1888
    x"04",x"0C",x"06",x"0F",x"0B",x"0F",x"0F",x"09", -- 0x1890
    x"0F",x"92",x"0F",x"0B",x"0D",x"09",x"0C",x"0D", -- 0x1898
    x"09",x"09",x"08",x"06",x"06",x"04",x"03",x"06", -- 0x18A0
    x"00",x"0B",x"00",x"0F",x"06",x"0F",x"52",x"00", -- 0x18A8
    x"04",x"02",x"06",x"03",x"02",x"06",x"06",x"07", -- 0x18B0
    x"09",x"09",x"0B",x"0C",x"09",x"0F",x"04",x"00", -- 0x18B8
    x"00",x"09",x"00",x"CD",x"48",x"1B",x"CD",x"E7", -- 0x18C0
    x"1D",x"3A",x"1E",x"40",x"E6",x"03",x"28",x"09", -- 0x18C8
    x"CD",x"D6",x"1C",x"CD",x"DD",x"0E",x"C3",x"B4", -- 0x18D0
    x"00",x"CD",x"81",x"1A",x"CD",x"FF",x"19",x"CD", -- 0x18D8
    x"AE",x"1A",x"CD",x"E7",x"1A",x"CD",x"CA",x"1D", -- 0x18E0
    x"C3",x"B4",x"00",x"DD",x"CB",x"00",x"46",x"C0", -- 0x18E8
    x"3A",x"AF",x"40",x"CB",x"57",x"C0",x"FD",x"E5", -- 0x18F0
    x"C5",x"47",x"FD",x"7E",x"01",x"D6",x"13",x"CB", -- 0x18F8
    x"27",x"5F",x"16",x"00",x"21",x"39",x"19",x"19", -- 0x1900
    x"5E",x"23",x"56",x"EB",x"CD",x"07",x"14",x"21", -- 0x1908
    x"AB",x"40",x"CB",x"68",x"F5",x"20",x"03",x"21", -- 0x1910
    x"AE",x"40",x"7B",x"86",x"27",x"77",x"2B",x"7A", -- 0x1918
    x"8E",x"27",x"77",x"2B",x"3E",x"00",x"8E",x"27", -- 0x1920
    x"77",x"21",x"4E",x"12",x"F1",x"20",x"03",x"21", -- 0x1928
    x"57",x"12",x"CD",x"07",x"14",x"C1",x"FD",x"E1", -- 0x1930
    x"C9",x"45",x"19",x"4E",x"19",x"57",x"19",x"00", -- 0x1938
    x"00",x"00",x"00",x"69",x"19",x"11",x"00",x"02", -- 0x1940
    x"21",x"EE",x"40",x"CB",x"DE",x"C9",x"11",x"53", -- 0x1948
    x"00",x"21",x"EE",x"40",x"CB",x"DE",x"C9",x"21", -- 0x1950
    x"EE",x"40",x"CB",x"D6",x"FD",x"7E",x"02",x"11", -- 0x1958
    x"00",x"01",x"FE",x"06",x"C8",x"11",x"50",x"01", -- 0x1960
    x"C9",x"11",x"00",x"01",x"21",x"EE",x"40",x"CB", -- 0x1968
    x"D6",x"C9",x"3A",x"AF",x"40",x"CB",x"57",x"C0", -- 0x1970
    x"47",x"FD",x"E5",x"C5",x"C3",x"0F",x"19",x"3A", -- 0x1978
    x"01",x"40",x"CB",x"47",x"C0",x"FD",x"21",x"24", -- 0x1980
    x"42",x"06",x"04",x"DD",x"21",x"00",x"42",x"C5", -- 0x1988
    x"FD",x"7E",x"01",x"DD",x"96",x"00",x"FE",x"10", -- 0x1990
    x"30",x"5C",x"4F",x"FD",x"7E",x"03",x"2F",x"D6", -- 0x1998
    x"50",x"47",x"DD",x"7E",x"03",x"90",x"FA",x"AE", -- 0x19A0
    x"19",x"FE",x"10",x"30",x"49",x"AF",x"47",x"FD", -- 0x19A8
    x"7E",x"03",x"2F",x"D6",x"70",x"DD",x"96",x"03", -- 0x19B0
    x"F2",x"F6",x"19",x"FE",x"10",x"38",x"02",x"3E", -- 0x19B8
    x"10",x"F5",x"21",x"D9",x"0C",x"3A",x"01",x"42", -- 0x19C0
    x"BE",x"28",x"05",x"23",x"23",x"23",x"18",x"F8", -- 0x19C8
    x"23",x"5E",x"23",x"56",x"EB",x"79",x"CB",x"27", -- 0x19D0
    x"85",x"6F",x"3E",x"00",x"8C",x"67",x"F1",x"5F", -- 0x19D8
    x"78",x"C6",x"20",x"BE",x"D2",x"F6",x"19",x"23", -- 0x19E0
    x"7B",x"C6",x"20",x"BE",x"DA",x"F6",x"19",x"21", -- 0x19E8
    x"01",x"40",x"CB",x"C6",x"C1",x"C9",x"11",x"08", -- 0x19F0
    x"00",x"FD",x"19",x"C1",x"10",x"91",x"C9",x"DD", -- 0x19F8
    x"21",x"24",x"42",x"FD",x"21",x"2C",x"42",x"01", -- 0x1A00
    x"09",x"02",x"3A",x"29",x"40",x"5F",x"DD",x"7E", -- 0x1A08
    x"01",x"A7",x"F5",x"C4",x"35",x"1A",x"F1",x"CC", -- 0x1A10
    x"57",x"1A",x"FD",x"7E",x"01",x"A7",x"F5",x"C4", -- 0x1A18
    x"46",x"1A",x"F1",x"CC",x"6C",x"1A",x"05",x"C8", -- 0x1A20
    x"D5",x"11",x"10",x"00",x"DD",x"19",x"FD",x"19", -- 0x1A28
    x"D1",x"0E",x"35",x"18",x"D9",x"DD",x"7E",x"03", -- 0x1A30
    x"93",x"DD",x"77",x"03",x"D0",x"DD",x"36",x"01", -- 0x1A38
    x"00",x"DD",x"36",x"03",x"00",x"C9",x"FD",x"7E", -- 0x1A40
    x"03",x"93",x"FD",x"77",x"03",x"D0",x"FD",x"36", -- 0x1A48
    x"01",x"00",x"FD",x"36",x"03",x"00",x"C9",x"FD", -- 0x1A50
    x"7E",x"03",x"FE",x"2C",x"D0",x"DD",x"36",x"03", -- 0x1A58
    x"5E",x"21",x"0C",x"42",x"7E",x"81",x"3C",x"3C", -- 0x1A60
    x"DD",x"77",x"01",x"C9",x"DD",x"7E",x"03",x"FE", -- 0x1A68
    x"2C",x"D0",x"FD",x"36",x"03",x"5E",x"21",x"0C", -- 0x1A70
    x"42",x"7E",x"81",x"3D",x"3D",x"FD",x"77",x"01", -- 0x1A78
    x"C9",x"11",x"D2",x"41",x"FD",x"21",x"20",x"40", -- 0x1A80
    x"21",x"D2",x"40",x"06",x"06",x"0E",x"01",x"35", -- 0x1A88
    x"28",x"10",x"13",x"13",x"13",x"13",x"13",x"13", -- 0x1A90
    x"79",x"ED",x"44",x"4F",x"23",x"FD",x"23",x"10", -- 0x1A98
    x"EE",x"C9",x"FD",x"7E",x"00",x"77",x"1A",x"81", -- 0x1AA0
    x"12",x"13",x"13",x"12",x"18",x"E6",x"21",x"D8", -- 0x1AA8
    x"40",x"35",x"C0",x"3A",x"26",x"40",x"77",x"FD", -- 0x1AB0
    x"21",x"04",x"42",x"11",x"04",x"00",x"06",x"04", -- 0x1AB8
    x"21",x"D1",x"40",x"4E",x"FD",x"7E",x"00",x"81", -- 0x1AC0
    x"FD",x"77",x"00",x"FE",x"10",x"DC",x"E0",x"1A", -- 0x1AC8
    x"FE",x"E0",x"D4",x"E0",x"1A",x"FD",x"19",x"10", -- 0x1AD0
    x"EB",x"21",x"CA",x"41",x"7E",x"81",x"77",x"C9", -- 0x1AD8
    x"F5",x"7E",x"ED",x"44",x"77",x"F1",x"C9",x"3A", -- 0x1AE0
    x"01",x"40",x"CB",x"47",x"C0",x"3A",x"B6",x"40", -- 0x1AE8
    x"A7",x"F0",x"3A",x"2B",x"40",x"32",x"B6",x"40", -- 0x1AF0
    x"3A",x"65",x"53",x"FE",x"18",x"28",x"11",x"21", -- 0x1AF8
    x"0C",x"1B",x"FD",x"21",x"65",x"53",x"06",x"04", -- 0x1B00
    x"CD",x"3F",x"12",x"C9",x"48",x"4F",x"4D",x"45", -- 0x1B08
    x"FD",x"21",x"05",x"53",x"21",x"28",x"40",x"7E", -- 0x1B10
    x"D6",x"99",x"27",x"77",x"F5",x"AF",x"ED",x"67", -- 0x1B18
    x"FD",x"77",x"00",x"ED",x"67",x"FD",x"77",x"20", -- 0x1B20
    x"ED",x"67",x"2B",x"F1",x"7E",x"DE",x"00",x"27", -- 0x1B28
    x"77",x"AF",x"ED",x"67",x"FD",x"77",x"40",x"ED", -- 0x1B30
    x"67",x"FD",x"77",x"60",x"ED",x"67",x"7E",x"23", -- 0x1B38
    x"B6",x"C0",x"21",x"01",x"40",x"CB",x"C6",x"C9", -- 0x1B40
    x"DD",x"21",x"00",x"40",x"FD",x"21",x"00",x"42", -- 0x1B48
    x"DD",x"CB",x"01",x"46",x"C2",x"FD",x"1B",x"CD", -- 0x1B50
    x"48",x"13",x"E6",x"0F",x"DD",x"BE",x"02",x"C4", -- 0x1B58
    x"90",x"1B",x"FD",x"7E",x"03",x"DD",x"86",x"03", -- 0x1B60
    x"21",x"CE",x"1C",x"F5",x"3A",x"1E",x"40",x"E6", -- 0x1B68
    x"03",x"20",x"03",x"21",x"D2",x"1C",x"F1",x"BE", -- 0x1B70
    x"D0",x"23",x"BE",x"D8",x"23",x"47",x"FD",x"7E", -- 0x1B78
    x"00",x"DD",x"86",x"04",x"BE",x"D0",x"23",x"BE", -- 0x1B80
    x"D8",x"FD",x"77",x"00",x"FD",x"70",x"03",x"C9", -- 0x1B88
    x"DD",x"4E",x"02",x"DD",x"77",x"02",x"21",x"D9", -- 0x1B90
    x"1B",x"11",x"E2",x"1B",x"06",x"09",x"BE",x"28", -- 0x1B98
    x"07",x"23",x"13",x"13",x"13",x"10",x"F7",x"C9", -- 0x1BA0
    x"1A",x"A7",x"28",x"03",x"FD",x"77",x"01",x"13", -- 0x1BA8
    x"1A",x"DD",x"77",x"03",x"13",x"1A",x"DD",x"77", -- 0x1BB0
    x"04",x"3A",x"1E",x"40",x"E6",x"03",x"C0",x"CB", -- 0x1BB8
    x"79",x"20",x"0D",x"DD",x"CB",x"03",x"26",x"DD", -- 0x1BC0
    x"CB",x"04",x"26",x"DD",x"CB",x"02",x"FE",x"C9", -- 0x1BC8
    x"DD",x"CB",x"03",x"2E",x"DD",x"CB",x"04",x"2E", -- 0x1BD0
    x"C9",x"00",x"01",x"02",x"04",x"08",x"05",x"09", -- 0x1BD8
    x"06",x"0A",x"00",x"00",x"00",x"50",x"02",x"00", -- 0x1BE0
    x"10",x"FE",x"00",x"11",x"00",x"02",x"91",x"00", -- 0x1BE8
    x"FE",x"52",x"02",x"02",x"D2",x"02",x"FE",x"12", -- 0x1BF0
    x"FE",x"02",x"92",x"FE",x"FE",x"DD",x"CB",x"01", -- 0x1BF8
    x"56",x"C0",x"DD",x"CB",x"01",x"4E",x"CA",x"6C", -- 0x1C00
    x"1C",x"DD",x"35",x"00",x"C0",x"DD",x"36",x"00", -- 0x1C08
    x"08",x"FD",x"7E",x"02",x"FE",x"06",x"28",x"28", -- 0x1C10
    x"3E",x"04",x"FD",x"86",x"01",x"FE",x"40",x"28", -- 0x1C18
    x"33",x"FD",x"77",x"01",x"FD",x"35",x"02",x"FD", -- 0x1C20
    x"21",x"14",x"42",x"06",x"03",x"11",x"04",x"00", -- 0x1C28
    x"FD",x"7E",x"01",x"C6",x"04",x"FD",x"77",x"01", -- 0x1C30
    x"FD",x"35",x"02",x"FD",x"19",x"10",x"F1",x"C9", -- 0x1C38
    x"FD",x"34",x"02",x"FD",x"21",x"14",x"42",x"11", -- 0x1C40
    x"04",x"00",x"06",x"03",x"FD",x"34",x"02",x"FD", -- 0x1C48
    x"19",x"10",x"F9",x"C9",x"AF",x"06",x"04",x"FD", -- 0x1C50
    x"77",x"00",x"FD",x"23",x"10",x"F9",x"21",x"14", -- 0x1C58
    x"42",x"06",x"0C",x"77",x"23",x"10",x"FC",x"DD", -- 0x1C60
    x"CB",x"01",x"D6",x"C9",x"FD",x"56",x"00",x"FD", -- 0x1C68
    x"5E",x"03",x"7A",x"C6",x"08",x"FD",x"77",x"00", -- 0x1C70
    x"7B",x"D6",x"08",x"FD",x"77",x"03",x"FD",x"36", -- 0x1C78
    x"01",x"34",x"FD",x"36",x"02",x"06",x"DD",x"CB", -- 0x1C80
    x"01",x"CE",x"DD",x"36",x"00",x"08",x"21",x"D9", -- 0x1C88
    x"40",x"CB",x"C6",x"DD",x"21",x"77",x"40",x"FD", -- 0x1C90
    x"21",x"14",x"42",x"21",x"C5",x"1C",x"06",x"03", -- 0x1C98
    x"7A",x"86",x"FD",x"77",x"00",x"23",x"7E",x"FD", -- 0x1CA0
    x"77",x"01",x"23",x"FD",x"36",x"02",x"06",x"7B", -- 0x1CA8
    x"86",x"FD",x"77",x"03",x"23",x"DD",x"CB",x"00", -- 0x1CB0
    x"8E",x"DD",x"CB",x"00",x"96",x"D5",x"CD",x"78", -- 0x1CB8
    x"09",x"D1",x"10",x"DC",x"C9",x"08",x"35",x"08", -- 0x1CC0
    x"F8",x"36",x"F8",x"F8",x"37",x"08",x"D8",x"20", -- 0x1CC8
    x"D8",x"20",x"E8",x"34",x"E0",x"18",x"DD",x"21", -- 0x1CD0
    x"37",x"40",x"FD",x"21",x"04",x"42",x"DD",x"7E", -- 0x1CD8
    x"FF",x"A7",x"28",x"03",x"DD",x"35",x"FF",x"06", -- 0x1CE0
    x"07",x"DD",x"CB",x"00",x"4E",x"C5",x"C4",x"F8", -- 0x1CE8
    x"1C",x"C1",x"CD",x"78",x"09",x"10",x"F2",x"C9", -- 0x1CF0
    x"DD",x"CB",x"00",x"46",x"C2",x"1A",x"1D",x"DD", -- 0x1CF8
    x"6E",x"01",x"DD",x"66",x"02",x"CD",x"07",x"14", -- 0x1D00
    x"78",x"FD",x"86",x"00",x"FD",x"77",x"00",x"79", -- 0x1D08
    x"FD",x"86",x"03",x"FD",x"77",x"03",x"DD",x"35", -- 0x1D10
    x"0E",x"C9",x"DD",x"CB",x"00",x"5E",x"28",x"22", -- 0x1D18
    x"DD",x"35",x"05",x"C0",x"FD",x"7E",x"01",x"3C", -- 0x1D20
    x"FE",x"20",x"28",x"08",x"FD",x"77",x"01",x"DD", -- 0x1D28
    x"36",x"05",x"04",x"C9",x"AF",x"DD",x"77",x"00", -- 0x1D30
    x"FD",x"77",x"00",x"FD",x"77",x"03",x"FD",x"77", -- 0x1D38
    x"01",x"C9",x"3A",x"A7",x"40",x"32",x"36",x"40", -- 0x1D40
    x"FD",x"36",x"01",x"1C",x"FD",x"36",x"02",x"07", -- 0x1D48
    x"DD",x"36",x"05",x"04",x"DD",x"CB",x"00",x"DE", -- 0x1D50
    x"C9",x"DD",x"7E",x"0D",x"A7",x"20",x"0A",x"3A", -- 0x1D58
    x"F4",x"40",x"DD",x"77",x"0D",x"01",x"00",x"00", -- 0x1D60
    x"C9",x"DD",x"35",x"0D",x"DD",x"6E",x"03",x"DD", -- 0x1D68
    x"66",x"04",x"DD",x"35",x"05",x"20",x"0F",x"DD", -- 0x1D70
    x"35",x"06",x"23",x"7E",x"DD",x"77",x"05",x"23", -- 0x1D78
    x"DD",x"75",x"03",x"DD",x"74",x"04",x"7E",x"CB", -- 0x1D80
    x"2F",x"CB",x"2F",x"CB",x"2F",x"CB",x"2F",x"47", -- 0x1D88
    x"7E",x"E6",x"0F",x"CB",x"5F",x"28",x"02",x"F6", -- 0x1D90
    x"F0",x"4F",x"C9",x"DD",x"46",x"03",x"DD",x"4E", -- 0x1D98
    x"04",x"C9",x"CD",x"59",x"1D",x"DD",x"CB",x"0F", -- 0x1DA0
    x"46",x"28",x"04",x"78",x"ED",x"44",x"47",x"DD", -- 0x1DA8
    x"CB",x"0F",x"4E",x"28",x"04",x"79",x"ED",x"44", -- 0x1DB0
    x"4F",x"DD",x"CB",x"0F",x"56",x"28",x"02",x"CB", -- 0x1DB8
    x"20",x"DD",x"CB",x"0F",x"5E",x"28",x"02",x"CB", -- 0x1DC0
    x"21",x"C9",x"3A",x"01",x"40",x"CB",x"47",x"C0", -- 0x1DC8
    x"FD",x"21",x"14",x"42",x"DD",x"21",x"77",x"40", -- 0x1DD0
    x"06",x"03",x"DD",x"CB",x"00",x"46",x"C4",x"1A", -- 0x1DD8
    x"1D",x"CD",x"78",x"09",x"10",x"F4",x"C9",x"DD", -- 0x1DE0
    x"21",x"06",x"40",x"FD",x"21",x"20",x"42",x"06", -- 0x1DE8
    x"04",x"DD",x"7E",x"00",x"A7",x"CC",x"49",x"1E", -- 0x1DF0
    x"C4",x"0B",x"1E",x"11",x"04",x"00",x"DD",x"19", -- 0x1DF8
    x"11",x"08",x"00",x"FD",x"19",x"10",x"EA",x"CD", -- 0x1E00
    x"E9",x"1E",x"C9",x"C5",x"D5",x"DD",x"35",x"00", -- 0x1E08
    x"20",x"0F",x"FD",x"36",x"01",x"00",x"FD",x"36", -- 0x1E10
    x"03",x"00",x"DD",x"36",x"00",x"00",x"D1",x"C1", -- 0x1E18
    x"C9",x"FD",x"7E",x"03",x"FE",x"E0",x"30",x"EA", -- 0x1E20
    x"FE",x"08",x"38",x"E6",x"FD",x"7E",x"01",x"FE", -- 0x1E28
    x"F8",x"30",x"DF",x"FE",x"16",x"38",x"DB",x"DD", -- 0x1E30
    x"86",x"02",x"FD",x"77",x"01",x"FD",x"7E",x"03", -- 0x1E38
    x"DD",x"86",x"01",x"FD",x"77",x"03",x"D1",x"C1", -- 0x1E40
    x"C9",x"C5",x"D5",x"3A",x"01",x"40",x"CB",x"47", -- 0x1E48
    x"C2",x"46",x"1E",x"CD",x"48",x"13",x"CB",x"6F", -- 0x1E50
    x"CA",x"46",x"1E",x"21",x"06",x"40",x"06",x"04", -- 0x1E58
    x"11",x"04",x"00",x"0E",x"1C",x"3A",x"1E",x"40", -- 0x1E60
    x"E6",x"03",x"20",x"02",x"0E",x"01",x"79",x"BE", -- 0x1E68
    x"38",x"D4",x"19",x"10",x"FA",x"21",x"BF",x"1E", -- 0x1E70
    x"11",x"C7",x"1E",x"06",x"08",x"3A",x"01",x"42", -- 0x1E78
    x"BE",x"28",x"07",x"23",x"13",x"13",x"13",x"13", -- 0x1E80
    x"10",x"F6",x"EB",x"3A",x"00",x"42",x"86",x"FD", -- 0x1E88
    x"77",x"01",x"23",x"3A",x"03",x"42",x"47",x"3E", -- 0x1E90
    x"F0",x"90",x"86",x"FD",x"77",x"03",x"23",x"7E", -- 0x1E98
    x"DD",x"77",x"02",x"23",x"7E",x"DD",x"77",x"01", -- 0x1EA0
    x"21",x"E7",x"1E",x"3A",x"1E",x"40",x"E6",x"03", -- 0x1EA8
    x"20",x"01",x"23",x"7E",x"DD",x"77",x"00",x"21", -- 0x1EB0
    x"D9",x"40",x"CB",x"CE",x"D1",x"C1",x"C9",x"50", -- 0x1EB8
    x"10",x"11",x"91",x"52",x"D2",x"12",x"92",x"09", -- 0x1EC0
    x"FD",x"00",x"FC",x"09",x"08",x"00",x"04",x"10", -- 0x1EC8
    x"02",x"04",x"00",x"00",x"02",x"FC",x"00",x"0F", -- 0x1ED0
    x"FA",x"04",x"FC",x"00",x"FA",x"FC",x"FC",x"0F", -- 0x1ED8
    x"09",x"04",x"04",x"00",x"09",x"FC",x"04",x"20", -- 0x1EE0
    x"0B",x"FD",x"21",x"20",x"42",x"06",x"04",x"11", -- 0x1EE8
    x"08",x"00",x"FD",x"7E",x"01",x"FD",x"E5",x"C5", -- 0x1EF0
    x"05",x"28",x"0A",x"FD",x"19",x"FD",x"BE",x"01", -- 0x1EF8
    x"CC",x"0D",x"1F",x"18",x"F3",x"C1",x"FD",x"E1", -- 0x1F00
    x"FD",x"19",x"10",x"E6",x"C9",x"FD",x"34",x"01", -- 0x1F08
    x"C9",x"3A",x"17",x"40",x"A7",x"C8",x"3E",x"13", -- 0x1F10
    x"21",x"1F",x"1F",x"CD",x"5C",x"09",x"C9",x"DD", -- 0x1F18
    x"CB",x"08",x"66",x"C4",x"41",x"1F",x"FD",x"7E", -- 0x1F20
    x"03",x"FE",x"10",x"DA",x"4F",x"0B",x"FE",x"F0", -- 0x1F28
    x"D2",x"4F",x"0B",x"FD",x"7E",x"00",x"FE",x"10", -- 0x1F30
    x"DA",x"4F",x"0B",x"FE",x"F0",x"D8",x"C3",x"4F", -- 0x1F38
    x"0B",x"DD",x"7E",x"0E",x"A7",x"F0",x"DD",x"36", -- 0x1F40
    x"0E",x"02",x"CD",x"E7",x"08",x"CB",x"28",x"CB", -- 0x1F48
    x"29",x"DD",x"70",x"03",x"DD",x"71",x"04",x"C9", -- 0x1F50
    x"CD",x"5F",x"1F",x"CD",x"2D",x"20",x"C9",x"DD", -- 0x1F58
    x"7E",x"FA",x"A7",x"C8",x"DD",x"7E",x"E2",x"DD", -- 0x1F60
    x"BE",x"F9",x"D0",x"21",x"72",x"1F",x"CD",x"3F", -- 0x1F68
    x"09",x"C9",x"FD",x"36",x"01",x"15",x"FD",x"36", -- 0x1F70
    x"02",x"06",x"CD",x"67",x"0B",x"FE",x"10",x"30", -- 0x1F78
    x"02",x"CB",x"E7",x"FE",x"F0",x"38",x"02",x"D6", -- 0x1F80
    x"10",x"57",x"26",x"10",x"CD",x"67",x"0B",x"CB", -- 0x1F88
    x"57",x"20",x"02",x"26",x"F0",x"CB",x"4F",x"20", -- 0x1F90
    x"01",x"EB",x"FD",x"72",x"00",x"FD",x"74",x"03", -- 0x1F98
    x"DD",x"E5",x"D1",x"13",x"21",x"75",x"20",x"01", -- 0x1FA0
    x"08",x"00",x"ED",x"B0",x"CD",x"E7",x"08",x"78", -- 0x1FA8
    x"A7",x"20",x"02",x"06",x"01",x"79",x"A7",x"20", -- 0x1FB0
    x"02",x"0E",x"01",x"DD",x"70",x"03",x"DD",x"71", -- 0x1FB8
    x"04",x"21",x"31",x"40",x"35",x"DD",x"CB",x"00", -- 0x1FC0
    x"CE",x"DD",x"CB",x"00",x"D6",x"21",x"DC",x"1F", -- 0x1FC8
    x"FD",x"E5",x"DD",x"E5",x"CD",x"3F",x"09",x"DD", -- 0x1FD0
    x"E1",x"FD",x"E1",x"C9",x"E1",x"DD",x"E5",x"D1", -- 0x1FD8
    x"FD",x"E5",x"E1",x"DD",x"E1",x"FD",x"E1",x"CD", -- 0x1FE0
    x"F8",x"1F",x"DD",x"7E",x"03",x"77",x"23",x"DD", -- 0x1FE8
    x"7E",x"04",x"77",x"DD",x"CB",x"08",x"DE",x"C9", -- 0x1FF0
    x"D5",x"E5",x"DD",x"72",x"0C",x"DD",x"73",x"0B", -- 0x1FF8
    x"DD",x"74",x"0A",x"DD",x"75",x"09",x"21",x"81", -- 0x2000
    x"29",x"13",x"01",x"08",x"00",x"ED",x"B0",x"E1", -- 0x2008
    x"D1",x"FD",x"7E",x"00",x"C6",x"02",x"77",x"23", -- 0x2010
    x"36",x"13",x"23",x"36",x"01",x"23",x"FD",x"7E", -- 0x2018
    x"03",x"C6",x"08",x"77",x"EB",x"CB",x"CE",x"CB", -- 0x2020
    x"D6",x"23",x"23",x"23",x"C9",x"DD",x"21",x"37", -- 0x2028
    x"40",x"DD",x"7E",x"E2",x"A7",x"C8",x"3E",x"15", -- 0x2030
    x"21",x"3F",x"20",x"CD",x"5C",x"09",x"C9",x"DD", -- 0x2038
    x"CB",x"08",x"5E",x"C8",x"DD",x"66",x"0C",x"DD", -- 0x2040
    x"6E",x"0B",x"CB",x"46",x"C8",x"21",x"5C",x"20", -- 0x2048
    x"FD",x"E5",x"DD",x"E5",x"CD",x"3F",x"09",x"DD", -- 0x2050
    x"E1",x"FD",x"E1",x"C9",x"E1",x"DD",x"E5",x"D1", -- 0x2058
    x"FD",x"E5",x"E1",x"DD",x"E1",x"FD",x"E1",x"CD", -- 0x2060
    x"F8",x"1F",x"CD",x"E7",x"08",x"70",x"23",x"71", -- 0x2068
    x"DD",x"CB",x"08",x"DE",x"C9",x"9B",x"1D",x"00", -- 0x2070
    x"00",x"00",x"00",x"00",x"00",x"DD",x"21",x"37", -- 0x2078
    x"40",x"DD",x"7E",x"E2",x"A7",x"C8",x"3E",x"15", -- 0x2080
    x"21",x"E4",x"20",x"CD",x"5C",x"09",x"DD",x"21", -- 0x2088
    x"37",x"40",x"DD",x"7E",x"E0",x"A7",x"C8",x"DD", -- 0x2090
    x"21",x"37",x"40",x"FD",x"21",x"04",x"42",x"06", -- 0x2098
    x"07",x"DD",x"CB",x"00",x"46",x"DD",x"E5",x"FD", -- 0x20A0
    x"E5",x"C5",x"C4",x"B8",x"20",x"C1",x"FD",x"E1", -- 0x20A8
    x"DD",x"E1",x"CD",x"78",x"09",x"10",x"EA",x"C9", -- 0x20B0
    x"DD",x"CB",x"08",x"5E",x"C8",x"DD",x"66",x"0C", -- 0x20B8
    x"DD",x"6E",x"0B",x"CB",x"46",x"C0",x"CB",x"4E", -- 0x20C0
    x"C8",x"DD",x"56",x"0A",x"DD",x"5E",x"09",x"13", -- 0x20C8
    x"1A",x"FE",x"13",x"C0",x"E5",x"D5",x"FD",x"E1", -- 0x20D0
    x"DD",x"E1",x"CD",x"E7",x"08",x"DD",x"70",x"03", -- 0x20D8
    x"DD",x"71",x"04",x"C9",x"FD",x"7E",x"00",x"FE", -- 0x20E0
    x"10",x"DA",x"4F",x"0B",x"FE",x"F0",x"D2",x"4F", -- 0x20E8
    x"0B",x"FD",x"7E",x"03",x"FE",x"10",x"DA",x"4F", -- 0x20F0
    x"0B",x"FE",x"F0",x"D2",x"4F",x"0B",x"DD",x"CB", -- 0x20F8
    x"00",x"46",x"C0",x"DD",x"7E",x"0E",x"E6",x"18", -- 0x2100
    x"20",x"05",x"FD",x"36",x"02",x"07",x"C9",x"FD", -- 0x2108
    x"36",x"02",x"06",x"C9",x"DD",x"21",x"C0",x"41", -- 0x2110
    x"DD",x"36",x"1B",x"06",x"DD",x"36",x"1A",x"04", -- 0x2118
    x"DD",x"36",x"1F",x"06",x"DD",x"36",x"1E",x"00", -- 0x2120
    x"DD",x"36",x"31",x"02",x"DD",x"36",x"30",x"00", -- 0x2128
    x"DD",x"36",x"35",x"02",x"DD",x"36",x"34",x"04", -- 0x2130
    x"21",x"20",x"22",x"FD",x"21",x"4D",x"53",x"06", -- 0x2138
    x"15",x"CD",x"3F",x"12",x"21",x"35",x"22",x"FD", -- 0x2140
    x"21",x"38",x"52",x"06",x"04",x"CD",x"3F",x"12", -- 0x2148
    x"11",x"00",x"03",x"3A",x"B0",x"40",x"A7",x"20", -- 0x2150
    x"29",x"D5",x"21",x"39",x"22",x"3A",x"B1",x"40", -- 0x2158
    x"DD",x"36",x"1E",x"04",x"3D",x"28",x"07",x"DD", -- 0x2160
    x"36",x"1E",x"00",x"21",x"47",x"22",x"FD",x"21", -- 0x2168
    x"CF",x"52",x"06",x"0E",x"CD",x"3F",x"12",x"D1", -- 0x2170
    x"CD",x"F5",x"21",x"C2",x"53",x"21",x"CD",x"17", -- 0x2178
    x"13",x"C9",x"D5",x"DD",x"36",x"1E",x"04",x"21", -- 0x2180
    x"55",x"22",x"FD",x"21",x"0F",x"53",x"06",x"11", -- 0x2188
    x"CD",x"3F",x"12",x"D1",x"AF",x"3D",x"08",x"CD", -- 0x2190
    x"48",x"13",x"CB",x"6F",x"08",x"20",x"03",x"08", -- 0x2198
    x"20",x"0A",x"CD",x"F5",x"21",x"C2",x"97",x"21", -- 0x21A0
    x"CD",x"17",x"13",x"C9",x"3A",x"B0",x"40",x"D6", -- 0x21A8
    x"01",x"27",x"32",x"B0",x"40",x"CD",x"9E",x"12", -- 0x21B0
    x"3A",x"00",x"68",x"06",x"03",x"CB",x"7F",x"28", -- 0x21B8
    x"02",x"06",x"05",x"78",x"32",x"1D",x"40",x"CD", -- 0x21C0
    x"17",x"13",x"3A",x"AF",x"40",x"CB",x"6F",x"28", -- 0x21C8
    x"12",x"21",x"A9",x"40",x"AF",x"77",x"23",x"77", -- 0x21D0
    x"23",x"77",x"CD",x"4E",x"12",x"21",x"BE",x"40", -- 0x21D8
    x"CB",x"C6",x"C9",x"21",x"AC",x"40",x"AF",x"77", -- 0x21E0
    x"23",x"77",x"23",x"77",x"CD",x"57",x"12",x"21", -- 0x21E8
    x"BE",x"40",x"CB",x"CE",x"C9",x"3E",x"05",x"CD", -- 0x21F0
    x"38",x"13",x"FD",x"21",x"3A",x"52",x"7B",x"D6", -- 0x21F8
    x"01",x"27",x"5F",x"7A",x"DE",x"00",x"27",x"57", -- 0x2200
    x"FD",x"77",x"00",x"7B",x"E6",x"0F",x"FD",x"77", -- 0x2208
    x"C0",x"7B",x"CB",x"3F",x"CB",x"3F",x"CB",x"3F", -- 0x2210
    x"CB",x"3F",x"FD",x"77",x"E0",x"7B",x"B2",x"C9", -- 0x2218
    x"54",x"4F",x"40",x"43",x"4F",x"4E",x"54",x"49", -- 0x2220
    x"4E",x"55",x"45",x"40",x"59",x"4F",x"55",x"52", -- 0x2228
    x"40",x"47",x"41",x"4D",x"45",x"54",x"49",x"4D", -- 0x2230
    x"45",x"49",x"4E",x"53",x"45",x"52",x"54",x"40", -- 0x2238
    x"41",x"40",x"43",x"4F",x"49",x"4E",x"40",x"49", -- 0x2240
    x"4E",x"53",x"45",x"52",x"54",x"40",x"32",x"40", -- 0x2248
    x"43",x"4F",x"49",x"4E",x"53",x"50",x"52",x"45", -- 0x2250
    x"53",x"53",x"40",x"46",x"49",x"52",x"45",x"40", -- 0x2258
    x"42",x"55",x"54",x"54",x"4F",x"4E",x"3A",x"EE", -- 0x2260
    x"40",x"A7",x"C2",x"72",x"23",x"21",x"D9",x"40", -- 0x2268
    x"46",x"CB",x"18",x"DC",x"EC",x"22",x"CB",x"18", -- 0x2270
    x"DC",x"FA",x"22",x"CB",x"18",x"DC",x"08",x"23", -- 0x2278
    x"CB",x"18",x"DC",x"21",x"23",x"CB",x"18",x"DC", -- 0x2280
    x"3A",x"23",x"CB",x"18",x"DC",x"53",x"23",x"3E", -- 0x2288
    x"FF",x"32",x"E2",x"40",x"3A",x"EF",x"40",x"CB", -- 0x2290
    x"67",x"C4",x"8F",x"24",x"E6",x"EF",x"C2",x"4F", -- 0x2298
    x"24",x"3A",x"EF",x"40",x"CB",x"7F",x"C4",x"E2", -- 0x22A0
    x"24",x"21",x"DA",x"40",x"46",x"CB",x"18",x"DC", -- 0x22A8
    x"98",x"23",x"CB",x"18",x"DC",x"A6",x"23",x"CB", -- 0x22B0
    x"18",x"DC",x"B1",x"23",x"CB",x"18",x"DC",x"C9", -- 0x22B8
    x"23",x"CB",x"18",x"DC",x"21",x"24",x"CB",x"18", -- 0x22C0
    x"DC",x"37",x"24",x"3A",x"E2",x"40",x"32",x"00", -- 0x22C8
    x"78",x"3A",x"E3",x"40",x"21",x"06",x"68",x"77", -- 0x22D0
    x"0F",x"77",x"3A",x"AF",x"40",x"CB",x"57",x"C0", -- 0x22D8
    x"21",x"03",x"68",x"3A",x"DA",x"40",x"77",x"0F", -- 0x22E0
    x"23",x"23",x"77",x"C9",x"21",x"D9",x"40",x"CB", -- 0x22E8
    x"86",x"23",x"CB",x"C6",x"3E",x"30",x"32",x"DB", -- 0x22F0
    x"40",x"C9",x"21",x"D9",x"40",x"CB",x"8E",x"23", -- 0x22F8
    x"CB",x"CE",x"3E",x"04",x"32",x"DC",x"40",x"C9", -- 0x2300
    x"21",x"D9",x"40",x"CB",x"96",x"23",x"CB",x"D6", -- 0x2308
    x"21",x"1C",x"23",x"11",x"DD",x"40",x"01",x"06", -- 0x2310
    x"00",x"ED",x"B0",x"C9",x"B9",x"23",x"08",x"01", -- 0x2318
    x"02",x"21",x"D9",x"40",x"CB",x"9E",x"23",x"CB", -- 0x2320
    x"DE",x"21",x"35",x"23",x"11",x"E4",x"40",x"01", -- 0x2328
    x"06",x"00",x"ED",x"B0",x"C9",x"D1",x"23",x"28", -- 0x2330
    x"01",x"02",x"21",x"D9",x"40",x"CB",x"A6",x"23", -- 0x2338
    x"CB",x"E6",x"21",x"4E",x"23",x"11",x"E9",x"40", -- 0x2340
    x"01",x"06",x"00",x"ED",x"B0",x"C9",x"29",x"24", -- 0x2348
    x"07",x"01",x"01",x"3A",x"AF",x"40",x"CB",x"57", -- 0x2350
    x"C0",x"21",x"D9",x"40",x"CB",x"AE",x"23",x"CB", -- 0x2358
    x"EE",x"21",x"6D",x"23",x"11",x"E4",x"40",x"01", -- 0x2360
    x"06",x"00",x"ED",x"B0",x"C9",x"3F",x"24",x"08", -- 0x2368
    x"01",x"03",x"21",x"EE",x"40",x"CB",x"56",x"20", -- 0x2370
    x"12",x"CB",x"5E",x"CA",x"6D",x"22",x"CB",x"9E", -- 0x2378
    x"23",x"CB",x"DE",x"21",x"F3",x"40",x"36",x"E0", -- 0x2380
    x"C3",x"6D",x"22",x"CB",x"96",x"23",x"CB",x"D6", -- 0x2388
    x"21",x"F2",x"40",x"36",x"00",x"C3",x"6D",x"22", -- 0x2390
    x"21",x"DB",x"40",x"35",x"C0",x"21",x"DA",x"40", -- 0x2398
    x"CB",x"86",x"2B",x"CB",x"EE",x"C9",x"21",x"DC", -- 0x23A0
    x"40",x"35",x"C0",x"21",x"DA",x"40",x"CB",x"8E", -- 0x23A8
    x"C9",x"FD",x"21",x"DD",x"40",x"0E",x"04",x"CD", -- 0x23B0
    x"AD",x"24",x"C9",x"4B",x"06",x"FF",x"03",x"4B", -- 0x23B8
    x"06",x"FF",x"03",x"4B",x"06",x"FF",x"03",x"1C", -- 0x23C0
    x"0C",x"FD",x"21",x"E4",x"40",x"0E",x"08",x"CD", -- 0x23C8
    x"AD",x"24",x"C9",x"68",x"05",x"FF",x"02",x"68", -- 0x23D0
    x"05",x"FF",x"02",x"68",x"05",x"FF",x"02",x"68", -- 0x23D8
    x"13",x"FF",x"02",x"68",x"05",x"FF",x"02",x"68", -- 0x23E0
    x"05",x"FF",x"02",x"68",x"05",x"FF",x"02",x"68", -- 0x23E8
    x"08",x"FF",x"02",x"4B",x"08",x"FF",x"02",x"1C", -- 0x23F0
    x"08",x"FF",x"02",x"4B",x"08",x"FF",x"02",x"68", -- 0x23F8
    x"08",x"FF",x"02",x"4B",x"08",x"FF",x"02",x"1C", -- 0x2400
    x"08",x"FF",x"02",x"4B",x"08",x"FF",x"02",x"68", -- 0x2408
    x"13",x"FF",x"02",x"68",x"05",x"FF",x"02",x"68", -- 0x2410
    x"05",x"FF",x"02",x"68",x"05",x"FF",x"02",x"68", -- 0x2418
    x"13",x"FD",x"21",x"E9",x"40",x"0E",x"10",x"CD", -- 0x2420
    x"AD",x"24",x"C9",x"9A",x"05",x"FF",x"04",x"9A", -- 0x2428
    x"05",x"FF",x"04",x"8E",x"03",x"9A",x"0C",x"FD", -- 0x2430
    x"21",x"E4",x"40",x"0E",x"20",x"CD",x"AD",x"24", -- 0x2438
    x"C9",x"80",x"10",x"FF",x"06",x"70",x"08",x"68", -- 0x2440
    x"10",x"FF",x"06",x"55",x"08",x"40",x"18",x"3A", -- 0x2448
    x"EF",x"40",x"CB",x"5F",x"20",x"1F",x"CB",x"57", -- 0x2450
    x"CA",x"A1",x"22",x"21",x"F2",x"40",x"3E",x"10", -- 0x2458
    x"86",x"77",x"32",x"E2",x"40",x"3E",x"03",x"32", -- 0x2460
    x"E3",x"40",x"D2",x"A1",x"22",x"21",x"EF",x"40", -- 0x2468
    x"CB",x"96",x"C3",x"A1",x"22",x"21",x"F3",x"40", -- 0x2470
    x"7E",x"D6",x"10",x"77",x"32",x"E2",x"40",x"3E", -- 0x2478
    x"03",x"32",x"E3",x"40",x"D2",x"A1",x"22",x"21", -- 0x2480
    x"EF",x"40",x"CB",x"9E",x"C3",x"A1",x"22",x"F5", -- 0x2488
    x"21",x"F0",x"40",x"7E",x"32",x"E2",x"40",x"3E", -- 0x2490
    x"03",x"32",x"E3",x"40",x"F1",x"23",x"35",x"C0", -- 0x2498
    x"36",x"0A",x"2B",x"CB",x"56",x"28",x"03",x"36", -- 0x24A0
    x"B8",x"C9",x"36",x"B4",x"C9",x"FD",x"35",x"03", -- 0x24A8
    x"20",x"1F",x"FD",x"35",x"02",x"20",x"07",x"21", -- 0x24B0
    x"DA",x"40",x"7E",x"A9",x"77",x"C9",x"FD",x"6E", -- 0x24B8
    x"00",x"FD",x"66",x"01",x"23",x"23",x"FD",x"75", -- 0x24C0
    x"00",x"FD",x"74",x"01",x"23",x"7E",x"FD",x"77", -- 0x24C8
    x"03",x"FD",x"6E",x"00",x"FD",x"66",x"01",x"7E", -- 0x24D0
    x"32",x"E2",x"40",x"FD",x"7E",x"04",x"32",x"E3", -- 0x24D8
    x"40",x"C9",x"3A",x"28",x"40",x"E6",x"0F",x"C6", -- 0x24E0
    x"80",x"32",x"E2",x"40",x"3E",x"03",x"32",x"E3", -- 0x24E8
    x"40",x"C9",x"3A",x"17",x"40",x"A7",x"20",x"08", -- 0x24F0
    x"21",x"EF",x"40",x"CB",x"A6",x"C3",x"21",x"25", -- 0x24F8
    x"3A",x"01",x"40",x"CB",x"47",x"20",x"F1",x"21", -- 0x2500
    x"EF",x"40",x"CB",x"66",x"20",x"13",x"3A",x"1E", -- 0x2508
    x"40",x"E6",x"03",x"FE",x"02",x"20",x"0A",x"CB", -- 0x2510
    x"E6",x"21",x"F0",x"40",x"36",x"B8",x"23",x"36", -- 0x2518
    x"0A",x"3A",x"AF",x"40",x"CB",x"57",x"C0",x"3A", -- 0x2520
    x"16",x"40",x"A7",x"20",x"0A",x"AF",x"21",x"00", -- 0x2528
    x"68",x"77",x"23",x"77",x"23",x"77",x"C9",x"CB", -- 0x2530
    x"27",x"3C",x"ED",x"44",x"06",x"04",x"21",x"04", -- 0x2538
    x"60",x"77",x"23",x"0F",x"10",x"FB",x"3E",x"01", -- 0x2540
    x"C3",x"2E",x"25",x"3A",x"AF",x"40",x"CB",x"57", -- 0x2548
    x"C0",x"3E",x"01",x"06",x"04",x"21",x"00",x"68", -- 0x2550
    x"77",x"23",x"10",x"FC",x"3A",x"27",x"40",x"E6", -- 0x2558
    x"F0",x"0F",x"0F",x"0F",x"0F",x"47",x"3E",x"0F", -- 0x2560
    x"90",x"06",x"04",x"21",x"04",x"60",x"77",x"0F", -- 0x2568
    x"23",x"10",x"FB",x"C9",x"DD",x"7E",x"DF",x"A7", -- 0x2570
    x"28",x"05",x"DD",x"7E",x"FF",x"A7",x"C0",x"CD", -- 0x2578
    x"67",x"0B",x"E6",x"3F",x"DD",x"77",x"FF",x"DD", -- 0x2580
    x"7E",x"F7",x"A7",x"C8",x"DD",x"7E",x"E1",x"DD", -- 0x2588
    x"BE",x"F8",x"D0",x"21",x"9A",x"25",x"CD",x"3F", -- 0x2590
    x"09",x"C9",x"FD",x"36",x"00",x"10",x"FD",x"36", -- 0x2598
    x"01",x"14",x"06",x"03",x"3A",x"2E",x"40",x"FE", -- 0x25A0
    x"03",x"30",x"02",x"06",x"05",x"FD",x"70",x"02", -- 0x25A8
    x"CD",x"67",x"0B",x"FD",x"77",x"03",x"DD",x"E5", -- 0x25B0
    x"D1",x"13",x"21",x"EE",x"25",x"01",x"08",x"00", -- 0x25B8
    x"ED",x"B0",x"CD",x"67",x"0B",x"6F",x"26",x"00", -- 0x25C0
    x"3A",x"1F",x"40",x"4F",x"06",x"08",x"29",x"7C", -- 0x25C8
    x"91",x"38",x"02",x"67",x"2C",x"10",x"F7",x"7C", -- 0x25D0
    x"DD",x"77",x"07",x"3A",x"F4",x"40",x"DD",x"77", -- 0x25D8
    x"0E",x"21",x"2E",x"40",x"35",x"DD",x"CB",x"00", -- 0x25E0
    x"CE",x"DD",x"CB",x"00",x"D6",x"C9",x"59",x"1D", -- 0x25E8
    x"79",x"0B",x"01",x"2C",x"00",x"01",x"DD",x"21", -- 0x25F0
    x"37",x"40",x"DD",x"7E",x"E1",x"A7",x"C8",x"3E", -- 0x25F8
    x"14",x"21",x"08",x"26",x"CD",x"5C",x"09",x"C9", -- 0x2600
    x"DD",x"CB",x"08",x"46",x"28",x"3E",x"DD",x"CB", -- 0x2608
    x"00",x"7E",x"20",x"1A",x"DD",x"7E",x"06",x"A7", -- 0x2610
    x"C0",x"DD",x"36",x"06",x"43",x"11",x"79",x"0B", -- 0x2618
    x"DD",x"73",x"03",x"DD",x"72",x"04",x"DD",x"36", -- 0x2620
    x"05",x"01",x"DD",x"35",x"07",x"C0",x"DD",x"CB", -- 0x2628
    x"08",x"26",x"AF",x"32",x"01",x"70",x"DD",x"36", -- 0x2630
    x"01",x"9B",x"DD",x"36",x"02",x"1D",x"3C",x"32", -- 0x2638
    x"01",x"70",x"CD",x"E7",x"08",x"DD",x"70",x"03", -- 0x2640
    x"DD",x"71",x"04",x"C9",x"FD",x"7E",x"00",x"FE", -- 0x2648
    x"10",x"38",x"0E",x"FE",x"F0",x"30",x"0A",x"FD", -- 0x2650
    x"7E",x"03",x"FE",x"02",x"38",x"03",x"FE",x"F0", -- 0x2658
    x"D8",x"DD",x"CB",x"00",x"46",x"C0",x"DD",x"CB", -- 0x2660
    x"00",x"8E",x"DD",x"CB",x"00",x"96",x"AF",x"FD", -- 0x2668
    x"77",x"00",x"FD",x"77",x"01",x"FD",x"77",x"03", -- 0x2670
    x"CD",x"67",x"0B",x"32",x"36",x"40",x"C9",x"3A", -- 0x2678
    x"1E",x"40",x"E6",x"1F",x"CB",x"2F",x"CB",x"2F", -- 0x2680
    x"A7",x"28",x"01",x"3D",x"6F",x"26",x"00",x"29", -- 0x2688
    x"29",x"29",x"E5",x"29",x"D1",x"19",x"11",x"A3", -- 0x2690
    x"26",x"19",x"11",x"1F",x"40",x"01",x"18",x"00", -- 0x2698
    x"ED",x"B0",x"C9",x"0E",x"10",x"0A",x"09",x"07", -- 0x26A0
    x"15",x"07",x"1C",x"99",x"99",x"02",x"00",x"3B", -- 0x26A8
    x"00",x"02",x"1E",x"04",x"04",x"32",x"02",x"0E", -- 0x26B0
    x"28",x"00",x"10",x"0D",x"0A",x"09",x"06",x"07", -- 0x26B8
    x"13",x"08",x"18",x"99",x"99",x"02",x"00",x"3A", -- 0x26C0
    x"00",x"02",x"23",x"05",x"05",x"3C",x"02",x"10", -- 0x26C8
    x"1E",x"00",x"10",x"0C",x"09",x"08",x"05",x"06", -- 0x26D0
    x"0C",x"07",x"16",x"99",x"99",x"02",x"00",x"39", -- 0x26D8
    x"00",x"03",x"23",x"05",x"05",x"46",x"02",x"12", -- 0x26E0
    x"14",x"00",x"10",x"0B",x"09",x"08",x"05",x"06", -- 0x26E8
    x"0C",x"04",x"14",x"99",x"99",x"02",x"00",x"38", -- 0x26F0
    x"00",x"03",x"28",x"06",x"05",x"50",x"03",x"14", -- 0x26F8
    x"0A",x"00",x"10",x"0A",x"0A",x"04",x"07",x"07", -- 0x2700
    x"06",x"04",x"13",x"99",x"99",x"02",x"00",x"37", -- 0x2708
    x"00",x"03",x"32",x"07",x"06",x"5A",x"03",x"16", -- 0x2710
    x"08",x"00",x"10",x"09",x"08",x"05",x"07",x"04", -- 0x2718
    x"06",x"03",x"12",x"99",x"99",x"02",x"00",x"36", -- 0x2720
    x"00",x"03",x"32",x"07",x"07",x"64",x"04",x"19", -- 0x2728
    x"06",x"00",x"10",x"07",x"08",x"05",x"07",x"04", -- 0x2730
    x"06",x"03",x"11",x"99",x"99",x"03",x"00",x"1A", -- 0x2738
    x"00",x"03",x"32",x"07",x"07",x"78",x"04",x"19", -- 0x2740
    x"04",x"00",x"10",x"DD",x"21",x"37",x"40",x"DD", -- 0x2748
    x"E5",x"CD",x"EC",x"27",x"DD",x"E1",x"DD",x"7E", -- 0x2750
    x"FB",x"DD",x"BE",x"E5",x"C8",x"DD",x"7E",x"FC", -- 0x2758
    x"A7",x"C8",x"DD",x"7E",x"DF",x"A7",x"28",x"05", -- 0x2760
    x"DD",x"7E",x"FF",x"A7",x"C0",x"DD",x"7E",x"FD", -- 0x2768
    x"DD",x"77",x"FF",x"21",x"7A",x"27",x"CD",x"3F", -- 0x2770
    x"09",x"C9",x"DD",x"E5",x"D1",x"13",x"21",x"DD", -- 0x2778
    x"27",x"01",x"0F",x"00",x"ED",x"B0",x"CD",x"67", -- 0x2780
    x"0B",x"DD",x"77",x"0F",x"06",x"10",x"16",x"02", -- 0x2788
    x"CB",x"7F",x"28",x"04",x"06",x"F0",x"16",x"FE", -- 0x2790
    x"0E",x"10",x"1E",x"02",x"CB",x"77",x"28",x"04", -- 0x2798
    x"0E",x"F0",x"1E",x"FE",x"FD",x"70",x"00",x"FD", -- 0x27A0
    x"71",x"03",x"DD",x"72",x"03",x"DD",x"73",x"04", -- 0x27A8
    x"CD",x"67",x"0B",x"E6",x"3F",x"F6",x"07",x"DD", -- 0x27B0
    x"77",x"0E",x"FD",x"36",x"01",x"18",x"06",x"00", -- 0x27B8
    x"3A",x"33",x"40",x"FE",x"03",x"30",x"02",x"06", -- 0x27C0
    x"01",x"FD",x"70",x"02",x"DD",x"CB",x"00",x"CE", -- 0x27C8
    x"DD",x"CB",x"00",x"D6",x"21",x"33",x"40",x"35", -- 0x27D0
    x"DD",x"CB",x"08",x"DE",x"C9",x"9B",x"1D",x"00", -- 0x27D8
    x"00",x"01",x"11",x"00",x"01",x"00",x"00",x"00", -- 0x27E0
    x"00",x"00",x"04",x"00",x"3E",x"18",x"21",x"3D", -- 0x27E8
    x"28",x"CD",x"5C",x"09",x"DD",x"21",x"37",x"40", -- 0x27F0
    x"DD",x"7E",x"FF",x"A7",x"C0",x"DD",x"7E",x"E0", -- 0x27F8
    x"DD",x"BE",x"F6",x"D0",x"CD",x"67",x"0B",x"6F", -- 0x2800
    x"26",x"00",x"3A",x"1C",x"40",x"4F",x"06",x"08", -- 0x2808
    x"29",x"7C",x"91",x"38",x"02",x"67",x"2C",x"10", -- 0x2810
    x"F7",x"4C",x"0C",x"DD",x"21",x"37",x"40",x"FD", -- 0x2818
    x"21",x"04",x"42",x"06",x"07",x"FD",x"7E",x"01", -- 0x2820
    x"FE",x"18",x"20",x"03",x"0D",x"28",x"06",x"CD", -- 0x2828
    x"78",x"09",x"10",x"F1",x"C9",x"DD",x"CB",x"08", -- 0x2830
    x"66",x"C0",x"C3",x"4B",x"28",x"DD",x"CB",x"00", -- 0x2838
    x"46",x"C8",x"DD",x"CB",x"08",x"66",x"C0",x"DD", -- 0x2840
    x"CB",x"08",x"E6",x"FD",x"E5",x"21",x"56",x"28", -- 0x2848
    x"CD",x"3F",x"09",x"FD",x"E1",x"C9",x"D1",x"D1", -- 0x2850
    x"1A",x"47",x"3A",x"00",x"42",x"B8",x"38",x"04", -- 0x2858
    x"78",x"C6",x"E0",x"47",x"78",x"C6",x"10",x"FD", -- 0x2860
    x"77",x"00",x"FD",x"36",x"01",x"13",x"FD",x"36", -- 0x2868
    x"02",x"06",x"13",x"13",x"13",x"1A",x"FD",x"77", -- 0x2870
    x"03",x"DD",x"E5",x"D1",x"13",x"21",x"81",x"29", -- 0x2878
    x"01",x"08",x"00",x"ED",x"B0",x"DD",x"36",x"0E", -- 0x2880
    x"0A",x"DD",x"CB",x"08",x"E6",x"DD",x"CB",x"00", -- 0x2888
    x"CE",x"DD",x"CB",x"00",x"D6",x"C9",x"DD",x"21", -- 0x2890
    x"37",x"40",x"DD",x"7E",x"FB",x"A7",x"C8",x"3E", -- 0x2898
    x"18",x"21",x"A8",x"28",x"CD",x"5C",x"09",x"C9", -- 0x28A0
    x"DD",x"CB",x"08",x"5E",x"C2",x"E4",x"28",x"DD", -- 0x28A8
    x"CB",x"00",x"7E",x"C2",x"5F",x"29",x"CD",x"2F", -- 0x28B0
    x"29",x"FD",x"7E",x"00",x"FE",x"20",x"47",x"30", -- 0x28B8
    x"04",x"FD",x"36",x"00",x"20",x"78",x"FE",x"E0", -- 0x28C0
    x"38",x"04",x"FD",x"36",x"00",x"DF",x"FD",x"7E", -- 0x28C8
    x"03",x"FE",x"20",x"47",x"30",x"04",x"FD",x"36", -- 0x28D0
    x"03",x"20",x"78",x"FE",x"E0",x"38",x"04",x"FD", -- 0x28D8
    x"36",x"03",x"DF",x"C9",x"FD",x"7E",x"00",x"FE", -- 0x28E0
    x"08",x"DA",x"4F",x"0B",x"FE",x"F8",x"D2",x"4F", -- 0x28E8
    x"0B",x"FD",x"7E",x"03",x"FE",x"08",x"DA",x"4F", -- 0x28F0
    x"0B",x"FE",x"F8",x"D2",x"4F",x"0B",x"DD",x"7E", -- 0x28F8
    x"0E",x"A7",x"C0",x"DD",x"CB",x"08",x"9E",x"CD", -- 0x2900
    x"67",x"0B",x"F6",x"0F",x"DD",x"77",x"0E",x"21", -- 0x2908
    x"2B",x"29",x"DD",x"E5",x"D1",x"13",x"3E",x"00", -- 0x2910
    x"32",x"01",x"70",x"01",x"04",x"00",x"ED",x"B0", -- 0x2918
    x"3C",x"32",x"01",x"70",x"CD",x"67",x"0B",x"DD", -- 0x2920
    x"77",x"07",x"C9",x"A2",x"1D",x"C1",x"0B",x"DD", -- 0x2928
    x"7E",x"06",x"A7",x"C0",x"DD",x"36",x"06",x"11", -- 0x2930
    x"11",x"C1",x"0B",x"DD",x"73",x"03",x"DD",x"72", -- 0x2938
    x"04",x"DD",x"36",x"05",x"01",x"DD",x"46",x"0F", -- 0x2940
    x"CB",x"60",x"28",x"04",x"3E",x"02",x"A8",x"47", -- 0x2948
    x"CB",x"68",x"28",x"04",x"3E",x"08",x"A8",x"47", -- 0x2950
    x"DD",x"70",x"0F",x"DD",x"35",x"07",x"C0",x"DD", -- 0x2958
    x"E5",x"D1",x"13",x"21",x"DD",x"27",x"01",x"04", -- 0x2960
    x"00",x"AF",x"32",x"01",x"70",x"ED",x"B0",x"3C", -- 0x2968
    x"32",x"01",x"70",x"CD",x"E7",x"08",x"DD",x"70", -- 0x2970
    x"03",x"DD",x"71",x"04",x"DD",x"CB",x"08",x"DE", -- 0x2978
    x"C9",x"9B",x"1D",x"00",x"00",x"00",x"00",x"00", -- 0x2980
    x"00",x"7F",x"7E",x"7F",x"7E",x"7F",x"7E",x"7F", -- 0x2988
    x"7E",x"7F",x"7E",x"7F",x"7E",x"7F",x"7E",x"7F", -- 0x2990
    x"7E",x"7F",x"7E",x"7F",x"7E",x"7F",x"7E",x"7F", -- 0x2998
    x"7E",x"5F",x"5E",x"5F",x"5E",x"5F",x"5E",x"5F", -- 0x29A0
    x"5E",x"5F",x"5E",x"5F",x"5E",x"5F",x"5E",x"5F", -- 0x29A8
    x"5E",x"5F",x"5E",x"5F",x"5E",x"5F",x"5E",x"5F", -- 0x29B0
    x"5E",x"5F",x"5E",x"5F",x"5E",x"5F",x"5E",x"5F", -- 0x29B8
    x"5E",x"3F",x"3E",x"3F",x"3E",x"3F",x"3E",x"3F", -- 0x29C0
    x"3E",x"3F",x"3E",x"3F",x"3E",x"3F",x"3E",x"3F", -- 0x29C8
    x"3E",x"3F",x"3E",x"3F",x"3E",x"3F",x"3E",x"3F", -- 0x29D0
    x"3E",x"3F",x"3E",x"3F",x"3E",x"3F",x"3E",x"3F", -- 0x29D8
    x"3E",x"1F",x"1E",x"1F",x"1E",x"1F",x"1E",x"1F", -- 0x29E0
    x"1E",x"1F",x"1E",x"1F",x"1E",x"1F",x"1E",x"1F", -- 0x29E8
    x"1E",x"1F",x"1E",x"1F",x"1E",x"1F",x"1E",x"1F", -- 0x29F0
    x"1E",x"1F",x"1E",x"1F",x"1E",x"1F",x"1E",x"1F", -- 0x29F8
    x"1E",x"FF",x"FF",x"FD",x"FD",x"FF",x"FF",x"FD", -- 0x2A00
    x"FD",x"FF",x"FF",x"FD",x"FD",x"FF",x"FF",x"FD", -- 0x2A08
    x"FD",x"FF",x"FF",x"FD",x"FD",x"FF",x"FF",x"FD", -- 0x2A10
    x"FD",x"FF",x"FF",x"FD",x"FD",x"FF",x"FF",x"FD", -- 0x2A18
    x"FD",x"DF",x"DF",x"DD",x"DD",x"DF",x"DF",x"DD", -- 0x2A20
    x"DD",x"DF",x"DF",x"DD",x"DD",x"DF",x"DF",x"DD", -- 0x2A28
    x"DD",x"DF",x"DF",x"DD",x"DD",x"DF",x"DF",x"DD", -- 0x2A30
    x"DD",x"DF",x"DF",x"DD",x"DD",x"DF",x"DF",x"DD", -- 0x2A38
    x"DD",x"BF",x"BF",x"BD",x"BD",x"BF",x"BF",x"BD", -- 0x2A40
    x"BD",x"BF",x"BF",x"BD",x"BD",x"BF",x"BF",x"BD", -- 0x2A48
    x"BD",x"BF",x"BF",x"BD",x"BD",x"BF",x"BF",x"BD", -- 0x2A50
    x"BD",x"BF",x"BF",x"BD",x"BD",x"BF",x"BF",x"BD", -- 0x2A58
    x"BD",x"9F",x"9F",x"9D",x"9D",x"9F",x"9F",x"9D", -- 0x2A60
    x"9D",x"9F",x"9F",x"9D",x"9D",x"9F",x"9F",x"9D", -- 0x2A68
    x"9D",x"9F",x"9F",x"9D",x"9D",x"9F",x"9F",x"9D", -- 0x2A70
    x"9D",x"9F",x"9F",x"9D",x"9D",x"9F",x"9F",x"9D", -- 0x2A78
    x"9D",x"7F",x"7F",x"7D",x"7D",x"7F",x"7F",x"7D", -- 0x2A80
    x"7D",x"7F",x"7F",x"7D",x"7D",x"7F",x"7F",x"7D", -- 0x2A88
    x"7D",x"7F",x"7F",x"7D",x"7D",x"7F",x"7F",x"7D", -- 0x2A90
    x"7D",x"7F",x"7F",x"7D",x"7D",x"7F",x"7F",x"7D", -- 0x2A98
    x"7D",x"5F",x"5F",x"5D",x"5D",x"5F",x"5F",x"5D", -- 0x2AA0
    x"5D",x"5F",x"5F",x"5D",x"5D",x"5F",x"5F",x"5D", -- 0x2AA8
    x"5D",x"5F",x"5F",x"5D",x"5D",x"5F",x"5F",x"5D", -- 0x2AB0
    x"5D",x"5F",x"5F",x"5D",x"5D",x"5F",x"5F",x"5D", -- 0x2AB8
    x"5D",x"3F",x"3F",x"3D",x"3D",x"3F",x"3F",x"3D", -- 0x2AC0
    x"3D",x"3F",x"3F",x"3D",x"3D",x"3F",x"3F",x"3D", -- 0x2AC8
    x"3D",x"3F",x"3F",x"3D",x"3D",x"3F",x"3F",x"3D", -- 0x2AD0
    x"3D",x"3F",x"3F",x"3D",x"3D",x"3F",x"3F",x"3D", -- 0x2AD8
    x"3D",x"1F",x"1F",x"1D",x"1D",x"1F",x"1F",x"1D", -- 0x2AE0
    x"1D",x"1F",x"1F",x"1D",x"1D",x"1F",x"1F",x"1D", -- 0x2AE8
    x"1D",x"1F",x"1F",x"1D",x"1D",x"1F",x"1F",x"1D", -- 0x2AF0
    x"1D",x"1F",x"1F",x"1D",x"1D",x"1F",x"1F",x"1D", -- 0x2AF8
    x"1D",x"FF",x"FE",x"FD",x"FC",x"FF",x"FE",x"FD", -- 0x2B00
    x"FC",x"FF",x"FE",x"FD",x"FC",x"FF",x"FE",x"FD", -- 0x2B08
    x"FC",x"FF",x"FE",x"FD",x"FC",x"FF",x"FE",x"FD", -- 0x2B10
    x"FC",x"FF",x"FE",x"FD",x"FC",x"FF",x"FE",x"FD", -- 0x2B18
    x"FC",x"DF",x"DE",x"DD",x"DC",x"DF",x"DE",x"DD", -- 0x2B20
    x"DC",x"DF",x"DE",x"DD",x"DC",x"DF",x"DE",x"DD", -- 0x2B28
    x"DC",x"DF",x"DE",x"DD",x"DC",x"DF",x"DE",x"DD", -- 0x2B30
    x"DC",x"DF",x"DE",x"DD",x"DC",x"DF",x"DE",x"DD", -- 0x2B38
    x"DC",x"BF",x"BE",x"BD",x"BC",x"BF",x"BE",x"BD", -- 0x2B40
    x"BC",x"BF",x"BE",x"BD",x"BC",x"BF",x"BE",x"BD", -- 0x2B48
    x"BC",x"BF",x"BE",x"BD",x"BC",x"BF",x"BE",x"BD", -- 0x2B50
    x"BC",x"BF",x"BE",x"BD",x"BC",x"BF",x"BE",x"BD", -- 0x2B58
    x"BC",x"9F",x"9E",x"9D",x"9C",x"9F",x"9E",x"9D", -- 0x2B60
    x"9C",x"9F",x"9E",x"9D",x"9C",x"9F",x"9E",x"9D", -- 0x2B68
    x"9C",x"9F",x"9E",x"9D",x"9C",x"9F",x"9E",x"9D", -- 0x2B70
    x"9C",x"9F",x"9E",x"9D",x"9C",x"9F",x"9E",x"9D", -- 0x2B78
    x"9C",x"7F",x"7E",x"7D",x"7C",x"7F",x"7E",x"7D", -- 0x2B80
    x"7C",x"7F",x"7E",x"7D",x"7C",x"7F",x"7E",x"7D", -- 0x2B88
    x"7C",x"7F",x"7E",x"7D",x"7C",x"7F",x"7E",x"7D", -- 0x2B90
    x"7C",x"7F",x"7E",x"7D",x"7C",x"7F",x"7E",x"7D", -- 0x2B98
    x"7C",x"5F",x"5E",x"5D",x"5C",x"5F",x"5E",x"5D", -- 0x2BA0
    x"5C",x"5F",x"5E",x"5D",x"5C",x"5F",x"5E",x"5D", -- 0x2BA8
    x"5C",x"5F",x"5E",x"5D",x"5C",x"5F",x"5E",x"5D", -- 0x2BB0
    x"5C",x"5F",x"5E",x"5D",x"5C",x"5F",x"5E",x"5D", -- 0x2BB8
    x"5C",x"3F",x"3E",x"3D",x"3C",x"3F",x"3E",x"3D", -- 0x2BC0
    x"3C",x"3F",x"3E",x"3D",x"3C",x"3F",x"3E",x"3D", -- 0x2BC8
    x"3C",x"3F",x"3E",x"3D",x"3C",x"3F",x"3E",x"3D", -- 0x2BD0
    x"3C",x"3F",x"3E",x"3D",x"3C",x"3F",x"3E",x"3D", -- 0x2BD8
    x"3C",x"1F",x"1E",x"1D",x"1C",x"1F",x"1E",x"1D", -- 0x2BE0
    x"1C",x"1F",x"1E",x"1D",x"1C",x"1F",x"1E",x"1D", -- 0x2BE8
    x"1C",x"1F",x"1E",x"1D",x"1C",x"1F",x"1E",x"1D", -- 0x2BF0
    x"1C",x"1F",x"1E",x"1D",x"1C",x"1F",x"1E",x"1D", -- 0x2BF8
    x"1C",x"FF",x"FF",x"FF",x"FF",x"FB",x"FB",x"FB", -- 0x2C00
    x"FB",x"FF",x"FF",x"FF",x"FF",x"FB",x"FB",x"FB", -- 0x2C08
    x"FB",x"FF",x"FF",x"FF",x"FF",x"FB",x"FB",x"FB", -- 0x2C10
    x"FB",x"FF",x"FF",x"FF",x"FF",x"FB",x"FB",x"FB", -- 0x2C18
    x"FB",x"DF",x"DF",x"DF",x"DF",x"DB",x"DB",x"DB", -- 0x2C20
    x"DB",x"DF",x"DF",x"DF",x"DF",x"DB",x"DB",x"DB", -- 0x2C28
    x"DB",x"DF",x"DF",x"DF",x"DF",x"DB",x"DB",x"DB", -- 0x2C30
    x"DB",x"DF",x"DF",x"DF",x"DF",x"DB",x"DB",x"DB", -- 0x2C38
    x"DB",x"BF",x"BF",x"BF",x"BF",x"BB",x"BB",x"BB", -- 0x2C40
    x"BB",x"BF",x"BF",x"BF",x"BF",x"BB",x"BB",x"BB", -- 0x2C48
    x"BB",x"BF",x"BF",x"BF",x"BF",x"BB",x"BB",x"BB", -- 0x2C50
    x"BB",x"BF",x"BF",x"BF",x"BF",x"BB",x"BB",x"BB", -- 0x2C58
    x"BB",x"9F",x"9F",x"9F",x"9F",x"9B",x"9B",x"9B", -- 0x2C60
    x"9B",x"9F",x"9F",x"9F",x"9F",x"9B",x"9B",x"9B", -- 0x2C68
    x"9B",x"9F",x"9F",x"9F",x"9F",x"9B",x"9B",x"9B", -- 0x2C70
    x"9B",x"9F",x"9F",x"9F",x"9F",x"9B",x"9B",x"9B", -- 0x2C78
    x"9B",x"7F",x"7F",x"7F",x"7F",x"7B",x"7B",x"7B", -- 0x2C80
    x"7B",x"7F",x"7F",x"7F",x"7F",x"7B",x"7B",x"7B", -- 0x2C88
    x"7B",x"7F",x"7F",x"7F",x"7F",x"7B",x"7B",x"7B", -- 0x2C90
    x"7B",x"7F",x"7F",x"7F",x"7F",x"7B",x"7B",x"7B", -- 0x2C98
    x"7B",x"5F",x"5F",x"5F",x"5F",x"5B",x"5B",x"5B", -- 0x2CA0
    x"5B",x"5F",x"5F",x"5F",x"5F",x"5B",x"5B",x"5B", -- 0x2CA8
    x"5B",x"5F",x"5F",x"5F",x"5F",x"5B",x"5B",x"5B", -- 0x2CB0
    x"5B",x"5F",x"5F",x"5F",x"5F",x"5B",x"5B",x"5B", -- 0x2CB8
    x"5B",x"3F",x"3F",x"3F",x"3F",x"3B",x"3B",x"3B", -- 0x2CC0
    x"3B",x"3F",x"3F",x"3F",x"3F",x"3B",x"3B",x"3B", -- 0x2CC8
    x"3B",x"3F",x"3F",x"3F",x"3F",x"3B",x"3B",x"3B", -- 0x2CD0
    x"3B",x"3F",x"3F",x"3F",x"3F",x"3B",x"3B",x"3B", -- 0x2CD8
    x"3B",x"1F",x"1F",x"1F",x"1F",x"1B",x"1B",x"1B", -- 0x2CE0
    x"1B",x"1F",x"1F",x"1F",x"1F",x"1B",x"1B",x"1B", -- 0x2CE8
    x"1B",x"1F",x"1F",x"1F",x"1F",x"1B",x"1B",x"1B", -- 0x2CF0
    x"1B",x"1F",x"1F",x"1F",x"1F",x"1B",x"1B",x"1B", -- 0x2CF8
    x"1B",x"FF",x"FE",x"FF",x"FE",x"FB",x"FA",x"FB", -- 0x2D00
    x"FA",x"FF",x"FE",x"FF",x"FE",x"FB",x"FA",x"FB", -- 0x2D08
    x"FA",x"FF",x"FE",x"FF",x"FE",x"FB",x"FA",x"FB", -- 0x2D10
    x"FA",x"FF",x"FE",x"FF",x"FE",x"FB",x"FA",x"FB", -- 0x2D18
    x"FA",x"DF",x"DE",x"DF",x"DE",x"DB",x"DA",x"DB", -- 0x2D20
    x"DA",x"DF",x"DE",x"DF",x"DE",x"DB",x"DA",x"DB", -- 0x2D28
    x"DA",x"DF",x"DE",x"DF",x"DE",x"DB",x"DA",x"DB", -- 0x2D30
    x"DA",x"DF",x"DE",x"DF",x"DE",x"DB",x"DA",x"DB", -- 0x2D38
    x"DA",x"BF",x"BE",x"BF",x"BE",x"BB",x"BA",x"BB", -- 0x2D40
    x"BA",x"BF",x"BE",x"BF",x"BE",x"BB",x"BA",x"BB", -- 0x2D48
    x"BA",x"BF",x"BE",x"BF",x"BE",x"BB",x"BA",x"BB", -- 0x2D50
    x"BA",x"BF",x"BE",x"BF",x"BE",x"BB",x"BA",x"BB", -- 0x2D58
    x"BA",x"9F",x"9E",x"9F",x"9E",x"9B",x"9A",x"9B", -- 0x2D60
    x"9A",x"9F",x"9E",x"9F",x"9E",x"9B",x"9A",x"9B", -- 0x2D68
    x"9A",x"9F",x"9E",x"9F",x"9E",x"9B",x"9A",x"9B", -- 0x2D70
    x"9A",x"9F",x"9E",x"9F",x"9E",x"9B",x"9A",x"9B", -- 0x2D78
    x"9A",x"7F",x"7E",x"7F",x"7E",x"7B",x"7A",x"7B", -- 0x2D80
    x"7A",x"7F",x"7E",x"7F",x"7E",x"7B",x"7A",x"7B", -- 0x2D88
    x"7A",x"7F",x"7E",x"7F",x"7E",x"7B",x"7A",x"7B", -- 0x2D90
    x"7A",x"7F",x"7E",x"7F",x"7E",x"7B",x"7A",x"7B", -- 0x2D98
    x"7A",x"5F",x"5E",x"5F",x"5E",x"5B",x"5A",x"5B", -- 0x2DA0
    x"5A",x"5F",x"5E",x"5F",x"5E",x"5B",x"5A",x"5B", -- 0x2DA8
    x"5A",x"5F",x"5E",x"5F",x"5E",x"5B",x"5A",x"5B", -- 0x2DB0
    x"5A",x"5F",x"5E",x"5F",x"5E",x"5B",x"5A",x"5B", -- 0x2DB8
    x"5A",x"3F",x"3E",x"3F",x"3E",x"3B",x"3A",x"3B", -- 0x2DC0
    x"3A",x"3F",x"3E",x"3F",x"3E",x"3B",x"3A",x"3B", -- 0x2DC8
    x"3A",x"3F",x"3E",x"3F",x"3E",x"3B",x"3A",x"3B", -- 0x2DD0
    x"3A",x"3F",x"3E",x"3F",x"3E",x"3B",x"3A",x"3B", -- 0x2DD8
    x"3A",x"1F",x"1E",x"1F",x"1E",x"1B",x"1A",x"1B", -- 0x2DE0
    x"1A",x"1F",x"1E",x"1F",x"1E",x"1B",x"1A",x"1B", -- 0x2DE8
    x"1A",x"1F",x"1E",x"1F",x"1E",x"1B",x"1A",x"1B", -- 0x2DF0
    x"1A",x"1F",x"1E",x"1F",x"1E",x"1B",x"1A",x"1B", -- 0x2DF8
    x"1A",x"FF",x"FF",x"FD",x"FD",x"FB",x"FB",x"F9", -- 0x2E00
    x"F9",x"FF",x"FF",x"FD",x"FD",x"FB",x"FB",x"F9", -- 0x2E08
    x"F9",x"FF",x"FF",x"FD",x"FD",x"FB",x"FB",x"F9", -- 0x2E10
    x"F9",x"FF",x"FF",x"FD",x"FD",x"FB",x"FB",x"F9", -- 0x2E18
    x"F9",x"DF",x"DF",x"DD",x"DD",x"DB",x"DB",x"D9", -- 0x2E20
    x"D9",x"DF",x"DF",x"DD",x"DD",x"DB",x"DB",x"D9", -- 0x2E28
    x"D9",x"DF",x"DF",x"DD",x"DD",x"DB",x"DB",x"D9", -- 0x2E30
    x"D9",x"DF",x"DF",x"DD",x"DD",x"DB",x"DB",x"D9", -- 0x2E38
    x"D9",x"BF",x"BF",x"BD",x"BD",x"BB",x"BB",x"B9", -- 0x2E40
    x"B9",x"BF",x"BF",x"BD",x"BD",x"BB",x"BB",x"B9", -- 0x2E48
    x"B9",x"BF",x"BF",x"BD",x"BD",x"BB",x"BB",x"B9", -- 0x2E50
    x"B9",x"BF",x"BF",x"BD",x"BD",x"BB",x"BB",x"B9", -- 0x2E58
    x"B9",x"9F",x"9F",x"9D",x"9D",x"9B",x"9B",x"99", -- 0x2E60
    x"99",x"9F",x"9F",x"9D",x"9D",x"9B",x"9B",x"99", -- 0x2E68
    x"99",x"9F",x"9F",x"9D",x"9D",x"9B",x"9B",x"99", -- 0x2E70
    x"99",x"9F",x"9F",x"9D",x"9D",x"9B",x"9B",x"99", -- 0x2E78
    x"99",x"7F",x"7F",x"7D",x"7D",x"7B",x"7B",x"79", -- 0x2E80
    x"79",x"7F",x"7F",x"7D",x"7D",x"7B",x"7B",x"79", -- 0x2E88
    x"79",x"7F",x"7F",x"7D",x"7D",x"7B",x"7B",x"79", -- 0x2E90
    x"79",x"7F",x"7F",x"7D",x"7D",x"7B",x"7B",x"79", -- 0x2E98
    x"79",x"5F",x"5F",x"5D",x"5D",x"5B",x"5B",x"59", -- 0x2EA0
    x"59",x"5F",x"5F",x"5D",x"5D",x"5B",x"5B",x"59", -- 0x2EA8
    x"59",x"5F",x"5F",x"5D",x"5D",x"5B",x"5B",x"59", -- 0x2EB0
    x"59",x"5F",x"5F",x"5D",x"5D",x"5B",x"5B",x"59", -- 0x2EB8
    x"59",x"3F",x"3F",x"3D",x"3D",x"3B",x"3B",x"39", -- 0x2EC0
    x"39",x"3F",x"3F",x"3D",x"3D",x"3B",x"3B",x"39", -- 0x2EC8
    x"39",x"3F",x"3F",x"3D",x"3D",x"3B",x"3B",x"39", -- 0x2ED0
    x"39",x"3F",x"3F",x"3D",x"3D",x"3B",x"3B",x"39", -- 0x2ED8
    x"39",x"1F",x"1F",x"1D",x"1D",x"1B",x"1B",x"19", -- 0x2EE0
    x"19",x"1F",x"1F",x"1D",x"1D",x"1B",x"1B",x"19", -- 0x2EE8
    x"19",x"1F",x"1F",x"1D",x"1D",x"1B",x"1B",x"19", -- 0x2EF0
    x"19",x"1F",x"1F",x"1D",x"1D",x"1B",x"1B",x"19", -- 0x2EF8
    x"19",x"FF",x"FE",x"FD",x"FC",x"FB",x"FA",x"F9", -- 0x2F00
    x"F8",x"FF",x"FE",x"FD",x"FC",x"FB",x"FA",x"F9", -- 0x2F08
    x"F8",x"FF",x"FE",x"FD",x"FC",x"FB",x"FA",x"F9", -- 0x2F10
    x"F8",x"FF",x"FE",x"FD",x"FC",x"FB",x"FA",x"F9", -- 0x2F18
    x"F8",x"DF",x"DE",x"DD",x"DC",x"DB",x"DA",x"D9", -- 0x2F20
    x"D8",x"DF",x"DE",x"DD",x"DC",x"DB",x"DA",x"D9", -- 0x2F28
    x"D8",x"DF",x"DE",x"DD",x"DC",x"DB",x"DA",x"D9", -- 0x2F30
    x"D8",x"DF",x"DE",x"DD",x"DC",x"DB",x"DA",x"D9", -- 0x2F38
    x"D8",x"BF",x"BE",x"BD",x"BC",x"BB",x"BA",x"B9", -- 0x2F40
    x"B8",x"BF",x"BE",x"BD",x"BC",x"BB",x"BA",x"B9", -- 0x2F48
    x"B8",x"BF",x"BE",x"BD",x"BC",x"BB",x"BA",x"B9", -- 0x2F50
    x"B8",x"BF",x"BE",x"BD",x"BC",x"BB",x"BA",x"B9", -- 0x2F58
    x"B8",x"9F",x"9E",x"9D",x"9C",x"9B",x"9A",x"99", -- 0x2F60
    x"98",x"9F",x"9E",x"9D",x"9C",x"9B",x"9A",x"99", -- 0x2F68
    x"98",x"9F",x"9E",x"9D",x"9C",x"9B",x"9A",x"99", -- 0x2F70
    x"98",x"9F",x"9E",x"9D",x"9C",x"9B",x"9A",x"99", -- 0x2F78
    x"98",x"7F",x"7E",x"7D",x"7C",x"7B",x"7A",x"79", -- 0x2F80
    x"78",x"7F",x"7E",x"7D",x"7C",x"7B",x"7A",x"79", -- 0x2F88
    x"78",x"7F",x"7E",x"7D",x"7C",x"7B",x"7A",x"79", -- 0x2F90
    x"78",x"7F",x"7E",x"7D",x"7C",x"7B",x"7A",x"79", -- 0x2F98
    x"78",x"5F",x"5E",x"5D",x"5C",x"5B",x"5A",x"59", -- 0x2FA0
    x"58",x"5F",x"5E",x"5D",x"5C",x"5B",x"5A",x"59", -- 0x2FA8
    x"58",x"5F",x"5E",x"5D",x"5C",x"5B",x"5A",x"59", -- 0x2FB0
    x"58",x"5F",x"5E",x"5D",x"5C",x"5B",x"5A",x"59", -- 0x2FB8
    x"58",x"3F",x"3E",x"3D",x"3C",x"3B",x"3A",x"39", -- 0x2FC0
    x"38",x"3F",x"3E",x"3D",x"3C",x"3B",x"3A",x"39", -- 0x2FC8
    x"38",x"3F",x"3E",x"3D",x"3C",x"3B",x"3A",x"39", -- 0x2FD0
    x"38",x"3F",x"3E",x"3D",x"3C",x"3B",x"3A",x"39", -- 0x2FD8
    x"38",x"1F",x"1E",x"1D",x"1C",x"1B",x"1A",x"19", -- 0x2FE0
    x"18",x"1F",x"1E",x"1D",x"1C",x"1B",x"1A",x"19", -- 0x2FE8
    x"18",x"1F",x"1E",x"1D",x"1C",x"1B",x"1A",x"19", -- 0x2FF0
    x"18",x"1F",x"1E",x"1D",x"1C",x"1B",x"1A",x"19"  -- 0x2FF8
  );
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;

