library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity jng_chr_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of jng_chr_rom is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"80",X"C0",X"20",X"20",X"60",X"C0",X"80",X"00",X"30",X"70",X"C0",X"80",X"80",X"70",X"30",X"00",
		X"20",X"20",X"E0",X"E0",X"20",X"20",X"00",X"00",X"00",X"00",X"F0",X"F0",X"40",X"00",X"00",X"00",
		X"20",X"20",X"A0",X"A0",X"E0",X"E0",X"60",X"00",X"60",X"F0",X"B0",X"90",X"90",X"C0",X"40",X"00",
		X"C0",X"E0",X"20",X"20",X"20",X"60",X"40",X"00",X"80",X"D0",X"F0",X"B0",X"90",X"80",X"00",X"00",
		X"80",X"E0",X"E0",X"80",X"80",X"80",X"80",X"00",X"00",X"F0",X"F0",X"C0",X"60",X"30",X"10",X"00",
		X"C0",X"E0",X"20",X"20",X"20",X"60",X"40",X"00",X"10",X"B0",X"A0",X"A0",X"A0",X"E0",X"E0",X"00",
		X"C0",X"E0",X"20",X"20",X"20",X"E0",X"C0",X"00",X"00",X"90",X"90",X"90",X"D0",X"70",X"30",X"00",
		X"00",X"00",X"00",X"E0",X"E0",X"00",X"00",X"00",X"C0",X"E0",X"B0",X"90",X"80",X"C0",X"C0",X"00",
		X"C0",X"E0",X"A0",X"A0",X"20",X"20",X"C0",X"00",X"00",X"60",X"90",X"90",X"B0",X"F0",X"60",X"00",
		X"80",X"C0",X"60",X"20",X"20",X"20",X"00",X"00",X"70",X"F0",X"90",X"90",X"90",X"F0",X"60",X"00",
		X"40",X"40",X"20",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"10",X"20",X"20",
		X"40",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"40",
		X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"40",
		X"00",X"00",X"00",X"00",X"90",X"F0",X"52",X"61",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"F0",X"A4",X"68",
		X"30",X"20",X"28",X"28",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"40",X"41",X"41",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"00",X"F0",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"E0",X"A4",X"78",
		X"10",X"F0",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"78",X"A4",X"E0",X"30",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"28",X"28",X"20",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"41",X"41",X"40",X"E0",
		X"61",X"52",X"F0",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"68",X"A4",X"F0",X"90",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"70",X"52",X"E1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"F0",X"80",
		X"E1",X"52",X"70",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"F0",X"00",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"81",X"F0",X"D2",X"61",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"F0",X"B4",X"68",
		X"30",X"10",X"18",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",X"81",X"81",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"00",X"10",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"E0",X"A4",X"69",
		X"F0",X"10",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"69",X"A4",X"E0",X"70",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"18",X"18",X"10",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"81",X"81",X"80",X"C0",
		X"61",X"D2",X"F0",X"81",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"68",X"B4",X"F0",X"18",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"E0",X"70",X"52",X"69",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"80",X"F0",
		X"69",X"52",X"70",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"80",X"00",X"03",X"00",X"00",X"00",X"00",
		X"00",X"77",X"44",X"44",X"77",X"00",X"77",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"22",X"22",X"EE",X"00",X"EE",X"22",
		X"44",X"77",X"00",X"55",X"55",X"55",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"EE",X"00",X"EE",X"22",X"22",X"22",X"00",
		X"00",X"E0",X"C0",X"C2",X"C2",X"C0",X"E0",X"00",X"00",X"04",X"10",X"61",X"61",X"10",X"04",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"80",X"80",X"80",X"E0",X"E0",X"00",X"30",X"70",X"C0",X"80",X"C0",X"70",X"30",X"00",
		X"C0",X"E0",X"20",X"20",X"20",X"E0",X"E0",X"00",X"60",X"F0",X"90",X"90",X"90",X"F0",X"F0",X"00",
		X"40",X"60",X"20",X"20",X"60",X"C0",X"80",X"00",X"40",X"C0",X"80",X"80",X"C0",X"70",X"30",X"00",
		X"80",X"C0",X"60",X"20",X"20",X"E0",X"E0",X"00",X"30",X"70",X"C0",X"80",X"80",X"F0",X"F0",X"00",
		X"20",X"20",X"20",X"20",X"E0",X"E0",X"00",X"00",X"80",X"90",X"90",X"90",X"F0",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"00",X"80",X"90",X"90",X"90",X"90",X"F0",X"F0",X"00",
		X"E0",X"E0",X"20",X"20",X"60",X"C0",X"80",X"00",X"90",X"90",X"90",X"80",X"C0",X"70",X"30",X"00",
		X"E0",X"E0",X"00",X"00",X"00",X"E0",X"E0",X"00",X"F0",X"F0",X"10",X"10",X"10",X"F0",X"F0",X"00",
		X"20",X"20",X"E0",X"E0",X"20",X"20",X"00",X"00",X"80",X"80",X"F0",X"F0",X"80",X"80",X"00",X"00",
		X"C0",X"E0",X"20",X"20",X"20",X"60",X"40",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"60",X"E0",X"C0",X"80",X"E0",X"E0",X"00",X"80",X"C0",X"60",X"30",X"10",X"F0",X"F0",X"00",
		X"20",X"20",X"20",X"20",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",
		X"E0",X"E0",X"00",X"80",X"00",X"E0",X"E0",X"00",X"F0",X"F0",X"70",X"30",X"70",X"F0",X"F0",X"00",
		X"E0",X"E0",X"C0",X"80",X"00",X"E0",X"E0",X"00",X"F0",X"F0",X"10",X"30",X"70",X"F0",X"F0",X"00",
		X"C0",X"E0",X"20",X"20",X"20",X"E0",X"C0",X"00",X"70",X"F0",X"80",X"80",X"80",X"F0",X"70",X"00",
		X"00",X"80",X"80",X"80",X"80",X"E0",X"E0",X"00",X"70",X"F0",X"80",X"80",X"80",X"F0",X"F0",X"00",
		X"A0",X"C0",X"E0",X"A0",X"20",X"E0",X"C0",X"00",X"70",X"F0",X"80",X"80",X"80",X"F0",X"70",X"00",
		X"20",X"60",X"E0",X"C0",X"80",X"E0",X"E0",X"00",X"70",X"F0",X"90",X"80",X"80",X"F0",X"F0",X"00",
		X"C0",X"E0",X"20",X"20",X"20",X"60",X"40",X"00",X"00",X"50",X"D0",X"90",X"90",X"F0",X"60",X"00",
		X"00",X"00",X"E0",X"E0",X"00",X"00",X"00",X"00",X"80",X"80",X"F0",X"F0",X"80",X"80",X"00",X"00",
		X"C0",X"E0",X"20",X"20",X"20",X"E0",X"C0",X"00",X"F0",X"F0",X"00",X"00",X"00",X"F0",X"F0",X"00",
		X"00",X"80",X"C0",X"E0",X"C0",X"80",X"00",X"00",X"F0",X"F0",X"10",X"00",X"10",X"F0",X"F0",X"00",
		X"E0",X"E0",X"C0",X"80",X"C0",X"E0",X"E0",X"00",X"F0",X"F0",X"10",X"30",X"10",X"F0",X"F0",X"00",
		X"60",X"E0",X"C0",X"80",X"C0",X"E0",X"60",X"00",X"C0",X"E0",X"70",X"30",X"70",X"E0",X"C0",X"00",
		X"00",X"00",X"E0",X"E0",X"00",X"00",X"00",X"00",X"E0",X"F0",X"10",X"10",X"F0",X"E0",X"00",X"00",
		X"20",X"20",X"20",X"A0",X"E0",X"E0",X"60",X"00",X"C0",X"E0",X"F0",X"B0",X"90",X"80",X"80",X"00",
		X"00",X"00",X"00",X"60",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"20",X"10",X"50",X"50",X"90",X"20",X"C0",X"30",X"40",X"80",X"A0",X"A0",X"90",X"40",X"30",
		X"C0",X"E8",X"E4",X"E0",X"E0",X"E0",X"C0",X"00",X"30",X"79",X"78",X"FC",X"78",X"78",X"30",X"00",
		X"E0",X"C0",X"68",X"E0",X"68",X"C0",X"E0",X"00",X"00",X"10",X"F0",X"21",X"F0",X"10",X"00",X"00",
		X"C0",X"20",X"80",X"C0",X"80",X"20",X"C0",X"00",X"10",X"30",X"70",X"F0",X"70",X"30",X"10",X"00",
		X"00",X"00",X"00",X"00",X"10",X"00",X"3F",X"56",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"4F",X"A6",
		X"25",X"2A",X"8B",X"26",X"15",X"00",X"00",X"00",X"11",X"11",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A2",X"4C",X"84",X"82",X"88",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"3B",X"AC",X"8A",X"98",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"08",X"88",X"88",X"00",X"00",X"00",X"00",X"04",X"15",X"8B",X"14",X"18",
		X"51",X"46",X"0D",X"A9",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",
		X"04",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"8B",X"E2",X"26",X"C6",X"09",X"08",X"00",X"00",
		X"00",X"00",X"11",X"2A",X"49",X"21",X"95",X"45",X"00",X"02",X"01",X"00",X"00",X"11",X"23",X"22",
		X"00",X"00",X"00",X"00",X"02",X"0C",X"88",X"88",X"00",X"02",X"8A",X"45",X"C6",X"11",X"AD",X"C4",
		X"5C",X"26",X"90",X"04",X"8A",X"01",X"01",X"00",X"11",X"01",X"02",X"13",X"04",X"00",X"00",X"00",
		X"00",X"06",X"08",X"00",X"00",X"08",X"08",X"00",X"A8",X"0A",X"91",X"66",X"81",X"00",X"00",X"00",
		X"00",X"18",X"AC",X"84",X"13",X"38",X"91",X"23",X"01",X"00",X"11",X"2E",X"47",X"54",X"40",X"06",
		X"09",X"0A",X"02",X"05",X"08",X"00",X"0C",X"03",X"04",X"04",X"05",X"CE",X"3E",X"31",X"39",X"89",
		X"2F",X"59",X"42",X"A8",X"6F",X"10",X"01",X"01",X"3A",X"32",X"11",X"05",X"08",X"01",X"01",X"01",
		X"88",X"C4",X"4C",X"8E",X"01",X"00",X"00",X"00",X"BA",X"32",X"4D",X"06",X"B3",X"4A",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"04",X"00",X"64",X"00",X"40",X"02",X"00",X"18",X"40",X"01",X"D5",X"01",X"04",X"18",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"18",X"F0",X"B4",X"68",X"C0",X"80",X"81",X"81",X"81",X"F0",X"D2",X"61",X"30",X"10",X"18",X"18",
		X"90",X"F0",X"A4",X"68",X"C0",X"40",X"41",X"41",X"90",X"F0",X"52",X"61",X"30",X"20",X"28",X"28",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"21",X"43",X"53",X"E1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"0C",X"0E",X"4F",
		X"D3",X"61",X"43",X"21",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"2E",X"8C",X"08",X"00",X"00",X"00",X"00",
		X"00",X"80",X"C0",X"E0",X"E0",X"C0",X"80",X"00",X"00",X"10",X"30",X"70",X"70",X"30",X"10",X"00",
		X"80",X"C0",X"E0",X"E0",X"C0",X"80",X"00",X"00",X"10",X"30",X"70",X"70",X"30",X"10",X"00",X"00",
		X"C0",X"E0",X"E0",X"E0",X"C0",X"00",X"00",X"08",X"70",X"70",X"70",X"30",X"10",X"00",X"00",X"03",
		X"E0",X"E0",X"E0",X"C0",X"00",X"00",X"08",X"0C",X"70",X"70",X"30",X"10",X"00",X"00",X"03",X"07",
		X"E0",X"C0",X"80",X"00",X"00",X"08",X"0C",X"0E",X"70",X"30",X"10",X"00",X"00",X"01",X"03",X"07",
		X"C0",X"80",X"00",X"00",X"08",X"0C",X"0E",X"0E",X"30",X"10",X"00",X"00",X"01",X"03",X"07",X"07",
		X"80",X"00",X"00",X"0C",X"0E",X"0E",X"0E",X"0C",X"30",X"00",X"00",X"01",X"03",X"07",X"07",X"07",
		X"00",X"00",X"0C",X"0E",X"0E",X"0E",X"0C",X"08",X"00",X"00",X"01",X"03",X"07",X"07",X"07",X"03",
		X"00",X"80",X"C0",X"E0",X"E0",X"C0",X"80",X"00",X"00",X"10",X"30",X"70",X"70",X"30",X"10",X"00",
		X"00",X"00",X"80",X"C0",X"C0",X"80",X"00",X"00",X"00",X"30",X"70",X"F0",X"F0",X"70",X"30",X"00",
		X"00",X"00",X"80",X"81",X"81",X"01",X"00",X"00",X"00",X"70",X"F0",X"F0",X"F0",X"F0",X"E0",X"00",
		X"00",X"00",X"01",X"03",X"03",X"03",X"01",X"00",X"00",X"E0",X"F0",X"F0",X"F0",X"E0",X"C0",X"00",
		X"00",X"01",X"03",X"07",X"07",X"03",X"01",X"00",X"00",X"80",X"C0",X"E0",X"E0",X"C0",X"80",X"00",
		X"00",X"03",X"07",X"0F",X"0F",X"07",X"03",X"00",X"00",X"00",X"80",X"C0",X"C0",X"80",X"00",X"00",
		X"00",X"0E",X"0F",X"0F",X"0F",X"0F",X"07",X"00",X"00",X"00",X"01",X"81",X"81",X"80",X"00",X"00",
		X"00",X"0C",X"0E",X"0F",X"0F",X"0F",X"0E",X"00",X"00",X"01",X"03",X"03",X"03",X"01",X"00",X"00",
		X"C0",X"E0",X"F0",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"10",X"30",X"30",X"10",X"00",X"00",X"00",
		X"80",X"C0",X"E0",X"E0",X"C0",X"80",X"00",X"00",X"10",X"30",X"70",X"70",X"30",X"10",X"00",X"00",
		X"C0",X"E0",X"E0",X"C1",X"81",X"00",X"00",X"00",X"30",X"70",X"70",X"30",X"10",X"00",X"00",X"00",
		X"E0",X"E0",X"C1",X"83",X"03",X"01",X"00",X"00",X"70",X"70",X"30",X"10",X"00",X"00",X"00",X"00",
		X"E0",X"C1",X"83",X"07",X"07",X"03",X"01",X"00",X"70",X"30",X"10",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"83",X"07",X"0F",X"0F",X"07",X"03",X"00",X"30",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"06",X"0F",X"0F",X"0F",X"0F",X"06",X"00",X"10",X"00",X"00",X"01",X"01",X"00",X"00",X"00",
		X"00",X"0C",X"0E",X"0F",X"0F",X"0E",X"0C",X"00",X"00",X"00",X"01",X"03",X"03",X"01",X"00",X"00",
		X"C0",X"E0",X"F0",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"10",X"30",X"30",X"10",X"00",X"00",X"00",
		X"00",X"C0",X"E0",X"F0",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"10",X"30",X"30",X"10",X"00",X"00",
		X"08",X"60",X"F0",X"F0",X"F0",X"F0",X"60",X"00",X"01",X"00",X"00",X"10",X"10",X"00",X"00",X"00",
		X"0C",X"38",X"70",X"F0",X"F0",X"70",X"30",X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"1C",X"38",X"70",X"70",X"30",X"10",X"00",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"0E",X"1C",X"38",X"30",X"10",X"00",X"00",X"07",X"07",X"03",X"01",X"00",X"00",X"00",X"00",
		X"0C",X"0E",X"0E",X"1C",X"18",X"00",X"00",X"00",X"03",X"07",X"07",X"03",X"01",X"00",X"00",X"00",
		X"08",X"0C",X"0E",X"0E",X"0C",X"08",X"00",X"00",X"01",X"03",X"07",X"07",X"03",X"01",X"00",X"00",
		X"00",X"80",X"C0",X"E0",X"E0",X"C0",X"80",X"00",X"00",X"10",X"30",X"70",X"70",X"30",X"10",X"00",
		X"80",X"C0",X"E0",X"E0",X"C0",X"80",X"00",X"00",X"10",X"30",X"70",X"70",X"30",X"10",X"00",X"00",
		X"C0",X"E0",X"E0",X"E0",X"C0",X"00",X"00",X"08",X"70",X"70",X"70",X"30",X"10",X"00",X"00",X"01",
		X"E0",X"E0",X"E0",X"C0",X"00",X"00",X"08",X"0C",X"70",X"70",X"30",X"10",X"00",X"00",X"01",X"03",
		X"E0",X"C0",X"80",X"00",X"00",X"08",X"0C",X"0E",X"70",X"30",X"10",X"00",X"00",X"01",X"03",X"07",
		X"C0",X"80",X"00",X"00",X"08",X"0C",X"0E",X"0F",X"30",X"10",X"00",X"00",X"01",X"03",X"07",X"0F",
		X"80",X"00",X"00",X"08",X"0C",X"0E",X"0F",X"0D",X"30",X"00",X"00",X"01",X"03",X"07",X"0F",X"0B",
		X"00",X"00",X"08",X"0C",X"0E",X"0F",X"0D",X"09",X"00",X"00",X"01",X"03",X"07",X"0F",X"0B",X"09",
		X"00",X"80",X"C0",X"E0",X"E0",X"C0",X"80",X"00",X"00",X"10",X"30",X"70",X"70",X"30",X"10",X"00",
		X"00",X"00",X"80",X"C0",X"C0",X"80",X"00",X"00",X"00",X"30",X"70",X"F0",X"F0",X"70",X"30",X"00",
		X"00",X"00",X"80",X"81",X"81",X"00",X"00",X"00",X"00",X"70",X"F0",X"F0",X"F0",X"F0",X"E0",X"00",
		X"00",X"00",X"01",X"03",X"03",X"01",X"00",X"00",X"00",X"E0",X"F0",X"F0",X"F0",X"E0",X"C0",X"00",
		X"00",X"01",X"03",X"07",X"07",X"03",X"01",X"00",X"00",X"80",X"C0",X"E0",X"E0",X"C0",X"80",X"00",
		X"01",X"03",X"07",X"0F",X"0F",X"07",X"03",X"01",X"00",X"00",X"80",X"C0",X"C0",X"80",X"00",X"00",
		X"03",X"06",X"0F",X"0F",X"0F",X"0F",X"06",X"03",X"00",X"00",X"00",X"81",X"81",X"80",X"00",X"00",
		X"07",X"0C",X"0E",X"0F",X"0F",X"0E",X"0C",X"07",X"00",X"00",X"01",X"03",X"03",X"01",X"00",X"00",
		X"C0",X"E0",X"F0",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"10",X"30",X"30",X"10",X"00",X"00",X"00",
		X"80",X"C0",X"E0",X"E0",X"C0",X"80",X"00",X"00",X"10",X"30",X"70",X"70",X"30",X"10",X"00",X"00",
		X"C0",X"E0",X"E0",X"C1",X"81",X"00",X"00",X"00",X"30",X"70",X"70",X"30",X"10",X"00",X"00",X"00",
		X"E0",X"E0",X"C1",X"83",X"03",X"01",X"00",X"00",X"70",X"70",X"30",X"10",X"00",X"00",X"00",X"00",
		X"E0",X"C1",X"83",X"07",X"07",X"03",X"01",X"00",X"70",X"30",X"10",X"00",X"00",X"00",X"00",X"00",
		X"C1",X"83",X"07",X"0F",X"0F",X"07",X"03",X"01",X"30",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"83",X"06",X"0F",X"0F",X"0F",X"0F",X"06",X"03",X"10",X"00",X"00",X"01",X"01",X"00",X"00",X"00",
		X"07",X"0C",X"0E",X"0F",X"0F",X"0E",X"0C",X"07",X"00",X"00",X"01",X"03",X"03",X"01",X"00",X"00",
		X"C0",X"E0",X"F0",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"10",X"30",X"30",X"10",X"00",X"00",X"00",
		X"00",X"C0",X"E0",X"F0",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"10",X"30",X"30",X"10",X"00",X"00",
		X"08",X"60",X"F0",X"F0",X"F0",X"F0",X"60",X"00",X"01",X"00",X"00",X"10",X"10",X"00",X"00",X"00",
		X"0C",X"38",X"70",X"F0",X"F0",X"70",X"30",X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"1C",X"38",X"70",X"70",X"30",X"10",X"00",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0E",X"1C",X"38",X"30",X"10",X"00",X"00",X"0F",X"07",X"03",X"01",X"00",X"00",X"00",X"00",
		X"0D",X"0F",X"0E",X"1C",X"18",X"00",X"00",X"00",X"0B",X"0F",X"07",X"03",X"01",X"00",X"00",X"00",
		X"09",X"0D",X"0F",X"0E",X"0C",X"08",X"00",X"00",X"09",X"0B",X"0F",X"07",X"03",X"01",X"00",X"00",
		X"00",X"80",X"C0",X"E0",X"F0",X"D0",X"90",X"20",X"00",X"10",X"30",X"70",X"F0",X"B0",X"90",X"40",
		X"80",X"C0",X"E0",X"F0",X"D0",X"90",X"20",X"00",X"10",X"30",X"70",X"F0",X"B0",X"90",X"40",X"00",
		X"C0",X"E0",X"F0",X"D0",X"90",X"20",X"00",X"00",X"30",X"70",X"F0",X"B0",X"90",X"40",X"00",X"00",
		X"E0",X"F0",X"D0",X"90",X"20",X"00",X"00",X"00",X"70",X"F0",X"B0",X"90",X"40",X"00",X"00",X"00",
		X"F0",X"D0",X"90",X"20",X"00",X"00",X"00",X"00",X"F0",X"B0",X"90",X"40",X"00",X"00",X"00",X"00",
		X"D0",X"90",X"20",X"00",X"00",X"00",X"00",X"00",X"B0",X"90",X"40",X"00",X"00",X"00",X"00",X"00",
		X"90",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"90",X"C0",X"E0",X"E0",X"C0",X"90",X"E0",X"00",X"10",X"30",X"70",X"70",X"30",X"10",X"00",
		X"C0",X"20",X"80",X"C0",X"C0",X"80",X"20",X"C0",X"10",X"30",X"70",X"F0",X"F0",X"70",X"30",X"10",
		X"80",X"40",X"00",X"80",X"80",X"00",X"40",X"80",X"30",X"60",X"F0",X"F0",X"F0",X"F0",X"60",X"30",
		X"00",X"80",X"00",X"00",X"00",X"00",X"80",X"00",X"70",X"C0",X"E0",X"F0",X"F0",X"E0",X"C0",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"90",X"C0",X"E0",X"E0",X"C0",X"90",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"20",X"80",X"C0",X"C0",X"80",X"20",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"00",X"80",X"80",X"00",X"40",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"80",X"00",
		X"80",X"C0",X"E0",X"F0",X"D0",X"90",X"20",X"00",X"10",X"30",X"70",X"F0",X"B0",X"90",X"40",X"00",
		X"80",X"C0",X"E0",X"F0",X"D0",X"90",X"20",X"00",X"10",X"30",X"70",X"F0",X"B0",X"90",X"40",X"00",
		X"C0",X"E0",X"F0",X"D0",X"90",X"20",X"00",X"00",X"30",X"70",X"F0",X"B0",X"90",X"40",X"00",X"00",
		X"E0",X"F0",X"D0",X"90",X"20",X"00",X"00",X"00",X"70",X"F0",X"B0",X"90",X"40",X"00",X"00",X"00",
		X"F0",X"D0",X"90",X"20",X"00",X"00",X"00",X"00",X"F0",X"B0",X"90",X"40",X"00",X"00",X"00",X"00",
		X"D0",X"90",X"20",X"00",X"00",X"00",X"00",X"00",X"B0",X"90",X"40",X"00",X"00",X"00",X"00",X"00",
		X"90",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"C0",X"E0",X"F0",X"F0",X"E0",X"C0",X"80",X"30",X"40",X"10",X"30",X"30",X"10",X"40",X"30",
		X"80",X"C0",X"E0",X"F0",X"F0",X"E0",X"C0",X"80",X"30",X"40",X"10",X"30",X"30",X"10",X"40",X"30",
		X"C0",X"60",X"F0",X"F0",X"F0",X"F0",X"60",X"C0",X"10",X"20",X"00",X"10",X"10",X"00",X"20",X"10",
		X"E0",X"30",X"70",X"F0",X"F0",X"70",X"30",X"E0",X"00",X"10",X"00",X"00",X"00",X"00",X"10",X"00",
		X"70",X"90",X"30",X"70",X"70",X"30",X"90",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"40",X"10",X"30",X"30",X"10",X"40",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"20",X"00",X"10",X"10",X"00",X"20",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"50",X"A0",X"50",X"A0",X"50",X"A0",X"F0",X"00",X"50",X"60",X"50",X"60",X"50",X"20",X"10",X"00",
		X"00",X"F0",X"A0",X"50",X"A0",X"50",X"A0",X"50",X"00",X"10",X"20",X"50",X"60",X"50",X"60",X"50",
		X"A0",X"60",X"A0",X"60",X"A0",X"40",X"80",X"00",X"A0",X"50",X"A0",X"50",X"A0",X"50",X"F0",X"00",
		X"00",X"80",X"40",X"A0",X"60",X"A0",X"60",X"A0",X"00",X"F0",X"50",X"A0",X"50",X"A0",X"50",X"A0",
		X"A0",X"50",X"A0",X"50",X"A0",X"50",X"F0",X"00",X"A0",X"50",X"A0",X"50",X"A0",X"50",X"F0",X"00",
		X"00",X"F0",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"00",X"F0",X"50",X"A0",X"50",X"A0",X"50",X"A0",
		X"A0",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"50",X"60",X"50",X"60",X"50",X"60",X"50",X"60",X"50",
		X"60",X"A0",X"60",X"A0",X"60",X"A0",X"60",X"A0",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"50",X"A0",
		X"50",X"A0",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"50",X"20",
		X"A0",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"50",X"20",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"50",
		X"A0",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"40",X"A0",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"50",
		X"40",X"A0",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"50",X"A0",
		X"A0",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"50",
		X"C0",X"20",X"50",X"90",X"90",X"50",X"20",X"C0",X"30",X"40",X"A0",X"90",X"90",X"A0",X"40",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"40",X"20",X"90",X"20",X"40",X"20",X"90",X"50",X"A0",X"50",X"20",X"50",X"A0",X"50",X"20",
		X"20",X"50",X"A0",X"50",X"80",X"20",X"50",X"80",X"20",X"50",X"A0",X"50",X"80",X"20",X"50",X"80",
		X"20",X"50",X"A0",X"50",X"00",X"20",X"10",X"A0",X"20",X"90",X"40",X"20",X"50",X"A0",X"50",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
