library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity guzzler_big_sprite_tile_bit0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of guzzler_big_sprite_tile_bit0 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",X"30",X"20",X"00",X"00",X"00",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"0C",X"04",X"00",X"00",X"00",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"C0",X"00",X"00",X"00",X"00",X"00",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"FF",X"F8",X"00",X"00",X"00",X"00",X"00",X"80",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E0",X"C0",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"80",X"E0",X"F8",X"FE",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"1F",X"0F",X"07",X"03",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"80",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"F8",X"FF",X"FC",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"38",X"70",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"3C",
		X"F8",X"FC",X"FF",X"FF",X"FC",X"F8",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"F8",X"F8",X"F0",X"F0",X"F0",
		X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F8",X"F8",X"FC",X"FE",X"FF",X"7F",
		X"F8",X"F8",X"00",X"00",X"00",X"00",X"00",X"F0",X"FC",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F8",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FC",X"F8",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FC",X"FF",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"7F",X"07",X"00",X"00",X"00",X"00",X"00",X"07",X"03",X"00",X"00",X"00",X"00",X"80",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"78",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FF",X"FF",X"0F",X"00",X"FC",X"FE",X"FF",X"0F",X"00",X"00",X"00",X"00",
		X"07",X"03",X"01",X"00",X"00",X"60",X"F0",X"F8",X"FC",X"FE",X"FF",X"FF",X"7F",X"3F",X"1F",X"0F",
		X"07",X"03",X"01",X"00",X"00",X"60",X"F0",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"0F",
		X"00",X"00",X"F0",X"3F",X"00",X"00",X"00",X"00",X"F0",X"F0",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"0F",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",
		X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"01",X"03",X"07",X"0F",X"7F",X"FF",X"FF",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"61",X"3F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"03",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"01",X"01",
		X"07",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",
		X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BF",X"BF",X"00",X"00",X"00",X"00",X"00",X"FF",X"81",X"CF",X"E7",X"F3",X"E7",X"CF",X"81",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"1F",X"0F",X"0F",X"07",X"03",X"01",X"00",
		X"3F",X"7F",X"7F",X"7F",X"7F",X"7F",X"3F",X"3F",X"00",X"00",X"03",X"07",X"0F",X"1F",X"3F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"3F",X"3F",X"7F",X"7F",X"7F",X"3F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",X"F8",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FE",X"E0",X"C0",X"C0",X"C0",X"E0",X"F0",X"00",X"70",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"1F",X"03",X"00",X"00",X"00",X"00",X"00",X"E0",X"FC",X"FF",X"FF",X"FF",
		X"01",X"03",X"07",X"07",X"07",X"03",X"03",X"01",X"07",X"03",X"01",X"00",X"80",X"80",X"80",X"80",
		X"01",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"07",X"03",X"00",X"01",X"03",X"07",X"07",X"03",
		X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"00",X"00",X"00",X"01",X"03",X"03",X"07",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"7E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"03",X"03",X"01",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"03",X"07",X"07",X"07",X"07",X"00",X"01",X"03",X"07",X"07",X"07",X"07",X"02",
		X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"07",X"07",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"00",X"7C",X"00",X"00",X"00",X"00",X"C0",X"FC",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"00",X"07",X"3F",X"FF",
		X"FF",X"01",X"00",X"00",X"00",X"E0",X"FE",X"FF",X"FE",X"FE",X"02",X"F8",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"00",X"00",X"F0",X"FC",X"FE",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"07",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F0",X"FF",X"FF",X"FF",X"FF",X"E0",X"F0",X"F8",X"FE",X"FF",X"3F",X"0F",X"03",
		X"FE",X"FF",X"FF",X"E0",X"C0",X"C0",X"C0",X"C0",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"1F",X"07",X"03",X"00",X"1F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"01",X"00",X"FF",X"FF",X"FF",X"00",X"7F",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"E0",X"FF",X"FF",X"FF",
		X"E0",X"F0",X"F8",X"FC",X"0F",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"7F",X"03",X"00",X"00",
		X"7F",X"07",X"00",X"00",X"80",X"FF",X"FF",X"FF",X"07",X"07",X"07",X"0F",X"FF",X"FF",X"FE",X"FF",
		X"1F",X"C0",X"F0",X"F8",X"3C",X"0E",X"06",X"07",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F8",X"C0",X"80",X"80",X"80",X"80",X"80",X"C0",X"00",X"F8",X"FC",X"FE",X"FE",X"FE",X"FE",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"80",X"00",X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FE",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"3F",X"3F",X"3F",X"3F",X"7F",X"FF",X"7F",X"3F",X"3F",X"3F",X"07",X"F0",X"FF",
		X"1F",X"1F",X"1F",X"3F",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"07",X"0F",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"F0",X"E0",X"00",X"00",
		X"CE",X"EF",X"0F",X"0F",X"1F",X"FF",X"FF",X"FF",X"87",X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"90",
		X"FF",X"00",X"1C",X"0F",X"07",X"07",X"07",X"07",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"F8",X"F0",X"E0",X"00",X"00",X"00",X"00",X"C0",X"F0",X"F8",X"FC",X"FE",X"FE",X"FE",X"FE",
		X"FC",X"FE",X"FE",X"FE",X"0C",X"00",X"00",X"80",X"FE",X"FC",X"FC",X"F8",X"00",X"E0",X"F0",X"F8",
		X"E0",X"F0",X"F8",X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"FC",X"F8",X"70",X"00",
		X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",X"00",X"00",X"00",X"00",X"F0",X"F8",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FC",X"FC",X"F8",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"F0",X"F8",X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FC",X"F8",X"F0",
		X"F8",X"00",X"00",X"80",X"E0",X"F8",X"FC",X"FE",X"00",X"F8",X"FC",X"FE",X"FE",X"FE",X"FE",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"78",X"78",X"30",X"00",X"00",X"00",X"00",X"3F",X"3F",X"7F",X"FF",X"9F",X"8F",X"86",X"C0",
		X"1F",X"1F",X"1F",X"0F",X"1F",X"3F",X"3F",X"3F",X"70",X"78",X"38",X"20",X"23",X"37",X"1F",X"1F",
		X"1F",X"19",X"18",X"08",X"0E",X"0F",X"0F",X"06",X"1F",X"1F",X"0F",X"07",X"03",X"07",X"07",X"0F",
		X"E1",X"C3",X"47",X"6F",X"7F",X"3F",X"1F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"F0",
		X"23",X"20",X"20",X"38",X"3C",X"3C",X"18",X"00",X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"37",
		X"47",X"6F",X"3F",X"3F",X"1F",X"1F",X"1F",X"0F",X"00",X"00",X"30",X"78",X"78",X"70",X"40",X"41",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"80",X"C0",X"71",X"10",X"E1",X"C0",X"80",X"00",X"80",X"C0",X"71",X"31",
		X"FF",X"FF",X"F9",X"F9",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F3",X"FF",X"7F",X"1F",X"0F",X"07",X"00",X"00",X"FF",X"E7",X"E7",X"FF",X"FF",X"FF",X"FF",X"F3",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"08",X"1C",X"3E",X"7E",X"7C",X"7F",
		X"FF",X"FF",X"3E",X"3F",X"3F",X"1F",X"0F",X"07",X"FF",X"FF",X"FF",X"FF",X"FC",X"FC",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FC",X"FC",X"FF",X"FF",X"07",X"0F",X"1F",X"3F",X"3F",X"3E",X"7F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F1",X"00",X"00",X"00",X"00",X"00",X"F1",X"10",X"C1",X"00",X"00",X"00",X"00",X"00",X"F1",X"F1",
		X"FF",X"FF",X"FF",X"C3",X"C3",X"C1",X"01",X"01",X"00",X"00",X"C0",X"E0",X"FC",X"FE",X"FF",X"FF",
		X"F7",X"F7",X"F9",X"80",X"80",X"00",X"00",X"00",X"EF",X"EF",X"F7",X"FB",X"FB",X"FB",X"F7",X"F7",
		X"FF",X"FF",X"F7",X"F7",X"F7",X"F7",X"EF",X"EF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"F3",X"01",X"00",X"00",X"00",X"00",X"00",X"F7",X"F7",X"F7",X"F3",X"FB",X"FB",X"FB",X"FB",
		X"FB",X"FB",X"FB",X"FB",X"F3",X"F7",X"F7",X"F7",X"00",X"00",X"00",X"00",X"00",X"01",X"F3",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"F1",X"10",X"F0",X"00",X"00",X"00",X"00",X"00",X"F1",X"F0",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"E0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"70",X"F8",X"F8",X"F8",
		X"F8",X"F8",X"F8",X"F8",X"70",X"00",X"00",X"00",X"E0",X"E0",X"E0",X"E0",X"F0",X"F8",X"F8",X"F8",
		X"F8",X"F8",X"F8",X"F0",X"E0",X"E0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"70",X"F8",X"F8",X"F8",
		X"F8",X"F0",X"C0",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C8",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"C8",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"C0",X"F0",X"F8",
		X"8F",X"87",X"E3",X"F0",X"F0",X"60",X"00",X"00",X"0F",X"1F",X"3F",X"3F",X"7F",X"FF",X"9F",X"9F",
		X"9F",X"9F",X"FF",X"7F",X"3F",X"3F",X"1F",X"0F",X"00",X"00",X"60",X"F0",X"F0",X"E3",X"87",X"8F",
		X"70",X"78",X"78",X"30",X"00",X"00",X"00",X"00",X"3E",X"3F",X"7C",X"5D",X"CE",X"87",X"C0",X"40",
		X"5F",X"7F",X"3F",X"3F",X"3E",X"3D",X"1D",X"3D",X"03",X"07",X"1F",X"33",X"60",X"C7",X"8F",X"DF",
		X"30",X"78",X"78",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"07",X"03",X"00",X"00",X"00",X"00",
		X"3C",X"3C",X"18",X"00",X"00",X"00",X"00",X"00",X"73",X"EB",X"AB",X"A8",X"90",X"CB",X"67",X"3B",
		X"3F",X"3C",X"3B",X"17",X"36",X"75",X"7B",X"7F",X"03",X"06",X"04",X"05",X"07",X"0F",X"1F",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"03",X"01",X"00",X"00",X"FF",X"FE",X"FE",X"CF",X"CE",X"FE",X"FE",X"FF",
		X"FF",X"FE",X"FE",X"CE",X"CF",X"FE",X"FE",X"FF",X"00",X"00",X"01",X"03",X"FF",X"FF",X"FF",X"FF",
		X"1F",X"1F",X"05",X"04",X"04",X"00",X"00",X"00",X"3E",X"FF",X"3E",X"CF",X"CF",X"1F",X"FF",X"1F",
		X"81",X"81",X"81",X"0B",X"EF",X"E7",X"E7",X"DF",X"00",X"80",X"80",X"1F",X"FF",X"FF",X"E3",X"C1",
		X"1F",X"1F",X"05",X"04",X"04",X"00",X"00",X"00",X"30",X"01",X"30",X"09",X"0D",X"1F",X"07",X"7F",
		X"00",X"00",X"00",X"08",X"0C",X"04",X"04",X"18",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"1F",X"0F",X"3F",X"1F",X"3F",X"3F",X"00",X"F1",X"E0",X"E0",X"FF",X"C6",X"CE",X"DE",X"9F",
		X"07",X"07",X"BF",X"7F",X"3F",X"38",X"F8",X"FC",X"FD",X"03",X"7F",X"FF",X"FF",X"FF",X"8F",X"07",
		X"C3",X"F3",X"FC",X"F8",X"F0",X"E0",X"00",X"00",X"03",X"01",X"07",X"81",X"01",X"01",X"03",X"03",
		X"03",X"03",X"01",X"01",X"81",X"07",X"01",X"03",X"00",X"00",X"E0",X"F0",X"F8",X"FC",X"F3",X"C3",
		X"FE",X"FE",X"3F",X"3E",X"0E",X"00",X"00",X"00",X"3F",X"9F",X"01",X"80",X"E0",X"E0",X"F9",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FE",X"3E",X"3E",X"0E",X"00",X"00",X"00",X"1E",X"9E",X"00",X"80",X"E0",X"E0",X"F8",X"FE",
		X"00",X"70",X"FC",X"FE",X"FE",X"7E",X"3E",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"FC",X"EC",X"E7",X"E1",X"E0",X"E0",X"00",X"3F",X"3F",X"3F",X"13",X"03",X"03",X"47",X"E7",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"80",X"C0",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",
		X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"04",X"3C",X"F0",X"C0",X"00",X"00",X"00",X"00",X"FE",X"FC",X"FC",X"FE",X"FE",X"F8",X"C0",X"00",
		X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"00",X"00",X"00",X"C0",X"F0",X"F8",X"FC",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"7C",X"E0",X"00",X"00",X"00",X"00",X"FE",X"FC",X"FC",X"FC",X"FC",X"F8",X"E0",X"00",
		X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"C0",X"F0",X"F8",X"FC",
		X"3C",X"3C",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"03",X"00",X"00",X"03",X"03",X"18",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"06",X"0F",X"0F",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"02",X"02",X"02",
		X"3C",X"3E",X"1B",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",
		X"00",X"30",X"78",X"7C",X"36",X"03",X"00",X"00",X"01",X"03",X"03",X"03",X"01",X"00",X"00",X"00",
		X"03",X"03",X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"08",X"0C",X"04",X"06",X"03",X"00",X"00",X"00",X"03",X"03",X"01",X"01",X"18",X"3C",X"3C",X"18",
		X"60",X"30",X"18",X"08",X"E0",X"38",X"04",X"76",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"1F",X"0F",X"3F",X"1F",X"3F",X"3F",X"00",X"01",X"00",X"00",X"9F",X"86",X"8E",X"1E",X"1F",
		X"00",X"00",X"31",X"71",X"31",X"20",X"C0",X"0C",X"01",X"03",X"03",X"01",X"00",X"00",X"00",X"00",
		X"01",X"03",X"03",X"07",X"07",X"03",X"01",X"00",X"1F",X"3F",X"7F",X"FF",X"7F",X"4B",X"01",X"01",
		X"01",X"01",X"4B",X"FF",X"FF",X"7F",X"3F",X"1F",X"00",X"01",X"03",X"07",X"07",X"03",X"03",X"01",
		X"3F",X"3F",X"1F",X"1F",X"0E",X"FC",X"00",X"00",X"80",X"A0",X"A0",X"FF",X"E7",X"8C",X"7F",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"F1",X"00",X"00",X"00",X"3F",X"3F",X"7F",X"FF",X"FF",
		X"7F",X"7F",X"3F",X"1F",X"8F",X"FE",X"00",X"00",X"E3",X"E3",X"FF",X"FF",X"FF",X"07",X"F3",X"7F",
		X"3F",X"3F",X"3F",X"7F",X"33",X"31",X"71",X"E3",X"00",X"00",X"00",X"3F",X"1F",X"1F",X"1F",X"1F",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"00",X"3C",X"38",X"38",X"10",X"00",X"00",X"40",X"E0",
		X"00",X"F0",X"FC",X"FE",X"FE",X"FE",X"7E",X"FC",X"80",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FD",X"F8",X"F0",X"00",X"FF",X"FF",X"E7",X"E7",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"E7",X"E7",X"FF",X"FF",X"00",X"00",X"F0",X"F8",X"FD",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"0C",X"07",X"0F",X"8F",X"9F",X"FF",X"E7",X"0F",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"1F",X"0F",X"00",X"00",X"00",X"03",X"C7",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"0C",X"07",X"FF",X"FF",X"FF",X"FF",X"07",X"F3",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"C1",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FC",X"FC",X"FC",X"7C",X"78",X"30",X"00",X"0E",X"8E",X"8E",X"1E",X"0C",X"0C",X"8C",X"DC",
		X"DC",X"8C",X"0C",X"0C",X"1E",X"8E",X"8E",X"0E",X"00",X"30",X"78",X"7C",X"FC",X"FC",X"FC",X"FC",
		X"C0",X"80",X"80",X"C0",X"82",X"0F",X"1F",X"F6",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",X"F8",
		X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"F0",X"F8",X"F8",X"FC",X"FC",
		X"C0",X"80",X"80",X"E0",X"D0",X"BC",X"3C",X"F8",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",X"F8",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FC",X"FC",X"FE",X"FE",X"FE",
		X"47",X"63",X"21",X"3C",X"1E",X"1E",X"0C",X"00",X"07",X"0F",X"1F",X"1F",X"3F",X"7F",X"4F",X"4F",
		X"67",X"3F",X"1F",X"1F",X"1F",X"1F",X"0F",X"07",X"18",X"3C",X"3C",X"78",X"C0",X"80",X"81",X"C3",
		X"70",X"78",X"78",X"30",X"00",X"00",X"00",X"00",X"3F",X"3F",X"7F",X"FF",X"9F",X"8F",X"86",X"C0",
		X"1F",X"1F",X"1F",X"0F",X"1F",X"3F",X"3F",X"3F",X"70",X"78",X"38",X"20",X"23",X"37",X"1F",X"1F",
		X"23",X"20",X"20",X"38",X"3C",X"3C",X"18",X"00",X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"37",
		X"47",X"6F",X"3F",X"3F",X"1F",X"1F",X"1F",X"0F",X"00",X"00",X"30",X"78",X"78",X"70",X"40",X"41",
		X"F1",X"F0",X"60",X"00",X"00",X"00",X"00",X"00",X"3F",X"3F",X"7F",X"FF",X"DF",X"CF",X"8F",X"E7",
		X"1F",X"1F",X"1F",X"0F",X"1F",X"3F",X"3F",X"3F",X"06",X"0F",X"0F",X"16",X"30",X"30",X"3B",X"3F",
		X"FF",X"FF",X"FF",X"7F",X"03",X"01",X"00",X"00",X"FF",X"FF",X"F9",X"F9",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FF",X"F9",X"F9",X"FF",X"FF",X"FF",X"FF",X"07",X"0F",X"0F",X"1F",X"1F",X"7F",X"FE",X"FE",
		X"11",X"00",X"00",X"00",X"80",X"C0",X"71",X"10",X"E1",X"C0",X"80",X"00",X"80",X"C0",X"71",X"31",
		X"F3",X"F3",X"FF",X"FF",X"FF",X"FF",X"FF",X"E7",X"00",X"00",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"3E",X"3F",X"3F",X"1F",X"0F",X"07",X"FF",X"FF",X"FC",X"FC",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FC",X"FC",X"FF",X"FF",X"FF",X"FF",X"07",X"0F",X"1F",X"3F",X"3F",X"3E",X"7F",X"FF",
		X"FF",X"7F",X"7F",X"7F",X"7F",X"3E",X"1C",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F3",X"FF",X"FF",X"FF",X"F3",X"F3",X"FF",X"FF",X"00",X"0F",X"1F",X"3F",X"3F",X"FF",X"FF",X"F3",
		X"F0",X"FD",X"FF",X"FC",X"F8",X"E0",X"00",X"00",X"F1",X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",X"E0",
		X"00",X"40",X"40",X"C1",X"F0",X"E0",X"E0",X"F1",X"00",X"80",X"C0",X"C0",X"9C",X"0F",X"0F",X"01",
		X"F1",X"00",X"00",X"00",X"00",X"00",X"F1",X"10",X"C1",X"00",X"00",X"00",X"00",X"00",X"F1",X"F1",
		X"FF",X"FF",X"FF",X"C3",X"C3",X"C1",X"01",X"01",X"00",X"00",X"C0",X"E0",X"FC",X"FE",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"0F",X"00",X"00",X"00",X"00",X"F7",X"FB",X"FB",X"FB",X"FB",X"FF",X"FF",X"FF",
		X"F7",X"F7",X"FB",X"FB",X"FB",X"F7",X"EF",X"EF",X"00",X"80",X"80",X"C0",X"C0",X"F1",X"FB",X"F7",
		X"F8",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"F8",X"78",X"78",X"78",X"78",X"F8",
		X"F8",X"78",X"78",X"F8",X"78",X"F8",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"F8",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"F1",X"10",X"F0",X"00",X"00",X"00",X"00",X"00",X"F1",X"F0",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"E0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"70",X"F8",X"F8",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"F8",X"F8",X"F8",X"F0",X"00",X"00",X"00",X"E0",X"E0",X"E0",X"E0",X"E0",X"F0",X"F8",X"F8",
		X"F8",X"F8",X"F8",X"F8",X"F0",X"E0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"70",X"F8",X"F8",X"F8");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
