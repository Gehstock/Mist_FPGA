library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity BLACKHOLE_ROM_PGM_0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of BLACKHOLE_ROM_PGM_0 is
	type rom is array(0 to  12287) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"AF",X"32",X"01",X"70",X"C3",X"50",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F5",X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",X"AF",X"32",
		X"01",X"70",X"21",X"00",X"42",X"11",X"00",X"58",X"01",X"80",X"00",X"ED",X"B0",X"CD",X"4F",X"01",
		X"3A",X"01",X"40",X"87",X"28",X"12",X"D6",X"02",X"5F",X"16",X"00",X"21",X"E3",X"00",X"19",X"5E",
		X"23",X"56",X"EB",X"11",X"98",X"00",X"D5",X"E9",X"CD",X"C4",X"26",X"CD",X"7F",X"01",X"21",X"07",
		X"40",X"35",X"3A",X"00",X"78",X"CD",X"CA",X"01",X"3A",X"00",X"60",X"32",X"05",X"40",X"3A",X"00",
		X"68",X"32",X"06",X"40",X"3A",X"00",X"40",X"87",X"28",X"1A",X"D6",X"02",X"5F",X"16",X"00",X"21",
		X"0B",X"01",X"19",X"5E",X"23",X"56",X"21",X"0C",X"00",X"39",X"73",X"23",X"72",X"AF",X"32",X"00",
		X"40",X"32",X"01",X"40",X"3E",X"FF",X"32",X"01",X"70",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",
		X"F1",X"ED",X"45",X"46",X"19",X"54",X"19",X"58",X"19",X"53",X"1E",X"67",X"1E",X"7B",X"1E",X"00",
		X"09",X"00",X"09",X"8C",X"20",X"9F",X"20",X"B2",X"20",X"27",X"10",X"49",X"10",X"46",X"10",X"53",
		X"10",X"96",X"18",X"A6",X"18",X"B0",X"18",X"00",X"09",X"C3",X"18",X"C7",X"18",X"00",X"09",X"CC",
		X"1B",X"4A",X"1C",X"9B",X"1C",X"18",X"1D",X"AD",X"1D",X"4E",X"1F",X"00",X"09",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"BC",X"0F",X"00",X"00",X"00",X"00",X"D7",
		X"1F",X"5E",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E6",X"11",X"00",X"00",X"25",
		X"14",X"00",X"00",X"00",X"00",X"49",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"B2",X"08",X"0E",
		X"06",X"21",X"FA",X"40",X"11",X"A1",X"53",X"CD",X"3C",X"07",X"21",X"40",X"41",X"11",X"41",X"52",
		X"CD",X"3C",X"07",X"3A",X"08",X"40",X"3D",X"CA",X"73",X"01",X"21",X"3A",X"41",X"11",X"E1",X"50",
		X"CD",X"3C",X"07",X"0E",X"02",X"21",X"0A",X"40",X"11",X"DF",X"52",X"CD",X"3C",X"07",X"C9",X"3A",
		X"00",X"60",X"E6",X"01",X"57",X"3A",X"02",X"40",X"CB",X"27",X"B2",X"E6",X"0F",X"32",X"02",X"40",
		X"FE",X"0C",X"C0",X"3A",X"00",X"68",X"E6",X"C0",X"07",X"07",X"FE",X"03",X"57",X"3A",X"03",X"60",
		X"7A",X"CA",X"BE",X"01",X"3C",X"21",X"03",X"40",X"86",X"27",X"57",X"77",X"AF",X"ED",X"6F",X"C6",
		X"58",X"32",X"0A",X"40",X"AF",X"ED",X"6F",X"C6",X"58",X"32",X"0B",X"40",X"72",X"C9",X"21",X"6F",
		X"40",X"34",X"CB",X"46",X"3E",X"00",X"CA",X"A4",X"01",X"C9",X"21",X"04",X"40",X"3A",X"00",X"40",
		X"A7",X"28",X"08",X"36",X"59",X"FE",X"06",X"38",X"02",X"36",X"4E",X"7E",X"FE",X"59",X"28",X"1A",
		X"21",X"00",X"40",X"7E",X"FE",X"22",X"28",X"69",X"3A",X"00",X"40",X"D6",X"01",X"D8",X"5F",X"16",
		X"00",X"21",X"67",X"02",X"19",X"7E",X"32",X"00",X"40",X"C9",X"3A",X"03",X"40",X"A7",X"28",X"E8",
		X"3E",X"4E",X"77",X"3E",X"06",X"32",X"00",X"40",X"C9",X"3A",X"06",X"40",X"2F",X"57",X"3A",X"00",
		X"68",X"A2",X"E6",X"03",X"C8",X"57",X"3D",X"28",X"05",X"3A",X"03",X"40",X"3D",X"C8",X"D5",X"AF",
		X"06",X"03",X"21",X"F7",X"40",X"11",X"37",X"41",X"77",X"12",X"23",X"13",X"10",X"FA",X"3E",X"58",
		X"06",X"06",X"21",X"FA",X"40",X"11",X"3A",X"41",X"77",X"12",X"23",X"13",X"10",X"FA",X"D1",X"7A",
		X"32",X"08",X"40",X"21",X"03",X"40",X"7E",X"92",X"27",X"CD",X"AA",X"01",X"21",X"00",X"40",X"18",
		X"97",X"3A",X"02",X"40",X"FE",X"0C",X"C2",X"09",X"02",X"3A",X"6F",X"40",X"E6",X"01",X"C2",X"09",
		X"02",X"3E",X"06",X"32",X"00",X"40",X"C9",X"03",X"03",X"04",X"05",X"01",X"22",X"08",X"09",X"0A",
		X"0B",X"1E",X"0E",X"14",X"10",X"19",X"1E",X"19",X"14",X"07",X"1E",X"01",X"3F",X"3F",X"3F",X"13",
		X"1B",X"14",X"13",X"1E",X"07",X"07",X"0E",X"19",X"07",X"3A",X"0F",X"40",X"3C",X"32",X"0F",X"40",
		X"CB",X"47",X"C8",X"0F",X"E6",X"07",X"57",X"0E",X"07",X"21",X"10",X"40",X"06",X"00",X"09",X"5E",
		X"AF",X"83",X"28",X"1B",X"CB",X"5B",X"28",X"0B",X"E6",X"07",X"5F",X"7A",X"BB",X"DC",X"C4",X"02",
		X"CD",X"C4",X"02",X"7B",X"E6",X"07",X"5F",X"7A",X"BB",X"DC",X"C4",X"02",X"CD",X"C4",X"02",X"0D",
		X"F2",X"99",X"02",X"C9",X"D5",X"21",X"28",X"40",X"09",X"7E",X"3C",X"E6",X"07",X"77",X"57",X"21",
		X"18",X"40",X"09",X"5E",X"7B",X"E6",X"C0",X"28",X"25",X"AF",X"82",X"28",X"1F",X"CB",X"47",X"28",
		X"1D",X"7B",X"E6",X"C0",X"FE",X"40",X"28",X"3A",X"FE",X"80",X"28",X"12",X"7B",X"E6",X"07",X"CB",
		X"57",X"C4",X"26",X"03",X"CD",X"63",X"21",X"83",X"5F",X"CD",X"4D",X"21",X"D1",X"C9",X"7B",X"E6",
		X"07",X"CB",X"57",X"C4",X"26",X"03",X"6F",X"7B",X"E6",X"38",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",
		X"CB",X"57",X"C4",X"26",X"03",X"CD",X"63",X"21",X"82",X"57",X"7D",X"83",X"5F",X"CD",X"4D",X"21",
		X"D1",X"C9",X"2E",X"00",X"18",X"E1",X"3E",X"FF",X"C9",X"06",X"07",X"21",X"20",X"40",X"58",X"16",
		X"00",X"19",X"7E",X"6F",X"CD",X"BC",X"21",X"30",X"11",X"7B",X"85",X"5F",X"CD",X"86",X"21",X"7B",
		X"FE",X"10",X"DC",X"B0",X"06",X"FE",X"F9",X"D4",X"B0",X"06",X"05",X"F2",X"2B",X"03",X"C9",X"3A",
		X"09",X"40",X"A7",X"CA",X"6C",X"03",X"3A",X"00",X"70",X"E6",X"02",X"C2",X"6C",X"03",X"3A",X"06",
		X"40",X"2F",X"21",X"00",X"68",X"A6",X"E6",X"10",X"C8",X"C3",X"77",X"03",X"3A",X"05",X"40",X"2F",
		X"21",X"00",X"60",X"A6",X"E6",X"10",X"C8",X"06",X"06",X"CD",X"BC",X"21",X"7B",X"FE",X"A0",X"D2",
		X"93",X"03",X"05",X"F2",X"79",X"03",X"06",X"06",X"CD",X"BC",X"21",X"D2",X"A0",X"03",X"05",X"F2",
		X"88",X"03",X"C9",X"21",X"20",X"40",X"16",X"00",X"58",X"19",X"7E",X"A7",X"F2",X"82",X"03",X"C9",
		X"3A",X"09",X"40",X"5F",X"16",X"00",X"21",X"F2",X"40",X"19",X"7E",X"3D",X"C2",X"C9",X"03",X"3A",
		X"38",X"42",X"C6",X"7F",X"57",X"1E",X"D4",X"CD",X"86",X"21",X"3E",X"01",X"32",X"30",X"40",X"21",
		X"20",X"40",X"58",X"16",X"00",X"19",X"36",X"FD",X"C9",X"3A",X"58",X"42",X"C6",X"08",X"C3",X"B4",
		X"03",X"3A",X"09",X"40",X"A7",X"CA",X"22",X"04",X"3A",X"00",X"70",X"E6",X"02",X"C2",X"22",X"04",
		X"3A",X"00",X"68",X"E6",X"0C",X"C8",X"CB",X"57",X"CA",X"2B",X"04",X"3E",X"FF",X"21",X"09",X"40",
		X"5E",X"16",X"00",X"21",X"F2",X"40",X"19",X"56",X"15",X"CA",X"0D",X"04",X"21",X"58",X"42",X"11",
		X"04",X"00",X"86",X"FE",X"10",X"C8",X"FE",X"E0",X"C8",X"77",X"19",X"77",X"C9",X"21",X"34",X"42",
		X"86",X"FE",X"6A",X"C8",X"FE",X"96",X"C8",X"11",X"02",X"00",X"77",X"19",X"77",X"19",X"77",X"19",
		X"77",X"C9",X"3A",X"00",X"60",X"E6",X"0C",X"C8",X"C3",X"E6",X"03",X"3E",X"01",X"C3",X"ED",X"03",
		X"3A",X"09",X"40",X"4F",X"06",X"00",X"21",X"C0",X"40",X"09",X"3A",X"73",X"40",X"3C",X"E6",X"03",
		X"32",X"73",X"40",X"C6",X"26",X"4F",X"09",X"11",X"FC",X"FF",X"06",X"04",X"7E",X"E5",X"CD",X"00",
		X"09",X"FE",X"FF",X"C4",X"39",X"08",X"CC",X"26",X"08",X"E1",X"19",X"79",X"90",X"4F",X"F2",X"4C",
		X"04",X"C9",X"0E",X"05",X"21",X"C0",X"40",X"3A",X"09",X"40",X"85",X"6F",X"5F",X"3E",X"00",X"8C",
		X"67",X"57",X"23",X"23",X"E5",X"7E",X"23",X"46",X"6F",X"60",X"B0",X"CA",X"87",X"04",X"CB",X"41",
		X"20",X"31",X"3E",X"DC",X"CD",X"39",X"08",X"E1",X"1A",X"BE",X"C2",X"9F",X"04",X"13",X"23",X"1A",
		X"BE",X"C2",X"B8",X"04",X"13",X"13",X"13",X"23",X"23",X"23",X"0D",X"F2",X"74",X"04",X"C9",X"E5",
		X"1A",X"6F",X"13",X"1A",X"67",X"CD",X"26",X"08",X"1B",X"E1",X"7E",X"12",X"23",X"13",X"7E",X"12",
		X"C3",X"94",X"04",X"3E",X"04",X"C3",X"84",X"04",X"1B",X"2B",X"C3",X"9F",X"04",X"21",X"7A",X"40",
		X"34",X"CA",X"05",X"05",X"21",X"7A",X"40",X"7E",X"E6",X"03",X"C6",X"A1",X"4F",X"21",X"50",X"41",
		X"06",X"00",X"09",X"EB",X"21",X"F0",X"21",X"09",X"09",X"7E",X"23",X"46",X"6F",X"60",X"E6",X"1F",
		X"47",X"3A",X"0D",X"40",X"80",X"FE",X"1E",X"D2",X"83",X"05",X"3A",X"0D",X"40",X"85",X"6F",X"3A",
		X"09",X"40",X"A7",X"C2",X"A4",X"05",X"1A",X"E6",X"0F",X"3C",X"ED",X"44",X"77",X"79",X"D6",X"04",
		X"4F",X"D2",X"CD",X"04",X"C9",X"11",X"0D",X"40",X"1A",X"C6",X"A7",X"6F",X"26",X"53",X"3E",X"FF",
		X"01",X"E0",X"FF",X"77",X"09",X"77",X"09",X"77",X"09",X"77",X"09",X"77",X"23",X"09",X"77",X"09",
		X"77",X"09",X"77",X"23",X"09",X"77",X"09",X"77",X"09",X"77",X"23",X"09",X"77",X"09",X"77",X"23",
		X"09",X"77",X"09",X"77",X"2B",X"09",X"77",X"09",X"77",X"2B",X"09",X"77",X"09",X"77",X"09",X"77",
		X"2B",X"09",X"77",X"09",X"77",X"09",X"77",X"2B",X"09",X"77",X"09",X"77",X"09",X"77",X"09",X"77",
		X"09",X"77",X"EB",X"34",X"21",X"71",X"05",X"11",X"60",X"53",X"0E",X"10",X"CD",X"3C",X"07",X"21",
		X"81",X"05",X"11",X"A0",X"50",X"0E",X"02",X"3A",X"08",X"40",X"3D",X"C4",X"3C",X"07",X"C3",X"C4",
		X"04",X"59",X"6B",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"66",X"67",X"FF",X"6D",X"63",X"6A",X"6C",
		X"65",X"5A",X"6B",X"3A",X"09",X"40",X"A7",X"C2",X"97",X"05",X"1A",X"E6",X"0F",X"C4",X"B5",X"05",
		X"1A",X"E6",X"F0",X"12",X"C3",X"FD",X"04",X"1A",X"E6",X"F0",X"C4",X"BA",X"05",X"1A",X"E6",X"0F",
		X"12",X"C3",X"FD",X"04",X"1A",X"E6",X"F0",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"3C",
		X"ED",X"44",X"C3",X"FC",X"04",X"21",X"C0",X"40",X"35",X"C9",X"21",X"00",X"41",X"35",X"C9",X"21",
		X"7B",X"40",X"34",X"CB",X"46",X"C8",X"3A",X"0C",X"40",X"FE",X"52",X"CA",X"E5",X"05",X"21",X"06",
		X"42",X"01",X"02",X"00",X"35",X"09",X"35",X"09",X"35",X"09",X"35",X"7E",X"FE",X"A0",X"C0",X"3E",
		X"52",X"32",X"0C",X"40",X"C9",X"21",X"06",X"42",X"01",X"02",X"00",X"34",X"09",X"34",X"09",X"34",
		X"09",X"34",X"7E",X"FE",X"60",X"C0",X"3E",X"4C",X"32",X"0C",X"40",X"C9",X"3A",X"09",X"40",X"4F",
		X"06",X"00",X"1E",X"5D",X"21",X"FC",X"40",X"3A",X"00",X"70",X"E6",X"01",X"CA",X"12",X"06",X"1E",
		X"59",X"2B",X"09",X"7B",X"BE",X"C0",X"21",X"7C",X"40",X"59",X"79",X"07",X"07",X"4F",X"09",X"7E",
		X"FE",X"4E",X"C8",X"3E",X"01",X"32",X"48",X"40",X"36",X"4E",X"21",X"F0",X"40",X"4B",X"09",X"34",
		X"C3",X"55",X"07",X"3A",X"0E",X"40",X"3D",X"FA",X"43",X"06",X"4F",X"06",X"00",X"21",X"92",X"40",
		X"09",X"36",X"21",X"0E",X"02",X"21",X"92",X"40",X"06",X"00",X"09",X"7E",X"A7",X"CA",X"7A",X"06",
		X"35",X"7E",X"16",X"0C",X"FE",X"20",X"28",X"13",X"FE",X"10",X"28",X"0F",X"16",X"10",X"FE",X"18",
		X"28",X"09",X"FE",X"08",X"28",X"05",X"A7",X"28",X"1A",X"18",X"0F",X"21",X"85",X"52",X"7A",X"11",
		X"C0",X"FF",X"41",X"04",X"19",X"10",X"FD",X"CD",X"39",X"08",X"0D",X"F2",X"45",X"06",X"AF",X"32",
		X"0E",X"40",X"C9",X"79",X"3D",X"3E",X"2E",X"21",X"05",X"52",X"CC",X"39",X"08",X"28",X"EB",X"79",
		X"A7",X"3E",X"32",X"21",X"25",X"52",X"28",X"05",X"3E",X"2C",X"21",X"C5",X"51",X"77",X"23",X"3C",
		X"77",X"79",X"A7",X"2E",X"45",X"28",X"02",X"2E",X"A5",X"3E",X"FF",X"77",X"23",X"77",X"18",X"CA",
		X"D5",X"11",X"00",X"00",X"CD",X"86",X"21",X"D1",X"C9",X"F5",X"C5",X"E5",X"21",X"02",X"50",X"3E",
		X"FF",X"0E",X"20",X"06",X"1D",X"77",X"23",X"10",X"FC",X"23",X"23",X"23",X"0D",X"C2",X"C3",X"06",
		X"E1",X"C1",X"F1",X"C9",X"F5",X"C5",X"D5",X"E5",X"3A",X"09",X"40",X"4F",X"06",X"00",X"21",X"F9",
		X"40",X"09",X"7E",X"83",X"27",X"77",X"2B",X"7E",X"8A",X"27",X"77",X"2B",X"7E",X"CE",X"00",X"27",
		X"77",X"11",X"FA",X"40",X"EB",X"09",X"EB",X"06",X"03",X"4E",X"AF",X"ED",X"6F",X"C6",X"58",X"12",
		X"13",X"AF",X"ED",X"6F",X"C6",X"58",X"12",X"13",X"71",X"23",X"10",X"ED",X"2B",X"D5",X"11",X"48",
		X"41",X"EB",X"1A",X"96",X"27",X"1B",X"2B",X"1A",X"9E",X"27",X"1B",X"2B",X"1A",X"9E",X"27",X"DA",
		X"36",X"07",X"01",X"03",X"00",X"EB",X"ED",X"B0",X"D1",X"1B",X"21",X"45",X"41",X"EB",X"01",X"06",
		X"00",X"ED",X"B8",X"C3",X"37",X"07",X"E1",X"E1",X"D1",X"C1",X"F1",X"C9",X"F5",X"C5",X"D5",X"E5",
		X"06",X"00",X"ED",X"A0",X"E2",X"50",X"07",X"7B",X"D6",X"21",X"5F",X"7A",X"98",X"57",X"18",X"F2",
		X"E1",X"D1",X"C1",X"F1",X"C9",X"3A",X"09",X"40",X"4F",X"06",X"00",X"21",X"F0",X"40",X"09",X"56",
		X"21",X"F2",X"40",X"09",X"7E",X"3D",X"C2",X"D2",X"07",X"15",X"CA",X"8A",X"07",X"15",X"CA",X"9F",
		X"07",X"15",X"CA",X"B4",X"07",X"3E",X"E8",X"21",X"1A",X"52",X"CD",X"39",X"08",X"3E",X"EC",X"21",
		X"1C",X"52",X"CD",X"39",X"08",X"16",X"02",X"C3",X"C6",X"07",X"3E",X"E0",X"21",X"1A",X"52",X"CD",
		X"39",X"08",X"3E",X"E4",X"21",X"1C",X"52",X"CD",X"39",X"08",X"16",X"01",X"C3",X"C6",X"07",X"3E",
		X"3C",X"21",X"1A",X"52",X"CD",X"39",X"08",X"3E",X"40",X"21",X"09",X"02",X"CD",X"39",X"08",X"16",
		X"02",X"C3",X"C6",X"07",X"3E",X"34",X"21",X"1A",X"52",X"CD",X"39",X"08",X"3E",X"38",X"21",X"1C",
		X"52",X"CD",X"39",X"08",X"16",X"07",X"06",X"1D",X"CD",X"ED",X"20",X"05",X"78",X"FE",X"19",X"20",
		X"F7",X"C9",X"15",X"CA",X"E4",X"07",X"15",X"CA",X"EA",X"07",X"15",X"CA",X"F0",X"07",X"01",X"02",
		X"3A",X"C3",X"F3",X"07",X"01",X"01",X"38",X"C3",X"F3",X"07",X"01",X"02",X"0F",X"C3",X"F3",X"07",
		X"01",X"07",X"0D",X"21",X"59",X"42",X"70",X"23",X"71",X"04",X"21",X"5D",X"42",X"70",X"23",X"71",
		X"23",X"7E",X"FE",X"E0",X"C2",X"10",X"08",X"3A",X"5B",X"42",X"FE",X"D0",X"C2",X"10",X"08",X"C9",
		X"3A",X"34",X"42",X"C6",X"78",X"32",X"58",X"42",X"32",X"5C",X"42",X"3E",X"D0",X"32",X"5B",X"42",
		X"3E",X"E0",X"32",X"5F",X"42",X"C9",X"F5",X"D5",X"E5",X"3E",X"FF",X"11",X"E0",X"FF",X"77",X"23",
		X"77",X"19",X"77",X"2B",X"77",X"E1",X"D1",X"F1",X"C9",X"F5",X"D5",X"E5",X"C6",X"02",X"77",X"3C",
		X"23",X"77",X"D6",X"02",X"11",X"E0",X"FF",X"19",X"77",X"3D",X"2B",X"77",X"E1",X"D1",X"F1",X"C9",
		X"01",X"04",X"00",X"21",X"00",X"40",X"77",X"23",X"10",X"FC",X"0D",X"20",X"F9",X"F9",X"06",X"80",
		X"21",X"00",X"58",X"77",X"23",X"10",X"FC",X"16",X"58",X"21",X"FA",X"40",X"3E",X"03",X"06",X"06",
		X"72",X"23",X"10",X"FC",X"3D",X"21",X"40",X"41",X"FE",X"02",X"28",X"F2",X"21",X"3A",X"41",X"FE",
		X"01",X"28",X"EB",X"21",X"0A",X"40",X"72",X"23",X"72",X"3E",X"FF",X"01",X"04",X"00",X"21",X"00",
		X"50",X"77",X"23",X"10",X"FC",X"0D",X"20",X"F9",X"ED",X"5F",X"32",X"91",X"40",X"AF",X"32",X"06",
		X"70",X"32",X"07",X"70",X"3E",X"FF",X"32",X"01",X"70",X"3E",X"05",X"32",X"00",X"40",X"00",X"18",
		X"FD",X"C9",X"3E",X"22",X"32",X"00",X"40",X"C3",X"B7",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CD",X"B9",X"06",X"AF",X"32",X"0D",X"40",X"21",X"C1",X"40",X"3A",X"09",X"40",X"06",X"00",X"4F",
		X"09",X"AF",X"06",X"0F",X"77",X"23",X"10",X"FC",X"3A",X"E3",X"51",X"FE",X"24",X"28",X"27",X"21",
		X"E3",X"51",X"3E",X"24",X"0E",X"02",X"06",X"02",X"CD",X"39",X"08",X"C6",X"08",X"23",X"23",X"10",
		X"F7",X"21",X"23",X"52",X"3E",X"28",X"0D",X"20",X"ED",X"21",X"06",X"42",X"06",X"04",X"36",X"00",
		X"23",X"36",X"02",X"23",X"10",X"F8",X"16",X"06",X"06",X"05",X"3E",X"1E",X"CD",X"ED",X"20",X"16",
		X"00",X"CD",X"DC",X"20",X"16",X"06",X"04",X"B8",X"C2",X"4C",X"09",X"16",X"05",X"06",X"1E",X"CD",
		X"ED",X"20",X"3A",X"09",X"40",X"4F",X"06",X"00",X"21",X"F2",X"40",X"09",X"36",X"02",X"21",X"F4",
		X"40",X"09",X"7E",X"FE",X"4E",X"CA",X"4C",X"0A",X"36",X"4E",X"21",X"C0",X"40",X"09",X"36",X"9E",
		X"21",X"50",X"41",X"11",X"A6",X"09",X"CB",X"71",X"01",X"00",X"A6",X"C2",X"9A",X"09",X"ED",X"67",
		X"1A",X"ED",X"6F",X"23",X"13",X"10",X"F7",X"C3",X"4C",X"0A",X"ED",X"6F",X"1A",X"ED",X"67",X"23",
		X"13",X"10",X"F7",X"C3",X"4C",X"0A",X"06",X"06",X"06",X"06",X"06",X"06",X"00",X"06",X"06",X"06",
		X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",
		X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",
		X"00",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",
		X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",
		X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"00",X"00",X"05",X"05",X"05",X"05",X"05",X"05",X"00",
		X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",
		X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",
		X"05",X"05",X"05",X"00",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",
		X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",
		X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"00",X"00",X"06",X"00",X"CD",X"FF",
		X"20",X"30",X"01",X"02",X"48",X"04",X"CD",X"FF",X"20",X"44",X"81",X"02",X"48",X"04",X"CD",X"FF",
		X"20",X"70",X"01",X"02",X"70",X"04",X"CD",X"FF",X"20",X"84",X"81",X"02",X"70",X"04",X"CD",X"FF",
		X"20",X"B4",X"01",X"06",X"40",X"04",X"CD",X"FF",X"20",X"C8",X"81",X"06",X"40",X"0E",X"00",X"CD",
		X"63",X"21",X"CD",X"4C",X"0D",X"0E",X"02",X"CD",X"63",X"21",X"CD",X"4C",X"0D",X"0E",X"04",X"CD",
		X"63",X"21",X"CD",X"4C",X"0D",X"3A",X"09",X"40",X"4F",X"06",X"00",X"21",X"F3",X"40",X"09",X"7E",
		X"87",X"C6",X"10",X"21",X"10",X"40",X"06",X"06",X"77",X"23",X"10",X"FC",X"21",X"00",X"00",X"22",
		X"28",X"40",X"22",X"2A",X"40",X"22",X"2C",X"40",X"22",X"C2",X"40",X"22",X"C4",X"40",X"22",X"C6",
		X"40",X"22",X"92",X"40",X"AF",X"32",X"94",X"40",X"06",X"07",X"CD",X"B0",X"06",X"05",X"F2",X"CA",
		X"0A",X"3E",X"FF",X"32",X"00",X"68",X"32",X"01",X"68",X"CD",X"55",X"07",X"3E",X"0C",X"32",X"01",
		X"40",X"06",X"06",X"3A",X"09",X"40",X"6F",X"26",X"00",X"0E",X"05",X"CD",X"BC",X"21",X"D2",X"FB",
		X"0A",X"CD",X"8B",X"26",X"DA",X"02",X"0B",X"0D",X"F2",X"EB",X"0A",X"05",X"F2",X"E9",X"0A",X"C3",
		X"22",X"0B",X"CD",X"B0",X"06",X"C5",X"11",X"C2",X"40",X"79",X"E6",X"0E",X"4F",X"06",X"00",X"09",
		X"19",X"7E",X"A7",X"C2",X"1C",X"0B",X"36",X"8C",X"C1",X"C3",X"FB",X"0A",X"36",X"8B",X"C1",X"C3",
		X"FB",X"0A",X"06",X"06",X"CD",X"BC",X"21",X"38",X"07",X"05",X"F2",X"24",X"0B",X"C3",X"F3",X"0B",
		X"7B",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"21",X"0D",X"40",X"96",X"FE",X"07",X"DA",X"29",X"0B",
		X"5F",X"C5",X"7A",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"D6",X"02",X"47",X"80",X"80",X"4F",X"21",
		X"9F",X"0B",X"06",X"00",X"09",X"7E",X"23",X"56",X"C1",X"4F",X"7B",X"B9",X"DA",X"29",X"0B",X"7A",
		X"93",X"DA",X"29",X"0B",X"23",X"86",X"21",X"50",X"41",X"16",X"00",X"5F",X"19",X"3A",X"09",X"40",
		X"0E",X"F0",X"A7",X"20",X"02",X"0E",X"0F",X"7E",X"A1",X"CA",X"29",X"0B",X"79",X"2F",X"A6",X"77",
		X"CD",X"B0",X"06",X"11",X"10",X"00",X"CD",X"D4",X"06",X"3E",X"01",X"32",X"64",X"40",X"3A",X"09",
		X"40",X"21",X"C0",X"40",X"5F",X"16",X"00",X"19",X"35",X"CA",X"AE",X"0E",X"C3",X"29",X"0B",X"07",
		X"08",X"A4",X"07",X"09",X"A1",X"07",X"0A",X"9D",X"07",X"0B",X"98",X"07",X"0C",X"92",X"08",X"0D",
		X"8C",X"08",X"0E",X"85",X"08",X"0E",X"7E",X"09",X"0F",X"76",X"09",X"0F",X"6F",X"09",X"0F",X"68",
		X"0A",X"10",X"61",X"0A",X"10",X"5A",X"0B",X"10",X"53",X"0B",X"10",X"00",X"0A",X"10",X"07",X"0A",
		X"10",X"0E",X"09",X"0F",X"15",X"09",X"0F",X"1C",X"09",X"0F",X"23",X"08",X"0E",X"2B",X"08",X"0E",
		X"32",X"08",X"0D",X"39",X"07",X"0C",X"3F",X"07",X"0B",X"45",X"07",X"0A",X"4A",X"07",X"09",X"4E",
		X"07",X"08",X"51",X"06",X"06",X"CD",X"29",X"26",X"DA",X"02",X"0C",X"05",X"F2",X"F5",X"0B",X"C3",
		X"33",X"0C",X"CD",X"BC",X"21",X"CD",X"2E",X"24",X"7C",X"D6",X"50",X"85",X"16",X"02",X"FE",X"30",
		X"38",X"0D",X"16",X"01",X"FE",X"50",X"38",X"07",X"16",X"03",X"FE",X"E0",X"38",X"01",X"15",X"21",
		X"0E",X"40",X"72",X"CD",X"B0",X"06",X"3E",X"FF",X"32",X"7A",X"40",X"3E",X"01",X"32",X"50",X"40",
		X"C3",X"FB",X"0B",X"06",X"05",X"CD",X"EB",X"25",X"DA",X"B5",X"0D",X"05",X"F2",X"35",X"0C",X"3A",
		X"0D",X"40",X"FE",X"0A",X"DA",X"79",X"0C",X"0E",X"06",X"CD",X"63",X"21",X"7A",X"CB",X"3F",X"CB",
		X"3F",X"CB",X"3F",X"D6",X"02",X"4F",X"81",X"81",X"4F",X"16",X"03",X"06",X"00",X"21",X"9F",X"0B",
		X"09",X"7E",X"23",X"96",X"ED",X"44",X"3C",X"23",X"46",X"CD",X"FE",X"25",X"DA",X"8A",X"0E",X"04",
		X"3D",X"C2",X"69",X"0C",X"23",X"15",X"C2",X"61",X"0C",X"01",X"06",X"00",X"CD",X"63",X"21",X"EB",
		X"0E",X"05",X"CD",X"63",X"21",X"7B",X"D6",X"E6",X"DA",X"B0",X"0C",X"D6",X"05",X"DA",X"A6",X"0C",
		X"D6",X"10",X"DA",X"B0",X"0C",X"E5",X"21",X"C2",X"40",X"09",X"3A",X"09",X"40",X"16",X"00",X"5F",
		X"19",X"70",X"E1",X"C3",X"B0",X"0C",X"7A",X"94",X"DA",X"B0",X"0C",X"D6",X"1E",X"DA",X"B8",X"0C",
		X"0D",X"0D",X"F2",X"82",X"0C",X"C3",X"00",X"0D",X"E5",X"21",X"C1",X"40",X"09",X"3A",X"09",X"40",
		X"16",X"00",X"5F",X"19",X"EB",X"E1",X"1A",X"A7",X"CA",X"B0",X"0C",X"13",X"1A",X"A7",X"C2",X"B0",
		X"0C",X"3C",X"12",X"3E",X"05",X"B9",X"11",X"00",X"01",X"C4",X"EA",X"0C",X"11",X"00",X"03",X"CC",
		X"EA",X"0C",X"3E",X"01",X"32",X"5C",X"40",X"C3",X"B0",X"0C",X"F5",X"E5",X"CD",X"D4",X"06",X"21",
		X"C8",X"40",X"3A",X"09",X"40",X"5F",X"7A",X"C6",X"1E",X"16",X"00",X"19",X"77",X"E1",X"F1",X"C9",
		X"3A",X"09",X"40",X"4F",X"06",X"00",X"21",X"C0",X"40",X"09",X"7E",X"A7",X"CA",X"AE",X"0E",X"0E",
		X"00",X"CD",X"63",X"21",X"3E",X"50",X"BB",X"CA",X"37",X"0D",X"3E",X"51",X"BB",X"CA",X"37",X"0D",
		X"3E",X"90",X"BB",X"CA",X"37",X"0D",X"3E",X"91",X"BB",X"CA",X"37",X"0D",X"0C",X"0C",X"3E",X"04",
		X"B9",X"D2",X"11",X"0D",X"C3",X"E1",X"0A",X"3E",X"2F",X"CD",X"A8",X"24",X"E6",X"F0",X"C4",X"4C",
		X"0D",X"21",X"58",X"40",X"7E",X"A7",X"20",X"E4",X"34",X"C3",X"2C",X"0D",X"F5",X"C5",X"D5",X"E5",
		X"EB",X"41",X"0C",X"CD",X"63",X"21",X"7A",X"CB",X"3F",X"57",X"7C",X"CB",X"3F",X"82",X"C6",X"08",
		X"67",X"0E",X"06",X"CD",X"63",X"21",X"7A",X"94",X"38",X"2F",X"16",X"49",X"FE",X"A0",X"D2",X"81",
		X"0D",X"16",X"89",X"FE",X"40",X"D2",X"81",X"0D",X"16",X"C9",X"FE",X"10",X"D2",X"81",X"0D",X"16",
		X"01",X"21",X"18",X"40",X"48",X"06",X"00",X"09",X"AF",X"32",X"01",X"40",X"72",X"23",X"72",X"3E",
		X"0C",X"32",X"01",X"40",X"E1",X"D1",X"C1",X"F1",X"C9",X"ED",X"44",X"16",X"79",X"FE",X"A0",X"D2",
		X"81",X"0D",X"16",X"B9",X"FE",X"40",X"D2",X"81",X"0D",X"16",X"F9",X"FE",X"10",X"D2",X"81",X"0D",
		X"16",X"01",X"C3",X"81",X"0D",X"3E",X"0D",X"32",X"01",X"40",X"AF",X"32",X"58",X"40",X"48",X"06",
		X"06",X"CD",X"B0",X"06",X"05",X"F2",X"C1",X"0D",X"3E",X"01",X"32",X"4C",X"40",X"79",X"E6",X"06",
		X"4F",X"CD",X"63",X"21",X"EB",X"0C",X"CD",X"63",X"21",X"06",X"06",X"CD",X"DF",X"0F",X"CD",X"EB",
		X"0F",X"CD",X"FD",X"0F",X"06",X"07",X"CD",X"DF",X"0F",X"CD",X"4D",X"21",X"0D",X"EB",X"CD",X"4D",
		X"21",X"CD",X"FD",X"0F",X"06",X"01",X"CD",X"DF",X"0F",X"CD",X"EB",X"0F",X"CD",X"FD",X"0F",X"04",
		X"CD",X"DF",X"0F",X"CD",X"4D",X"21",X"0C",X"EB",X"CD",X"4D",X"21",X"CD",X"FD",X"0F",X"06",X"06",
		X"CD",X"DF",X"0F",X"CD",X"EB",X"0F",X"CD",X"FD",X"0F",X"04",X"CD",X"DF",X"0F",X"CD",X"4D",X"21",
		X"0D",X"EB",X"CD",X"4D",X"21",X"CD",X"FD",X"0F",X"06",X"01",X"CD",X"DF",X"0F",X"CD",X"EB",X"0F",
		X"CD",X"FD",X"0F",X"04",X"CD",X"DF",X"0F",X"CD",X"4D",X"21",X"0C",X"EB",X"CD",X"4D",X"21",X"CD",
		X"FD",X"0F",X"04",X"CD",X"DF",X"0F",X"CD",X"EB",X"0F",X"CD",X"FD",X"0F",X"04",X"CD",X"DF",X"0F",
		X"CD",X"4D",X"21",X"0D",X"EB",X"CD",X"4D",X"21",X"CD",X"FD",X"0F",X"11",X"00",X"00",X"0E",X"07",
		X"CD",X"4D",X"21",X"0D",X"F2",X"60",X"0E",X"3A",X"09",X"40",X"4F",X"06",X"00",X"21",X"F0",X"40",
		X"09",X"35",X"CD",X"B9",X"06",X"AF",X"32",X"00",X"68",X"32",X"01",X"68",X"06",X"0A",X"CD",X"FD",
		X"0F",X"10",X"FB",X"3E",X"0E",X"32",X"00",X"40",X"18",X"FE",X"3E",X"0D",X"32",X"01",X"40",X"AF",
		X"32",X"58",X"40",X"06",X"06",X"CD",X"B0",X"06",X"05",X"F2",X"95",X"0E",X"11",X"00",X"00",X"0E",
		X"05",X"CD",X"4D",X"21",X"0D",X"F2",X"A1",X"0E",X"CD",X"09",X"11",X"C3",X"72",X"0E",X"AF",X"32",
		X"01",X"40",X"06",X"06",X"CD",X"B0",X"06",X"05",X"F2",X"B4",X"0E",X"11",X"00",X"00",X"0E",X"05",
		X"CD",X"4D",X"21",X"0D",X"F2",X"C0",X"0E",X"3E",X"0E",X"32",X"01",X"40",X"3A",X"06",X"42",X"A7",
		X"20",X"FA",X"AF",X"32",X"01",X"40",X"06",X"00",X"CD",X"FF",X"20",X"80",X"09",X"02",X"18",X"04",
		X"CD",X"FF",X"20",X"70",X"0A",X"02",X"18",X"04",X"CD",X"FF",X"20",X"80",X"0B",X"06",X"28",X"04",
		X"CD",X"FF",X"20",X"70",X"0C",X"06",X"28",X"CD",X"B9",X"06",X"21",X"18",X"18",X"22",X"10",X"40",
		X"22",X"12",X"40",X"21",X"00",X"00",X"22",X"14",X"40",X"21",X"01",X"01",X"22",X"18",X"40",X"22",
		X"1A",X"40",X"3E",X"0F",X"32",X"01",X"40",X"3A",X"43",X"42",X"FE",X"50",X"38",X"F9",X"AF",X"32",
		X"01",X"40",X"CD",X"FD",X"0F",X"CD",X"FD",X"0F",X"06",X"0F",X"16",X"05",X"CD",X"ED",X"20",X"21",
		X"AE",X"0F",X"11",X"2F",X"52",X"0E",X"04",X"CD",X"3C",X"07",X"06",X"06",X"CD",X"FD",X"0F",X"10",
		X"FB",X"CD",X"B9",X"06",X"3E",X"9F",X"CD",X"A8",X"24",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",
		X"3F",X"21",X"B2",X"0F",X"4F",X"06",X"00",X"09",X"7E",X"67",X"6F",X"22",X"18",X"40",X"22",X"1A",
		X"40",X"21",X"1F",X"1F",X"22",X"10",X"40",X"22",X"12",X"40",X"3E",X"0F",X"32",X"01",X"40",X"06",
		X"04",X"0E",X"03",X"CD",X"63",X"21",X"7A",X"FE",X"F0",X"D2",X"89",X"0F",X"7B",X"FE",X"03",X"DA",
		X"89",X"0F",X"0D",X"F2",X"73",X"0F",X"C3",X"71",X"0F",X"11",X"10",X"00",X"CD",X"4D",X"21",X"21",
		X"10",X"40",X"16",X"00",X"59",X"19",X"36",X"00",X"05",X"C2",X"82",X"0F",X"AF",X"32",X"01",X"40",
		X"06",X"03",X"CD",X"FD",X"0F",X"10",X"FB",X"3E",X"0F",X"32",X"00",X"40",X"18",X"FE",X"FC",X"6A",
		X"6A",X"64",X"79",X"49",X"38",X"08",X"7F",X"BF",X"8F",X"FF",X"CF",X"4F",X"3A",X"09",X"40",X"4F",
		X"06",X"00",X"21",X"F0",X"40",X"09",X"7E",X"A7",X"16",X"12",X"CA",X"D9",X"0F",X"3A",X"0D",X"40",
		X"FE",X"18",X"16",X"11",X"CA",X"D9",X"0F",X"16",X"10",X"21",X"00",X"40",X"72",X"18",X"FE",X"C5",
		X"0E",X"06",X"CD",X"1B",X"24",X"0C",X"CD",X"1B",X"24",X"C1",X"C9",X"D5",X"C5",X"F5",X"4F",X"11",
		X"00",X"00",X"CD",X"4D",X"21",X"0C",X"CD",X"4D",X"21",X"F1",X"C1",X"D1",X"C9",X"F5",X"3E",X"0D",
		X"32",X"07",X"40",X"3A",X"07",X"40",X"A7",X"C2",X"03",X"10",X"F1",X"C9",X"F5",X"C5",X"E5",X"21",
		X"50",X"41",X"06",X"00",X"09",X"06",X"0F",X"3A",X"09",X"40",X"A7",X"C2",X"20",X"10",X"06",X"F0",
		X"7E",X"A0",X"77",X"E1",X"C1",X"F1",X"C9",X"CD",X"BD",X"04",X"CD",X"BF",X"10",X"CD",X"33",X"06",
		X"CD",X"29",X"03",X"CD",X"4F",X"03",X"CD",X"FC",X"05",X"CD",X"89",X"02",X"CD",X"56",X"10",X"CD",
		X"D1",X"03",X"CD",X"BF",X"05",X"C9",X"CD",X"BD",X"04",X"CD",X"33",X"06",X"CD",X"FC",X"05",X"CD",
		X"BF",X"05",X"C9",X"C3",X"89",X"02",X"0E",X"05",X"21",X"C6",X"40",X"3A",X"09",X"40",X"5F",X"16",
		X"00",X"19",X"7E",X"A7",X"CA",X"72",X"10",X"FE",X"8C",X"CA",X"7A",X"10",X"FE",X"01",X"CA",X"9B",
		X"10",X"35",X"2B",X"2B",X"0D",X"0D",X"F2",X"62",X"10",X"C9",X"79",X"CB",X"3F",X"CB",X"3F",X"CB",
		X"27",X"ED",X"44",X"C6",X"0A",X"47",X"CD",X"63",X"21",X"82",X"57",X"CD",X"4D",X"21",X"0D",X"90",
		X"90",X"D6",X"14",X"57",X"CD",X"4D",X"21",X"0C",X"C3",X"71",X"10",X"CD",X"63",X"21",X"E5",X"EB",
		X"0D",X"CD",X"63",X"21",X"79",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"ED",X"44",X"C6",X"10",X"82",
		X"57",X"CD",X"4D",X"21",X"0C",X"C6",X"14",X"57",X"CD",X"4D",X"21",X"E1",X"C3",X"71",X"10",X"21",
		X"C8",X"40",X"3A",X"09",X"40",X"4F",X"06",X"00",X"09",X"7E",X"A7",X"C8",X"FE",X"1F",X"30",X"07",
		X"FE",X"01",X"CC",X"F2",X"10",X"35",X"C9",X"CD",X"F2",X"10",X"36",X"1E",X"D6",X"21",X"ED",X"44",
		X"0E",X"06",X"CD",X"63",X"21",X"1E",X"F0",X"CD",X"2E",X"24",X"11",X"E0",X"FF",X"77",X"3C",X"19",
		X"77",X"C9",X"F5",X"C5",X"D5",X"E5",X"21",X"1E",X"50",X"11",X"20",X"00",X"3E",X"FF",X"06",X"20",
		X"77",X"19",X"10",X"FC",X"E1",X"D1",X"C1",X"F1",X"C9",X"3E",X"01",X"32",X"3A",X"40",X"21",X"09",
		X"40",X"4E",X"06",X"00",X"21",X"F0",X"40",X"09",X"35",X"21",X"07",X"40",X"77",X"DD",X"21",X"50",
		X"42",X"FD",X"21",X"7F",X"40",X"D6",X"02",X"FD",X"77",X"00",X"3E",X"02",X"CD",X"C9",X"11",X"3E",
		X"05",X"CD",X"D6",X"11",X"DD",X"7E",X"08",X"FE",X"18",X"38",X"16",X"FE",X"D8",X"30",X"24",X"D6",
		X"08",X"DD",X"77",X"00",X"DD",X"77",X"04",X"C6",X"10",X"DD",X"77",X"08",X"DD",X"77",X"0C",X"18",
		X"22",X"3E",X"10",X"DD",X"77",X"00",X"DD",X"77",X"04",X"3E",X"20",X"DD",X"77",X"08",X"DD",X"77",
		X"0C",X"18",X"10",X"3E",X"D0",X"DD",X"77",X"00",X"DD",X"77",X"04",X"3E",X"E0",X"DD",X"77",X"08",
		X"DD",X"77",X"0C",X"DD",X"7E",X"0B",X"DD",X"77",X"03",X"DD",X"7E",X"0F",X"DD",X"77",X"07",X"CD",
		X"FD",X"0F",X"FD",X"34",X"00",X"FD",X"7E",X"00",X"FE",X"0C",X"C8",X"E6",X"03",X"FE",X"01",X"28",
		X"14",X"FE",X"02",X"28",X"1C",X"FE",X"03",X"28",X"24",X"3E",X"02",X"CD",X"C9",X"11",X"3E",X"05",
		X"CD",X"D6",X"11",X"18",X"DA",X"3E",X"01",X"CD",X"C9",X"11",X"3E",X"11",X"CD",X"D6",X"11",X"18",
		X"CE",X"3E",X"06",X"CD",X"C9",X"11",X"3E",X"05",X"CD",X"D6",X"11",X"18",X"C2",X"3E",X"07",X"CD",
		X"C9",X"11",X"3E",X"11",X"CD",X"D6",X"11",X"18",X"B6",X"DD",X"77",X"02",X"DD",X"77",X"06",X"DD",
		X"77",X"0A",X"DD",X"77",X"0E",X"C9",X"DD",X"77",X"09",X"3C",X"DD",X"77",X"0D",X"3C",X"DD",X"77",
		X"01",X"3C",X"DD",X"77",X"05",X"C9",X"CD",X"B9",X"06",X"0E",X"07",X"11",X"00",X"00",X"CD",X"4D",
		X"21",X"0D",X"F2",X"EE",X"11",X"21",X"F2",X"40",X"06",X"00",X"3A",X"09",X"40",X"4F",X"09",X"3E",
		X"03",X"77",X"21",X"F3",X"40",X"09",X"46",X"3E",X"0A",X"3D",X"10",X"FD",X"32",X"95",X"40",X"3E",
		X"18",X"32",X"75",X"40",X"3E",X"01",X"32",X"96",X"40",X"3E",X"0E",X"32",X"77",X"40",X"3E",X"0F",
		X"32",X"78",X"40",X"CD",X"55",X"07",X"06",X"00",X"CD",X"FF",X"20",X"80",X"0B",X"06",X"28",X"04",
		X"CD",X"FF",X"20",X"80",X"09",X"02",X"18",X"04",X"CD",X"FF",X"20",X"70",X"0C",X"06",X"28",X"04",
		X"CD",X"FF",X"20",X"70",X"0A",X"02",X"18",X"11",X"05",X"0E",X"CD",X"7A",X"18",X"16",X"06",X"06",
		X"1D",X"04",X"CD",X"ED",X"20",X"05",X"05",X"20",X"F8",X"AF",X"DD",X"21",X"00",X"42",X"DD",X"77",
		X"06",X"DD",X"77",X"08",X"DD",X"77",X"0A",X"DD",X"77",X"0C",X"21",X"F1",X"40",X"06",X"00",X"3A",
		X"09",X"40",X"4F",X"09",X"7E",X"CD",X"B4",X"13",X"21",X"FF",X"FF",X"22",X"00",X"68",X"22",X"01",
		X"68",X"3E",X"01",X"32",X"72",X"40",X"32",X"79",X"40",X"3E",X"10",X"32",X"01",X"40",X"3E",X"0A",
		X"CD",X"6F",X"18",X"BB",X"30",X"FA",X"AF",X"32",X"01",X"40",X"3E",X"06",X"CD",X"12",X"13",X"C6",
		X"05",X"CD",X"0C",X"14",X"06",X"00",X"21",X"F1",X"40",X"3A",X"09",X"40",X"4F",X"09",X"7E",X"3D",
		X"3E",X"12",X"28",X"02",X"3D",X"3D",X"32",X"01",X"40",X"CD",X"6F",X"18",X"7A",X"CB",X"7F",X"20",
		X"17",X"FE",X"08",X"38",X"13",X"FE",X"15",X"30",X"10",X"7B",X"CB",X"7F",X"20",X"2B",X"FE",X"08",
		X"38",X"27",X"FE",X"1A",X"30",X"24",X"18",X"4A",X"AF",X"F5",X"7B",X"FE",X"15",X"38",X"07",X"3E",
		X"02",X"CD",X"12",X"13",X"18",X"05",X"3E",X"06",X"CD",X"12",X"13",X"3C",X"CD",X"0C",X"14",X"47",
		X"F1",X"A7",X"78",X"28",X"18",X"C6",X"30",X"18",X"14",X"AF",X"F5",X"3E",X"06",X"CD",X"12",X"13",
		X"C6",X"05",X"CD",X"0C",X"14",X"47",X"F1",X"A7",X"78",X"28",X"02",X"C6",X"06",X"32",X"72",X"40",
		X"18",X"10",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"CD",X"A8",X"24",X"CB",X"3F",X"CB",X"3F",X"CB",
		X"3F",X"C9",X"06",X"07",X"0E",X"13",X"05",X"CD",X"B4",X"26",X"DC",X"64",X"13",X"04",X"0D",X"3E",
		X"0D",X"B9",X"20",X"02",X"0E",X"07",X"3E",X"FF",X"B9",X"20",X"EB",X"10",X"E7",X"06",X"07",X"05",
		X"CD",X"32",X"26",X"DA",X"8F",X"13",X"04",X"10",X"F6",X"06",X"0E",X"05",X"CD",X"0F",X"26",X"DA",
		X"E5",X"13",X"04",X"10",X"F6",X"06",X"07",X"05",X"CD",X"20",X"26",X"DA",X"E5",X"13",X"04",X"10",
		X"F6",X"C3",X"B9",X"12",X"21",X"20",X"40",X"58",X"16",X"00",X"19",X"7E",X"CB",X"7F",X"28",X"0B",
		X"F5",X"3E",X"01",X"32",X"60",X"40",X"F1",X"ED",X"44",X"77",X"C9",X"57",X"79",X"FE",X"11",X"C8",
		X"FE",X"10",X"C8",X"FE",X"05",X"C8",X"FE",X"04",X"C8",X"FE",X"03",X"C8",X"7A",X"18",X"E1",X"3E",
		X"01",X"32",X"50",X"40",X"11",X"00",X"00",X"CD",X"86",X"21",X"21",X"F1",X"40",X"06",X"00",X"3A",
		X"09",X"40",X"4F",X"09",X"34",X"7E",X"FE",X"02",X"28",X"31",X"CD",X"B4",X"13",X"FE",X"01",X"28",
		X"1E",X"C3",X"46",X"13",X"21",X"C5",X"13",X"4F",X"09",X"46",X"DD",X"21",X"42",X"42",X"DD",X"70",
		X"00",X"DD",X"70",X"08",X"C9",X"06",X"06",X"07",X"01",X"06",X"07",X"01",X"03",X"04",X"06",X"AF",
		X"32",X"7F",X"40",X"3E",X"12",X"32",X"01",X"40",X"C3",X"46",X"13",X"CD",X"FB",X"13",X"CD",X"C1",
		X"14",X"3E",X"19",X"18",X"08",X"CD",X"FB",X"13",X"CD",X"09",X"11",X"3E",X"1A",X"21",X"00",X"00",
		X"22",X"00",X"68",X"22",X"01",X"68",X"32",X"00",X"40",X"18",X"FE",X"AF",X"32",X"01",X"40",X"11",
		X"00",X"00",X"06",X"07",X"05",X"CD",X"86",X"21",X"04",X"10",X"F9",X"C9",X"21",X"15",X"14",X"16",
		X"00",X"5F",X"19",X"7E",X"C9",X"07",X"CF",X"8F",X"4F",X"08",X"49",X"89",X"C9",X"01",X"F9",X"B9",
		X"79",X"38",X"7F",X"BF",X"FF",X"21",X"F0",X"40",X"06",X"00",X"3A",X"09",X"40",X"4F",X"09",X"7E",
		X"FE",X"00",X"28",X"0D",X"23",X"7E",X"FE",X"0A",X"28",X"0B",X"3E",X"1D",X"32",X"00",X"40",X"18",
		X"FE",X"3E",X"1B",X"18",X"F7",X"3E",X"1C",X"18",X"F3",X"3A",X"08",X"40",X"3D",X"28",X"3E",X"3A",
		X"09",X"40",X"A7",X"20",X"03",X"3E",X"40",X"CB",X"AF",X"32",X"09",X"40",X"21",X"F0",X"40",X"4F",
		X"06",X"00",X"09",X"7E",X"A7",X"79",X"28",X"E1",X"21",X"00",X"70",X"CB",X"4E",X"20",X"0F",X"A7",
		X"28",X"05",X"01",X"01",X"01",X"18",X"03",X"01",X"00",X"00",X"ED",X"43",X"06",X"70",X"CD",X"B9",
		X"06",X"11",X"00",X"00",X"0E",X"07",X"CD",X"4D",X"21",X"0D",X"F2",X"86",X"14",X"21",X"F2",X"40",
		X"06",X"00",X"4F",X"09",X"46",X"3E",X"1E",X"80",X"32",X"00",X"40",X"18",X"FE",X"21",X"7F",X"40",
		X"34",X"7E",X"E6",X"F0",X"BE",X"C0",X"DD",X"E5",X"7E",X"E6",X"E0",X"BE",X"DD",X"21",X"42",X"42",
		X"28",X"0B",X"3E",X"02",X"DD",X"77",X"00",X"DD",X"77",X"08",X"DD",X"E1",X"C9",X"3E",X"04",X"18",
		X"F3",X"3E",X"01",X"32",X"3A",X"40",X"21",X"07",X"40",X"77",X"DD",X"21",X"40",X"42",X"FD",X"21",
		X"7F",X"40",X"D6",X"02",X"FD",X"77",X"00",X"3E",X"02",X"CD",X"41",X"15",X"3E",X"05",X"CD",X"4E",
		X"15",X"DD",X"7E",X"00",X"DD",X"77",X"10",X"D6",X"10",X"DD",X"77",X"14",X"DD",X"7E",X"03",X"C6",
		X"10",X"DD",X"77",X"13",X"DD",X"77",X"17",X"CD",X"FD",X"0F",X"FD",X"34",X"00",X"FD",X"7E",X"00",
		X"FE",X"0C",X"C8",X"E6",X"03",X"FE",X"01",X"28",X"14",X"FE",X"02",X"28",X"1C",X"FE",X"03",X"28",
		X"24",X"3E",X"02",X"CD",X"41",X"15",X"3E",X"05",X"CD",X"4E",X"15",X"18",X"DA",X"3E",X"01",X"CD",
		X"41",X"15",X"3E",X"11",X"CD",X"4E",X"15",X"18",X"CE",X"3E",X"06",X"CD",X"41",X"15",X"3E",X"05",
		X"CD",X"4E",X"15",X"18",X"C2",X"3E",X"07",X"CD",X"41",X"15",X"3E",X"11",X"CD",X"4E",X"15",X"18",
		X"B6",X"DD",X"77",X"12",X"DD",X"77",X"16",X"DD",X"77",X"0A",X"DD",X"77",X"02",X"C9",X"DD",X"77",
		X"01",X"3C",X"DD",X"77",X"11",X"3C",X"DD",X"77",X"09",X"3C",X"DD",X"77",X"15",X"C9",X"CD",X"B9",
		X"06",X"06",X"08",X"11",X"00",X"00",X"48",X"0D",X"CD",X"4D",X"21",X"10",X"F9",X"3E",X"1F",X"3D",
		X"47",X"16",X"00",X"CD",X"DC",X"20",X"16",X"03",X"CD",X"ED",X"20",X"FE",X"02",X"20",X"F0",X"3A",
		X"09",X"40",X"FE",X"00",X"28",X"05",X"21",X"AA",X"16",X"18",X"03",X"21",X"A1",X"16",X"22",X"8E",
		X"40",X"3E",X"0C",X"32",X"7F",X"40",X"AF",X"32",X"8A",X"40",X"3E",X"18",X"32",X"8B",X"40",X"3E",
		X"E0",X"32",X"8C",X"40",X"3E",X"E8",X"32",X"8D",X"40",X"3E",X"14",X"32",X"01",X"40",X"3A",X"01",
		X"40",X"FE",X"00",X"20",X"F9",X"3E",X"7D",X"32",X"07",X"40",X"3A",X"07",X"40",X"A7",X"20",X"FA",
		X"3A",X"F0",X"40",X"A7",X"20",X"1D",X"3A",X"08",X"40",X"3D",X"28",X"06",X"3A",X"30",X"41",X"A7",
		X"20",X"11",X"21",X"00",X"00",X"22",X"06",X"70",X"AF",X"32",X"F2",X"40",X"32",X"32",X"41",X"3E",
		X"05",X"18",X"02",X"3E",X"14",X"32",X"00",X"40",X"18",X"FE",X"21",X"07",X"40",X"7E",X"E6",X"F8",
		X"BE",X"C0",X"3A",X"8A",X"40",X"32",X"82",X"40",X"3A",X"8B",X"40",X"32",X"83",X"40",X"CD",X"51",
		X"16",X"3A",X"8C",X"40",X"32",X"82",X"40",X"CD",X"51",X"16",X"3E",X"60",X"32",X"82",X"40",X"3A",
		X"8D",X"40",X"32",X"83",X"40",X"CD",X"51",X"16",X"21",X"8A",X"40",X"CD",X"5A",X"16",X"21",X"8B",
		X"40",X"CD",X"66",X"16",X"21",X"99",X"16",X"CD",X"54",X"16",X"21",X"8C",X"40",X"CD",X"62",X"16",
		X"21",X"9D",X"16",X"CD",X"54",X"16",X"3E",X"60",X"32",X"82",X"40",X"21",X"8D",X"40",X"CD",X"6E",
		X"16",X"2A",X"8E",X"40",X"CD",X"54",X"16",X"21",X"7F",X"40",X"35",X"C0",X"AF",X"32",X"01",X"40",
		X"C9",X"21",X"90",X"16",X"22",X"80",X"40",X"C3",X"72",X"16",X"3E",X"08",X"86",X"77",X"32",X"82",
		X"40",X"C9",X"3E",X"F8",X"18",X"F6",X"3E",X"08",X"86",X"77",X"32",X"83",X"40",X"C9",X"3E",X"F8",
		X"18",X"F6",X"2A",X"80",X"40",X"3A",X"82",X"40",X"57",X"3A",X"83",X"40",X"5F",X"E5",X"CD",X"2E",
		X"24",X"EB",X"E1",X"01",X"E0",X"FF",X"7E",X"A7",X"C8",X"12",X"EB",X"09",X"EB",X"23",X"18",X"F6",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"6E",X"66",X"65",X"00",X"65",X"69",X"64",
		X"00",X"6B",X"68",X"62",X"70",X"65",X"6C",X"FF",X"59",X"00",X"6B",X"68",X"62",X"70",X"65",X"6C",
		X"FF",X"5A",X"00",X"3A",X"71",X"40",X"CB",X"7F",X"20",X"44",X"FE",X"1C",X"30",X"40",X"3A",X"70",
		X"40",X"CB",X"7F",X"20",X"39",X"FE",X"02",X"38",X"35",X"FE",X"1F",X"30",X"31",X"3A",X"71",X"40",
		X"CB",X"27",X"CB",X"27",X"CB",X"27",X"57",X"3A",X"70",X"40",X"CB",X"27",X"CB",X"27",X"CB",X"27",
		X"5F",X"0E",X"02",X"CD",X"4D",X"21",X"C6",X"F0",X"5F",X"0C",X"CD",X"4D",X"21",X"7A",X"C6",X"10",
		X"57",X"0D",X"0D",X"CD",X"4D",X"21",X"7B",X"C6",X"10",X"5F",X"0D",X"C3",X"4D",X"21",X"11",X"00",
		X"00",X"0E",X"00",X"CD",X"4D",X"21",X"0C",X"CD",X"4D",X"21",X"0C",X"CD",X"4D",X"21",X"0C",X"C3",
		X"4D",X"21",X"21",X"96",X"40",X"35",X"7E",X"A7",X"28",X"14",X"21",X"77",X"40",X"46",X"21",X"78",
		X"40",X"4E",X"CD",X"6F",X"18",X"7A",X"B8",X"20",X"32",X"7B",X"B9",X"C8",X"18",X"2D",X"3A",X"95",
		X"40",X"CB",X"27",X"CB",X"27",X"77",X"3A",X"7E",X"40",X"A7",X"20",X"04",X"3E",X"30",X"18",X"01",
		X"AF",X"32",X"7E",X"40",X"21",X"74",X"40",X"34",X"7E",X"FE",X"0E",X"20",X"02",X"AF",X"77",X"21",
		X"75",X"40",X"35",X"7E",X"FE",X"0D",X"20",X"03",X"3E",X"17",X"77",X"3A",X"76",X"40",X"06",X"00",
		X"4F",X"DD",X"21",X"83",X"23",X"DD",X"09",X"3A",X"09",X"40",X"4F",X"21",X"C0",X"40",X"09",X"7E",
		X"CB",X"7F",X"20",X"13",X"3A",X"77",X"40",X"DD",X"86",X"01",X"57",X"3A",X"78",X"40",X"DD",X"86",
		X"00",X"5F",X"3E",X"FF",X"CD",X"83",X"18",X"DD",X"23",X"DD",X"23",X"23",X"04",X"3E",X"18",X"B8",
		X"20",X"DD",X"CD",X"6F",X"18",X"06",X"00",X"3A",X"7E",X"40",X"32",X"76",X"40",X"4F",X"DD",X"21",
		X"83",X"23",X"DD",X"09",X"7A",X"32",X"77",X"40",X"7B",X"32",X"78",X"40",X"3A",X"09",X"40",X"4F",
		X"21",X"C0",X"40",X"09",X"3A",X"77",X"40",X"DD",X"86",X"01",X"57",X"FA",X"F0",X"17",X"FE",X"02",
		X"38",X"2E",X"FE",X"1E",X"30",X"2A",X"3A",X"78",X"40",X"DD",X"86",X"00",X"5F",X"FA",X"F0",X"17",
		X"FE",X"02",X"38",X"1C",X"FE",X"1F",X"30",X"18",X"3A",X"74",X"40",X"B8",X"28",X"0A",X"3A",X"75",
		X"40",X"B8",X"28",X"04",X"3E",X"54",X"18",X"02",X"3E",X"56",X"77",X"CD",X"83",X"18",X"18",X"03",
		X"3E",X"FF",X"77",X"DD",X"23",X"DD",X"23",X"23",X"04",X"3E",X"18",X"B8",X"20",X"B6",X"C9",X"21",
		X"79",X"40",X"35",X"7E",X"A7",X"C0",X"3A",X"95",X"40",X"77",X"21",X"90",X"40",X"7E",X"3C",X"E6",
		X"07",X"77",X"57",X"21",X"72",X"40",X"5E",X"7B",X"E6",X"C0",X"28",X"27",X"AF",X"82",X"CA",X"B3",
		X"16",X"CB",X"47",X"28",X"1E",X"7B",X"E6",X"C0",X"FE",X"40",X"28",X"3C",X"FE",X"80",X"28",X"13",
		X"7B",X"E6",X"07",X"CB",X"57",X"C4",X"6C",X"18",X"CD",X"6F",X"18",X"83",X"5F",X"CD",X"7A",X"18",
		X"C3",X"B3",X"16",X"7B",X"E6",X"07",X"CB",X"57",X"C4",X"6C",X"18",X"6F",X"7B",X"E6",X"38",X"CB",
		X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"57",X"C4",X"6C",X"18",X"CD",X"6F",X"18",X"82",X"57",X"7D",
		X"83",X"5F",X"CD",X"7A",X"18",X"C3",X"B3",X"16",X"2E",X"00",X"18",X"E0",X"3E",X"FF",X"C9",X"E5",
		X"21",X"71",X"40",X"56",X"21",X"70",X"40",X"5E",X"E1",X"C9",X"21",X"71",X"40",X"72",X"21",X"70",
		X"40",X"73",X"C9",X"CB",X"22",X"CB",X"22",X"CB",X"22",X"CB",X"23",X"CB",X"23",X"CB",X"23",X"E5",
		X"CD",X"2E",X"24",X"77",X"E1",X"C9",X"CD",X"FF",X"17",X"CD",X"12",X"17",X"CD",X"D1",X"03",X"CD",
		X"4F",X"03",X"CD",X"29",X"03",X"C9",X"CD",X"D1",X"03",X"CD",X"4F",X"03",X"CD",X"29",X"03",X"C9",
		X"CD",X"FF",X"17",X"CD",X"12",X"17",X"CD",X"D1",X"03",X"CD",X"4F",X"03",X"CD",X"29",X"03",X"CD",
		X"9D",X"14",X"C9",X"CD",X"EA",X"15",X"C9",X"CD",X"95",X"24",X"CD",X"C5",X"20",X"21",X"06",X"70",
		X"AF",X"77",X"23",X"77",X"06",X"1F",X"16",X"06",X"CD",X"ED",X"20",X"06",X"16",X"16",X"02",X"CD",
		X"ED",X"20",X"04",X"CD",X"ED",X"20",X"21",X"C1",X"1A",X"22",X"88",X"40",X"21",X"C6",X"52",X"22",
		X"BE",X"40",X"3E",X"01",X"32",X"04",X"70",X"CD",X"BB",X"19",X"CD",X"92",X"19",X"3E",X"01",X"32",
		X"01",X"40",X"3A",X"0C",X"42",X"FE",X"4F",X"20",X"F9",X"3E",X"02",X"32",X"01",X"40",X"3A",X"0C",
		X"42",X"A7",X"20",X"FA",X"06",X"7D",X"CD",X"06",X"1A",X"21",X"C6",X"52",X"22",X"BE",X"40",X"3E",
		X"02",X"32",X"01",X"40",X"3A",X"0C",X"42",X"FE",X"B7",X"20",X"F9",X"3E",X"03",X"32",X"01",X"40",
		X"3A",X"0C",X"42",X"FE",X"57",X"20",X"F9",X"06",X"82",X"CD",X"06",X"1A",X"AF",X"32",X"01",X"40",
		X"3C",X"32",X"00",X"40",X"18",X"FE",X"3A",X"12",X"42",X"E6",X"07",X"20",X"03",X"CD",X"66",X"19",
		X"CD",X"81",X"19",X"C9",X"CD",X"81",X"19",X"C9",X"3A",X"0C",X"42",X"E6",X"07",X"20",X"03",X"CD",
		X"A0",X"19",X"CD",X"81",X"19",X"C9",X"2A",X"88",X"40",X"ED",X"5B",X"BE",X"40",X"06",X"08",X"7E",
		X"12",X"23",X"13",X"10",X"FA",X"22",X"88",X"40",X"EB",X"11",X"D8",X"FF",X"19",X"22",X"BE",X"40",
		X"C9",X"3A",X"0C",X"42",X"57",X"15",X"0E",X"08",X"06",X"06",X"CD",X"DC",X"20",X"04",X"0D",X"20",
		X"F9",X"C9",X"0E",X"08",X"06",X"06",X"16",X"B0",X"CD",X"DC",X"20",X"04",X"0D",X"20",X"F9",X"C9",
		X"2A",X"BE",X"40",X"06",X"08",X"36",X"FF",X"23",X"10",X"FB",X"11",X"D8",X"FF",X"19",X"22",X"BE",
		X"40",X"C9",X"06",X"08",X"0A",X"0C",X"01",X"07",X"09",X"0B",X"0D",X"21",X"B2",X"19",X"0E",X"04",
		X"16",X"01",X"46",X"CD",X"ED",X"20",X"0D",X"23",X"20",X"F8",X"0E",X"05",X"16",X"03",X"46",X"CD",
		X"ED",X"20",X"0D",X"23",X"20",X"F8",X"11",X"2C",X"1A",X"21",X"60",X"53",X"CD",X"FB",X"19",X"11",
		X"29",X"1B",X"21",X"D6",X"52",X"CD",X"FB",X"19",X"11",X"33",X"1B",X"21",X"17",X"53",X"CD",X"FB",
		X"19",X"11",X"45",X"1A",X"21",X"BF",X"53",X"CD",X"FB",X"19",X"C9",X"01",X"E0",X"FF",X"1A",X"A7",
		X"C8",X"77",X"09",X"13",X"18",X"F5",X"AF",X"32",X"01",X"40",X"78",X"32",X"07",X"40",X"3A",X"07",
		X"40",X"A7",X"20",X"FA",X"C9",X"E5",X"D5",X"C5",X"21",X"00",X"50",X"06",X"00",X"09",X"11",X"20",
		X"00",X"06",X"20",X"36",X"FF",X"19",X"10",X"FB",X"C1",X"D1",X"E1",X"C9",X"59",X"6B",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"66",X"67",X"FF",X"6D",X"63",X"6A",X"6C",X"65",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"5A",X"6B",X"00",X"63",X"6C",X"65",X"64",X"67",X"6E",X"00",X"6B",X"6A",X"67",X"69",
		X"6E",X"6D",X"FF",X"00",X"6F",X"68",X"62",X"63",X"55",X"FF",X"66",X"6A",X"68",X"65",X"00",X"6F",
		X"6A",X"69",X"FD",X"6D",X"FF",X"6B",X"6A",X"67",X"69",X"6E",X"00",X"62",X"64",X"64",X"FF",X"59",
		X"FF",X"6C",X"6A",X"63",X"55",X"65",X"6E",X"00",X"63",X"67",X"6E",X"70",X"FF",X"6C",X"65",X"6D",
		X"63",X"FD",X"65",X"FF",X"00",X"67",X"69",X"6D",X"65",X"6C",X"6E",X"FF",X"63",X"6A",X"67",X"69",
		X"00",X"59",X"FF",X"6A",X"6C",X"FF",X"5A",X"FF",X"6B",X"68",X"62",X"70",X"65",X"6C",X"6D",X"FF",
		X"00",X"6B",X"FD",X"6D",X"66",X"00",X"6B",X"68",X"62",X"70",X"00",X"6A",X"69",X"68",X"70",X"FF",
		X"59",X"FF",X"6B",X"68",X"62",X"70",X"65",X"6C",X"FF",X"00",X"6F",X"FD",X"6E",X"6E",X"6A",X"69",
		X"00",X"FF",X"8A",X"8B",X"8C",X"8D",X"8E",X"8F",X"90",X"FF",X"FF",X"91",X"92",X"93",X"94",X"95",
		X"96",X"FF",X"97",X"98",X"99",X"9A",X"9B",X"9C",X"9D",X"FF",X"9E",X"9F",X"A0",X"A1",X"A2",X"A3",
		X"A4",X"FF",X"A5",X"A6",X"A7",X"A8",X"A9",X"AA",X"AB",X"FF",X"AC",X"AD",X"AE",X"AF",X"B0",X"B1",
		X"B2",X"FF",X"B3",X"B4",X"B5",X"B6",X"B7",X"B8",X"FF",X"B9",X"BA",X"BB",X"BC",X"BD",X"BE",X"BF",
		X"FF",X"C0",X"C1",X"C2",X"C3",X"C4",X"C5",X"FF",X"FF",X"C6",X"C7",X"C8",X"C9",X"CA",X"CB",X"FF",
		X"FF",X"CC",X"CD",X"CE",X"CF",X"D0",X"D1",X"FF",X"FF",X"D2",X"D3",X"D4",X"D5",X"D6",X"FF",X"FF",
		X"FF",X"D7",X"D8",X"D9",X"DA",X"DB",X"FF",X"FF",X"FF",X"78",X"7A",X"7C",X"7E",X"80",X"82",X"84",
		X"86",X"88",X"00",X"71",X"FF",X"79",X"7B",X"7D",X"7F",X"81",X"83",X"85",X"87",X"89",X"FF",X"72",
		X"73",X"74",X"75",X"76",X"77",X"00",X"FD",X"FE",X"6A",X"00",X"59",X"58",X"FF",X"00",X"5A",X"58",
		X"FF",X"00",X"5B",X"58",X"FF",X"00",X"5D",X"58",X"FF",X"00",X"5E",X"58",X"FF",X"00",X"59",X"58",
		X"58",X"FF",X"00",X"5B",X"58",X"58",X"FF",X"00",X"5D",X"58",X"58",X"FF",X"00",X"FF",X"5D",X"58",
		X"58",X"58",X"FF",X"00",X"59",X"58",X"58",X"58",X"58",X"FF",X"00",X"59",X"FF",X"63",X"6A",X"67",
		X"69",X"FF",X"FF",X"59",X"FF",X"6B",X"68",X"62",X"70",X"00",X"59",X"FF",X"63",X"6A",X"67",X"69",
		X"FF",X"FF",X"5A",X"FF",X"6B",X"68",X"62",X"70",X"6D",X"00",X"59",X"FF",X"63",X"6A",X"67",X"69",
		X"FF",X"FF",X"5B",X"FF",X"6B",X"68",X"62",X"70",X"6D",X"00",X"5A",X"FF",X"63",X"6A",X"67",X"69",
		X"6D",X"FF",X"FF",X"59",X"FF",X"6B",X"68",X"62",X"70",X"00",X"F1",X"F2",X"F3",X"F4",X"F5",X"F6",
		X"F7",X"00",X"F0",X"F4",X"F4",X"F4",X"F4",X"F4",X"F4",X"F4",X"F8",X"00",X"CD",X"95",X"24",X"CD",
		X"96",X"1F",X"CD",X"A9",X"1F",X"CD",X"D0",X"20",X"CD",X"B6",X"1F",X"11",X"54",X"1A",X"21",X"8A",
		X"52",X"CD",X"C1",X"1F",X"06",X"04",X"CD",X"FF",X"20",X"68",X"02",X"02",X"68",X"11",X"4A",X"1B",
		X"21",X"CD",X"51",X"CD",X"C1",X"1F",X"11",X"4C",X"1A",X"CD",X"C1",X"1F",X"06",X"00",X"CD",X"FF",
		X"20",X"38",X"01",X"01",X"80",X"06",X"01",X"CD",X"FF",X"20",X"60",X"37",X"01",X"80",X"11",X"5E",
		X"1B",X"21",X"F1",X"51",X"CD",X"C1",X"1F",X"11",X"4C",X"1A",X"CD",X"C1",X"1F",X"06",X"02",X"CD",
		X"FF",X"20",X"3A",X"01",X"06",X"A0",X"06",X"03",X"CD",X"FF",X"20",X"5E",X"37",X"06",X"A0",X"11",
		X"63",X"1B",X"21",X"F5",X"51",X"CD",X"C1",X"1F",X"11",X"4C",X"1A",X"CD",X"C1",X"1F",X"06",X"82",
		X"CD",X"06",X"1A",X"3E",X"03",X"32",X"00",X"40",X"18",X"FE",X"CD",X"B9",X"06",X"CD",X"B6",X"1F",
		X"11",X"5F",X"1A",X"21",X"AD",X"52",X"CD",X"C1",X"1F",X"3A",X"00",X"70",X"CB",X"47",X"28",X"05",
		X"11",X"74",X"1B",X"18",X"03",X"11",X"6D",X"1B",X"21",X"6F",X"53",X"CD",X"C1",X"1F",X"11",X"4C",
		X"1A",X"CD",X"C1",X"1F",X"11",X"6B",X"1A",X"CD",X"C1",X"1F",X"11",X"78",X"1A",X"21",X"51",X"53",
		X"CD",X"C1",X"1F",X"11",X"68",X"1B",X"CD",X"C1",X"1F",X"11",X"4C",X"1A",X"CD",X"C1",X"1F",X"06",
		X"41",X"CD",X"06",X"1A",X"3E",X"04",X"32",X"00",X"40",X"18",X"FE",X"0E",X"0D",X"CD",X"15",X"1A",
		X"0E",X"0F",X"CD",X"15",X"1A",X"0E",X"11",X"CD",X"15",X"1A",X"11",X"85",X"1A",X"21",X"AA",X"52",
		X"CD",X"C1",X"1F",X"11",X"91",X"1A",X"21",X"CC",X"52",X"CD",X"C1",X"1F",X"21",X"D1",X"1C",X"3A",
		X"00",X"68",X"CB",X"07",X"CB",X"07",X"E6",X"03",X"47",X"87",X"87",X"80",X"4F",X"06",X"00",X"09",
		X"E9",X"11",X"7B",X"1B",X"18",X"0D",X"11",X"8A",X"1B",X"18",X"08",X"11",X"9A",X"1B",X"18",X"03",
		X"11",X"AA",X"1B",X"21",X"CF",X"52",X"CD",X"C1",X"1F",X"06",X"82",X"CD",X"06",X"1A",X"06",X"06",
		X"C5",X"0E",X"0A",X"CD",X"15",X"1A",X"06",X"19",X"CD",X"06",X"1A",X"11",X"85",X"1A",X"21",X"AA",
		X"52",X"CD",X"FB",X"19",X"06",X"19",X"CD",X"06",X"1A",X"C1",X"10",X"E4",X"06",X"82",X"CD",X"06",
		X"1A",X"3E",X"05",X"32",X"00",X"40",X"18",X"FE",X"31",X"00",X"44",X"AF",X"21",X"06",X"70",X"77",
		X"23",X"77",X"32",X"F1",X"40",X"32",X"31",X"41",X"3E",X"59",X"32",X"F4",X"40",X"32",X"34",X"41",
		X"3E",X"01",X"32",X"F3",X"40",X"32",X"33",X"41",X"3C",X"3C",X"32",X"F0",X"40",X"32",X"30",X"41",
		X"21",X"09",X"40",X"36",X"00",X"21",X"7C",X"40",X"36",X"59",X"23",X"36",X"59",X"CD",X"95",X"24",
		X"06",X"80",X"21",X"00",X"42",X"36",X"00",X"23",X"10",X"FB",X"CD",X"96",X"1F",X"06",X"01",X"16",
		X"03",X"CD",X"ED",X"20",X"06",X"1F",X"16",X"06",X"CD",X"ED",X"20",X"16",X"03",X"06",X"0C",X"CD",
		X"ED",X"20",X"06",X"0E",X"CD",X"ED",X"20",X"11",X"A1",X"1A",X"21",X"2C",X"52",X"CD",X"FB",X"19",
		X"3A",X"03",X"40",X"3D",X"28",X"11",X"11",X"91",X"1A",X"21",X"2E",X"53",X"CD",X"FB",X"19",X"11",
		X"BA",X"1A",X"CD",X"FB",X"19",X"18",X"0F",X"11",X"AB",X"1A",X"21",X"2E",X"53",X"CD",X"FB",X"19",
		X"11",X"BA",X"1A",X"CD",X"FB",X"19",X"3E",X"06",X"32",X"00",X"40",X"18",X"FE",X"CD",X"95",X"24",
		X"CD",X"96",X"1F",X"21",X"C0",X"40",X"3A",X"09",X"40",X"16",X"00",X"5F",X"19",X"06",X"2A",X"36",
		X"FF",X"23",X"10",X"FB",X"3E",X"59",X"21",X"F4",X"40",X"19",X"77",X"AF",X"21",X"F1",X"40",X"19",
		X"77",X"CD",X"B6",X"1F",X"06",X"03",X"16",X"02",X"CD",X"ED",X"20",X"04",X"CD",X"ED",X"20",X"16",
		X"06",X"04",X"CD",X"ED",X"20",X"04",X"CD",X"ED",X"20",X"06",X"03",X"16",X"00",X"CD",X"DC",X"20",
		X"04",X"CD",X"DC",X"20",X"04",X"CD",X"DC",X"20",X"04",X"CD",X"DC",X"20",X"3E",X"01",X"32",X"40",
		X"40",X"AF",X"32",X"3F",X"40",X"3A",X"08",X"40",X"3D",X"20",X"0F",X"21",X"A0",X"50",X"36",X"FF",
		X"21",X"80",X"50",X"36",X"FF",X"0E",X"01",X"CD",X"15",X"1A",X"CD",X"97",X"1E",X"3E",X"04",X"32",
		X"01",X"40",X"3A",X"43",X"42",X"FE",X"E0",X"20",X"F9",X"AF",X"32",X"01",X"40",X"3E",X"05",X"32",
		X"01",X"40",X"3A",X"4B",X"42",X"FE",X"D0",X"20",X"F9",X"3E",X"06",X"32",X"01",X"40",X"3A",X"4B",
		X"42",X"FE",X"18",X"20",X"F9",X"AF",X"32",X"01",X"40",X"CD",X"D7",X"1E",X"3E",X"07",X"32",X"00",
		X"40",X"18",X"FE",X"0E",X"00",X"CD",X"63",X"21",X"1C",X"1C",X"CD",X"4D",X"21",X"0C",X"CD",X"63",
		X"21",X"1C",X"1C",X"CD",X"4D",X"21",X"C9",X"0E",X"02",X"CD",X"63",X"21",X"1D",X"1D",X"CD",X"4D",
		X"21",X"0C",X"CD",X"63",X"21",X"1D",X"1D",X"CD",X"4D",X"21",X"C9",X"01",X"00",X"04",X"CD",X"63",
		X"21",X"1D",X"1D",X"CD",X"4D",X"21",X"0C",X"10",X"F5",X"3A",X"3F",X"40",X"21",X"45",X"1F",X"4F",
		X"09",X"7E",X"BB",X"CC",X"05",X"1F",X"C9",X"06",X"00",X"CD",X"FF",X"20",X"70",X"0C",X"06",X"18",
		X"06",X"01",X"CD",X"FF",X"20",X"80",X"0B",X"06",X"18",X"06",X"02",X"CD",X"FF",X"20",X"70",X"0A",
		X"02",X"E0",X"06",X"03",X"CD",X"FF",X"20",X"80",X"09",X"02",X"E0",X"06",X"1E",X"16",X"06",X"CD",
		X"ED",X"20",X"04",X"CD",X"ED",X"20",X"11",X"BA",X"1B",X"21",X"7E",X"52",X"CD",X"FB",X"19",X"13",
		X"21",X"9F",X"52",X"CD",X"FB",X"19",X"C9",X"21",X"E3",X"51",X"3E",X"24",X"CD",X"39",X"08",X"21",
		X"E5",X"51",X"3E",X"2C",X"CD",X"39",X"08",X"21",X"23",X"52",X"3E",X"28",X"CD",X"39",X"08",X"21",
		X"25",X"52",X"3E",X"30",X"CD",X"39",X"08",X"11",X"00",X"00",X"0E",X"00",X"06",X"04",X"CD",X"4D",
		X"21",X"0C",X"10",X"FA",X"C9",X"21",X"21",X"1F",X"3A",X"3F",X"40",X"87",X"87",X"5F",X"16",X"00",
		X"19",X"3E",X"FF",X"5E",X"23",X"56",X"12",X"23",X"5E",X"23",X"56",X"12",X"21",X"3F",X"40",X"34",
		X"C9",X"7E",X"52",X"BE",X"51",X"5E",X"52",X"DE",X"51",X"3E",X"52",X"FE",X"51",X"1E",X"52",X"1E",
		X"52",X"9F",X"52",X"9F",X"51",X"7F",X"52",X"BF",X"51",X"5F",X"52",X"DF",X"51",X"3F",X"52",X"FF",
		X"51",X"1F",X"52",X"1F",X"52",X"C8",X"B8",X"A8",X"90",X"78",X"60",X"48",X"30",X"18",X"06",X"0E",
		X"16",X"03",X"CD",X"ED",X"20",X"06",X"10",X"CD",X"ED",X"20",X"11",X"A6",X"1A",X"21",X"2E",X"52",
		X"CD",X"FB",X"19",X"11",X"B2",X"1A",X"21",X"50",X"52",X"CD",X"FB",X"19",X"21",X"70",X"51",X"3A",
		X"09",X"40",X"A7",X"28",X"04",X"36",X"5A",X"18",X"02",X"36",X"59",X"06",X"28",X"CD",X"06",X"1A",
		X"0E",X"0E",X"CD",X"15",X"1A",X"0E",X"10",X"CD",X"15",X"1A",X"01",X"04",X"1A",X"16",X"07",X"3E",
		X"08",X"32",X"00",X"40",X"18",X"FE",X"11",X"2C",X"1A",X"21",X"60",X"53",X"CD",X"FB",X"19",X"11",
		X"45",X"1A",X"21",X"BF",X"53",X"CD",X"FB",X"19",X"C9",X"01",X"0E",X"09",X"16",X"03",X"CD",X"ED",
		X"20",X"04",X"0D",X"20",X"F9",X"C9",X"06",X"20",X"21",X"40",X"42",X"36",X"00",X"23",X"10",X"FB",
		X"C9",X"01",X"E0",X"FF",X"1A",X"A7",X"C8",X"77",X"3E",X"0B",X"32",X"07",X"40",X"3A",X"07",X"40",
		X"A7",X"20",X"FA",X"09",X"13",X"18",X"ED",X"06",X"41",X"CD",X"06",X"1A",X"CD",X"B9",X"06",X"11",
		X"00",X"00",X"0E",X"00",X"CD",X"4D",X"21",X"0E",X"02",X"CD",X"4D",X"21",X"0E",X"04",X"CD",X"4D",
		X"21",X"0C",X"CD",X"4D",X"21",X"3A",X"4C",X"42",X"C6",X"07",X"47",X"3A",X"58",X"42",X"B8",X"28",
		X"1A",X"38",X"0D",X"3E",X"09",X"32",X"01",X"40",X"3A",X"58",X"42",X"B8",X"20",X"FA",X"18",X"0B",
		X"3E",X"0A",X"32",X"01",X"40",X"3A",X"58",X"42",X"B8",X"20",X"FA",X"3A",X"47",X"42",X"C6",X"0B",
		X"47",X"3E",X"0B",X"32",X"01",X"40",X"3E",X"01",X"32",X"68",X"40",X"3A",X"5B",X"42",X"B8",X"20",
		X"FA",X"3E",X"01",X"32",X"44",X"40",X"AF",X"32",X"68",X"40",X"32",X"01",X"40",X"06",X"96",X"CD",
		X"06",X"1A",X"CD",X"B6",X"1F",X"06",X"01",X"CD",X"06",X"1A",X"06",X"0F",X"16",X"03",X"CD",X"ED",
		X"20",X"06",X"11",X"CD",X"ED",X"20",X"11",X"5F",X"1A",X"21",X"8F",X"52",X"CD",X"FB",X"19",X"11",
		X"68",X"1B",X"21",X"11",X"52",X"CD",X"FB",X"19",X"11",X"00",X"05",X"CD",X"D4",X"06",X"06",X"41",
		X"CD",X"06",X"1A",X"21",X"F3",X"40",X"3A",X"09",X"40",X"B7",X"28",X"03",X"21",X"33",X"41",X"3E",
		X"07",X"BE",X"28",X"01",X"34",X"3E",X"13",X"32",X"00",X"40",X"18",X"FE",X"0E",X"06",X"CD",X"63",
		X"21",X"15",X"CD",X"4D",X"21",X"0E",X"07",X"CD",X"63",X"21",X"15",X"CD",X"4D",X"21",X"C9",X"0E",
		X"06",X"CD",X"63",X"21",X"14",X"CD",X"4D",X"21",X"0E",X"07",X"CD",X"63",X"21",X"14",X"CD",X"4D",
		X"21",X"C9",X"0E",X"06",X"CD",X"63",X"21",X"1D",X"CD",X"4D",X"21",X"0E",X"07",X"CD",X"63",X"21",
		X"1D",X"CD",X"4D",X"21",X"C9",X"06",X"80",X"21",X"00",X"42",X"36",X"00",X"23",X"10",X"FB",X"C9",
		X"06",X"20",X"21",X"00",X"42",X"36",X"00",X"23",X"23",X"10",X"FA",X"C9",X"F5",X"E5",X"D5",X"78",
		X"87",X"5F",X"16",X"00",X"21",X"00",X"42",X"19",X"D1",X"72",X"E1",X"F1",X"C9",X"F5",X"E5",X"D5",
		X"78",X"87",X"3C",X"5F",X"16",X"00",X"21",X"00",X"42",X"19",X"D1",X"72",X"E1",X"F1",X"C9",X"F5",
		X"C5",X"D5",X"E5",X"21",X"40",X"42",X"16",X"00",X"78",X"87",X"87",X"5F",X"19",X"EB",X"21",X"08",
		X"00",X"39",X"D5",X"5E",X"23",X"56",X"EB",X"D1",X"78",X"FE",X"03",X"30",X"18",X"7E",X"F5",X"3A",
		X"09",X"40",X"B7",X"28",X"0B",X"3A",X"00",X"70",X"CB",X"4F",X"20",X"04",X"F1",X"3D",X"18",X"02",
		X"F1",X"3C",X"12",X"18",X"02",X"7E",X"12",X"06",X"03",X"13",X"23",X"7E",X"12",X"10",X"FA",X"23",
		X"EB",X"21",X"08",X"00",X"39",X"73",X"23",X"72",X"E1",X"D1",X"C1",X"F1",X"C9",X"F5",X"DD",X"E5",
		X"D5",X"DD",X"21",X"40",X"42",X"CD",X"B3",X"21",X"D1",X"DD",X"72",X"00",X"DD",X"73",X"03",X"DD",
		X"E1",X"F1",X"C9",X"DD",X"E5",X"F5",X"DD",X"21",X"40",X"42",X"CD",X"B3",X"21",X"DD",X"7E",X"00",
		X"DD",X"B6",X"03",X"28",X"0B",X"DD",X"56",X"00",X"DD",X"5E",X"03",X"F1",X"DD",X"E1",X"37",X"C9",
		X"F1",X"37",X"3F",X"DD",X"E1",X"C9",X"F5",X"DD",X"E5",X"D5",X"C5",X"48",X"DD",X"21",X"60",X"42",
		X"CD",X"B3",X"21",X"C1",X"D1",X"D5",X"3A",X"09",X"40",X"A7",X"28",X"07",X"3A",X"00",X"70",X"CB",
		X"4F",X"28",X"05",X"7B",X"C6",X"05",X"2F",X"5F",X"DD",X"72",X"01",X"DD",X"73",X"03",X"D1",X"DD",
		X"E1",X"F1",X"C9",X"79",X"87",X"87",X"5F",X"16",X"00",X"DD",X"19",X"C9",X"DD",X"E5",X"F5",X"C5",
		X"48",X"DD",X"21",X"60",X"42",X"CD",X"B3",X"21",X"C1",X"DD",X"56",X"01",X"DD",X"5E",X"03",X"3A",
		X"09",X"40",X"B7",X"28",X"07",X"3A",X"00",X"70",X"CB",X"4F",X"28",X"05",X"7B",X"C6",X"05",X"2F",
		X"5F",X"7A",X"B3",X"28",X"05",X"F1",X"DD",X"E1",X"37",X"C9",X"F1",X"DD",X"E1",X"37",X"3F",X"C9",
		X"F0",X"51",X"EF",X"51",X"EE",X"51",X"ED",X"51",X"EC",X"51",X"EB",X"51",X"EA",X"51",X"D0",X"51",
		X"CF",X"51",X"CE",X"51",X"CD",X"51",X"CC",X"51",X"CB",X"51",X"CA",X"51",X"B0",X"51",X"AF",X"51",
		X"AE",X"51",X"AD",X"51",X"AC",X"51",X"AB",X"51",X"AA",X"51",X"8F",X"51",X"8E",X"51",X"8D",X"51",
		X"8C",X"51",X"8B",X"51",X"8A",X"51",X"89",X"51",X"6F",X"51",X"6E",X"51",X"6D",X"51",X"6C",X"51",
		X"6B",X"51",X"6A",X"51",X"69",X"51",X"4F",X"51",X"4E",X"51",X"4D",X"51",X"4C",X"51",X"4B",X"51",
		X"4A",X"51",X"49",X"51",X"2F",X"51",X"2E",X"51",X"2D",X"51",X"2C",X"51",X"2B",X"51",X"2A",X"51",
		X"29",X"51",X"28",X"51",X"0E",X"51",X"0D",X"51",X"0C",X"51",X"0B",X"51",X"0A",X"51",X"09",X"51",
		X"08",X"51",X"ED",X"50",X"EC",X"50",X"EB",X"50",X"EA",X"50",X"E9",X"50",X"E8",X"50",X"CC",X"50",
		X"CB",X"50",X"CA",X"50",X"C9",X"50",X"C8",X"50",X"C7",X"50",X"AB",X"50",X"AA",X"50",X"A9",X"50",
		X"A8",X"50",X"A7",X"50",X"8A",X"50",X"89",X"50",X"88",X"50",X"87",X"50",X"69",X"50",X"68",X"50",
		X"67",X"50",X"48",X"50",X"47",X"50",X"10",X"52",X"0F",X"52",X"0E",X"52",X"0D",X"52",X"0C",X"52",
		X"0B",X"52",X"0A",X"52",X"30",X"52",X"2F",X"52",X"2E",X"52",X"2D",X"52",X"2C",X"52",X"2B",X"52",
		X"2A",X"52",X"50",X"52",X"4F",X"52",X"4E",X"52",X"4D",X"52",X"4C",X"52",X"4B",X"52",X"4A",X"52",
		X"6F",X"52",X"6E",X"52",X"6D",X"52",X"6C",X"52",X"6B",X"52",X"6A",X"52",X"69",X"52",X"8F",X"52",
		X"8E",X"52",X"8D",X"52",X"8C",X"52",X"8B",X"52",X"8A",X"52",X"89",X"52",X"AF",X"52",X"AE",X"52",
		X"AD",X"52",X"AC",X"52",X"AB",X"52",X"AA",X"52",X"A9",X"52",X"CF",X"52",X"CE",X"52",X"CD",X"52",
		X"CC",X"52",X"CB",X"52",X"CA",X"52",X"C9",X"52",X"C8",X"52",X"EE",X"52",X"ED",X"52",X"EC",X"52",
		X"EB",X"52",X"EA",X"52",X"E9",X"52",X"E8",X"52",X"0D",X"53",X"0C",X"53",X"0B",X"53",X"0A",X"53",
		X"09",X"53",X"08",X"53",X"2C",X"53",X"2B",X"53",X"2A",X"53",X"29",X"53",X"28",X"53",X"27",X"53",
		X"4B",X"53",X"4A",X"53",X"49",X"53",X"48",X"53",X"47",X"53",X"6A",X"53",X"69",X"53",X"68",X"53",
		X"67",X"53",X"89",X"53",X"88",X"53",X"87",X"53",X"A8",X"53",X"A7",X"53",X"F5",X"D5",X"DD",X"E5",
		X"DD",X"21",X"F0",X"21",X"59",X"16",X"00",X"EB",X"29",X"EB",X"DD",X"19",X"DD",X"6E",X"00",X"DD",
		X"66",X"01",X"3A",X"0D",X"40",X"5F",X"16",X"00",X"19",X"DD",X"E1",X"D1",X"F1",X"C9",X"E5",X"16",
		X"00",X"59",X"21",X"50",X"41",X"19",X"3A",X"09",X"40",X"A7",X"7E",X"28",X"08",X"E6",X"F0",X"0F",
		X"0F",X"0F",X"0F",X"18",X"02",X"E6",X"0F",X"A7",X"28",X"07",X"CD",X"3C",X"23",X"CD",X"5B",X"24",
		X"37",X"E1",X"C9",X"FF",X"08",X"01",X"07",X"03",X"05",X"04",X"03",X"04",X"01",X"04",X"FF",X"02",
		X"FD",X"00",X"FB",X"FE",X"FC",X"FC",X"FE",X"FB",X"00",X"FB",X"02",X"FB",X"04",X"FD",X"06",X"00",
		X"05",X"02",X"04",X"03",X"02",X"03",X"00",X"01",X"FE",X"FF",X"FE",X"FD",X"FF",X"FC",X"01",X"FC",
		X"03",X"FE",X"05",X"00",X"08",X"02",X"06",X"04",X"04",X"04",X"02",X"04",X"00",X"03",X"FE",X"01",
		X"FC",X"FF",X"FB",X"FD",X"FD",X"FB",X"FF",X"FB",X"01",X"FB",X"03",X"FC",X"05",X"FE",X"07",X"00",
		X"05",X"02",X"04",X"03",X"02",X"03",X"00",X"01",X"FE",X"FF",X"FE",X"FD",X"FF",X"FC",X"01",X"FC",
		X"03",X"FE",X"05",X"E5",X"21",X"C0",X"40",X"3A",X"09",X"40",X"5F",X"16",X"00",X"19",X"59",X"19",
		X"7E",X"3C",X"20",X"03",X"A7",X"E1",X"C9",X"21",X"83",X"23",X"3A",X"7E",X"40",X"5F",X"19",X"79",
		X"87",X"5F",X"19",X"7E",X"5F",X"3A",X"70",X"40",X"83",X"87",X"87",X"87",X"5F",X"23",X"7E",X"57",
		X"3A",X"71",X"40",X"82",X"87",X"87",X"87",X"57",X"37",X"E1",X"C9",X"F5",X"DD",X"E5",X"D5",X"DD",
		X"21",X"42",X"42",X"CD",X"B3",X"21",X"D1",X"DD",X"70",X"00",X"DD",X"E1",X"F1",X"C9",X"F5",X"D5",
		X"C5",X"7A",X"C6",X"04",X"57",X"CB",X"3A",X"CB",X"3A",X"CB",X"3A",X"3E",X"1F",X"92",X"26",X"00",
		X"6F",X"06",X"05",X"29",X"10",X"FD",X"7B",X"C6",X"04",X"5F",X"CB",X"3B",X"CB",X"3B",X"CB",X"3B",
		X"16",X"00",X"19",X"11",X"00",X"50",X"19",X"C1",X"D1",X"F1",X"C9",X"F5",X"C5",X"E5",X"11",X"00",
		X"50",X"A7",X"ED",X"52",X"E5",X"7D",X"E6",X"1F",X"5F",X"D5",X"21",X"00",X"42",X"87",X"5F",X"16",
		X"00",X"19",X"7E",X"D1",X"F5",X"7B",X"87",X"87",X"87",X"5F",X"06",X"05",X"F1",X"E1",X"E5",X"F5",
		X"CB",X"3C",X"CB",X"1D",X"10",X"FA",X"3E",X"1F",X"95",X"87",X"87",X"87",X"57",X"F1",X"82",X"57",
		X"E1",X"E1",X"C1",X"F1",X"C9",X"E5",X"C5",X"21",X"00",X"50",X"01",X"00",X"04",X"36",X"FF",X"0D",
		X"23",X"20",X"FA",X"10",X"F8",X"C1",X"E1",X"C9",X"C5",X"E5",X"47",X"CD",X"B7",X"24",X"90",X"28",
		X"03",X"30",X"FB",X"80",X"E1",X"C1",X"C9",X"21",X"91",X"40",X"3A",X"91",X"40",X"4F",X"CB",X"27",
		X"CB",X"27",X"81",X"3C",X"32",X"91",X"40",X"C9",X"CD",X"A8",X"24",X"FE",X"FF",X"28",X"01",X"3C",
		X"C9",X"21",X"34",X"42",X"7E",X"C6",X"78",X"67",X"2E",X"D0",X"C9",X"21",X"58",X"42",X"7E",X"67",
		X"2E",X"D0",X"C9",X"21",X"0A",X"42",X"7E",X"C6",X"70",X"67",X"2E",X"28",X"C9",X"21",X"40",X"42",
		X"78",X"87",X"87",X"4F",X"06",X"00",X"09",X"46",X"23",X"7E",X"23",X"23",X"4E",X"E6",X"3F",X"C9",
		X"C1",X"E1",X"F1",X"37",X"C9",X"C1",X"E1",X"F1",X"37",X"3F",X"C9",X"CD",X"D1",X"24",X"78",X"C6",
		X"0C",X"94",X"DA",X"05",X"25",X"D6",X"18",X"D2",X"05",X"25",X"79",X"C6",X"05",X"95",X"DA",X"05",
		X"25",X"D6",X"15",X"D2",X"05",X"25",X"C3",X"00",X"25",X"CD",X"DB",X"24",X"C3",X"0E",X"25",X"CD",
		X"D1",X"24",X"78",X"C6",X"04",X"94",X"DA",X"05",X"25",X"D6",X"10",X"D2",X"05",X"25",X"79",X"C6",
		X"07",X"95",X"DA",X"05",X"25",X"D6",X"20",X"D2",X"05",X"25",X"C3",X"00",X"25",X"CD",X"DB",X"24",
		X"C3",X"32",X"25",X"D5",X"CD",X"BC",X"21",X"7A",X"4B",X"D1",X"D2",X"05",X"25",X"D6",X"06",X"94",
		X"DA",X"05",X"25",X"D6",X"0A",X"D2",X"05",X"25",X"79",X"D6",X"13",X"95",X"DA",X"05",X"25",X"D6",
		X"0F",X"D2",X"05",X"25",X"C3",X"00",X"25",X"D5",X"CD",X"BC",X"21",X"7A",X"4B",X"D1",X"D2",X"05",
		X"25",X"94",X"DA",X"05",X"25",X"D6",X"1E",X"D2",X"05",X"25",X"79",X"C6",X"07",X"95",X"DA",X"05",
		X"25",X"D6",X"15",X"D2",X"05",X"25",X"C3",X"00",X"25",X"D5",X"CD",X"BC",X"21",X"7A",X"4B",X"D1",
		X"D2",X"05",X"25",X"94",X"DA",X"05",X"25",X"D6",X"0E",X"D2",X"05",X"25",X"79",X"C6",X"07",X"95",
		X"DA",X"05",X"25",X"D6",X"15",X"D2",X"05",X"25",X"C3",X"00",X"25",X"D5",X"CD",X"BC",X"21",X"7A",
		X"4B",X"D1",X"D2",X"05",X"25",X"94",X"DA",X"05",X"25",X"D6",X"0A",X"D2",X"05",X"25",X"79",X"C6",
		X"07",X"95",X"DA",X"05",X"25",X"D6",X"0D",X"D2",X"05",X"25",X"C3",X"00",X"25",X"F5",X"E5",X"C5",
		X"CD",X"ED",X"24",X"FE",X"02",X"CA",X"0B",X"25",X"C3",X"05",X"25",X"F5",X"E5",X"C5",X"CD",X"ED",
		X"24",X"FE",X"01",X"CA",X"29",X"25",X"FE",X"37",X"CA",X"29",X"25",X"C3",X"05",X"25",X"F5",X"E5",
		X"C5",X"D5",X"48",X"CD",X"5E",X"23",X"42",X"4B",X"D1",X"D2",X"05",X"25",X"C3",X"4D",X"25",X"F5",
		X"E5",X"C5",X"D5",X"48",X"CD",X"E3",X"23",X"42",X"4B",X"D1",X"D2",X"05",X"25",X"C3",X"4D",X"25",
		X"F5",X"E5",X"C5",X"CD",X"DB",X"24",X"C3",X"53",X"25",X"F5",X"E5",X"C5",X"CD",X"E3",X"24",X"C3",
		X"77",X"25",X"F5",X"E5",X"C5",X"06",X"02",X"CD",X"ED",X"24",X"60",X"69",X"FE",X"0C",X"C2",X"05",
		X"25",X"C1",X"C5",X"C3",X"77",X"25",X"F5",X"E5",X"C5",X"D5",X"CD",X"00",X"09",X"62",X"6B",X"D1",
		X"D2",X"05",X"25",X"C3",X"99",X"25",X"F5",X"E5",X"C5",X"D5",X"CD",X"00",X"09",X"62",X"6B",X"D1",
		X"D2",X"05",X"25",X"C3",X"99",X"25",X"F5",X"E5",X"C5",X"41",X"CD",X"ED",X"24",X"FE",X"02",X"28",
		X"03",X"C3",X"05",X"25",X"60",X"69",X"C1",X"C5",X"C3",X"99",X"25",X"F5",X"E5",X"C5",X"D5",X"CD",
		X"00",X"09",X"62",X"6B",X"D1",X"D2",X"05",X"25",X"C3",X"99",X"25",X"F5",X"E5",X"C5",X"41",X"CD",
		X"ED",X"24",X"FE",X"01",X"28",X"07",X"FE",X"37",X"28",X"03",X"C3",X"05",X"25",X"60",X"69",X"C1",
		X"C5",X"C3",X"99",X"25",X"F5",X"E5",X"C5",X"D5",X"CD",X"5E",X"23",X"62",X"6B",X"D1",X"D2",X"05",
		X"25",X"C3",X"BB",X"25",X"F5",X"E5",X"C5",X"D5",X"CD",X"E3",X"23",X"62",X"6B",X"D1",X"D2",X"05",
		X"25",X"C3",X"BB",X"25",X"F5",X"C5",X"E5",X"DD",X"E5",X"21",X"FF",X"FF",X"22",X"06",X"68",X"DD",
		X"21",X"30",X"40",X"DD",X"CB",X"00",X"46",X"28",X"13",X"3E",X"03",X"DD",X"77",X"01",X"21",X"05",
		X"68",X"DD",X"75",X"03",X"DD",X"74",X"04",X"CD",X"E1",X"27",X"18",X"04",X"AF",X"32",X"05",X"68",
		X"DD",X"21",X"35",X"40",X"DD",X"CB",X"00",X"46",X"28",X"10",X"3E",X"08",X"DD",X"77",X"01",X"21",
		X"03",X"68",X"DD",X"75",X"03",X"DD",X"74",X"04",X"18",X"18",X"DD",X"21",X"3A",X"40",X"DD",X"CB",
		X"00",X"46",X"28",X"14",X"3E",X"0C",X"DD",X"77",X"01",X"21",X"03",X"68",X"DD",X"75",X"03",X"DD",
		X"74",X"04",X"CD",X"E1",X"27",X"C3",X"2C",X"27",X"AF",X"32",X"03",X"68",X"DD",X"21",X"40",X"40",
		X"DD",X"CB",X"00",X"46",X"28",X"06",X"21",X"CB",X"28",X"C3",X"D1",X"27",X"DD",X"21",X"44",X"40",
		X"DD",X"CB",X"00",X"46",X"28",X"06",X"21",X"08",X"29",X"C3",X"D1",X"27",X"DD",X"21",X"48",X"40",
		X"DD",X"CB",X"00",X"46",X"28",X"05",X"21",X"1C",X"29",X"18",X"76",X"DD",X"21",X"4C",X"40",X"DD",
		X"CB",X"00",X"46",X"28",X"05",X"21",X"35",X"29",X"18",X"67",X"DD",X"21",X"50",X"40",X"DD",X"CB",
		X"00",X"46",X"28",X"05",X"21",X"5C",X"29",X"18",X"58",X"DD",X"21",X"54",X"40",X"DD",X"CB",X"00",
		X"46",X"28",X"05",X"21",X"6A",X"29",X"18",X"49",X"DD",X"21",X"68",X"40",X"DD",X"CB",X"00",X"46",
		X"28",X"05",X"21",X"C4",X"29",X"18",X"3A",X"DD",X"21",X"58",X"40",X"DD",X"CB",X"00",X"46",X"28",
		X"05",X"21",X"78",X"29",X"18",X"2B",X"DD",X"21",X"5C",X"40",X"DD",X"CB",X"00",X"46",X"28",X"05",
		X"21",X"8D",X"29",X"18",X"1C",X"DD",X"21",X"60",X"40",X"DD",X"CB",X"00",X"46",X"28",X"05",X"21",
		X"9A",X"29",X"18",X"0D",X"DD",X"21",X"64",X"40",X"DD",X"CB",X"00",X"46",X"28",X"08",X"21",X"B3",
		X"29",X"CD",X"0B",X"28",X"18",X"05",X"3E",X"FF",X"32",X"00",X"78",X"DD",X"E1",X"E1",X"C1",X"F1",
		X"C9",X"DD",X"CB",X"00",X"4E",X"20",X"14",X"DD",X"CB",X"00",X"CE",X"DD",X"7E",X"01",X"DD",X"77",
		X"02",X"DD",X"6E",X"03",X"DD",X"66",X"04",X"3E",X"FF",X"77",X"C9",X"DD",X"35",X"02",X"C0",X"DD",
		X"6E",X"03",X"DD",X"66",X"04",X"AF",X"77",X"DD",X"77",X"00",X"C9",X"DD",X"CB",X"00",X"4E",X"20",
		X"3A",X"DD",X"CB",X"00",X"CE",X"DD",X"75",X"01",X"DD",X"74",X"02",X"DD",X"6E",X"01",X"DD",X"66",
		X"02",X"7E",X"23",X"DD",X"75",X"01",X"DD",X"74",X"02",X"FE",X"FF",X"28",X"24",X"F5",X"21",X"AB",
		X"28",X"E6",X"1F",X"4F",X"06",X"00",X"09",X"7E",X"32",X"00",X"78",X"F1",X"E6",X"E0",X"CB",X"3F",
		X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"3C",X"DD",X"77",X"03",X"C9",X"DD",X"35",X"03",X"28",X"CB",
		X"C9",X"AF",X"DD",X"77",X"00",X"2F",X"32",X"00",X"78",X"C9",X"DD",X"CB",X"00",X"4E",X"20",X"1E",
		X"DD",X"CB",X"00",X"CE",X"DD",X"75",X"01",X"DD",X"74",X"02",X"AF",X"DD",X"77",X"04",X"3E",X"A0",
		X"DD",X"77",X"05",X"DD",X"36",X"06",X"01",X"DD",X"7E",X"05",X"32",X"00",X"78",X"C9",X"DD",X"CB",
		X"04",X"46",X"20",X"23",X"DD",X"7E",X"06",X"3D",X"DD",X"77",X"06",X"C0",X"DD",X"7E",X"05",X"3D",
		X"DD",X"77",X"05",X"FE",X"55",X"20",X"DC",X"3E",X"FF",X"DD",X"77",X"04",X"2F",X"DD",X"CB",X"00",
		X"8E",X"DD",X"6E",X"01",X"DD",X"66",X"02",X"CD",X"0B",X"28",X"C9",X"00",X"0E",X"1B",X"28",X"34",
		X"40",X"4A",X"55",X"5E",X"67",X"70",X"78",X"80",X"87",X"8D",X"94",X"9A",X"A0",X"A5",X"AA",X"AF",
		X"B3",X"B8",X"BC",X"C0",X"C3",X"C6",X"CA",X"CD",X"D0",X"D2",X"FF",X"31",X"30",X"2B",X"27",X"30",
		X"2C",X"29",X"25",X"2E",X"2A",X"27",X"24",X"2C",X"29",X"25",X"22",X"20",X"22",X"24",X"25",X"22",
		X"24",X"25",X"27",X"24",X"25",X"27",X"29",X"25",X"27",X"29",X"2A",X"27",X"29",X"2A",X"2C",X"2A",
		X"2C",X"2E",X"30",X"28",X"2A",X"2C",X"2E",X"2A",X"2C",X"2E",X"30",X"2C",X"2E",X"30",X"31",X"2C",
		X"2E",X"30",X"31",X"2C",X"2E",X"30",X"91",X"FF",X"EC",X"CB",X"47",X"89",X"87",X"85",X"84",X"E0",
		X"84",X"42",X"44",X"E2",X"40",X"42",X"44",X"45",X"47",X"49",X"EB",X"FF",X"30",X"3F",X"30",X"3F",
		X"30",X"3F",X"30",X"3F",X"32",X"3F",X"32",X"3F",X"32",X"3F",X"32",X"3F",X"30",X"3F",X"30",X"3F",
		X"30",X"3F",X"30",X"3F",X"FF",X"67",X"EB",X"0B",X"09",X"07",X"05",X"04",X"02",X"0B",X"09",X"07",
		X"05",X"04",X"02",X"0B",X"09",X"07",X"05",X"04",X"02",X"0B",X"09",X"07",X"05",X"04",X"02",X"0B",
		X"09",X"07",X"05",X"04",X"02",X"0B",X"09",X"07",X"05",X"04",X"02",X"FF",X"00",X"0C",X"00",X"00",
		X"0C",X"00",X"00",X"01",X"03",X"05",X"07",X"09",X"0B",X"FF",X"00",X"0C",X"00",X"00",X"0C",X"00",
		X"00",X"01",X"03",X"05",X"07",X"09",X"0B",X"FF",X"00",X"02",X"04",X"05",X"07",X"04",X"06",X"08",
		X"09",X"0B",X"07",X"09",X"0B",X"0C",X"0E",X"0C",X"0E",X"10",X"11",X"13",X"FF",X"03",X"05",X"0B",
		X"03",X"05",X"0B",X"03",X"05",X"0B",X"03",X"05",X"0B",X"FF",X"04",X"05",X"07",X"09",X"0B",X"1F",
		X"0B",X"1F",X"0B",X"1F",X"0B",X"1F",X"0C",X"0E",X"10",X"11",X"10",X"1F",X"10",X"1F",X"10",X"1F",
		X"10",X"1F",X"FF",X"0A",X"09",X"08",X"07",X"0A",X"09",X"08",X"07",X"0A",X"09",X"08",X"07",X"0A",
		X"09",X"08",X"07",X"FF",X"90",X"87",X"89",X"80",X"90",X"87",X"89",X"80",X"90",X"87",X"89",X"80",
		X"90",X"87",X"89",X"80",X"90",X"87",X"89",X"80",X"90",X"87",X"89",X"80",X"90",X"87",X"89",X"80",
		X"90",X"87",X"89",X"80",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
