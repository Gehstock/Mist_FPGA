library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity berzerk_program2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of berzerk_program2 is
	type rom is array(0 to  10239) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"10",X"D1",X"10",X"DE",X"10",X"EB",X"10",X"F8",X"10",X"F8",X"10",X"F8",X"11",X"05",X"11",X"12",
		X"00",X"00",X"10",X"11",X"2C",X"11",X"1F",X"11",X"1F",X"00",X"13",X"10",X"10",X"D1",X"11",X"39",
		X"10",X"D1",X"11",X"47",X"00",X"1C",X"10",X"11",X"55",X"11",X"62",X"11",X"62",X"00",X"27",X"10",
		X"11",X"6F",X"11",X"7C",X"11",X"6F",X"11",X"8A",X"00",X"30",X"10",X"11",X"98",X"11",X"BC",X"11",
		X"E0",X"12",X"08",X"00",X"41",X"10",X"10",X"BF",X"00",X"46",X"10",X"10",X"AD",X"10",X"9B",X"10",
		X"89",X"10",X"9B",X"00",X"4B",X"10",X"13",X"B5",X"13",X"A3",X"13",X"91",X"13",X"A3",X"00",X"56",
		X"10",X"13",X"09",X"00",X"61",X"10",X"13",X"1A",X"00",X"66",X"10",X"13",X"2B",X"00",X"6B",X"10",
		X"13",X"3C",X"00",X"70",X"10",X"13",X"4D",X"00",X"75",X"10",X"13",X"5E",X"00",X"7A",X"10",X"13",
		X"6F",X"00",X"7F",X"10",X"13",X"80",X"00",X"84",X"10",X"01",X"10",X"18",X"18",X"00",X"3C",X"5A",
		X"99",X"58",X"18",X"18",X"24",X"22",X"41",X"41",X"81",X"81",X"00",X"01",X"10",X"00",X"18",X"18",
		X"00",X"3C",X"5C",X"5C",X"3E",X"18",X"18",X"14",X"12",X"F2",X"82",X"02",X"03",X"01",X"10",X"18",
		X"18",X"00",X"3C",X"5C",X"5C",X"5A",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"1C",X"10",X"01",
		X"10",X"18",X"18",X"00",X"3C",X"5A",X"5A",X"5A",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"1C",
		X"10",X"01",X"0B",X"3C",X"66",X"FF",X"BD",X"BD",X"BD",X"3C",X"24",X"24",X"24",X"66",X"01",X"0B",
		X"3C",X"4E",X"FF",X"BD",X"BD",X"BD",X"3C",X"24",X"24",X"24",X"66",X"01",X"0B",X"3C",X"1E",X"FF",
		X"BD",X"BD",X"BD",X"3C",X"24",X"24",X"24",X"66",X"01",X"0B",X"3C",X"7E",X"FF",X"BD",X"BD",X"BD",
		X"3C",X"24",X"24",X"24",X"66",X"01",X"0B",X"3C",X"78",X"FF",X"BD",X"BD",X"BD",X"3C",X"24",X"24",
		X"24",X"66",X"01",X"0B",X"3C",X"71",X"FF",X"BD",X"BD",X"BD",X"3C",X"24",X"24",X"24",X"66",X"01",
		X"0B",X"3C",X"78",X"FF",X"BD",X"BD",X"BD",X"3C",X"18",X"18",X"18",X"1C",X"01",X"0B",X"3C",X"78",
		X"FF",X"BD",X"BD",X"BD",X"3C",X"24",X"24",X"24",X"36",X"01",X"0C",X"3C",X"66",X"FF",X"BD",X"BD",
		X"BD",X"3C",X"24",X"24",X"26",X"20",X"60",X"01",X"0C",X"3C",X"66",X"FF",X"BD",X"BD",X"BD",X"3C",
		X"24",X"24",X"64",X"04",X"06",X"01",X"0B",X"3C",X"1E",X"FF",X"BD",X"BD",X"BD",X"3C",X"24",X"24",
		X"24",X"6C",X"01",X"0B",X"3C",X"1E",X"FF",X"BD",X"BD",X"BD",X"3C",X"18",X"18",X"18",X"38",X"01",
		X"0B",X"3C",X"7E",X"FF",X"BD",X"BD",X"BD",X"3C",X"24",X"24",X"24",X"66",X"01",X"0C",X"3C",X"7E",
		X"FF",X"BD",X"BD",X"BD",X"3C",X"24",X"24",X"26",X"20",X"60",X"01",X"0C",X"3C",X"7E",X"FF",X"BD",
		X"BD",X"BD",X"3C",X"24",X"24",X"64",X"04",X"06",X"02",X"11",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"C0",X"07",X"E0",X"0F",X"F0",X"13",X"C8",X"22",X"C4",
		X"03",X"40",X"03",X"C0",X"02",X"40",X"02",X"40",X"02",X"40",X"06",X"60",X"02",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"C0",X"06",X"60",X"12",X"48",X"08",X"10",X"10",X"08",
		X"22",X"44",X"44",X"42",X"02",X"10",X"03",X"C0",X"02",X"40",X"04",X"20",X"02",X"40",X"06",X"60",
		X"02",X"13",X"00",X"00",X"02",X"00",X"00",X"40",X"00",X"08",X"10",X"00",X"03",X"00",X"00",X"12",
		X"08",X"01",X"80",X"00",X"08",X"02",X"40",X"02",X"04",X"10",X"23",X"C0",X"40",X"04",X"20",X"02",
		X"00",X"00",X"80",X"00",X"10",X"08",X"18",X"0C",X"01",X"01",X"00",X"12",X"2E",X"12",X"34",X"12",
		X"3B",X"12",X"43",X"12",X"4C",X"12",X"56",X"12",X"A7",X"12",X"6D",X"12",X"79",X"12",X"85",X"12",
		X"91",X"12",X"9D",X"12",X"91",X"12",X"85",X"12",X"79",X"12",X"6D",X"00",X"17",X"12",X"84",X"00",
		X"01",X"02",X"18",X"18",X"84",X"00",X"01",X"03",X"10",X"38",X"10",X"84",X"00",X"01",X"04",X"18",
		X"3C",X"3C",X"18",X"84",X"00",X"01",X"05",X"38",X"7C",X"7C",X"7C",X"38",X"84",X"00",X"01",X"06",
		X"3C",X"7E",X"7E",X"7E",X"7E",X"3C",X"84",X"00",X"01",X"07",X"38",X"7C",X"FE",X"FE",X"FE",X"7C",
		X"38",X"84",X"00",X"01",X"08",X"3C",X"7E",X"FF",X"FF",X"FF",X"FF",X"7E",X"3C",X"82",X"00",X"01",
		X"08",X"3C",X"7E",X"DB",X"FF",X"FF",X"BD",X"42",X"3C",X"81",X"00",X"01",X"08",X"3C",X"7E",X"DB",
		X"FF",X"FF",X"BD",X"42",X"3C",X"80",X"80",X"01",X"08",X"3C",X"7E",X"DB",X"FF",X"FF",X"BD",X"42",
		X"3C",X"80",X"40",X"01",X"08",X"3C",X"7E",X"DB",X"FF",X"FF",X"BD",X"42",X"3C",X"01",X"08",X"3C",
		X"7E",X"DB",X"FF",X"FF",X"BD",X"42",X"3C",X"84",X"00",X"01",X"08",X"00",X"00",X"00",X"3C",X"7E",
		X"DB",X"FF",X"7E",X"12",X"D0",X"12",X"BE",X"12",X"E3",X"12",X"F6",X"00",X"B3",X"12",X"01",X"10",
		X"00",X"18",X"18",X"00",X"3C",X"5A",X"5A",X"5A",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"3C",
		X"01",X"11",X"18",X"24",X"24",X"42",X"81",X"81",X"81",X"81",X"81",X"42",X"24",X"24",X"24",X"24",
		X"24",X"42",X"3C",X"01",X"11",X"3C",X"24",X"24",X"7E",X"C3",X"A5",X"A5",X"A5",X"E7",X"66",X"24",
		X"24",X"24",X"24",X"66",X"42",X"7E",X"01",X"11",X"3C",X"3C",X"3C",X"7E",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"7E",X"3C",X"3C",X"3C",X"3C",X"7E",X"7E",X"7E",X"01",X"0F",X"18",X"19",X"04",X"1C",X"18",
		X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"1C",X"01",X"0F",X"18",X"18",X"00",X"1F",
		X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"1C",X"01",X"0F",X"18",X"18",X"00",
		X"18",X"18",X"1C",X"1A",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"1C",X"01",X"0F",X"18",X"18",
		X"00",X"3C",X"3C",X"3A",X"3A",X"3A",X"18",X"18",X"18",X"18",X"18",X"18",X"1C",X"01",X"0F",X"18",
		X"18",X"00",X"3C",X"3C",X"5C",X"9C",X"1C",X"18",X"18",X"18",X"18",X"18",X"18",X"38",X"01",X"0F",
		X"18",X"18",X"00",X"F8",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"38",X"01",
		X"0F",X"98",X"58",X"20",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"38",
		X"01",X"0F",X"18",X"18",X"00",X"1D",X"1B",X"19",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",
		X"38",X"01",X"10",X"18",X"18",X"00",X"3C",X"5A",X"99",X"9A",X"18",X"18",X"24",X"44",X"42",X"42",
		X"41",X"41",X"80",X"01",X"10",X"00",X"18",X"18",X"00",X"3C",X"3A",X"3A",X"7C",X"18",X"18",X"28",
		X"48",X"4F",X"41",X"40",X"80",X"01",X"10",X"18",X"18",X"00",X"3C",X"3A",X"3A",X"7A",X"18",X"18",
		X"18",X"18",X"18",X"18",X"18",X"18",X"38",X"72",X"20",X"62",X"6F",X"75",X"74",X"6F",X"6E",X"20",
		X"73",X"74",X"61",X"72",X"74",X"20",X"31",X"20",X"6F",X"75",X"20",X"32",X"00",X"C9",X"CD",X"7B",
		X"29",X"90",X"20",X"BE",X"53",X"74",X"61",X"72",X"74",X"6B",X"6E",X"6F",X"65",X"70",X"66",X"65",
		X"20",X"64",X"72",X"75",X"65",X"63",X"6B",X"65",X"6E",X"00",X"C9",X"CD",X"7B",X"29",X"90",X"44",
		X"BE",X"50",X"75",X"6C",X"73",X"61",X"72",X"20",X"53",X"74",X"61",X"72",X"74",X"00",X"C9",X"CD",
		X"7B",X"29",X"90",X"58",X"BE",X"49",X"6E",X"73",X"65",X"72",X"74",X"20",X"43",X"6F",X"69",X"6E",
		X"00",X"C9",X"CD",X"7B",X"29",X"90",X"30",X"BE",X"49",X"6E",X"74",X"72",X"6F",X"64",X"75",X"69",
		X"72",X"65",X"20",X"6C",X"61",X"20",X"6D",X"6F",X"6E",X"6E",X"61",X"69",X"65",X"00",X"C9",X"CD",
		X"7B",X"29",X"90",X"48",X"BE",X"4D",X"75",X"6E",X"7A",X"65",X"20",X"65",X"69",X"6E",X"77",X"65",
		X"72",X"66",X"65",X"6E",X"00",X"C9",X"CD",X"7B",X"29",X"90",X"48",X"BE",X"50",X"6F",X"6E",X"67",
		X"61",X"20",X"6C",X"61",X"20",X"6D",X"6F",X"6E",X"65",X"64",X"61",X"00",X"C9",X"00",X"C5",X"F5",
		X"FD",X"2A",X"76",X"08",X"FD",X"66",X"07",X"FD",X"6E",X"09",X"CD",X"E7",X"1C",X"D5",X"DD",X"66",
		X"07",X"DD",X"6E",X"09",X"2D",X"2D",X"2D",X"2D",X"25",X"25",X"25",X"25",X"CD",X"E7",X"1C",X"D9",
		X"47",X"D9",X"C1",X"79",X"BB",X"20",X"03",X"F1",X"C1",X"C9",X"7C",X"E5",X"C6",X"10",X"67",X"CD",
		X"E7",X"1C",X"D9",X"4F",X"D9",X"7D",X"C6",X"13",X"6F",X"CD",X"E7",X"1C",X"D9",X"57",X"D9",X"7D",
		X"E1",X"6F",X"CD",X"E7",X"1C",X"D9",X"5F",X"F1",X"67",X"2E",X"00",X"CB",X"5C",X"28",X"06",X"78",
		X"B1",X"E6",X"08",X"B5",X"6F",X"CB",X"54",X"28",X"06",X"7A",X"B3",X"E6",X"04",X"B5",X"6F",X"CB",
		X"4C",X"28",X"06",X"78",X"B3",X"E6",X"02",X"B5",X"6F",X"CB",X"44",X"28",X"06",X"79",X"B2",X"E6",
		X"01",X"B5",X"6F",X"2F",X"A4",X"C1",X"C9",X"7D",X"1E",X"00",X"FE",X"46",X"38",X"08",X"1E",X"05",
		X"FE",X"8A",X"EA",X"06",X"02",X"CD",X"05",X"15",X"3A",X"7A",X"43",X"C6",X"02",X"E6",X"07",X"47",
		X"CD",X"05",X"15",X"06",X"07",X"FD",X"21",X"7B",X"43",X"C5",X"FD",X"E5",X"CD",X"1A",X"15",X"FD",
		X"E1",X"C1",X"11",X"08",X"00",X"FD",X"19",X"10",X"F0",X"C9",X"FD",X"7E",X"00",X"B7",X"28",X"0C",
		X"FD",X"34",X"01",X"CD",X"53",X"15",X"DC",X"A0",X"15",X"CD",X"7E",X"15",X"01",X"04",X"00",X"FD",
		X"09",X"FD",X"35",X"01",X"C0",X"FD",X"34",X"01",X"AF",X"FD",X"B6",X"FD",X"C8",X"AF",X"FD",X"B6",
		X"00",X"CA",X"4A",X"15",X"CD",X"53",X"15",X"CD",X"7E",X"15",X"FD",X"35",X"FD",X"C0",X"FD",X"36",
		X"00",X"00",X"C9",X"0F",X"D2",X"5A",X"15",X"FD",X"35",X"02",X"0F",X"D2",X"61",X"15",X"FD",X"34",
		X"02",X"0F",X"D2",X"68",X"15",X"FD",X"35",X"03",X"0F",X"D2",X"6F",X"15",X"FD",X"34",X"03",X"FD",
		X"66",X"03",X"FD",X"6E",X"02",X"CD",X"A1",X"29",X"36",X"80",X"DB",X"4E",X"07",X"C9",X"FD",X"7E",
		X"02",X"FD",X"46",X"00",X"11",X"FF",X"03",X"CD",X"97",X"15",X"FD",X"7E",X"03",X"11",X"D0",X"0C",
		X"CD",X"97",X"15",X"FD",X"70",X"00",X"C9",X"FE",X"00",X"28",X"02",X"BB",X"C0",X"06",X"00",X"C9",
		X"FD",X"36",X"00",X"00",X"DD",X"2A",X"76",X"08",X"CD",X"CB",X"15",X"ED",X"4B",X"70",X"08",X"78",
		X"B1",X"28",X"17",X"C5",X"DD",X"E1",X"CD",X"CB",X"15",X"DD",X"66",X"FF",X"DD",X"6E",X"FE",X"E5",
		X"DD",X"E1",X"7D",X"B9",X"20",X"F0",X"7C",X"B8",X"20",X"EC",X"C9",X"DD",X"CB",X"00",X"56",X"C8",
		X"DD",X"66",X"0B",X"DD",X"6E",X"0A",X"56",X"23",X"5E",X"EB",X"56",X"23",X"5E",X"1C",X"FD",X"7E",
		X"03",X"DD",X"96",X"09",X"3C",X"F8",X"BB",X"D0",X"FD",X"7E",X"02",X"DD",X"96",X"07",X"F8",X"CB",
		X"22",X"CB",X"22",X"CB",X"22",X"14",X"BA",X"D0",X"DD",X"CB",X"00",X"FE",X"DD",X"CB",X"FA",X"C6",
		X"E1",X"C9",X"F3",X"31",X"00",X"43",X"DB",X"60",X"CB",X"4F",X"C2",X"3A",X"07",X"21",X"70",X"08",
		X"06",X"34",X"36",X"00",X"23",X"10",X"FB",X"21",X"00",X"40",X"01",X"00",X"04",X"AF",X"77",X"23",
		X"0D",X"20",X"FB",X"10",X"F9",X"CD",X"21",X"17",X"21",X"DC",X"08",X"11",X"02",X"43",X"06",X"1E",
		X"7E",X"23",X"E6",X"F0",X"4F",X"7E",X"23",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"B1",X"12",X"13",
		X"10",X"EE",X"DB",X"49",X"2F",X"21",X"9F",X"08",X"77",X"23",X"77",X"CD",X"66",X"16",X"CD",X"AC",
		X"19",X"CD",X"8B",X"18",X"CD",X"98",X"1A",X"CD",X"8B",X"18",X"CD",X"85",X"16",X"CA",X"4B",X"16",
		X"CD",X"66",X"16",X"CD",X"B2",X"18",X"F3",X"E1",X"22",X"00",X"44",X"32",X"02",X"44",X"31",X"00",
		X"43",X"CD",X"22",X"1E",X"FD",X"2A",X"72",X"08",X"CD",X"F1",X"22",X"CD",X"AB",X"26",X"2A",X"00",
		X"44",X"3A",X"02",X"44",X"E9",X"2A",X"3E",X"43",X"22",X"73",X"43",X"3A",X"40",X"43",X"32",X"75",
		X"43",X"21",X"00",X"00",X"22",X"3E",X"43",X"22",X"3F",X"43",X"2A",X"5C",X"43",X"E5",X"21",X"D9",
		X"16",X"22",X"6F",X"43",X"3E",X"FF",X"32",X"6E",X"43",X"01",X"0C",X"00",X"11",X"44",X"43",X"21",
		X"CD",X"16",X"ED",X"B0",X"CD",X"9D",X"20",X"E1",X"F5",X"22",X"5C",X"43",X"CD",X"78",X"26",X"2A",
		X"73",X"43",X"22",X"3E",X"43",X"2A",X"74",X"43",X"22",X"3F",X"43",X"F1",X"C9",X"01",X"02",X"02",
		X"1E",X"64",X"01",X"70",X"00",X"01",X"1E",X"02",X"00",X"0A",X"8F",X"12",X"8F",X"14",X"8F",X"19",
		X"8F",X"02",X"9F",X"19",X"8F",X"06",X"8F",X"18",X"8F",X"02",X"FF",X"00",X"FF",X"02",X"FF",X"BF",
		X"08",X"AF",X"09",X"BF",X"01",X"BF",X"09",X"FF",X"09",X"C1",X"12",X"8F",X"00",X"FF",X"01",X"D4",
		X"08",X"BF",X"18",X"BF",X"18",X"8F",X"08",X"FF",X"08",X"B6",X"02",X"C0",X"06",X"9C",X"12",X"8F",
		X"08",X"BF",X"00",X"FF",X"14",X"8F",X"14",X"8F",X"14",X"8F",X"14",X"8F",X"14",X"8F",X"00",X"FF",
		X"FF",X"ED",X"73",X"5E",X"08",X"31",X"5E",X"08",X"F5",X"C5",X"D5",X"E5",X"DD",X"E5",X"DB",X"65",
		X"CB",X"7F",X"C2",X"05",X"06",X"3A",X"6E",X"43",X"B7",X"CC",X"12",X"1D",X"CD",X"76",X"17",X"3A",
		X"6E",X"43",X"B7",X"20",X"1D",X"2A",X"98",X"08",X"7C",X"B5",X"28",X"19",X"DB",X"44",X"E6",X"C0",
		X"FE",X"40",X"20",X"11",X"7E",X"CB",X"7F",X"20",X"09",X"23",X"D3",X"44",X"CB",X"77",X"28",X"05",
		X"18",X"E6",X"21",X"00",X"00",X"22",X"98",X"08",X"DD",X"E1",X"E1",X"D1",X"C1",X"F1",X"ED",X"7B",
		X"5E",X"08",X"D3",X"4C",X"ED",X"45",X"21",X"78",X"08",X"46",X"23",X"56",X"23",X"5E",X"23",X"0E",
		X"41",X"CB",X"80",X"CB",X"C2",X"ED",X"51",X"0D",X"ED",X"41",X"0C",X"CB",X"82",X"ED",X"51",X"0D",
		X"ED",X"59",X"0C",X"0C",X"06",X"03",X"79",X"0C",X"51",X"5E",X"23",X"4F",X"7E",X"23",X"ED",X"79",
		X"79",X"4A",X"ED",X"59",X"14",X"14",X"10",X"F1",X"0D",X"3E",X"00",X"06",X"04",X"B6",X"23",X"ED",
		X"79",X"E6",X"C0",X"C6",X"40",X"10",X"F6",X"C9",X"06",X"06",X"21",X"BE",X"08",X"CD",X"B3",X"2D",
		X"3A",X"76",X"43",X"FE",X"02",X"CC",X"B3",X"2D",X"CD",X"51",X"18",X"01",X"0C",X"00",X"11",X"44",
		X"43",X"21",X"7F",X"18",X"ED",X"B0",X"CD",X"78",X"26",X"2A",X"5C",X"43",X"22",X"45",X"43",X"AF",
		X"32",X"6E",X"43",X"32",X"9A",X"08",X"3C",X"32",X"9B",X"08",X"CD",X"A7",X"33",X"21",X"44",X"43",
		X"11",X"50",X"43",X"01",X"0C",X"00",X"ED",X"B0",X"3E",X"02",X"77",X"3A",X"76",X"43",X"FE",X"02",
		X"28",X"04",X"AF",X"32",X"55",X"43",X"FB",X"21",X"1E",X"64",X"22",X"47",X"43",X"3A",X"44",X"43",
		X"3D",X"28",X"0B",X"DB",X"4A",X"CB",X"7F",X"28",X"05",X"3E",X"E0",X"32",X"47",X"43",X"CD",X"9D",
		X"20",X"CD",X"78",X"26",X"2A",X"5C",X"43",X"22",X"45",X"43",X"3E",X"5A",X"CD",X"6D",X"1E",X"CD",
		X"F1",X"22",X"21",X"49",X"43",X"35",X"08",X"CD",X"6A",X"18",X"7E",X"B7",X"C2",X"06",X"18",X"08",
		X"20",X"F5",X"CD",X"6A",X"18",X"CD",X"51",X"2C",X"CD",X"6A",X"18",X"CD",X"51",X"2C",X"C3",X"4B",
		X"16",X"21",X"00",X"00",X"22",X"3E",X"43",X"22",X"40",X"43",X"22",X"42",X"43",X"22",X"A1",X"08",
		X"22",X"A2",X"08",X"21",X"DB",X"1A",X"22",X"98",X"08",X"C9",X"E5",X"21",X"44",X"43",X"11",X"50",
		X"43",X"06",X"0C",X"1A",X"4E",X"EB",X"12",X"71",X"EB",X"23",X"13",X"10",X"F6",X"E1",X"C9",X"01",
		X"00",X"00",X"1E",X"64",X"03",X"60",X"00",X"05",X"5A",X"00",X"00",X"06",X"03",X"2A",X"72",X"08",
		X"23",X"36",X"3C",X"2B",X"CB",X"CE",X"DB",X"65",X"CB",X"47",X"28",X"04",X"3E",X"01",X"18",X"21",
		X"CD",X"7B",X"19",X"CD",X"97",X"19",X"20",X"0A",X"2A",X"72",X"08",X"CB",X"4E",X"20",X"E7",X"10",
		X"DC",X"C9",X"6F",X"CD",X"F1",X"18",X"CB",X"4D",X"3E",X"01",X"28",X"05",X"CD",X"F1",X"18",X"3E",
		X"02",X"32",X"76",X"43",X"2A",X"72",X"08",X"36",X"01",X"E1",X"C3",X"B8",X"17",X"E5",X"21",X"00",
		X"00",X"39",X"CD",X"E0",X"18",X"77",X"06",X"02",X"11",X"78",X"D5",X"CD",X"40",X"2A",X"E1",X"C9",
		X"3A",X"A5",X"08",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"4F",X"3A",X"A4",X"08",X"E6",X"F0",X"B1",
		X"C9",X"CD",X"E0",X"18",X"C6",X"99",X"27",X"4F",X"E6",X"F0",X"32",X"A4",X"08",X"79",X"07",X"07",
		X"07",X"07",X"E6",X"F0",X"32",X"A5",X"08",X"C9",X"7E",X"B7",X"C8",X"C5",X"E5",X"35",X"78",X"3D",
		X"87",X"87",X"87",X"5F",X"16",X"00",X"21",X"A6",X"08",X"19",X"06",X"08",X"CD",X"B3",X"2D",X"E1",
		X"E5",X"11",X"05",X"00",X"19",X"7E",X"57",X"3C",X"E6",X"03",X"77",X"ED",X"78",X"E6",X"0F",X"CB",
		X"1A",X"17",X"4F",X"06",X"00",X"21",X"5B",X"19",X"09",X"7E",X"CB",X"42",X"28",X"04",X"07",X"07",
		X"07",X"07",X"E6",X"0F",X"C6",X"00",X"27",X"57",X"CD",X"E0",X"18",X"FE",X"99",X"28",X"09",X"82",
		X"27",X"30",X"02",X"3E",X"99",X"CD",X"F7",X"18",X"E1",X"C1",X"C9",X"11",X"11",X"22",X"22",X"33",
		X"33",X"44",X"44",X"55",X"55",X"66",X"66",X"77",X"77",X"AA",X"AA",X"EE",X"EE",X"00",X"11",X"11",
		X"22",X"00",X"55",X"00",X"77",X"00",X"21",X"11",X"21",X"11",X"32",X"C5",X"21",X"9C",X"08",X"CD",
		X"E0",X"18",X"F5",X"01",X"62",X"03",X"CD",X"08",X"19",X"23",X"0C",X"10",X"F9",X"CD",X"E0",X"18",
		X"C1",X"B8",X"C4",X"CD",X"18",X"C1",X"C9",X"CD",X"E0",X"18",X"2E",X"00",X"B7",X"28",X"08",X"FE",
		X"01",X"2E",X"01",X"28",X"02",X"2E",X"03",X"DB",X"49",X"2F",X"A5",X"C9",X"CD",X"4E",X"1A",X"CD",
		X"AF",X"35",X"CD",X"7B",X"29",X"90",X"0C",X"BE",X"1F",X"31",X"39",X"38",X"30",X"20",X"53",X"54",
		X"45",X"52",X"4E",X"20",X"45",X"6C",X"65",X"63",X"74",X"72",X"6F",X"6E",X"69",X"63",X"73",X"2C",
		X"20",X"49",X"6E",X"63",X"2E",X"00",X"CD",X"CD",X"18",X"CD",X"14",X"23",X"CD",X"ED",X"1A",X"04",
		X"1B",X"2D",X"1B",X"17",X"1B",X"45",X"1B",X"21",X"02",X"43",X"3E",X"01",X"32",X"00",X"43",X"11",
		X"38",X"18",X"D5",X"E5",X"7E",X"23",X"B6",X"23",X"B6",X"E1",X"E5",X"20",X"04",X"E1",X"D1",X"18",
		X"35",X"21",X"00",X"43",X"06",X"02",X"CD",X"40",X"2A",X"13",X"E1",X"06",X"06",X"CD",X"4A",X"2A",
		X"13",X"AF",X"4E",X"CD",X"DB",X"29",X"13",X"23",X"4E",X"CD",X"DB",X"29",X"13",X"23",X"4E",X"CD",
		X"DB",X"29",X"23",X"D1",X"7A",X"C6",X"10",X"57",X"3A",X"00",X"43",X"C6",X"01",X"27",X"32",X"00",
		X"43",X"FE",X"11",X"C2",X"F2",X"19",X"21",X"00",X"46",X"CD",X"45",X"1A",X"21",X"00",X"5B",X"CD",
		X"45",X"1A",X"21",X"80",X"5D",X"3E",X"FF",X"06",X"40",X"77",X"23",X"10",X"FC",X"C9",X"21",X"00",
		X"81",X"01",X"00",X"07",X"AF",X"77",X"23",X"0D",X"20",X"FB",X"10",X"F9",X"F3",X"ED",X"73",X"00",
		X"43",X"31",X"00",X"60",X"06",X"E0",X"11",X"00",X"00",X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",
		X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",X"10",X"EE",X"ED",X"7B",X"00",X"43",X"FB",
		X"DB",X"4A",X"CB",X"7F",X"20",X"0D",X"3A",X"44",X"43",X"FE",X"02",X"20",X"06",X"3E",X"08",X"32",
		X"79",X"43",X"C9",X"AF",X"32",X"79",X"43",X"C9",X"CD",X"DD",X"1A",X"CD",X"E0",X"18",X"28",X"21",
		X"3D",X"28",X"0F",X"CD",X"13",X"36",X"CD",X"ED",X"1A",X"94",X"1B",X"DE",X"1B",X"BB",X"1B",X"FB",
		X"1B",X"C9",X"CD",X"0A",X"36",X"CD",X"ED",X"1A",X"54",X"1B",X"DE",X"1B",X"76",X"1B",X"FB",X"1B",
		X"C9",X"CD",X"01",X"36",X"CD",X"ED",X"1A",X"0F",X"1C",X"3F",X"1C",X"22",X"1C",X"56",X"1C",X"21",
		X"D6",X"1A",X"22",X"98",X"08",X"C9",X"65",X"10",X"09",X"0B",X"11",X"45",X"FF",X"21",X"C0",X"5B",
		X"01",X"C0",X"02",X"AF",X"77",X"23",X"0D",X"C2",X"E4",X"1A",X"10",X"F8",X"C9",X"E1",X"54",X"5D",
		X"01",X"08",X"00",X"09",X"E5",X"EB",X"DB",X"60",X"E6",X"C0",X"07",X"07",X"07",X"4F",X"09",X"7E",
		X"23",X"66",X"6F",X"E9",X"CD",X"7B",X"29",X"90",X"58",X"00",X"48",X"69",X"67",X"68",X"20",X"53",
		X"63",X"6F",X"72",X"65",X"73",X"00",X"C9",X"CD",X"7B",X"29",X"90",X"48",X"00",X"4D",X"65",X"69",
		X"6C",X"6C",X"65",X"75",X"72",X"20",X"53",X"63",X"6F",X"72",X"65",X"00",X"C9",X"CD",X"7B",X"29",
		X"90",X"40",X"00",X"48",X"6F",X"65",X"63",X"68",X"73",X"74",X"65",X"72",X"20",X"47",X"65",X"62",
		X"6E",X"69",X"73",X"00",X"C9",X"CD",X"7B",X"29",X"90",X"5C",X"00",X"52",X"65",X"63",X"6F",X"72",
		X"64",X"73",X"00",X"C9",X"CD",X"7B",X"29",X"90",X"14",X"BE",X"50",X"75",X"73",X"68",X"20",X"31",
		X"20",X"50",X"6C",X"61",X"79",X"65",X"72",X"20",X"53",X"74",X"61",X"72",X"74",X"20",X"42",X"75",
		X"74",X"74",X"6F",X"6E",X"00",X"C9",X"CD",X"7B",X"29",X"90",X"24",X"BE",X"50",X"6F",X"75",X"73",
		X"73",X"65",X"72",X"20",X"62",X"6F",X"75",X"74",X"6F",X"6E",X"20",X"73",X"74",X"61",X"72",X"74",
		X"20",X"31",X"00",X"C9",X"CD",X"7B",X"29",X"90",X"04",X"BE",X"50",X"75",X"73",X"68",X"20",X"31",
		X"20",X"6F",X"72",X"20",X"32",X"20",X"50",X"6C",X"61",X"79",X"65",X"72",X"20",X"53",X"74",X"61",
		X"72",X"74",X"20",X"42",X"75",X"74",X"74",X"6F",X"6E",X"00",X"C9",X"CD",X"7B",X"29",X"90",X"10",
		X"BE",X"50",X"6F",X"75",X"73",X"73",X"65",X"72",X"20",X"62",X"6F",X"75",X"74",X"6F",X"6E",X"20",
		X"73",X"74",X"61",X"72",X"74",X"20",X"31",X"20",X"6F",X"75",X"20",X"32",X"00",X"C9",X"CD",X"7B",
		X"29",X"90",X"20",X"BE",X"53",X"74",X"61",X"72",X"74",X"6B",X"6E",X"6F",X"65",X"70",X"66",X"65",
		X"20",X"64",X"72",X"75",X"65",X"63",X"6B",X"65",X"6E",X"00",X"C9",X"CD",X"7B",X"29",X"90",X"44",
		X"BE",X"50",X"75",X"6C",X"73",X"61",X"72",X"20",X"53",X"74",X"61",X"72",X"74",X"00",X"C9",X"CD",
		X"7B",X"29",X"90",X"58",X"BE",X"49",X"6E",X"73",X"65",X"72",X"74",X"20",X"43",X"6F",X"69",X"6E",
		X"00",X"C9",X"CD",X"7B",X"29",X"90",X"30",X"BE",X"49",X"6E",X"74",X"72",X"6F",X"64",X"75",X"69",
		X"72",X"65",X"20",X"6C",X"61",X"20",X"6D",X"6F",X"6E",X"6E",X"61",X"69",X"65",X"00",X"C9",X"CD",
		X"7B",X"29",X"90",X"48",X"BE",X"4D",X"75",X"6E",X"7A",X"65",X"20",X"65",X"69",X"6E",X"77",X"65",
		X"72",X"66",X"65",X"6E",X"00",X"C9",X"CD",X"7B",X"29",X"90",X"48",X"BE",X"50",X"6F",X"6E",X"67",
		X"61",X"20",X"6C",X"61",X"20",X"6D",X"6F",X"6E",X"65",X"64",X"61",X"00",X"C9",X"A3",X"C5",X"F5",
		X"FD",X"2A",X"76",X"08",X"FD",X"66",X"07",X"FD",X"6E",X"09",X"CD",X"E7",X"1C",X"D5",X"DD",X"66",
		X"07",X"DD",X"6E",X"09",X"2D",X"2D",X"2D",X"2D",X"25",X"25",X"25",X"25",X"CD",X"E7",X"1C",X"D9",
		X"47",X"D9",X"C1",X"79",X"BB",X"20",X"03",X"F1",X"C1",X"C9",X"7C",X"E5",X"C6",X"10",X"67",X"CD",
		X"E7",X"1C",X"D9",X"4F",X"D9",X"7D",X"C6",X"13",X"6F",X"CD",X"E7",X"1C",X"D9",X"57",X"D9",X"7D",
		X"E1",X"6F",X"CD",X"E7",X"1C",X"D9",X"5F",X"F1",X"67",X"2E",X"00",X"CB",X"5C",X"28",X"06",X"78",
		X"B1",X"E6",X"08",X"B5",X"6F",X"CB",X"54",X"28",X"06",X"7A",X"B3",X"E6",X"04",X"B5",X"6F",X"CB",
		X"4C",X"28",X"06",X"78",X"B3",X"E6",X"02",X"B5",X"6F",X"CB",X"44",X"28",X"06",X"79",X"B2",X"E6",
		X"01",X"B5",X"6F",X"2F",X"A4",X"C1",X"C9",X"7D",X"1E",X"00",X"FE",X"46",X"38",X"08",X"1E",X"05",
		X"FE",X"8A",X"38",X"02",X"1E",X"0A",X"7C",X"06",X"05",X"0E",X"3A",X"16",X"30",X"B9",X"38",X"08",
		X"1C",X"08",X"79",X"82",X"4F",X"08",X"10",X"F5",X"EB",X"01",X"5E",X"43",X"26",X"00",X"09",X"7E",
		X"EB",X"C9",X"DD",X"21",X"22",X"1D",X"ED",X"4B",X"85",X"08",X"CD",X"22",X"1D",X"ED",X"43",X"85",
		X"08",X"C9",X"0A",X"03",X"26",X"00",X"87",X"6F",X"11",X"31",X"1D",X"19",X"7E",X"23",X"66",X"6F",
		X"E9",X"51",X"1D",X"5C",X"1D",X"5D",X"1D",X"68",X"1D",X"74",X"1D",X"7E",X"1D",X"8A",X"1D",X"96",
		X"1D",X"A7",X"1D",X"B1",X"1D",X"BD",X"1D",X"CB",X"1D",X"E4",X"1D",X"F4",X"1D",X"09",X"1E",X"1C",
		X"1E",X"0B",X"21",X"00",X"00",X"22",X"87",X"08",X"22",X"89",X"08",X"C9",X"C9",X"0A",X"03",X"6F",
		X"87",X"9F",X"67",X"09",X"44",X"4D",X"DD",X"E9",X"0A",X"03",X"6F",X"0A",X"03",X"67",X"35",X"20",
		X"EC",X"03",X"DD",X"E9",X"0A",X"03",X"6F",X"0A",X"03",X"67",X"5E",X"C3",X"8D",X"1D",X"0A",X"03",
		X"6F",X"0A",X"03",X"67",X"5E",X"23",X"56",X"C3",X"9C",X"1D",X"0A",X"03",X"5F",X"0A",X"03",X"6F",
		X"0A",X"03",X"67",X"73",X"DD",X"E9",X"0A",X"03",X"5F",X"0A",X"03",X"57",X"0A",X"03",X"6F",X"0A",
		X"03",X"67",X"73",X"23",X"72",X"DD",X"E9",X"0A",X"03",X"6F",X"0A",X"03",X"67",X"5E",X"C3",X"C0",
		X"1D",X"0A",X"03",X"6F",X"0A",X"03",X"67",X"5E",X"23",X"56",X"C3",X"D1",X"1D",X"0A",X"03",X"5F",
		X"0A",X"03",X"6F",X"0A",X"03",X"67",X"7E",X"83",X"77",X"DD",X"E9",X"0A",X"03",X"5F",X"0A",X"03",
		X"57",X"0A",X"03",X"6F",X"0A",X"03",X"67",X"E5",X"7E",X"23",X"66",X"6F",X"19",X"EB",X"E1",X"73",
		X"23",X"72",X"DD",X"E9",X"0A",X"03",X"5F",X"0A",X"03",X"6F",X"0A",X"03",X"67",X"CB",X"2E",X"1D",
		X"20",X"FB",X"DD",X"E9",X"0A",X"03",X"5F",X"0A",X"03",X"6F",X"0A",X"03",X"67",X"23",X"CB",X"2E",
		X"2B",X"CB",X"1E",X"23",X"1D",X"20",X"F7",X"DD",X"E9",X"0A",X"03",X"5F",X"0A",X"03",X"6F",X"0A",
		X"03",X"67",X"0A",X"77",X"23",X"03",X"1D",X"C2",X"12",X"1E",X"DD",X"E9",X"0A",X"03",X"87",X"C3",
		X"0B",X"1E",X"E1",X"D9",X"21",X"01",X"00",X"E5",X"E5",X"21",X"00",X"00",X"39",X"3A",X"73",X"08",
		X"B7",X"20",X"06",X"E5",X"22",X"72",X"08",X"18",X"1E",X"FD",X"E5",X"C1",X"FD",X"2A",X"72",X"08",
		X"EB",X"FD",X"66",X"FF",X"FD",X"6E",X"FE",X"E5",X"F3",X"FD",X"72",X"FF",X"FD",X"73",X"FE",X"FB",
		X"ED",X"53",X"72",X"08",X"C5",X"FD",X"E1",X"D9",X"E9",X"21",X"00",X"00",X"39",X"EB",X"21",X"E8",
		X"FF",X"39",X"F9",X"2A",X"72",X"08",X"23",X"23",X"73",X"23",X"72",X"FD",X"E9",X"FD",X"2A",X"72",
		X"08",X"FD",X"77",X"01",X"FD",X"36",X"00",X"82",X"FD",X"2A",X"72",X"08",X"21",X"00",X"00",X"39",
		X"31",X"70",X"08",X"FD",X"75",X"02",X"FD",X"74",X"03",X"18",X"04",X"FD",X"2A",X"72",X"08",X"FD",
		X"66",X"FF",X"FD",X"6E",X"FE",X"E5",X"FD",X"E1",X"CB",X"46",X"CA",X"8F",X"1E",X"FD",X"6E",X"02",
		X"FD",X"66",X"03",X"FD",X"22",X"72",X"08",X"F9",X"C9",X"CD",X"D4",X"1F",X"DD",X"36",X"00",X"16",
		X"CD",X"22",X"1E",X"C5",X"FD",X"21",X"8B",X"1E",X"CD",X"59",X"1E",X"C1",X"DD",X"2A",X"76",X"08",
		X"DD",X"CB",X"00",X"7E",X"C2",X"A7",X"1F",X"3A",X"6E",X"43",X"B7",X"28",X"14",X"2A",X"6F",X"43",
		X"7E",X"23",X"22",X"6F",X"43",X"CB",X"7F",X"28",X"16",X"CB",X"BF",X"C5",X"CD",X"6D",X"1E",X"18",
		X"DA",X"3A",X"79",X"43",X"B7",X"28",X"04",X"DB",X"4A",X"18",X"02",X"DB",X"48",X"EE",X"1F",X"CB",
		X"67",X"57",X"20",X"0D",X"E6",X"0F",X"B9",X"C4",X"91",X"1F",X"C5",X"CD",X"78",X"1E",X"C3",X"BB",
		X"1E",X"FD",X"CB",X"00",X"4E",X"20",X"F3",X"AF",X"FD",X"21",X"7B",X"43",X"FD",X"B6",X"04",X"28",
		X"0A",X"FD",X"21",X"83",X"43",X"AF",X"FD",X"B6",X"04",X"20",X"DF",X"7A",X"E6",X"0F",X"CA",X"FA",
		X"1E",X"CD",X"BD",X"33",X"4F",X"21",X"42",X"20",X"06",X"00",X"50",X"09",X"5E",X"21",X"67",X"20",
		X"19",X"19",X"19",X"DD",X"36",X"06",X"00",X"DD",X"36",X"08",X"00",X"7E",X"23",X"F3",X"DD",X"77",
		X"0A",X"7E",X"23",X"DD",X"77",X"0B",X"FB",X"DD",X"36",X"0C",X"01",X"00",X"DD",X"7E",X"0C",X"FE",
		X"02",X"20",X"F8",X"0E",X"FF",X"C5",X"46",X"23",X"4E",X"23",X"56",X"DD",X"7E",X"07",X"80",X"6F",
		X"DD",X"7E",X"09",X"81",X"67",X"FD",X"75",X"02",X"FD",X"74",X"03",X"FD",X"75",X"06",X"FD",X"74",
		X"07",X"F3",X"FD",X"72",X"00",X"FD",X"36",X"01",X"00",X"FD",X"72",X"04",X"FD",X"36",X"05",X"08",
		X"FB",X"3E",X"08",X"CD",X"6D",X"1E",X"FD",X"CB",X"00",X"CE",X"FD",X"36",X"01",X"0C",X"C3",X"BB",
		X"1E",X"4F",X"E6",X"0F",X"CD",X"3D",X"2B",X"21",X"53",X"20",X"19",X"7E",X"23",X"66",X"F3",X"DD",
		X"77",X"0A",X"DD",X"74",X"0B",X"FB",X"C9",X"CD",X"39",X"34",X"3E",X"10",X"CD",X"94",X"1F",X"DD",
		X"CB",X"00",X"EE",X"CD",X"1F",X"2C",X"3E",X"2D",X"CD",X"6D",X"1E",X"FD",X"7E",X"01",X"B7",X"28",
		X"05",X"CD",X"78",X"1E",X"18",X"F5",X"2A",X"76",X"08",X"36",X"09",X"FD",X"CB",X"00",X"86",X"CD",
		X"78",X"1E",X"18",X"FB",X"FD",X"E1",X"21",X"00",X"00",X"06",X"07",X"E5",X"10",X"FD",X"DD",X"21",
		X"00",X"00",X"DD",X"39",X"E5",X"DD",X"22",X"76",X"08",X"3A",X"44",X"43",X"FE",X"01",X"3E",X"AA",
		X"28",X"02",X"3E",X"DD",X"32",X"78",X"43",X"2A",X"47",X"43",X"DD",X"75",X"07",X"DD",X"74",X"09",
		X"AF",X"CD",X"91",X"1F",X"DD",X"36",X"0D",X"02",X"DD",X"36",X"0C",X"01",X"FD",X"E9",X"E1",X"D9",
		X"06",X"07",X"11",X"00",X"00",X"D5",X"10",X"FD",X"21",X"00",X"00",X"39",X"EB",X"3A",X"71",X"08",
		X"B7",X"20",X"07",X"D5",X"ED",X"53",X"70",X"08",X"18",X"13",X"DD",X"2A",X"70",X"08",X"DD",X"66",
		X"FF",X"DD",X"6E",X"FE",X"E5",X"F3",X"DD",X"72",X"FF",X"DD",X"73",X"FE",X"FB",X"D5",X"DD",X"E1",
		X"D9",X"E9",X"00",X"0C",X"04",X"00",X"10",X"0E",X"02",X"10",X"08",X"0A",X"06",X"08",X"00",X"0C",
		X"04",X"00",X"12",X"46",X"10",X"4B",X"10",X"4B",X"10",X"4B",X"10",X"4B",X"10",X"56",X"10",X"56",
		X"10",X"56",X"10",X"4B",X"10",X"B3",X"12",X"46",X"10",X"00",X"00",X"00",X"00",X"61",X"10",X"07",
		X"01",X"06",X"00",X"66",X"10",X"07",X"03",X"02",X"00",X"6B",X"10",X"06",X"06",X"0A",X"00",X"70",
		X"10",X"06",X"07",X"08",X"00",X"75",X"10",X"00",X"06",X"09",X"00",X"7A",X"10",X"00",X"03",X"01",
		X"00",X"7F",X"10",X"00",X"00",X"05",X"00",X"84",X"10",X"07",X"02",X"04",X"00",X"CD",X"4E",X"1A",
		X"CD",X"40",X"25",X"3A",X"6E",X"43",X"B7",X"20",X"2E",X"CD",X"D4",X"1F",X"01",X"12",X"18",X"3A",
		X"76",X"43",X"FE",X"02",X"28",X"02",X"06",X"08",X"DD",X"71",X"00",X"C5",X"DD",X"E5",X"3E",X"0A",
		X"CD",X"6D",X"1E",X"DD",X"E1",X"C1",X"3E",X"1B",X"A9",X"4F",X"10",X"EC",X"21",X"00",X"00",X"22",
		X"76",X"08",X"06",X"08",X"D1",X"10",X"FD",X"FB",X"3A",X"4A",X"43",X"C6",X"60",X"27",X"32",X"4A",
		X"43",X"3A",X"4C",X"43",X"FE",X"01",X"28",X"04",X"3D",X"32",X"4C",X"43",X"AF",X"32",X"71",X"43",
		X"FD",X"2A",X"72",X"08",X"FD",X"77",X"01",X"3A",X"4D",X"43",X"FE",X"14",X"38",X"05",X"D6",X"0A",
		X"32",X"4D",X"43",X"FD",X"21",X"17",X"21",X"21",X"F0",X"FF",X"39",X"F9",X"CD",X"59",X"1E",X"21",
		X"10",X"00",X"39",X"F9",X"C3",X"57",X"21",X"3E",X"16",X"32",X"00",X"43",X"4F",X"3A",X"4A",X"43",
		X"47",X"CD",X"78",X"26",X"B8",X"38",X"1E",X"21",X"A0",X"23",X"06",X"00",X"09",X"46",X"23",X"4E",
		X"CD",X"78",X"26",X"E6",X"1F",X"80",X"47",X"CD",X"78",X"26",X"E6",X"1F",X"81",X"4F",X"FD",X"21",
		X"45",X"21",X"C3",X"B8",X"23",X"3A",X"00",X"43",X"3D",X"3D",X"32",X"00",X"43",X"4F",X"20",X"CD",
		X"FD",X"21",X"A9",X"1E",X"C3",X"8E",X"2A",X"DD",X"2A",X"76",X"08",X"DD",X"CB",X"00",X"56",X"C8",
		X"DD",X"7E",X"09",X"32",X"48",X"43",X"47",X"DD",X"7E",X"07",X"32",X"47",X"43",X"DD",X"CB",X"00",
		X"7E",X"C2",X"8D",X"21",X"B7",X"F2",X"82",X"21",X"FE",X"FC",X"D2",X"AC",X"22",X"FE",X"F6",X"D2",
		X"5D",X"22",X"78",X"FE",X"02",X"DA",X"20",X"22",X"FE",X"BE",X"D2",X"CF",X"21",X"3A",X"6D",X"43",
		X"B7",X"28",X"03",X"CD",X"14",X"23",X"3A",X"6E",X"43",X"B7",X"28",X"07",X"CD",X"7B",X"19",X"CD",
		X"97",X"19",X"C0",X"FD",X"2A",X"72",X"08",X"FD",X"CB",X"00",X"CE",X"FD",X"7E",X"01",X"B7",X"20",
		X"18",X"FD",X"36",X"01",X"3B",X"06",X"0C",X"21",X"D0",X"08",X"3A",X"6E",X"43",X"B7",X"20",X"06",
		X"CD",X"B3",X"2D",X"CD",X"97",X"2B",X"CD",X"78",X"26",X"CD",X"78",X"1E",X"C3",X"57",X"21",X"3E",
		X"06",X"32",X"48",X"43",X"21",X"46",X"43",X"34",X"CD",X"EB",X"22",X"28",X"09",X"21",X"AD",X"5F",
		X"11",X"DF",X"5F",X"C3",X"3D",X"22",X"21",X"2D",X"44",X"11",X"00",X"44",X"E5",X"3E",X"1B",X"21",
		X"00",X"01",X"19",X"01",X"00",X"19",X"D5",X"ED",X"B0",X"D1",X"01",X"00",X"01",X"2B",X"36",X"00",
		X"0D",X"C2",X"FD",X"21",X"10",X"F7",X"3D",X"20",X"E6",X"CD",X"40",X"25",X"E1",X"11",X"1A",X"00",
		X"0E",X"02",X"06",X"06",X"36",X"FF",X"23",X"10",X"FB",X"19",X"0D",X"20",X"F5",X"C3",X"D7",X"20",
		X"3E",X"B9",X"32",X"48",X"43",X"21",X"46",X"43",X"35",X"CD",X"EB",X"22",X"28",X"09",X"21",X"2D",
		X"46",X"11",X"00",X"46",X"C3",X"EC",X"21",X"21",X"AD",X"5D",X"11",X"FF",X"5D",X"E5",X"3E",X"1A",
		X"01",X"00",X"19",X"21",X"00",X"FF",X"19",X"D5",X"ED",X"B8",X"D1",X"01",X"00",X"01",X"23",X"36",
		X"00",X"0D",X"C2",X"4E",X"22",X"10",X"F7",X"3D",X"20",X"E6",X"C3",X"09",X"22",X"3E",X"08",X"32",
		X"47",X"43",X"21",X"45",X"43",X"34",X"CD",X"EB",X"22",X"28",X"09",X"21",X"1F",X"4F",X"11",X"E0",
		X"5F",X"C3",X"C9",X"22",X"21",X"00",X"4D",X"11",X"00",X"44",X"E5",X"3E",X"20",X"01",X"FF",X"19",
		X"21",X"01",X"00",X"19",X"D5",X"ED",X"B0",X"06",X"D0",X"11",X"E1",X"FF",X"36",X"00",X"2B",X"36",
		X"00",X"19",X"10",X"F8",X"D1",X"3D",X"20",X"E5",X"3E",X"06",X"F5",X"CD",X"40",X"25",X"F1",X"E1",
		X"11",X"20",X"00",X"06",X"40",X"77",X"19",X"10",X"FC",X"C3",X"D7",X"20",X"3E",X"E6",X"32",X"47",
		X"43",X"21",X"45",X"43",X"35",X"CD",X"EB",X"22",X"28",X"09",X"21",X"00",X"4F",X"11",X"00",X"46",
		X"C3",X"7A",X"22",X"21",X"1F",X"4D",X"11",X"00",X"5E",X"E5",X"3E",X"20",X"01",X"00",X"1A",X"21",
		X"FF",X"FF",X"19",X"D5",X"ED",X"B8",X"11",X"1F",X"00",X"36",X"00",X"23",X"36",X"00",X"19",X"10",
		X"F8",X"D1",X"3D",X"20",X"E7",X"3E",X"60",X"F5",X"C3",X"9B",X"22",X"CD",X"E4",X"2B",X"CD",X"4E",
		X"36",X"FD",X"E5",X"E1",X"FD",X"74",X"FF",X"FD",X"75",X"FE",X"21",X"00",X"00",X"F3",X"22",X"70",
		X"08",X"22",X"76",X"08",X"AF",X"21",X"7B",X"43",X"06",X"38",X"77",X"23",X"10",X"FC",X"3A",X"79",
		X"43",X"B7",X"FB",X"C9",X"AF",X"32",X"6D",X"43",X"11",X"00",X"D5",X"21",X"3E",X"43",X"06",X"06",
		X"CD",X"40",X"2A",X"3A",X"76",X"43",X"FE",X"02",X"C0",X"11",X"B0",X"D5",X"21",X"41",X"43",X"06",
		X"06",X"C3",X"40",X"2A",X"3A",X"44",X"43",X"FE",X"02",X"21",X"41",X"43",X"C8",X"21",X"3E",X"43",
		X"C9",X"3E",X"FF",X"32",X"6D",X"43",X"1E",X"04",X"CD",X"34",X"23",X"23",X"23",X"23",X"CB",X"38",
		X"08",X"04",X"2B",X"1D",X"10",X"FC",X"08",X"30",X"08",X"CB",X"21",X"CB",X"21",X"CB",X"21",X"CB",
		X"21",X"79",X"86",X"27",X"77",X"30",X"08",X"2B",X"1D",X"28",X"04",X"0E",X"01",X"18",X"F2",X"CD",
		X"34",X"23",X"44",X"4D",X"21",X"4F",X"43",X"11",X"49",X"43",X"DB",X"61",X"CB",X"7F",X"28",X"11",
		X"0A",X"B7",X"28",X"0D",X"CB",X"4E",X"C0",X"CB",X"CE",X"EB",X"34",X"CD",X"38",X"35",X"C3",X"9A",
		X"25",X"DB",X"61",X"CB",X"77",X"C8",X"03",X"0A",X"FE",X"50",X"D8",X"CB",X"46",X"C0",X"CB",X"C6",
		X"18",X"E7",X"0C",X"0C",X"40",X"0C",X"A0",X"0C",X"CE",X"0C",X"40",X"50",X"70",X"50",X"9E",X"50",
		X"0C",X"96",X"40",X"96",X"A0",X"96",X"CE",X"96",X"C5",X"D1",X"21",X"71",X"43",X"34",X"7E",X"32",
		X"72",X"43",X"CD",X"0E",X"20",X"DD",X"72",X"07",X"DD",X"73",X"09",X"AF",X"CD",X"36",X"24",X"DD",
		X"36",X"0C",X"01",X"DD",X"36",X"00",X"06",X"CD",X"22",X"1E",X"DD",X"E5",X"CD",X"59",X"1E",X"3A",
		X"4D",X"43",X"FE",X"1E",X"30",X"02",X"3E",X"1E",X"CD",X"6D",X"1E",X"DD",X"E1",X"0E",X"00",X"FD",
		X"2A",X"76",X"08",X"C5",X"FD",X"7E",X"07",X"DD",X"96",X"07",X"57",X"06",X"00",X"28",X"06",X"06",
		X"01",X"38",X"02",X"06",X"02",X"FD",X"7E",X"09",X"C6",X"02",X"DD",X"96",X"09",X"5F",X"0E",X"00",
		X"28",X"06",X"0E",X"04",X"38",X"02",X"0E",X"08",X"78",X"81",X"F5",X"4F",X"CD",X"7F",X"28",X"F1",
		X"C1",X"CD",X"36",X"24",X"DD",X"E5",X"C5",X"CD",X"78",X"1E",X"C1",X"DD",X"E1",X"DD",X"CB",X"00",
		X"7E",X"CA",X"EF",X"23",X"18",X"21",X"E6",X"0F",X"C4",X"6E",X"1C",X"B9",X"C8",X"4F",X"CD",X"3D",
		X"2B",X"21",X"2D",X"25",X"19",X"7E",X"23",X"66",X"F3",X"DD",X"77",X"0A",X"DD",X"74",X"0B",X"FB",
		X"3A",X"4C",X"43",X"DD",X"77",X"0D",X"C9",X"E5",X"DD",X"E5",X"CD",X"8A",X"34",X"E1",X"11",X"06",
		X"00",X"19",X"F3",X"72",X"23",X"7E",X"D6",X"04",X"77",X"23",X"72",X"23",X"7E",X"D6",X"06",X"77",
		X"23",X"01",X"3B",X"10",X"71",X"23",X"70",X"FB",X"23",X"36",X"01",X"23",X"36",X"01",X"DD",X"E5",
		X"01",X"05",X"01",X"CD",X"41",X"23",X"21",X"4E",X"43",X"34",X"34",X"21",X"71",X"43",X"35",X"20",
		X"3A",X"3A",X"72",X"43",X"F5",X"01",X"01",X"01",X"CD",X"41",X"23",X"F1",X"3D",X"20",X"F5",X"CD",
		X"7B",X"29",X"00",X"60",X"D5",X"42",X"4F",X"4E",X"55",X"53",X"00",X"F5",X"3A",X"72",X"43",X"C6",
		X"00",X"27",X"0F",X"0F",X"0F",X"0F",X"6F",X"E6",X"F0",X"67",X"3E",X"0F",X"A5",X"6F",X"F1",X"22",
		X"00",X"43",X"08",X"21",X"00",X"43",X"06",X"04",X"CD",X"4A",X"2A",X"3E",X"1E",X"CD",X"6D",X"1E",
		X"DD",X"E1",X"21",X"08",X"12",X"DD",X"7E",X"04",X"BD",X"20",X"06",X"DD",X"7E",X"05",X"BC",X"28",
		X"09",X"DD",X"E5",X"CD",X"78",X"1E",X"DD",X"E1",X"18",X"E8",X"CD",X"F7",X"24",X"2A",X"72",X"08",
		X"CB",X"86",X"CD",X"78",X"1E",X"18",X"F6",X"DD",X"E5",X"C1",X"50",X"59",X"EB",X"2B",X"56",X"2B",
		X"5E",X"78",X"BA",X"20",X"F7",X"79",X"BB",X"20",X"F3",X"F3",X"DD",X"7E",X"FE",X"77",X"23",X"DD",
		X"7E",X"FF",X"77",X"23",X"22",X"70",X"08",X"FB",X"C9",X"00",X"00",X"01",X"FF",X"01",X"00",X"01",
		X"01",X"00",X"01",X"FF",X"01",X"FF",X"00",X"FF",X"FF",X"00",X"FF",X"00",X"00",X"00",X"10",X"13",
		X"10",X"13",X"10",X"13",X"10",X"1C",X"10",X"27",X"10",X"27",X"10",X"27",X"10",X"30",X"10",X"41",
		X"2A",X"45",X"43",X"22",X"5C",X"43",X"3A",X"79",X"43",X"B7",X"20",X"05",X"21",X"6A",X"5E",X"18",
		X"03",X"21",X"4A",X"44",X"11",X"14",X"00",X"AF",X"0E",X"0C",X"06",X"0C",X"77",X"23",X"10",X"FC",
		X"19",X"0D",X"20",X"F6",X"01",X"0F",X"00",X"11",X"5E",X"43",X"21",X"8C",X"26",X"ED",X"B0",X"21",
		X"08",X"00",X"CD",X"D4",X"25",X"21",X"08",X"CC",X"CD",X"D4",X"25",X"21",X"04",X"00",X"CD",X"CA",
		X"25",X"21",X"F8",X"00",X"CD",X"CA",X"25",X"DD",X"21",X"5E",X"43",X"21",X"38",X"44",X"CD",X"EB",
		X"25",X"21",X"38",X"88",X"CD",X"EB",X"25",X"CD",X"9F",X"36",X"3A",X"44",X"43",X"FE",X"02",X"21",
		X"38",X"D5",X"20",X"02",X"2E",X"E8",X"06",X"00",X"CD",X"A3",X"29",X"EB",X"08",X"3A",X"49",X"43",
		X"47",X"08",X"05",X"28",X"0A",X"C5",X"0E",X"80",X"CD",X"DB",X"29",X"13",X"C1",X"10",X"F6",X"3A",
		X"6E",X"43",X"B7",X"C4",X"CD",X"18",X"CD",X"14",X"23",X"C9",X"CD",X"62",X"26",X"3E",X"40",X"84",
		X"67",X"C3",X"62",X"26",X"CD",X"4C",X"26",X"CD",X"4C",X"26",X"3E",X"30",X"85",X"6F",X"CD",X"4C",
		X"26",X"C3",X"4C",X"26",X"06",X"10",X"CD",X"A3",X"29",X"EB",X"C9",X"CD",X"78",X"26",X"E5",X"CD",
		X"78",X"26",X"01",X"06",X"26",X"C5",X"E6",X"03",X"CA",X"30",X"26",X"3D",X"CA",X"40",X"26",X"3D",
		X"CA",X"14",X"26",X"C3",X"20",X"26",X"E1",X"DD",X"23",X"3E",X"30",X"85",X"6F",X"FE",X"DC",X"38",
		X"DA",X"DD",X"23",X"C9",X"CD",X"4C",X"26",X"DD",X"CB",X"01",X"DE",X"DD",X"CB",X"06",X"D6",X"C9",
		X"7D",X"D6",X"30",X"6F",X"CD",X"4C",X"26",X"DD",X"CB",X"00",X"DE",X"DD",X"CB",X"05",X"D6",X"C9",
		X"7C",X"D6",X"44",X"67",X"CD",X"62",X"26",X"DD",X"CB",X"00",X"CE",X"DD",X"CB",X"01",X"C6",X"C9",
		X"CD",X"62",X"26",X"DD",X"CB",X"05",X"CE",X"DD",X"CB",X"06",X"C6",X"C9",X"06",X"0C",X"C5",X"E5",
		X"CD",X"E4",X"25",X"21",X"9B",X"26",X"CD",X"17",X"28",X"E1",X"C1",X"3E",X"04",X"85",X"6F",X"10",
		X"ED",X"C9",X"06",X"12",X"C5",X"E5",X"CD",X"E4",X"25",X"21",X"9B",X"26",X"CD",X"17",X"28",X"E1",
		X"C1",X"3E",X"04",X"84",X"67",X"10",X"ED",X"C9",X"E5",X"2A",X"5C",X"43",X"54",X"5D",X"29",X"19",
		X"29",X"19",X"11",X"53",X"31",X"19",X"22",X"5C",X"43",X"7C",X"E1",X"C9",X"05",X"04",X"04",X"04",
		X"06",X"01",X"00",X"00",X"00",X"02",X"09",X"08",X"08",X"08",X"0A",X"01",X"04",X"F0",X"F0",X"F0",
		X"F0",X"02",X"04",X"FF",X"F0",X"FF",X"F0",X"FF",X"F0",X"FF",X"F0",X"F3",X"ED",X"73",X"74",X"08",
		X"31",X"40",X"08",X"F5",X"DB",X"4E",X"1F",X"38",X"20",X"E5",X"C5",X"21",X"9F",X"08",X"7E",X"23",
		X"46",X"A8",X"4F",X"DB",X"49",X"2F",X"77",X"2B",X"70",X"A1",X"E6",X"E0",X"2B",X"87",X"30",X"03",
		X"34",X"18",X"F9",X"20",X"F7",X"C1",X"E1",X"18",X"43",X"FD",X"E5",X"DD",X"E5",X"E5",X"D5",X"C5",
		X"08",X"F5",X"2A",X"70",X"08",X"E5",X"2A",X"76",X"08",X"CD",X"2D",X"27",X"CD",X"19",X"37",X"E1",
		X"E5",X"CD",X"2D",X"27",X"CD",X"F3",X"14",X"2A",X"76",X"08",X"CD",X"A9",X"27",X"E1",X"CD",X"A9",
		X"27",X"2A",X"70",X"08",X"7C",X"B5",X"28",X"08",X"2B",X"56",X"2B",X"5E",X"ED",X"53",X"70",X"08",
		X"CD",X"F5",X"27",X"F1",X"08",X"C1",X"D1",X"E1",X"DD",X"E1",X"FD",X"E1",X"3E",X"01",X"D3",X"4F",
		X"3E",X"37",X"ED",X"47",X"ED",X"5E",X"F1",X"ED",X"7B",X"74",X"08",X"FB",X"C9",X"22",X"70",X"08",
		X"E5",X"FD",X"E1",X"CB",X"46",X"CA",X"4D",X"27",X"CB",X"86",X"23",X"7E",X"D3",X"4B",X"23",X"5E",
		X"23",X"56",X"23",X"7E",X"23",X"66",X"6F",X"CD",X"17",X"28",X"2A",X"70",X"08",X"CB",X"4E",X"C8",
		X"CB",X"8E",X"11",X"07",X"00",X"19",X"5E",X"23",X"23",X"56",X"23",X"06",X"90",X"EB",X"CD",X"A3",
		X"29",X"FD",X"77",X"01",X"EB",X"7E",X"23",X"66",X"6F",X"7E",X"23",X"6E",X"67",X"7E",X"CB",X"7F",
		X"28",X"19",X"23",X"E6",X"7F",X"47",X"7E",X"23",X"4F",X"EB",X"3A",X"79",X"43",X"B7",X"CA",X"86",
		X"27",X"ED",X"42",X"C3",X"8A",X"27",X"09",X"C3",X"8A",X"27",X"EB",X"FD",X"75",X"04",X"FD",X"74",
		X"05",X"FD",X"73",X"02",X"FD",X"72",X"03",X"CD",X"17",X"28",X"2A",X"70",X"08",X"DB",X"4E",X"CB",
		X"7F",X"C8",X"CB",X"FE",X"FD",X"CB",X"FA",X"C6",X"C9",X"22",X"70",X"08",X"CB",X"56",X"C8",X"E5",
		X"FD",X"E1",X"11",X"0C",X"00",X"19",X"35",X"C0",X"23",X"7E",X"2B",X"77",X"11",X"FA",X"FF",X"19",
		X"7E",X"23",X"86",X"77",X"23",X"7E",X"23",X"86",X"77",X"23",X"5E",X"23",X"56",X"13",X"13",X"EB",
		X"7E",X"B7",X"C2",X"DA",X"27",X"23",X"7E",X"23",X"66",X"6F",X"EB",X"72",X"2B",X"73",X"3E",X"1B",
		X"FD",X"B6",X"00",X"FD",X"77",X"00",X"FD",X"CB",X"00",X"6E",X"C8",X"3A",X"78",X"43",X"07",X"EE",
		X"11",X"32",X"78",X"43",X"C9",X"2A",X"72",X"08",X"7C",X"B5",X"C8",X"54",X"5D",X"CB",X"4E",X"28",
		X"09",X"23",X"35",X"2B",X"20",X"04",X"CB",X"8E",X"CB",X"C6",X"2B",X"7E",X"2B",X"6E",X"67",X"BA",
		X"20",X"EB",X"7D",X"BB",X"20",X"E7",X"C9",X"06",X"00",X"7E",X"23",X"3D",X"CA",X"53",X"28",X"3A",
		X"79",X"43",X"B7",X"7E",X"23",X"C2",X"3D",X"28",X"01",X"1E",X"00",X"EB",X"08",X"1A",X"13",X"77",
		X"23",X"1A",X"13",X"77",X"23",X"70",X"08",X"09",X"3D",X"C2",X"2C",X"28",X"C9",X"01",X"E2",X"FF",
		X"EB",X"08",X"1A",X"13",X"77",X"2B",X"1A",X"13",X"77",X"2B",X"36",X"00",X"08",X"09",X"3D",X"C2",
		X"41",X"28",X"C9",X"3A",X"79",X"43",X"B7",X"7E",X"23",X"C2",X"6D",X"28",X"01",X"1F",X"00",X"EB",
		X"08",X"1A",X"13",X"77",X"23",X"70",X"08",X"09",X"3D",X"C2",X"60",X"28",X"C9",X"01",X"E1",X"FF",
		X"EB",X"08",X"1A",X"13",X"77",X"2B",X"36",X"00",X"08",X"09",X"3D",X"C2",X"71",X"28",X"C9",X"2A",
		X"72",X"08",X"23",X"7E",X"B7",X"C0",X"C5",X"D5",X"11",X"08",X"00",X"21",X"8F",X"43",X"3A",X"4B",
		X"43",X"B7",X"28",X"08",X"47",X"7E",X"B7",X"28",X"06",X"19",X"10",X"F9",X"D1",X"C1",X"C9",X"D1",
		X"C1",X"2B",X"2B",X"2B",X"2B",X"7A",X"FE",X"FE",X"D2",X"D8",X"28",X"FE",X"06",X"38",X"29",X"7B",
		X"FE",X"FC",X"30",X"1E",X"FE",X"07",X"38",X"1A",X"7A",X"CB",X"41",X"28",X"03",X"ED",X"44",X"57",
		X"7B",X"CB",X"51",X"28",X"03",X"ED",X"44",X"5F",X"92",X"FE",X"F6",X"30",X"11",X"FE",X"06",X"D0",
		X"18",X"0C",X"79",X"E6",X"03",X"4F",X"18",X"06",X"79",X"E6",X"0C",X"4F",X"18",X"00",X"06",X"00",
		X"E5",X"CD",X"E7",X"34",X"21",X"42",X"20",X"09",X"4E",X"21",X"44",X"29",X"09",X"09",X"09",X"DD",
		X"70",X"06",X"DD",X"70",X"08",X"7E",X"23",X"F3",X"DD",X"77",X"0A",X"7E",X"DD",X"77",X"0B",X"FB",
		X"23",X"DD",X"36",X"0C",X"01",X"46",X"23",X"4E",X"23",X"56",X"DD",X"7E",X"07",X"80",X"47",X"DD",
		X"7E",X"09",X"81",X"4F",X"E1",X"F3",X"72",X"23",X"36",X"00",X"23",X"70",X"23",X"71",X"23",X"72",
		X"23",X"36",X"05",X"23",X"70",X"23",X"71",X"FB",X"DD",X"E5",X"3E",X"0A",X"CD",X"6D",X"1E",X"DD",
		X"E1",X"2A",X"72",X"08",X"23",X"3A",X"4D",X"43",X"77",X"2B",X"CB",X"CE",X"E1",X"23",X"23",X"F1",
		X"C1",X"0E",X"10",X"E9",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"10",X"07",X"06",X"06",X"00",
		X"00",X"10",X"07",X"06",X"02",X"00",X"00",X"10",X"07",X"06",X"0A",X"00",X"00",X"10",X"07",X"06",
		X"08",X"00",X"00",X"10",X"00",X"06",X"09",X"00",X"00",X"10",X"00",X"06",X"01",X"00",X"00",X"10",
		X"00",X"06",X"05",X"00",X"00",X"10",X"07",X"01",X"04",X"00",X"CA",X"E1",X"46",X"23",X"5E",X"23",
		X"56",X"23",X"EB",X"CD",X"A3",X"29",X"EB",X"4E",X"CB",X"B9",X"CD",X"DB",X"29",X"47",X"3A",X"79",
		X"43",X"B7",X"20",X"03",X"13",X"18",X"01",X"1B",X"23",X"7E",X"B7",X"78",X"C2",X"87",X"29",X"23",
		X"E9",X"06",X"90",X"3A",X"79",X"43",X"B7",X"3E",X"07",X"20",X"15",X"A5",X"B0",X"D3",X"4B",X"CB",
		X"3C",X"CB",X"1D",X"CB",X"3C",X"CB",X"1D",X"CB",X"3C",X"CB",X"1D",X"01",X"00",X"64",X"09",X"C9",
		X"A5",X"B0",X"CB",X"DF",X"D3",X"4B",X"CB",X"3C",X"CB",X"1D",X"CB",X"3C",X"CB",X"1D",X"CB",X"3C",
		X"CB",X"1D",X"44",X"4D",X"21",X"FF",X"7F",X"B7",X"ED",X"42",X"C9",X"E5",X"21",X"00",X"00",X"06",
		X"00",X"09",X"29",X"29",X"29",X"09",X"01",X"1E",X"2F",X"09",X"D5",X"F5",X"EB",X"3A",X"79",X"43",
		X"B7",X"1A",X"20",X"26",X"B7",X"F2",X"FC",X"29",X"01",X"60",X"00",X"09",X"3E",X"09",X"01",X"1F",
		X"00",X"08",X"F1",X"F5",X"F3",X"D3",X"4B",X"1A",X"E6",X"7F",X"13",X"77",X"23",X"36",X"00",X"FB",
		X"09",X"08",X"3D",X"C2",X"01",X"2A",X"F1",X"D1",X"E1",X"C9",X"B7",X"F2",X"22",X"2A",X"01",X"A0",
		X"FF",X"09",X"3E",X"09",X"01",X"E1",X"FF",X"08",X"F1",X"F5",X"F3",X"D3",X"4B",X"1A",X"E6",X"7F",
		X"13",X"77",X"2B",X"36",X"00",X"FB",X"09",X"08",X"3D",X"C2",X"27",X"2A",X"F1",X"D1",X"E1",X"C9",
		X"C5",X"06",X"00",X"EB",X"CD",X"A3",X"29",X"EB",X"08",X"C1",X"CB",X"81",X"78",X"3D",X"20",X"02",
		X"CB",X"C1",X"7E",X"CB",X"40",X"20",X"09",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"2B",
		X"23",X"E6",X"0F",X"20",X"08",X"CB",X"41",X"20",X"06",X"3E",X"20",X"18",X"0A",X"CB",X"C1",X"C6",
		X"30",X"FE",X"3A",X"38",X"02",X"C6",X"07",X"E5",X"C5",X"4F",X"08",X"CD",X"DB",X"29",X"08",X"C1",
		X"E1",X"3A",X"79",X"43",X"B7",X"20",X"03",X"13",X"18",X"01",X"1B",X"10",X"BF",X"C9",X"C5",X"D1",
		X"CD",X"0E",X"20",X"CD",X"22",X"1E",X"DD",X"E5",X"CD",X"59",X"1E",X"DD",X"E1",X"2A",X"47",X"43",
		X"7D",X"FE",X"18",X"30",X"04",X"2E",X"02",X"18",X"06",X"FE",X"E6",X"38",X"02",X"2E",X"F8",X"7C",
		X"FE",X"B4",X"38",X"02",X"26",X"A0",X"DD",X"75",X"07",X"DD",X"74",X"09",X"3A",X"4C",X"43",X"47",
		X"3A",X"72",X"43",X"80",X"47",X"3A",X"4B",X"43",X"80",X"32",X"4E",X"43",X"DD",X"E5",X"3E",X"28",
		X"CD",X"6D",X"1E",X"DD",X"E1",X"21",X"4E",X"43",X"35",X"20",X"F1",X"CD",X"DE",X"2B",X"21",X"0B",
		X"12",X"DD",X"75",X"0A",X"DD",X"74",X"0B",X"DD",X"36",X"0C",X"01",X"DD",X"36",X"0D",X"02",X"DD",
		X"36",X"00",X"06",X"AF",X"CD",X"39",X"2B",X"DD",X"E5",X"C5",X"3E",X"28",X"CD",X"6D",X"1E",X"C1",
		X"DD",X"E1",X"FD",X"2A",X"76",X"08",X"C5",X"FD",X"7E",X"07",X"C6",X"02",X"DD",X"96",X"07",X"57",
		X"06",X"00",X"28",X"06",X"06",X"01",X"38",X"02",X"06",X"02",X"FD",X"7E",X"09",X"DD",X"96",X"09",
		X"5F",X"0E",X"00",X"28",X"06",X"0E",X"04",X"38",X"02",X"0E",X"08",X"78",X"81",X"C1",X"CD",X"39",
		X"2B",X"3E",X"04",X"CD",X"54",X"2B",X"C3",X"02",X"2B",X"E6",X"0F",X"B9",X"C8",X"4F",X"06",X"00",
		X"50",X"21",X"42",X"20",X"09",X"5E",X"21",X"19",X"25",X"19",X"7E",X"23",X"DD",X"77",X"06",X"7E",
		X"DD",X"77",X"08",X"C9",X"2A",X"72",X"08",X"36",X"82",X"23",X"77",X"DD",X"E5",X"E5",X"C5",X"CD",
		X"78",X"1E",X"C1",X"E1",X"DD",X"E1",X"DD",X"CB",X"00",X"7E",X"C9",X"D5",X"CD",X"78",X"26",X"D1",
		X"07",X"07",X"EE",X"09",X"E6",X"0F",X"90",X"FA",X"7C",X"2B",X"18",X"FA",X"80",X"28",X"0C",X"47",
		X"7E",X"CB",X"7F",X"20",X"03",X"23",X"18",X"F8",X"23",X"10",X"F5",X"7E",X"47",X"E6",X"7F",X"12",
		X"13",X"CB",X"78",X"23",X"28",X"F5",X"C9",X"2A",X"98",X"08",X"7C",X"B5",X"C0",X"21",X"9B",X"08",
		X"35",X"C0",X"CD",X"78",X"26",X"07",X"07",X"E6",X"0C",X"C6",X"04",X"77",X"21",X"18",X"09",X"CD",
		X"78",X"26",X"E6",X"1F",X"F6",X"60",X"77",X"23",X"EB",X"21",X"2C",X"2C",X"06",X"06",X"CD",X"6B",
		X"2B",X"21",X"25",X"2C",X"06",X"04",X"3A",X"9A",X"08",X"B7",X"20",X"03",X"23",X"23",X"05",X"CD",
		X"6B",X"2B",X"EB",X"36",X"47",X"23",X"36",X"FF",X"21",X"18",X"09",X"C3",X"1B",X"2C",X"21",X"4A",
		X"2C",X"C3",X"1B",X"2C",X"3A",X"71",X"43",X"B7",X"20",X"29",X"21",X"18",X"09",X"CD",X"78",X"26",
		X"E6",X"07",X"F6",X"70",X"77",X"23",X"EB",X"21",X"28",X"2C",X"06",X"02",X"CD",X"6B",X"2B",X"21",
		X"32",X"2C",X"06",X"01",X"CD",X"6B",X"2B",X"EB",X"36",X"44",X"23",X"36",X"FF",X"21",X"18",X"09",
		X"AF",X"18",X"05",X"21",X"35",X"2C",X"3E",X"FF",X"32",X"9A",X"08",X"22",X"98",X"08",X"C9",X"21",
		X"40",X"2C",X"AF",X"18",X"F3",X"0A",X"98",X"8C",X"0A",X"8F",X"0A",X"92",X"86",X"83",X"82",X"95",
		X"85",X"81",X"16",X"17",X"94",X"73",X"18",X"47",X"1B",X"73",X"19",X"1A",X"1B",X"1C",X"47",X"FF",
		X"7B",X"04",X"0A",X"0F",X"7D",X"04",X"0A",X"12",X"47",X"FF",X"7B",X"12",X"08",X"12",X"08",X"47",
		X"FF",X"CD",X"34",X"23",X"E5",X"23",X"23",X"EB",X"21",X"C4",X"08",X"0E",X"03",X"06",X"0C",X"1A",
		X"E6",X"0F",X"28",X"06",X"CD",X"B3",X"2D",X"3D",X"20",X"FA",X"05",X"1A",X"E6",X"F0",X"28",X"07",
		X"CD",X"B3",X"2D",X"D6",X"10",X"20",X"F9",X"05",X"1B",X"0D",X"20",X"E3",X"0E",X"0A",X"11",X"02",
		X"43",X"E1",X"E5",X"D5",X"06",X"03",X"1A",X"BE",X"38",X"11",X"20",X"04",X"13",X"23",X"10",X"F6",
		X"D1",X"21",X"06",X"00",X"19",X"EB",X"E1",X"0D",X"20",X"E8",X"C9",X"D1",X"D5",X"06",X"00",X"0D",
		X"28",X"14",X"21",X"00",X"00",X"09",X"29",X"09",X"29",X"E5",X"19",X"2B",X"54",X"5D",X"01",X"06",
		X"00",X"09",X"EB",X"C1",X"ED",X"B8",X"D1",X"E1",X"06",X"03",X"7E",X"23",X"12",X"13",X"10",X"FA",
		X"EB",X"E5",X"CD",X"4E",X"1A",X"CD",X"1C",X"36",X"CD",X"ED",X"1A",X"1B",X"00",X"D8",X"2D",X"3A",
		X"00",X"F4",X"2D",X"08",X"06",X"01",X"21",X"44",X"43",X"CD",X"4A",X"2A",X"CD",X"ED",X"1A",X"93",
		X"07",X"71",X"2E",X"13",X"2E",X"CB",X"2E",X"CD",X"7B",X"29",X"90",X"78",X"62",X"5F",X"5F",X"5F",
		X"00",X"CD",X"ED",X"1A",X"1B",X"2F",X"1B",X"2F",X"61",X"2F",X"BC",X"2F",X"06",X"00",X"21",X"78",
		X"60",X"CD",X"A3",X"29",X"EB",X"E1",X"E5",X"06",X"03",X"36",X"20",X"23",X"10",X"FB",X"E1",X"3E",
		X"1E",X"32",X"49",X"43",X"06",X"03",X"0E",X"41",X"C5",X"3A",X"79",X"43",X"CD",X"DB",X"29",X"D5",
		X"E5",X"3E",X"0F",X"CD",X"6D",X"1E",X"E1",X"D1",X"C1",X"FD",X"CB",X"00",X"CE",X"FD",X"36",X"01",
		X"3C",X"FD",X"7E",X"01",X"B7",X"20",X"0B",X"3A",X"49",X"43",X"3D",X"32",X"49",X"43",X"28",X"3A",
		X"18",X"E7",X"CD",X"CE",X"2D",X"CB",X"67",X"20",X"46",X"71",X"C5",X"3A",X"79",X"43",X"B7",X"01",
		X"40",X"00",X"28",X"03",X"01",X"C0",X"FF",X"D5",X"EB",X"09",X"EB",X"3A",X"79",X"43",X"F6",X"90",
		X"0E",X"5F",X"CD",X"DB",X"29",X"D1",X"C1",X"23",X"3A",X"79",X"43",X"B7",X"13",X"28",X"02",X"1B",
		X"1B",X"CD",X"CE",X"2D",X"CB",X"67",X"28",X"F9",X"10",X"9E",X"21",X"02",X"43",X"11",X"DC",X"08",
		X"06",X"1E",X"7E",X"23",X"12",X"13",X"07",X"07",X"07",X"07",X"12",X"13",X"10",X"F4",X"C9",X"CD",
		X"CE",X"2D",X"2F",X"CB",X"47",X"28",X"04",X"3E",X"FF",X"18",X"07",X"CB",X"4F",X"CA",X"31",X"2D",
		X"3E",X"01",X"81",X"FE",X"40",X"20",X"02",X"3E",X"5A",X"FE",X"5B",X"20",X"02",X"3E",X"41",X"4F",
		X"C3",X"18",X"2D",X"F5",X"C5",X"D5",X"E5",X"16",X"00",X"58",X"1D",X"19",X"0E",X"10",X"7E",X"E6",
		X"F0",X"81",X"27",X"77",X"30",X"03",X"2B",X"10",X"F5",X"E1",X"D1",X"C1",X"F1",X"C9",X"3A",X"79",
		X"43",X"B7",X"DB",X"48",X"C8",X"DB",X"4A",X"C9",X"CD",X"7B",X"29",X"90",X"20",X"08",X"47",X"72",
		X"61",X"74",X"75",X"6C",X"69",X"65",X"72",X"65",X"2C",X"20",X"53",X"70",X"69",X"65",X"6C",X"65",
		X"72",X"20",X"00",X"C9",X"CD",X"7B",X"29",X"90",X"20",X"08",X"46",X"65",X"6C",X"69",X"63",X"69",
		X"74",X"61",X"63",X"69",X"6F",X"6E",X"65",X"73",X"20",X"6A",X"75",X"67",X"61",X"64",X"6F",X"72",
		X"20",X"00",X"C9",X"CD",X"7B",X"29",X"90",X"08",X"20",X"56",X"6F",X"75",X"73",X"20",X"61",X"76",
		X"65",X"7A",X"20",X"6A",X"6F",X"69",X"6E",X"74",X"20",X"6C",X"65",X"73",X"20",X"69",X"6D",X"6D",
		X"6F",X"72",X"74",X"65",X"6C",X"73",X"00",X"CD",X"7B",X"29",X"90",X"08",X"30",X"64",X"75",X"20",
		X"70",X"61",X"6E",X"74",X"68",X"65",X"6F",X"6E",X"20",X"42",X"45",X"52",X"5A",X"45",X"52",X"4B",
		X"2E",X"00",X"CD",X"7B",X"29",X"90",X"08",X"50",X"49",X"6E",X"73",X"63",X"72",X"69",X"72",X"65",
		X"20",X"76",X"6F",X"73",X"20",X"69",X"6E",X"69",X"74",X"69",X"61",X"6C",X"65",X"73",X"3A",X"00",
		X"C9",X"CD",X"7B",X"29",X"90",X"08",X"20",X"44",X"61",X"73",X"20",X"57",X"61",X"72",X"20",X"65",
		X"69",X"6E",X"20",X"52",X"75",X"68",X"6D",X"76",X"6F",X"6C",X"6C",X"65",X"72",X"20",X"53",X"69",
		X"65",X"67",X"21",X"00",X"CD",X"7B",X"29",X"90",X"08",X"40",X"54",X"72",X"61",X"67",X"20",X"44",
		X"65",X"69",X"6E",X"65",X"6E",X"20",X"4E",X"61",X"6D",X"65",X"6E",X"20",X"69",X"6E",X"20",X"64",
		X"69",X"65",X"00",X"CD",X"7B",X"29",X"90",X"08",X"50",X"48",X"65",X"6C",X"64",X"65",X"6E",X"6C",
		X"69",X"73",X"74",X"65",X"20",X"65",X"69",X"6E",X"21",X"00",X"C9",X"CD",X"7B",X"29",X"90",X"04",
		X"20",X"53",X"65",X"20",X"70",X"75",X"6E",X"74",X"61",X"6A",X"65",X"20",X"65",X"73",X"74",X"61",
		X"20",X"65",X"6E",X"74",X"72",X"65",X"20",X"6C",X"6F",X"73",X"20",X"64",X"69",X"65",X"7A",X"00",
		X"CD",X"7B",X"29",X"90",X"08",X"30",X"6D",X"65",X"6A",X"6F",X"72",X"65",X"73",X"2E",X"00",X"CD",
		X"7B",X"29",X"90",X"18",X"50",X"45",X"6E",X"74",X"72",X"65",X"20",X"73",X"75",X"73",X"20",X"69",
		X"6E",X"69",X"63",X"69",X"61",X"6C",X"65",X"73",X"3A",X"00",X"C9",X"CD",X"7B",X"29",X"90",X"08",
		X"80",X"4D",X"6F",X"76",X"65",X"20",X"73",X"74",X"69",X"63",X"6B",X"20",X"74",X"6F",X"20",X"63",
		X"68",X"61",X"6E",X"67",X"65",X"20",X"6C",X"65",X"74",X"74",X"65",X"72",X"00",X"CD",X"7B",X"29",
		X"90",X"08",X"90",X"74",X"68",X"65",X"6E",X"20",X"70",X"72",X"65",X"73",X"73",X"20",X"46",X"49",
		X"52",X"45",X"20",X"74",X"6F",X"20",X"73",X"74",X"6F",X"72",X"65",X"20",X"69",X"74",X"2E",X"00",
		X"C9",X"CD",X"7B",X"29",X"90",X"04",X"80",X"50",X"6F",X"75",X"73",X"73",X"65",X"7A",X"20",X"62",
		X"61",X"74",X"6F",X"6E",X"6E",X"65",X"74",X"20",X"70",X"6F",X"75",X"72",X"20",X"76",X"6F",X"73",
		X"00",X"CD",X"7B",X"29",X"90",X"04",X"90",X"69",X"6E",X"69",X"74",X"69",X"61",X"6C",X"65",X"73",
		X"2E",X"20",X"50",X"6F",X"75",X"73",X"73",X"65",X"7A",X"20",X"46",X"49",X"52",X"45",X"20",X"71",
		X"75",X"61",X"6E",X"64",X"00",X"CD",X"7B",X"29",X"90",X"04",X"A0",X"6C",X"65",X"74",X"74",X"72",
		X"65",X"20",X"63",X"6F",X"72",X"72",X"65",X"63",X"74",X"65",X"00",X"C9",X"CD",X"7B",X"29",X"90",
		X"04",X"80",X"4D",X"6F",X"76",X"69",X"65",X"6E",X"64",X"6F",X"20",X"6C",X"61",X"20",X"70",X"61",
		X"6C",X"61",X"6E",X"63",X"61",X"20",X"70",X"61",X"72",X"61",X"00",X"CD",X"7B",X"29",X"90",X"04",
		X"90",X"63",X"61",X"6D",X"62",X"69",X"61",X"72",X"20",X"6C",X"61",X"73",X"20",X"6C",X"65",X"74",
		X"72",X"61",X"73",X"2C",X"20",X"6C",X"75",X"65",X"67",X"6F",X"00",X"CD",X"7B",X"29",X"90",X"04",
		X"A0",X"61",X"70",X"6C",X"61",X"73",X"74",X"65",X"20",X"65",X"6C",X"20",X"62",X"6F",X"74",X"6F",
		X"6E",X"20",X"64",X"65",X"20",X"64",X"69",X"73",X"70",X"61",X"72",X"6F",X"00",X"CD",X"7B",X"29",
		X"90",X"04",X"B0",X"70",X"61",X"72",X"61",X"20",X"72",X"65",X"74",X"65",X"6E",X"65",X"72",X"6C",
		X"61",X"73",X"2E",X"00",X"C9",X"00",X"3E",X"41",X"5D",X"51",X"5D",X"41",X"3E",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"10",
		X"14",X"14",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"14",X"14",X"14",X"7F",X"14",X"7F",X"14",
		X"14",X"14",X"14",X"7F",X"54",X"54",X"7F",X"15",X"15",X"7F",X"14",X"20",X"51",X"22",X"04",X"08",
		X"10",X"22",X"45",X"02",X"00",X"18",X"24",X"28",X"10",X"29",X"46",X"46",X"39",X"08",X"08",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"08",X"10",X"10",X"10",X"10",X"10",X"08",X"04",X"10",
		X"08",X"04",X"04",X"04",X"04",X"04",X"08",X"10",X"00",X"00",X"08",X"2A",X"1C",X"1C",X"2A",X"08",
		X"00",X"00",X"00",X"08",X"08",X"3E",X"08",X"08",X"00",X"00",X"80",X"00",X"00",X"00",X"18",X"18",
		X"08",X"10",X"00",X"00",X"00",X"00",X"00",X"3E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"18",X"18",X"00",X"00",X"01",X"02",X"04",X"08",X"10",X"20",X"40",X"1C",X"22",
		X"41",X"41",X"41",X"41",X"41",X"22",X"1C",X"08",X"18",X"08",X"08",X"08",X"08",X"08",X"08",X"1C",
		X"3E",X"41",X"01",X"01",X"3E",X"40",X"40",X"40",X"7F",X"3E",X"41",X"01",X"01",X"1E",X"01",X"01",
		X"41",X"3E",X"02",X"06",X"0A",X"12",X"22",X"7F",X"02",X"02",X"02",X"7F",X"40",X"40",X"40",X"7E",
		X"01",X"01",X"41",X"3E",X"3E",X"41",X"40",X"40",X"7E",X"41",X"41",X"41",X"3E",X"7F",X"01",X"02",
		X"02",X"04",X"04",X"08",X"08",X"08",X"3E",X"41",X"41",X"41",X"3E",X"41",X"41",X"41",X"3E",X"3E",
		X"41",X"41",X"41",X"3F",X"01",X"01",X"41",X"3E",X"00",X"00",X"00",X"18",X"18",X"00",X"00",X"18",
		X"18",X"98",X"18",X"00",X"00",X"18",X"18",X"08",X"10",X"00",X"02",X"04",X"08",X"10",X"20",X"10",
		X"08",X"04",X"02",X"00",X"00",X"00",X"3E",X"00",X"3E",X"00",X"00",X"00",X"20",X"10",X"08",X"04",
		X"02",X"04",X"08",X"10",X"20",X"1C",X"22",X"02",X"02",X"04",X"08",X"08",X"00",X"08",X"3E",X"41",
		X"4F",X"49",X"49",X"4F",X"40",X"40",X"3F",X"3E",X"41",X"41",X"41",X"7F",X"41",X"41",X"41",X"41",
		X"7E",X"41",X"41",X"41",X"7E",X"41",X"41",X"41",X"7E",X"3E",X"41",X"40",X"40",X"40",X"40",X"40",
		X"41",X"3E",X"7E",X"41",X"41",X"41",X"41",X"41",X"41",X"41",X"7E",X"7F",X"40",X"40",X"40",X"7C",
		X"40",X"40",X"40",X"7F",X"7F",X"40",X"40",X"40",X"7C",X"40",X"40",X"40",X"40",X"3E",X"41",X"40",
		X"40",X"47",X"41",X"41",X"41",X"3F",X"41",X"41",X"41",X"41",X"7F",X"41",X"41",X"41",X"41",X"1C",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"1C",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"41",
		X"3E",X"41",X"42",X"44",X"48",X"50",X"68",X"44",X"42",X"41",X"40",X"40",X"40",X"40",X"40",X"40",
		X"40",X"40",X"7F",X"41",X"63",X"55",X"49",X"41",X"41",X"41",X"41",X"41",X"41",X"61",X"51",X"49",
		X"45",X"43",X"41",X"41",X"41",X"3E",X"41",X"41",X"41",X"41",X"41",X"41",X"41",X"3E",X"7E",X"41",
		X"41",X"41",X"7E",X"40",X"40",X"40",X"40",X"3E",X"41",X"41",X"41",X"41",X"41",X"45",X"42",X"3D",
		X"7E",X"41",X"41",X"41",X"7E",X"48",X"44",X"42",X"41",X"3E",X"41",X"40",X"40",X"3E",X"01",X"01",
		X"41",X"3E",X"7F",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"41",X"41",X"41",X"41",X"41",
		X"41",X"41",X"41",X"3E",X"41",X"41",X"41",X"22",X"22",X"14",X"14",X"08",X"08",X"41",X"41",X"41",
		X"41",X"41",X"49",X"55",X"63",X"41",X"41",X"41",X"22",X"14",X"08",X"14",X"22",X"41",X"41",X"41",
		X"41",X"22",X"14",X"08",X"08",X"08",X"08",X"08",X"7F",X"01",X"02",X"04",X"08",X"10",X"20",X"40",
		X"7F",X"3C",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"3C",X"00",X"00",X"40",X"20",X"10",X"08",
		X"04",X"02",X"01",X"3C",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"3C",X"08",X"14",X"22",X"41",
		X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"18",X"18",
		X"10",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3A",X"46",X"42",X"42",X"46",X"3A",
		X"40",X"40",X"40",X"5C",X"62",X"42",X"42",X"62",X"5C",X"00",X"00",X"00",X"3C",X"42",X"40",X"40",
		X"42",X"3C",X"02",X"02",X"02",X"3A",X"46",X"42",X"42",X"46",X"3A",X"00",X"00",X"00",X"3C",X"42",
		X"7E",X"40",X"40",X"3C",X"0C",X"12",X"10",X"10",X"38",X"10",X"10",X"10",X"10",X"BA",X"46",X"42",
		X"42",X"46",X"3A",X"02",X"42",X"3C",X"40",X"40",X"40",X"7C",X"42",X"42",X"42",X"42",X"42",X"00",
		X"08",X"00",X"08",X"08",X"08",X"08",X"08",X"08",X"84",X"04",X"04",X"04",X"04",X"04",X"04",X"44",
		X"38",X"40",X"40",X"40",X"44",X"48",X"50",X"70",X"48",X"44",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"00",X"00",X"00",X"76",X"49",X"49",X"49",X"49",X"49",X"00",X"00",X"00",X"7C",
		X"42",X"42",X"42",X"42",X"42",X"00",X"00",X"00",X"3C",X"42",X"42",X"42",X"42",X"3C",X"DC",X"62",
		X"42",X"42",X"62",X"5C",X"40",X"40",X"40",X"BA",X"46",X"42",X"42",X"46",X"3A",X"02",X"02",X"02",
		X"00",X"00",X"00",X"5C",X"62",X"40",X"40",X"40",X"40",X"00",X"00",X"00",X"3C",X"42",X"30",X"0C",
		X"42",X"3C",X"00",X"10",X"10",X"7C",X"10",X"10",X"10",X"10",X"10",X"00",X"00",X"00",X"42",X"42",
		X"42",X"42",X"42",X"3C",X"00",X"00",X"00",X"44",X"44",X"44",X"44",X"28",X"10",X"00",X"00",X"00",
		X"41",X"41",X"41",X"49",X"49",X"36",X"00",X"00",X"00",X"42",X"24",X"18",X"18",X"24",X"42",X"C2",
		X"42",X"42",X"42",X"46",X"3A",X"02",X"42",X"3C",X"00",X"00",X"00",X"7E",X"04",X"08",X"10",X"20",
		X"7E",X"0C",X"10",X"10",X"10",X"20",X"10",X"10",X"10",X"0C",X"08",X"08",X"08",X"00",X"00",X"08",
		X"08",X"08",X"00",X"18",X"04",X"04",X"04",X"02",X"04",X"04",X"04",X"18",X"30",X"49",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"55",X"2A",X"55",X"2A",X"55",X"2A",X"55",X"2A",X"55",X"08",X"00",
		X"1C",X"2A",X"08",X"08",X"14",X"22",X"00",X"21",X"89",X"08",X"F5",X"3E",X"FF",X"BE",X"38",X"09",
		X"D3",X"4D",X"77",X"21",X"29",X"34",X"22",X"85",X"08",X"F1",X"D3",X"4C",X"C9",X"21",X"89",X"08",
		X"F5",X"3E",X"00",X"BE",X"38",X"09",X"D3",X"4D",X"77",X"21",X"D3",X"33",X"22",X"85",X"08",X"F1",
		X"D3",X"4C",X"C9",X"0E",X"04",X"81",X"08",X"00",X"05",X"06",X"06",X"0E",X"03",X"78",X"08",X"92",
		X"92",X"92",X"0F",X"03",X"7B",X"08",X"32",X"00",X"32",X"00",X"32",X"00",X"06",X"04",X"95",X"08",
		X"06",X"32",X"93",X"08",X"01",X"0B",X"0F",X"00",X"7B",X"08",X"0B",X"11",X"00",X"7D",X"08",X"0B",
		X"10",X"00",X"7F",X"08",X"03",X"93",X"08",X"EC",X"07",X"32",X"00",X"7B",X"08",X"03",X"95",X"08",
		X"DF",X"06",X"FA",X"93",X"08",X"01",X"0B",X"0A",X"00",X"7B",X"08",X"0B",X"0D",X"00",X"7D",X"08",
		X"0B",X"0F",X"00",X"7F",X"08",X"03",X"93",X"08",X"EC",X"0E",X"03",X"78",X"08",X"00",X"00",X"00",
		X"0E",X"04",X"82",X"08",X"00",X"00",X"00",X"00",X"00",X"21",X"89",X"08",X"F5",X"3E",X"03",X"BE",
		X"38",X"09",X"D3",X"4D",X"77",X"21",X"4F",X"34",X"22",X"85",X"08",X"F1",X"D3",X"4C",X"C9",X"0E",
		X"04",X"81",X"08",X"00",X"06",X"07",X"07",X"0E",X"03",X"78",X"08",X"90",X"90",X"90",X"06",X"10",
		X"93",X"08",X"07",X"AC",X"00",X"7B",X"08",X"0F",X"02",X"7D",X"08",X"14",X"00",X"0A",X"00",X"06",
		X"19",X"95",X"08",X"01",X"0A",X"05",X"7D",X"08",X"0A",X"1E",X"7F",X"08",X"03",X"95",X"08",X"F3",
		X"0A",X"FC",X"7B",X"08",X"03",X"93",X"08",X"DF",X"02",X"9F",X"21",X"89",X"08",X"F5",X"3E",X"01",
		X"BE",X"38",X"09",X"D3",X"4D",X"77",X"21",X"A0",X"34",X"22",X"85",X"08",X"F1",X"D3",X"4C",X"C9",
		X"0E",X"03",X"78",X"08",X"82",X"80",X"80",X"0E",X"04",X"81",X"08",X"03",X"07",X"07",X"07",X"0F",
		X"03",X"7B",X"08",X"01",X"00",X"01",X"00",X"05",X"00",X"01",X"0E",X"03",X"78",X"08",X"92",X"90",
		X"90",X"06",X"37",X"95",X"08",X"06",X"06",X"93",X"08",X"01",X"03",X"93",X"08",X"FB",X"0B",X"01",
		X"00",X"7B",X"08",X"03",X"95",X"08",X"EE",X"0E",X"03",X"78",X"08",X"00",X"00",X"00",X"0E",X"04",
		X"81",X"08",X"00",X"00",X"00",X"00",X"00",X"21",X"89",X"08",X"F5",X"3E",X"01",X"BE",X"38",X"09",
		X"D3",X"4D",X"77",X"21",X"FD",X"34",X"22",X"85",X"08",X"F1",X"D3",X"4C",X"C9",X"0E",X"03",X"78",
		X"08",X"92",X"92",X"92",X"0E",X"04",X"81",X"08",X"00",X"06",X"06",X"07",X"0F",X"03",X"7B",X"08",
		X"14",X"00",X"2D",X"00",X"5A",X"00",X"06",X"04",X"95",X"08",X"06",X"50",X"93",X"08",X"01",X"0B",
		X"08",X"00",X"7B",X"08",X"0B",X"11",X"00",X"7D",X"08",X"0B",X"2F",X"00",X"7F",X"08",X"03",X"93",
		X"08",X"EC",X"03",X"95",X"08",X"E4",X"02",X"9F",X"21",X"89",X"08",X"F5",X"3E",X"02",X"BE",X"38",
		X"09",X"D3",X"4D",X"77",X"21",X"4E",X"35",X"22",X"85",X"08",X"F1",X"D3",X"4C",X"C9",X"0E",X"04",
		X"81",X"08",X"00",X"07",X"07",X"07",X"0E",X"03",X"78",X"08",X"92",X"92",X"92",X"0F",X"03",X"7B",
		X"08",X"C8",X"00",X"3C",X"00",X"28",X"00",X"06",X"14",X"95",X"08",X"06",X"14",X"93",X"08",X"01",
		X"0B",X"14",X"00",X"7B",X"08",X"0B",X"06",X"00",X"7D",X"08",X"0B",X"04",X"00",X"7F",X"08",X"03",
		X"93",X"08",X"EC",X"06",X"14",X"93",X"08",X"01",X"0B",X"EC",X"FF",X"7B",X"08",X"0B",X"FA",X"FF",
		X"7D",X"08",X"0B",X"FC",X"FF",X"7F",X"08",X"03",X"93",X"08",X"EC",X"03",X"95",X"08",X"CC",X"0E",
		X"03",X"78",X"08",X"00",X"00",X"00",X"0E",X"04",X"81",X"08",X"00",X"00",X"00",X"00",X"00",X"CD",
		X"57",X"36",X"00",X"00",X"04",X"20",X"AA",X"CD",X"57",X"36",X"80",X"00",X"01",X"20",X"FF",X"CD",
		X"57",X"36",X"A0",X"00",X"29",X"20",X"11",X"CD",X"57",X"36",X"A0",X"00",X"29",X"09",X"99",X"CD",
		X"57",X"36",X"A9",X"00",X"29",X"08",X"BB",X"CD",X"57",X"36",X"B0",X"00",X"29",X"10",X"55",X"CD",
		X"57",X"36",X"C0",X"05",X"0A",X"20",X"77",X"CD",X"57",X"36",X"80",X"06",X"04",X"0A",X"AA",X"CD",
		X"57",X"36",X"96",X"06",X"04",X"0A",X"DD",X"C9",X"CD",X"57",X"36",X"00",X"00",X"38",X"20",X"FF",
		X"C9",X"CD",X"57",X"36",X"E0",X"05",X"04",X"20",X"33",X"C9",X"CD",X"57",X"36",X"E0",X"05",X"04",
		X"20",X"99",X"C9",X"CD",X"57",X"36",X"E0",X"05",X"04",X"20",X"66",X"C9",X"CD",X"57",X"36",X"00",
		X"00",X"08",X"20",X"BB",X"CD",X"57",X"36",X"00",X"01",X"10",X"20",X"66",X"CD",X"57",X"36",X"00",
		X"03",X"04",X"20",X"FF",X"CD",X"57",X"36",X"80",X"03",X"1C",X"20",X"AA",X"C9",X"CD",X"57",X"36",
		X"00",X"00",X"2F",X"20",X"CC",X"CD",X"57",X"36",X"E0",X"05",X"09",X"20",X"AA",X"C9",X"CD",X"57",
		X"36",X"00",X"00",X"34",X"20",X"44",X"C9",X"E1",X"5E",X"23",X"56",X"23",X"E5",X"3A",X"79",X"43",
		X"B7",X"20",X"06",X"21",X"00",X"81",X"19",X"18",X"05",X"21",X"FF",X"87",X"ED",X"52",X"EB",X"E1",
		X"4E",X"23",X"08",X"7E",X"23",X"08",X"B7",X"7E",X"23",X"E5",X"EB",X"20",X"11",X"11",X"20",X"00",
		X"08",X"47",X"08",X"E5",X"77",X"23",X"10",X"FC",X"E1",X"19",X"0D",X"20",X"F3",X"C9",X"11",X"E0",
		X"FF",X"08",X"47",X"08",X"E5",X"77",X"2B",X"10",X"FC",X"E1",X"19",X"0D",X"20",X"F3",X"C9",X"CD",
		X"57",X"36",X"80",X"06",X"04",X"20",X"77",X"CD",X"E7",X"35",X"CD",X"34",X"23",X"EB",X"01",X"05",
		X"00",X"13",X"1A",X"08",X"1B",X"1A",X"B7",X"21",X"94",X"37",X"28",X"0F",X"E6",X"0F",X"67",X"08",
		X"E6",X"F0",X"B4",X"07",X"07",X"07",X"07",X"21",X"BC",X"37",X"08",X"08",X"BE",X"38",X"06",X"08",
		X"09",X"7E",X"B7",X"20",X"F6",X"23",X"7E",X"23",X"32",X"4B",X"43",X"7E",X"23",X"32",X"7A",X"43",
		X"7E",X"23",X"32",X"4D",X"43",X"4E",X"3A",X"79",X"43",X"B7",X"DD",X"21",X"00",X"81",X"21",X"00",
		X"44",X"28",X"07",X"DD",X"21",X"80",X"81",X"21",X"00",X"46",X"3E",X"34",X"08",X"06",X"20",X"7E",
		X"23",X"5F",X"E6",X"44",X"57",X"7B",X"2F",X"A1",X"B2",X"DD",X"77",X"00",X"DD",X"23",X"10",X"EF",
		X"11",X"60",X"00",X"19",X"08",X"3D",X"20",X"E4",X"C9",X"CB",X"5E",X"CA",X"3C",X"37",X"CB",X"9E",
		X"E5",X"2A",X"40",X"09",X"11",X"42",X"09",X"3E",X"05",X"08",X"06",X"02",X"1A",X"13",X"77",X"23",
		X"10",X"FA",X"01",X"1E",X"00",X"09",X"08",X"3D",X"C2",X"29",X"37",X"E1",X"CB",X"66",X"C8",X"CB",
		X"DE",X"E5",X"11",X"07",X"00",X"19",X"5E",X"23",X"23",X"3A",X"79",X"43",X"B7",X"7E",X"28",X"0A",
		X"ED",X"44",X"C6",X"D0",X"08",X"3E",X"F7",X"93",X"5F",X"08",X"CB",X"3F",X"CB",X"3F",X"67",X"6B",
		X"CB",X"3C",X"CB",X"1D",X"CB",X"3C",X"CB",X"1D",X"CB",X"3C",X"CB",X"1D",X"01",X"00",X"81",X"09",
		X"22",X"40",X"09",X"3A",X"78",X"43",X"11",X"1E",X"00",X"FD",X"21",X"42",X"09",X"0E",X"05",X"06",
		X"02",X"08",X"7E",X"FD",X"77",X"00",X"FD",X"23",X"08",X"77",X"23",X"10",X"F4",X"19",X"0D",X"C2",
		X"7F",X"37",X"E1",X"C9",X"03",X"00",X"00",X"50",X"33",X"15",X"01",X"00",X"50",X"99",X"30",X"02",
		X"00",X"14",X"66",X"45",X"03",X"00",X"0A",X"AA",X"60",X"04",X"00",X"0A",X"55",X"75",X"05",X"00",
		X"0F",X"BB",X"90",X"01",X"01",X"3C",X"FF",X"00",X"01",X"01",X"32",X"FF",X"10",X"01",X"01",X"2D",
		X"FF",X"11",X"02",X"02",X"23",X"66",X"13",X"03",X"03",X"19",X"DD",X"15",X"04",X"04",X"14",X"77",
		X"17",X"05",X"05",X"0F",X"33",X"19",X"05",X"05",X"0A",X"99",X"00",X"05",X"05",X"05",X"EE",X"81",
		X"94",X"0C",X"02",X"AD",X"20",X"75",X"7A",X"0D",X"5F",X"40",X"93",X"D5",X"67",X"8A",X"49",X"14",
		X"F5",X"74",X"CF",X"80",X"21",X"2B",X"CA",X"CC",X"2B",X"3C",X"04",X"FB",X"AB",X"26",X"F8",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
