library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity MOONCR_1H is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of MOONCR_1H is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",X"00",X"02",X"02",X"FE",X"FE",X"42",X"02",X"00",X"00",
		X"62",X"F2",X"BA",X"9A",X"9E",X"CE",X"46",X"00",X"8C",X"DE",X"F2",X"B2",X"92",X"86",X"04",X"00",
		X"08",X"FE",X"FE",X"C8",X"68",X"38",X"18",X"00",X"1C",X"BE",X"A2",X"A2",X"A2",X"E6",X"E4",X"00",
		X"0C",X"9E",X"92",X"92",X"D2",X"7E",X"3C",X"00",X"C0",X"E0",X"B0",X"9E",X"8E",X"C0",X"C0",X"00",
		X"0C",X"6E",X"9A",X"9A",X"B2",X"F2",X"6C",X"00",X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",X"00",
		X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",
		X"44",X"C6",X"82",X"82",X"C6",X"7C",X"38",X"00",X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",
		X"82",X"92",X"92",X"92",X"FE",X"FE",X"00",X"00",X"80",X"90",X"90",X"90",X"90",X"FE",X"FE",X"00",
		X"9E",X"9E",X"92",X"82",X"C6",X"7C",X"38",X"00",X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",
		X"82",X"82",X"FE",X"FE",X"82",X"82",X"00",X"00",X"FC",X"FE",X"02",X"02",X"02",X"06",X"04",X"00",
		X"82",X"C6",X"6E",X"3C",X"18",X"FE",X"FE",X"00",X"02",X"02",X"02",X"02",X"FE",X"FE",X"00",X"00",
		X"FE",X"FE",X"70",X"38",X"70",X"FE",X"FE",X"00",X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",
		X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",X"00",X"70",X"F8",X"88",X"88",X"88",X"FE",X"FE",X"00",
		X"7A",X"FC",X"8E",X"8A",X"82",X"FE",X"7C",X"00",X"72",X"F6",X"9E",X"8C",X"88",X"FE",X"FE",X"00",
		X"0C",X"5E",X"D2",X"92",X"92",X"F6",X"64",X"00",X"80",X"80",X"FE",X"FE",X"80",X"80",X"00",X"00",
		X"FC",X"FE",X"02",X"02",X"02",X"FE",X"FC",X"00",X"F0",X"F8",X"1C",X"0E",X"1C",X"F8",X"F0",X"00",
		X"F8",X"FE",X"1C",X"38",X"1C",X"FE",X"F8",X"00",X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",
		X"C0",X"F0",X"1E",X"1E",X"F0",X"C0",X"00",X"00",X"C2",X"E2",X"F2",X"BA",X"9E",X"8E",X"86",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"F0",X"FB",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"D0",X"00",X"00",
		X"81",X"42",X"24",X"18",X"18",X"24",X"42",X"81",X"00",X"18",X"18",X"18",X"18",X"18",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",X"00",
		X"00",X"28",X"28",X"28",X"28",X"28",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"0A",X"08",X"08",X"10",X"20",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"10",X"08",X"08",X"0A",X"07",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"06",X"0C",X"18",X"3C",X"3E",X"BE",X"DE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BE",X"3E",X"3C",X"18",X"0C",X"06",X"02",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"01",X"00",X"C0",X"E0",X"E0",X"A0",X"C0",X"60",X"A0",
		X"01",X"03",X"03",X"01",X"07",X"0F",X"3F",X"FF",X"E0",X"80",X"60",X"F0",X"F8",X"FC",X"FE",X"FF",
		X"3F",X"0F",X"07",X"01",X"03",X"03",X"01",X"01",X"FE",X"FC",X"F8",X"F0",X"60",X"80",X"E0",X"A0",
		X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"60",X"C0",X"A0",X"E0",X"E0",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"54",X"D8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"3B",X"7D",X"E8",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",
		X"74",X"3F",X"08",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"00",X"3A",X"7D",X"EA",X"00",X"00",X"04",X"40",X"80",X"24",X"02",X"40",
		X"74",X"1A",X"00",X"00",X"02",X"00",X"00",X"00",X"28",X"14",X"00",X"10",X"00",X"20",X"00",X"00",
		X"00",X"40",X"80",X"20",X"40",X"11",X"19",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"16",X"10",X"00",X"18",X"0E",X"06",X"03",X"33",X"20",X"21",X"7E",X"7F",X"09",X"06",X"00",X"10",
		X"33",X"00",X"10",X"38",X"3C",X"66",X"6A",X"31",X"3D",X"3D",X"11",X"3F",X"3E",X"10",X"00",X"40",
		X"11",X"40",X"80",X"20",X"56",X"10",X"7F",X"7F",X"80",X"20",X"40",X"10",X"38",X"3C",X"6E",X"66",
		X"10",X"16",X"00",X"00",X"01",X"09",X"3B",X"0F",X"33",X"11",X"00",X"18",X"0E",X"06",X"03",X"33",
		X"06",X"00",X"0C",X"0C",X"0C",X"0C",X"0C",X"40",X"33",X"00",X"28",X"28",X"7F",X"7E",X"28",X"28",
		X"80",X"23",X"4F",X"1E",X"38",X"00",X"1E",X"07",X"00",X"0C",X"02",X"09",X"00",X"08",X"00",X"20",
		X"00",X"08",X"04",X"06",X"03",X"7F",X"7F",X"00",X"40",X"10",X"26",X"0C",X"18",X"7F",X"7F",X"00",
		X"00",X"02",X"07",X"0C",X"0B",X"03",X"03",X"17",X"00",X"20",X"20",X"00",X"80",X"C8",X"C8",X"E4",
		X"23",X"03",X"13",X"09",X"08",X"03",X"00",X"00",X"F0",X"E0",X"C4",X"E8",X"C0",X"20",X"C0",X"00",
		X"00",X"00",X"02",X"09",X"01",X"02",X"04",X"00",X"00",X"00",X"00",X"10",X"00",X"48",X"30",X"20",
		X"0E",X"14",X"01",X"03",X"04",X"01",X"00",X"00",X"68",X"04",X"40",X"20",X"10",X"00",X"00",X"00",
		X"00",X"04",X"04",X"00",X"02",X"65",X"1A",X"07",X"00",X"40",X"82",X"84",X"08",X"20",X"60",X"C0",
		X"09",X"05",X"06",X"21",X"02",X"12",X"24",X"00",X"90",X"C6",X"80",X"61",X"10",X"08",X"40",X"00",
		X"90",X"40",X"20",X"19",X"86",X"44",X"03",X"03",X"55",X"02",X"95",X"2A",X"44",X"C8",X"90",X"C3",
		X"77",X"CB",X"1B",X"0D",X"50",X"21",X"41",X"81",X"E0",X"E8",X"D4",X"86",X"01",X"48",X"24",X"02",
		X"04",X"10",X"48",X"20",X"00",X"81",X"43",X"07",X"20",X"08",X"12",X"04",X"00",X"81",X"C2",X"E0",
		X"07",X"43",X"81",X"00",X"20",X"48",X"10",X"04",X"E0",X"C2",X"81",X"00",X"04",X"12",X"08",X"20",
		X"04",X"10",X"48",X"20",X"00",X"81",X"43",X"07",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"A0",
		X"07",X"43",X"81",X"00",X"20",X"48",X"10",X"04",X"A0",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"09",X"24",X"10",X"00",X"40",X"21",X"03",X"07",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"00",
		X"47",X"83",X"01",X"40",X"90",X"20",X"00",X"08",X"A0",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"01",X"09",X"08",X"20",X"20",X"01",X"03",X"C7",X"40",X"00",X"00",X"00",X"00",X"80",X"C0",X"80",
		X"07",X"02",X"C1",X"00",X"40",X"80",X"00",X"20",X"80",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"09",X"08",X"00",X"60",X"01",X"03",X"C7",X"20",X"28",X"00",X"00",X"00",X"80",X"C0",X"A0",
		X"07",X"02",X"C1",X"00",X"40",X"00",X"00",X"00",X"80",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"04",X"20",X"10",X"80",X"41",X"03",X"07",X"48",X"90",X"04",X"00",X"00",X"80",X"C0",X"A0",
		X"C7",X"02",X"00",X"80",X"00",X"00",X"00",X"00",X"80",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"22",X"10",X"80",X"40",X"01",X"83",X"07",X"50",X"54",X"08",X"02",X"00",X"80",X"C0",X"E0",
		X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"22",X"10",X"40",X"20",X"81",X"03",X"07",X"20",X"44",X"08",X"02",X"04",X"81",X"C0",X"E0",
		X"05",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"04",X"10",X"48",X"20",X"00",X"81",X"43",X"07",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"80",
		X"07",X"43",X"81",X"00",X"20",X"48",X"10",X"04",X"80",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"02",X"08",X"24",X"10",X"00",X"40",X"21",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"03",X"21",X"40",X"00",X"10",X"24",X"08",X"02",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"08",X"24",X"10",X"40",X"21",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"03",X"21",X"40",X"10",X"24",X"08",X"02",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"08",X"14",X"08",X"31",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"31",X"08",X"14",X"08",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"04",X"08",X"10",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"10",X"08",X"04",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"04",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"04",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0F",X"0B",X"0B",
		X"07",X"0F",X"0D",X"04",X"0E",X"01",X"01",X"01",X"BF",X"9F",X"07",X"60",X"7C",X"7E",X"FE",X"FE",
		X"02",X"06",X"06",X"03",X"01",X"00",X"00",X"00",X"F7",X"7F",X"FF",X"F3",X"FF",X"7F",X"13",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"40",X"20",X"10",X"08",X"04",X"03",X"00",X"10",X"08",X"08",X"1C",X"0C",X"C0",X"20",
		X"01",X"02",X"02",X"01",X"00",X"00",X"00",X"00",X"E0",X"F0",X"70",X"06",X"0A",X"10",X"60",X"20",
		X"31",X"08",X"00",X"00",X"00",X"00",X"01",X"01",X"C1",X"20",X"18",X"08",X"48",X"C4",X"7B",X"00",
		X"01",X"06",X"0C",X"08",X"08",X"10",X"20",X"00",X"00",X"10",X"20",X"20",X"13",X"0C",X"00",X"00",
		X"00",X"80",X"40",X"30",X"08",X"05",X"07",X"01",X"80",X"40",X"20",X"10",X"63",X"90",X"0E",X"21",
		X"01",X"01",X"03",X"06",X"04",X"04",X"0B",X"3A",X"48",X"38",X"0E",X"1F",X"0F",X"07",X"01",X"D9",
		X"C5",X"02",X"00",X"06",X"02",X"05",X"0E",X"0E",X"3F",X"8F",X"07",X"02",X"08",X"15",X"C7",X"F5",
		X"0E",X"07",X"0F",X"18",X"30",X"20",X"40",X"00",X"74",X"A2",X"D9",X"0C",X"02",X"0C",X"0C",X"12",
		X"00",X"00",X"20",X"08",X"02",X"00",X"00",X"02",X"00",X"00",X"04",X"08",X"08",X"80",X"65",X"32",
		X"11",X"04",X"03",X"00",X"00",X"00",X"00",X"AA",X"18",X"0C",X"4B",X"20",X"03",X"80",X"C0",X"80",
		X"02",X"0C",X"00",X"01",X"00",X"04",X"10",X"42",X"58",X"83",X"32",X"10",X"21",X"80",X"02",X"08",
		X"01",X"00",X"04",X"00",X"10",X"00",X"40",X"00",X"00",X"17",X"09",X"16",X"20",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"81",X"C7",X"E9",X"E8",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"60",
		X"FE",X"FF",X"E7",X"C3",X"0F",X"1F",X"03",X"0F",X"30",X"30",X"30",X"B0",X"30",X"60",X"C0",X"C0",
		X"83",X"A2",X"18",X"0E",X"8F",X"9F",X"9F",X"FE",X"80",X"A0",X"D0",X"48",X"68",X"B0",X"00",X"00",
		X"FE",X"FE",X"7C",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"00",X"04",X"08",X"18",X"30",X"20",X"E0",X"40",
		X"00",X"00",X"71",X"12",X"11",X"16",X"04",X"84",X"00",X"00",X"80",X"60",X"10",X"08",X"08",X"10",
		X"40",X"21",X"22",X"40",X"20",X"CA",X"0F",X"03",X"78",X"9E",X"10",X"08",X"04",X"08",X"10",X"C0",
		X"23",X"41",X"00",X"A4",X"28",X"10",X"00",X"00",X"B0",X"30",X"30",X"1C",X"0C",X"04",X"02",X"00",
		X"00",X"0C",X"32",X"41",X"00",X"06",X"04",X"09",X"01",X"02",X"06",X"0C",X"38",X"3C",X"5C",X"A8",
		X"D3",X"C6",X"87",X"6B",X"F4",X"A0",X"08",X"CC",X"C0",X"C0",X"10",X"40",X"80",X"80",X"00",X"CF",
		X"EF",X"EE",X"79",X"28",X"84",X"91",X"0B",X"15",X"98",X"30",X"20",X"20",X"C0",X"00",X"40",X"F8",
		X"94",X"C4",X"28",X"D0",X"30",X"30",X"C0",X"00",X"70",X"28",X"64",X"C2",X"C1",X"00",X"00",X"00",
		X"00",X"01",X"00",X"42",X"04",X"20",X"84",X"60",X"00",X"00",X"10",X"00",X"00",X"00",X"80",X"00",
		X"22",X"50",X"1D",X"1D",X"01",X"C6",X"06",X"19",X"10",X"80",X"60",X"10",X"60",X"00",X"00",X"B2",
		X"38",X"84",X"01",X"22",X"00",X"10",X"08",X"02",X"00",X"00",X"40",X"10",X"80",X"20",X"00",X"08",
		X"10",X"00",X"08",X"82",X"00",X"41",X"00",X"80",X"00",X"08",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"7F",X"00",X"00",X"06",X"00",X"00",X"0C",X"C0",X"C0",
		X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"0C",X"00",X"00",X"06",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"65",X"1F",X"0B",X"00",X"00",X"00",X"03",X"00",X"00",X"CC",X"C0",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"18",X"00",X"00",X"18",X"00",X"00",
		X"00",X"00",X"00",X"20",X"1A",X"04",X"0A",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"C3",X"E0",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"80",X"00",X"20",X"10",X"00",X"40",X"20",
		X"00",X"00",X"00",X"10",X"1A",X"04",X"0A",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"01",X"08",X"04",X"20",X"10",X"80",X"40",
		X"00",X"00",X"10",X"08",X"0A",X"04",X"0A",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"03",X"03",X"01",X"00",X"00",X"00",X"02",X"02",X"C0",X"82",X"11",X"08",X"80",X"80",X"00",X"00",
		X"00",X"04",X"04",X"02",X"03",X"06",X"03",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"03",X"03",X"00",X"00",X"02",X"02",X"10",X"10",X"80",X"00",X"00",X"24",X"24",X"00",X"00",X"00",
		X"00",X"01",X"01",X"01",X"01",X"03",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"80",
		X"03",X"03",X"00",X"00",X"04",X"24",X"20",X"00",X"80",X"80",X"00",X"00",X"40",X"48",X"08",X"00",
		X"02",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"06",X"00",X"00",X"0C",X"00",X"00",
		X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"06",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"03",X"00",X"02",X"28",X"00",X"00",
		X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"28",X"02",X"00",X"03",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"84",X"00",X"00",
		X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"84",X"00",X"01",X"00",X"01",X"00",X"00",
		X"00",X"00",X"00",X"02",X"20",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"02",X"00",X"00",X"00",
		X"00",X"00",X"20",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"06",X"00",
		X"00",X"08",X"00",X"40",X"00",X"00",X"00",X"00",X"08",X"00",X"09",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"40",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"08",X"00",
		X"20",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"00",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"22",X"00",X"00",X"00",
		X"00",X"C0",X"00",X"01",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"01",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",
		X"20",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"05",X"1F",X"36",X"39",X"72",X"E0",X"E8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"04",X"02",X"02",X"35",X"10",X"72",X"25",X"2A",X"80",X"58",X"50",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"11",X"4C",X"60",X"01",X"86",
		X"00",X"00",X"18",X"1A",X"10",X"02",X"19",X"0A",X"10",X"42",X"40",X"00",X"10",X"40",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"01",X"80",X"61",X"0C",X"10",X"84",X"80",
		X"00",X"20",X"28",X"20",X"04",X"42",X"10",X"10",X"00",X"00",X"00",X"10",X"00",X"40",X"00",X"00",
		X"00",X"01",X"00",X"00",X"02",X"81",X"00",X"40",X"00",X"0D",X"68",X"10",X"00",X"82",X"00",X"00",
		X"40",X"10",X"00",X"00",X"00",X"A0",X"20",X"00",X"00",X"00",X"00",X"20",X"00",X"80",X"00",X"00",
		X"00",X"08",X"01",X"00",X"00",X"80",X"80",X"20",X"19",X"00",X"80",X"00",X"02",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"80",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"01",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"80",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"00",X"80",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"40",X"00",X"00",X"00",X"00",X"08",
		X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"09",X"30",X"1F",X"63",X"4E",X"D9",X"00",X"90",X"F4",X"E6",X"28",X"CC",X"46",X"B3",
		X"E3",X"7B",X"7C",X"1F",X"25",X"30",X"0F",X"02",X"C6",X"F6",X"DC",X"68",X"9E",X"24",X"80",X"80",
		X"00",X"00",X"04",X"19",X"08",X"3F",X"2F",X"6C",X"00",X"C0",X"E0",X"F4",X"26",X"88",X"8E",X"E7",
		X"E1",X"3D",X"0E",X"23",X"80",X"0F",X"02",X"00",X"EE",X"DC",X"68",X"9C",X"28",X"00",X"00",X"00",
		X"00",X"00",X"00",X"05",X"01",X"00",X"1F",X"3E",X"00",X"00",X"C0",X"E0",X"FC",X"38",X"9C",X"1E",
		X"38",X"1D",X"16",X"10",X"0F",X"02",X"00",X"00",X"D4",X"B8",X"D0",X"18",X"80",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"01",X"0C",X"1E",X"00",X"00",X"00",X"80",X"D0",X"F8",X"10",X"CC",
		X"0C",X"06",X"0C",X"07",X"01",X"00",X"00",X"00",X"B0",X"D0",X"00",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"07",X"04",X"0E",X"00",X"00",X"00",X"40",X"D0",X"B0",X"50",X"E8",
		X"06",X"04",X"01",X"01",X"00",X"00",X"00",X"00",X"A0",X"80",X"00",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"06",X"00",X"00",X"00",X"00",X"40",X"E0",X"60",X"70",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"12",X"06",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",
		X"07",X"0F",X"06",X"12",X"0E",X"00",X"00",X"00",X"F0",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"07",X"09",X"06",X"0F",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",
		X"1F",X"0F",X"25",X"1C",X"00",X"00",X"00",X"00",X"F0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"05",X"00",X"07",X"03",X"0F",X"00",X"00",X"00",X"80",X"80",X"00",X"C0",X"C0",
		X"0F",X"2D",X"1C",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"70",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"02",X"01",X"0B",X"27",X"00",X"00",X"80",X"40",X"40",X"80",X"80",X"C0",
		X"27",X"19",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"60",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"15",X"27",X"00",X"00",X"00",X"40",X"20",X"E0",X"E0",X"80",
		X"17",X"1B",X"03",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"E0",X"E0",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"05",X"0B",X"0B",X"00",X"00",X"00",X"10",X"48",X"68",X"F8",X"C0",
		X"0D",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"E0",X"E0",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"09",X"0B",X"0F",X"01",X"00",X"00",X"00",X"10",X"48",X"E8",X"F8",X"C0",
		X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"E0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"0E",X"12",X"06",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",
		X"07",X"0F",X"06",X"12",X"0E",X"00",X"00",X"00",X"F0",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"0A",X"06",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",
		X"07",X"0F",X"06",X"0A",X"06",X"00",X"00",X"00",X"F0",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"0A",X"06",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"07",X"0F",X"06",X"0A",X"04",X"00",X"00",X"00",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"06",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"07",X"03",X"06",X"02",X"00",X"00",X"00",X"00",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"03",X"03",X"06",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"06",X"02",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"F0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"FE",X"1E",X"06",X"06",X"06",X"06",X"06",X"06",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"F0",X"FF",X"00",X"06",X"06",X"06",X"06",X"06",X"1E",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"08",X"DF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"DF",X"08",X"06",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"37",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"37",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"00",X"00",X"40",X"80",X"FF",
		X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"80",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"7F",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"20",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"DF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DF",X"10",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"2F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2F",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"28",X"54",X"7C",X"00",X"78",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"78",X"00",X"6C",X"50",X"7C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"1E",X"3E",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"3E",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"1C",X"3C",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"3C",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"38",X"78",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"78",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"30",X"70",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"70",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"60",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"60",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
