library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity rom6t31 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of rom6t31 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"10",X"13",X"03",X"01",X"00",X"05",X"05",X"06",X"08",X"14",X"00",X"05",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"04",X"01",X"12",X"09",X"14",X"0E",X"0F",
		X"57",X"21",X"36",X"22",X"21",X"00",X"2E",X"88",X"00",X"1B",X"00",X"1B",X"00",X"1B",X"00",X"00",
		X"32",X"00",X"22",X"5B",X"1C",X"C2",X"C3",X"49",X"13",X"C3",X"21",X"49",X"22",X"57",X"3E",X"34",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"05",X"18",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C2",X"0D",X"4A",X"55",X"18",X"11",X"19",X"00",X"0C",X"21",X"0E",X"2E",X"36",X"08",X"23",X"00",
		X"FF",X"04",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"7C",X"C2",X"37",X"4A",X"53",X"D3",X"C3",
		X"CA",X"81",X"4A",X"83",X"01",X"3E",X"59",X"32",X"03",X"DB",X"7F",X"EE",X"E6",X"F3",X"FE",X"81",
		X"32",X"AF",X"22",X"59",X"00",X"DB",X"80",X"E6",X"AF",X"22",X"3A",X"C9",X"22",X"59",X"C8",X"A7",
		X"22",X"5A",X"CA",X"A7",X"4A",X"A5",X"32",X"AF",X"97",X"CA",X"3E",X"4A",X"A7",X"01",X"3A",X"C9",
		X"22",X"5A",X"C9",X"AF",X"18",X"01",X"1A",X"04",X"22",X"5A",X"93",X"C3",X"3E",X"4A",X"32",X"01",
		X"06",X"C8",X"D5",X"04",X"1C",X"11",X"19",X"00",X"13",X"77",X"05",X"23",X"AF",X"C2",X"0D",X"4A",
		X"4B",X"E0",X"AC",X"CD",X"21",X"4A",X"2A",X"16",X"C3",X"D1",X"4A",X"AF",X"16",X"21",X"11",X"26",
		X"11",X"2E",X"4D",X"00",X"AC",X"CD",X"21",X"4A",X"A0",X"11",X"CD",X"4C",X"4A",X"AC",X"16",X"21",
		X"60",X"11",X"21",X"4D",X"36",X"16",X"AC",X"CD",X"32",X"16",X"40",X"11",X"CD",X"4C",X"4A",X"AC",
		X"4A",X"AC",X"DF",X"DF",X"DF",X"DF",X"C9",X"DF",X"11",X"4A",X"4D",X"C0",X"16",X"21",X"CD",X"3A",
		X"1F",X"00",X"44",X"24",X"1F",X"24",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3E",X"00",X"41",X"41",X"22",X"41",X"00",X"00",X"7F",X"00",X"49",X"49",X"36",X"49",X"00",X"00",
		X"7F",X"00",X"49",X"49",X"41",X"49",X"00",X"00",X"7F",X"00",X"41",X"41",X"3E",X"41",X"00",X"00",
		X"3E",X"00",X"41",X"41",X"47",X"45",X"00",X"00",X"7F",X"00",X"48",X"48",X"40",X"48",X"00",X"00",
		X"00",X"00",X"7F",X"41",X"00",X"41",X"00",X"00",X"7F",X"00",X"08",X"08",X"7F",X"08",X"00",X"00",
		X"7F",X"00",X"14",X"08",X"41",X"22",X"00",X"00",X"02",X"00",X"01",X"01",X"7E",X"01",X"00",X"00",
		X"7F",X"00",X"18",X"20",X"7F",X"20",X"00",X"00",X"7F",X"00",X"01",X"01",X"01",X"01",X"00",X"00",
		X"3E",X"00",X"41",X"41",X"3E",X"41",X"00",X"00",X"7F",X"00",X"08",X"10",X"7F",X"04",X"00",X"00",
		X"3E",X"00",X"45",X"41",X"3D",X"42",X"00",X"00",X"7F",X"00",X"48",X"48",X"30",X"48",X"00",X"00",
		X"32",X"00",X"49",X"49",X"26",X"49",X"00",X"00",X"7F",X"00",X"4C",X"48",X"31",X"4A",X"00",X"00",
		X"7E",X"00",X"01",X"01",X"7E",X"01",X"00",X"00",X"40",X"00",X"7F",X"40",X"40",X"40",X"00",X"00",
		X"7F",X"00",X"0C",X"02",X"7F",X"02",X"00",X"00",X"7C",X"00",X"01",X"02",X"7C",X"02",X"00",X"00",
		X"60",X"00",X"0F",X"10",X"60",X"10",X"00",X"00",X"63",X"00",X"08",X"14",X"63",X"14",X"00",X"00",
		X"08",X"00",X"08",X"08",X"08",X"08",X"00",X"00",X"43",X"00",X"49",X"45",X"61",X"51",X"00",X"00",
		X"00",X"00",X"FF",X"C0",X"00",X"00",X"FF",X"F8",X"00",X"00",X"F8",X"00",X"00",X"00",X"FF",X"00",
		X"FC",X"00",X"00",X"FF",X"FF",X"80",X"00",X"1F",X"00",X"00",X"FF",X"FF",X"F0",X"00",X"07",X"FF",
		X"C2",X"23",X"48",X"03",X"A0",X"3E",X"43",X"32",X"00",X"21",X"36",X"00",X"23",X"00",X"FE",X"7C",
		X"32",X"3D",X"22",X"4C",X"CA",X"A7",X"48",X"22",X"C3",X"22",X"40",X"CD",X"3A",X"F5",X"22",X"4C",
		X"C3",X"33",X"1F",X"9F",X"D5",X"1A",X"11",X"E5",X"C9",X"F1",X"03",X"3E",X"4C",X"32",X"33",X"22",
		X"0D",X"13",X"2C",X"C2",X"C9",X"48",X"FF",X"FF",X"4B",X"00",X"AA",X"CD",X"E1",X"0B",X"24",X"D1",
		X"46",X"1A",X"DA",X"B8",X"48",X"57",X"7E",X"C2",X"AB",X"11",X"21",X"20",X"20",X"A7",X"03",X"0E",
		X"50",X"32",X"11",X"22",X"20",X"A5",X"4D",X"21",X"1B",X"48",X"0D",X"2B",X"48",X"C2",X"AF",X"48",
		X"22",X"4F",X"03",X"0E",X"46",X"1A",X"DA",X"B8",X"06",X"22",X"EF",X"03",X"A3",X"11",X"21",X"20",
		X"6C",X"C2",X"C3",X"48",X"05",X"18",X"20",X"3E",X"48",X"89",X"18",X"C2",X"1B",X"05",X"0D",X"2B",
		X"21",X"48",X"20",X"A1",X"4D",X"11",X"06",X"22",X"50",X"32",X"11",X"22",X"20",X"A9",X"5E",X"C3",
		X"07",X"D3",X"51",X"21",X"3E",X"22",X"77",X"01",X"EF",X"03",X"80",X"C3",X"3A",X"49",X"22",X"50",
		X"49",X"A0",X"0F",X"0E",X"2C",X"CD",X"3A",X"48",X"77",X"23",X"77",X"23",X"99",X"21",X"11",X"29",
		X"11",X"49",X"0B",X"90",X"08",X"0E",X"F1",X"CD",X"22",X"50",X"21",X"A7",X"2D",X"17",X"76",X"C2",
		X"CD",X"11",X"48",X"2C",X"93",X"21",X"11",X"29",X"21",X"09",X"28",X"95",X"B0",X"11",X"0E",X"49",
		X"29",X"91",X"D8",X"11",X"0E",X"49",X"CD",X"0F",X"49",X"C8",X"0F",X"0E",X"2C",X"CD",X"21",X"48",
		X"12",X"0E",X"2C",X"CD",X"21",X"48",X"2F",X"8D",X"48",X"2C",X"0F",X"21",X"11",X"28",X"49",X"E8",
		X"0B",X"21",X"11",X"29",X"4A",X"08",X"10",X"0E",X"00",X"11",X"0E",X"4A",X"CD",X"03",X"48",X"2C",
		X"0E",X"4A",X"CD",X"05",X"48",X"2C",X"03",X"3E",X"2C",X"CD",X"21",X"48",X"2E",X"88",X"20",X"11",
		X"22",X"22",X"22",X"55",X"55",X"2A",X"0E",X"22",X"28",X"C3",X"11",X"4A",X"22",X"51",X"54",X"32",
		X"22",X"50",X"C2",X"A7",X"49",X"4F",X"03",X"DB",X"D5",X"01",X"2C",X"CD",X"DF",X"48",X"3A",X"D1",
		X"C4",X"20",X"49",X"6D",X"03",X"DB",X"10",X"E6",X"40",X"E6",X"64",X"C4",X"DB",X"49",X"E6",X"03",
		X"C2",X"00",X"49",X"16",X"92",X"C3",X"DB",X"49",X"33",X"CA",X"C3",X"4A",X"4E",X"50",X"22",X"54",
		X"20",X"E6",X"6D",X"C4",X"DB",X"49",X"E6",X"00",X"E6",X"00",X"C4",X"40",X"49",X"64",X"00",X"DB",
		X"C0",X"1B",X"12",X"AF",X"1A",X"C9",X"12",X"3D",X"C3",X"10",X"49",X"40",X"3C",X"1A",X"FE",X"12",
		X"C3",X"0B",X"48",X"BC",X"FF",X"FF",X"FF",X"FF",X"F0",X"A7",X"1A",X"3E",X"C9",X"12",X"98",X"11",
		X"48",X"94",X"01",X"3E",X"E2",X"32",X"C3",X"20",X"11",X"CD",X"3A",X"40",X"22",X"50",X"CA",X"A7",
		X"FF",X"05",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"48",X"95",X"32",X"AF",X"20",X"E2",X"18",X"C3",
		X"01",X"0C",X"09",X"14",X"0E",X"0F",X"00",X"13",X"0F",X"03",X"07",X"0E",X"01",X"12",X"15",X"14",
		X"01",X"00",X"08",X"03",X"09",X"05",X"05",X"16",X"0F",X"19",X"00",X"15",X"01",X"08",X"05",X"16",
		X"0F",X"14",X"01",X"04",X"13",X"19",X"08",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"10",X"01",X"05",X"05",X"13",X"12",X"00",X"1B",X"09",X"03",X"13",X"12",X"0F",X"00",X"05",
		X"0F",X"19",X"12",X"15",X"09",X"00",X"09",X"0E",X"07",X"05",X"13",X"09",X"05",X"14",X"00",X"12",
		X"08",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"14",X"0C",X"01",X"00",X"13",X"09",X"17",
		X"07",X"E0",X"07",X"E0",X"03",X"FF",X"FF",X"C0",X"1F",X"80",X"01",X"F8",X"0F",X"C0",X"03",X"F0",
		X"00",X"7F",X"FE",X"00",X"00",X"3F",X"FC",X"00",X"01",X"FF",X"FF",X"80",X"00",X"FF",X"FF",X"00",
		X"06",X"06",X"EE",X"7E",X"77",X"FF",X"05",X"23",X"0F",X"0E",X"15",X"21",X"11",X"25",X"00",X"1A",
		X"19",X"4E",X"28",X"C3",X"0D",X"4E",X"C5",X"F5",X"2A",X"C2",X"7C",X"4E",X"3E",X"FE",X"3D",X"CA",
		X"FF",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"DF",X"C1",X"00",X"C2",X"F1",X"4E",X"22",
		X"3A",X"24",X"22",X"54",X"CA",X"3D",X"49",X"92",X"5B",X"3A",X"A7",X"22",X"1C",X"C2",X"13",X"49",
		X"C3",X"3D",X"49",X"16",X"FF",X"FF",X"FF",X"FF",X"01",X"3E",X"5B",X"32",X"3A",X"22",X"22",X"54",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"FF",X"00",X"00",X"0F",X"FF",X"00",X"00",X"FF",X"F0",X"00",X"03",X"FF",X"FC",X"00",X"00",
		X"FF",X"FC",X"00",X"00",X"FF",X"F0",X"00",X"03",X"0F",X"FF",X"00",X"00",X"3F",X"FF",X"00",X"00",
		X"F0",X"00",X"07",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"80",X"00",X"1F",X"FC",X"00",X"00",X"FF",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"F8",X"00",X"00",X"00",X"FF",X"F8",X"00",X"00",X"FF",X"C0",
		X"00",X"00",X"F8",X"00",X"00",X"00",X"F8",X"00",X"00",X"00",X"F8",X"00",X"00",X"00",X"F8",X"00",
		X"00",X"00",X"F8",X"00",X"00",X"00",X"F8",X"00",X"00",X"00",X"F8",X"00",X"00",X"00",X"F8",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"F8",X"00",X"00",X"00",X"F8",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"F8",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"F8",X"00",X"00",X"00",X"F8",X"00",X"00",X"00",X"F8",X"00",X"00",X"00",X"F8",X"00",
		X"00",X"00",X"F8",X"00",X"00",X"00",X"F8",X"00",X"00",X"00",X"F8",X"00",X"00",X"00",X"F8",X"00",
		X"FF",X"FC",X"3F",X"FF",X"FF",X"FE",X"7F",X"FF",X"FF",X"F0",X"0F",X"FF",X"FF",X"F8",X"1F",X"FF",
		X"00",X"3F",X"FC",X"00",X"00",X"1F",X"F8",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"7F",X"FE",X"00",
		X"00",X"1F",X"F8",X"00",X"00",X"1F",X"F8",X"00",X"00",X"1F",X"F8",X"00",X"00",X"1F",X"F8",X"00",
		X"00",X"1F",X"F8",X"00",X"00",X"1F",X"F8",X"00",X"00",X"1F",X"F8",X"00",X"00",X"1F",X"F8",X"00",
		X"00",X"7F",X"FE",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"1F",X"F8",X"00",X"00",X"3F",X"FC",X"00",
		X"FF",X"F8",X"1F",X"FF",X"FF",X"F0",X"0F",X"FF",X"FF",X"FE",X"7F",X"FF",X"FF",X"FC",X"3F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E0",X"00",X"F8",X"03",X"E0",X"00",X"F8",X"03",X"FF",X"FF",X"FF",X"FF",X"E0",X"00",X"F8",X"03",
		X"FE",X"00",X"F8",X"03",X"FF",X"80",X"F8",X"03",X"F0",X"00",X"F8",X"03",X"FC",X"00",X"F8",X"03",
		X"EF",X"F8",X"F8",X"03",X"E3",X"FC",X"F8",X"03",X"FF",X"C0",X"F8",X"03",X"FF",X"E0",X"F8",X"03",
		X"C0",X"3F",X"7F",X"FF",X"80",X"0F",X"7F",X"FF",X"E1",X"FF",X"FC",X"07",X"C0",X"FF",X"FE",X"0F",
		X"00",X"01",X"07",X"F8",X"00",X"00",X"00",X"00",X"00",X"07",X"3F",X"FF",X"00",X"03",X"1F",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E0",X"1F",X"F8",X"03",X"E0",X"1F",X"F8",X"03",X"FF",X"FF",X"FF",X"FF",X"E0",X"1F",X"F8",X"03",
		X"E0",X"1F",X"F8",X"03",X"E0",X"1F",X"F8",X"03",X"E0",X"1F",X"F8",X"03",X"E0",X"1F",X"F8",X"03",
		X"E0",X"1F",X"F8",X"03",X"E0",X"1F",X"F8",X"03",X"E0",X"1F",X"F8",X"03",X"E0",X"1F",X"F8",X"03",
		X"E0",X"1F",X"F8",X"03",X"00",X"1F",X"F8",X"00",X"E0",X"1F",X"F8",X"03",X"E0",X"1F",X"F8",X"03",
		X"00",X"1F",X"F8",X"00",X"00",X"1F",X"F8",X"00",X"00",X"1F",X"F8",X"00",X"00",X"1F",X"F8",X"00",
		X"00",X"FF",X"FF",X"00",X"01",X"FF",X"FF",X"80",X"00",X"3F",X"FC",X"00",X"00",X"7F",X"FE",X"00",
		X"0F",X"C0",X"03",X"F0",X"1F",X"80",X"01",X"F8",X"03",X"FF",X"FF",X"C0",X"07",X"E0",X"07",X"E0",
		X"FC",X"00",X"00",X"3F",X"F8",X"00",X"00",X"1F",X"3F",X"00",X"00",X"FC",X"FE",X"00",X"00",X"7F",
		X"FE",X"00",X"00",X"7F",X"3F",X"00",X"00",X"FC",X"F8",X"00",X"00",X"1F",X"FC",X"00",X"00",X"3F");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
