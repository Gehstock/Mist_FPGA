library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity PROG is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of PROG is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"4C",X"4B",X"3B",X"1B",X"31",X"39",X"38",X"30",X"20",X"41",X"54",X"41",X"52",X"C9",X"20",X"76",
		X"28",X"58",X"20",X"60",X"2D",X"46",X"8A",X"90",X"FC",X"8D",X"00",X"20",X"AD",X"00",X"0C",X"29",
		X"20",X"F0",X"FE",X"20",X"66",X"25",X"20",X"79",X"30",X"20",X"45",X"27",X"10",X"E7",X"20",X"07",
		X"3B",X"20",X"19",X"21",X"20",X"27",X"33",X"20",X"55",X"29",X"20",X"01",X"27",X"20",X"D2",X"2A",
		X"20",X"02",X"22",X"20",X"D7",X"2E",X"20",X"DD",X"2B",X"20",X"1C",X"2E",X"20",X"59",X"20",X"20",
		X"DA",X"23",X"20",X"F3",X"2C",X"4C",X"15",X"20",X"55",X"A5",X"43",X"29",X"AF",X"D0",X"08",X"A5",
		X"40",X"45",X"EF",X"C9",X"20",X"90",X"01",X"60",X"A5",X"70",X"45",X"F0",X"C9",X"F8",X"90",X"20",
		X"A6",X"88",X"B5",X"9A",X"C9",X"0C",X"B0",X"6B",X"B5",X"AB",X"C9",X"02",X"A0",X"05",X"90",X"02",
		X"A0",X"09",X"C9",X"12",X"90",X"05",X"4A",X"18",X"69",X"06",X"A8",X"98",X"D5",X"D7",X"90",X"53",
		X"A5",X"00",X"29",X"03",X"D0",X"0F",X"E6",X"40",X"A5",X"40",X"18",X"69",X"01",X"29",X"03",X"09",
		X"1C",X"45",X"EF",X"85",X"40",X"A5",X"60",X"85",X"8B",X"A5",X"70",X"A4",X"EF",X"F0",X"06",X"18",
		X"65",X"80",X"4C",X"B8",X"20",X"38",X"E5",X"80",X"85",X"70",X"45",X"F0",X"C9",X"04",X"90",X"24",
		X"A2",X"0C",X"20",X"9A",X"2C",X"90",X"1C",X"A5",X"00",X"29",X"03",X"D0",X"16",X"AD",X"0A",X"10",
		X"29",X"03",X"D0",X"0F",X"A9",X"04",X"45",X"F3",X"18",X"65",X"70",X"A0",X"00",X"20",X"2F",X"2C",
		X"20",X"AC",X"2B",X"60",X"20",X"E8",X"20",X"60",X"A9",X"1C",X"45",X"EF",X"85",X"40",X"A9",X"F8",
		X"45",X"F0",X"85",X"70",X"AD",X"0A",X"10",X"29",X"F8",X"F0",X"F9",X"C9",X"10",X"90",X"F5",X"38",
		X"E9",X"04",X"85",X"60",X"A0",X"03",X"A6",X"88",X"B5",X"AB",X"C9",X"06",X"B0",X"02",X"A0",X"02",
		X"84",X"80",X"A9",X"00",X"85",X"50",X"85",X"B8",X"60",X"A5",X"86",X"10",X"6F",X"20",X"95",X"21",
		X"A9",X"03",X"85",X"93",X"A9",X"20",X"85",X"94",X"A9",X"40",X"85",X"91",X"A9",X"05",X"85",X"92",
		X"20",X"74",X"38",X"A5",X"00",X"D0",X"05",X"A9",X"84",X"20",X"24",X"38",X"A5",X"00",X"AE",X"00",
		X"06",X"86",X"FF",X"29",X"80",X"D0",X"45",X"A5",X"43",X"29",X"AF",X"D0",X"30",X"A5",X"63",X"A0",
		X"01",X"C9",X"1C",X"90",X"08",X"A0",X"FF",X"C9",X"E4",X"B0",X"02",X"A4",X"53",X"98",X"84",X"53",
		X"18",X"20",X"EF",X"2A",X"A5",X"73",X"85",X"8D",X"A0",X"FF",X"C9",X"30",X"B0",X"08",X"A0",X"01",
		X"C9",X"09",X"90",X"02",X"A4",X"83",X"98",X"84",X"83",X"18",X"20",X"28",X"2B",X"20",X"64",X"2B",
		X"A2",X"13",X"A9",X"AB",X"5D",X"20",X"21",X"CA",X"10",X"FA",X"85",X"FE",X"60",X"02",X"BB",X"5A",
		X"30",X"5F",X"EE",X"7D",X"A8",X"20",X"B3",X"21",X"85",X"AE",X"B9",X"C0",X"21",X"85",X"B0",X"A9",
		X"06",X"20",X"24",X"38",X"A5",X"B0",X"20",X"AB",X"38",X"A5",X"AE",X"20",X"9E",X"38",X"A9",X"00",
		X"4C",X"9E",X"38",X"A5",X"FD",X"29",X"30",X"4A",X"4A",X"4A",X"A8",X"B9",X"BF",X"21",X"60",X"00",
		X"01",X"20",X"01",X"50",X"01",X"00",X"02",X"A6",X"88",X"A0",X"02",X"B5",X"AB",X"D0",X"0C",X"A5",
		X"FD",X"29",X"40",X"09",X"10",X"D5",X"A9",X"90",X"02",X"A0",X"01",X"84",X"81",X"AD",X"0A",X"10",
		X"29",X"04",X"F0",X"05",X"98",X"20",X"7C",X"38",X"A8",X"84",X"51",X"A9",X"60",X"45",X"F0",X"85",
		X"71",X"A9",X"FF",X"85",X"61",X"A9",X"F8",X"85",X"41",X"A9",X"60",X"85",X"A1",X"A9",X"00",X"85",
		X"B5",X"60",X"A5",X"43",X"29",X"AF",X"F0",X"01",X"60",X"A2",X"0D",X"A5",X"41",X"A8",X"29",X"20",
		X"F0",X"07",X"C0",X"F8",X"90",X"F2",X"4C",X"FA",X"22",X"A5",X"00",X"29",X"03",X"D0",X"10",X"E6",
		X"41",X"A5",X"41",X"45",X"F2",X"C9",X"1C",X"90",X"06",X"A9",X"14",X"45",X"F2",X"85",X"41",X"C6",
		X"A1",X"D0",X"35",X"AD",X"0A",X"10",X"29",X"80",X"F0",X"18",X"A5",X"51",X"F0",X"10",X"A4",X"61",
		X"C0",X"FB",X"B0",X"0E",X"C0",X"05",X"90",X"0A",X"85",X"BE",X"A9",X"00",X"F0",X"02",X"A5",X"BE",
		X"85",X"51",X"A5",X"FD",X"29",X"40",X"09",X"20",X"2D",X"0A",X"10",X"F0",X"07",X"A5",X"81",X"20",
		X"7C",X"38",X"85",X"81",X"A9",X"30",X"85",X"A1",X"A5",X"61",X"38",X"E5",X"51",X"85",X"61",X"85",
		X"8B",X"A5",X"71",X"A4",X"EF",X"F0",X"06",X"18",X"65",X"81",X"4C",X"80",X"22",X"38",X"E5",X"81",
		X"85",X"71",X"A0",X"00",X"20",X"2F",X"2C",X"F0",X"13",X"A0",X"00",X"B1",X"32",X"29",X"3F",X"C9",
		X"38",X"90",X"09",X"A9",X"00",X"91",X"32",X"20",X"95",X"2B",X"A2",X"0D",X"A5",X"61",X"C9",X"FF",
		X"B0",X"54",X"A5",X"71",X"45",X"F0",X"C9",X"09",X"B0",X"06",X"A5",X"81",X"10",X"3D",X"30",X"32",
		X"A6",X"88",X"B5",X"AB",X"F8",X"38",X"E9",X"06",X"D8",X"10",X"02",X"A9",X"00",X"4A",X"C9",X"06",
		X"90",X"02",X"A9",X"05",X"0A",X"0A",X"0A",X"85",X"8D",X"A9",X"60",X"45",X"F0",X"38",X"E5",X"8D",
		X"A6",X"EF",X"F0",X"06",X"C5",X"71",X"90",X"0A",X"B0",X"04",X"C5",X"71",X"B0",X"04",X"A5",X"81",
		X"30",X"09",X"A2",X"0D",X"20",X"6F",X"2C",X"90",X"07",X"A5",X"81",X"20",X"7C",X"38",X"85",X"81",
		X"A2",X"0D",X"20",X"9A",X"2C",X"60",X"20",X"C7",X"21",X"60",X"C6",X"A1",X"D0",X"11",X"AD",X"0A",
		X"10",X"29",X"2F",X"09",X"0F",X"85",X"A1",X"A9",X"14",X"85",X"B5",X"45",X"F2",X"85",X"41",X"60",
		X"B5",X"54",X"85",X"8B",X"A0",X"FF",X"B5",X"44",X"30",X"02",X"A0",X"01",X"B5",X"64",X"60",X"A6",
		X"88",X"B5",X"94",X"D0",X"20",X"B5",X"C2",X"09",X"80",X"95",X"C2",X"B5",X"9C",X"C9",X"03",X"90",
		X"14",X"D6",X"9A",X"D0",X"04",X"A9",X"0C",X"95",X"9A",X"A9",X"02",X"B4",X"AB",X"C0",X"04",X"B0",
		X"02",X"A9",X"01",X"95",X"9C",X"A9",X"03",X"85",X"34",X"B5",X"9C",X"85",X"74",X"A8",X"A5",X"00",
		X"29",X"02",X"D0",X"05",X"98",X"20",X"7C",X"38",X"A8",X"84",X"44",X"A9",X"F8",X"45",X"F0",X"85",
		X"64",X"A9",X"80",X"85",X"54",X"B5",X"9A",X"85",X"8B",X"C9",X"01",X"F0",X"35",X"A0",X"42",X"A2",
		X"01",X"94",X"34",X"A9",X"F8",X"45",X"F0",X"95",X"64",X"B5",X"73",X"95",X"74",X"B5",X"43",X"95",
		X"44",X"10",X"04",X"A9",X"08",X"D0",X"02",X"A9",X"F8",X"18",X"75",X"53",X"95",X"54",X"88",X"C0",
		X"3F",X"D0",X"02",X"A0",X"47",X"E8",X"E4",X"8B",X"90",X"D7",X"A6",X"88",X"B5",X"9A",X"C9",X"0C",
		X"F0",X"2D",X"A9",X"F8",X"45",X"F0",X"A6",X"8B",X"95",X"64",X"A9",X"00",X"95",X"34",X"A9",X"02",
		X"A4",X"F4",X"F0",X"01",X"98",X"95",X"74",X"2C",X"0A",X"10",X"10",X"03",X"20",X"7C",X"38",X"95",
		X"44",X"AD",X"0A",X"10",X"29",X"F8",X"95",X"54",X"B5",X"64",X"E8",X"E0",X"0C",X"90",X"D9",X"A9",
		X"0C",X"A6",X"88",X"95",X"94",X"A5",X"FE",X"85",X"97",X"60",X"A5",X"86",X"30",X"38",X"AD",X"01",
		X"08",X"29",X"1C",X"F0",X"31",X"A5",X"AB",X"05",X"AD",X"F0",X"1B",X"C6",X"A9",X"D0",X"27",X"A9",
		X"3C",X"85",X"A9",X"F8",X"A5",X"AB",X"38",X"E9",X"01",X"D8",X"85",X"AB",X"10",X"18",X"C6",X"AD",
		X"A9",X"59",X"85",X"AB",X"D0",X"10",X"A9",X"00",X"85",X"A5",X"20",X"BC",X"26",X"A5",X"43",X"29",
		X"AF",X"D0",X"03",X"20",X"C8",X"2C",X"A5",X"87",X"D0",X"01",X"60",X"A5",X"DB",X"D0",X"FB",X"C6",
		X"87",X"D0",X"F7",X"A5",X"D6",X"F0",X"0F",X"A9",X"80",X"20",X"24",X"38",X"A9",X"00",X"A8",X"91",
		X"91",X"85",X"D6",X"4C",X"36",X"29",X"A5",X"43",X"29",X"AF",X"D0",X"03",X"4C",X"41",X"25",X"20",
		X"36",X"29",X"A5",X"86",X"10",X"11",X"A5",X"01",X"10",X"0A",X"29",X"7F",X"85",X"01",X"20",X"FE",
		X"31",X"20",X"60",X"2D",X"4C",X"3B",X"25",X"A5",X"A5",X"05",X"A6",X"D0",X"46",X"C6",X"86",X"20",
		X"67",X"32",X"A5",X"EF",X"F0",X"18",X"A5",X"C2",X"10",X"14",X"A9",X"80",X"85",X"EE",X"20",X"45",
		X"25",X"20",X"36",X"29",X"20",X"FE",X"31",X"A5",X"C1",X"10",X"03",X"20",X"60",X"2D",X"20",X"C7",
		X"21",X"20",X"1F",X"23",X"20",X"E8",X"20",X"A9",X"01",X"85",X"00",X"A9",X"04",X"20",X"24",X"38",
		X"A6",X"89",X"A9",X"FF",X"9D",X"02",X"1C",X"20",X"4F",X"3A",X"A9",X"3D",X"85",X"F9",X"A9",X"00",
		X"85",X"FA",X"60",X"A6",X"89",X"CA",X"D0",X"03",X"4C",X"34",X"25",X"A6",X"88",X"B5",X"A4",X"D0",
		X"24",X"A5",X"A7",X"D0",X"1E",X"E6",X"A7",X"A9",X"80",X"85",X"87",X"A9",X"F9",X"85",X"43",X"85",
		X"42",X"A9",X"04",X"20",X"24",X"38",X"A9",X"00",X"20",X"24",X"38",X"A5",X"88",X"09",X"20",X"20",
		X"85",X"38",X"60",X"C6",X"A7",X"A5",X"88",X"49",X"03",X"AA",X"B5",X"A4",X"F0",X"56",X"86",X"88",
		X"A9",X"80",X"25",X"EE",X"05",X"88",X"85",X"EE",X"C9",X"82",X"D0",X"03",X"20",X"65",X"25",X"B5",
		X"A1",X"85",X"A0",X"A6",X"88",X"E0",X"01",X"D0",X"03",X"20",X"45",X"25",X"20",X"FE",X"31",X"A6",
		X"88",X"E0",X"02",X"D0",X"11",X"B5",X"A4",X"C5",X"A4",X"D0",X"0B",X"A5",X"AD",X"D0",X"07",X"A9",
		X"0C",X"95",X"94",X"20",X"C3",X"28",X"B5",X"C2",X"09",X"40",X"95",X"C2",X"A9",X"A0",X"85",X"87",
		X"A9",X"00",X"20",X"24",X"38",X"A5",X"88",X"09",X"20",X"20",X"85",X"38",X"A9",X"F9",X"85",X"43",
		X"85",X"42",X"85",X"D6",X"A6",X"88",X"D6",X"A4",X"20",X"BC",X"26",X"20",X"C7",X"21",X"20",X"E8",
		X"20",X"20",X"1F",X"23",X"60",X"A5",X"FE",X"85",X"BD",X"85",X"BF",X"8D",X"07",X"1C",X"8D",X"00",
		X"24",X"85",X"F5",X"85",X"F7",X"85",X"F6",X"85",X"F0",X"85",X"EF",X"85",X"F1",X"85",X"F2",X"85",
		X"F3",X"85",X"F4",X"85",X"F8",X"60",X"AD",X"01",X"08",X"29",X"E3",X"85",X"D3",X"29",X"03",X"85",
		X"8D",X"D0",X"04",X"A9",X"02",X"85",X"C8",X"A5",X"FD",X"29",X"0C",X"4A",X"4A",X"69",X"02",X"85",
		X"A4",X"A5",X"86",X"30",X"01",X"60",X"A5",X"8D",X"F0",X"03",X"20",X"24",X"38",X"A5",X"00",X"29",
		X"20",X"0A",X"0A",X"85",X"8D",X"A5",X"C8",X"05",X"C9",X"F0",X"10",X"A6",X"DC",X"10",X"29",X"C9",
		X"02",X"90",X"1E",X"A9",X"00",X"85",X"DC",X"A9",X"8A",X"D0",X"1A",X"A5",X"FD",X"29",X"80",X"85",
		X"DC",X"49",X"8A",X"20",X"24",X"38",X"A2",X"FF",X"8E",X"03",X"1C",X"A2",X"FF",X"8E",X"04",X"1C",
		X"60",X"A9",X"0A",X"05",X"8D",X"20",X"24",X"38",X"A9",X"09",X"20",X"24",X"38",X"A5",X"C8",X"C9",
		X"0A",X"90",X"0A",X"A9",X"21",X"20",X"85",X"38",X"A5",X"C8",X"38",X"E9",X"0A",X"09",X"20",X"20",
		X"85",X"38",X"A5",X"C9",X"F0",X"02",X"A9",X"1E",X"20",X"85",X"38",X"A6",X"C8",X"F0",X"CC",X"A5",
		X"DC",X"30",X"C8",X"A5",X"8D",X"8D",X"03",X"1C",X"AD",X"01",X"0C",X"A6",X"FF",X"4A",X"B0",X"BB",
		X"C6",X"C8",X"A9",X"FF",X"8D",X"03",X"1C",X"8D",X"04",X"1C",X"A9",X"00",X"85",X"FB",X"85",X"FC",
		X"85",X"9A",X"85",X"CB",X"85",X"CA",X"86",X"89",X"9D",X"02",X"1C",X"A6",X"A4",X"CA",X"86",X"A5",
		X"E6",X"86",X"20",X"A4",X"26",X"20",X"B3",X"21",X"85",X"AE",X"85",X"AF",X"B9",X"C0",X"21",X"85",
		X"B0",X"85",X"B1",X"AD",X"00",X"0C",X"29",X"10",X"F0",X"07",X"A9",X"80",X"85",X"EE",X"20",X"45",
		X"25",X"20",X"76",X"28",X"AD",X"01",X"08",X"29",X"1C",X"F0",X"0C",X"4A",X"4A",X"85",X"AD",X"A9",
		X"00",X"85",X"AB",X"A9",X"3C",X"85",X"A9",X"4C",X"BC",X"26",X"BD",X"7A",X"26",X"48",X"BD",X"7B",
		X"26",X"A8",X"BD",X"7C",X"26",X"AA",X"68",X"8E",X"0E",X"14",X"8E",X"06",X"14",X"8D",X"0F",X"14",
		X"8D",X"05",X"14",X"8C",X"0D",X"14",X"8C",X"07",X"14",X"60",X"0D",X"00",X"0E",X"02",X"04",X"01",
		X"0E",X"01",X"0C",X"04",X"01",X"0B",X"01",X"0C",X"0A",X"09",X"0B",X"04",X"0C",X"0D",X"0A",X"09",
		X"0C",X"0E",X"0A",X"0E",X"01",X"0B",X"01",X"04",X"01",X"00",X"06",X"0D",X"0E",X"0A",X"0E",X"0C",
		X"0B",X"00",X"0D",X"02",X"A9",X"FF",X"85",X"C1",X"85",X"C2",X"A2",X"08",X"B5",X"02",X"9D",X"78",
		X"01",X"B5",X"1A",X"9D",X"81",X"01",X"CA",X"10",X"F3",X"4C",X"4F",X"3A",X"A9",X"06",X"85",X"8B",
		X"A9",X"04",X"45",X"F7",X"29",X"06",X"85",X"92",X"A9",X"DF",X"45",X"F6",X"85",X"91",X"A6",X"A5",
		X"A9",X"1F",X"CA",X"10",X"02",X"A9",X"00",X"20",X"85",X"38",X"C6",X"8B",X"D0",X"F2",X"A9",X"06",
		X"45",X"F7",X"85",X"92",X"A9",X"5F",X"45",X"F6",X"85",X"91",X"A9",X"06",X"85",X"8B",X"38",X"E5",
		X"A6",X"AA",X"A9",X"00",X"CA",X"10",X"02",X"A9",X"1F",X"20",X"85",X"38",X"C6",X"8B",X"D0",X"F2",
		X"60",X"A2",X"0D",X"B4",X"34",X"C0",X"F9",X"90",X"18",X"C0",X"FA",X"90",X"04",X"D6",X"34",X"D0",
		X"10",X"E0",X"0D",X"D0",X"0C",X"A5",X"43",X"29",X"AF",X"D0",X"06",X"A5",X"D7",X"45",X"EF",X"85",
		X"41",X"CA",X"10",X"DF",X"A5",X"43",X"29",X"AF",X"F0",X"1A",X"A5",X"00",X"29",X"03",X"D0",X"14",
		X"A5",X"43",X"C9",X"28",X"B0",X"0E",X"E6",X"43",X"C9",X"27",X"D0",X"08",X"A9",X"00",X"85",X"DA",
		X"A9",X"04",X"85",X"DB",X"60",X"A5",X"C1",X"25",X"C2",X"10",X"01",X"60",X"A5",X"C2",X"30",X"18",
		X"A5",X"EE",X"10",X"14",X"A5",X"EF",X"D0",X"10",X"A9",X"82",X"85",X"EE",X"20",X"65",X"25",X"20",
		X"FE",X"31",X"20",X"27",X"33",X"20",X"36",X"29",X"A5",X"89",X"4A",X"F0",X"14",X"A9",X"00",X"20",
		X"24",X"38",X"A0",X"02",X"A6",X"C2",X"10",X"01",X"88",X"84",X"88",X"98",X"09",X"20",X"20",X"85",
		X"38",X"A9",X"08",X"20",X"24",X"38",X"A9",X"05",X"20",X"24",X"38",X"A9",X"89",X"45",X"F5",X"85",
		X"91",X"A9",X"05",X"45",X"F7",X"85",X"92",X"A6",X"88",X"B4",X"C0",X"84",X"8D",X"98",X"18",X"65",
		X"C0",X"85",X"8E",X"20",X"82",X"38",X"A4",X"8D",X"C8",X"20",X"82",X"38",X"A4",X"8D",X"C8",X"C8",
		X"20",X"82",X"38",X"AD",X"01",X"0C",X"A6",X"EF",X"F0",X"01",X"4A",X"4A",X"4A",X"4A",X"26",X"9A",
		X"A5",X"9A",X"29",X"1F",X"C9",X"18",X"D0",X"46",X"E6",X"C0",X"A5",X"C0",X"C9",X"03",X"90",X"32",
		X"A6",X"88",X"A9",X"FF",X"95",X"C0",X"A5",X"EF",X"F0",X"1D",X"A9",X"80",X"85",X"EE",X"20",X"45",
		X"25",X"20",X"FE",X"31",X"20",X"36",X"29",X"20",X"27",X"33",X"20",X"1F",X"23",X"20",X"C7",X"21",
		X"20",X"E8",X"20",X"A5",X"C1",X"30",X"32",X"A5",X"C1",X"25",X"C2",X"30",X"17",X"A2",X"00",X"86",
		X"C0",X"60",X"E6",X"8E",X"A6",X"8E",X"A9",X"F4",X"85",X"01",X"A9",X"01",X"95",X"1A",X"A5",X"01",
		X"F0",X"BE",X"D0",X"2E",X"A9",X"88",X"20",X"24",X"38",X"A9",X"85",X"20",X"24",X"38",X"A9",X"00",
		X"8D",X"89",X"05",X"8D",X"A9",X"05",X"8D",X"C9",X"05",X"20",X"A4",X"26",X"20",X"60",X"2D",X"A6",
		X"89",X"86",X"01",X"CA",X"F0",X"C7",X"A9",X"80",X"20",X"24",X"38",X"A9",X"00",X"A8",X"91",X"91",
		X"F0",X"BB",X"A5",X"00",X"29",X"07",X"D0",X"2B",X"A2",X"FF",X"A9",X"00",X"A4",X"B9",X"85",X"B9",
		X"10",X"07",X"A2",X"01",X"98",X"20",X"7C",X"38",X"A8",X"C0",X"04",X"90",X"16",X"8A",X"45",X"F4",
		X"A6",X"8E",X"18",X"75",X"1A",X"30",X"08",X"C9",X"1B",X"90",X"06",X"A9",X"00",X"F0",X"02",X"A9",
		X"1A",X"95",X"1A",X"A9",X"00",X"60",X"A9",X"20",X"8D",X"08",X"10",X"A9",X"0C",X"85",X"9B",X"85",
		X"9C",X"A5",X"FF",X"85",X"88",X"85",X"53",X"85",X"83",X"A9",X"02",X"85",X"9D",X"85",X"9E",X"A2",
		X"06",X"A9",X"00",X"8D",X"0F",X"10",X"95",X"B2",X"CA",X"10",X"FB",X"A2",X"05",X"95",X"A8",X"CA",
		X"10",X"FB",X"AD",X"0A",X"10",X"4D",X"0A",X"10",X"18",X"65",X"C8",X"85",X"C8",X"A9",X"03",X"8D",
		X"0F",X"10",X"20",X"1F",X"23",X"A9",X"C0",X"85",X"A0",X"85",X"A2",X"85",X"A3",X"20",X"C7",X"21",
		X"20",X"E8",X"20",X"A9",X"0F",X"8D",X"04",X"14",X"A6",X"88",X"A9",X"00",X"95",X"C2",X"AA",X"20",
		X"5A",X"26",X"A2",X"00",X"8A",X"9D",X"00",X"04",X"9D",X"00",X"05",X"9D",X"00",X"06",X"9D",X"00",
		X"07",X"E8",X"D0",X"F1",X"A6",X"88",X"95",X"D7",X"A2",X"1B",X"86",X"8B",X"A2",X"2D",X"AD",X"0A",
		X"10",X"29",X"E0",X"05",X"8B",X"85",X"8D",X"AD",X"0A",X"10",X"29",X"03",X"09",X"04",X"85",X"8E",
		X"86",X"8F",X"A0",X"00",X"A5",X"8D",X"29",X"1F",X"A6",X"EF",X"F0",X"06",X"C9",X"14",X"90",X"0E",
		X"B0",X"04",X"C9",X"0C",X"B0",X"08",X"B1",X"8D",X"D0",X"04",X"A6",X"88",X"F6",X"D7",X"A9",X"3F",
		X"45",X"EF",X"91",X"8D",X"A5",X"8B",X"38",X"E9",X"01",X"C9",X"02",X"B0",X"02",X"A9",X"1B",X"85",
		X"8B",X"A6",X"8F",X"CA",X"10",X"B8",X"A9",X"10",X"45",X"F2",X"85",X"43",X"A9",X"80",X"85",X"63",
		X"85",X"62",X"A9",X"08",X"45",X"F0",X"85",X"73",X"A9",X"0C",X"45",X"F1",X"85",X"72",X"A9",X"11",
		X"45",X"F2",X"85",X"42",X"60",X"A5",X"87",X"F0",X"01",X"60",X"A2",X"0B",X"A5",X"00",X"29",X"0F",
		X"D0",X"04",X"A9",X"07",X"85",X"B3",X"B5",X"34",X"10",X"03",X"4C",X"CB",X"2A",X"A5",X"00",X"29",
		X"01",X"D0",X"09",X"B5",X"34",X"18",X"69",X"01",X"29",X"F7",X"95",X"34",X"A0",X"01",X"B5",X"64",
		X"45",X"F0",X"C9",X"09",X"B0",X"0A",X"B5",X"34",X"C9",X"10",X"B0",X"02",X"84",X"97",X"B5",X"64",
		X"29",X"07",X"D0",X"73",X"98",X"A4",X"88",X"D9",X"94",X"00",X"D0",X"14",X"A9",X"02",X"B4",X"44",
		X"10",X"02",X"A9",X"FE",X"95",X"44",X"A9",X"02",X"B4",X"74",X"10",X"02",X"A9",X"FE",X"95",X"74",
		X"B5",X"34",X"29",X"40",X"F0",X"0F",X"B5",X"63",X"38",X"F5",X"64",X"20",X"7A",X"38",X"C9",X"08",
		X"B0",X"45",X"4C",X"96",X"2A",X"B5",X"34",X"29",X"20",X"D0",X"3C",X"B5",X"54",X"C9",X"F0",X"90",
		X"0A",X"B4",X"74",X"F0",X"0E",X"B4",X"44",X"10",X"2E",X"30",X"0F",X"C9",X"10",X"B0",X"0B",X"B4",
		X"74",X"D0",X"03",X"4C",X"AA",X"2A",X"B4",X"44",X"30",X"1D",X"20",X"10",X"23",X"20",X"2F",X"2C",
		X"F0",X"10",X"C9",X"38",X"90",X"11",X"C9",X"3C",X"B0",X"0D",X"B5",X"34",X"09",X"20",X"95",X"34",
		X"90",X"05",X"20",X"6F",X"2C",X"90",X"BB",X"B5",X"64",X"45",X"F0",X"B4",X"74",X"F0",X"D4",X"10",
		X"12",X"A4",X"EF",X"F0",X"08",X"45",X"F0",X"C9",X"C9",X"90",X"63",X"B0",X"68",X"C9",X"30",X"B0",
		X"5D",X"90",X"62",X"C9",X"09",X"B0",X"5E",X"B5",X"34",X"29",X"40",X"D0",X"51",X"B5",X"34",X"29",
		X"DF",X"95",X"34",X"E0",X"0B",X"F0",X"47",X"8A",X"A8",X"C8",X"B9",X"34",X"00",X"30",X"3F",X"29",
		X"40",X"F0",X"3B",X"C0",X"0B",X"F0",X"09",X"B9",X"35",X"00",X"30",X"04",X"29",X"40",X"D0",X"29",
		X"B9",X"64",X"00",X"45",X"F0",X"C9",X"09",X"B0",X"25",X"B9",X"34",X"00",X"29",X"07",X"99",X"34",
		X"00",X"B9",X"44",X"00",X"20",X"7C",X"38",X"99",X"44",X"00",X"B9",X"64",X"00",X"29",X"F8",X"99",
		X"64",X"00",X"A9",X"00",X"99",X"74",X"00",X"F0",X"05",X"C8",X"C0",X"0C",X"90",X"C5",X"B5",X"74",
		X"20",X"7C",X"38",X"95",X"74",X"B5",X"64",X"A4",X"EF",X"F0",X"06",X"18",X"75",X"74",X"4C",X"94",
		X"2A",X"38",X"F5",X"74",X"95",X"64",X"B5",X"44",X"18",X"75",X"54",X"95",X"54",X"20",X"9A",X"2C",
		X"90",X"2F",X"B5",X"64",X"29",X"07",X"C9",X"04",X"D0",X"21",X"B5",X"44",X"20",X"7C",X"38",X"95",
		X"44",X"B4",X"74",X"D0",X"16",X"09",X"00",X"30",X"03",X"20",X"7C",X"38",X"95",X"74",X"A9",X"04",
		X"B4",X"44",X"10",X"02",X"A9",X"FC",X"18",X"75",X"54",X"95",X"54",X"CA",X"30",X"03",X"4C",X"66",
		X"29",X"60",X"A5",X"86",X"10",X"01",X"60",X"A5",X"43",X"29",X"AF",X"D0",X"F9",X"A5",X"73",X"85",
		X"8D",X"A4",X"FE",X"A5",X"B9",X"84",X"B9",X"20",X"4F",X"32",X"65",X"84",X"85",X"84",X"98",X"65",
		X"63",X"AA",X"85",X"8B",X"A0",X"00",X"A5",X"73",X"20",X"2F",X"2C",X"D0",X"11",X"8A",X"C9",X"F4",
		X"90",X"04",X"A9",X"F4",X"D0",X"0A",X"C9",X"0B",X"B0",X"06",X"A9",X"0B",X"D0",X"02",X"A5",X"63",
		X"85",X"63",X"A4",X"86",X"10",X"01",X"60",X"A0",X"00",X"A5",X"BB",X"84",X"BB",X"20",X"7C",X"38",
		X"20",X"4F",X"32",X"65",X"85",X"85",X"85",X"98",X"65",X"73",X"AA",X"A4",X"63",X"84",X"8B",X"A0",
		X"00",X"20",X"2F",X"2C",X"D0",X"25",X"8A",X"C9",X"08",X"90",X"1C",X"C9",X"F1",X"B0",X"14",X"C9",
		X"80",X"90",X"08",X"C9",X"C8",X"B0",X"16",X"A9",X"C8",X"D0",X"12",X"C9",X"31",X"90",X"0E",X"A9",
		X"30",X"D0",X"0A",X"A9",X"F0",X"D0",X"06",X"A9",X"08",X"D0",X"02",X"A5",X"73",X"85",X"73",X"A4",
		X"86",X"10",X"01",X"60",X"A5",X"72",X"A6",X"EF",X"F0",X"07",X"38",X"E5",X"8D",X"B0",X"0E",X"90",
		X"05",X"38",X"E5",X"8D",X"90",X"07",X"20",X"7A",X"38",X"C9",X"05",X"B0",X"0D",X"A9",X"04",X"45",
		X"F0",X"18",X"65",X"73",X"85",X"72",X"A5",X"63",X"85",X"62",X"A5",X"43",X"29",X"AF",X"F0",X"04",
		X"A9",X"28",X"85",X"42",X"60",X"A5",X"32",X"29",X"1F",X"A6",X"EF",X"F0",X"06",X"C9",X"14",X"90",
		X"0A",X"B0",X"04",X"C9",X"0C",X"B0",X"04",X"A6",X"88",X"D6",X"D7",X"60",X"A0",X"00",X"B1",X"32",
		X"D0",X"2A",X"A5",X"32",X"29",X"1F",X"F0",X"24",X"C9",X"1F",X"F0",X"20",X"A6",X"EF",X"F0",X"0A",
		X"C9",X"1E",X"F0",X"18",X"C9",X"14",X"90",X"0E",X"B0",X"08",X"C9",X"01",X"F0",X"0E",X"C9",X"0C",
		X"B0",X"04",X"A6",X"88",X"F6",X"D7",X"A9",X"3F",X"45",X"EF",X"91",X"32",X"60",X"A5",X"97",X"F0",
		X"4D",X"A5",X"87",X"D0",X"49",X"A5",X"A0",X"F0",X"03",X"C6",X"A0",X"60",X"A6",X"88",X"A0",X"0B",
		X"B9",X"34",X"00",X"30",X"04",X"88",X"10",X"F8",X"60",X"A9",X"00",X"99",X"34",X"00",X"A9",X"40",
		X"45",X"F0",X"99",X"64",X"00",X"A9",X"FC",X"99",X"54",X"00",X"A9",X"02",X"99",X"74",X"00",X"B5",
		X"A1",X"C9",X"60",X"90",X"04",X"E9",X"08",X"95",X"A1",X"85",X"A0",X"AD",X"0A",X"10",X"29",X"02",
		X"D0",X"07",X"A9",X"04",X"99",X"54",X"00",X"A9",X"FE",X"99",X"44",X"00",X"F6",X"94",X"60",X"4A",
		X"4A",X"4A",X"69",X"00",X"85",X"32",X"A9",X"01",X"85",X"33",X"98",X"0A",X"0A",X"0A",X"18",X"65",
		X"8B",X"85",X"8B",X"A9",X"F7",X"38",X"E5",X"8B",X"B0",X"02",X"A9",X"00",X"29",X"F8",X"0A",X"26",
		X"33",X"0A",X"26",X"33",X"05",X"32",X"A4",X"33",X"C0",X"07",X"D0",X"08",X"C9",X"C0",X"90",X"04",
		X"29",X"1F",X"09",X"A0",X"85",X"32",X"A0",X"00",X"B1",X"32",X"F0",X"02",X"45",X"EF",X"60",X"86",
		X"8B",X"86",X"8C",X"E6",X"8C",X"A0",X"0C",X"B9",X"64",X"00",X"D5",X"64",X"D0",X"17",X"B9",X"34",
		X"00",X"C9",X"F4",X"B0",X"10",X"C4",X"8B",X"F0",X"0C",X"B5",X"54",X"38",X"F9",X"54",X"00",X"55",
		X"44",X"C9",X"F4",X"B0",X"04",X"88",X"10",X"DF",X"18",X"60",X"B5",X"54",X"38",X"E5",X"63",X"20",
		X"7A",X"38",X"E0",X"0D",X"D0",X"05",X"C9",X"0A",X"90",X"05",X"60",X"C9",X"07",X"B0",X"FB",X"85",
		X"8D",X"B5",X"64",X"38",X"E5",X"73",X"20",X"7A",X"38",X"C9",X"07",X"B0",X"ED",X"18",X"65",X"8D",
		X"E0",X"0D",X"F0",X"2A",X"C9",X"0C",X"B0",X"E2",X"A9",X"30",X"85",X"87",X"A9",X"20",X"85",X"43",
		X"A9",X"FF",X"95",X"34",X"A9",X"28",X"85",X"42",X"A5",X"86",X"30",X"04",X"A9",X"13",X"85",X"B7",
		X"A9",X"00",X"85",X"B2",X"85",X"B3",X"85",X"B4",X"85",X"B5",X"85",X"B8",X"18",X"60",X"C9",X"0E",
		X"4C",X"C6",X"2C",X"A0",X"00",X"A5",X"00",X"29",X"07",X"D0",X"14",X"A5",X"B7",X"D0",X"10",X"A5",
		X"DB",X"F0",X"0C",X"C9",X"07",X"D0",X"09",X"A5",X"DA",X"C9",X"C0",X"90",X"03",X"84",X"DB",X"60",
		X"B1",X"DA",X"29",X"3F",X"C9",X"38",X"90",X"40",X"C9",X"3F",X"B0",X"3C",X"A9",X"3F",X"45",X"EF",
		X"91",X"DA",X"A9",X"00",X"85",X"8B",X"A9",X"05",X"20",X"BA",X"2D",X"A9",X"FF",X"85",X"3F",X"A5",
		X"DB",X"85",X"8B",X"A5",X"DA",X"0A",X"26",X"8B",X"0A",X"26",X"8B",X"0A",X"26",X"8B",X"85",X"6F",
		X"A5",X"8B",X"29",X"1F",X"49",X"1F",X"0A",X"0A",X"0A",X"E9",X"03",X"85",X"5F",X"E6",X"DA",X"D0",
		X"02",X"E6",X"DB",X"A9",X"13",X"85",X"B2",X"60",X"E6",X"DA",X"D0",X"A3",X"E6",X"DB",X"D0",X"B0",
		X"A9",X"07",X"20",X"24",X"38",X"A0",X"00",X"A2",X"5C",X"86",X"91",X"A9",X"05",X"85",X"92",X"B9",
		X"04",X"00",X"84",X"8D",X"38",X"20",X"9E",X"38",X"A4",X"8D",X"B9",X"03",X"00",X"20",X"9E",X"38",
		X"A4",X"8D",X"B9",X"02",X"00",X"18",X"20",X"9E",X"38",X"A9",X"00",X"20",X"85",X"38",X"A4",X"8D",
		X"20",X"82",X"38",X"E6",X"8D",X"A4",X"8D",X"20",X"82",X"38",X"E6",X"8D",X"A4",X"8D",X"20",X"82",
		X"38",X"A5",X"91",X"29",X"1F",X"09",X"40",X"AA",X"CA",X"A4",X"8D",X"C8",X"C0",X"18",X"90",X"B9",
		X"60",X"C9",X"86",X"8D",X"A6",X"88",X"D6",X"94",X"A6",X"8D",X"A4",X"86",X"30",X"5D",X"86",X"8D",
		X"F8",X"A6",X"88",X"18",X"75",X"A7",X"95",X"A7",X"B5",X"A9",X"65",X"8B",X"95",X"A9",X"90",X"0D",
		X"B5",X"A1",X"E9",X"02",X"95",X"A1",X"B5",X"AB",X"18",X"69",X"01",X"95",X"AB",X"D8",X"A6",X"88",
		X"B5",X"A9",X"D5",X"AD",X"B5",X"AB",X"F5",X"AF",X"90",X"2F",X"20",X"B3",X"21",X"F8",X"18",X"75",
		X"AD",X"95",X"AD",X"B9",X"C0",X"21",X"75",X"AF",X"95",X"AF",X"D8",X"AD",X"01",X"08",X"29",X"1C",
		X"F0",X"06",X"A5",X"AD",X"05",X"AB",X"F0",X"11",X"B5",X"A4",X"C9",X"06",X"F0",X"0B",X"B0",X"FE",
		X"F6",X"A4",X"A9",X"11",X"85",X"B6",X"20",X"BC",X"26",X"A6",X"8D",X"60",X"A5",X"40",X"45",X"EF",
		X"C9",X"34",X"90",X"03",X"4C",X"A5",X"2E",X"C9",X"30",X"B0",X"5D",X"A5",X"70",X"45",X"F0",X"C9",
		X"F8",X"90",X"04",X"A5",X"00",X"F0",X"03",X"4C",X"D6",X"2E",X"A6",X"88",X"B5",X"9A",X"C9",X"0B",
		X"B0",X"F5",X"AD",X"0A",X"10",X"29",X"03",X"D0",X"EE",X"A9",X"14",X"85",X"B8",X"A9",X"30",X"45",
		X"EF",X"85",X"40",X"B5",X"AB",X"C9",X"02",X"90",X"12",X"AD",X"0A",X"10",X"29",X"03",X"F0",X"0B",
		X"A9",X"02",X"2C",X"0A",X"10",X"10",X"0D",X"A9",X"FE",X"D0",X"09",X"A9",X"01",X"2C",X"0A",X"10",
		X"10",X"02",X"A9",X"FF",X"85",X"50",X"A9",X"00",X"85",X"60",X"85",X"80",X"AD",X"0A",X"10",X"29",
		X"78",X"18",X"69",X"70",X"45",X"F0",X"85",X"70",X"A5",X"43",X"29",X"AF",X"D0",X"1D",X"A5",X"60",
		X"A4",X"EF",X"F0",X"06",X"38",X"E5",X"50",X"4C",X"9D",X"2E",X"18",X"65",X"50",X"85",X"60",X"85",
		X"8B",X"D0",X"0B",X"F0",X"06",X"45",X"EF",X"C9",X"FA",X"B0",X"2B",X"4C",X"E8",X"20",X"A5",X"00",
		X"29",X"03",X"D0",X"0D",X"A5",X"40",X"18",X"69",X"01",X"29",X"03",X"09",X"30",X"45",X"EF",X"85",
		X"40",X"A0",X"00",X"A5",X"70",X"20",X"2F",X"2C",X"C9",X"40",X"B0",X"0A",X"C9",X"3C",X"90",X"06",
		X"29",X"FB",X"45",X"EF",X"91",X"32",X"60",X"A5",X"72",X"A4",X"EF",X"F0",X"05",X"18",X"69",X"07",
		X"49",X"FF",X"C9",X"F3",X"B0",X"75",X"A9",X"04",X"45",X"F0",X"18",X"65",X"73",X"C5",X"72",X"D0",
		X"25",X"A5",X"43",X"29",X"AF",X"D0",X"18",X"AD",X"01",X"0C",X"A6",X"86",X"10",X"03",X"AD",X"0A",
		X"10",X"C0",X"C0",X"D0",X"06",X"29",X"08",X"F0",X"09",X"D0",X"04",X"29",X"04",X"F0",X"03",X"4C",
		X"5A",X"30",X"A9",X"0B",X"85",X"B4",X"A5",X"62",X"85",X"8B",X"A9",X"07",X"45",X"F4",X"A4",X"72",
		X"18",X"65",X"72",X"85",X"72",X"84",X"8D",X"A9",X"01",X"45",X"F3",X"18",X"65",X"8D",X"A0",X"00",
		X"20",X"2F",X"2C",X"F0",X"29",X"29",X"3F",X"C9",X"38",X"90",X"20",X"E9",X"01",X"C9",X"3B",X"F0",
		X"04",X"C9",X"37",X"D0",X"0D",X"A9",X"00",X"85",X"8B",X"A9",X"01",X"20",X"BA",X"2D",X"A0",X"00",
		X"A5",X"EF",X"45",X"EF",X"91",X"32",X"D0",X"03",X"20",X"95",X"2B",X"4C",X"57",X"30",X"A2",X"0D",
		X"B5",X"34",X"C9",X"76",X"90",X"08",X"C9",X"B9",X"90",X"69",X"C9",X"F8",X"B0",X"65",X"B5",X"64",
		X"45",X"F0",X"C9",X"F8",X"B0",X"5D",X"45",X"F0",X"38",X"E5",X"72",X"20",X"7A",X"38",X"A8",X"E0",
		X"0C",X"D0",X"16",X"B5",X"34",X"45",X"EF",X"C9",X"20",X"B0",X"0E",X"A5",X"80",X"45",X"F0",X"C9",
		X"04",X"90",X"06",X"C0",X"07",X"B0",X"3C",X"90",X"04",X"C0",X"05",X"B0",X"36",X"B5",X"54",X"38",
		X"E5",X"62",X"20",X"7A",X"38",X"A8",X"E0",X"0D",X"F0",X"25",X"E0",X"0C",X"90",X"60",X"B5",X"34",
		X"45",X"EF",X"C9",X"20",X"B0",X"10",X"C0",X"06",X"B0",X"19",X"A0",X"02",X"A9",X"04",X"C5",X"80",
		X"F0",X"0A",X"85",X"80",X"D0",X"95",X"C0",X"0A",X"B0",X"09",X"A0",X"10",X"4C",X"48",X"30",X"C0",
		X"0A",X"90",X"03",X"4C",X"42",X"30",X"A0",X"B6",X"84",X"D7",X"A0",X"03",X"A5",X"71",X"38",X"E5",
		X"73",X"20",X"7A",X"38",X"C9",X"40",X"B0",X"0C",X"E6",X"D7",X"A0",X"09",X"C9",X"16",X"90",X"04",
		X"E6",X"D7",X"A0",X"06",X"A9",X"80",X"85",X"9F",X"85",X"A1",X"A9",X"00",X"85",X"B5",X"A9",X"F0",
		X"C5",X"61",X"90",X"06",X"A9",X"10",X"C5",X"61",X"90",X"3E",X"85",X"61",X"D0",X"3A",X"C0",X"06",
		X"B0",X"30",X"A9",X"00",X"85",X"8B",X"A0",X"10",X"B5",X"34",X"29",X"40",X"D0",X"04",X"A0",X"00",
		X"E6",X"8B",X"98",X"20",X"B2",X"2D",X"E0",X"0B",X"F0",X"08",X"B5",X"35",X"30",X"04",X"29",X"BF",
		X"95",X"35",X"20",X"10",X"23",X"20",X"2F",X"2C",X"86",X"8D",X"20",X"AC",X"2B",X"A6",X"8D",X"4C",
		X"4F",X"30",X"CA",X"30",X"15",X"4C",X"60",X"2F",X"84",X"8B",X"A9",X"00",X"20",X"BA",X"2D",X"A9",
		X"13",X"85",X"B2",X"A9",X"FF",X"95",X"34",X"20",X"7D",X"2B",X"A6",X"88",X"B5",X"94",X"05",X"87",
		X"F0",X"10",X"A5",X"41",X"45",X"EF",X"C9",X"9C",X"90",X"07",X"C6",X"9F",X"D0",X"03",X"20",X"C7",
		X"21",X"60",X"F6",X"9C",X"A9",X"40",X"85",X"87",X"60",X"A6",X"86",X"10",X"0F",X"A2",X"00",X"8E",
		X"01",X"10",X"8E",X"03",X"10",X"8E",X"05",X"10",X"8E",X"07",X"10",X"60",X"A5",X"00",X"4A",X"90",
		X"19",X"A4",X"B5",X"98",X"F0",X"11",X"C6",X"B5",X"D0",X"04",X"A9",X"14",X"85",X"B5",X"B9",X"B0",
		X"31",X"8D",X"06",X"10",X"B9",X"C4",X"31",X"8D",X"07",X"10",X"A4",X"B4",X"98",X"F0",X"0A",X"C6",
		X"B4",X"B9",X"A5",X"31",X"8D",X"04",X"10",X"A9",X"64",X"8D",X"05",X"10",X"A5",X"AD",X"D0",X"14",
		X"A5",X"AB",X"C9",X"16",X"B0",X"0E",X"C9",X"14",X"90",X"0A",X"A5",X"00",X"29",X"04",X"F0",X"16",
		X"A9",X"10",X"D0",X"12",X"A4",X"B6",X"F0",X"28",X"A5",X"00",X"29",X"07",X"D0",X"73",X"C6",X"B6",
		X"88",X"F0",X"1D",X"B9",X"D8",X"31",X"8D",X"02",X"10",X"A9",X"A4",X"D0",X"61",X"A4",X"B8",X"88",
		X"D0",X"02",X"A0",X"14",X"84",X"B8",X"B9",X"E9",X"31",X"8D",X"02",X"10",X"A9",X"A4",X"D0",X"4E",
		X"A5",X"70",X"45",X"F0",X"C9",X"F8",X"B0",X"36",X"A5",X"43",X"29",X"AF",X"D0",X"30",X"A5",X"40",
		X"45",X"EF",X"C9",X"34",X"B0",X"28",X"C9",X"20",X"B0",X"D3",X"A5",X"70",X"45",X"F4",X"4A",X"49",
		X"FF",X"09",X"80",X"8D",X"02",X"10",X"A9",X"A4",X"D0",X"24",X"A4",X"B2",X"98",X"F0",X"0B",X"C6",
		X"B2",X"B9",X"71",X"31",X"8D",X"00",X"10",X"B9",X"84",X"31",X"8D",X"01",X"10",X"60",X"A4",X"B3",
		X"98",X"F0",X"0B",X"C6",X"B3",X"B9",X"97",X"31",X"8D",X"02",X"10",X"B9",X"9E",X"31",X"8D",X"03",
		X"10",X"A4",X"B7",X"F0",X"D5",X"A5",X"00",X"29",X"03",X"D0",X"16",X"C6",X"B7",X"88",X"F0",X"11",
		X"B9",X"71",X"31",X"8D",X"00",X"10",X"B9",X"84",X"31",X"F0",X"03",X"18",X"69",X"02",X"8D",X"01",
		X"10",X"60",X"00",X"00",X"00",X"00",X"F0",X"E0",X"D0",X"C0",X"B0",X"A0",X"90",X"80",X"70",X"60",
		X"50",X"40",X"30",X"20",X"10",X"00",X"00",X"00",X"00",X"81",X"81",X"81",X"82",X"82",X"82",X"82",
		X"83",X"83",X"83",X"83",X"84",X"84",X"84",X"84",X"70",X"00",X"00",X"A0",X"00",X"C0",X"E0",X"A1",
		X"00",X"00",X"A2",X"00",X"A2",X"A4",X"F0",X"E0",X"D0",X"C0",X"B0",X"A0",X"90",X"80",X"70",X"60",
		X"50",X"05",X"05",X"20",X"20",X"30",X"30",X"35",X"35",X"30",X"30",X"20",X"20",X"05",X"05",X"20",
		X"20",X"30",X"30",X"35",X"35",X"A1",X"00",X"A2",X"00",X"A3",X"00",X"A4",X"00",X"A3",X"00",X"A2",
		X"00",X"A1",X"00",X"A2",X"00",X"A3",X"00",X"A2",X"00",X"28",X"28",X"30",X"28",X"28",X"30",X"3C",
		X"51",X"50",X"50",X"60",X"50",X"50",X"60",X"74",X"A2",X"00",X"60",X"60",X"70",X"70",X"60",X"60",
		X"60",X"70",X"70",X"70",X"50",X"50",X"80",X"80",X"50",X"50",X"50",X"80",X"80",X"80",X"A0",X"00",
		X"84",X"32",X"A9",X"04",X"85",X"33",X"84",X"8D",X"A9",X"00",X"85",X"8B",X"84",X"8E",X"A2",X"08",
		X"B1",X"32",X"29",X"3F",X"C9",X"38",X"26",X"8B",X"C8",X"CA",X"D0",X"F4",X"A6",X"8D",X"BD",X"00",
		X"01",X"E6",X"8D",X"A8",X"A5",X"8B",X"9D",X"00",X"01",X"84",X"8B",X"A4",X"8E",X"A2",X"08",X"A9",
		X"00",X"26",X"8B",X"90",X"04",X"A9",X"3F",X"45",X"EF",X"91",X"32",X"C8",X"CA",X"D0",X"F0",X"98",
		X"D0",X"02",X"E6",X"33",X"C0",X"C0",X"D0",X"C0",X"A5",X"33",X"C9",X"07",X"D0",X"BA",X"60",X"C9",
		X"08",X"90",X"0C",X"C9",X"F8",X"B0",X"08",X"C9",X"80",X"A9",X"08",X"90",X"02",X"A9",X"F8",X"C9",
		X"80",X"6A",X"A8",X"A9",X"00",X"6A",X"60",X"A9",X"FF",X"A2",X"00",X"85",X"C1",X"85",X"C2",X"F8",
		X"A5",X"FB",X"18",X"6D",X"8E",X"01",X"8D",X"8E",X"01",X"A5",X"FC",X"6D",X"8F",X"01",X"8D",X"8F",
		X"01",X"AD",X"90",X"01",X"69",X"00",X"8D",X"90",X"01",X"AD",X"91",X"01",X"69",X"00",X"B0",X"1C",
		X"8D",X"91",X"01",X"AD",X"8B",X"01",X"18",X"65",X"89",X"8D",X"8B",X"01",X"AD",X"8C",X"01",X"69",
		X"00",X"8D",X"8C",X"01",X"AD",X"8D",X"01",X"69",X"00",X"8D",X"8D",X"01",X"D8",X"A0",X"00",X"B9",
		X"02",X"00",X"D5",X"A8",X"B9",X"03",X"00",X"F5",X"AA",X"B9",X"04",X"00",X"F5",X"AC",X"90",X"2E",
		X"C8",X"C8",X"C8",X"C0",X"18",X"90",X"E8",X"CA",X"10",X"E3",X"A5",X"C2",X"30",X"0E",X"C5",X"C1",
		X"90",X"0A",X"69",X"02",X"C9",X"18",X"90",X"02",X"A9",X"FF",X"85",X"C2",X"A9",X"00",X"85",X"C0",
		X"A5",X"C2",X"25",X"C1",X"10",X"07",X"A9",X"00",X"85",X"01",X"20",X"60",X"2D",X"60",X"86",X"8D",
		X"84",X"8E",X"94",X"C1",X"A2",X"17",X"B5",X"17",X"95",X"1A",X"BD",X"FF",X"FF",X"95",X"02",X"CA",
		X"E4",X"8E",X"D0",X"F2",X"A9",X"01",X"95",X"1A",X"A9",X"00",X"95",X"1B",X"95",X"1C",X"85",X"B9",
		X"A6",X"8D",X"B5",X"AC",X"99",X"04",X"00",X"B5",X"AA",X"99",X"03",X"00",X"B5",X"A8",X"99",X"02",
		X"00",X"A9",X"F0",X"85",X"01",X"D0",X"A0",X"A9",X"1F",X"45",X"F5",X"85",X"91",X"A9",X"04",X"45",
		X"F7",X"85",X"92",X"A5",X"AC",X"38",X"20",X"9E",X"38",X"A5",X"AA",X"20",X"9E",X"38",X"A5",X"A8",
		X"18",X"20",X"9E",X"38",X"AD",X"01",X"08",X"29",X"1C",X"F0",X"1D",X"A9",X"07",X"45",X"F7",X"85",
		X"92",X"A9",X"1F",X"45",X"F5",X"85",X"91",X"A5",X"AD",X"38",X"20",X"9E",X"38",X"A9",X"2E",X"20",
		X"85",X"38",X"A5",X"AB",X"18",X"20",X"9E",X"38",X"A9",X"9F",X"45",X"F5",X"85",X"91",X"A9",X"05",
		X"45",X"F7",X"85",X"92",X"A5",X"04",X"38",X"20",X"9E",X"38",X"A5",X"03",X"20",X"9E",X"38",X"A5",
		X"02",X"18",X"4C",X"9E",X"38",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F5",X"A2",X"02",X"AD",
		X"01",X"0C",X"E0",X"01",X"F0",X"03",X"B0",X"02",X"0A",X"0A",X"0A",X"B5",X"CF",X"29",X"1F",X"B0",
		X"37",X"F0",X"10",X"C9",X"1B",X"B0",X"0A",X"A8",X"A5",X"D4",X"29",X"07",X"C9",X"07",X"98",X"90",
		X"02",X"E9",X"01",X"95",X"CF",X"AD",X"01",X"0C",X"29",X"10",X"D0",X"04",X"A9",X"F0",X"85",X"D2",
		X"A5",X"D2",X"F0",X"08",X"C6",X"D2",X"A9",X"00",X"95",X"CF",X"95",X"CC",X"18",X"B5",X"CC",X"F0",
		X"23",X"D6",X"CC",X"D0",X"1F",X"38",X"B0",X"1C",X"C9",X"1B",X"B0",X"09",X"B5",X"CF",X"69",X"20",
		X"90",X"D1",X"F0",X"01",X"18",X"A9",X"1F",X"B0",X"CA",X"95",X"CF",X"B5",X"CC",X"F0",X"01",X"38",
		X"A9",X"78",X"95",X"CC",X"90",X"2A",X"A9",X"00",X"E0",X"01",X"90",X"16",X"F0",X"0C",X"A5",X"D3",
		X"29",X"0C",X"4A",X"4A",X"F0",X"0C",X"69",X"02",X"D0",X"08",X"A5",X"D3",X"29",X"10",X"F0",X"02",
		X"A9",X"01",X"38",X"48",X"65",X"CA",X"85",X"CA",X"68",X"38",X"65",X"C9",X"85",X"C9",X"F6",X"C5",
		X"CA",X"30",X"03",X"4C",X"AF",X"33",X"A5",X"D3",X"4A",X"4A",X"4A",X"4A",X"4A",X"A8",X"A5",X"CA",
		X"38",X"F9",X"62",X"34",X"30",X"14",X"85",X"CA",X"E6",X"CB",X"C0",X"03",X"D0",X"0C",X"E6",X"CB",
		X"D0",X"08",X"7F",X"02",X"04",X"04",X"05",X"03",X"7F",X"7F",X"A5",X"D3",X"29",X"03",X"A8",X"F0",
		X"1A",X"4A",X"69",X"00",X"49",X"FF",X"38",X"65",X"C9",X"B0",X"08",X"65",X"CB",X"30",X"0E",X"85",
		X"CB",X"A9",X"00",X"C0",X"02",X"B0",X"02",X"E6",X"C8",X"E6",X"C8",X"85",X"C9",X"E6",X"D4",X"A5",
		X"D4",X"4A",X"B0",X"27",X"A0",X"00",X"A2",X"02",X"B5",X"C5",X"F0",X"09",X"C9",X"10",X"90",X"05",
		X"69",X"EF",X"C8",X"95",X"C5",X"CA",X"10",X"F0",X"98",X"D0",X"10",X"A2",X"02",X"B5",X"C5",X"F0",
		X"07",X"18",X"69",X"EF",X"95",X"C5",X"30",X"03",X"CA",X"10",X"F2",X"60",X"14",X"35",X"1F",X"35",
		X"2B",X"35",X"36",X"35",X"42",X"35",X"54",X"35",X"69",X"35",X"7E",X"35",X"92",X"35",X"A3",X"35",
		X"B7",X"35",X"CB",X"35",X"DE",X"35",X"F0",X"35",X"05",X"36",X"1A",X"36",X"2E",X"36",X"3B",X"36",
		X"48",X"36",X"59",X"36",X"6C",X"36",X"83",X"36",X"A3",X"36",X"BB",X"36",X"D2",X"36",X"E2",X"36",
		X"F1",X"36",X"02",X"37",X"11",X"37",X"20",X"37",X"35",X"37",X"48",X"37",X"53",X"37",X"62",X"37",
		X"7B",X"37",X"8E",X"37",X"9E",X"37",X"AA",X"37",X"B6",X"37",X"C2",X"37",X"CF",X"37",X"E3",X"37",
		X"FF",X"37",X"11",X"38",X"6E",X"05",X"51",X"06",X"50",X"4C",X"41",X"59",X"45",X"52",X"A0",X"6E",
		X"05",X"51",X"06",X"53",X"50",X"49",X"45",X"4C",X"45",X"52",X"A0",X"6E",X"05",X"51",X"06",X"4A",
		X"4F",X"55",X"45",X"55",X"52",X"A0",X"6E",X"05",X"51",X"06",X"4A",X"55",X"47",X"41",X"44",X"4F",
		X"52",X"A0",X"13",X"05",X"AC",X"06",X"31",X"20",X"43",X"4F",X"49",X"4E",X"20",X"32",X"20",X"50",
		X"4C",X"41",X"59",X"D3",X"F3",X"04",X"CC",X"06",X"31",X"20",X"4D",X"55",X"45",X"4E",X"5A",X"45",
		X"20",X"32",X"20",X"53",X"50",X"49",X"45",X"4C",X"C5",X"F3",X"04",X"CC",X"06",X"31",X"20",X"50",
		X"49",X"45",X"43",X"45",X"20",X"32",X"20",X"4A",X"4F",X"55",X"45",X"55",X"52",X"D3",X"F3",X"04",
		X"CC",X"06",X"31",X"20",X"46",X"49",X"43",X"48",X"41",X"20",X"32",X"20",X"4A",X"55",X"45",X"47",
		X"4F",X"D3",X"13",X"05",X"AC",X"06",X"31",X"20",X"43",X"4F",X"49",X"4E",X"20",X"31",X"20",X"50",
		X"4C",X"41",X"D9",X"F3",X"04",X"CC",X"06",X"31",X"20",X"4D",X"55",X"45",X"4E",X"5A",X"45",X"20",
		X"31",X"20",X"53",X"50",X"49",X"45",X"CC",X"F3",X"04",X"CC",X"06",X"31",X"20",X"50",X"49",X"45",
		X"43",X"45",X"20",X"31",X"20",X"4A",X"4F",X"55",X"45",X"55",X"D2",X"F3",X"04",X"CC",X"06",X"31",
		X"20",X"46",X"49",X"43",X"48",X"41",X"20",X"31",X"20",X"4A",X"55",X"45",X"47",X"CF",X"13",X"05",
		X"AC",X"06",X"32",X"20",X"43",X"4F",X"49",X"4E",X"53",X"20",X"31",X"20",X"50",X"4C",X"41",X"D9",
		X"F3",X"04",X"CC",X"06",X"32",X"20",X"4D",X"55",X"45",X"4E",X"5A",X"45",X"4E",X"20",X"31",X"20",
		X"53",X"50",X"49",X"45",X"CC",X"F3",X"04",X"CC",X"06",X"32",X"20",X"50",X"49",X"45",X"43",X"45",
		X"53",X"20",X"31",X"20",X"4A",X"4F",X"55",X"45",X"55",X"D2",X"F3",X"04",X"CC",X"06",X"32",X"20",
		X"46",X"49",X"43",X"48",X"41",X"53",X"20",X"31",X"20",X"4A",X"55",X"45",X"47",X"CF",X"6F",X"05",
		X"50",X"06",X"47",X"41",X"4D",X"45",X"20",X"4F",X"56",X"45",X"D2",X"6F",X"05",X"50",X"06",X"53",
		X"50",X"49",X"45",X"4C",X"45",X"4E",X"44",X"C5",X"0F",X"05",X"B0",X"06",X"46",X"49",X"4E",X"20",
		X"44",X"45",X"20",X"50",X"41",X"52",X"54",X"49",X"C5",X"EF",X"04",X"D0",X"06",X"4A",X"55",X"45",
		X"47",X"4F",X"20",X"54",X"45",X"52",X"4D",X"49",X"4E",X"41",X"44",X"CF",X"AB",X"04",X"14",X"07",
		X"45",X"4E",X"54",X"45",X"52",X"20",X"59",X"4F",X"55",X"52",X"20",X"49",X"4E",X"49",X"54",X"49",
		X"41",X"4C",X"D3",X"2B",X"04",X"94",X"07",X"47",X"45",X"42",X"45",X"4E",X"20",X"53",X"49",X"45",
		X"20",X"49",X"48",X"52",X"45",X"20",X"49",X"4E",X"49",X"54",X"49",X"41",X"4C",X"45",X"4E",X"20",
		X"45",X"49",X"CE",X"8B",X"04",X"34",X"07",X"45",X"4E",X"54",X"52",X"45",X"5A",X"20",X"56",X"4F",
		X"53",X"20",X"49",X"4E",X"49",X"54",X"49",X"41",X"4C",X"45",X"D3",X"8B",X"04",X"34",X"07",X"45",
		X"4E",X"54",X"52",X"45",X"20",X"53",X"55",X"53",X"20",X"49",X"4E",X"49",X"43",X"49",X"41",X"4C",
		X"45",X"D3",X"F1",X"04",X"CE",X"06",X"42",X"4F",X"4E",X"55",X"53",X"20",X"45",X"56",X"45",X"52",
		X"59",X"A0",X"F1",X"04",X"CE",X"06",X"42",X"4F",X"4E",X"55",X"53",X"20",X"4A",X"45",X"44",X"45",
		X"A0",X"D1",X"04",X"EE",X"06",X"42",X"4F",X"4E",X"55",X"53",X"20",X"43",X"48",X"41",X"51",X"55",
		X"45",X"A0",X"F1",X"04",X"CE",X"06",X"45",X"58",X"54",X"52",X"41",X"20",X"43",X"41",X"44",X"41",
		X"A0",X"5D",X"05",X"62",X"06",X"48",X"49",X"47",X"48",X"20",X"53",X"43",X"4F",X"52",X"45",X"D3",
		X"DD",X"04",X"E2",X"06",X"48",X"4F",X"45",X"43",X"48",X"53",X"54",X"45",X"52",X"47",X"45",X"42",
		X"4E",X"49",X"53",X"53",X"C5",X"1D",X"05",X"A2",X"06",X"4D",X"45",X"49",X"4C",X"4C",X"45",X"55",
		X"52",X"53",X"20",X"53",X"43",X"4F",X"52",X"C5",X"9D",X"05",X"22",X"06",X"52",X"45",X"43",X"4F",
		X"52",X"44",X"D3",X"2C",X"05",X"93",X"06",X"47",X"52",X"45",X"41",X"54",X"20",X"53",X"43",X"4F",
		X"52",X"C5",X"8C",X"04",X"33",X"07",X"47",X"52",X"4F",X"53",X"53",X"41",X"52",X"54",X"49",X"47",
		X"45",X"53",X"20",X"45",X"52",X"47",X"45",X"42",X"4E",X"49",X"D3",X"EC",X"04",X"D3",X"06",X"53",
		X"50",X"4C",X"45",X"4E",X"44",X"49",X"44",X"45",X"20",X"53",X"43",X"4F",X"52",X"C5",X"0C",X"05",
		X"B3",X"06",X"47",X"52",X"41",X"4E",X"20",X"50",X"55",X"4E",X"54",X"41",X"4A",X"C5",X"52",X"05",
		X"6D",X"06",X"43",X"52",X"45",X"44",X"49",X"54",X"53",X"A0",X"52",X"05",X"6D",X"06",X"4B",X"52",
		X"45",X"44",X"49",X"54",X"45",X"A0",X"52",X"05",X"6D",X"06",X"43",X"52",X"45",X"44",X"49",X"54",
		X"53",X"A0",X"52",X"05",X"6D",X"06",X"43",X"52",X"45",X"44",X"49",X"54",X"4F",X"53",X"A0",X"F0",
		X"04",X"CF",X"06",X"32",X"20",X"43",X"52",X"45",X"44",X"49",X"54",X"20",X"4D",X"49",X"4E",X"49",
		X"4D",X"55",X"CD",X"30",X"04",X"8F",X"07",X"47",X"45",X"4C",X"44",X"45",X"49",X"4E",X"57",X"55",
		X"52",X"46",X"20",X"46",X"55",X"52",X"20",X"32",X"20",X"53",X"50",X"49",X"45",X"4C",X"C5",X"F0",
		X"04",X"CF",X"06",X"32",X"20",X"4A",X"55",X"45",X"58",X"20",X"4D",X"49",X"4E",X"49",X"4D",X"55",
		X"CD",X"F0",X"04",X"CF",X"06",X"32",X"20",X"4A",X"55",X"45",X"47",X"41",X"53",X"20",X"4D",X"49",
		X"4E",X"49",X"4D",X"B0",X"0A",X"66",X"8C",X"A8",X"0A",X"85",X"8B",X"A5",X"FD",X"29",X"03",X"05",
		X"8B",X"0A",X"AA",X"BD",X"BC",X"34",X"85",X"93",X"BD",X"BD",X"34",X"85",X"94",X"A0",X"00",X"A6",
		X"EF",X"F0",X"02",X"A0",X"02",X"B1",X"93",X"85",X"91",X"C8",X"B1",X"93",X"85",X"92",X"A0",X"04",
		X"84",X"8B",X"A4",X"8B",X"B1",X"93",X"29",X"3F",X"C9",X"20",X"F0",X"04",X"A6",X"8C",X"10",X"02",
		X"A9",X"00",X"C9",X"30",X"90",X"02",X"29",X"2F",X"20",X"85",X"38",X"A4",X"8B",X"E6",X"8B",X"B1",
		X"93",X"10",X"DF",X"60",X"A0",X"00",X"84",X"8C",X"F0",X"D6",X"10",X"05",X"49",X"FF",X"18",X"69",
		X"01",X"60",X"B9",X"1A",X"00",X"A8",X"F0",X"02",X"45",X"EF",X"A0",X"00",X"91",X"91",X"A9",X"20",
		X"45",X"EF",X"18",X"65",X"91",X"85",X"91",X"A5",X"F3",X"65",X"92",X"85",X"92",X"60",X"48",X"08",
		X"4A",X"4A",X"4A",X"4A",X"28",X"20",X"AB",X"38",X"68",X"29",X"0F",X"90",X"04",X"29",X"0F",X"F0",
		X"03",X"18",X"09",X"20",X"08",X"C9",X"2A",X"90",X"02",X"E9",X"29",X"20",X"85",X"38",X"28",X"60",
		X"48",X"8A",X"48",X"98",X"48",X"D8",X"A5",X"D2",X"F0",X"0A",X"A9",X"10",X"8D",X"02",X"10",X"A9",
		X"AF",X"8D",X"03",X"10",X"2C",X"00",X"0C",X"70",X"03",X"4C",X"B4",X"39",X"E6",X"8A",X"E6",X"00",
		X"D0",X"11",X"E6",X"01",X"F8",X"A5",X"FB",X"18",X"69",X"01",X"85",X"FB",X"A5",X"FC",X"69",X"00",
		X"85",X"FC",X"D8",X"A5",X"8A",X"C9",X"08",X"B0",X"FE",X"A5",X"C8",X"C9",X"25",X"B0",X"FE",X"C9",
		X"13",X"90",X"04",X"A9",X"12",X"85",X"C8",X"AD",X"03",X"0C",X"A6",X"88",X"AC",X"B8",X"01",X"20",
		X"31",X"3A",X"8C",X"B8",X"01",X"48",X"98",X"18",X"65",X"B9",X"85",X"B9",X"68",X"AC",X"B9",X"01",
		X"20",X"31",X"3A",X"8C",X"B9",X"01",X"98",X"20",X"7C",X"38",X"18",X"65",X"BB",X"85",X"BB",X"B5",
		X"C2",X"30",X"08",X"C9",X"40",X"90",X"15",X"29",X"3F",X"10",X"0B",X"29",X"3F",X"18",X"69",X"03",
		X"C9",X"2A",X"90",X"02",X"A9",X"00",X"95",X"C2",X"AA",X"20",X"5A",X"26",X"A2",X"0F",X"B5",X"64",
		X"9D",X"E0",X"07",X"B5",X"54",X"A0",X"00",X"E0",X"0D",X"F0",X"07",X"B4",X"44",X"10",X"03",X"18",
		X"69",X"01",X"9D",X"D0",X"07",X"98",X"29",X"80",X"85",X"99",X"AD",X"00",X"0C",X"29",X"20",X"D0",
		X"05",X"B5",X"34",X"4C",X"9D",X"39",X"B5",X"34",X"E0",X"0C",X"B0",X"1F",X"29",X"3F",X"C9",X"30",
		X"B0",X"19",X"29",X"0F",X"85",X"98",X"B5",X"64",X"29",X"07",X"F0",X"0D",X"A8",X"A9",X"08",X"C0",
		X"06",X"B0",X"06",X"C0",X"03",X"90",X"02",X"A9",X"0C",X"45",X"98",X"45",X"99",X"9D",X"C0",X"07",
		X"B5",X"34",X"29",X"40",X"F0",X"06",X"E0",X"0C",X"B0",X"02",X"A9",X"0C",X"09",X"39",X"9D",X"F0",
		X"07",X"CA",X"10",X"9A",X"AD",X"00",X"0C",X"29",X"20",X"D0",X"1F",X"A5",X"D5",X"30",X"3B",X"E6",
		X"D5",X"2C",X"00",X"0C",X"50",X"04",X"A9",X"00",X"85",X"D5",X"A5",X"D5",X"0A",X"0A",X"A2",X"03",
		X"9D",X"04",X"14",X"69",X"01",X"CA",X"10",X"F8",X"30",X"20",X"20",X"AD",X"33",X"A2",X"02",X"B5",
		X"C5",X"9D",X"00",X"1C",X"CA",X"10",X"F8",X"A2",X"0A",X"A9",X"F4",X"5D",X"03",X"20",X"CA",X"10",
		X"FA",X"AA",X"F0",X"06",X"BA",X"A9",X"03",X"9D",X"04",X"01",X"A2",X"02",X"BD",X"00",X"0C",X"A8",
		X"38",X"F5",X"BD",X"94",X"BD",X"29",X"0F",X"C9",X"08",X"90",X"02",X"09",X"F0",X"A8",X"F0",X"14",
		X"55",X"BA",X"10",X"08",X"98",X"5D",X"00",X"0C",X"10",X"02",X"B4",X"BA",X"98",X"95",X"BA",X"18",
		X"75",X"B9",X"95",X"B9",X"CA",X"CA",X"10",X"D4",X"8D",X"00",X"18",X"68",X"A8",X"68",X"AA",X"68",
		X"40",X"0A",X"90",X"06",X"0A",X"90",X"0E",X"A0",X"00",X"60",X"C0",X"FA",X"F0",X"05",X"B0",X"02",
		X"A0",X"00",X"88",X"0A",X"60",X"C0",X"06",X"F0",X"05",X"90",X"02",X"A0",X"00",X"C8",X"60",X"A0",
		X"3C",X"A9",X"FF",X"59",X"78",X"01",X"88",X"10",X"FA",X"AC",X"B5",X"01",X"8D",X"B5",X"01",X"98",
		X"4D",X"B5",X"01",X"60",X"A2",X"2F",X"BD",X"B0",X"3A",X"95",X"02",X"CA",X"10",X"F8",X"20",X"4F",
		X"3A",X"D0",X"2B",X"A5",X"FD",X"29",X"7C",X"CD",X"8A",X"01",X"8D",X"8A",X"01",X"D0",X"1E",X"AD",
		X"7A",X"01",X"F0",X"1A",X"A2",X"08",X"BD",X"78",X"01",X"95",X"02",X"C9",X"9A",X"B0",X"0F",X"29",
		X"0F",X"C9",X"0A",X"B0",X"09",X"BD",X"81",X"01",X"95",X"1A",X"CA",X"10",X"E9",X"60",X"A9",X"00",
		X"A2",X"3E",X"9D",X"78",X"01",X"CA",X"10",X"FA",X"A5",X"FD",X"29",X"7C",X"8D",X"8A",X"01",X"60",
		X"43",X"65",X"01",X"32",X"54",X"01",X"20",X"43",X"01",X"10",X"32",X"01",X"10",X"30",X"01",X"05",
		X"28",X"01",X"01",X"22",X"01",X"02",X"21",X"01",X"05",X"0A",X"04",X"04",X"06",X"14",X"03",X"01",
		X"04",X"04",X"03",X"02",X"05",X"04",X"00",X"04",X"05",X"17",X"04",X"06",X"17",X"07",X"0A",X"12",
		X"A2",X"3F",X"20",X"EE",X"3A",X"9D",X"78",X"01",X"CA",X"10",X"F7",X"86",X"F9",X"60",X"9D",X"00",
		X"16",X"A0",X"08",X"8C",X"80",X"16",X"C8",X"8C",X"80",X"16",X"88",X"8C",X"80",X"16",X"A0",X"00",
		X"BD",X"00",X"17",X"8C",X"80",X"16",X"60",X"A5",X"00",X"29",X"03",X"D0",X"17",X"8D",X"80",X"16",
		X"A6",X"F9",X"30",X"10",X"46",X"FA",X"90",X"0D",X"A9",X"02",X"8D",X"80",X"16",X"A9",X"0A",X"8D",
		X"80",X"16",X"C6",X"F9",X"60",X"78",X"20",X"EE",X"3A",X"DD",X"78",X"01",X"D0",X"07",X"CA",X"10",
		X"F5",X"58",X"86",X"F9",X"60",X"58",X"86",X"F9",X"A9",X"06",X"8D",X"80",X"16",X"BD",X"78",X"01",
		X"9D",X"00",X"16",X"A9",X"0E",X"8D",X"80",X"16",X"E6",X"FA",X"60",X"D8",X"A2",X"FF",X"9A",X"E8",
		X"8A",X"95",X"00",X"9D",X"00",X"01",X"9D",X"00",X"04",X"9D",X"00",X"05",X"9D",X"00",X"06",X"9D",
		X"00",X"07",X"CA",X"D0",X"EC",X"8D",X"0F",X"10",X"8D",X"08",X"10",X"8D",X"00",X"24",X"8D",X"07",
		X"1C",X"AD",X"00",X"0C",X"29",X"20",X"F0",X"19",X"AD",X"00",X"08",X"85",X"FD",X"CA",X"86",X"86",
		X"86",X"C1",X"86",X"C2",X"A9",X"01",X"85",X"FF",X"20",X"E0",X"3A",X"20",X"64",X"3A",X"4C",X"0E",
		X"20",X"8E",X"04",X"14",X"8E",X"01",X"10",X"8E",X"03",X"10",X"8E",X"05",X"10",X"8E",X"07",X"10",
		X"E8",X"8E",X"05",X"14",X"8E",X"0D",X"14",X"E8",X"8E",X"06",X"14",X"8E",X"0E",X"14",X"E8",X"8E",
		X"07",X"14",X"8E",X"0F",X"14",X"A2",X"00",X"B5",X"00",X"D0",X"43",X"A9",X"11",X"95",X"00",X"A8",
		X"55",X"00",X"D0",X"3A",X"98",X"0A",X"90",X"F5",X"E8",X"D0",X"EC",X"8D",X"00",X"20",X"8A",X"85",
		X"8B",X"2A",X"85",X"8C",X"A0",X"00",X"A2",X"11",X"B1",X"8B",X"D0",X"28",X"8A",X"91",X"8B",X"51",
		X"8B",X"D0",X"21",X"8A",X"0A",X"AA",X"90",X"F4",X"C8",X"D0",X"EB",X"8D",X"00",X"20",X"E6",X"8C",
		X"A5",X"8C",X"C9",X"02",X"D0",X"02",X"A9",X"04",X"C9",X"08",X"90",X"D6",X"B0",X"5F",X"C9",X"10",
		X"A9",X"00",X"10",X"12",X"A6",X"8C",X"E0",X"04",X"90",X"F4",X"AA",X"98",X"29",X"30",X"4A",X"4A",
		X"4A",X"4A",X"69",X"01",X"E0",X"10",X"2A",X"A8",X"A9",X"40",X"8D",X"00",X"10",X"A2",X"03",X"8E",
		X"0F",X"10",X"A2",X"10",X"A9",X"AF",X"8D",X"01",X"10",X"2C",X"00",X"0C",X"50",X"FB",X"2C",X"00",
		X"0C",X"70",X"FB",X"8D",X"00",X"20",X"CA",X"D0",X"F0",X"8E",X"01",X"10",X"A2",X"10",X"2C",X"00",
		X"0C",X"50",X"FB",X"2C",X"00",X"0C",X"70",X"FB",X"8D",X"00",X"20",X"CA",X"D0",X"F0",X"88",X"10",
		X"D1",X"8D",X"00",X"20",X"AD",X"00",X"0C",X"29",X"20",X"F0",X"F6",X"D0",X"FE",X"AD",X"01",X"0C",
		X"29",X"10",X"F0",X"03",X"4C",X"DE",X"3C",X"AA",X"95",X"00",X"E8",X"D0",X"FB",X"A2",X"0F",X"A9",
		X"F8",X"95",X"64",X"CA",X"10",X"FB",X"A9",X"07",X"85",X"8C",X"A0",X"BF",X"A9",X"2D",X"A2",X"08",
		X"91",X"8B",X"88",X"CA",X"D0",X"FA",X"38",X"E9",X"01",X"C9",X"2A",X"B0",X"F1",X"C0",X"FF",X"D0",
		X"EB",X"C6",X"8C",X"A5",X"8C",X"C9",X"04",X"B0",X"E3",X"58",X"AD",X"00",X"0C",X"29",X"20",X"D0",
		X"F9",X"46",X"8A",X"8D",X"00",X"20",X"AD",X"01",X"0C",X"29",X"E0",X"49",X"E0",X"F0",X"EB",X"A9",
		X"1D",X"78",X"9D",X"00",X"04",X"9D",X"00",X"05",X"9D",X"00",X"06",X"E8",X"D0",X"F4",X"9D",X"00",
		X"07",X"E8",X"E0",X"C0",X"90",X"F8",X"A2",X"08",X"8E",X"05",X"14",X"A2",X"0F",X"8E",X"04",X"14",
		X"AD",X"00",X"0C",X"29",X"20",X"D0",X"F9",X"8D",X"00",X"20",X"46",X"8A",X"10",X"F2",X"A2",X"00",
		X"8A",X"9D",X"00",X"07",X"A9",X"00",X"95",X"00",X"9D",X"00",X"04",X"9D",X"00",X"05",X"9D",X"00",
		X"06",X"E8",X"D0",X"EC",X"CA",X"86",X"D5",X"86",X"E3",X"8D",X"03",X"1C",X"8D",X"04",X"1C",X"A2",
		X"0F",X"8A",X"09",X"80",X"95",X"54",X"95",X"64",X"CA",X"10",X"F6",X"AD",X"0A",X"10",X"4D",X"0A",
		X"10",X"85",X"E5",X"A9",X"03",X"8D",X"0F",X"10",X"A2",X"00",X"86",X"8B",X"A9",X"20",X"85",X"8C",
		X"A2",X"1F",X"A9",X"FF",X"A0",X"00",X"8E",X"00",X"20",X"51",X"8B",X"C8",X"D0",X"FB",X"A8",X"8A",
		X"29",X"07",X"C9",X"01",X"98",X"B0",X"03",X"48",X"A9",X"FF",X"E6",X"8C",X"CA",X"10",X"E5",X"A9",
		X"04",X"85",X"92",X"A2",X"03",X"8A",X"49",X"3F",X"85",X"91",X"68",X"F0",X"11",X"48",X"8A",X"09",
		X"20",X"20",X"85",X"38",X"A9",X"00",X"20",X"85",X"38",X"68",X"18",X"20",X"9E",X"38",X"CA",X"10",
		X"E4",X"20",X"E0",X"3A",X"A0",X"06",X"B9",X"8B",X"01",X"99",X"8E",X"00",X"88",X"10",X"F7",X"F8",
		X"AD",X"8B",X"01",X"0D",X"8C",X"01",X"0D",X"8D",X"01",X"F0",X"1F",X"C8",X"C8",X"F0",X"1B",X"A5",
		X"91",X"38",X"E5",X"8E",X"85",X"91",X"A5",X"92",X"E5",X"8F",X"85",X"92",X"A5",X"93",X"E5",X"90",
		X"85",X"93",X"A5",X"94",X"E9",X"00",X"85",X"94",X"10",X"E2",X"D8",X"84",X"8D",X"58",X"46",X"8A",
		X"90",X"FC",X"AD",X"00",X"0C",X"29",X"20",X"D0",X"FE",X"8D",X"00",X"20",X"AD",X"01",X"0C",X"4A",
		X"26",X"EA",X"A5",X"EA",X"29",X"03",X"C9",X"02",X"D0",X"24",X"A5",X"E6",X"AA",X"18",X"69",X"02",
		X"29",X"06",X"85",X"E6",X"A9",X"00",X"9D",X"01",X"10",X"A5",X"E7",X"18",X"69",X"01",X"29",X"0F",
		X"85",X"E7",X"A6",X"E8",X"E8",X"8A",X"29",X"0F",X"AA",X"8E",X"04",X"14",X"86",X"E8",X"AD",X"01",
		X"0C",X"4A",X"4A",X"26",X"EB",X"A5",X"EB",X"29",X"03",X"C9",X"02",X"D0",X"16",X"E6",X"E9",X"A5",
		X"E9",X"A0",X"01",X"18",X"69",X"01",X"29",X"0F",X"99",X"04",X"14",X"99",X"0C",X"14",X"C8",X"C0",
		X"04",X"90",X"F0",X"AD",X"01",X"0C",X"4A",X"4A",X"4A",X"26",X"EC",X"A5",X"EC",X"29",X"03",X"49",
		X"02",X"D0",X"07",X"A2",X"0F",X"F6",X"34",X"CA",X"10",X"FB",X"A9",X"05",X"85",X"92",X"A9",X"38",
		X"85",X"91",X"AD",X"00",X"08",X"29",X"0C",X"4A",X"4A",X"69",X"01",X"85",X"8B",X"A2",X"05",X"A9",
		X"1F",X"24",X"8B",X"10",X"02",X"A9",X"00",X"20",X"85",X"38",X"C6",X"8B",X"CA",X"D0",X"F0",X"A9",
		X"37",X"85",X"91",X"A9",X"21",X"20",X"85",X"38",X"A9",X"21",X"20",X"85",X"38",X"A9",X"21",X"20",
		X"85",X"38",X"A9",X"36",X"85",X"91",X"A9",X"00",X"A8",X"91",X"91",X"A0",X"40",X"91",X"91",X"AD",
		X"01",X"08",X"4A",X"4A",X"4A",X"4A",X"4A",X"F0",X"1B",X"AA",X"C9",X"06",X"B0",X"16",X"BD",X"D8",
		X"3F",X"20",X"85",X"38",X"A9",X"00",X"20",X"85",X"38",X"A9",X"21",X"E0",X"03",X"D0",X"02",X"A9",
		X"22",X"20",X"85",X"38",X"A9",X"3F",X"85",X"94",X"A9",X"EE",X"2C",X"00",X"08",X"50",X"02",X"A9",
		X"F2",X"85",X"93",X"A9",X"35",X"85",X"91",X"20",X"74",X"38",X"AD",X"01",X"0C",X"85",X"DF",X"AD",
		X"00",X"08",X"85",X"DD",X"AD",X"01",X"08",X"85",X"DE",X"AD",X"00",X"0C",X"29",X"8F",X"85",X"E0",
		X"AD",X"02",X"0C",X"29",X"8F",X"85",X"E1",X"AD",X"03",X"0C",X"85",X"E2",X"AD",X"0A",X"10",X"48",
		X"25",X"E3",X"85",X"E3",X"68",X"05",X"E4",X"85",X"E4",X"A2",X"00",X"AD",X"01",X"0C",X"38",X"2A",
		X"B0",X"01",X"E8",X"0A",X"D0",X"FA",X"8A",X"A4",X"E6",X"0A",X"0A",X"0A",X"99",X"00",X"10",X"8A",
		X"09",X"A0",X"99",X"01",X"10",X"A6",X"E7",X"A0",X"00",X"A5",X"B9",X"84",X"B9",X"18",X"75",X"54",
		X"95",X"54",X"B5",X"64",X"38",X"E5",X"BB",X"84",X"BB",X"95",X"64",X"A0",X"D0",X"A2",X"05",X"9A",
		X"A2",X"07",X"8A",X"BA",X"36",X"DD",X"AA",X"A9",X"21",X"B0",X"02",X"A9",X"20",X"C8",X"99",X"00",
		X"04",X"CA",X"10",X"EE",X"98",X"38",X"E9",X"28",X"A8",X"BA",X"CA",X"10",X"E2",X"A9",X"04",X"85",
		X"92",X"A9",X"3A",X"85",X"91",X"A5",X"E4",X"49",X"FF",X"05",X"E3",X"05",X"E5",X"F0",X"02",X"A9",
		X"25",X"20",X"85",X"38",X"20",X"07",X"3B",X"20",X"4F",X"3A",X"8C",X"B5",X"01",X"F0",X"16",X"48",
		X"A9",X"3B",X"85",X"91",X"A9",X"24",X"20",X"85",X"38",X"A9",X"00",X"20",X"85",X"38",X"68",X"20",
		X"9E",X"38",X"4C",X"D6",X"3F",X"A9",X"04",X"85",X"92",X"A9",X"E9",X"85",X"91",X"38",X"AD",X"8D",
		X"01",X"20",X"9E",X"38",X"AD",X"8C",X"01",X"20",X"9E",X"38",X"AD",X"8B",X"01",X"18",X"20",X"9E",
		X"38",X"A9",X"DE",X"85",X"93",X"A9",X"3F",X"85",X"94",X"20",X"74",X"38",X"A9",X"05",X"85",X"92",
		X"A9",X"08",X"85",X"91",X"A5",X"8D",X"4A",X"4A",X"4A",X"4A",X"F8",X"18",X"69",X"00",X"D8",X"38",
		X"20",X"9E",X"38",X"A9",X"2E",X"20",X"85",X"38",X"A5",X"8D",X"29",X"0F",X"F8",X"18",X"69",X"00",
		X"85",X"8E",X"65",X"8E",X"85",X"8E",X"65",X"8E",X"D8",X"C9",X"60",X"90",X"02",X"A9",X"59",X"18",
		X"20",X"9E",X"38",X"A9",X"E4",X"85",X"93",X"A9",X"3F",X"85",X"94",X"20",X"74",X"38",X"A5",X"EA",
		X"05",X"EB",X"05",X"EC",X"D0",X"10",X"AD",X"B5",X"01",X"49",X"FF",X"8D",X"B5",X"01",X"A9",X"3D",
		X"85",X"F9",X"A9",X"00",X"85",X"FA",X"4C",X"9E",X"3D",X"22",X"24",X"24",X"25",X"23",X"20",X"50",
		X"4C",X"41",X"59",X"D3",X"20",X"47",X"41",X"4D",X"45",X"20",X"54",X"49",X"4D",X"C5",X"48",X"41",
		X"52",X"C4",X"45",X"41",X"53",X"D9",X"4C",X"F6",X"3F",X"13",X"F6",X"3F",X"4B",X"3B",X"C0",X"38");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
