library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity obj1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of obj1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"11",X"11",X"22",X"22",X"22",X"44",X"44",X"8E",X"01",X"11",X"22",X"22",X"22",X"44",X"44",
		X"E8",X"10",X"19",X"2A",X"26",X"26",X"46",X"46",X"EE",X"11",X"91",X"A2",X"62",X"62",X"64",X"64",
		X"44",X"44",X"44",X"88",X"88",X"88",X"88",X"88",X"44",X"44",X"44",X"88",X"88",X"88",X"88",X"88",
		X"46",X"46",X"46",X"89",X"89",X"89",X"89",X"89",X"64",X"64",X"64",X"98",X"98",X"98",X"98",X"98",
		X"88",X"00",X"99",X"AA",X"66",X"66",X"66",X"66",X"8E",X"01",X"11",X"22",X"22",X"22",X"44",X"44",
		X"E8",X"10",X"08",X"08",X"04",X"04",X"02",X"02",X"00",X"00",X"80",X"80",X"40",X"40",X"20",X"20",
		X"66",X"66",X"66",X"99",X"99",X"99",X"99",X"99",X"44",X"44",X"44",X"88",X"88",X"88",X"88",X"88",
		X"02",X"02",X"02",X"01",X"01",X"01",X"01",X"01",X"20",X"20",X"20",X"10",X"10",X"10",X"10",X"10",
		X"88",X"88",X"88",X"88",X"88",X"44",X"44",X"44",X"88",X"88",X"88",X"88",X"88",X"44",X"44",X"44",
		X"89",X"89",X"89",X"89",X"89",X"46",X"46",X"46",X"98",X"98",X"98",X"98",X"98",X"64",X"64",X"64",
		X"44",X"44",X"22",X"22",X"22",X"11",X"11",X"00",X"44",X"44",X"22",X"22",X"22",X"11",X"01",X"8E",
		X"46",X"46",X"26",X"26",X"2A",X"19",X"10",X"E8",X"64",X"64",X"62",X"62",X"A2",X"91",X"11",X"EE",
		X"99",X"99",X"99",X"99",X"99",X"66",X"66",X"66",X"88",X"88",X"88",X"88",X"88",X"44",X"44",X"44",
		X"01",X"01",X"01",X"01",X"01",X"02",X"02",X"02",X"10",X"10",X"10",X"10",X"10",X"20",X"20",X"20",
		X"66",X"66",X"66",X"66",X"AA",X"99",X"00",X"88",X"44",X"44",X"22",X"22",X"22",X"11",X"01",X"8E",
		X"02",X"02",X"04",X"04",X"08",X"08",X"10",X"E8",X"20",X"20",X"40",X"40",X"80",X"80",X"00",X"00",
		X"00",X"11",X"11",X"22",X"22",X"22",X"44",X"44",X"8E",X"01",X"11",X"22",X"22",X"22",X"44",X"44",
		X"E8",X"10",X"19",X"2A",X"26",X"26",X"46",X"46",X"EE",X"11",X"91",X"A2",X"62",X"62",X"64",X"64",
		X"44",X"44",X"44",X"88",X"88",X"88",X"88",X"88",X"44",X"44",X"44",X"88",X"88",X"88",X"88",X"88",
		X"46",X"46",X"46",X"89",X"89",X"89",X"89",X"89",X"64",X"64",X"64",X"98",X"98",X"98",X"98",X"98",
		X"88",X"00",X"99",X"AA",X"66",X"66",X"66",X"66",X"8E",X"01",X"11",X"22",X"22",X"22",X"44",X"44",
		X"E8",X"10",X"08",X"08",X"15",X"15",X"02",X"02",X"00",X"00",X"86",X"81",X"40",X"40",X"20",X"31",
		X"66",X"66",X"66",X"99",X"99",X"99",X"99",X"99",X"44",X"44",X"44",X"88",X"88",X"88",X"88",X"88",
		X"02",X"02",X"02",X"23",X"23",X"23",X"23",X"23",X"31",X"31",X"31",X"32",X"32",X"32",X"32",X"32",
		X"88",X"88",X"88",X"88",X"88",X"44",X"44",X"44",X"88",X"88",X"88",X"88",X"88",X"44",X"44",X"44",
		X"89",X"89",X"89",X"89",X"89",X"46",X"46",X"46",X"98",X"98",X"98",X"98",X"98",X"64",X"64",X"64",
		X"44",X"44",X"22",X"22",X"22",X"11",X"11",X"00",X"44",X"44",X"22",X"22",X"22",X"11",X"01",X"8E",
		X"46",X"46",X"26",X"26",X"2A",X"19",X"10",X"E8",X"64",X"64",X"62",X"62",X"A2",X"91",X"11",X"EE",
		X"99",X"99",X"99",X"99",X"99",X"66",X"66",X"66",X"88",X"88",X"88",X"88",X"88",X"44",X"44",X"44",
		X"23",X"23",X"23",X"23",X"23",X"02",X"02",X"02",X"32",X"32",X"32",X"32",X"32",X"31",X"31",X"31",
		X"66",X"66",X"66",X"66",X"AA",X"99",X"00",X"88",X"44",X"44",X"22",X"22",X"22",X"11",X"01",X"8E",
		X"02",X"02",X"15",X"15",X"08",X"08",X"10",X"E8",X"31",X"20",X"40",X"40",X"81",X"86",X"00",X"00",
		X"00",X"00",X"00",X"00",X"68",X"18",X"9C",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E6",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"04",X"15",X"13",X"13",X"13",X"13",X"13",X"91",X"91",X"40",X"40",X"40",X"40",X"40",X"40",
		X"00",X"00",X"88",X"88",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"11",X"22",X"22",X"22",X"44",X"44",X"8E",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"08",X"04",X"04",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"44",X"44",X"88",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"02",X"02",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"13",X"13",X"13",X"13",X"13",X"15",X"04",X"04",X"40",X"40",X"40",X"40",X"40",X"40",X"91",X"91",
		X"88",X"88",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"9C",X"18",X"68",X"00",X"00",X"00",X"00",X"E6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"88",X"88",X"88",X"88",X"44",X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"01",X"01",X"02",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"44",X"22",X"22",X"22",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"8E",
		X"02",X"02",X"04",X"04",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"00",X"06",X"89",X"89",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"22",X"22",X"22",X"22",X"22",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"04",X"04",X"04",X"04",X"04",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"89",X"89",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"08",X"08",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"22",X"22",X"22",X"22",X"11",X"11",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"04",X"04",X"04",X"04",X"08",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"89",X"89",X"06",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"11",X"11",X"11",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"89",X"89",
		X"08",X"08",X"08",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"88",X"01",X"89",X"05",X"00",X"44",X"23",X"23",X"1D",X"1F",X"16",X"1C",X"10",
		X"00",X"08",X"0F",X"B4",X"D2",X"F8",X"F8",X"50",X"01",X"16",X"78",X"E0",X"E0",X"C0",X"40",X"40",
		X"33",X"05",X"89",X"01",X"88",X"00",X"00",X"00",X"EF",X"2F",X"16",X"1F",X"1D",X"23",X"23",X"46",
		X"AF",X"F8",X"F8",X"D2",X"B4",X"0F",X"08",X"00",X"BF",X"AE",X"C0",X"E0",X"E0",X"78",X"16",X"01",
		X"00",X"00",X"11",X"00",X"01",X"8B",X"02",X"8B",X"00",X"00",X"0F",X"FC",X"7A",X"3D",X"3D",X"58",
		X"03",X"3C",X"1E",X"78",X"D2",X"E0",X"D0",X"63",X"00",X"80",X"C0",X"E0",X"A0",X"D0",X"37",X"BE",
		X"04",X"33",X"23",X"05",X"44",X"00",X"22",X"00",X"23",X"EF",X"1E",X"0B",X"0F",X"17",X"11",X"11",
		X"AF",X"E9",X"D2",X"F8",X"CB",X"C3",X"0C",X"08",X"BC",X"F0",X"F0",X"3C",X"87",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"21",X"03",X"02",X"00",X"01",X"12",X"16",X"DE",X"F5",X"79",X"3C",
		X"2C",X"F0",X"96",X"3C",X"E0",X"E0",X"A1",X"36",X"00",X"00",X"80",X"00",X"A2",X"A6",X"AE",X"F0",
		X"8B",X"12",X"46",X"11",X"01",X"11",X"00",X"00",X"09",X"77",X"CF",X"0F",X"0D",X"07",X"00",X"88",
		X"F8",X"7C",X"D2",X"D6",X"CF",X"00",X"00",X"00",X"96",X"3C",X"E1",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"01",X"03",X"16",X"FE",X"F9",X"2C",
		X"06",X"3C",X"2C",X"58",X"D1",X"93",X"B6",X"BC",X"00",X"00",X"44",X"CC",X"6C",X"E9",X"87",X"0E",
		X"02",X"8B",X"01",X"46",X"00",X"00",X"00",X"00",X"0D",X"3B",X"67",X"CF",X"8E",X"0B",X"88",X"22",
		X"FC",X"6B",X"6B",X"6E",X"0C",X"08",X"00",X"00",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"11",X"11",X"34",X"69",X"4B",X"5A",X"F0",X"3C",X"FA",X"D3",
		X"80",X"F7",X"86",X"F4",X"84",X"F8",X"38",X"70",X"00",X"00",X"00",X"40",X"E0",X"B4",X"2D",X"69",
		X"03",X"02",X"03",X"89",X"23",X"00",X"00",X"00",X"2F",X"2E",X"6E",X"4D",X"89",X"07",X"44",X"11",
		X"F6",X"E1",X"7B",X"3D",X"06",X"2C",X"00",X"00",X"C2",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"12",X"03",X"03",X"34",X"3D",X"F0",X"F0",X"69",X"79",X"C3",X"B5",X"E1",X"FB",
		X"E4",X"DC",X"2C",X"B8",X"58",X"A9",X"F0",X"70",X"00",X"80",X"C0",X"E0",X"E1",X"A5",X"86",X"0E",
		X"EF",X"03",X"03",X"01",X"00",X"44",X"11",X"00",X"4B",X"3F",X"26",X"2E",X"2E",X"66",X"09",X"00",
		X"F6",X"71",X"96",X"0F",X"0B",X"0E",X"00",X"AA",X"84",X"84",X"8C",X"8C",X"44",X"00",X"00",X"00",
		X"68",X"34",X"34",X"12",X"12",X"12",X"03",X"16",X"11",X"B3",X"C3",X"F3",X"E1",X"79",X"E1",X"F7",
		X"00",X"10",X"F0",X"30",X"F0",X"61",X"F0",X"76",X"61",X"C2",X"C2",X"84",X"84",X"84",X"0C",X"86",
		X"17",X"6E",X"89",X"01",X"00",X"00",X"00",X"11",X"CB",X"3F",X"1F",X"1B",X"1F",X"11",X"02",X"44",
		X"F1",X"03",X"07",X"05",X"07",X"00",X"04",X"22",X"8E",X"66",X"19",X"08",X"00",X"00",X"00",X"88",
		X"00",X"10",X"30",X"70",X"78",X"5A",X"16",X"07",X"72",X"E6",X"9E",X"A6",X"D6",X"7B",X"E1",X"F1",
		X"F0",X"F0",X"E1",X"61",X"B4",X"52",X"F0",X"75",X"08",X"08",X"08",X"84",X"0C",X"0C",X"C2",X"CB",
		X"12",X"12",X"13",X"13",X"22",X"00",X"00",X"00",X"E7",X"F9",X"96",X"0F",X"0D",X"07",X"00",X"55",
		X"69",X"8B",X"8A",X"8B",X"8B",X"CC",X"09",X"00",X"7F",X"0C",X"0C",X"08",X"00",X"22",X"88",X"00",
		X"00",X"11",X"11",X"31",X"70",X"D2",X"4B",X"69",X"10",X"98",X"F8",X"1C",X"FC",X"86",X"F2",X"D3",
		X"C2",X"69",X"2D",X"A5",X"F0",X"C3",X"F5",X"70",X"00",X"00",X"00",X"00",X"08",X"08",X"88",X"88",
		X"34",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"E7",X"78",X"ED",X"CB",X"06",X"43",X"00",X"00",
		X"0B",X"8B",X"CD",X"4D",X"6E",X"0E",X"22",X"88",X"0C",X"04",X"0C",X"19",X"4C",X"00",X"00",X"00",
		X"00",X"00",X"22",X"33",X"63",X"79",X"1E",X"07",X"06",X"C3",X"43",X"A1",X"B8",X"9C",X"D6",X"D3",
		X"00",X"00",X"08",X"0C",X"86",X"F7",X"F9",X"43",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0C",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"F3",X"6D",X"6D",X"67",X"03",X"01",X"00",X"00",
		X"0B",X"CD",X"6E",X"3F",X"17",X"0D",X"11",X"44",X"04",X"1D",X"08",X"26",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"00",X"54",X"56",X"57",X"F0",X"43",X"F0",X"96",X"C3",X"70",X"70",X"58",X"C6",
		X"00",X"08",X"84",X"86",X"B7",X"FA",X"E9",X"C3",X"00",X"00",X"00",X"00",X"00",X"48",X"0C",X"04",
		X"96",X"C3",X"78",X"07",X"00",X"00",X"00",X"00",X"F1",X"E3",X"B4",X"B6",X"3F",X"00",X"00",X"00",
		X"09",X"EE",X"3F",X"0F",X"0B",X"0E",X"00",X"11",X"1D",X"04",X"26",X"88",X"08",X"88",X"00",X"00",
		X"00",X"10",X"30",X"70",X"50",X"B0",X"CE",X"D7",X"0C",X"C3",X"87",X"E1",X"B4",X"70",X"B0",X"6C",
		X"00",X"00",X"0F",X"F3",X"E5",X"CB",X"CB",X"A1",X"00",X"00",X"88",X"00",X"08",X"1D",X"04",X"1D",
		X"D3",X"F0",X"F0",X"C3",X"1E",X"01",X"00",X"00",X"5F",X"79",X"B4",X"F1",X"3D",X"3C",X"03",X"01",
		X"4C",X"7F",X"87",X"0D",X"0F",X"8E",X"88",X"88",X"02",X"CC",X"4C",X"0A",X"22",X"00",X"44",X"00",
		X"00",X"00",X"00",X"88",X"01",X"89",X"05",X"00",X"00",X"47",X"23",X"1D",X"1F",X"16",X"1C",X"10",
		X"00",X"01",X"1E",X"87",X"F0",X"CB",X"F8",X"50",X"07",X"78",X"F0",X"68",X"E0",X"C0",X"40",X"40",
		X"33",X"05",X"89",X"01",X"88",X"00",X"00",X"00",X"EF",X"2F",X"16",X"1F",X"1D",X"23",X"47",X"00",
		X"AF",X"F8",X"CB",X"F0",X"87",X"1E",X"01",X"00",X"BF",X"AE",X"C0",X"E0",X"68",X"F0",X"78",X"07",
		X"00",X"00",X"00",X"88",X"01",X"89",X"05",X"00",X"00",X"00",X"00",X"3F",X"1F",X"16",X"1C",X"10",
		X"00",X"01",X"1E",X"3C",X"4B",X"F8",X"F8",X"50",X"00",X"0E",X"F0",X"F0",X"2C",X"E0",X"40",X"40",
		X"33",X"05",X"89",X"01",X"88",X"00",X"00",X"00",X"EF",X"2F",X"16",X"1F",X"3F",X"00",X"00",X"00",
		X"AF",X"F8",X"F8",X"C3",X"3C",X"1E",X"01",X"00",X"BF",X"AE",X"E0",X"2C",X"F0",X"F0",X"0E",X"00",
		X"00",X"00",X"00",X"88",X"01",X"89",X"05",X"00",X"00",X"00",X"00",X"0D",X"3F",X"16",X"1C",X"10",
		X"00",X"00",X"00",X"0F",X"0F",X"F8",X"F8",X"50",X"00",X"00",X"00",X"0F",X"96",X"E0",X"40",X"40",
		X"33",X"05",X"89",X"01",X"88",X"00",X"00",X"00",X"EF",X"2F",X"16",X"3F",X"0D",X"00",X"00",X"00",
		X"AF",X"F8",X"F8",X"0F",X"0F",X"00",X"00",X"00",X"BF",X"AE",X"E0",X"96",X"0F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"88",X"01",X"89",X"05",X"00",X"00",X"00",X"00",X"0C",X"0F",X"37",X"1C",X"10",
		X"00",X"00",X"00",X"00",X"0F",X"0F",X"8F",X"50",X"00",X"00",X"00",X"00",X"0F",X"1E",X"2C",X"40",
		X"33",X"05",X"89",X"01",X"88",X"00",X"00",X"00",X"EF",X"2F",X"37",X"0F",X"0C",X"00",X"00",X"00",
		X"AF",X"8F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"BF",X"2C",X"1E",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"40",X"44",X"23",X"2A",X"00",X"00",X"00",X"00",X"06",X"0B",X"0E",X"00",
		X"00",X"00",X"10",X"31",X"71",X"73",X"64",X"A0",X"00",X"00",X"C0",X"EC",X"EE",X"EE",X"C4",X"80",
		X"75",X"39",X"21",X"44",X"40",X"02",X"00",X"00",X"FF",X"FF",X"1F",X"0B",X"17",X"33",X"00",X"00",
		X"5F",X"5F",X"EC",X"FB",X"F9",X"31",X"10",X"00",X"6E",X"4C",X"C4",X"EE",X"EE",X"EC",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"41",X"00",X"00",X"00",X"00",X"00",X"9F",X"0B",X"0E",
		X"00",X"30",X"70",X"73",X"F3",X"D1",X"20",X"93",X"00",X"80",X"C0",X"C8",X"CC",X"44",X"A2",X"4C",
		X"3B",X"75",X"10",X"14",X"20",X"02",X"00",X"00",X"DD",X"FF",X"FF",X"0F",X"05",X"00",X"00",X"00",
		X"5F",X"7E",X"F3",X"FC",X"88",X"00",X"00",X"00",X"4C",X"FF",X"FE",X"EC",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",
		X"00",X"00",X"70",X"F0",X"F3",X"F2",X"40",X"31",X"00",X"00",X"80",X"88",X"88",X"00",X"6E",X"AE",
		X"00",X"13",X"11",X"11",X"12",X"02",X"00",X"00",X"03",X"8F",X"8D",X"9F",X"F7",X"F3",X"A3",X"08",
		X"E7",X"BF",X"DF",X"DE",X"EE",X"8C",X"08",X"00",X"BF",X"7E",X"EC",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"32",X"36",X"68",X"80",
		X"00",X"60",X"F0",X"F3",X"E6",X"F6",X"C0",X"13",X"00",X"00",X"00",X"00",X"00",X"EE",X"7E",X"AC",
		X"10",X"00",X"00",X"01",X"11",X"00",X"01",X"00",X"33",X"67",X"47",X"46",X"47",X"FB",X"20",X"04",
		X"E7",X"3E",X"4E",X"6E",X"CE",X"8C",X"00",X"00",X"C8",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"12",X"76",X"06",X"0E",X"0C",
		X"00",X"F0",X"E2",X"E6",X"F6",X"E0",X"D4",X"11",X"00",X"00",X"00",X"00",X"6E",X"AE",X"CC",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"3B",X"33",X"33",X"33",X"36",X"30",X"02",
		X"EF",X"9F",X"0F",X"0D",X"1F",X"F7",X"00",X"08",X"88",X"08",X"C8",X"8C",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"07",X"0F",X"1E",X"1E",X"DE",X"3E",X"2C",
		X"00",X"20",X"60",X"E0",X"F0",X"E0",X"D0",X"73",X"00",X"00",X"00",X"CC",X"0C",X"CC",X"08",X"00",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"2C",X"59",X"59",X"11",X"00",X"00",X"00",X"00",
		X"CF",X"EF",X"8F",X"8E",X"8F",X"57",X"E8",X"0A",X"08",X"4C",X"4C",X"4C",X"CC",X"88",X"00",X"00",
		X"00",X"00",X"01",X"21",X"21",X"21",X"33",X"21",X"00",X"62",X"F7",X"F7",X"F7",X"F3",X"F8",X"2C",
		X"00",X"22",X"77",X"87",X"77",X"86",X"44",X"CB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"21",X"21",X"01",X"00",X"00",X"00",X"00",X"00",X"3D",X"3D",X"1D",X"19",X"00",X"11",X"11",X"00",
		X"FF",X"CF",X"CF",X"CF",X"EF",X"C0",X"23",X"08",X"08",X"0C",X"04",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"03",X"03",X"11",X"00",X"30",X"30",X"78",X"78",X"78",X"3F",X"EC",
		X"44",X"22",X"C3",X"B3",X"C2",X"B3",X"C7",X"67",X"00",X"00",X"00",X"00",X"00",X"00",X"4C",X"2E",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"2C",X"2C",X"2C",X"06",X"00",X"00",X"00",X"00",
		X"CF",X"EF",X"77",X"33",X"10",X"11",X"01",X"00",X"26",X"2E",X"AE",X"CC",X"C8",X"42",X"00",X"00",
		X"00",X"00",X"00",X"30",X"30",X"34",X"34",X"12",X"00",X"11",X"11",X"ED",X"D5",X"E5",X"C0",X"E0",
		X"00",X"88",X"4C",X"CC",X"0C",X"CF",X"BF",X"C7",X"00",X"00",X"00",X"00",X"00",X"00",X"8C",X"CE",
		X"13",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"C8",X"2C",X"2C",X"1E",X"16",X"00",X"00",X"00",
		X"8E",X"8F",X"CF",X"FF",X"77",X"00",X"00",X"00",X"6E",X"6E",X"6D",X"C8",X"CE",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"33",X"70",X"70",X"30",X"00",X"66",X"67",X"57",X"73",X"AB",X"A0",X"E0",
		X"00",X"00",X"00",X"00",X"08",X"DF",X"BF",X"87",X"00",X"00",X"00",X"00",X"00",X"08",X"8C",X"CC",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C4",X"D9",X"15",X"13",X"01",X"00",X"00",X"00",
		X"8E",X"8F",X"CF",X"FF",X"CD",X"00",X"00",X"00",X"4C",X"6D",X"C8",X"CA",X"04",X"00",X"00",X"00",
		X"00",X"00",X"11",X"00",X"00",X"33",X"77",X"71",X"F0",X"77",X"BF",X"AF",X"E7",X"93",X"A8",X"CC",
		X"00",X"80",X"80",X"C8",X"AF",X"BF",X"F7",X"17",X"00",X"00",X"00",X"00",X"08",X"0C",X"EF",X"EC",
		X"70",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"C6",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0D",X"0F",X"17",X"00",X"00",X"00",X"00",X"00",X"EC",X"6D",X"44",X"82",X"08",X"00",X"00",X"00",
		X"00",X"10",X"31",X"11",X"33",X"67",X"10",X"10",X"00",X"C0",X"EC",X"EC",X"7E",X"DF",X"BF",X"41",
		X"00",X"00",X"00",X"00",X"CF",X"6F",X"7F",X"FF",X"00",X"00",X"00",X"00",X"00",X"09",X"AC",X"C8",
		X"76",X"FF",X"F7",X"70",X"00",X"00",X"00",X"00",X"54",X"CC",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"17",X"0D",X"0F",X"33",X"00",X"00",X"00",X"00",X"EB",X"4C",X"CE",X"40",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"40",X"44",X"23",X"2A",X"00",X"00",X"00",X"00",X"06",X"0B",X"0E",X"00",
		X"00",X"00",X"00",X"00",X"32",X"77",X"64",X"A0",X"00",X"00",X"00",X"00",X"C0",X"E8",X"C4",X"80",
		X"75",X"39",X"21",X"40",X"40",X"02",X"00",X"00",X"FF",X"FF",X"1F",X"0B",X"17",X"33",X"00",X"00",
		X"5F",X"5F",X"EC",X"FF",X"BA",X"00",X"00",X"00",X"6E",X"4C",X"C4",X"E8",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"40",X"44",X"23",X"2A",X"00",X"00",X"00",X"00",X"06",X"0B",X"0E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"73",X"70",X"B0",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"C4",
		X"75",X"39",X"21",X"40",X"40",X"02",X"00",X"00",X"FF",X"FF",X"1F",X"0B",X"17",X"33",X"00",X"00",
		X"4E",X"5E",X"F8",X"FB",X"88",X"00",X"00",X"00",X"2A",X"C4",X"EE",X"EE",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"FE",
		X"00",X"11",X"30",X"00",X"F0",X"00",X"10",X"F0",X"00",X"FF",X"F0",X"00",X"86",X"00",X"F0",X"00",
		X"0F",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"E1",X"11",X"11",X"01",X"00",X"00",X"00",
		X"02",X"0F",X"EF",X"FF",X"0F",X"33",X"03",X"10",X"0C",X"00",X"0F",X"CC",X"0E",X"EE",X"0F",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"67",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"8F",X"67",X"00",X"00",X"00",X"00",X"00",X"00",X"2D",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"06",X"0F",X"0B",X"0E",X"00",
		X"00",X"62",X"F1",X"F1",X"F3",X"E3",X"E6",X"A0",X"00",X"00",X"0C",X"0C",X"08",X"00",X"00",X"A0",
		X"11",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"FF",X"1F",X"0B",X"0F",X"06",X"00",X"00",X"00",
		X"5F",X"6E",X"E3",X"F3",X"F1",X"F1",X"62",X"00",X"4E",X"00",X"00",X"08",X"0C",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"16",X"0F",X"0B",
		X"00",X"00",X"C4",X"E3",X"E3",X"E3",X"E2",X"F7",X"00",X"00",X"00",X"08",X"08",X"20",X"C6",X"08",
		X"40",X"11",X"00",X"00",X"20",X"00",X"00",X"00",X"9F",X"FF",X"EF",X"07",X"05",X"03",X"00",X"00",
		X"5F",X"DF",X"78",X"78",X"38",X"00",X"00",X"00",X"00",X"0E",X"CE",X"C4",X"88",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"06",X"0F",
		X"00",X"00",X"CF",X"E3",X"E3",X"E3",X"F2",X"B3",X"00",X"00",X"08",X"08",X"20",X"46",X"C4",X"0C",
		X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"0B",X"1F",X"BB",X"FF",X"46",X"81",X"00",X"00",
		X"B7",X"DE",X"FC",X"1C",X"0C",X"08",X"00",X"00",X"8E",X"8C",X"80",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"76",
		X"00",X"00",X"02",X"86",X"C6",X"F6",X"D5",X"5B",X"00",X"00",X"00",X"40",X"8C",X"08",X"0C",X"08",
		X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"8F",X"8F",X"8D",X"FF",X"45",X"80",X"00",X"00",
		X"F6",X"BC",X"CC",X"8C",X"08",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",
		X"00",X"00",X"12",X"9F",X"E5",X"F7",X"C2",X"A2",X"00",X"00",X"08",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"67",X"47",X"67",X"33",X"80",X"00",X"00",
		X"84",X"08",X"0C",X"04",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",
		X"00",X"42",X"26",X"0C",X"6C",X"E8",X"E2",X"84",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"23",X"23",X"33",X"11",X"00",X"20",X"00",
		X"C8",X"0C",X"28",X"0C",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"10",X"00",X"10",X"00",X"30",
		X"00",X"08",X"8A",X"0E",X"8E",X"3E",X"7C",X"68",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"33",X"11",X"00",X"00",X"00",X"00",
		X"CE",X"0F",X"0D",X"8E",X"CC",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"12",X"01",X"03",X"01",X"11",X"10",X"30",
		X"00",X"00",X"00",X"88",X"80",X"C0",X"C0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"00",X"00",X"00",X"00",X"00",
		X"8F",X"0E",X"8F",X"EE",X"00",X"00",X"20",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"08",X"C4",X"46",X"7D",X"79",X"70",X"74",
		X"00",X"00",X"00",X"00",X"00",X"08",X"C8",X"A6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"31",X"33",X"33",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0D",X"9F",X"EE",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"00",X"00",X"03",X"13",X"11",X"00",X"00",X"0A",X"9E",X"72",X"09",X"FF",X"E1",
		X"00",X"00",X"00",X"00",X"80",X"8C",X"AF",X"F7",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"D1",X"11",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"0D",X"0F",X"9F",X"00",X"10",X"00",X"00",X"88",X"88",X"88",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"31",X"13",X"10",X"03",X"17",X"00",X"00",X"3E",X"36",X"3B",X"DF",X"40",X"FE",
		X"00",X"00",X"00",X"80",X"80",X"0B",X"6E",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",
		X"32",X"30",X"10",X"00",X"00",X"00",X"00",X"00",X"E0",X"C1",X"81",X"00",X"00",X"00",X"00",X"00",
		X"1D",X"1B",X"1F",X"1F",X"00",X"00",X"00",X"00",X"A8",X"88",X"00",X"00",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"00",X"62",X"05",X"10",X"00",X"00",X"74",X"7C",X"7E",X"33",X"AF",X"63",
		X"00",X"00",X"00",X"80",X"87",X"86",X"CF",X"FF",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"A8",
		X"00",X"01",X"03",X"01",X"00",X"00",X"00",X"00",X"76",X"7C",X"FC",X"F8",X"F8",X"64",X"00",X"00",
		X"33",X"17",X"0D",X"0F",X"06",X"00",X"00",X"00",X"88",X"88",X"00",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"06",X"0F",X"0B",X"0E",X"00",
		X"00",X"00",X"E3",X"F1",X"F1",X"F1",X"E7",X"A0",X"00",X"00",X"00",X"08",X"08",X"08",X"00",X"A0",
		X"11",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"FF",X"1F",X"0B",X"0F",X"06",X"00",X"00",X"00",
		X"5F",X"6F",X"F1",X"F1",X"F1",X"E3",X"00",X"00",X"4E",X"00",X"08",X"08",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"06",X"0F",X"0B",X"0E",X"00",
		X"00",X"00",X"00",X"00",X"30",X"F0",X"F0",X"A0",X"00",X"00",X"00",X"00",X"C4",X"C6",X"8C",X"A0",
		X"11",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"FF",X"1F",X"0B",X"0F",X"06",X"00",X"00",X"00",
		X"5F",X"78",X"F0",X"30",X"00",X"00",X"00",X"00",X"4E",X"8C",X"C6",X"C4",X"00",X"00",X"00",X"00",
		X"00",X"9F",X"6F",X"9F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"9F",X"66",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"9F",X"6F",X"9F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"9F",X"66",
		X"00",X"66",X"9F",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9F",X"6F",X"9F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"66",X"9F",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9F",X"6F",X"9F",
		X"00",X"00",X"00",X"00",X"04",X"44",X"32",X"10",X"00",X"00",X"00",X"06",X"0F",X"0B",X"1E",X"F0",
		X"00",X"33",X"44",X"44",X"44",X"80",X"90",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"01",X"23",X"44",X"04",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0B",X"0F",X"06",X"00",X"00",X"00",
		X"0F",X"4D",X"C4",X"44",X"77",X"77",X"33",X"00",X"0C",X"80",X"00",X"00",X"00",X"88",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"76",X"00",X"00",X"00",X"00",X"00",X"06",X"0F",X"1A",
		X"00",X"00",X"44",X"CC",X"88",X"DC",X"D4",X"C5",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"0C",
		X"10",X"01",X"11",X"22",X"02",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"07",X"05",X"12",X"00",X"00",
		X"0F",X"0E",X"6A",X"3B",X"91",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"88",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"11",X"11",X"00",X"B4",X"0F",
		X"00",X"00",X"88",X"88",X"00",X"98",X"F4",X"E1",X"00",X"00",X"00",X"00",X"80",X"84",X"08",X"08",
		X"10",X"14",X"33",X"00",X"00",X"11",X"00",X"00",X"1A",X"2D",X"4B",X"0F",X"8A",X"01",X"08",X"00",
		X"86",X"7B",X"59",X"0C",X"48",X"08",X"00",X"00",X"00",X"44",X"88",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"70",X"F0",
		X"00",X"00",X"00",X"98",X"A9",X"B8",X"A9",X"D7",X"00",X"00",X"00",X"00",X"08",X"08",X"00",X"00",
		X"10",X"10",X"10",X"02",X"11",X"00",X"00",X"00",X"C3",X"87",X"85",X"0F",X"8D",X"08",X"00",X"00",
		X"97",X"68",X"0C",X"0C",X"48",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"70",
		X"00",X"00",X"00",X"61",X"A9",X"89",X"8A",X"D3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"E1",X"C3",X"C3",X"47",X"08",X"00",X"00",
		X"C2",X"48",X"0C",X"40",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"20",X"70",
		X"00",X"00",X"84",X"C2",X"42",X"46",X"8C",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"F0",X"F0",X"70",X"70",X"11",X"02",X"00",
		X"C0",X"2C",X"0A",X"2C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"30",X"30",X"30",X"30",
		X"00",X"00",X"08",X"84",X"95",X"91",X"A2",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"70",X"70",X"70",X"30",X"00",X"00",X"00",
		X"C2",X"87",X"85",X"0E",X"84",X"88",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"70",X"41",X"60",X"20",X"30",
		X"00",X"00",X"00",X"08",X"08",X"08",X"8C",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"70",X"70",X"30",X"10",X"00",X"00",X"00",
		X"87",X"85",X"87",X"C2",X"C0",X"44",X"02",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"86",X"81",X"88",X"FF",X"70",
		X"00",X"00",X"00",X"00",X"88",X"08",X"48",X"96",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"70",X"70",X"30",X"10",X"00",X"00",X"00",
		X"0F",X"0D",X"87",X"D2",X"E2",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"00",X"33",X"11",X"00",X"00",X"00",X"0C",X"97",X"90",X"11",X"FE",
		X"00",X"00",X"00",X"00",X"88",X"68",X"4B",X"87",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"30",X"30",X"10",X"00",X"00",X"00",X"00",
		X"0F",X"0D",X"87",X"F0",X"E0",X"01",X"00",X"00",X"08",X"08",X"08",X"8C",X"88",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"30",X"10",X"00",X"00",X"00",X"11",X"11",X"0E",X"C3",X"F0",X"32",
		X"00",X"00",X"00",X"88",X"88",X"83",X"0E",X"87",X"00",X"00",X"00",X"00",X"00",X"80",X"08",X"08",
		X"00",X"22",X"11",X"00",X"00",X"00",X"00",X"00",X"74",X"CD",X"98",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"1A",X"1E",X"F0",X"00",X"00",X"00",X"00",X"2B",X"4C",X"00",X"88",X"88",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"30",X"00",X"44",X"22",X"33",X"11",X"1D",X"0F",X"C3",
		X"00",X"00",X"00",X"00",X"07",X"86",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"08",X"01",X"2A",
		X"10",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"F2",X"76",X"CD",X"DC",X"88",X"00",X"00",X"00",
		X"87",X"0F",X"1A",X"0E",X"C0",X"00",X"00",X"00",X"4C",X"80",X"88",X"44",X"44",X"04",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"44",X"32",X"10",X"00",X"00",X"00",X"06",X"0F",X"0B",X"1E",X"F0",
		X"00",X"00",X"00",X"33",X"44",X"C4",X"90",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"01",X"23",X"44",X"04",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0B",X"0F",X"06",X"00",X"00",X"00",
		X"0F",X"5C",X"C4",X"77",X"33",X"00",X"00",X"00",X"0C",X"80",X"00",X"44",X"88",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"44",X"32",X"10",X"00",X"00",X"00",X"06",X"0F",X"0B",X"1E",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"F7",X"C4",X"F0",X"00",X"00",X"00",X"00",X"00",X"88",X"44",X"C0",
		X"01",X"23",X"44",X"04",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0B",X"0F",X"06",X"00",X"00",X"00",
		X"1E",X"4C",X"F7",X"00",X"00",X"00",X"00",X"00",X"48",X"44",X"88",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"73",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"73",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"BC",X"9E",X"8F",
		X"00",X"00",X"00",X"00",X"EE",X"F1",X"F3",X"F7",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"8F",X"9E",X"BC",X"77",X"00",X"00",X"00",X"00",
		X"F7",X"F3",X"F1",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"22",X"10",X"10",X"00",X"00",X"00",X"06",X"0F",X"0B",X"1E",X"F0",
		X"00",X"33",X"44",X"44",X"44",X"80",X"90",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"01",X"01",X"22",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0B",X"0F",X"06",X"00",X"00",X"00",
		X"AF",X"CD",X"C4",X"44",X"77",X"77",X"33",X"00",X"8C",X"80",X"00",X"00",X"00",X"88",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"30",X"00",X"00",X"00",X"00",X"0C",X"1E",X"16",X"3C",
		X"00",X"00",X"22",X"44",X"88",X"98",X"F0",X"A7",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C8",
		X"32",X"01",X"01",X"11",X"00",X"00",X"00",X"00",X"C3",X"0F",X"0F",X"0D",X"03",X"00",X"00",X"00",
		X"CD",X"CC",X"7B",X"19",X"00",X"00",X"00",X"00",X"80",X"00",X"88",X"CC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"10",X"00",X"00",X"00",X"00",X"0C",X"1E",X"16",X"3C",
		X"00",X"00",X"00",X"33",X"CC",X"B8",X"C3",X"AE",X"00",X"00",X"00",X"00",X"80",X"80",X"CC",X"44",
		X"23",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"C3",X"0F",X"0F",X"0D",X"8B",X"00",X"00",X"00",
		X"FF",X"7B",X"08",X"08",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"11",X"22",X"22",X"22",X"3D",X"3C",X"34",
		X"00",X"00",X"00",X"30",X"71",X"43",X"A7",X"8C",X"00",X"00",X"00",X"00",X"80",X"88",X"22",X"22",
		X"01",X"00",X"23",X"00",X"00",X"00",X"00",X"00",X"2D",X"4B",X"87",X"87",X"05",X"44",X"00",X"00",
		X"7F",X"3D",X"0E",X"06",X"0C",X"00",X"00",X"00",X"EE",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"11",X"11",X"00",X"00",X"01",X"03",X"00",X"88",X"00",X"00",X"88",X"44",X"78",X"3C",
		X"00",X"00",X"00",X"F0",X"F2",X"96",X"C4",X"BF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"01",X"00",X"11",X"00",X"00",X"00",X"00",X"34",X"2D",X"4B",X"87",X"03",X"01",X"11",X"00",
		X"7D",X"0E",X"0F",X"0B",X"0E",X"00",X"00",X"00",X"FF",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"DC",X"CD",X"44",X"73",X"3F",
		X"00",X"00",X"C0",X"E8",X"68",X"C8",X"48",X"F3",X"00",X"00",X"00",X"00",X"00",X"44",X"88",X"00",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"07",X"1E",X"1E",X"9E",X"11",X"00",X"00",
		X"E0",X"86",X"0F",X"0B",X"86",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"23",X"55",X"45",X"55",X"67",X"73",
		X"00",X"00",X"C4",X"A2",X"A2",X"A2",X"E6",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0B",X"0F",X"03",X"44",X"00",X"00",
		X"C3",X"87",X"85",X"87",X"C0",X"22",X"00",X"00",X"00",X"08",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"22",X"11",X"00",X"00",X"00",X"30",X"71",X"61",X"31",X"21",X"FC",
		X"00",X"00",X"11",X"B3",X"3B",X"22",X"EC",X"CF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"16",X"0F",X"0D",X"16",X"10",X"00",X"00",
		X"0F",X"0E",X"87",X"87",X"97",X"88",X"00",X"00",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F4",X"96",X"32",X"DF",
		X"00",X"11",X"00",X"00",X"11",X"22",X"E1",X"C3",X"00",X"00",X"88",X"88",X"00",X"00",X"08",X"0C",
		X"FF",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"EB",X"07",X"0F",X"0D",X"07",X"00",X"00",X"00",
		X"C2",X"4B",X"2D",X"1E",X"0C",X"08",X"88",X"00",X"0C",X"08",X"00",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"33",X"00",X"C4",X"8E",X"A6",X"C3",X"31",
		X"00",X"88",X"CC",X"CC",X"CC",X"CB",X"8F",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",
		X"44",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"74",X"F8",X"07",X"06",X"03",X"00",X"00",X"00",
		X"0F",X"87",X"4B",X"3C",X"0A",X"22",X"00",X"00",X"08",X"00",X"4C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"10",X"33",X"22",X"00",X"00",X"00",X"CC",X"33",X"D1",X"3C",X"57",
		X"00",X"00",X"00",X"00",X"03",X"87",X"86",X"C3",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"80",
		X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"ED",X"01",X"01",X"00",X"00",X"00",X"00",
		X"3C",X"0F",X"0F",X"0B",X"1D",X"00",X"00",X"00",X"4C",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"31",X"00",X"00",X"44",X"22",X"11",X"91",X"F0",X"5E",
		X"00",X"00",X"00",X"00",X"03",X"87",X"86",X"C3",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"C0",
		X"10",X"00",X"11",X"33",X"00",X"00",X"00",X"00",X"3B",X"33",X"ED",X"89",X"00",X"00",X"00",X"00",
		X"3C",X"0F",X"0F",X"0B",X"0C",X"00",X"00",X"00",X"C4",X"08",X"08",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"22",X"10",X"10",X"00",X"00",X"00",X"06",X"0F",X"0B",X"1E",X"F0",
		X"00",X"00",X"00",X"33",X"44",X"C4",X"90",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"01",X"01",X"22",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0B",X"0F",X"06",X"00",X"00",X"00",
		X"AF",X"DC",X"C4",X"77",X"33",X"00",X"00",X"00",X"8C",X"80",X"00",X"44",X"88",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"22",X"10",X"10",X"00",X"00",X"00",X"06",X"0F",X"0B",X"1E",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"F7",X"C4",X"F0",X"00",X"00",X"00",X"00",X"00",X"88",X"44",X"C0",
		X"01",X"01",X"22",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0B",X"0F",X"06",X"00",X"00",X"00",
		X"BE",X"4C",X"F7",X"00",X"00",X"00",X"00",X"00",X"C8",X"44",X"88",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"23",
		X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"4C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"23",X"11",X"00",X"00",X"00",X"00",X"00",X"00",
		X"4C",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"32",X"74",X"F8",X"F0",
		X"00",X"00",X"00",X"88",X"CC",X"EE",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",
		X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"8F",X"47",X"23",X"11",X"00",X"00",X"00",
		X"F0",X"F1",X"E2",X"C4",X"88",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"07",X"03",X"01",X"06",X"46",X"68",X"00",X"00",X"0C",X"1E",X"1E",X"2D",X"78",X"20",
		X"00",X"03",X"0F",X"0F",X"0E",X"0C",X"80",X"00",X"00",X"0C",X"0E",X"08",X"00",X"00",X"00",X"00",
		X"77",X"79",X"46",X"06",X"01",X"03",X"07",X"0F",X"FF",X"EC",X"78",X"2D",X"1E",X"1E",X"0C",X"00",
		X"FF",X"77",X"80",X"48",X"0E",X"0F",X"0F",X"03",X"DA",X"00",X"00",X"00",X"00",X"08",X"0E",X"0C",
		X"00",X"00",X"00",X"07",X"0F",X"0F",X"01",X"06",X"00",X"00",X"01",X"0B",X"2D",X"2D",X"3C",X"2C",
		X"43",X"0F",X"1E",X"0C",X"0C",X"08",X"80",X"77",X"08",X"80",X"00",X"00",X"00",X"00",X"52",X"88",
		X"46",X"7B",X"31",X"27",X"03",X"00",X"01",X"01",X"33",X"FC",X"DE",X"16",X"07",X"0F",X"0F",X"0E",
		X"FF",X"00",X"0C",X"0F",X"87",X"87",X"03",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0C",X"00",
		X"00",X"00",X"00",X"00",X"07",X"0F",X"0F",X"09",X"10",X"03",X"07",X"07",X"4B",X"4B",X"2D",X"68",
		X"0C",X"0C",X"08",X"08",X"00",X"00",X"33",X"FF",X"00",X"00",X"00",X"00",X"42",X"84",X"88",X"00",
		X"06",X"56",X"31",X"36",X"03",X"11",X"00",X"00",X"19",X"FE",X"FE",X"83",X"0B",X"0F",X"03",X"07",
		X"AA",X"0E",X"87",X"4B",X"2D",X"0C",X"0C",X"08",X"00",X"00",X"0F",X"0F",X"0E",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"0F",X"07",X"07",X"0E",X"0E",X"0E",X"87",X"87",X"68",
		X"08",X"00",X"00",X"00",X"10",X"BB",X"FF",X"66",X"00",X"00",X"40",X"08",X"00",X"00",X"00",X"01",
		X"0F",X"0C",X"16",X"32",X"13",X"01",X"00",X"00",X"39",X"32",X"FF",X"EF",X"C1",X"8D",X"07",X"03",
		X"06",X"87",X"87",X"69",X"0E",X"0E",X"0C",X"08",X"03",X"0F",X"0F",X"0C",X"00",X"00",X"00",X"00",
		X"00",X"01",X"01",X"01",X"01",X"10",X"07",X"0F",X"0C",X"0C",X"0C",X"0C",X"0C",X"1F",X"86",X"59",
		X"00",X"01",X"12",X"64",X"CC",X"CC",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0F",
		X"0F",X"0F",X"0A",X"03",X"23",X"01",X"00",X"00",X"79",X"6E",X"66",X"E7",X"E4",X"CB",X"2B",X"00",
		X"07",X"C3",X"B4",X"0F",X"0F",X"07",X"07",X"0E",X"0F",X"0E",X"0C",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"07",X"07",X"07",X"07",X"03",X"30",X"00",X"00",X"00",X"00",X"19",X"19",X"1D",X"1D",
		X"40",X"04",X"40",X"88",X"88",X"88",X"89",X"43",X"00",X"00",X"00",X"21",X"43",X"07",X"1E",X"0E",
		X"07",X"0F",X"0F",X"0E",X"0D",X"01",X"00",X"00",X"F1",X"3D",X"6E",X"66",X"6E",X"EB",X"39",X"02",
		X"43",X"F0",X"0F",X"0F",X"07",X"0B",X"0B",X"03",X"0C",X"08",X"00",X"08",X"08",X"08",X"08",X"00",
		X"00",X"02",X"06",X"07",X"07",X"07",X"03",X"03",X"00",X"00",X"00",X"00",X"11",X"19",X"59",X"2C",
		X"80",X"08",X"80",X"88",X"88",X"88",X"89",X"A9",X"00",X"02",X"03",X"07",X"07",X"0F",X"0E",X"0E",
		X"10",X"01",X"03",X"03",X"07",X"07",X"06",X"04",X"A4",X"78",X"3D",X"1F",X"19",X"16",X"36",X"01",
		X"A9",X"F8",X"A9",X"8B",X"88",X"CB",X"EB",X"04",X"C0",X"0C",X"0E",X"0E",X"0F",X"07",X"03",X"01",
		X"00",X"00",X"00",X"0C",X"0E",X"0E",X"0F",X"07",X"20",X"02",X"20",X"11",X"11",X"11",X"19",X"2C",
		X"00",X"00",X"00",X"00",X"89",X"89",X"8B",X"8B",X"0C",X"0C",X"0E",X"0E",X"0E",X"0E",X"0C",X"C0",
		X"03",X"01",X"00",X"01",X"01",X"01",X"01",X"00",X"2C",X"F0",X"0F",X"0F",X"0E",X"0D",X"0D",X"0C",
		X"F8",X"CB",X"67",X"66",X"67",X"7D",X"C9",X"04",X"0E",X"0F",X"0F",X"07",X"0B",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0F",X"00",X"08",X"84",X"40",X"EE",X"66",X"77",X"33",
		X"03",X"03",X"03",X"03",X"03",X"07",X"16",X"A9",X"00",X"08",X"08",X"08",X"08",X"80",X"0E",X"0F",
		X"0F",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"0E",X"3C",X"D2",X"0F",X"0F",X"0E",X"0E",X"07",
		X"E9",X"CD",X"CC",X"7E",X"72",X"3D",X"4D",X"00",X"0F",X"0F",X"05",X"0C",X"4C",X"08",X"00",X"00",
		X"00",X"00",X"20",X"01",X"00",X"00",X"00",X"08",X"01",X"00",X"00",X"00",X"80",X"DD",X"FF",X"66",
		X"0E",X"0E",X"07",X"07",X"07",X"1E",X"1E",X"61",X"00",X"00",X"00",X"00",X"00",X"0C",X"0E",X"0F",
		X"0C",X"0F",X"0F",X"03",X"00",X"00",X"00",X"00",X"06",X"1E",X"1E",X"69",X"07",X"07",X"03",X"01",
		X"C9",X"C4",X"FF",X"7F",X"3C",X"1B",X"0A",X"0C",X"0F",X"09",X"86",X"C4",X"8C",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"24",X"12",X"11",X"00",X"03",X"03",X"01",X"01",X"00",X"00",X"CC",X"FF",
		X"80",X"0C",X"0E",X"0E",X"2D",X"2D",X"4B",X"61",X"00",X"00",X"00",X"00",X"0E",X"0F",X"0F",X"09",
		X"00",X"00",X"0F",X"0F",X"07",X"00",X"00",X"00",X"55",X"06",X"1E",X"2D",X"4B",X"03",X"03",X"01",
		X"89",X"F7",X"F7",X"1C",X"0D",X"0F",X"0C",X"0E",X"06",X"A6",X"C8",X"C6",X"0C",X"88",X"00",X"00",
		X"01",X"10",X"00",X"00",X"00",X"00",X"A4",X"11",X"2C",X"0F",X"87",X"03",X"03",X"01",X"10",X"EE",
		X"00",X"00",X"08",X"0D",X"4B",X"4B",X"C3",X"43",X"00",X"00",X"00",X"0E",X"0F",X"0F",X"08",X"06",
		X"00",X"00",X"00",X"00",X"0F",X"0F",X"03",X"00",X"FF",X"00",X"03",X"0F",X"1E",X"1E",X"0C",X"00",
		X"CC",X"F3",X"B7",X"86",X"0E",X"0F",X"0F",X"07",X"26",X"ED",X"C8",X"4E",X"0C",X"00",X"08",X"08",
		X"00",X"00",X"0F",X"07",X"01",X"06",X"46",X"68",X"00",X"00",X"0C",X"1E",X"1E",X"2D",X"78",X"20",
		X"00",X"03",X"87",X"0F",X"0E",X"0C",X"80",X"00",X"00",X"0C",X"0E",X"08",X"00",X"00",X"00",X"00",
		X"77",X"79",X"46",X"06",X"01",X"07",X"0F",X"00",X"FF",X"EC",X"F8",X"2D",X"1E",X"1E",X"0C",X"00",
		X"FF",X"77",X"80",X"48",X"0E",X"0F",X"0F",X"03",X"DA",X"00",X"00",X"00",X"00",X"08",X"0E",X"0C",
		X"00",X"00",X"00",X"0F",X"03",X"06",X"46",X"68",X"00",X"00",X"00",X"0C",X"1E",X"2D",X"78",X"20",
		X"00",X"00",X"07",X"0F",X"0F",X"0C",X"80",X"00",X"00",X"00",X"0C",X"0E",X"00",X"00",X"00",X"00",
		X"77",X"79",X"46",X"06",X"03",X"0F",X"00",X"00",X"FF",X"EC",X"F8",X"2D",X"1E",X"0C",X"00",X"00",
		X"FF",X"77",X"80",X"48",X"0F",X"0F",X"07",X"00",X"DA",X"00",X"00",X"00",X"00",X"0E",X"0C",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"06",X"46",X"68",X"00",X"00",X"00",X"00",X"1E",X"2D",X"70",X"20",
		X"00",X"00",X"00",X"0F",X"0F",X"0C",X"80",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",
		X"77",X"79",X"46",X"06",X"0F",X"00",X"00",X"00",X"FF",X"EC",X"70",X"2D",X"1E",X"00",X"00",X"00",
		X"FF",X"77",X"80",X"48",X"87",X"0F",X"00",X"00",X"DA",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"46",X"68",X"00",X"00",X"00",X"00",X"00",X"0C",X"0F",X"02",
		X"00",X"00",X"00",X"00",X"00",X"87",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"C0",X"00",
		X"77",X"79",X"46",X"0F",X"00",X"00",X"00",X"00",X"FF",X"CE",X"0F",X"0C",X"00",X"00",X"00",X"00",
		X"FF",X"77",X"3C",X"0F",X"00",X"00",X"00",X"00",X"DA",X"00",X"C0",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"24",X"12",X"01",X"00",X"22",X"22",X"11",X"00",X"00",X"C0",X"78",X"16",X"10",X"70",X"F0",
		X"00",X"00",X"10",X"E0",X"C0",X"91",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",
		X"00",X"11",X"22",X"22",X"00",X"01",X"03",X"06",X"F0",X"B4",X"70",X"10",X"07",X"0F",X"0C",X"00",
		X"22",X"77",X"00",X"91",X"C0",X"2C",X"01",X"00",X"10",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",
		X"00",X"00",X"00",X"78",X"07",X"00",X"00",X"22",X"00",X"00",X"00",X"F0",X"F0",X"1E",X"10",X"70",
		X"00",X"60",X"40",X"91",X"A2",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"10",X"00",
		X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"00",X"F0",X"B4",X"F8",X"30",X"01",X"03",X"07",X"0E",
		X"77",X"00",X"80",X"68",X"0F",X"0E",X"00",X"00",X"00",X"00",X"AA",X"44",X"80",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"30",X"78",X"06",X"00",X"00",X"00",X"10",X"30",X"F0",X"E0",X"68",X"70",
		X"00",X"80",X"22",X"44",X"44",X"00",X"00",X"33",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",
		X"44",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"F0",X"52",X"F8",X"88",X"88",X"01",X"03",
		X"66",X"80",X"C0",X"78",X"0F",X"0E",X"08",X"08",X"00",X"EE",X"00",X"E0",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"70",X"4B",X"0C",X"00",X"20",X"20",X"60",X"E0",X"E0",X"40",X"60",
		X"00",X"88",X"88",X"88",X"00",X"00",X"33",X"66",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"EE",
		X"00",X"22",X"11",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"DA",X"74",X"44",X"22",X"00",X"00",
		X"00",X"B0",X"C3",X"12",X"06",X"06",X"0E",X"0C",X"00",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"70",X"00",X"91",X"A2",X"D1",X"C0",X"C0",X"C0",X"60",
		X"00",X"10",X"00",X"00",X"00",X"00",X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"22",X"CC",X"00",
		X"C3",X"0C",X"00",X"33",X"00",X"00",X"00",X"00",X"70",X"70",X"61",X"98",X"22",X"11",X"11",X"00",
		X"80",X"F0",X"C1",X"83",X"03",X"03",X"03",X"21",X"F0",X"0C",X"08",X"08",X"00",X"80",X"00",X"00",
		X"00",X"00",X"00",X"10",X"00",X"00",X"10",X"10",X"00",X"22",X"44",X"22",X"80",X"C0",X"C0",X"E0",
		X"20",X"00",X"00",X"00",X"00",X"88",X"CC",X"00",X"00",X"00",X"00",X"44",X"44",X"88",X"10",X"E0",
		X"12",X"34",X"24",X"68",X"08",X"00",X"00",X"00",X"B0",X"B0",X"21",X"30",X"CC",X"00",X"00",X"00",
		X"D0",X"C3",X"E1",X"81",X"88",X"44",X"44",X"00",X"C0",X"C0",X"48",X"48",X"48",X"0C",X"0C",X"04",
		X"00",X"00",X"00",X"00",X"02",X"10",X"10",X"01",X"00",X"00",X"88",X"88",X"55",X"11",X"91",X"C0",
		X"80",X"00",X"00",X"00",X"11",X"88",X"00",X"10",X"00",X"00",X"88",X"88",X"20",X"40",X"C0",X"C0",
		X"01",X"01",X"12",X"12",X"12",X"24",X"04",X"00",X"F0",X"B0",X"A1",X"10",X"11",X"66",X"00",X"00",
		X"F0",X"E0",X"E0",X"C0",X"44",X"33",X"00",X"00",X"48",X"48",X"2C",X"24",X"24",X"12",X"10",X"00",
		X"00",X"00",X"00",X"11",X"11",X"04",X"06",X"01",X"20",X"00",X"00",X"00",X"00",X"BB",X"11",X"80",
		X"00",X"22",X"11",X"22",X"00",X"10",X"10",X"30",X"00",X"00",X"40",X"80",X"80",X"C0",X"C0",X"48",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"F0",X"D0",X"D0",X"C0",X"80",X"91",X"80",X"00",
		X"F0",X"F0",X"68",X"E2",X"99",X"00",X"00",X"00",X"2C",X"16",X"12",X"01",X"88",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"22",X"11",X"04",X"00",X"80",X"00",X"00",X"00",X"66",X"BB",X"22",
		X"00",X"54",X"54",X"54",X"01",X"01",X"03",X"61",X"00",X"00",X"00",X"80",X"80",X"C0",X"48",X"3C",
		X"12",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"F0",X"78",X"68",X"48",X"68",X"24",X"04",
		X"F0",X"78",X"F0",X"51",X"44",X"44",X"88",X"00",X"12",X"01",X"00",X"CC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"00",X"00",X"11",X"00",X"77",X"00",X"11",X"11",X"11",X"00",X"88",X"CC",X"44",
		X"00",X"40",X"40",X"24",X"34",X"07",X"02",X"60",X"00",X"00",X"00",X"00",X"00",X"E0",X"3C",X"12",
		X"00",X"16",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"F0",X"48",X"24",X"24",X"34",X"12",
		X"F0",X"F0",X"79",X"E2",X"22",X"44",X"00",X"00",X"00",X"44",X"88",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"00",X"11",X"00",X"00",X"44",X"22",X"22",X"00",X"00",X"88",X"CC",
		X"80",X"80",X"C0",X"78",X"16",X"05",X"60",X"F0",X"00",X"00",X"00",X"40",X"F0",X"0F",X"00",X"00",
		X"55",X"22",X"10",X"07",X"00",X"00",X"00",X"00",X"00",X"10",X"F0",X"68",X"34",X"12",X"01",X"00",
		X"F0",X"A4",X"E0",X"11",X"91",X"91",X"C0",X"48",X"66",X"88",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"11",X"00",X"00",X"80",X"33",X"11",X"02",X"10",X"89",X"45",X"00",X"00",X"00",X"88",
		X"00",X"00",X"F0",X"0F",X"0F",X"60",X"E0",X"F0",X"00",X"00",X"F0",X"0E",X"00",X"00",X"66",X"88",
		X"00",X"55",X"22",X"00",X"01",X"00",X"00",X"00",X"00",X"10",X"70",X"3C",X"03",X"00",X"00",X"00",
		X"B4",X"F0",X"00",X"C0",X"C0",X"78",X"16",X"01",X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"07",X"32",X"22",X"11",X"00",X"00",X"00",X"00",X"2C",X"F0",X"70",X"F0",
		X"00",X"00",X"00",X"00",X"30",X"B4",X"E0",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",
		X"00",X"11",X"22",X"32",X"07",X"00",X"00",X"00",X"F0",X"B4",X"70",X"F0",X"2C",X"00",X"00",X"00",
		X"22",X"77",X"E0",X"96",X"30",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"34",X"03",X"11",X"00",X"00",X"00",X"00",X"00",X"F0",X"1E",X"C3",
		X"00",X"00",X"00",X"00",X"00",X"91",X"96",X"48",X"00",X"00",X"00",X"00",X"00",X"CC",X"08",X"00",
		X"00",X"11",X"03",X"34",X"00",X"00",X"00",X"00",X"F0",X"87",X"1E",X"F0",X"00",X"00",X"00",X"00",
		X"22",X"48",X"96",X"91",X"00",X"00",X"00",X"00",X"10",X"00",X"08",X"CC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"21",X"00",X"00",X"00",X"30",X"16",X"00",X"F0",X"0F",X"FF",X"70",X"70",X"F7",X"E0",
		X"00",X"F0",X"3D",X"FF",X"C0",X"80",X"00",X"00",X"00",X"98",X"10",X"70",X"00",X"00",X"00",X"00",
		X"E9",X"56",X"33",X"00",X"00",X"00",X"21",X"00",X"1F",X"0E",X"7E",X"70",X"77",X"F0",X"0F",X"FF",
		X"0F",X"00",X"00",X"80",X"CC",X"F0",X"3D",X"FF",X"4C",X"00",X"00",X"00",X"00",X"98",X"10",X"70",
		X"00",X"00",X"00",X"10",X"00",X"00",X"10",X"03",X"00",X"00",X"70",X"0F",X"77",X"30",X"F3",X"E0",
		X"00",X"00",X"F0",X"3D",X"FF",X"80",X"00",X"00",X"00",X"00",X"A8",X"20",X"60",X"00",X"00",X"00",
		X"74",X"23",X"11",X"00",X"00",X"10",X"00",X"00",X"1F",X"86",X"BE",X"33",X"70",X"0F",X"77",X"00",
		X"0F",X"00",X"00",X"88",X"F0",X"3D",X"FF",X"00",X"88",X"00",X"00",X"00",X"A8",X"20",X"60",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
