library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity nrx_nprg_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of nrx_nprg_rom is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"C3",X"00",X"38",X"31",X"00",X"84",X"18",X"32",X"C3",X"80",X"25",X"00",X"00",X"00",X"00",X"00",
		X"D6",X"03",X"D0",X"DD",X"36",X"CA",X"64",X"3C",X"C8",X"DD",X"36",X"AA",X"64",X"DD",X"36",X"88",
		X"0F",X"AF",X"C9",X"98",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C3",X"F0",X"01",X"00",X"00",X"00",X"00",X"00",X"18",X"C6",X"ED",X"46",X"FB",X"3E",X"F7",X"D3",
		X"00",X"21",X"00",X"80",X"11",X"01",X"80",X"01",X"00",X"08",X"36",X"00",X"ED",X"B0",X"E5",X"0E",
		X"08",X"36",X"60",X"ED",X"B0",X"0E",X"18",X"36",X"00",X"ED",X"B0",X"EB",X"E1",X"01",X"E0",X"07",
		X"ED",X"B0",X"C3",X"F7",X"04",X"00",X"C3",X"00",X"00",X"32",X"80",X"A0",X"FD",X"26",X"01",X"2A",
		X"69",X"80",X"ED",X"4B",X"50",X"80",X"3A",X"6B",X"80",X"A7",X"28",X"27",X"3A",X"48",X"80",X"CB",
		X"47",X"C2",X"CE",X"00",X"ED",X"5B",X"4C",X"80",X"19",X"22",X"4C",X"80",X"7A",X"94",X"21",X"73",
		X"80",X"CD",X"3E",X"0F",X"81",X"32",X"50",X"80",X"FD",X"7C",X"A7",X"28",X"31",X"2A",X"5A",X"80",
		X"FD",X"26",X"00",X"3A",X"48",X"80",X"CB",X"4F",X"C2",X"CE",X"00",X"ED",X"5B",X"4E",X"80",X"19",
		X"22",X"4E",X"80",X"7A",X"94",X"21",X"75",X"80",X"CD",X"3E",X"0F",X"ED",X"44",X"80",X"32",X"51",
		X"80",X"FD",X"7C",X"A7",X"28",X"08",X"FD",X"26",X"00",X"2A",X"5A",X"80",X"18",X"B6",X"DD",X"21",
		X"68",X"80",X"3A",X"4E",X"82",X"3C",X"47",X"FD",X"2E",X"01",X"CD",X"E0",X"00",X"C3",X"78",X"01",
		X"DD",X"7E",X"00",X"A7",X"28",X"0D",X"DD",X"7E",X"15",X"A7",X"C2",X"85",X"01",X"DD",X"34",X"00",
		X"C3",X"5A",X"01",X"DD",X"66",X"02",X"DD",X"6E",X"01",X"DD",X"7E",X"03",X"DD",X"E5",X"DD",X"23",
		X"4F",X"A7",X"20",X"04",X"DD",X"23",X"DD",X"23",X"DD",X"56",X"04",X"DD",X"5E",X"03",X"19",X"DD",
		X"75",X"03",X"DD",X"74",X"04",X"7C",X"C6",X"18",X"6F",X"3D",X"FA",X"51",X"01",X"D6",X"2F",X"6F",
		X"FA",X"2D",X"01",X"79",X"A1",X"20",X"2D",X"DD",X"35",X"07",X"DD",X"75",X"04",X"7C",X"92",X"CB",
		X"7F",X"28",X"03",X"DD",X"34",X"0A",X"DD",X"86",X"0B",X"DD",X"77",X"0B",X"30",X"03",X"DD",X"34",
		X"0A",X"DD",X"E1",X"FD",X"2D",X"20",X"13",X"DD",X"7E",X"03",X"2F",X"2A",X"5A",X"80",X"C3",X"FC",
		X"00",X"A1",X"20",X"D3",X"DD",X"34",X"07",X"C3",X"2A",X"01",X"DD",X"7E",X"08",X"87",X"87",X"87",
		X"DD",X"56",X"0A",X"CB",X"3A",X"1F",X"CB",X"3A",X"1F",X"CB",X"3A",X"1F",X"DD",X"77",X"11",X"7A",
		X"E6",X"07",X"F6",X"98",X"DD",X"77",X"12",X"C9",X"11",X"20",X"00",X"DD",X"19",X"FD",X"2E",X"00",
		X"05",X"C2",X"DA",X"00",X"C9",X"DD",X"7E",X"0F",X"21",X"3A",X"25",X"BE",X"23",X"20",X"FC",X"DD",
		X"7E",X"00",X"E6",X"03",X"20",X"04",X"7E",X"DD",X"77",X"0F",X"DD",X"35",X"00",X"C2",X"5A",X"01",
		X"DD",X"36",X"15",X"00",X"C5",X"DD",X"46",X"0C",X"DD",X"4E",X"0E",X"C5",X"CD",X"31",X"10",X"C1",
		X"7E",X"D6",X"BD",X"28",X"14",X"FE",X"09",X"30",X"33",X"FE",X"03",X"38",X"06",X"79",X"C6",X"08",
		X"4F",X"18",X"E8",X"78",X"D6",X"08",X"47",X"18",X"E2",X"06",X"03",X"54",X"5D",X"CB",X"DC",X"0E",
		X"03",X"E5",X"D5",X"1A",X"D6",X"BD",X"FE",X"09",X"30",X"05",X"3E",X"81",X"12",X"36",X"15",X"CD",
		X"0F",X"10",X"0D",X"20",X"EE",X"D1",X"E1",X"CD",X"1E",X"10",X"10",X"E3",X"C1",X"C3",X"5A",X"01",
		X"E5",X"D5",X"C5",X"F5",X"DD",X"E5",X"FD",X"E5",X"AF",X"32",X"81",X"A1",X"32",X"80",X"A0",X"CD",
		X"B3",X"16",X"CD",X"3B",X"17",X"3A",X"20",X"80",X"A7",X"28",X"05",X"FE",X"02",X"C2",X"C3",X"03",
		X"3A",X"4D",X"80",X"32",X"30",X"A1",X"3A",X"4F",X"80",X"ED",X"44",X"32",X"40",X"A1",X"DD",X"21",
		X"14",X"88",X"21",X"15",X"80",X"FD",X"21",X"02",X"80",X"06",X"06",X"FD",X"E5",X"FD",X"5E",X"00",
		X"FD",X"56",X"01",X"7A",X"B3",X"28",X"6E",X"D5",X"FD",X"E1",X"D5",X"CD",X"A0",X"04",X"FD",X"7E",
		X"00",X"0F",X"30",X"07",X"DD",X"CB",X"01",X"FE",X"C3",X"4F",X"02",X"DD",X"CB",X"01",X"BE",X"FD",
		X"7E",X"01",X"77",X"FD",X"7E",X"03",X"DD",X"77",X"00",X"FD",X"7E",X"04",X"2B",X"77",X"23",X"FD",
		X"7E",X"05",X"E6",X"7F",X"57",X"DD",X"7E",X"01",X"E6",X"80",X"B2",X"DD",X"77",X"01",X"78",X"FD",
		X"E1",X"FE",X"06",X"28",X"30",X"ED",X"5B",X"52",X"80",X"3A",X"55",X"80",X"0F",X"E6",X"01",X"ED",
		X"44",X"FD",X"86",X"FF",X"92",X"FE",X"0B",X"30",X"2E",X"57",X"3A",X"54",X"80",X"0F",X"E6",X"01",
		X"ED",X"44",X"FD",X"86",X"FD",X"93",X"FE",X"0B",X"30",X"1D",X"FE",X"0A",X"CC",X"C7",X"02",X"7A",
		X"FE",X"0A",X"CC",X"D8",X"02",X"FD",X"E1",X"FD",X"23",X"FD",X"23",X"DD",X"23",X"DD",X"23",X"23",
		X"23",X"05",X"C2",X"2B",X"02",X"18",X"34",X"FD",X"E1",X"AF",X"FD",X"77",X"00",X"FD",X"77",X"01",
		X"2B",X"3E",X"EC",X"77",X"23",X"18",X"E0",X"3A",X"54",X"80",X"A7",X"28",X"04",X"3D",X"C8",X"18",
		X"16",X"FD",X"CB",X"FA",X"7E",X"C0",X"18",X"0F",X"3A",X"55",X"80",X"A7",X"28",X"04",X"3D",X"C8",
		X"18",X"05",X"FD",X"CB",X"FC",X"7E",X"C8",X"F1",X"C3",X"B7",X"02",X"CD",X"69",X"00",X"CD",X"64",
		X"0F",X"CD",X"CC",X"1E",X"DD",X"21",X"68",X"80",X"06",X"09",X"21",X"94",X"82",X"11",X"34",X"80",
		X"3A",X"6F",X"82",X"E6",X"0F",X"20",X"04",X"36",X"0E",X"18",X"06",X"E6",X"07",X"20",X"02",X"36",
		X"08",X"3A",X"A8",X"81",X"A7",X"20",X"39",X"DD",X"7E",X"08",X"87",X"C6",X"E0",X"CB",X"86",X"38",
		X"02",X"CB",X"C6",X"12",X"DD",X"7E",X"0A",X"D6",X"64",X"28",X"07",X"C6",X"64",X"87",X"ED",X"44",
		X"C6",X"9D",X"CB",X"DA",X"12",X"78",X"23",X"CB",X"9A",X"13",X"01",X"20",X"00",X"DD",X"09",X"47",
		X"10",X"CF",X"21",X"94",X"82",X"11",X"04",X"A0",X"01",X"09",X"00",X"ED",X"B0",X"C3",X"6D",X"03",
		X"DD",X"7E",X"08",X"87",X"ED",X"44",X"C6",X"41",X"CB",X"C6",X"12",X"DD",X"7E",X"0A",X"D6",X"64",
		X"28",X"05",X"C6",X"64",X"87",X"C6",X"5F",X"CB",X"DA",X"12",X"C3",X"35",X"03",X"06",X"05",X"3A",
		X"B3",X"82",X"A7",X"20",X"4E",X"DD",X"21",X"68",X"80",X"FD",X"21",X"04",X"80",X"21",X"4C",X"82",
		X"7E",X"35",X"FE",X"32",X"30",X"3D",X"A7",X"20",X"3A",X"77",X"FD",X"66",X"01",X"FD",X"6E",X"00",
		X"7D",X"B4",X"28",X"29",X"7E",X"CB",X"47",X"20",X"24",X"DD",X"7E",X"0C",X"23",X"96",X"30",X"02",
		X"ED",X"44",X"FE",X"0B",X"30",X"17",X"DD",X"7E",X"0E",X"23",X"23",X"96",X"30",X"02",X"ED",X"44",
		X"FE",X"0B",X"30",X"09",X"3E",X"01",X"32",X"81",X"A1",X"FB",X"C3",X"C1",X"18",X"FD",X"23",X"FD",
		X"23",X"10",X"C7",X"3A",X"4B",X"82",X"3C",X"32",X"4B",X"82",X"CD",X"24",X"0F",X"3A",X"6F",X"82",
		X"3C",X"32",X"6F",X"82",X"E6",X"1F",X"CC",X"8E",X"1F",X"FE",X"0E",X"CC",X"9C",X"1F",X"C6",X"08",
		X"E6",X"0F",X"CC",X"D7",X"04",X"3A",X"4D",X"82",X"3C",X"32",X"4D",X"82",X"E6",X"3F",X"CC",X"82",
		X"04",X"E6",X"07",X"CC",X"72",X"04",X"3A",X"69",X"82",X"3C",X"32",X"69",X"82",X"2A",X"9A",X"89",
		X"3A",X"8C",X"82",X"A7",X"20",X"03",X"3A",X"88",X"82",X"3D",X"32",X"8C",X"82",X"20",X"2F",X"34",
		X"7E",X"21",X"8A",X"82",X"36",X"04",X"FE",X"28",X"38",X"17",X"36",X"03",X"28",X"10",X"FE",X"50",
		X"38",X"0F",X"36",X"02",X"28",X"08",X"FE",X"C8",X"38",X"07",X"36",X"01",X"20",X"03",X"CD",X"1F",
		X"1B",X"3A",X"69",X"82",X"47",X"3A",X"6E",X"82",X"B8",X"30",X"03",X"32",X"69",X"82",X"00",X"21",
		X"F4",X"89",X"3A",X"21",X"80",X"A7",X"20",X"03",X"77",X"23",X"77",X"CD",X"80",X"25",X"3A",X"24",
		X"80",X"FE",X"09",X"3E",X"00",X"30",X"01",X"3C",X"32",X"86",X"A1",X"3A",X"00",X"A1",X"E6",X"01",
		X"CA",X"00",X"38",X"3E",X"01",X"32",X"81",X"A1",X"FD",X"E1",X"DD",X"E1",X"F1",X"C1",X"D1",X"E1",
		X"FB",X"C9",X"2A",X"2D",X"80",X"ED",X"5B",X"69",X"80",X"19",X"CB",X"2C",X"CB",X"1D",X"22",X"69",
		X"80",X"C9",X"47",X"3A",X"92",X"82",X"A7",X"78",X"C8",X"2A",X"27",X"80",X"11",X"E0",X"FF",X"19",
		X"7C",X"A7",X"20",X"07",X"3A",X"2B",X"80",X"BD",X"38",X"01",X"6F",X"22",X"27",X"80",X"78",X"C9",
		X"3A",X"A8",X"81",X"A7",X"C8",X"E5",X"FD",X"56",X"00",X"FD",X"5E",X"01",X"21",X"14",X"01",X"A7",
		X"ED",X"52",X"FD",X"7E",X"03",X"ED",X"44",X"D6",X"10",X"57",X"FD",X"7E",X"04",X"EE",X"03",X"FD",
		X"5E",X"05",X"FD",X"21",X"88",X"81",X"FD",X"74",X"00",X"FD",X"75",X"01",X"FD",X"72",X"03",X"FD",
		X"77",X"04",X"FD",X"73",X"05",X"E1",X"C9",X"3A",X"20",X"80",X"06",X"04",X"2A",X"98",X"89",X"FE",
		X"02",X"C0",X"7E",X"FE",X"66",X"3E",X"67",X"28",X"02",X"3E",X"66",X"77",X"23",X"10",X"FC",X"C9",
		X"06",X"04",X"2A",X"98",X"89",X"18",X"EB",X"21",X"2F",X"22",X"11",X"40",X"80",X"0E",X"66",X"CD",
		X"AF",X"1E",X"CD",X"8A",X"1D",X"3A",X"00",X"A1",X"47",X"21",X"AA",X"82",X"E6",X"C0",X"28",X"0E",
		X"34",X"CB",X"7F",X"28",X"09",X"23",X"34",X"CB",X"77",X"20",X"03",X"34",X"2B",X"34",X"78",X"0F",
		X"0F",X"0F",X"E6",X"01",X"C6",X"02",X"3C",X"32",X"0E",X"80",X"21",X"45",X"23",X"3E",X"15",X"11",
		X"C5",X"24",X"22",X"D2",X"82",X"32",X"D8",X"82",X"21",X"60",X"80",X"0E",X"70",X"EB",X"CD",X"AF",
		X"1E",X"3A",X"0E",X"80",X"3D",X"87",X"87",X"87",X"4F",X"78",X"E6",X"06",X"B1",X"21",X"85",X"24",
		X"85",X"6F",X"30",X"01",X"24",X"5E",X"23",X"56",X"ED",X"53",X"B3",X"81",X"11",X"1F",X"00",X"19",
		X"5E",X"23",X"56",X"ED",X"53",X"B9",X"81",X"3A",X"80",X"A0",X"F6",X"FE",X"2F",X"32",X"A9",X"81",
		X"CD",X"B3",X"16",X"3A",X"A9",X"81",X"32",X"83",X"A1",X"32",X"A8",X"81",X"CD",X"8A",X"1D",X"3A",
		X"24",X"80",X"A7",X"C2",X"5A",X"07",X"32",X"21",X"80",X"3C",X"32",X"81",X"A1",X"32",X"20",X"80",
		X"3E",X"F7",X"D3",X"00",X"3E",X"49",X"CD",X"E5",X"20",X"21",X"A0",X"85",X"06",X"07",X"36",X"81",
		X"23",X"10",X"FB",X"21",X"A0",X"85",X"11",X"C0",X"85",X"01",X"60",X"01",X"ED",X"B0",X"21",X"A0",
		X"8D",X"06",X"07",X"36",X"56",X"23",X"10",X"FB",X"21",X"A0",X"8D",X"11",X"C0",X"8D",X"01",X"C0",
		X"00",X"ED",X"B0",X"06",X"07",X"36",X"55",X"23",X"10",X"FB",X"21",X"60",X"8E",X"01",X"60",X"00",
		X"ED",X"B0",X"06",X"07",X"36",X"45",X"23",X"10",X"FB",X"21",X"C0",X"8E",X"01",X"40",X"00",X"ED",
		X"B0",X"21",X"40",X"8C",X"11",X"41",X"8C",X"01",X"7F",X"00",X"36",X"4A",X"ED",X"B0",X"21",X"40",
		X"8F",X"11",X"41",X"8F",X"01",X"BF",X"00",X"36",X"47",X"ED",X"B0",X"FB",X"21",X"C8",X"22",X"11",
		X"88",X"84",X"CD",X"19",X"07",X"11",X"CA",X"84",X"CD",X"19",X"07",X"DD",X"21",X"14",X"80",X"FD",
		X"21",X"14",X"88",X"DD",X"36",X"00",X"F3",X"DD",X"36",X"01",X"F4",X"FD",X"36",X"00",X"44",X"FD",
		X"36",X"01",X"01",X"3A",X"A8",X"81",X"A7",X"CC",X"DC",X"06",X"11",X"27",X"85",X"CD",X"19",X"07",
		X"DD",X"36",X"02",X"F3",X"DD",X"36",X"03",X"F4",X"FD",X"36",X"02",X"56",X"FD",X"36",X"03",X"02",
		X"3A",X"A8",X"81",X"A7",X"CC",X"E9",X"06",X"11",X"67",X"85",X"CD",X"19",X"07",X"DD",X"21",X"A4",
		X"85",X"DD",X"36",X"00",X"87",X"DD",X"36",X"1F",X"88",X"DD",X"36",X"20",X"89",X"11",X"A7",X"85",
		X"CD",X"19",X"07",X"DD",X"36",X"3F",X"8A",X"DD",X"36",X"40",X"87",X"DD",X"36",X"5F",X"88",X"DD",
		X"36",X"60",X"89",X"11",X"E7",X"85",X"CD",X"19",X"07",X"DD",X"21",X"23",X"86",X"DD",X"36",X"00",
		X"8B",X"DD",X"36",X"01",X"87",X"DD",X"36",X"20",X"88",X"DD",X"36",X"21",X"89",X"11",X"27",X"86",
		X"CD",X"19",X"07",X"E5",X"3E",X"94",X"21",X"63",X"86",X"CD",X"2C",X"07",X"E1",X"11",X"87",X"86",
		X"CD",X"19",X"07",X"E5",X"21",X"C3",X"86",X"3E",X"BD",X"CD",X"2C",X"07",X"E1",X"11",X"E7",X"86",
		X"CD",X"19",X"07",X"11",X"6B",X"87",X"CD",X"19",X"07",X"3E",X"01",X"32",X"4B",X"82",X"3A",X"4B",
		X"82",X"E6",X"3F",X"20",X"F9",X"3E",X"01",X"32",X"0F",X"80",X"32",X"B0",X"81",X"21",X"3F",X"E0",
		X"22",X"F2",X"82",X"21",X"AB",X"81",X"36",X"03",X"AF",X"C3",X"5E",X"08",X"DD",X"36",X"00",X"F0",
		X"DD",X"36",X"01",X"1E",X"FD",X"36",X"00",X"AE",X"C9",X"DD",X"36",X"02",X"F0",X"DD",X"36",X"03",
		X"1E",X"FD",X"36",X"02",X"9C",X"C9",X"DD",X"36",X"00",X"F0",X"DD",X"36",X"01",X"58",X"FD",X"36",
		X"00",X"64",X"C9",X"06",X"00",X"FE",X"0A",X"38",X"05",X"04",X"D6",X"0A",X"18",X"F7",X"4F",X"78",
		X"A7",X"28",X"02",X"12",X"13",X"79",X"12",X"13",X"C9",X"76",X"76",X"76",X"7E",X"23",X"FE",X"20",
		X"28",X"05",X"12",X"13",X"C3",X"19",X"07",X"76",X"3D",X"20",X"FC",X"C9",X"0E",X"03",X"11",X"1D",
		X"00",X"06",X"03",X"77",X"3C",X"23",X"10",X"FB",X"19",X"0D",X"20",X"F5",X"C9",X"21",X"4B",X"82",
		X"36",X"88",X"7E",X"A7",X"20",X"FC",X"21",X"14",X"80",X"11",X"02",X"80",X"06",X"0C",X"AF",X"0E",
		X"EC",X"71",X"23",X"12",X"13",X"10",X"FA",X"C3",X"73",X"05",X"31",X"00",X"84",X"3E",X"02",X"32",
		X"21",X"80",X"3D",X"32",X"20",X"80",X"32",X"81",X"A1",X"FB",X"32",X"B0",X"81",X"32",X"B1",X"81",
		X"21",X"0E",X"80",X"7E",X"23",X"77",X"23",X"77",X"3E",X"66",X"CD",X"E5",X"20",X"21",X"93",X"21",
		X"11",X"66",X"85",X"CD",X"3D",X"1E",X"E5",X"2A",X"B3",X"81",X"7E",X"E1",X"FE",X"49",X"28",X"67",
		X"3A",X"0E",X"80",X"FE",X"03",X"28",X"20",X"11",X"E3",X"85",X"CD",X"3D",X"1E",X"2A",X"B3",X"81",
		X"01",X"07",X"00",X"09",X"11",X"F1",X"85",X"0E",X"01",X"CD",X"3F",X"1E",X"2A",X"B3",X"81",X"0E",
		X"04",X"CD",X"3F",X"1E",X"C3",X"F7",X"07",X"11",X"C2",X"85",X"21",X"F9",X"21",X"CD",X"3D",X"1E",
		X"2A",X"B3",X"81",X"01",X"07",X"00",X"09",X"11",X"D1",X"85",X"0E",X"01",X"CD",X"3F",X"1E",X"2A",
		X"B3",X"81",X"0E",X"04",X"CD",X"3F",X"1E",X"11",X"02",X"86",X"21",X"14",X"22",X"CD",X"3D",X"1E",
		X"2A",X"B9",X"81",X"01",X"06",X"00",X"09",X"11",X"10",X"86",X"0E",X"02",X"CD",X"3F",X"1E",X"2A",
		X"B9",X"81",X"0E",X"04",X"CD",X"3F",X"1E",X"21",X"BD",X"21",X"11",X"6A",X"86",X"CD",X"3D",X"1E",
		X"3A",X"AA",X"82",X"A7",X"C4",X"35",X"21",X"11",X"25",X"87",X"21",X"D1",X"21",X"CD",X"29",X"1D",
		X"11",X"65",X"87",X"21",X"E5",X"21",X"CD",X"29",X"1D",X"3A",X"4B",X"82",X"E6",X"1F",X"CC",X"44",
		X"1E",X"E6",X"0F",X"CC",X"4E",X"1E",X"3A",X"00",X"A0",X"E6",X"40",X"28",X"18",X"3A",X"80",X"A0",
		X"E6",X"40",X"20",X"E5",X"3A",X"24",X"80",X"D6",X"02",X"38",X"DE",X"32",X"24",X"80",X"21",X"AB",
		X"81",X"36",X"03",X"18",X"09",X"21",X"24",X"80",X"35",X"21",X"AB",X"81",X"36",X"01",X"AF",X"E5",
		X"21",X"14",X"80",X"11",X"15",X"80",X"01",X"0B",X"00",X"36",X"EC",X"ED",X"B0",X"E1",X"32",X"81",
		X"A1",X"32",X"80",X"A0",X"3E",X"F7",X"D3",X"00",X"FB",X"3E",X"80",X"32",X"F5",X"89",X"CD",X"33",
		X"19",X"CD",X"4E",X"1E",X"21",X"3F",X"22",X"11",X"80",X"80",X"0E",X"66",X"CD",X"AF",X"1E",X"0E",
		X"72",X"21",X"37",X"22",X"CD",X"BA",X"0C",X"CD",X"AF",X"1E",X"3A",X"AB",X"81",X"47",X"0E",X"66",
		X"FE",X"01",X"21",X"5F",X"22",X"28",X"03",X"21",X"47",X"22",X"CD",X"BA",X"0C",X"CD",X"AF",X"1E",
		X"0E",X"72",X"21",X"37",X"22",X"10",X"03",X"21",X"5F",X"22",X"CD",X"BA",X"0C",X"CD",X"AF",X"1E",
		X"21",X"5F",X"22",X"CD",X"AF",X"1E",X"AF",X"32",X"B2",X"81",X"3E",X"01",X"32",X"B7",X"81",X"2A",
		X"8A",X"89",X"34",X"AF",X"2A",X"8C",X"89",X"77",X"32",X"92",X"82",X"CD",X"1F",X"1B",X"CD",X"43",
		X"13",X"CD",X"79",X"13",X"3E",X"03",X"32",X"81",X"A1",X"FB",X"32",X"20",X"80",X"32",X"4B",X"82",
		X"3A",X"4B",X"82",X"E6",X"3F",X"20",X"F9",X"AF",X"32",X"92",X"82",X"32",X"B4",X"82",X"21",X"90",
		X"82",X"77",X"23",X"77",X"2A",X"9C",X"89",X"77",X"2A",X"9A",X"89",X"77",X"2A",X"8E",X"89",X"77",
		X"23",X"36",X"3C",X"21",X"8A",X"82",X"36",X"04",X"CD",X"8A",X"1D",X"CD",X"1F",X"1B",X"21",X"00",
		X"00",X"11",X"00",X"98",X"0E",X"38",X"06",X"20",X"CD",X"B3",X"14",X"12",X"13",X"24",X"10",X"F8",
		X"32",X"80",X"A0",X"60",X"2C",X"0D",X"20",X"EE",X"2A",X"92",X"89",X"06",X"09",X"3E",X"01",X"5E",
		X"23",X"56",X"23",X"12",X"10",X"F9",X"3E",X"04",X"12",X"5E",X"23",X"56",X"3E",X"02",X"12",X"3A",
		X"51",X"82",X"A7",X"28",X"0D",X"47",X"3E",X"03",X"2A",X"96",X"89",X"5E",X"23",X"56",X"23",X"12",
		X"10",X"F9",X"21",X"4F",X"22",X"11",X"20",X"81",X"0E",X"6B",X"CD",X"AF",X"1E",X"11",X"40",X"81",
		X"0E",X"66",X"06",X"02",X"21",X"5F",X"22",X"CD",X"AF",X"1E",X"10",X"F8",X"06",X"0E",X"0E",X"63",
		X"21",X"67",X"22",X"CD",X"AF",X"1E",X"10",X"F8",X"3A",X"B7",X"81",X"A7",X"C4",X"0F",X"0B",X"11",
		X"80",X"83",X"0E",X"66",X"21",X"57",X"22",X"3A",X"83",X"83",X"A7",X"28",X"06",X"3A",X"21",X"80",
		X"A7",X"28",X"1D",X"CD",X"AF",X"1E",X"2A",X"8A",X"89",X"7E",X"3D",X"21",X"83",X"83",X"06",X"00",
		X"FE",X"0A",X"38",X"05",X"04",X"D6",X"0A",X"18",X"F7",X"77",X"78",X"2B",X"A7",X"28",X"01",X"77",
		X"3A",X"A8",X"81",X"32",X"83",X"A1",X"CD",X"6F",X"14",X"CD",X"7C",X"1F",X"AF",X"32",X"D0",X"82",
		X"21",X"14",X"80",X"06",X"0C",X"36",X"EC",X"23",X"10",X"FB",X"2A",X"8A",X"89",X"7E",X"E6",X"03",
		X"C2",X"92",X"0A",X"21",X"F5",X"89",X"36",X"40",X"3E",X"49",X"CD",X"E5",X"20",X"21",X"40",X"8C",
		X"11",X"41",X"8C",X"01",X"DF",X"00",X"36",X"4A",X"ED",X"B0",X"3A",X"A8",X"81",X"32",X"83",X"A1",
		X"21",X"7F",X"22",X"11",X"E4",X"84",X"CD",X"19",X"07",X"11",X"4B",X"85",X"CD",X"19",X"07",X"E5",
		X"2A",X"8A",X"89",X"7E",X"0F",X"0F",X"E6",X"3F",X"CD",X"03",X"07",X"3E",X"01",X"32",X"20",X"80",
		X"3E",X"94",X"21",X"AA",X"85",X"CD",X"2C",X"07",X"21",X"AA",X"8D",X"36",X"55",X"2C",X"36",X"55",
		X"2C",X"36",X"55",X"11",X"1E",X"00",X"19",X"36",X"55",X"2C",X"36",X"55",X"2C",X"36",X"55",X"19",
		X"36",X"55",X"2C",X"36",X"55",X"2C",X"36",X"55",X"E1",X"11",X"CE",X"85",X"CD",X"19",X"07",X"3A",
		X"51",X"82",X"CD",X"03",X"07",X"DD",X"21",X"14",X"80",X"FD",X"21",X"14",X"88",X"DD",X"36",X"00",
		X"F3",X"DD",X"36",X"01",X"BA",X"FD",X"36",X"00",X"8C",X"FD",X"36",X"01",X"02",X"3A",X"A8",X"81",
		X"A7",X"CC",X"F6",X"06",X"11",X"4E",X"86",X"CD",X"19",X"07",X"3A",X"4E",X"82",X"CD",X"03",X"07",
		X"11",X"A4",X"86",X"CD",X"19",X"07",X"11",X"E3",X"86",X"CD",X"19",X"07",X"3E",X"03",X"32",X"20",
		X"80",X"32",X"81",X"A1",X"FB",X"06",X"40",X"76",X"76",X"10",X"FD",X"21",X"F5",X"89",X"CB",X"46",
		X"28",X"FC",X"CD",X"6C",X"0C",X"21",X"0A",X"2D",X"22",X"52",X"80",X"3E",X"03",X"32",X"20",X"80",
		X"32",X"81",X"A1",X"FB",X"AF",X"32",X"40",X"A1",X"32",X"30",X"A1",X"CD",X"E3",X"12",X"21",X"F5",
		X"89",X"CB",X"46",X"28",X"FC",X"06",X"05",X"11",X"20",X"00",X"0E",X"0D",X"2A",X"27",X"80",X"22",
		X"2D",X"80",X"2A",X"25",X"80",X"AF",X"DD",X"19",X"DD",X"36",X"00",X"88",X"DD",X"77",X"03",X"DD",
		X"77",X"04",X"DD",X"77",X"05",X"DD",X"77",X"06",X"DD",X"77",X"07",X"DD",X"77",X"13",X"DD",X"77",
		X"15",X"DD",X"71",X"08",X"0C",X"0C",X"DD",X"36",X"0A",X"34",X"DD",X"36",X"0F",X"F0",X"DD",X"36",
		X"10",X"02",X"DD",X"75",X"01",X"DD",X"74",X"02",X"10",X"CC",X"3A",X"4E",X"82",X"D7",X"00",X"20",
		X"05",X"DD",X"36",X"EA",X"64",X"3C",X"3D",X"20",X"5A",X"DD",X"36",X"0A",X"64",X"18",X"58",X"D5",
		X"AF",X"32",X"B7",X"81",X"11",X"40",X"83",X"06",X"02",X"0E",X"63",X"21",X"5F",X"22",X"CD",X"AF",
		X"1E",X"10",X"F8",X"D1",X"DD",X"21",X"44",X"83",X"2A",X"88",X"89",X"4E",X"0C",X"18",X"17",X"DD",
		X"21",X"44",X"83",X"11",X"40",X"83",X"06",X"02",X"0E",X"63",X"21",X"5F",X"22",X"CD",X"AF",X"1E",
		X"10",X"F8",X"2A",X"88",X"89",X"4E",X"0D",X"C8",X"3E",X"B0",X"DD",X"77",X"00",X"3C",X"DD",X"77",
		X"01",X"3C",X"DD",X"77",X"20",X"3C",X"DD",X"77",X"21",X"DD",X"7D",X"3C",X"3C",X"E6",X"F7",X"DD",
		X"6F",X"18",X"E3",X"DD",X"36",X"08",X"0B",X"AF",X"0E",X"0F",X"06",X"03",X"CD",X"2B",X"21",X"DD",
		X"19",X"DD",X"36",X"00",X"88",X"DD",X"77",X"03",X"DD",X"77",X"04",X"DD",X"77",X"05",X"DD",X"77",
		X"06",X"DD",X"77",X"07",X"DD",X"71",X"08",X"0C",X"0C",X"DD",X"77",X"13",X"DD",X"77",X"15",X"DD",
		X"36",X"0A",X"64",X"DD",X"36",X"0F",X"F2",X"DD",X"36",X"10",X"02",X"DD",X"75",X"01",X"DD",X"74",
		X"02",X"10",X"CC",X"DD",X"36",X"08",X"0D",X"3A",X"4E",X"82",X"D6",X"06",X"38",X"0E",X"47",X"04",
		X"DD",X"21",X"08",X"81",X"DD",X"19",X"DD",X"36",X"0A",X"01",X"10",X"F8",X"21",X"02",X"80",X"06",
		X"0C",X"11",X"14",X"88",X"AF",X"77",X"12",X"23",X"13",X"10",X"FA",X"21",X"73",X"80",X"22",X"02",
		X"80",X"3E",X"03",X"32",X"20",X"80",X"32",X"81",X"A1",X"32",X"4B",X"82",X"3A",X"4B",X"82",X"E6",
		X"3F",X"20",X"F9",X"21",X"95",X"82",X"06",X"08",X"3E",X"0C",X"77",X"23",X"10",X"FC",X"3E",X"08",
		X"06",X"03",X"77",X"23",X"10",X"FC",X"AF",X"32",X"8C",X"82",X"2A",X"9A",X"89",X"7E",X"FE",X"64",
		X"38",X"02",X"36",X"64",X"3A",X"21",X"80",X"32",X"20",X"80",X"3E",X"5A",X"32",X"4C",X"82",X"3E",
		X"01",X"32",X"81",X"A1",X"21",X"F4",X"89",X"36",X"40",X"23",X"36",X"10",X"2A",X"9C",X"89",X"36",
		X"01",X"CD",X"2F",X"0B",X"CD",X"64",X"20",X"CD",X"69",X"00",X"18",X"39",X"31",X"00",X"84",X"3A",
		X"50",X"80",X"C6",X"07",X"FE",X"0F",X"D4",X"BF",X"11",X"3A",X"51",X"80",X"C6",X"07",X"FE",X"0F",
		X"D4",X"07",X"12",X"3A",X"4B",X"82",X"FE",X"04",X"D4",X"DF",X"1D",X"3A",X"22",X"80",X"A7",X"CA",
		X"52",X"10",X"3D",X"CA",X"D6",X"0C",X"3D",X"CA",X"52",X"10",X"3D",X"CA",X"74",X"17",X"3D",X"CA",
		X"52",X"10",X"CD",X"BD",X"15",X"AF",X"32",X"22",X"80",X"C3",X"2C",X"0C",X"DD",X"21",X"68",X"80",
		X"AF",X"32",X"23",X"80",X"21",X"48",X"80",X"06",X"18",X"77",X"23",X"10",X"FC",X"32",X"81",X"A1",
		X"32",X"50",X"82",X"DD",X"77",X"00",X"DD",X"77",X"01",X"DD",X"77",X"02",X"DD",X"77",X"03",X"DD",
		X"77",X"04",X"DD",X"77",X"05",X"DD",X"77",X"06",X"DD",X"77",X"07",X"DD",X"36",X"08",X"0F",X"DD",
		X"36",X"0A",X"32",X"DD",X"77",X"0B",X"DD",X"36",X"0C",X"70",X"DD",X"36",X"0E",X"74",X"DD",X"36",
		X"0F",X"F0",X"DD",X"36",X"10",X"01",X"DD",X"77",X"13",X"C9",X"3A",X"21",X"80",X"A7",X"C0",X"D5",
		X"13",X"1A",X"A7",X"D1",X"C8",X"C5",X"01",X"08",X"00",X"09",X"EB",X"0E",X"20",X"09",X"EB",X"C1",
		X"E3",X"23",X"23",X"23",X"E3",X"C9",X"DD",X"21",X"88",X"80",X"FD",X"21",X"68",X"80",X"3A",X"4E",
		X"82",X"47",X"A7",X"CA",X"43",X"0E",X"DD",X"7E",X"00",X"A7",X"C2",X"3A",X"0E",X"AF",X"32",X"B5",
		X"81",X"DD",X"7E",X"13",X"DD",X"35",X"13",X"A7",X"C2",X"01",X"0E",X"DD",X"77",X"13",X"FD",X"7E",
		X"08",X"DD",X"96",X"08",X"57",X"30",X"02",X"ED",X"44",X"5F",X"DD",X"7E",X"0A",X"FD",X"96",X"0A",
		X"67",X"30",X"02",X"ED",X"44",X"6F",X"7D",X"FE",X"07",X"30",X"33",X"7B",X"FE",X"07",X"30",X"2E",
		X"7D",X"B3",X"CC",X"4A",X"0E",X"D9",X"DD",X"46",X"0C",X"DD",X"4E",X"0E",X"CD",X"31",X"10",X"7E",
		X"D9",X"FE",X"BD",X"38",X"10",X"FE",X"C6",X"30",X"0C",X"DD",X"36",X"00",X"88",X"DD",X"36",X"15",
		X"01",X"DD",X"36",X"13",X"82",X"0E",X"01",X"78",X"E6",X"03",X"28",X"0C",X"18",X"3E",X"78",X"32",
		X"B5",X"81",X"CB",X"47",X"28",X"36",X"0E",X"03",X"FD",X"7E",X"03",X"A7",X"20",X"18",X"FD",X"CB",
		X"02",X"7E",X"28",X"03",X"79",X"18",X"02",X"AF",X"91",X"84",X"67",X"CB",X"7C",X"6C",X"28",X"1C",
		X"7D",X"ED",X"44",X"6F",X"18",X"16",X"FD",X"CB",X"02",X"7E",X"28",X"04",X"AF",X"91",X"18",X"01",
		X"79",X"82",X"57",X"CB",X"7A",X"5A",X"28",X"04",X"7A",X"ED",X"44",X"5F",X"DD",X"7E",X"05",X"C6",
		X"03",X"FE",X"07",X"D2",X"01",X"0E",X"DD",X"7E",X"07",X"C6",X"03",X"FE",X"07",X"D2",X"01",X"0E",
		X"7D",X"BB",X"30",X"05",X"4C",X"3E",X"FF",X"18",X"03",X"4A",X"54",X"AF",X"F5",X"3A",X"B5",X"81",
		X"A7",X"2A",X"25",X"80",X"28",X"03",X"2A",X"29",X"80",X"F1",X"CB",X"7A",X"C4",X"2B",X"21",X"DD",
		X"36",X"14",X"02",X"5F",X"DD",X"BE",X"03",X"20",X"0D",X"DD",X"7E",X"02",X"AC",X"CB",X"7F",X"7B",
		X"20",X"09",X"DD",X"36",X"14",X"00",X"CD",X"63",X"0E",X"30",X"56",X"2F",X"F5",X"79",X"AC",X"CB",
		X"7F",X"C4",X"2B",X"21",X"F1",X"DD",X"36",X"14",X"02",X"DD",X"BE",X"03",X"20",X"0E",X"DD",X"36",
		X"14",X"00",X"5F",X"DD",X"7E",X"02",X"AC",X"CB",X"7F",X"20",X"06",X"7B",X"CD",X"63",X"0E",X"30",
		X"30",X"2A",X"25",X"80",X"3A",X"B5",X"81",X"A7",X"28",X"03",X"2A",X"29",X"80",X"DD",X"7E",X"02",
		X"AC",X"CB",X"7F",X"C4",X"2B",X"21",X"DD",X"7E",X"03",X"CD",X"63",X"0E",X"30",X"13",X"DD",X"36",
		X"14",X"02",X"2F",X"CD",X"63",X"0E",X"30",X"09",X"CD",X"2B",X"21",X"CD",X"63",X"0E",X"30",X"01",
		X"2F",X"DD",X"77",X"03",X"DD",X"74",X"02",X"DD",X"75",X"01",X"11",X"20",X"00",X"DD",X"19",X"05",
		X"C2",X"E6",X"0C",X"21",X"22",X"80",X"34",X"C3",X"2C",X"0C",X"FD",X"7E",X"0C",X"DD",X"96",X"0C",
		X"57",X"30",X"02",X"ED",X"44",X"5F",X"FD",X"7E",X"0E",X"DD",X"96",X"0E",X"67",X"30",X"02",X"ED",
		X"44",X"6F",X"C9",X"C5",X"4F",X"E5",X"EB",X"DD",X"66",X"08",X"DD",X"6E",X"0A",X"06",X"00",X"1E",
		X"00",X"79",X"A7",X"20",X"40",X"DD",X"7E",X"05",X"C6",X"18",X"FE",X"2B",X"30",X"1C",X"FE",X"06",
		X"38",X"15",X"FE",X"1E",X"30",X"04",X"FE",X"13",X"30",X"11",X"3A",X"5B",X"80",X"A7",X"CA",X"0C",
		X"0F",X"3C",X"CA",X"0C",X"0F",X"18",X"04",X"25",X"18",X"01",X"24",X"CB",X"7A",X"20",X"0B",X"DD",
		X"7E",X"07",X"1D",X"A7",X"FA",X"EE",X"0E",X"2D",X"18",X"44",X"DD",X"7E",X"07",X"1C",X"3D",X"F2",
		X"EE",X"0E",X"2C",X"18",X"39",X"DD",X"7E",X"07",X"C6",X"18",X"FE",X"2B",X"30",X"1A",X"FE",X"06",
		X"38",X"13",X"FE",X"1E",X"30",X"04",X"FE",X"13",X"30",X"0F",X"3A",X"5B",X"80",X"A7",X"28",X"3C",
		X"3C",X"28",X"39",X"18",X"04",X"2C",X"18",X"01",X"2D",X"DD",X"7E",X"05",X"CB",X"7A",X"20",X"08",
		X"04",X"A7",X"FA",X"EE",X"0E",X"24",X"18",X"06",X"05",X"3D",X"F2",X"EE",X"0E",X"25",X"EB",X"CD",
		X"E0",X"14",X"08",X"7A",X"80",X"57",X"7B",X"85",X"5F",X"CD",X"E0",X"14",X"38",X"09",X"7A",X"80",
		X"57",X"7B",X"85",X"5F",X"CD",X"E0",X"14",X"08",X"E1",X"79",X"C1",X"C9",X"E1",X"79",X"C1",X"37",
		X"C9",X"2B",X"7D",X"F6",X"E0",X"3C",X"C0",X"21",X"00",X"9F",X"C9",X"23",X"7D",X"E6",X"1F",X"C0",
		X"21",X"00",X"9F",X"C9",X"E5",X"D5",X"F5",X"2A",X"00",X"80",X"29",X"30",X"01",X"2C",X"7D",X"E6",
		X"49",X"20",X"04",X"11",X"80",X"40",X"19",X"22",X"00",X"80",X"F1",X"D1",X"E1",X"C9",X"57",X"1E",
		X"09",X"23",X"CB",X"7F",X"28",X"03",X"2B",X"34",X"23",X"86",X"77",X"30",X"03",X"2B",X"34",X"23",
		X"7D",X"C6",X"20",X"30",X"01",X"24",X"6F",X"7A",X"1D",X"20",X"E7",X"C9",X"E5",X"21",X"F4",X"89",
		X"CB",X"EE",X"E1",X"C9",X"E5",X"D5",X"C5",X"2A",X"9E",X"89",X"7E",X"21",X"90",X"82",X"0F",X"0F",
		X"CB",X"16",X"7E",X"E6",X"0F",X"FE",X"0C",X"23",X"20",X"2C",X"7E",X"A7",X"20",X"28",X"ED",X"5B",
		X"8A",X"89",X"1A",X"E6",X"03",X"28",X"1F",X"3A",X"21",X"80",X"A7",X"28",X"19",X"ED",X"5B",X"8E",
		X"89",X"13",X"1A",X"A7",X"28",X"10",X"06",X"02",X"3D",X"28",X"0B",X"FE",X"0A",X"CC",X"5C",X"0F",
		X"10",X"F6",X"12",X"34",X"34",X"34",X"7E",X"A7",X"28",X"61",X"DD",X"21",X"68",X"80",X"DD",X"7E",
		X"0F",X"06",X"08",X"0E",X"F0",X"FE",X"F0",X"28",X"14",X"0E",X"18",X"FE",X"F2",X"28",X"0E",X"0E",
		X"08",X"06",X"20",X"FE",X"FC",X"28",X"06",X"06",X"F0",X"FE",X"FD",X"20",X"3E",X"DD",X"7E",X"0C",
		X"90",X"47",X"DD",X"7E",X"0E",X"81",X"4F",X"CD",X"31",X"10",X"54",X"5D",X"CB",X"DC",X"CB",X"7E",
		X"28",X"29",X"1A",X"FE",X"81",X"20",X"24",X"CB",X"BE",X"06",X"03",X"3E",X"BD",X"0E",X"03",X"E5",
		X"D5",X"12",X"3C",X"36",X"45",X"CD",X"0F",X"10",X"0D",X"20",X"F6",X"D1",X"E1",X"CD",X"1E",X"10",
		X"10",X"EB",X"21",X"91",X"82",X"35",X"21",X"F4",X"89",X"CB",X"E6",X"C1",X"D1",X"E1",X"C9",X"F5",
		X"7B",X"F6",X"E0",X"3C",X"20",X"04",X"7B",X"D6",X"20",X"5F",X"1C",X"6B",X"F1",X"C9",X"C5",X"F5",
		X"01",X"20",X"00",X"09",X"7C",X"E6",X"03",X"F6",X"8C",X"67",X"E6",X"F7",X"57",X"5D",X"F1",X"C1",
		X"C9",X"3A",X"4D",X"80",X"80",X"C6",X"03",X"0F",X"0F",X"0F",X"E6",X"1F",X"47",X"3A",X"4F",X"80",
		X"ED",X"44",X"91",X"D6",X"08",X"26",X"21",X"17",X"CB",X"14",X"17",X"CB",X"14",X"E6",X"E0",X"B0",
		X"6F",X"C9",X"11",X"00",X"00",X"DD",X"21",X"68",X"80",X"DD",X"7E",X"13",X"DD",X"35",X"13",X"A7",
		X"C2",X"58",X"11",X"DD",X"77",X"13",X"21",X"F4",X"89",X"CB",X"F6",X"2A",X"27",X"80",X"ED",X"4B",
		X"9E",X"89",X"0A",X"47",X"F3",X"22",X"2D",X"80",X"AF",X"32",X"68",X"80",X"32",X"48",X"80",X"2A",
		X"69",X"80",X"3A",X"20",X"80",X"A7",X"CC",X"A2",X"1D",X"CD",X"8A",X"11",X"30",X"79",X"3A",X"6B",
		X"80",X"2A",X"69",X"80",X"CD",X"63",X"0E",X"30",X"2F",X"2F",X"57",X"3A",X"4B",X"80",X"A7",X"3E",
		X"00",X"32",X"4B",X"80",X"7A",X"28",X"0B",X"2A",X"49",X"80",X"CD",X"63",X"0E",X"30",X"19",X"2A",
		X"69",X"80",X"A7",X"CC",X"2B",X"21",X"CD",X"63",X"0E",X"30",X"0D",X"CD",X"2B",X"21",X"CD",X"63",
		X"0E",X"30",X"05",X"A7",X"CC",X"2B",X"21",X"2F",X"32",X"6B",X"80",X"22",X"69",X"80",X"EB",X"2A",
		X"2D",X"80",X"F5",X"7A",X"AC",X"CB",X"7F",X"C4",X"2B",X"21",X"F1",X"22",X"2D",X"80",X"FB",X"21",
		X"80",X"00",X"A7",X"CA",X"2A",X"11",X"CB",X"68",X"CA",X"62",X"11",X"CB",X"60",X"CA",X"6C",X"11",
		X"3A",X"6F",X"80",X"A7",X"CA",X"4B",X"11",X"FE",X"13",X"F2",X"4E",X"11",X"FE",X"EE",X"FA",X"46",
		X"11",X"CB",X"7F",X"20",X"49",X"18",X"3F",X"08",X"38",X"04",X"08",X"C3",X"C8",X"10",X"08",X"C5",
		X"DD",X"46",X"03",X"B8",X"C1",X"CA",X"C8",X"10",X"08",X"3E",X"01",X"32",X"4B",X"80",X"08",X"ED",
		X"5B",X"69",X"80",X"ED",X"53",X"49",X"80",X"C3",X"C8",X"10",X"CB",X"58",X"28",X"48",X"CB",X"50",
		X"28",X"4E",X"3A",X"6D",X"80",X"A7",X"28",X"13",X"FE",X"13",X"F2",X"4E",X"11",X"FE",X"EE",X"FA",
		X"46",X"11",X"CB",X"7F",X"20",X"08",X"21",X"80",X"FF",X"18",X"03",X"21",X"00",X"00",X"22",X"5A",
		X"80",X"3A",X"20",X"80",X"A7",X"CC",X"D9",X"1D",X"3A",X"22",X"80",X"3C",X"32",X"22",X"80",X"C3",
		X"2C",X"0C",X"3A",X"6F",X"80",X"FE",X"03",X"FA",X"4E",X"11",X"18",X"DF",X"3A",X"6F",X"80",X"FE",
		X"FE",X"F2",X"46",X"11",X"18",X"D5",X"3A",X"6D",X"80",X"FE",X"03",X"FA",X"4E",X"11",X"18",X"CB",
		X"3A",X"6D",X"80",X"FE",X"FE",X"F2",X"46",X"11",X"18",X"C1",X"78",X"CB",X"6F",X"28",X"0E",X"CB",
		X"67",X"28",X"17",X"CB",X"5F",X"28",X"20",X"CB",X"57",X"28",X"20",X"37",X"C9",X"3E",X"00",X"CB",
		X"7C",X"CA",X"63",X"0E",X"CD",X"2B",X"21",X"C3",X"63",X"0E",X"3E",X"00",X"CB",X"7C",X"C2",X"63",
		X"0E",X"CD",X"2B",X"21",X"C3",X"63",X"0E",X"3E",X"FF",X"18",X"E4",X"3E",X"FF",X"18",X"ED",X"F3",
		X"CB",X"7F",X"28",X"22",X"3A",X"50",X"80",X"C6",X"08",X"32",X"50",X"80",X"3A",X"54",X"80",X"3C",
		X"32",X"54",X"80",X"FE",X"03",X"C2",X"7E",X"12",X"AF",X"32",X"54",X"80",X"3A",X"52",X"80",X"3C",
		X"32",X"52",X"80",X"C3",X"7E",X"12",X"3A",X"50",X"80",X"D6",X"08",X"32",X"50",X"80",X"3A",X"54",
		X"80",X"3D",X"32",X"54",X"80",X"F2",X"A8",X"12",X"3E",X"02",X"32",X"54",X"80",X"3A",X"52",X"80",
		X"3D",X"32",X"52",X"80",X"C3",X"A8",X"12",X"F3",X"CB",X"7F",X"28",X"22",X"3A",X"51",X"80",X"C6",
		X"08",X"32",X"51",X"80",X"3A",X"55",X"80",X"3C",X"32",X"55",X"80",X"FE",X"03",X"C2",X"4F",X"12",
		X"AF",X"32",X"55",X"80",X"3A",X"53",X"80",X"3C",X"32",X"53",X"80",X"C3",X"4F",X"12",X"3A",X"51",
		X"80",X"D6",X"08",X"32",X"51",X"80",X"3A",X"55",X"80",X"3D",X"32",X"55",X"80",X"F2",X"73",X"12",
		X"3E",X"02",X"32",X"55",X"80",X"3A",X"53",X"80",X"3D",X"32",X"53",X"80",X"C3",X"73",X"12",X"CD",
		X"D9",X"12",X"ED",X"5B",X"54",X"80",X"14",X"7A",X"FE",X"03",X"20",X"03",X"24",X"16",X"00",X"7C",
		X"C6",X"0A",X"32",X"59",X"80",X"2A",X"56",X"80",X"01",X"E0",X"FF",X"09",X"CB",X"D4",X"22",X"56",
		X"80",X"18",X"07",X"CD",X"D9",X"12",X"ED",X"5B",X"54",X"80",X"FB",X"C3",X"14",X"13",X"CD",X"D9",
		X"12",X"ED",X"5B",X"54",X"80",X"1C",X"7B",X"FE",X"03",X"20",X"03",X"1E",X"00",X"2C",X"7D",X"C6",
		X"0A",X"32",X"58",X"80",X"2A",X"56",X"80",X"7D",X"E6",X"1F",X"20",X"06",X"7D",X"F6",X"1F",X"6F",
		X"18",X"01",X"2B",X"22",X"56",X"80",X"18",X"07",X"CD",X"D9",X"12",X"ED",X"5B",X"54",X"80",X"FB",
		X"06",X"20",X"48",X"2A",X"58",X"80",X"CD",X"0C",X"15",X"14",X"05",X"C8",X"E5",X"2A",X"56",X"80",
		X"78",X"06",X"00",X"09",X"47",X"7C",X"E6",X"03",X"F6",X"84",X"67",X"22",X"56",X"80",X"E1",X"7A",
		X"FE",X"03",X"20",X"E2",X"16",X"00",X"24",X"18",X"DD",X"CD",X"85",X"16",X"2A",X"52",X"80",X"22",
		X"58",X"80",X"C9",X"CD",X"D9",X"12",X"ED",X"5B",X"54",X"80",X"06",X"20",X"CD",X"14",X"13",X"32",
		X"80",X"A0",X"2A",X"56",X"80",X"78",X"01",X"20",X"00",X"09",X"47",X"CB",X"D4",X"CB",X"9C",X"22",
		X"56",X"80",X"7A",X"05",X"C8",X"FE",X"03",X"20",X"E3",X"3A",X"59",X"80",X"3C",X"32",X"59",X"80",
		X"16",X"00",X"18",X"D8",X"C5",X"D5",X"06",X"20",X"2A",X"58",X"80",X"CD",X"0C",X"15",X"1C",X"E5",
		X"2A",X"56",X"80",X"23",X"7D",X"E6",X"1F",X"20",X"05",X"2B",X"7D",X"E6",X"E0",X"6F",X"22",X"56",
		X"80",X"E1",X"05",X"28",X"0A",X"7B",X"FE",X"03",X"20",X"E1",X"1E",X"00",X"2C",X"18",X"DC",X"D1",
		X"C1",X"14",X"C9",X"2A",X"96",X"89",X"11",X"20",X"00",X"19",X"ED",X"5B",X"94",X"89",X"3E",X"FF",
		X"06",X"18",X"77",X"12",X"13",X"23",X"10",X"FA",X"3A",X"51",X"82",X"A7",X"C8",X"47",X"DD",X"2A",
		X"96",X"89",X"0E",X"00",X"CD",X"24",X"0F",X"3A",X"00",X"80",X"E6",X"1E",X"C6",X"E0",X"6F",X"3A",
		X"8F",X"82",X"67",X"5E",X"23",X"56",X"EB",X"18",X"37",X"00",X"DD",X"2A",X"96",X"89",X"11",X"20",
		X"00",X"DD",X"19",X"0E",X"01",X"06",X"0A",X"DD",X"2A",X"92",X"89",X"3A",X"20",X"80",X"A7",X"20",
		X"05",X"3E",X"34",X"32",X"8F",X"82",X"79",X"A7",X"28",X"CA",X"CD",X"24",X"0F",X"3A",X"01",X"80",
		X"E6",X"3F",X"67",X"3A",X"00",X"80",X"E6",X"1F",X"6F",X"5C",X"55",X"CD",X"E0",X"14",X"38",X"E6",
		X"C5",X"0E",X"0A",X"ED",X"5B",X"94",X"89",X"06",X"04",X"CD",X"1B",X"14",X"C1",X"38",X"D7",X"3A",
		X"51",X"82",X"A7",X"28",X"14",X"C5",X"4F",X"E5",X"2A",X"96",X"89",X"11",X"20",X"00",X"19",X"EB",
		X"E1",X"06",X"03",X"CD",X"1B",X"14",X"C1",X"38",X"BD",X"C5",X"11",X"17",X"14",X"01",X"02",X"05",
		X"CD",X"1B",X"14",X"C1",X"38",X"B0",X"DD",X"74",X"21",X"DD",X"75",X"20",X"7D",X"87",X"87",X"87",
		X"CB",X"3C",X"1F",X"CB",X"3C",X"1F",X"CB",X"3C",X"1F",X"6F",X"7C",X"E6",X"07",X"F6",X"98",X"67",
		X"DD",X"74",X"01",X"DD",X"75",X"00",X"DD",X"23",X"DD",X"23",X"10",X"8A",X"3A",X"20",X"80",X"A7",
		X"C0",X"3E",X"28",X"32",X"8F",X"82",X"C9",X"0F",X"00",X"0F",X"32",X"1A",X"13",X"FE",X"FF",X"28",
		X"16",X"95",X"F2",X"27",X"14",X"ED",X"44",X"B8",X"30",X"0D",X"1A",X"FE",X"FF",X"28",X"08",X"94",
		X"F2",X"35",X"14",X"ED",X"44",X"B8",X"D8",X"13",X"0D",X"20",X"E0",X"AF",X"C9",X"0E",X"80",X"E5",
		X"7B",X"0F",X"0F",X"C6",X"04",X"E6",X"07",X"6F",X"7A",X"26",X"40",X"17",X"17",X"17",X"CB",X"14",
		X"E6",X"E0",X"B5",X"24",X"C6",X"80",X"30",X"01",X"24",X"6F",X"71",X"CB",X"DC",X"7E",X"E6",X"3F",
		X"CB",X"4B",X"28",X"02",X"F6",X"40",X"CB",X"4A",X"28",X"02",X"F6",X"80",X"77",X"E1",X"C9",X"2A",
		X"94",X"89",X"AF",X"32",X"B4",X"82",X"0E",X"C6",X"06",X"0A",X"5E",X"7B",X"23",X"56",X"23",X"A2",
		X"3C",X"28",X"03",X"CD",X"3F",X"14",X"10",X"F2",X"2B",X"56",X"2B",X"5E",X"7B",X"A2",X"3C",X"C8",
		X"7B",X"0F",X"0F",X"C6",X"04",X"E6",X"07",X"6F",X"7A",X"26",X"40",X"17",X"17",X"17",X"CB",X"14",
		X"E6",X"E0",X"B5",X"24",X"C6",X"80",X"30",X"01",X"24",X"6F",X"22",X"B5",X"82",X"3E",X"01",X"32",
		X"B4",X"82",X"C9",X"E5",X"D5",X"C5",X"AF",X"EB",X"CD",X"E0",X"14",X"30",X"1F",X"15",X"1D",X"21",
		X"31",X"25",X"0E",X"03",X"06",X"03",X"CD",X"E0",X"14",X"30",X"01",X"B6",X"23",X"14",X"10",X"F6",
		X"15",X"15",X"15",X"1C",X"0D",X"20",X"ED",X"A7",X"20",X"02",X"F6",X"87",X"C1",X"D1",X"E1",X"C9",
		X"D5",X"C5",X"4F",X"7A",X"FE",X"20",X"30",X"1F",X"E6",X"07",X"47",X"04",X"7B",X"FE",X"38",X"30",
		X"16",X"7A",X"87",X"87",X"87",X"87",X"CB",X"13",X"87",X"CB",X"13",X"3A",X"8F",X"82",X"57",X"1A",
		X"87",X"10",X"FD",X"79",X"C1",X"D1",X"C9",X"79",X"C1",X"D1",X"37",X"C9",X"C5",X"D5",X"E5",X"7C",
		X"FE",X"38",X"D2",X"A3",X"15",X"7D",X"FE",X"20",X"D2",X"A3",X"15",X"87",X"87",X"87",X"CB",X"3C",
		X"1F",X"CB",X"3C",X"1F",X"CB",X"3C",X"1F",X"6F",X"7C",X"E6",X"07",X"F6",X"98",X"67",X"4E",X"79",
		X"E6",X"F8",X"CA",X"74",X"15",X"7A",X"87",X"82",X"83",X"87",X"87",X"21",X"05",X"25",X"85",X"30",
		X"01",X"24",X"6F",X"1E",X"00",X"46",X"23",X"7E",X"A1",X"28",X"02",X"CB",X"D3",X"23",X"7E",X"A1",
		X"28",X"02",X"CB",X"CB",X"23",X"7E",X"A1",X"28",X"02",X"CB",X"C3",X"7B",X"21",X"29",X"25",X"85",
		X"30",X"01",X"24",X"6F",X"4E",X"2A",X"56",X"80",X"71",X"CB",X"DC",X"3A",X"B1",X"82",X"B0",X"77",
		X"E1",X"D1",X"C1",X"C9",X"AF",X"47",X"67",X"69",X"29",X"29",X"29",X"09",X"4A",X"09",X"09",X"09",
		X"4B",X"09",X"01",X"52",X"25",X"09",X"ED",X"5B",X"56",X"80",X"7E",X"E6",X"C0",X"F6",X"15",X"47",
		X"7E",X"CB",X"6F",X"28",X"01",X"04",X"E6",X"1F",X"CB",X"FF",X"12",X"EB",X"CB",X"DC",X"70",X"E1",
		X"D1",X"C1",X"C9",X"3A",X"D6",X"82",X"82",X"82",X"82",X"83",X"ED",X"5B",X"56",X"80",X"12",X"06",
		X"51",X"3A",X"D6",X"82",X"FE",X"5F",X"38",X"E3",X"D6",X"09",X"04",X"18",X"F7",X"3A",X"4E",X"82",
		X"A7",X"C8",X"21",X"F8",X"01",X"F3",X"ED",X"5B",X"54",X"80",X"3A",X"50",X"80",X"06",X"00",X"4F",
		X"CB",X"7F",X"28",X"01",X"05",X"09",X"01",X"F8",X"FF",X"1C",X"1D",X"28",X"03",X"09",X"18",X"FA",
		X"22",X"48",X"82",X"3A",X"51",X"80",X"C6",X"14",X"ED",X"44",X"14",X"15",X"28",X"03",X"91",X"18",
		X"FA",X"32",X"4A",X"82",X"3A",X"4E",X"82",X"47",X"DD",X"21",X"93",X"80",X"2A",X"52",X"80",X"DD",
		X"7E",X"FD",X"95",X"FE",X"0B",X"30",X"0A",X"4F",X"DD",X"7E",X"FF",X"94",X"FE",X"0B",X"57",X"38",
		X"09",X"11",X"20",X"00",X"DD",X"19",X"10",X"E4",X"FB",X"C9",X"DD",X"E5",X"E1",X"FD",X"21",X"02",
		X"80",X"1E",X"06",X"FD",X"7E",X"00",X"BD",X"20",X"06",X"FD",X"7E",X"01",X"BC",X"28",X"E2",X"FD",
		X"23",X"FD",X"23",X"1D",X"20",X"ED",X"1E",X"06",X"FD",X"2B",X"FD",X"2B",X"FD",X"7E",X"00",X"FD",
		X"B6",X"01",X"28",X"10",X"1D",X"20",X"F1",X"11",X"F5",X"FF",X"DD",X"19",X"CD",X"85",X"18",X"11",
		X"2B",X"00",X"18",X"C0",X"FD",X"75",X"00",X"FD",X"74",X"01",X"7A",X"87",X"82",X"87",X"87",X"87",
		X"57",X"3A",X"4A",X"82",X"92",X"DD",X"77",X"03",X"79",X"87",X"81",X"87",X"87",X"87",X"5F",X"16",
		X"00",X"2A",X"48",X"82",X"19",X"DD",X"74",X"00",X"DD",X"75",X"01",X"AF",X"DD",X"77",X"FC",X"DD",
		X"77",X"FA",X"C3",X"11",X"16",X"E5",X"F5",X"3A",X"4D",X"80",X"6F",X"3A",X"4F",X"80",X"ED",X"44",
		X"67",X"3A",X"50",X"80",X"85",X"E6",X"F8",X"D6",X"10",X"0F",X"0F",X"0F",X"6F",X"3A",X"51",X"80",
		X"84",X"26",X"21",X"07",X"CB",X"14",X"07",X"CB",X"14",X"E6",X"E0",X"B5",X"6F",X"22",X"56",X"80",
		X"F1",X"E1",X"C9",X"00",X"E5",X"D5",X"C5",X"F5",X"3A",X"AA",X"82",X"A7",X"20",X"07",X"21",X"24",
		X"80",X"36",X"FF",X"18",X"3C",X"21",X"AC",X"82",X"3A",X"00",X"A0",X"47",X"1F",X"CB",X"16",X"23",
		X"CB",X"10",X"CB",X"16",X"23",X"3A",X"80",X"A0",X"17",X"CB",X"16",X"7E",X"E6",X"0F",X"FE",X"0C",
		X"CC",X"06",X"17",X"2B",X"7E",X"E6",X"0F",X"FE",X"0C",X"CC",X"06",X"17",X"2B",X"7E",X"E6",X"0F",
		X"06",X"01",X"FE",X"0C",X"20",X"0B",X"3A",X"F6",X"89",X"CB",X"F7",X"32",X"F6",X"89",X"CD",X"18",
		X"17",X"F1",X"C1",X"D1",X"E1",X"C9",X"EB",X"21",X"A8",X"82",X"34",X"23",X"34",X"CB",X"46",X"23",
		X"28",X"01",X"23",X"46",X"EB",X"78",X"A7",X"C8",X"EB",X"21",X"24",X"80",X"34",X"20",X"01",X"35",
		X"10",X"FA",X"EB",X"3A",X"21",X"80",X"A7",X"28",X"09",X"3A",X"20",X"80",X"FE",X"01",X"CC",X"35",
		X"21",X"C9",X"21",X"F4",X"89",X"77",X"23",X"77",X"C3",X"5A",X"07",X"3A",X"A8",X"82",X"A7",X"C8",
		X"E5",X"D5",X"C5",X"21",X"AF",X"82",X"11",X"87",X"A1",X"7E",X"23",X"A7",X"20",X"0B",X"AF",X"77",
		X"3C",X"12",X"2B",X"36",X"01",X"C1",X"D1",X"E1",X"C9",X"34",X"7E",X"FE",X"10",X"20",X"0E",X"2B",
		X"36",X"00",X"21",X"A8",X"82",X"35",X"21",X"F6",X"89",X"36",X"80",X"18",X"E8",X"D6",X"08",X"20",
		X"E4",X"12",X"18",X"E1",X"DD",X"21",X"68",X"80",X"DD",X"6E",X"11",X"DD",X"66",X"12",X"DD",X"7E",
		X"05",X"C6",X"0C",X"FE",X"19",X"38",X"08",X"CB",X"7F",X"20",X"03",X"23",X"18",X"01",X"2B",X"DD",
		X"7E",X"07",X"11",X"20",X"00",X"C6",X"0C",X"FE",X"19",X"38",X"0A",X"CB",X"7F",X"28",X"03",X"19",
		X"18",X"03",X"A7",X"ED",X"52",X"EB",X"2A",X"92",X"89",X"06",X"0A",X"7B",X"BE",X"23",X"20",X"02",
		X"7A",X"BE",X"23",X"CA",X"A1",X"19",X"10",X"F3",X"3A",X"4C",X"82",X"A7",X"C2",X"61",X"18",X"1A",
		X"FE",X"03",X"CA",X"AA",X"1B",X"DD",X"21",X"88",X"80",X"FD",X"21",X"A8",X"80",X"06",X"07",X"C5",
		X"FD",X"E5",X"DD",X"7E",X"13",X"A7",X"28",X"05",X"DD",X"35",X"13",X"18",X"2C",X"DD",X"7E",X"08",
		X"FD",X"96",X"08",X"6F",X"DD",X"7E",X"05",X"FD",X"96",X"05",X"CD",X"B1",X"18",X"20",X"13",X"DD",
		X"7E",X"0A",X"FD",X"96",X"0A",X"6F",X"FD",X"7E",X"07",X"DD",X"96",X"07",X"CD",X"B1",X"18",X"CC",
		X"68",X"18",X"11",X"20",X"00",X"FD",X"19",X"10",X"C9",X"11",X"20",X"00",X"FD",X"E1",X"C1",X"DD",
		X"19",X"FD",X"19",X"10",X"BA",X"06",X"08",X"DD",X"21",X"88",X"80",X"DD",X"7E",X"13",X"A7",X"20",
		X"37",X"DD",X"66",X"12",X"DD",X"6E",X"11",X"DD",X"7E",X"05",X"C6",X"0C",X"FE",X"19",X"38",X"0C",
		X"CB",X"7F",X"20",X"05",X"CD",X"1B",X"0F",X"18",X"03",X"CD",X"11",X"0F",X"DD",X"7E",X"07",X"11",
		X"20",X"00",X"C6",X"0C",X"FE",X"19",X"38",X"0A",X"CB",X"7F",X"28",X"03",X"19",X"18",X"03",X"A7",
		X"ED",X"52",X"7E",X"FE",X"03",X"CC",X"85",X"18",X"11",X"20",X"00",X"DD",X"19",X"05",X"C2",X"1B",
		X"18",X"21",X"22",X"80",X"34",X"C3",X"2C",X"0C",X"DD",X"E5",X"FD",X"E5",X"DD",X"E1",X"CD",X"85",
		X"18",X"DD",X"E1",X"FD",X"7E",X"02",X"DD",X"AE",X"02",X"CB",X"7F",X"DD",X"7E",X"02",X"28",X"02",
		X"ED",X"44",X"DD",X"77",X"02",X"E5",X"DD",X"36",X"00",X"E0",X"DD",X"36",X"13",X"32",X"21",X"00",
		X"01",X"DD",X"CB",X"02",X"7E",X"20",X"02",X"26",X"FF",X"DD",X"74",X"02",X"DD",X"75",X"01",X"06",
		X"08",X"FD",X"E5",X"FD",X"2E",X"00",X"CD",X"F3",X"00",X"10",X"FB",X"FD",X"E1",X"06",X"01",X"E1",
		X"C9",X"2D",X"2D",X"C6",X"23",X"CB",X"7F",X"20",X"05",X"2C",X"D6",X"18",X"18",X"F7",X"7D",X"A7",
		X"C9",X"3E",X"03",X"32",X"20",X"80",X"3E",X"EC",X"32",X"14",X"80",X"21",X"F4",X"89",X"36",X"80",
		X"23",X"36",X"08",X"CD",X"60",X"19",X"AF",X"32",X"B4",X"82",X"3A",X"21",X"80",X"A7",X"CA",X"3D",
		X"07",X"2A",X"88",X"89",X"35",X"CA",X"CD",X"1B",X"21",X"AA",X"81",X"7E",X"47",X"23",X"A6",X"CA",
		X"1C",X"19",X"78",X"FE",X"02",X"28",X"0B",X"CD",X"33",X"19",X"3E",X"01",X"32",X"B7",X"81",X"C3",
		X"1C",X"19",X"CD",X"46",X"19",X"3E",X"01",X"32",X"B7",X"81",X"21",X"0E",X"80",X"3A",X"B2",X"81",
		X"CB",X"47",X"C2",X"1C",X"19",X"7E",X"23",X"23",X"BE",X"CA",X"BF",X"08",X"2A",X"8A",X"89",X"7E",
		X"E6",X"03",X"CA",X"BF",X"08",X"AF",X"32",X"4B",X"82",X"3A",X"4B",X"82",X"FE",X"78",X"20",X"F9",
		X"C3",X"E7",X"08",X"2B",X"36",X"02",X"2B",X"7E",X"2B",X"77",X"21",X"63",X"21",X"11",X"88",X"89",
		X"01",X"18",X"00",X"ED",X"B0",X"C9",X"2B",X"36",X"01",X"2B",X"46",X"2B",X"AF",X"77",X"21",X"7B",
		X"21",X"11",X"88",X"89",X"78",X"01",X"16",X"00",X"A7",X"28",X"02",X"03",X"03",X"ED",X"B0",X"C9",
		X"3E",X"20",X"90",X"90",X"6F",X"26",X"80",X"36",X"EC",X"DD",X"7E",X"0C",X"D6",X"08",X"47",X"DD",
		X"7E",X"0E",X"C6",X"08",X"4F",X"CD",X"31",X"10",X"54",X"5D",X"CB",X"DC",X"3E",X"B4",X"0E",X"03",
		X"E5",X"D5",X"06",X"03",X"12",X"36",X"46",X"CD",X"0F",X"10",X"3C",X"10",X"F7",X"D1",X"E1",X"CD",
		X"1E",X"10",X"0D",X"20",X"EB",X"2A",X"98",X"89",X"06",X"04",X"3E",X"66",X"77",X"23",X"10",X"FC",
		X"C9",X"E5",X"3E",X"01",X"32",X"B3",X"82",X"AF",X"12",X"05",X"21",X"F4",X"89",X"0E",X"04",X"28",
		X"06",X"05",X"CC",X"62",X"1E",X"18",X"09",X"0E",X"08",X"3A",X"23",X"80",X"3C",X"32",X"23",X"80",
		X"7E",X"B1",X"77",X"E1",X"AF",X"2B",X"77",X"2B",X"77",X"11",X"20",X"00",X"19",X"3D",X"5E",X"77",
		X"23",X"56",X"77",X"CD",X"3D",X"14",X"CD",X"6F",X"14",X"DD",X"7E",X"05",X"C6",X"0C",X"FE",X"19",
		X"38",X"08",X"D6",X"18",X"FE",X"1E",X"38",X"02",X"C6",X"30",X"D6",X"0C",X"ED",X"44",X"DD",X"86",
		X"0C",X"47",X"DD",X"7E",X"07",X"C6",X"0C",X"FE",X"19",X"38",X"08",X"D6",X"18",X"FE",X"1E",X"38",
		X"02",X"C6",X"30",X"D6",X"0C",X"ED",X"44",X"DD",X"86",X"0E",X"4F",X"C5",X"CD",X"31",X"10",X"36",
		X"81",X"C1",X"E5",X"C5",X"78",X"D6",X"08",X"47",X"C5",X"CD",X"31",X"10",X"36",X"81",X"C1",X"79",
		X"D6",X"08",X"4F",X"C5",X"CD",X"31",X"10",X"36",X"81",X"C1",X"79",X"C1",X"4F",X"CD",X"31",X"10",
		X"36",X"81",X"E1",X"7D",X"E6",X"1F",X"11",X"20",X"00",X"20",X"01",X"19",X"2B",X"3A",X"50",X"82",
		X"3C",X"32",X"50",X"82",X"FE",X"0A",X"20",X"02",X"3E",X"01",X"C6",X"9F",X"77",X"CD",X"8D",X"1A",
		X"CD",X"9C",X"1B",X"36",X"AA",X"CD",X"8D",X"1A",X"3A",X"50",X"82",X"FE",X"0A",X"20",X"08",X"CD",
		X"9C",X"1B",X"36",X"AB",X"CD",X"8D",X"1A",X"3A",X"23",X"80",X"E6",X"01",X"28",X"28",X"E5",X"CD",
		X"9C",X"1B",X"7E",X"FE",X"81",X"20",X"08",X"36",X"AC",X"CD",X"8D",X"1A",X"E1",X"18",X"17",X"E1",
		X"11",X"20",X"00",X"19",X"7C",X"E6",X"07",X"F6",X"84",X"67",X"E5",X"18",X"E5",X"CB",X"DC",X"CB",
		X"F6",X"CB",X"BE",X"CB",X"9C",X"C9",X"2A",X"8C",X"89",X"34",X"7E",X"FE",X"0A",X"20",X"05",X"3E",
		X"03",X"32",X"20",X"80",X"3A",X"50",X"82",X"47",X"3A",X"23",X"80",X"E6",X"01",X"28",X"09",X"4F",
		X"78",X"CB",X"20",X"0D",X"28",X"02",X"80",X"47",X"0E",X"0A",X"C5",X"CD",X"64",X"20",X"CD",X"0F",
		X"21",X"C1",X"0D",X"20",X"F5",X"10",X"F1",X"CD",X"64",X"20",X"3A",X"23",X"80",X"CB",X"4F",X"C4",
		X"6B",X"1E",X"CD",X"1F",X"1B",X"2A",X"8C",X"89",X"AF",X"32",X"B3",X"82",X"7E",X"FE",X"0A",X"C2",
		X"C5",X"17",X"3A",X"21",X"80",X"A7",X"CA",X"3D",X"07",X"CD",X"95",X"19",X"21",X"F4",X"89",X"7E",
		X"E6",X"3F",X"77",X"23",X"36",X"28",X"3E",X"EC",X"32",X"14",X"80",X"3E",X"03",X"32",X"20",X"80",
		X"32",X"4B",X"82",X"3A",X"4B",X"82",X"E6",X"3F",X"20",X"F9",X"CB",X"46",X"28",X"FC",X"CD",X"A9",
		X"1F",X"3E",X"E0",X"32",X"4B",X"82",X"3A",X"4B",X"82",X"A7",X"20",X"FA",X"C3",X"BF",X"08",X"3A",
		X"92",X"82",X"A7",X"C0",X"2A",X"8A",X"89",X"7E",X"3D",X"0F",X"0F",X"E6",X"03",X"47",X"04",X"F6",
		X"30",X"32",X"8F",X"82",X"D6",X"23",X"32",X"B1",X"82",X"3E",X"53",X"C6",X"09",X"10",X"FC",X"32",
		X"D6",X"82",X"3A",X"D8",X"82",X"57",X"7E",X"BA",X"38",X"04",X"D6",X"04",X"18",X"F9",X"D6",X"02",
		X"87",X"87",X"87",X"6F",X"26",X"00",X"ED",X"5B",X"D2",X"82",X"19",X"7E",X"32",X"4E",X"82",X"23",
		X"7E",X"32",X"6E",X"82",X"23",X"7E",X"32",X"88",X"82",X"23",X"7E",X"32",X"51",X"82",X"23",X"3A",
		X"8A",X"82",X"47",X"ED",X"5B",X"8C",X"89",X"1A",X"05",X"28",X"11",X"23",X"05",X"28",X"0D",X"FE",
		X"08",X"30",X"09",X"23",X"05",X"28",X"05",X"FE",X"05",X"30",X"01",X"23",X"5E",X"16",X"00",X"21",
		X"DD",X"23",X"19",X"11",X"25",X"80",X"01",X"08",X"00",X"ED",X"B0",X"C9",X"23",X"47",X"7D",X"E6",
		X"1F",X"78",X"C0",X"2B",X"7D",X"E6",X"E0",X"6F",X"78",X"C9",X"3E",X"03",X"32",X"20",X"80",X"3E",
		X"EC",X"32",X"14",X"80",X"21",X"F4",X"89",X"36",X"80",X"23",X"36",X"08",X"CD",X"60",X"19",X"3A",
		X"21",X"80",X"A7",X"CA",X"3D",X"07",X"2A",X"88",X"89",X"35",X"C2",X"E8",X"18",X"3E",X"A0",X"32",
		X"4B",X"82",X"3A",X"4B",X"82",X"A7",X"20",X"FA",X"AF",X"32",X"F4",X"89",X"DD",X"7E",X"0C",X"D6",
		X"08",X"47",X"DD",X"7E",X"0E",X"C6",X"08",X"4F",X"CD",X"31",X"10",X"54",X"5D",X"06",X"03",X"3E",
		X"81",X"E5",X"D5",X"0E",X"03",X"12",X"CD",X"0F",X"10",X"0D",X"20",X"F9",X"D1",X"E1",X"CD",X"1E",
		X"10",X"10",X"EE",X"DD",X"21",X"14",X"80",X"FD",X"21",X"14",X"88",X"3A",X"A8",X"81",X"A7",X"20",
		X"22",X"DD",X"36",X"00",X"E0",X"DD",X"36",X"01",X"68",X"FD",X"36",X"00",X"74",X"FD",X"36",X"01",
		X"66",X"DD",X"36",X"02",X"E4",X"DD",X"36",X"03",X"78",X"FD",X"36",X"02",X"74",X"FD",X"36",X"03",
		X"66",X"18",X"20",X"DD",X"36",X"00",X"E3",X"DD",X"36",X"01",X"AC",X"DD",X"36",X"02",X"E7",X"DD",
		X"36",X"03",X"9C",X"FD",X"36",X"00",X"7C",X"FD",X"36",X"01",X"66",X"FD",X"36",X"02",X"7C",X"FD",
		X"36",X"03",X"66",X"3E",X"01",X"32",X"4B",X"82",X"3A",X"4B",X"82",X"E6",X"3F",X"20",X"F9",X"3A",
		X"D0",X"82",X"A7",X"CA",X"EC",X"1C",X"3E",X"75",X"CD",X"E5",X"20",X"21",X"3D",X"1D",X"11",X"07",
		X"85",X"CD",X"29",X"1D",X"11",X"86",X"85",X"CD",X"29",X"1D",X"11",X"C9",X"85",X"CD",X"29",X"1D",
		X"11",X"86",X"86",X"CD",X"29",X"1D",X"11",X"C8",X"86",X"CD",X"29",X"1D",X"3E",X"83",X"32",X"2F",
		X"86",X"21",X"F5",X"89",X"CB",X"D6",X"3E",X"01",X"32",X"4B",X"82",X"3A",X"4B",X"82",X"E6",X"0F",
		X"20",X"F9",X"CB",X"46",X"20",X"46",X"11",X"60",X"88",X"1A",X"EE",X"1F",X"06",X"08",X"12",X"13",
		X"10",X"FC",X"E5",X"11",X"2F",X"86",X"1A",X"11",X"28",X"86",X"FE",X"40",X"20",X"1D",X"21",X"64",
		X"80",X"01",X"04",X"00",X"ED",X"B0",X"0E",X"04",X"21",X"60",X"80",X"ED",X"B0",X"3E",X"22",X"12",
		X"1B",X"1A",X"FE",X"40",X"20",X"FA",X"3E",X"22",X"12",X"18",X"08",X"06",X"09",X"3E",X"40",X"12",
		X"13",X"10",X"FC",X"CD",X"F0",X"04",X"CD",X"09",X"1D",X"E1",X"18",X"AA",X"CD",X"95",X"19",X"CD",
		X"1A",X"1D",X"21",X"60",X"88",X"06",X"08",X"36",X"70",X"23",X"10",X"FB",X"21",X"AA",X"81",X"7E",
		X"23",X"A6",X"77",X"C2",X"E8",X"18",X"C3",X"3D",X"07",X"2A",X"98",X"89",X"01",X"1C",X"00",X"09",
		X"06",X"08",X"7E",X"EE",X"15",X"77",X"23",X"10",X"FC",X"C9",X"2A",X"98",X"89",X"01",X"1C",X"00",
		X"09",X"06",X"08",X"36",X"72",X"23",X"10",X"FB",X"C9",X"F5",X"C5",X"D5",X"7E",X"CB",X"DA",X"23",
		X"46",X"12",X"13",X"10",X"FC",X"4E",X"D1",X"23",X"ED",X"B0",X"C1",X"F1",X"C9",X"75",X"0D",X"59",
		X"4F",X"55",X"40",X"44",X"49",X"44",X"40",X"49",X"54",X"40",X"21",X"21",X"74",X"0E",X"54",X"48",
		X"45",X"40",X"48",X"49",X"47",X"48",X"40",X"53",X"43",X"4F",X"52",X"45",X"74",X"0B",X"4F",X"46",
		X"40",X"54",X"48",X"45",X"40",X"44",X"41",X"59",X"2E",X"76",X"10",X"47",X"4F",X"40",X"46",X"4F",
		X"52",X"40",X"54",X"48",X"45",X"40",X"57",X"4F",X"52",X"4C",X"44",X"76",X"0D",X"52",X"45",X"43",
		X"4F",X"52",X"44",X"40",X"4E",X"4F",X"57",X"40",X"21",X"21",X"E5",X"C5",X"21",X"34",X"88",X"06",
		X"0C",X"0E",X"00",X"71",X"23",X"10",X"FC",X"C1",X"E1",X"C9",X"E5",X"21",X"91",X"82",X"36",X"03",
		X"E1",X"C9",X"D9",X"06",X"FF",X"FD",X"21",X"88",X"80",X"3A",X"4E",X"82",X"47",X"DD",X"7E",X"08",
		X"FD",X"96",X"08",X"30",X"02",X"ED",X"44",X"57",X"FD",X"7E",X"0A",X"DD",X"96",X"0A",X"30",X"02",
		X"ED",X"44",X"B2",X"FE",X"04",X"DC",X"9A",X"1D",X"11",X"20",X"00",X"FD",X"19",X"10",X"DE",X"3E",
		X"34",X"32",X"8F",X"82",X"3E",X"FF",X"D9",X"47",X"C9",X"3E",X"30",X"32",X"8F",X"82",X"C9",X"DD",
		X"21",X"68",X"80",X"06",X"09",X"21",X"3A",X"25",X"DD",X"7E",X"15",X"A7",X"20",X"43",X"DD",X"4E",
		X"02",X"79",X"DD",X"B6",X"01",X"28",X"3A",X"DD",X"7E",X"03",X"A7",X"28",X"08",X"CB",X"79",X"28",
		X"0E",X"0E",X"FD",X"18",X"0C",X"CB",X"79",X"28",X"03",X"0E",X"F2",X"11",X"0E",X"F0",X"11",X"0E",
		X"FC",X"DD",X"7E",X"0F",X"B9",X"28",X"1A",X"79",X"BE",X"23",X"20",X"FC",X"DD",X"7E",X"0F",X"0E",
		X"00",X"0C",X"BE",X"23",X"20",X"FB",X"79",X"FE",X"06",X"30",X"02",X"2B",X"2B",X"7E",X"DD",X"77",
		X"0F",X"11",X"20",X"00",X"DD",X"19",X"10",X"AD",X"AF",X"32",X"4B",X"82",X"C9",X"4E",X"23",X"06",
		X"00",X"ED",X"B0",X"C9",X"3A",X"24",X"80",X"A7",X"28",X"04",X"06",X"01",X"18",X"02",X"06",X"00",
		X"21",X"84",X"A1",X"70",X"23",X"3A",X"24",X"80",X"FE",X"01",X"20",X"02",X"06",X"00",X"70",X"3E",
		X"01",X"C9",X"3A",X"23",X"80",X"C6",X"02",X"32",X"23",X"80",X"C9",X"CB",X"8F",X"32",X"23",X"80",
		X"2A",X"8C",X"89",X"7E",X"FE",X"0A",X"C8",X"3A",X"20",X"80",X"A7",X"C8",X"F5",X"3E",X"03",X"32",
		X"20",X"80",X"DD",X"E5",X"DD",X"2A",X"8E",X"89",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"E5",X"CD",
		X"A9",X"1F",X"E1",X"2C",X"DD",X"75",X"00",X"DD",X"74",X"01",X"CD",X"13",X"1F",X"DD",X"E1",X"2A",
		X"9A",X"89",X"AF",X"77",X"32",X"92",X"82",X"32",X"8A",X"82",X"F1",X"32",X"20",X"80",X"C9",X"D5",
		X"C5",X"01",X"08",X"00",X"ED",X"B0",X"C1",X"D1",X"E5",X"D5",X"EB",X"CB",X"DC",X"16",X"08",X"71",
		X"23",X"15",X"20",X"FB",X"D1",X"21",X"20",X"00",X"19",X"EB",X"E1",X"C9",X"00",X"3A",X"21",X"80",
		X"A7",X"C8",X"2A",X"9C",X"89",X"7E",X"A7",X"C8",X"3A",X"69",X"82",X"47",X"3A",X"6E",X"82",X"B8",
		X"C0",X"AF",X"32",X"69",X"82",X"DD",X"2A",X"8E",X"89",X"DD",X"7E",X"01",X"21",X"6F",X"22",X"FE",
		X"0A",X"30",X"03",X"21",X"77",X"22",X"11",X"40",X"89",X"01",X"08",X"00",X"ED",X"B0",X"DD",X"7E",
		X"00",X"A7",X"20",X"0F",X"DD",X"7E",X"01",X"FE",X"0A",X"20",X"08",X"3A",X"F4",X"89",X"F6",X"20",
		X"32",X"F4",X"89",X"DD",X"2A",X"8E",X"89",X"DD",X"66",X"01",X"DD",X"6E",X"00",X"7C",X"B5",X"C8",
		X"2D",X"CB",X"7D",X"28",X"03",X"2E",X"09",X"25",X"DD",X"75",X"00",X"DD",X"74",X"01",X"7C",X"DD",
		X"5E",X"01",X"21",X"44",X"81",X"16",X"36",X"0E",X"C7",X"3E",X"05",X"93",X"FE",X"CF",X"38",X"02",
		X"3E",X"CF",X"77",X"2C",X"06",X"07",X"7A",X"BB",X"30",X"01",X"5A",X"D6",X"08",X"57",X"7B",X"92",
		X"CB",X"7F",X"28",X"01",X"AF",X"81",X"77",X"7D",X"3C",X"E6",X"F7",X"6F",X"10",X"E8",X"DD",X"7E",
		X"01",X"A7",X"C0",X"DD",X"7E",X"00",X"FE",X"01",X"28",X"07",X"A7",X"C0",X"3C",X"32",X"92",X"82",
		X"C9",X"2A",X"9A",X"89",X"36",X"C7",X"21",X"8C",X"82",X"36",X"01",X"C9",X"DD",X"2A",X"8E",X"89",
		X"21",X"6F",X"22",X"11",X"40",X"89",X"01",X"08",X"00",X"ED",X"B0",X"C3",X"2F",X"1F",X"47",X"3A",
		X"B4",X"82",X"FE",X"00",X"78",X"C8",X"2A",X"B5",X"82",X"36",X"80",X"C9",X"47",X"3A",X"B4",X"82",
		X"A7",X"78",X"C8",X"2A",X"B5",X"82",X"36",X"C6",X"C9",X"DD",X"2A",X"8E",X"89",X"3A",X"20",X"80",
		X"A7",X"C8",X"06",X"03",X"DD",X"7E",X"00",X"DD",X"B6",X"01",X"C8",X"3A",X"F4",X"89",X"E6",X"03",
		X"F6",X"02",X"32",X"F4",X"89",X"AF",X"32",X"69",X"82",X"E5",X"2A",X"8A",X"89",X"7E",X"E1",X"FE",
		X"0D",X"38",X"2A",X"06",X"05",X"DD",X"7E",X"00",X"DD",X"B6",X"01",X"C8",X"C5",X"CD",X"13",X"1F",
		X"CD",X"0F",X"21",X"CD",X"64",X"20",X"CD",X"13",X"1F",X"CD",X"0F",X"21",X"CD",X"64",X"20",X"76",
		X"C1",X"10",X"E2",X"3A",X"69",X"82",X"FE",X"05",X"38",X"F9",X"C3",X"A9",X"1F",X"FE",X"09",X"38",
		X"24",X"DD",X"7E",X"00",X"DD",X"B6",X"01",X"C8",X"C5",X"CD",X"13",X"1F",X"CD",X"13",X"1F",X"CD",
		X"13",X"1F",X"CD",X"0F",X"21",X"CD",X"64",X"20",X"76",X"CD",X"0F",X"21",X"CD",X"64",X"20",X"C1",
		X"10",X"DF",X"C3",X"F3",X"1F",X"FE",X"05",X"38",X"1D",X"06",X"05",X"DD",X"7E",X"00",X"DD",X"B6",
		X"01",X"C8",X"C5",X"CD",X"13",X"1F",X"CD",X"13",X"1F",X"CD",X"0F",X"21",X"CD",X"64",X"20",X"76",
		X"C1",X"10",X"E8",X"C3",X"F3",X"1F",X"DD",X"7E",X"00",X"DD",X"B6",X"01",X"C8",X"C5",X"CD",X"13",
		X"1F",X"CD",X"13",X"1F",X"CD",X"13",X"1F",X"CD",X"0F",X"21",X"CD",X"64",X"20",X"76",X"C1",X"10",
		X"E5",X"C3",X"F3",X"1F",X"3A",X"20",X"80",X"A7",X"C8",X"3A",X"D0",X"82",X"11",X"60",X"80",X"2A",
		X"90",X"89",X"01",X"08",X"00",X"FE",X"01",X"20",X"04",X"ED",X"B0",X"18",X"12",X"1A",X"FE",X"40",
		X"28",X"03",X"BE",X"20",X"0A",X"23",X"13",X"0D",X"20",X"F3",X"3E",X"01",X"32",X"D0",X"82",X"3A",
		X"B2",X"81",X"4F",X"3A",X"AA",X"81",X"A1",X"20",X"29",X"2A",X"90",X"89",X"ED",X"5B",X"B3",X"81",
		X"06",X"08",X"1A",X"BE",X"20",X"1C",X"23",X"13",X"10",X"F8",X"3A",X"AA",X"81",X"B1",X"32",X"B2",
		X"81",X"2A",X"88",X"89",X"34",X"DD",X"E5",X"CD",X"2F",X"0B",X"DD",X"E1",X"21",X"F4",X"89",X"CB",
		X"C6",X"C9",X"3A",X"AA",X"81",X"87",X"87",X"A1",X"C0",X"ED",X"5B",X"B9",X"81",X"2A",X"90",X"89",
		X"06",X"08",X"1A",X"BE",X"C0",X"23",X"13",X"10",X"F9",X"3A",X"AA",X"81",X"87",X"87",X"B1",X"32",
		X"B2",X"81",X"C3",X"B1",X"20",X"21",X"00",X"84",X"11",X"01",X"84",X"01",X"FF",X"03",X"36",X"40",
		X"ED",X"B0",X"21",X"00",X"8C",X"11",X"01",X"8C",X"01",X"FF",X"03",X"77",X"ED",X"B0",X"AF",X"32",
		X"40",X"A1",X"32",X"30",X"A1",X"21",X"4C",X"80",X"06",X"04",X"77",X"23",X"10",X"FC",X"C9",X"2A",
		X"90",X"89",X"3A",X"20",X"80",X"A7",X"C8",X"23",X"23",X"7E",X"3C",X"E6",X"0F",X"77",X"FE",X"0A",
		X"D8",X"D6",X"0A",X"77",X"CB",X"DD",X"2D",X"CB",X"9D",X"18",X"EE",X"F5",X"7C",X"2F",X"67",X"7D",
		X"2F",X"6F",X"23",X"F1",X"C9",X"E5",X"D5",X"C5",X"21",X"C7",X"21",X"11",X"6A",X"86",X"CD",X"3D",
		X"1E",X"3A",X"24",X"80",X"21",X"72",X"86",X"06",X"00",X"FE",X"63",X"38",X"02",X"3E",X"63",X"FE",
		X"0A",X"38",X"05",X"04",X"D6",X"0A",X"18",X"F7",X"77",X"78",X"A7",X"28",X"02",X"2B",X"77",X"C1",
		X"D1",X"E1",X"C9",X"0F",X"80",X"B0",X"81",X"71",X"82",X"6A",X"82",X"A0",X"80",X"C8",X"81",X"E8",
		X"81",X"08",X"82",X"84",X"88",X"89",X"82",X"8B",X"82",X"00",X"A0",X"10",X"80",X"B1",X"81",X"72",
		X"82",X"6C",X"82",X"E0",X"80",X"08",X"89",X"28",X"89",X"48",X"89",X"C4",X"88",X"8D",X"82",X"8E",
		X"82",X"80",X"A0",X"11",X"50",X"55",X"53",X"48",X"40",X"53",X"54",X"41",X"52",X"54",X"40",X"42",
		X"55",X"54",X"54",X"4F",X"4E",X"17",X"42",X"4F",X"4E",X"55",X"53",X"40",X"43",X"41",X"52",X"40",
		X"46",X"4F",X"52",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"50",X"54",X"53",X"09",X"46",X"52",
		X"45",X"45",X"40",X"50",X"4C",X"41",X"59",X"09",X"43",X"52",X"45",X"44",X"49",X"54",X"40",X"40",
		X"40",X"73",X"12",X"18",X"40",X"19",X"1A",X"1B",X"1C",X"1D",X"1E",X"1F",X"40",X"31",X"39",X"38",
		X"30",X"40",X"31",X"53",X"54",X"73",X"12",X"18",X"40",X"19",X"1A",X"1B",X"1C",X"1D",X"1E",X"1F",
		X"40",X"31",X"39",X"38",X"31",X"40",X"32",X"4E",X"44",X"18",X"31",X"53",X"54",X"40",X"42",X"4F",
		X"4E",X"55",X"53",X"40",X"46",X"4F",X"52",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"50",
		X"54",X"53",X"40",X"40",X"18",X"32",X"4E",X"44",X"40",X"42",X"4F",X"4E",X"55",X"53",X"40",X"46",
		X"4F",X"52",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"50",X"54",X"53",X"40",X"40",X"43",
		X"4F",X"52",X"45",X"48",X"49",X"2D",X"53",X"40",X"40",X"30",X"30",X"40",X"40",X"40",X"40",X"40",
		X"40",X"40",X"40",X"31",X"55",X"50",X"40",X"40",X"40",X"40",X"40",X"32",X"55",X"50",X"40",X"D4",
		X"D5",X"D6",X"D7",X"D0",X"D1",X"D2",X"D3",X"44",X"40",X"40",X"40",X"52",X"4F",X"55",X"4E",X"40",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"29",
		X"29",X"29",X"2A",X"68",X"29",X"29",X"29",X"30",X"30",X"30",X"31",X"6F",X"30",X"30",X"30",X"43",
		X"48",X"41",X"4C",X"4C",X"45",X"4E",X"47",X"49",X"4E",X"47",X"40",X"53",X"54",X"41",X"47",X"45",
		X"20",X"4E",X"4F",X"2E",X"20",X"3D",X"40",X"20",X"3D",X"40",X"20",X"52",X"45",X"44",X"40",X"43",
		X"41",X"52",X"53",X"40",X"44",X"4F",X"4E",X"27",X"54",X"40",X"4D",X"4F",X"56",X"45",X"20",X"55",
		X"4E",X"54",X"49",X"4C",X"40",X"46",X"55",X"45",X"4C",X"40",X"52",X"55",X"4E",X"53",X"40",X"4F",
		X"55",X"54",X"2E",X"20",X"20",X"20",X"20",X"20",X"4E",X"45",X"57",X"40",X"52",X"41",X"4C",X"4C",
		X"59",X"2D",X"58",X"20",X"40",X"43",X"41",X"53",X"54",X"40",X"40",X"40",X"20",X"4D",X"59",X"40",
		X"43",X"41",X"52",X"20",X"52",X"45",X"44",X"40",X"43",X"41",X"52",X"20",X"43",X"48",X"45",X"43",
		X"4B",X"40",X"50",X"4F",X"49",X"4E",X"54",X"20",X"53",X"50",X"45",X"43",X"49",X"41",X"4C",X"40",
		X"43",X"48",X"45",X"43",X"4B",X"40",X"50",X"4F",X"49",X"4E",X"54",X"20",X"4C",X"55",X"43",X"4B",
		X"59",X"40",X"43",X"48",X"45",X"43",X"4B",X"40",X"50",X"4F",X"49",X"4E",X"54",X"20",X"52",X"4F",
		X"43",X"4B",X"40",X"28",X"40",X"44",X"41",X"4E",X"47",X"45",X"52",X"40",X"21",X"40",X"29",X"20",
		X"53",X"4D",X"4F",X"4B",X"45",X"40",X"53",X"43",X"52",X"45",X"45",X"4E",X"20",X"19",X"1A",X"1B",
		X"1C",X"1D",X"1E",X"1F",X"20",X"01",X"09",X"64",X"00",X"A0",X"08",X"08",X"00",X"02",X"09",X"64",
		X"02",X"A0",X"18",X"18",X"10",X"07",X"07",X"50",X"05",X"A0",X"80",X"80",X"80",X"03",X"08",X"5A",
		X"02",X"A0",X"20",X"20",X"10",X"03",X"08",X"5A",X"03",X"A0",X"30",X"30",X"28",X"04",X"07",X"50",
		X"03",X"A0",X"38",X"38",X"30",X"07",X"07",X"50",X"07",X"A0",X"88",X"88",X"88",X"04",X"07",X"50",
		X"05",X"A0",X"40",X"40",X"38",X"05",X"06",X"46",X"05",X"A0",X"50",X"50",X"48",X"05",X"06",X"46",
		X"06",X"A0",X"58",X"58",X"48",X"07",X"06",X"46",X"0A",X"A0",X"90",X"90",X"90",X"06",X"06",X"46",
		X"06",X"A0",X"48",X"48",X"60",X"06",X"06",X"46",X"07",X"A0",X"70",X"70",X"68",X"06",X"06",X"46",
		X"07",X"A0",X"70",X"70",X"70",X"07",X"06",X"46",X"0A",X"A0",X"90",X"90",X"90",X"06",X"05",X"3C",
		X"08",X"A0",X"70",X"70",X"70",X"06",X"05",X"3C",X"08",X"A0",X"78",X"78",X"78",X"07",X"05",X"3C",
		X"08",X"A0",X"78",X"78",X"78",X"07",X"05",X"3C",X"0C",X"A0",X"98",X"98",X"98",X"20",X"02",X"20",
		X"02",X"50",X"02",X"C0",X"00",X"40",X"02",X"20",X"02",X"70",X"02",X"C0",X"00",X"60",X"02",X"40",
		X"02",X"90",X"02",X"C0",X"00",X"70",X"02",X"40",X"02",X"A0",X"02",X"C0",X"00",X"80",X"02",X"40",
		X"02",X"B0",X"02",X"C0",X"00",X"80",X"02",X"50",X"02",X"B0",X"02",X"C0",X"00",X"90",X"02",X"50",
		X"02",X"C0",X"02",X"C0",X"00",X"A0",X"02",X"50",X"02",X"D0",X"02",X"C0",X"00",X"B0",X"02",X"50",
		X"02",X"E0",X"02",X"C0",X"00",X"B0",X"02",X"60",X"02",X"E0",X"02",X"C0",X"00",X"C0",X"02",X"60",
		X"02",X"F0",X"02",X"C0",X"00",X"D0",X"02",X"60",X"02",X"F0",X"02",X"C0",X"00",X"A0",X"02",X"60",
		X"02",X"D0",X"02",X"C0",X"00",X"C0",X"02",X"70",X"02",X"F0",X"02",X"C0",X"00",X"D0",X"02",X"70",
		X"02",X"F0",X"02",X"C0",X"00",X"E0",X"02",X"70",X"02",X"F0",X"02",X"C0",X"00",X"00",X"00",X"A0",
		X"02",X"00",X"00",X"C0",X"00",X"00",X"00",X"B0",X"02",X"00",X"00",X"C0",X"00",X"00",X"00",X"C0",
		X"02",X"00",X"00",X"C0",X"00",X"00",X"00",X"D0",X"02",X"00",X"00",X"C0",X"00",X"00",X"03",X"20",
		X"02",X"00",X"03",X"C0",X"00",X"E5",X"24",X"E5",X"24",X"E5",X"24",X"E5",X"24",X"E5",X"24",X"C5",
		X"24",X"C5",X"24",X"CD",X"24",X"E5",X"24",X"C5",X"24",X"C5",X"24",X"C5",X"24",X"E5",X"24",X"C5",
		X"24",X"D5",X"24",X"DD",X"24",X"E5",X"24",X"E5",X"24",X"E5",X"24",X"E5",X"24",X"E5",X"24",X"CD",
		X"24",X"DD",X"24",X"FD",X"24",X"E5",X"24",X"ED",X"24",X"F5",X"24",X"FD",X"24",X"E5",X"24",X"E5",
		X"24",X"E5",X"24",X"E5",X"24",X"00",X"00",X"00",X"30",X"40",X"40",X"40",X"02",X"00",X"00",X"00",
		X"30",X"40",X"40",X"40",X"03",X"00",X"00",X"00",X"30",X"40",X"40",X"40",X"04",X"00",X"00",X"00",
		X"30",X"40",X"40",X"40",X"06",X"49",X"4E",X"47",X"40",X"4E",X"4F",X"54",X"48",X"00",X"00",X"00",
		X"30",X"40",X"40",X"40",X"08",X"00",X"00",X"00",X"30",X"40",X"40",X"01",X"00",X"00",X"00",X"00",
		X"30",X"40",X"40",X"01",X"02",X"40",X"80",X"08",X"40",X"40",X"FF",X"FF",X"40",X"00",X"04",X"20",
		X"40",X"40",X"FF",X"08",X"FF",X"40",X"FF",X"FF",X"FF",X"00",X"FF",X"20",X"FF",X"C0",X"01",X"08",
		X"10",X"80",X"FF",X"FF",X"10",X"80",X"02",X"20",X"10",X"90",X"91",X"92",X"93",X"90",X"91",X"92",
		X"80",X"80",X"40",X"04",X"08",X"00",X"20",X"01",X"10",X"02",X"F0",X"F4",X"F8",X"FC",X"FA",X"F6",
		X"F2",X"F7",X"FB",X"FD",X"F9",X"F5",X"F0",X"F4",X"F8",X"FC",X"FA",X"F6",X"F2",X"F7",X"FB",X"FD",
		X"F9",X"F5",X"E1",X"61",X"61",X"61",X"61",X"61",X"61",X"61",X"61",X"21",X"21",X"21",X"21",X"67",
		X"21",X"68",X"69",X"21",X"21",X"21",X"21",X"6A",X"67",X"21",X"68",X"69",X"21",X"54",X"55",X"56",
		X"57",X"58",X"59",X"5A",X"5B",X"5C",X"21",X"21",X"21",X"6B",X"67",X"21",X"68",X"69",X"21",X"06",
		X"3A",X"AE",X"8B",X"A7",X"CC",X"17",X"2B",X"CD",X"31",X"2B",X"21",X"F5",X"89",X"CB",X"46",X"28",
		X"07",X"21",X"AF",X"8B",X"36",X"00",X"18",X"02",X"CB",X"C6",X"21",X"F6",X"89",X"CB",X"7E",X"28",
		X"04",X"21",X"14",X"8A",X"34",X"CB",X"76",X"28",X"04",X"21",X"13",X"8A",X"34",X"21",X"28",X"8A",
		X"06",X"18",X"34",X"23",X"10",X"FC",X"3A",X"F5",X"89",X"CB",X"67",X"CA",X"5C",X"26",X"2A",X"8A",
		X"89",X"7E",X"E6",X"03",X"28",X"45",X"21",X"54",X"2B",X"3A",X"AF",X"8B",X"CD",X"F8",X"2A",X"7E",
		X"FE",X"FF",X"20",X"07",X"21",X"AF",X"8B",X"36",X"00",X"18",X"EB",X"21",X"A8",X"8B",X"77",X"3A",
		X"08",X"8A",X"A7",X"20",X"14",X"3C",X"32",X"08",X"8A",X"CD",X"D5",X"2A",X"36",X"00",X"23",X"36",
		X"00",X"CD",X"DF",X"2A",X"36",X"01",X"23",X"36",X"01",X"CD",X"15",X"2A",X"CD",X"52",X"2A",X"21",
		X"A8",X"8B",X"34",X"CD",X"28",X"2A",X"CD",X"52",X"2A",X"18",X"40",X"3A",X"AF",X"8B",X"CB",X"4F",
		X"20",X"04",X"3E",X"17",X"18",X"02",X"3E",X"0E",X"21",X"A8",X"8B",X"77",X"3A",X"08",X"8A",X"A7",
		X"20",X"18",X"3C",X"32",X"08",X"8A",X"CD",X"D5",X"2A",X"36",X"00",X"21",X"55",X"8A",X"36",X"00",
		X"CD",X"DF",X"2A",X"36",X"01",X"21",X"35",X"8A",X"36",X"01",X"CD",X"28",X"2A",X"CD",X"52",X"2A",
		X"21",X"A8",X"8B",X"36",X"0D",X"CD",X"15",X"2A",X"CD",X"52",X"2A",X"3A",X"A9",X"8B",X"A7",X"28",
		X"12",X"AF",X"32",X"A9",X"8B",X"32",X"08",X"8A",X"21",X"AF",X"8B",X"34",X"AF",X"32",X"08",X"8A",
		X"C3",X"AC",X"26",X"3A",X"F4",X"89",X"CB",X"77",X"28",X"42",X"21",X"A8",X"8B",X"36",X"02",X"CD",
		X"02",X"2A",X"21",X"69",X"80",X"FE",X"20",X"28",X"04",X"3E",X"00",X"18",X"02",X"3E",X"02",X"F5",
		X"CD",X"D5",X"2A",X"F1",X"77",X"CD",X"52",X"2A",X"3A",X"6A",X"80",X"CB",X"7F",X"20",X"0E",X"3A",
		X"6B",X"80",X"A7",X"28",X"04",X"3E",X"00",X"18",X"10",X"3E",X"01",X"18",X"0C",X"3A",X"6B",X"80",
		X"A7",X"28",X"04",X"3E",X"02",X"18",X"02",X"3E",X"03",X"32",X"97",X"8B",X"3A",X"F4",X"89",X"CB",
		X"67",X"28",X"36",X"21",X"A8",X"8B",X"36",X"05",X"3A",X"0B",X"8A",X"A7",X"20",X"0E",X"3C",X"32",
		X"0B",X"8A",X"CD",X"D5",X"2A",X"36",X"00",X"CD",X"DF",X"2A",X"36",X"01",X"CD",X"02",X"2A",X"CD",
		X"52",X"2A",X"3E",X"0F",X"32",X"94",X"8B",X"3A",X"A9",X"8B",X"A7",X"28",X"0C",X"AF",X"32",X"A9",
		X"8B",X"32",X"0B",X"8A",X"21",X"F4",X"89",X"CB",X"A6",X"21",X"F4",X"89",X"CB",X"56",X"28",X"16",
		X"CB",X"96",X"3E",X"01",X"32",X"09",X"8A",X"21",X"A8",X"8B",X"36",X"03",X"CD",X"D5",X"2A",X"36",
		X"00",X"CD",X"DF",X"2A",X"36",X"01",X"3A",X"09",X"8A",X"A7",X"28",X"18",X"21",X"A8",X"8B",X"36",
		X"03",X"CD",X"02",X"2A",X"CD",X"52",X"2A",X"3A",X"A9",X"8B",X"A7",X"28",X"07",X"AF",X"32",X"A9",
		X"8B",X"32",X"09",X"8A",X"3A",X"F4",X"89",X"CB",X"5F",X"28",X"31",X"21",X"A8",X"8B",X"36",X"04",
		X"3A",X"0A",X"8A",X"A7",X"20",X"0E",X"3C",X"32",X"0A",X"8A",X"CD",X"D5",X"2A",X"36",X"00",X"CD",
		X"DF",X"2A",X"36",X"01",X"CD",X"02",X"2A",X"CD",X"52",X"2A",X"3A",X"A9",X"8B",X"A7",X"28",X"0C",
		X"AF",X"32",X"A9",X"8B",X"32",X"0A",X"8A",X"21",X"F4",X"89",X"CB",X"9E",X"3A",X"F4",X"89",X"CB",
		X"6F",X"28",X"36",X"21",X"A8",X"8B",X"36",X"06",X"3A",X"0C",X"8A",X"A7",X"20",X"0E",X"3C",X"32",
		X"0C",X"8A",X"CD",X"D5",X"2A",X"36",X"00",X"CD",X"DF",X"2A",X"36",X"01",X"CD",X"02",X"2A",X"CD",
		X"52",X"2A",X"3E",X"0C",X"32",X"94",X"8B",X"3A",X"A9",X"8B",X"A7",X"28",X"0C",X"AF",X"32",X"A9",
		X"8B",X"32",X"0C",X"8A",X"21",X"F4",X"89",X"CB",X"AE",X"3A",X"F4",X"89",X"CB",X"47",X"28",X"36",
		X"21",X"A8",X"8B",X"36",X"07",X"3A",X"0D",X"8A",X"A7",X"20",X"0E",X"3C",X"32",X"0D",X"8A",X"CD",
		X"D5",X"2A",X"36",X"00",X"CD",X"DF",X"2A",X"36",X"01",X"CD",X"28",X"2A",X"CD",X"52",X"2A",X"3E",
		X"0C",X"32",X"94",X"8B",X"3A",X"A9",X"8B",X"A7",X"28",X"0C",X"AF",X"32",X"A9",X"8B",X"32",X"0D",
		X"8A",X"21",X"F4",X"89",X"CB",X"86",X"3A",X"F5",X"89",X"CB",X"6F",X"28",X"40",X"21",X"A8",X"8B",
		X"36",X"08",X"3A",X"0E",X"8A",X"A7",X"20",X"07",X"3C",X"32",X"0E",X"8A",X"CD",X"3B",X"2A",X"CD",
		X"02",X"2A",X"CD",X"52",X"2A",X"21",X"A8",X"8B",X"36",X"09",X"CD",X"15",X"2A",X"CD",X"52",X"2A",
		X"21",X"A8",X"8B",X"36",X"0A",X"CD",X"28",X"2A",X"CD",X"52",X"2A",X"3A",X"A9",X"8B",X"A7",X"28",
		X"0C",X"AF",X"32",X"A9",X"8B",X"32",X"0E",X"8A",X"21",X"F5",X"89",X"CB",X"AE",X"3A",X"F4",X"89",
		X"CB",X"4F",X"28",X"39",X"21",X"A8",X"8B",X"36",X"0B",X"3A",X"0F",X"8A",X"A7",X"20",X"11",X"3C",
		X"32",X"0F",X"8A",X"32",X"AD",X"8B",X"CD",X"D5",X"2A",X"36",X"00",X"CD",X"DF",X"2A",X"36",X"01",
		X"21",X"AC",X"8B",X"36",X"00",X"CD",X"02",X"2A",X"CD",X"52",X"2A",X"21",X"F4",X"89",X"CB",X"8E",
		X"3A",X"A9",X"8B",X"A7",X"28",X"07",X"AF",X"32",X"0F",X"8A",X"32",X"A9",X"8B",X"3A",X"AD",X"8B",
		X"A7",X"28",X"10",X"21",X"AC",X"8B",X"34",X"3E",X"06",X"BE",X"30",X"07",X"AF",X"32",X"AD",X"8B",
		X"32",X"0F",X"8A",X"3A",X"F5",X"89",X"CB",X"77",X"28",X"31",X"21",X"A8",X"8B",X"36",X"0F",X"3A",
		X"10",X"8A",X"A7",X"20",X"08",X"3E",X"02",X"32",X"10",X"8A",X"CD",X"3B",X"2A",X"CD",X"02",X"2A",
		X"CD",X"52",X"2A",X"3A",X"A9",X"8B",X"A7",X"28",X"12",X"AF",X"32",X"A9",X"8B",X"CD",X"3B",X"2A",
		X"21",X"10",X"8A",X"35",X"20",X"05",X"21",X"F5",X"89",X"CB",X"B6",X"3A",X"F4",X"89",X"CB",X"7F",
		X"28",X"0F",X"21",X"80",X"A1",X"3E",X"FF",X"77",X"3D",X"20",X"FC",X"77",X"21",X"F4",X"89",X"CB",
		X"BE",X"3A",X"F5",X"89",X"CB",X"7F",X"28",X"40",X"21",X"A8",X"8B",X"36",X"12",X"3A",X"11",X"8A",
		X"A7",X"20",X"07",X"3C",X"32",X"11",X"8A",X"CD",X"3B",X"2A",X"CD",X"02",X"2A",X"CD",X"52",X"2A",
		X"21",X"A8",X"8B",X"36",X"13",X"CD",X"15",X"2A",X"CD",X"52",X"2A",X"21",X"A8",X"8B",X"36",X"14",
		X"CD",X"28",X"2A",X"CD",X"52",X"2A",X"3A",X"A9",X"8B",X"A7",X"28",X"0C",X"AF",X"32",X"A9",X"8B",
		X"32",X"11",X"8A",X"21",X"F5",X"89",X"CB",X"BE",X"3A",X"F5",X"89",X"CB",X"57",X"CA",X"46",X"29",
		X"21",X"A8",X"8B",X"36",X"15",X"3A",X"12",X"8A",X"A7",X"20",X"07",X"3C",X"32",X"12",X"8A",X"CD",
		X"3B",X"2A",X"CD",X"02",X"2A",X"CD",X"52",X"2A",X"21",X"A8",X"8B",X"36",X"16",X"CD",X"15",X"2A",
		X"CD",X"52",X"2A",X"3A",X"A9",X"8B",X"A7",X"CA",X"46",X"29",X"AF",X"32",X"A9",X"8B",X"32",X"12",
		X"8A",X"21",X"F5",X"89",X"CB",X"96",X"AF",X"32",X"F6",X"89",X"3A",X"14",X"8A",X"A7",X"28",X"36",
		X"21",X"A8",X"8B",X"36",X"00",X"3A",X"16",X"8A",X"A7",X"20",X"0E",X"3C",X"32",X"16",X"8A",X"CD",
		X"D5",X"2A",X"36",X"00",X"CD",X"DF",X"2A",X"36",X"01",X"CD",X"02",X"2A",X"CD",X"52",X"2A",X"21",
		X"29",X"8A",X"35",X"3A",X"A9",X"8B",X"A7",X"28",X"43",X"AF",X"32",X"A9",X"8B",X"32",X"16",X"8A",
		X"21",X"14",X"8A",X"35",X"18",X"36",X"3A",X"13",X"8A",X"A7",X"28",X"30",X"21",X"A8",X"8B",X"36",
		X"01",X"3A",X"15",X"8A",X"A7",X"20",X"0E",X"3C",X"32",X"15",X"8A",X"CD",X"D5",X"2A",X"36",X"00",
		X"CD",X"DF",X"2A",X"36",X"01",X"CD",X"02",X"2A",X"CD",X"52",X"2A",X"3A",X"A9",X"8B",X"A7",X"28",
		X"0B",X"AF",X"32",X"A9",X"8B",X"32",X"15",X"8A",X"21",X"13",X"8A",X"35",X"21",X"88",X"8B",X"11",
		X"11",X"A1",X"01",X"04",X"00",X"ED",X"B0",X"3A",X"94",X"8B",X"32",X"15",X"A1",X"3A",X"97",X"8B",
		X"32",X"05",X"A1",X"21",X"8C",X"8B",X"11",X"16",X"A1",X"01",X"04",X"00",X"ED",X"B0",X"3A",X"95",
		X"8B",X"32",X"1A",X"A1",X"3A",X"98",X"8B",X"32",X"0A",X"A1",X"21",X"90",X"8B",X"11",X"1B",X"A1",
		X"01",X"04",X"00",X"ED",X"B0",X"3A",X"96",X"8B",X"32",X"1F",X"A1",X"3A",X"99",X"8B",X"32",X"0F",
		X"A1",X"C9",X"21",X"97",X"8B",X"22",X"9E",X"8B",X"21",X"88",X"8B",X"22",X"9A",X"8B",X"21",X"94",
		X"8B",X"22",X"9C",X"8B",X"C9",X"21",X"98",X"8B",X"22",X"9E",X"8B",X"21",X"8C",X"8B",X"22",X"9A",
		X"8B",X"21",X"95",X"8B",X"22",X"9C",X"8B",X"C9",X"21",X"99",X"8B",X"22",X"9E",X"8B",X"21",X"90",
		X"8B",X"22",X"9A",X"8B",X"21",X"96",X"8B",X"22",X"9C",X"8B",X"C9",X"CD",X"D5",X"2A",X"36",X"00",
		X"23",X"36",X"00",X"23",X"36",X"00",X"CD",X"DF",X"2A",X"36",X"01",X"23",X"36",X"01",X"23",X"36",
		X"01",X"C9",X"21",X"F5",X"89",X"CB",X"86",X"3A",X"A8",X"8B",X"21",X"58",X"2B",X"CD",X"F4",X"2A",
		X"5E",X"23",X"56",X"CD",X"D5",X"2A",X"7E",X"EB",X"CD",X"F8",X"2A",X"7E",X"FE",X"FF",X"CA",X"E9",
		X"2A",X"E6",X"0F",X"EB",X"21",X"FD",X"2A",X"CD",X"F4",X"2A",X"4E",X"23",X"46",X"EB",X"7E",X"E6",
		X"F0",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"A7",X"28",X"05",X"CB",X"38",X"CB",X"19",
		X"3D",X"20",X"F9",X"ED",X"5B",X"9A",X"8B",X"79",X"12",X"0F",X"0F",X"0F",X"0F",X"13",X"12",X"78",
		X"13",X"12",X"0F",X"0F",X"0F",X"0F",X"13",X"12",X"EB",X"CD",X"DF",X"2A",X"4E",X"EB",X"3E",X"08",
		X"ED",X"5B",X"9C",X"8B",X"12",X"E5",X"21",X"68",X"8A",X"3A",X"A8",X"8B",X"CD",X"F8",X"2A",X"7E",
		X"ED",X"5B",X"9E",X"8B",X"12",X"E1",X"79",X"23",X"BE",X"D8",X"CD",X"D5",X"2A",X"34",X"34",X"CD",
		X"DF",X"2A",X"36",X"00",X"C9",X"21",X"48",X"8A",X"3A",X"A8",X"8B",X"CD",X"F8",X"2A",X"C9",X"21",
		X"28",X"8A",X"3A",X"A8",X"8B",X"CD",X"F8",X"2A",X"C9",X"2A",X"9C",X"8B",X"36",X"00",X"3E",X"01",
		X"32",X"A9",X"8B",X"C9",X"87",X"30",X"01",X"24",X"85",X"6F",X"D0",X"24",X"C9",X"50",X"81",X"00",
		X"89",X"26",X"91",X"C8",X"99",X"EC",X"A2",X"9D",X"AC",X"E0",X"B6",X"C0",X"C1",X"45",X"CD",X"7A",
		X"D9",X"69",X"E6",X"1C",X"F4",X"00",X"00",X"21",X"3C",X"2B",X"11",X"68",X"8A",X"01",X"18",X"00",
		X"ED",X"B0",X"3E",X"01",X"32",X"AE",X"8B",X"21",X"08",X"8A",X"06",X"18",X"36",X"00",X"23",X"10",
		X"FB",X"AF",X"32",X"94",X"8B",X"32",X"95",X"8B",X"32",X"96",X"8B",X"C9",X"06",X"07",X"00",X"07",
		X"07",X"04",X"07",X"07",X"07",X"07",X"07",X"07",X"00",X"07",X"07",X"04",X"07",X"07",X"06",X"05",
		X"07",X"04",X"07",X"07",X"10",X"0D",X"0D",X"FF",X"05",X"2D",X"FC",X"2C",X"6F",X"2C",X"8E",X"2C",
		X"72",X"2C",X"9D",X"2C",X"A6",X"2C",X"BD",X"2C",X"D6",X"2C",X"D8",X"2C",X"DA",X"2C",X"EB",X"2C",
		X"00",X"00",X"88",X"2B",X"09",X"2C",X"0E",X"2D",X"45",X"2D",X"42",X"2E",X"D4",X"2E",X"06",X"2F",
		X"26",X"2F",X"4B",X"2F",X"BB",X"2F",X"39",X"2C",X"93",X"08",X"0C",X"04",X"93",X"08",X"0C",X"04",
		X"83",X"08",X"0C",X"04",X"83",X"08",X"0C",X"04",X"93",X"08",X"0C",X"04",X"93",X"08",X"0C",X"04",
		X"83",X"08",X"0C",X"04",X"83",X"08",X"0C",X"04",X"93",X"08",X"0C",X"04",X"93",X"08",X"0C",X"04",
		X"83",X"08",X"0C",X"04",X"83",X"08",X"0C",X"04",X"93",X"08",X"0C",X"04",X"93",X"08",X"0C",X"04",
		X"83",X"08",X"0C",X"04",X"83",X"08",X"0C",X"04",X"A8",X"08",X"0C",X"04",X"A8",X"08",X"0C",X"04",
		X"98",X"08",X"0C",X"04",X"98",X"08",X"0C",X"04",X"A8",X"08",X"0C",X"04",X"A8",X"08",X"0C",X"04",
		X"98",X"08",X"0C",X"04",X"98",X"08",X"0C",X"04",X"93",X"08",X"0C",X"04",X"93",X"08",X"0C",X"04",
		X"83",X"08",X"0C",X"04",X"83",X"08",X"0C",X"04",X"93",X"08",X"0C",X"04",X"93",X"08",X"0C",X"04",
		X"83",X"08",X"0C",X"04",X"83",X"08",X"0C",X"04",X"FF",X"7A",X"18",X"77",X"0C",X"7A",X"0C",X"60",
		X"0C",X"77",X"0C",X"7A",X"0C",X"60",X"0C",X"77",X"0C",X"75",X"0C",X"73",X"0C",X"70",X"0C",X"73",
		X"30",X"70",X"0C",X"73",X"0C",X"75",X"0C",X"73",X"0C",X"77",X"0C",X"75",X"0C",X"73",X"0C",X"75",
		X"0C",X"77",X"0C",X"73",X"18",X"70",X"0C",X"8A",X"30",X"73",X"0C",X"71",X"0C",X"8A",X"0C",X"73",
		X"0C",X"72",X"0C",X"8A",X"0C",X"88",X"0C",X"8A",X"0C",X"88",X"0C",X"86",X"0C",X"83",X"0C",X"88",
		X"0C",X"87",X"0C",X"83",X"24",X"88",X"0C",X"86",X"0C",X"83",X"0C",X"81",X"0C",X"83",X"0C",X"86",
		X"0C",X"88",X"0C",X"89",X"0C",X"8A",X"0C",X"72",X"0C",X"8A",X"0C",X"88",X"0C",X"87",X"30",X"A1",
		X"04",X"A6",X"78",X"02",X"7B",X"02",X"61",X"02",X"63",X"02",X"66",X"02",X"68",X"02",X"6B",X"02",
		X"78",X"02",X"7B",X"02",X"61",X"02",X"63",X"02",X"66",X"02",X"68",X"02",X"6B",X"02",X"7B",X"02",
		X"61",X"02",X"63",X"02",X"66",X"02",X"68",X"02",X"6B",X"02",X"51",X"02",X"FF",X"96",X"01",X"97",
		X"01",X"98",X"01",X"99",X"01",X"FF",X"89",X"0C",X"0C",X"03",X"89",X"0C",X"0C",X"03",X"89",X"0C",
		X"0C",X"03",X"89",X"0C",X"0C",X"03",X"89",X"0C",X"0C",X"03",X"89",X"0C",X"FF",X"68",X"04",X"6A",
		X"04",X"68",X"04",X"6A",X"04",X"68",X"04",X"6A",X"04",X"68",X"04",X"6A",X"04",X"68",X"04",X"6A",
		X"04",X"68",X"04",X"6A",X"04",X"FF",X"0C",X"08",X"0C",X"08",X"76",X"0C",X"7A",X"0C",X"61",X"0C",
		X"78",X"0C",X"7B",X"0C",X"7A",X"0C",X"66",X"12",X"0C",X"10",X"FF",X"63",X"01",X"65",X"05",X"67",
		X"05",X"68",X"05",X"6A",X"05",X"50",X"05",X"52",X"05",X"53",X"05",X"FF",X"79",X"04",X"61",X"04",
		X"7B",X"04",X"62",X"04",X"FF",X"64",X"04",X"61",X"04",X"63",X"04",X"7B",X"04",X"FF",X"93",X"0C",
		X"AA",X"06",X"91",X"06",X"93",X"06",X"96",X"06",X"98",X"06",X"9A",X"06",X"83",X"06",X"81",X"06",
		X"83",X"06",X"0C",X"06",X"86",X"0C",X"83",X"06",X"81",X"06",X"93",X"0C",X"AA",X"06",X"91",X"06",
		X"93",X"06",X"96",X"06",X"98",X"06",X"9A",X"06",X"83",X"06",X"81",X"06",X"99",X"06",X"9A",X"06",
		X"97",X"0C",X"0C",X"0C",X"FF",X"93",X"08",X"0C",X"04",X"93",X"08",X"0C",X"04",X"83",X"08",X"0C",
		X"04",X"83",X"08",X"0C",X"04",X"93",X"08",X"0C",X"04",X"93",X"08",X"0C",X"04",X"83",X"08",X"0C",
		X"04",X"83",X"08",X"0C",X"04",X"93",X"08",X"0C",X"04",X"93",X"08",X"0C",X"04",X"83",X"08",X"0C",
		X"04",X"83",X"08",X"0C",X"04",X"93",X"08",X"0C",X"04",X"93",X"08",X"0C",X"04",X"83",X"08",X"0C",
		X"04",X"83",X"08",X"0C",X"04",X"93",X"08",X"0C",X"04",X"93",X"08",X"0C",X"04",X"83",X"08",X"0C",
		X"04",X"83",X"08",X"0C",X"04",X"93",X"08",X"0C",X"04",X"93",X"08",X"0C",X"04",X"83",X"08",X"0C",
		X"04",X"83",X"08",X"0C",X"04",X"AA",X"08",X"0C",X"04",X"AA",X"08",X"0C",X"04",X"9A",X"08",X"0C",
		X"04",X"9A",X"08",X"0C",X"04",X"9A",X"08",X"0C",X"04",X"AA",X"08",X"0C",X"04",X"90",X"08",X"0C",
		X"04",X"92",X"08",X"0C",X"04",X"93",X"08",X"0C",X"04",X"93",X"08",X"0C",X"04",X"83",X"08",X"0C",
		X"04",X"83",X"08",X"0C",X"04",X"93",X"08",X"0C",X"04",X"93",X"08",X"0C",X"04",X"83",X"08",X"0C",
		X"04",X"83",X"08",X"0C",X"04",X"93",X"08",X"0C",X"04",X"93",X"08",X"0C",X"04",X"83",X"08",X"0C",
		X"04",X"83",X"08",X"0C",X"04",X"93",X"08",X"0C",X"04",X"93",X"08",X"0C",X"04",X"83",X"08",X"0C",
		X"04",X"83",X"08",X"0C",X"04",X"93",X"08",X"0C",X"04",X"93",X"08",X"0C",X"04",X"83",X"08",X"0C",
		X"04",X"83",X"08",X"0C",X"04",X"93",X"08",X"0C",X"04",X"93",X"08",X"0C",X"04",X"83",X"08",X"0C",
		X"04",X"83",X"08",X"0C",X"04",X"A8",X"09",X"0C",X"04",X"98",X"08",X"0C",X"04",X"AA",X"09",X"0C",
		X"04",X"9A",X"08",X"0C",X"04",X"93",X"08",X"0C",X"04",X"83",X"08",X"0C",X"04",X"83",X"0C",X"0C",
		X"0C",X"FF",X"73",X"0A",X"0C",X"02",X"73",X"0C",X"70",X"0C",X"8A",X"0C",X"73",X"0C",X"0C",X"0C",
		X"76",X"18",X"73",X"0A",X"0C",X"02",X"73",X"0C",X"70",X"0C",X"8A",X"0C",X"73",X"0C",X"0C",X"0C",
		X"70",X"18",X"73",X"0A",X"0C",X"02",X"73",X"0C",X"70",X"0C",X"8A",X"0C",X"73",X"0C",X"76",X"0C",
		X"78",X"0C",X"79",X"0C",X"7A",X"0C",X"79",X"06",X"7A",X"06",X"79",X"06",X"7A",X"06",X"79",X"06",
		X"7A",X"04",X"0C",X"02",X"7A",X"14",X"0C",X"04",X"7A",X"06",X"78",X"06",X"77",X"06",X"75",X"06",
		X"73",X"0A",X"0C",X"02",X"73",X"0C",X"70",X"0C",X"8A",X"0C",X"73",X"0C",X"0C",X"0C",X"76",X"18",
		X"73",X"0A",X"0C",X"02",X"73",X"0C",X"70",X"0C",X"8A",X"0C",X"73",X"0C",X"0C",X"0C",X"70",X"18",
		X"73",X"0A",X"0C",X"02",X"73",X"0C",X"70",X"0C",X"8A",X"0C",X"73",X"0C",X"76",X"0C",X"78",X"0C",
		X"79",X"0C",X"63",X"0C",X"7A",X"06",X"78",X"06",X"76",X"0C",X"73",X"0C",X"71",X"0C",X"72",X"0C",
		X"73",X"0C",X"0C",X"0C",X"78",X"0C",X"7A",X"04",X"61",X"0C",X"65",X"10",X"61",X"04",X"7A",X"10",
		X"78",X"0C",X"7A",X"04",X"61",X"0C",X"64",X"10",X"61",X"04",X"7A",X"10",X"78",X"0C",X"7A",X"04",
		X"61",X"0C",X"65",X"10",X"61",X"04",X"65",X"0C",X"66",X"04",X"68",X"0C",X"66",X"04",X"64",X"0C",
		X"61",X"04",X"64",X"0C",X"61",X"04",X"78",X"1C",X"75",X"10",X"71",X"14",X"78",X"1C",X"74",X"10",
		X"71",X"14",X"78",X"1C",X"75",X"10",X"71",X"10",X"78",X"04",X"74",X"0C",X"71",X"04",X"8B",X"0C",
		X"88",X"04",X"70",X"0C",X"71",X"04",X"91",X"10",X"81",X"10",X"91",X"10",X"81",X"10",X"91",X"10",
		X"81",X"10",X"91",X"10",X"81",X"10",X"91",X"10",X"81",X"10",X"91",X"10",X"81",X"10",X"A6",X"0C",
		X"96",X"04",X"A8",X"0C",X"98",X"04",X"91",X"0C",X"81",X"04",X"FF",X"88",X"10",X"85",X"0C",X"88",
		X"04",X"71",X"10",X"88",X"0C",X"85",X"04",X"86",X"0A",X"0C",X"02",X"86",X"03",X"0C",X"01",X"86",
		X"0C",X"85",X"04",X"86",X"10",X"0C",X"10",X"86",X"10",X"83",X"0C",X"86",X"04",X"70",X"10",X"8A",
		X"0C",X"88",X"04",X"85",X"0A",X"0C",X"02",X"85",X"03",X"0C",X"01",X"85",X"0C",X"84",X"04",X"85",
		X"10",X"0C",X"10",X"81",X"10",X"85",X"0C",X"88",X"04",X"71",X"10",X"88",X"0C",X"85",X"04",X"86",
		X"0A",X"0C",X"02",X"86",X"03",X"0C",X"01",X"86",X"0C",X"88",X"04",X"8A",X"10",X"0C",X"10",X"8A",
		X"0A",X"0C",X"02",X"8A",X"04",X"73",X"0C",X"71",X"04",X"70",X"0C",X"71",X"04",X"88",X"0C",X"85",
		X"04",X"88",X"0C",X"86",X"04",X"85",X"0C",X"83",X"04",X"81",X"10",X"81",X"10",X"88",X"10",X"81",
		X"10",X"88",X"10",X"80",X"10",X"88",X"10",X"80",X"10",X"88",X"10",X"80",X"10",X"86",X"10",X"83",
		X"10",X"80",X"10",X"81",X"10",X"85",X"0C",X"86",X"04",X"88",X"10",X"98",X"10",X"81",X"10",X"88",
		X"10",X"81",X"10",X"88",X"10",X"86",X"10",X"71",X"10",X"86",X"10",X"71",X"10",X"86",X"10",X"8A",
		X"10",X"88",X"10",X"81",X"10",X"83",X"10",X"98",X"10",X"81",X"10",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"01",X"FE",X"00",X"77",X"D8",X"1E",X"FE",X"77",X"D8",X"9E",X"00",X"00",X"00",X"80",X"EE",
		X"7E",X"F8",X"1E",X"EE",X"00",X"01",X"DE",X"00",X"0F",X"D7",X"DE",X"FE",X"20",X"57",X"00",X"00",
		X"2F",X"57",X"77",X"FD",X"28",X"57",X"70",X"05",X"2B",X"50",X"74",X"05",X"2B",X"57",X"75",X"F5",
		X"68",X"57",X"75",X"F5",X"6B",X"D0",X"04",X"05",X"08",X"17",X"67",X"3D",X"6B",X"F7",X"67",X"3D",
		X"60",X"07",X"67",X"3D",X"7F",X"F7",X"00",X"01",X"03",X"00",X"00",X"3B",X"7B",X"7F",X"3F",X"3B",
		X"78",X"07",X"3F",X"03",X"7B",X"77",X"03",X"39",X"03",X"70",X"33",X"39",X"BF",X"7F",X"33",X"3D",
		X"80",X"00",X"30",X"01",X"BF",X"7F",X"3F",X"3D",X"BF",X"7F",X"3F",X"3D",X"80",X"00",X"00",X"01",
		X"BB",X"7B",X"3B",X"3D",X"BB",X"7B",X"3B",X"3D",X"BB",X"60",X"03",X"31",X"BB",X"6B",X"3B",X"35",
		X"80",X"03",X"38",X"35",X"B7",X"7B",X"03",X"04",X"37",X"7B",X"3B",X"3E",X"00",X"1B",X"3B",X"3E",
		X"3D",X"C0",X"00",X"00",X"3D",X"C0",X"00",X"00",X"00",X"76",X"EF",X"36",X"37",X"76",X"EF",X"36",
		X"37",X"70",X"0F",X"36",X"37",X"76",X"E0",X"30",X"30",X"06",X"0B",X"36",X"37",X"DE",X"EB",X"36",
		X"37",X"DE",X"EB",X"36",X"00",X"00",X"08",X"06",X"DD",X"BE",X"EB",X"36",X"DD",X"BE",X"EB",X"36",
		X"C0",X"00",X"03",X"36",X"DD",X"AA",X"AB",X"36",X"DD",X"AA",X"AB",X"00",X"0C",X"2A",X"A8",X"3E",
		X"61",X"AA",X"AB",X"3E",X"6F",X"AA",X"AB",X"06",X"6F",X"AA",X"AB",X"36",X"00",X"00",X"00",X"30",
		X"0B",X"05",X"17",X"05",X"17",X"05",X"15",X"09",X"15",X"09",X"01",X"0E",X"01",X"0E",X"05",X"0F",
		X"18",X"11",X"18",X"11",X"06",X"14",X"14",X"16",X"11",X"1B",X"0B",X"20",X"01",X"23",X"1C",X"2B",
		X"FF",X"F8",X"00",X"00",X"80",X"0A",X"AF",X"DE",X"BD",X"EA",X"AF",X"DE",X"A0",X"2A",X"A0",X"02",
		X"AD",X"AA",X"AE",X"DA",X"A8",X"AA",X"AE",X"DA",X"A8",X"A8",X"00",X"00",X"AA",X"AA",X"DB",X"FA",
		X"AA",X"AA",X"DA",X"02",X"8A",X"82",X"DA",X"FA",X"AA",X"AA",X"DA",X"82",X"A8",X"A8",X"00",X"3A",
		X"A8",X"AA",X"DA",X"82",X"AD",X"AA",X"DA",X"FA",X"A0",X"2A",X"DA",X"02",X"BD",X"EA",X"DB",X"FA",
		X"80",X"08",X"00",X"00",X"FD",X"FA",X"DB",X"7A",X"00",X"02",X"DB",X"7A",X"AD",X"EE",X"C0",X"02",
		X"AD",X"EE",X"FB",X"DA",X"AD",X"EE",X"FB",X"DA",X"AD",X"EE",X"FB",X"DA",X"20",X"00",X"03",X"DA",
		X"2E",X"F7",X"E0",X"00",X"2E",X"C1",X"00",X"00",X"20",X"DD",X"7B",X"BE",X"2E",X"DD",X"7B",X"BE",
		X"2E",X"DC",X"7B",X"BE",X"00",X"00",X"71",X"B0",X"2E",X"7C",X"75",X"B6",X"2E",X"7C",X"75",X"B6",
		X"28",X"1C",X"00",X"06",X"08",X"1C",X"75",X"B6",X"29",X"9C",X"75",X"B6",X"29",X"9C",X"71",X"B0",
		X"28",X"00",X"7B",X"BE",X"2F",X"EC",X"7B",X"BE",X"00",X"0C",X"78",X"00",X"6D",X"AC",X"7B",X"FE",
		X"6D",X"A0",X"03",X"00",X"00",X"0E",X"DB",X"76",X"6D",X"AE",X"18",X"06",X"6D",X"AE",X"FB",X"FE",
		X"00",X"20",X"00",X"00",X"6D",X"AE",X"EF",X"BB",X"6D",X"AE",X"EF",X"BB",X"00",X"00",X"03",X"BB",
		X"EF",X"6A",X"A8",X"00",X"EF",X"2A",X"AB",X"BE",X"EF",X"AA",X"A8",X"00",X"01",X"AA",X"AB",X"F6",
		X"6D",X"AA",X"AA",X"06",X"6C",X"00",X"02",X"F6",X"6D",X"BE",X"FA",X"F6",X"00",X"00",X"00",X"00",
		X"18",X"03",X"16",X"0B",X"1F",X"0B",X"14",X"10",X"14",X"10",X"01",X"18",X"01",X"18",X"16",X"20",
		X"16",X"20",X"1F",X"20",X"0C",X"24",X"1A",X"28",X"03",X"29",X"17",X"30",X"07",X"35",X"07",X"35",
		X"00",X"00",X"0E",X"00",X"3F",X"7A",X"AE",X"EE",X"20",X"7A",X"A0",X"E0",X"20",X"7A",X"AE",X"EE",
		X"20",X"02",X"AE",X"0E",X"3F",X"DA",X"AF",X"BE",X"0F",X"D8",X"0F",X"BE",X"2F",X"DE",X"E0",X"00",
		X"20",X"00",X"EF",X"B2",X"2D",X"DE",X"EF",X"B2",X"2D",X"DE",X"00",X"32",X"01",X"DE",X"AF",X"B2",
		X"7D",X"DE",X"AF",X"B2",X"7D",X"C0",X"AF",X"B0",X"7D",X"DE",X"AC",X"02",X"7D",X"DE",X"2D",X"F2",
		X"00",X"1E",X"AD",X"F2",X"7D",X"DE",X"AD",X"F2",X"7D",X"DE",X"AD",X"F2",X"7D",X"C0",X"00",X"00",
		X"7D",X"F6",X"0F",X"6C",X"60",X"37",X"FF",X"6C",X"67",X"34",X"01",X"6D",X"07",X"05",X"9D",X"6D",
		X"60",X"34",X"01",X"61",X"7D",X"F5",X"9D",X"7D",X"7D",X"F4",X"01",X"7D",X"7D",X"F7",X"9F",X"01",
		X"00",X"07",X"9F",X"7D",X"00",X"07",X"9F",X"7D",X"6D",X"B0",X"00",X"00",X"6D",X"B0",X"00",X"00",
		X"6D",X"B7",X"DE",X"FE",X"0D",X"87",X"DE",X"FE",X"7D",X"EF",X"DE",X"1E",X"7D",X"EF",X"06",X"DE",
		X"00",X"00",X"76",X"C6",X"7D",X"EF",X"70",X"F6",X"7D",X"EF",X"06",X"F0",X"0D",X"8F",X"76",X"FE",
		X"6D",X"B8",X"76",X"FE",X"6D",X"83",X"00",X"00",X"6D",X"B7",X"7B",X"DE",X"60",X"37",X"7B",X"DE",
		X"7D",X"80",X"1B",X"DE",X"7D",X"AE",X"D8",X"00",X"00",X"2E",X"DB",X"FE",X"7F",X"A0",X"00",X"00",
		X"7F",X"AA",X"AB",X"BE",X"70",X"2A",X"AA",X"20",X"77",X"AA",X"AA",X"AA",X"07",X"AA",X"AA",X"AA",
		X"7F",X"AA",X"AA",X"AA",X"70",X"00",X"02",X"82",X"77",X"BF",X"BA",X"FA",X"00",X"00",X"00",X"00",
		X"1B",X"02",X"08",X"03",X"08",X"03",X"0C",X"08",X"00",X"0A",X"1E",X"0D",X"11",X"0E",X"11",X"0E",
		X"06",X"13",X"1E",X"14",X"0C",X"21",X"0C",X"21",X"14",X"25",X"14",X"25",X"1C",X"2D",X"07",X"2E",
		X"00",X"00",X"00",X"00",X"7F",X"78",X"1D",X"FE",X"1F",X"78",X"1D",X"FE",X"4F",X"78",X"1C",X"00",
		X"67",X"7A",X"5E",X"F4",X"70",X"1A",X"5E",X"F4",X"7B",X"DA",X"5E",X"F4",X"7B",X"82",X"40",X"74",
		X"7B",X"BA",X"5F",X"74",X"7B",X"9A",X"5F",X"74",X"03",X"DA",X"5F",X"74",X"77",X"D8",X"1F",X"04",
		X"70",X"1E",X"7F",X"B4",X"7D",X"DE",X"7F",X"B4",X"7D",X"D0",X"0F",X"B4",X"7D",X"D0",X"0F",X"B0",
		X"7D",X"D3",X"CF",X"BC",X"00",X"03",X"C0",X"00",X"00",X"03",X"C0",X"5E",X"DD",X"F3",X"CD",X"1E",
		X"DD",X"F0",X"0D",X"DE",X"DD",X"F0",X"08",X"42",X"00",X"1E",X"7B",X"7A",X"DD",X"DE",X"63",X"00",
		X"DD",X"DE",X"6F",X"DA",X"DD",X"DE",X"6E",X"1A",X"C0",X"00",X"6E",X"FA",X"DD",X"D6",X"6E",X"FA",
		X"DD",X"D6",X"6E",X"FA",X"0D",X"D6",X"6E",X"FA",X"60",X"00",X"00",X"F0",X"60",X"0E",X"6E",X"F6",
		X"6F",X"EE",X"6E",X"F0",X"20",X"2E",X"6E",X"F7",X"27",X"2E",X"6C",X"37",X"20",X"2E",X"6D",X"87",
		X"2F",X"20",X"6D",X"BF",X"01",X"2E",X"01",X"BF",X"2D",X"2E",X"6C",X"00",X"2D",X"2E",X"6D",X"BE",
		X"25",X"2E",X"6D",X"B8",X"35",X"2E",X"60",X"3A",X"35",X"2E",X"6D",X"BA",X"71",X"2E",X"6D",X"80",
		X"7D",X"2E",X"6F",X"BE",X"7D",X"2E",X"6F",X"A2",X"40",X"00",X"00",X"0A",X"55",X"2A",X"AB",X"6A",
		X"55",X"2A",X"AB",X"6A",X"15",X"2A",X"AB",X"62",X"75",X"2A",X"AB",X"6A",X"05",X"2A",X"AB",X"6A",
		X"7D",X"20",X"03",X"6A",X"7D",X"2F",X"FB",X"60",X"01",X"20",X"00",X"7E",X"00",X"00",X"00",X"00",
		X"1F",X"04",X"1F",X"04",X"1F",X"0F",X"18",X"11",X"18",X"11",X"06",X"14",X"10",X"16",X"10",X"16",
		X"0B",X"1E",X"0F",X"21",X"00",X"22",X"08",X"23",X"08",X"23",X"17",X"26",X"17",X"36",X"05",X"37",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"01",X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",X"F7",X"07",X"FF",
		X"FF",X"F7",X"77",X"FF",X"FF",X"F7",X"77",X"FF",X"FF",X"F0",X"77",X"FF",X"FF",X"F7",X"77",X"FF",
		X"FF",X"F7",X"77",X"FF",X"FF",X"F0",X"07",X"FF",X"FF",X"F7",X"7F",X"FF",X"FF",X"F7",X"7F",X"FF",
		X"FF",X"F7",X"7F",X"FF",X"FF",X"F7",X"00",X"3F",X"FF",X"00",X"00",X"3F",X"FF",X"7F",X"3F",X"3F",
		X"F8",X"7F",X"FF",X"3F",X"FB",X"7F",X"07",X"3F",X"83",X"7F",X"37",X"3F",X"BF",X"7F",X"33",X"3F",
		X"80",X"00",X"30",X"01",X"FF",X"FF",X"3F",X"FD",X"FF",X"FF",X"3F",X"FD",X"FF",X"00",X"03",X"81",
		X"FF",X"7F",X"FB",X"BD",X"FF",X"7F",X"FB",X"BD",X"FF",X"60",X"7B",X"BD",X"FF",X"6F",X"7B",X"BD",
		X"87",X"0F",X"78",X"3D",X"B7",X"FF",X"7F",X"BC",X"37",X"FF",X"7F",X"BE",X"70",X"1F",X"7F",X"FE",
		X"7F",X"C0",X"00",X"06",X"7F",X"FF",X"00",X"30",X"7F",X"FF",X"FF",X"B6",X"7F",X"FF",X"FF",X"B6",
		X"7F",X"FF",X"FF",X"B6",X"7F",X"FF",X"FF",X"B0",X"7F",X"FF",X"FF",X"BF",X"7F",X"FF",X"FF",X"BF",
		X"7F",X"FF",X"FF",X"BF",X"00",X"00",X"FF",X"87",X"FD",X"FE",X"FF",X"F7",X"FD",X"FE",X"FF",X"F7",
		X"FD",X"80",X"0F",X"F7",X"FD",X"BE",X"EF",X"F7",X"FD",X"BE",X"EF",X"F0",X"FD",X"BF",X"EF",X"FE",
		X"E1",X"BF",X"EF",X"FE",X"EF",X"BF",X"EF",X"86",X"EF",X"BF",X"EF",X"B6",X"E0",X"3F",X"E0",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"00",X"1F",X"00",X"0C",X"08",X"05",X"0A",X"1C",X"0B",X"09",X"10",X"0C",X"15",X"18",X"18",
		X"08",X"1B",X"1C",X"1F",X"10",X"20",X"05",X"26",X"0C",X"28",X"16",X"29",X"1F",X"2D",X"01",X"33",
		X"17",X"00",X"01",X"01",X"11",X"05",X"07",X"09",X"0A",X"09",X"19",X"0B",X"17",X"13",X"1F",X"14",
		X"09",X"17",X"15",X"1D",X"01",X"1E",X"05",X"24",X"06",X"26",X"1C",X"2C",X"03",X"33",X"19",X"34",
		X"19",X"00",X"01",X"01",X"04",X"03",X"17",X"0A",X"1F",X"10",X"11",X"14",X"0E",X"16",X"03",X"18",
		X"12",X"1B",X"1B",X"1F",X"06",X"20",X"1B",X"24",X"12",X"29",X"18",X"2D",X"06",X"31",X"1B",X"35",
		X"03",X"00",X"1A",X"03",X"0A",X"0A",X"00",X"0C",X"10",X"0F",X"0D",X"11",X"12",X"12",X"0F",X"14",
		X"1F",X"1B",X"06",X"1C",X"0C",X"1C",X"00",X"25",X"13",X"26",X"04",X"28",X"1D",X"31",X"02",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"31",X"4C",X"38",X"C9",X"E5",X"D5",X"C5",X"F5",X"DD",X"E5",X"FD",X"E5",X"AF",X"32",X"81",X"A1",
		X"32",X"80",X"A0",X"3C",X"32",X"81",X"A1",X"CD",X"52",X"3A",X"CD",X"E1",X"3A",X"CD",X"4A",X"3B",
		X"CD",X"6B",X"3B",X"CD",X"F6",X"3B",X"CD",X"0C",X"3C",X"CD",X"38",X"3C",X"CF",X"CD",X"DD",X"3D",
		X"3A",X"00",X"A0",X"21",X"80",X"A0",X"B6",X"2F",X"0F",X"E6",X"01",X"21",X"05",X"80",X"AE",X"32",
		X"83",X"A1",X"FD",X"E1",X"DD",X"E1",X"F1",X"C1",X"D1",X"E1",X"FB",X"C9",X"11",X"39",X"67",X"39",
		X"B1",X"39",X"00",X"9C",X"0F",X"04",X"B1",X"39",X"00",X"9C",X"F0",X"04",X"B1",X"39",X"00",X"98",
		X"0F",X"04",X"B1",X"39",X"00",X"98",X"F0",X"04",X"B1",X"39",X"00",X"88",X"0F",X"04",X"B1",X"39",
		X"00",X"88",X"F0",X"04",X"B1",X"39",X"00",X"80",X"0F",X"04",X"B1",X"39",X"00",X"80",X"F0",X"04",
		X"B1",X"39",X"00",X"8C",X"0F",X"04",X"B1",X"39",X"00",X"8C",X"F0",X"04",X"46",X"3A",X"B1",X"39",
		X"00",X"84",X"0F",X"04",X"B1",X"39",X"00",X"84",X"F0",X"04",X"32",X"3A",X"9E",X"38",X"31",X"00",
		X"84",X"21",X"00",X"80",X"11",X"01",X"80",X"01",X"FF",X"03",X"36",X"00",X"ED",X"B0",X"21",X"00",
		X"88",X"11",X"01",X"88",X"01",X"FF",X"03",X"36",X"00",X"ED",X"B0",X"CD",X"1E",X"39",X"3E",X"01",
		X"32",X"84",X"A1",X"32",X"85",X"A1",X"21",X"A0",X"02",X"22",X"69",X"80",X"ED",X"5E",X"3E",X"3F",
		X"ED",X"47",X"3E",X"FE",X"D3",X"00",X"3E",X"01",X"32",X"81",X"A1",X"32",X"82",X"A1",X"FB",X"3A",
		X"00",X"A1",X"CB",X"47",X"28",X"F9",X"F3",X"AF",X"32",X"81",X"A1",X"32",X"82",X"A1",X"CD",X"1D",
		X"3E",X"01",X"00",X"00",X"3E",X"02",X"32",X"80",X"A0",X"3D",X"20",X"FA",X"0D",X"20",X"F5",X"10",
		X"F3",X"32",X"80",X"A0",X"3A",X"00",X"A1",X"CB",X"47",X"28",X"F6",X"CD",X"59",X"39",X"C3",X"03",
		X"00",X"21",X"00",X"84",X"11",X"01",X"84",X"01",X"FF",X"03",X"36",X"40",X"ED",X"B0",X"21",X"00",
		X"8C",X"11",X"01",X"8C",X"01",X"FF",X"03",X"36",X"66",X"ED",X"B0",X"21",X"40",X"80",X"01",X"08",
		X"1C",X"3E",X"40",X"57",X"3E",X"20",X"91",X"5F",X"7A",X"51",X"77",X"23",X"15",X"20",X"FB",X"19",
		X"10",X"F7",X"21",X"40",X"88",X"01",X"08",X"1C",X"3E",X"66",X"57",X"3E",X"20",X"91",X"5F",X"7A",
		X"51",X"77",X"23",X"15",X"20",X"FB",X"19",X"10",X"F7",X"21",X"00",X"A0",X"01",X"00",X"02",X"71",
		X"2C",X"20",X"FC",X"24",X"10",X"F9",X"C9",X"11",X"F9",X"3F",X"21",X"00",X"00",X"01",X"00",X"10",
		X"32",X"80",X"A0",X"79",X"86",X"4F",X"2C",X"20",X"FA",X"24",X"10",X"F4",X"1A",X"B9",X"20",X"0F",
		X"13",X"7B",X"FE",X"FD",X"38",X"E7",X"3E",X"4F",X"32",X"8B",X"84",X"3E",X"4B",X"18",X"03",X"7B",
		X"D6",X"F8",X"32",X"8C",X"84",X"06",X"4F",X"21",X"86",X"84",X"36",X"4D",X"2D",X"70",X"2D",X"36",
		X"52",X"FE",X"4B",X"C8",X"32",X"80",X"A0",X"3A",X"00",X"A1",X"CB",X"47",X"28",X"F6",X"C3",X"00",
		X"00",X"16",X"0F",X"E1",X"C1",X"5A",X"32",X"80",X"A0",X"7B",X"0F",X"0F",X"0F",X"0F",X"83",X"80",
		X"A1",X"77",X"7B",X"87",X"87",X"83",X"3C",X"5F",X"2C",X"20",X"EE",X"24",X"10",X"E8",X"3B",X"3B",
		X"3B",X"3B",X"E1",X"C1",X"5A",X"32",X"80",X"A0",X"7B",X"0F",X"0F",X"0F",X"0F",X"83",X"80",X"AE",
		X"A1",X"20",X"17",X"7B",X"87",X"87",X"83",X"3C",X"5F",X"2C",X"20",X"EC",X"24",X"10",X"E6",X"3B",
		X"3B",X"3B",X"3B",X"15",X"F2",X"B3",X"39",X"E1",X"C1",X"C9",X"7C",X"0F",X"E6",X"0E",X"FE",X"0C",
		X"38",X"02",X"D6",X"04",X"CB",X"41",X"20",X"01",X"3C",X"FE",X"04",X"30",X"0F",X"FE",X"02",X"38",
		X"0B",X"21",X"00",X"9C",X"11",X"00",X"84",X"01",X"00",X"04",X"ED",X"B0",X"CB",X"3F",X"32",X"CB",
		X"84",X"3E",X"4C",X"30",X"02",X"3E",X"48",X"32",X"CC",X"84",X"06",X"0A",X"21",X"C6",X"84",X"C3",
		X"9A",X"39",X"21",X"00",X"9C",X"11",X"00",X"84",X"01",X"00",X"04",X"ED",X"B0",X"3E",X"4F",X"32",
		X"CB",X"84",X"3E",X"4B",X"18",X"E1",X"21",X"00",X"84",X"11",X"00",X"9C",X"01",X"00",X"04",X"ED",
		X"B0",X"C9",X"3A",X"00",X"A1",X"07",X"07",X"07",X"E6",X"06",X"5F",X"16",X"00",X"21",X"AB",X"3A",
		X"19",X"5E",X"23",X"56",X"ED",X"53",X"00",X"80",X"3A",X"00",X"A1",X"0F",X"0F",X"E6",X"0E",X"5F",
		X"16",X"00",X"21",X"B3",X"3A",X"19",X"5E",X"23",X"56",X"ED",X"53",X"02",X"80",X"7B",X"3D",X"3D",
		X"87",X"5F",X"16",X"00",X"21",X"C3",X"3A",X"19",X"5E",X"23",X"56",X"3A",X"00",X"A1",X"0F",X"E6",
		X"03",X"6F",X"26",X"00",X"19",X"7E",X"32",X"04",X"80",X"11",X"0C",X"00",X"19",X"7E",X"32",X"07",
		X"80",X"3A",X"80",X"A0",X"2F",X"E6",X"01",X"32",X"05",X"80",X"C9",X"00",X"00",X"02",X"01",X"01",
		X"02",X"01",X"01",X"03",X"41",X"04",X"41",X"01",X"42",X"02",X"42",X"03",X"42",X"01",X"43",X"02",
		X"43",X"03",X"43",X"C9",X"3A",X"CD",X"3A",X"D1",X"3A",X"FF",X"10",X"20",X"30",X"FF",X"20",X"20",
		X"20",X"FF",X"20",X"40",X"60",X"FF",X"FF",X"FF",X"FF",X"FF",X"08",X"10",X"12",X"FF",X"FF",X"FF",
		X"FF",X"3A",X"00",X"80",X"A7",X"20",X"1D",X"21",X"F3",X"3A",X"11",X"04",X"85",X"01",X"11",X"00",
		X"ED",X"B0",X"C9",X"46",X"52",X"45",X"45",X"40",X"50",X"4C",X"41",X"59",X"40",X"40",X"40",X"40",
		X"40",X"40",X"40",X"40",X"21",X"3E",X"3B",X"11",X"05",X"85",X"01",X"05",X"00",X"ED",X"B0",X"21",
		X"43",X"3B",X"11",X"0D",X"85",X"01",X"07",X"00",X"ED",X"B0",X"3A",X"00",X"80",X"FE",X"01",X"32",
		X"04",X"85",X"21",X"40",X"40",X"28",X"02",X"2E",X"53",X"22",X"0A",X"85",X"3A",X"01",X"80",X"FE",
		X"01",X"32",X"0C",X"85",X"3E",X"40",X"28",X"02",X"3E",X"53",X"32",X"14",X"85",X"C9",X"40",X"43",
		X"4F",X"49",X"4E",X"40",X"43",X"52",X"45",X"44",X"49",X"54",X"21",X"67",X"3B",X"11",X"45",X"85",
		X"01",X"04",X"00",X"ED",X"B0",X"3A",X"02",X"80",X"FE",X"01",X"32",X"44",X"85",X"3E",X"40",X"28",
		X"02",X"3E",X"53",X"32",X"49",X"85",X"C9",X"40",X"43",X"41",X"52",X"21",X"EA",X"3B",X"11",X"84",
		X"85",X"01",X"05",X"00",X"ED",X"B0",X"3A",X"04",X"80",X"3C",X"20",X"11",X"21",X"EF",X"3B",X"11",
		X"8B",X"85",X"01",X"07",X"00",X"ED",X"B0",X"EB",X"36",X"40",X"C3",X"E1",X"3B",X"21",X"8B",X"85",
		X"36",X"40",X"2C",X"3A",X"04",X"80",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"20",X"02",X"3E",X"40",
		X"77",X"2C",X"3A",X"04",X"80",X"E6",X"0F",X"77",X"2C",X"36",X"00",X"2C",X"36",X"00",X"2C",X"36",
		X"00",X"2C",X"36",X"40",X"3A",X"07",X"80",X"3C",X"CA",X"E1",X"3B",X"0F",X"0F",X"0F",X"0F",X"E6",
		X"0F",X"20",X"02",X"3E",X"40",X"2C",X"36",X"2C",X"2C",X"36",X"40",X"2C",X"77",X"3A",X"07",X"80",
		X"E6",X"0F",X"2C",X"77",X"2C",X"36",X"00",X"2C",X"36",X"00",X"2C",X"36",X"00",X"2C",X"36",X"00",
		X"C9",X"3E",X"0A",X"2C",X"36",X"40",X"3D",X"20",X"FA",X"C9",X"42",X"4F",X"4E",X"55",X"53",X"4E",
		X"4F",X"54",X"48",X"49",X"4E",X"47",X"21",X"08",X"3C",X"11",X"C4",X"85",X"01",X"04",X"00",X"ED",
		X"B0",X"3A",X"03",X"80",X"32",X"CC",X"85",X"C9",X"52",X"41",X"4E",X"4B",X"3A",X"05",X"80",X"A7",
		X"20",X"0C",X"21",X"31",X"3C",X"11",X"04",X"86",X"01",X"07",X"00",X"ED",X"B0",X"C9",X"21",X"2A",
		X"3C",X"11",X"04",X"86",X"01",X"07",X"00",X"ED",X"B0",X"C9",X"54",X"41",X"42",X"4C",X"45",X"40",
		X"40",X"55",X"50",X"52",X"49",X"47",X"48",X"54",X"3A",X"00",X"A0",X"01",X"03",X"00",X"21",X"13",
		X"80",X"11",X"14",X"80",X"ED",X"B8",X"23",X"77",X"23",X"B6",X"2F",X"23",X"A6",X"23",X"A6",X"23",
		X"77",X"CD",X"A9",X"3C",X"CD",X"BA",X"3C",X"CD",X"CB",X"3C",X"CD",X"DC",X"3C",X"CD",X"ED",X"3C",
		X"CD",X"FE",X"3C",X"CD",X"0F",X"3D",X"CD",X"25",X"3D",X"3A",X"80",X"A0",X"01",X"03",X"00",X"21",
		X"1B",X"80",X"11",X"1C",X"80",X"ED",X"B8",X"23",X"77",X"23",X"B6",X"2F",X"23",X"A6",X"23",X"A6",
		X"23",X"77",X"2B",X"7E",X"2B",X"B6",X"2F",X"2B",X"A6",X"2B",X"A6",X"2B",X"77",X"CD",X"36",X"3D",
		X"CD",X"47",X"3D",X"CD",X"58",X"3D",X"CD",X"69",X"3D",X"CD",X"7C",X"3D",X"CD",X"8A",X"3D",X"CD",
		X"9B",X"3D",X"CD",X"AC",X"3D",X"CD",X"BD",X"3D",X"C9",X"3A",X"15",X"80",X"CB",X"7F",X"C8",X"21",
		X"F6",X"89",X"CB",X"FE",X"3E",X"37",X"CD",X"C9",X"3D",X"C9",X"3A",X"15",X"80",X"CB",X"77",X"C8",
		X"21",X"F5",X"89",X"CB",X"FE",X"3E",X"36",X"CD",X"C9",X"3D",X"C9",X"3A",X"15",X"80",X"CB",X"6F",
		X"C8",X"21",X"F4",X"89",X"CB",X"EE",X"3E",X"35",X"CD",X"C9",X"3D",X"C9",X"3A",X"15",X"80",X"CB",
		X"67",X"C8",X"21",X"F4",X"89",X"CB",X"CE",X"3E",X"34",X"CD",X"C9",X"3D",X"C9",X"3A",X"15",X"80",
		X"CB",X"5F",X"C8",X"21",X"F4",X"89",X"CB",X"DE",X"3E",X"33",X"CD",X"C9",X"3D",X"C9",X"3A",X"15",
		X"80",X"CB",X"57",X"C8",X"21",X"F4",X"89",X"CB",X"D6",X"3E",X"32",X"CD",X"C9",X"3D",X"C9",X"3A",
		X"15",X"80",X"CB",X"4F",X"C8",X"21",X"F4",X"89",X"CB",X"76",X"28",X"03",X"CB",X"E6",X"C9",X"21",
		X"F4",X"89",X"CB",X"C6",X"C9",X"3A",X"15",X"80",X"CB",X"47",X"C8",X"21",X"F6",X"89",X"CB",X"F6",
		X"3E",X"30",X"CD",X"C9",X"3D",X"C9",X"3A",X"1D",X"80",X"CB",X"7F",X"C8",X"21",X"F6",X"89",X"CB",
		X"FE",X"3E",X"46",X"CD",X"C9",X"3D",X"C9",X"3A",X"1D",X"80",X"CB",X"77",X"C8",X"21",X"F5",X"89",
		X"CB",X"F6",X"3E",X"45",X"CD",X"C9",X"3D",X"C9",X"3A",X"1D",X"80",X"CB",X"6F",X"C8",X"21",X"F5",
		X"89",X"CB",X"EE",X"3E",X"44",X"CD",X"C9",X"3D",X"C9",X"3A",X"1D",X"80",X"CB",X"67",X"C8",X"21",
		X"F5",X"89",X"CB",X"E6",X"CB",X"9E",X"3E",X"43",X"CD",X"C9",X"3D",X"C9",X"3A",X"18",X"80",X"CB",
		X"67",X"C8",X"21",X"F5",X"89",X"CB",X"DE",X"CB",X"A6",X"C9",X"3A",X"1D",X"80",X"CB",X"5F",X"C8",
		X"21",X"F4",X"89",X"CB",X"FE",X"3E",X"42",X"CD",X"C9",X"3D",X"C9",X"3A",X"1D",X"80",X"CB",X"57",
		X"C8",X"21",X"F5",X"89",X"CB",X"D6",X"3E",X"41",X"CD",X"C9",X"3D",X"C9",X"3A",X"1D",X"80",X"CB",
		X"4F",X"C8",X"21",X"F4",X"89",X"CB",X"F6",X"3E",X"39",X"CD",X"C9",X"3D",X"C9",X"3A",X"18",X"80",
		X"CB",X"4F",X"C8",X"21",X"F4",X"89",X"CB",X"B6",X"C9",X"21",X"00",X"A0",X"CB",X"4E",X"C0",X"21",
		X"21",X"80",X"11",X"20",X"80",X"01",X"0F",X"00",X"ED",X"B0",X"2B",X"77",X"C9",X"21",X"20",X"80",
		X"11",X"0D",X"3E",X"06",X"10",X"1A",X"FE",X"FF",X"28",X"02",X"BE",X"C0",X"23",X"13",X"10",X"F5",
		X"21",X"FC",X"3D",X"11",X"84",X"86",X"01",X"11",X"00",X"ED",X"B0",X"C9",X"18",X"40",X"4E",X"41",
		X"4D",X"43",X"4F",X"40",X"4C",X"54",X"44",X"2E",X"40",X"31",X"39",X"38",X"30",X"35",X"35",X"34",
		X"34",X"34",X"34",X"34",X"34",X"34",X"33",X"32",X"32",X"32",X"32",X"32",X"32",X"3E",X"03",X"32",
		X"30",X"A1",X"21",X"00",X"84",X"11",X"01",X"84",X"01",X"FF",X"03",X"36",X"5B",X"ED",X"B0",X"21",
		X"40",X"80",X"01",X"08",X"1C",X"3E",X"5B",X"CD",X"6F",X"3E",X"21",X"00",X"8C",X"01",X"00",X"04",
		X"CD",X"5F",X"3E",X"23",X"0B",X"79",X"B0",X"20",X"F7",X"21",X"40",X"88",X"01",X"08",X"1C",X"3E",
		X"20",X"91",X"5F",X"51",X"CD",X"5F",X"3E",X"23",X"15",X"20",X"F9",X"19",X"10",X"F5",X"C9",X"CB",
		X"45",X"CB",X"F6",X"28",X"02",X"CB",X"B6",X"CB",X"6D",X"CB",X"BE",X"C8",X"CB",X"FE",X"C9",X"57",
		X"3E",X"20",X"91",X"5F",X"7A",X"51",X"77",X"23",X"15",X"20",X"FB",X"19",X"10",X"F7",X"C9",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"75",X"C3",X"C8",X"AE",X"52",X"04",X"38");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
