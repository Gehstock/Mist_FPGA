library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity gfx_3j is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of gfx_3j is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"3C",X"62",X"C8",X"84",X"84",X"94",X"4C",X"20",X"FE",X"80",X"20",X"20",X"20",X"24",X"20",X"20",
		X"FF",X"80",X"38",X"60",X"C0",X"87",X"9C",X"40",X"7E",X"C1",X"84",X"9C",X"00",X"60",X"CE",X"80",
		X"70",X"40",X"CF",X"80",X"4C",X"48",X"40",X"40",X"7E",X"C1",X"80",X"80",X"9F",X"00",X"7C",X"40",
		X"7E",X"C1",X"84",X"9C",X"00",X"0C",X"78",X"40",X"1C",X"10",X"10",X"30",X"60",X"C7",X"9C",X"80",
		X"7E",X"C1",X"82",X"86",X"61",X"48",X"5C",X"20",X"3E",X"60",X"C0",X"9E",X"81",X"84",X"9C",X"40",
		X"00",X"00",X"00",X"00",X"6C",X"5A",X"48",X"48",X"00",X"00",X"00",X"7E",X"40",X"00",X"00",X"00",
		X"78",X"40",X"20",X"10",X"18",X"30",X"60",X"40",X"00",X"00",X"7E",X"40",X"00",X"7E",X"40",X"00",
		X"1E",X"30",X"60",X"C0",X"80",X"40",X"20",X"10",X"38",X"20",X"38",X"60",X"C7",X"84",X"9C",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E7",X"84",X"9C",X"80",X"84",X"8C",X"48",X"20",
		X"7F",X"C0",X"84",X"9C",X"40",X"84",X"9C",X"40",X"7C",X"C2",X"89",X"04",X"04",X"EC",X"98",X"00",
		X"3F",X"60",X"C4",X"84",X"84",X"94",X"4C",X"20",X"FF",X"80",X"04",X"7C",X"40",X"04",X"FC",X"80",
		X"07",X"04",X"04",X"7C",X"40",X"04",X"FC",X"80",X"FC",X"82",X"89",X"94",X"84",X"04",X"F8",X"80",
		X"E7",X"84",X"84",X"9C",X"80",X"84",X"84",X"84",X"FE",X"80",X"20",X"20",X"20",X"20",X"E6",X"80",
		X"7E",X"C1",X"84",X"84",X"80",X"80",X"80",X"80",X"F7",X"84",X"04",X"00",X"30",X"64",X"C4",X"84",
		X"FE",X"80",X"08",X"08",X"08",X"08",X"08",X"08",X"E7",X"84",X"9C",X"94",X"80",X"80",X"88",X"84",
		X"E7",X"84",X"84",X"84",X"80",X"90",X"88",X"84",X"3E",X"41",X"84",X"84",X"84",X"84",X"9C",X"40",
		X"07",X"04",X"7C",X"C0",X"84",X"84",X"9C",X"40",X"DE",X"A1",X"CC",X"84",X"84",X"84",X"9C",X"40",
		X"F7",X"84",X"04",X"E0",X"84",X"84",X"9C",X"40",X"7E",X"C1",X"84",X"9E",X"41",X"74",X"4C",X"20",
		X"38",X"20",X"20",X"20",X"20",X"20",X"E6",X"80",X"7E",X"C1",X"84",X"84",X"84",X"84",X"84",X"84",
		X"18",X"30",X"60",X"C0",X"88",X"84",X"84",X"84",X"E7",X"8C",X"88",X"80",X"80",X"94",X"84",X"84",
		X"E7",X"8C",X"88",X"00",X"60",X"C0",X"88",X"84",X"38",X"20",X"20",X"64",X"C2",X"88",X"88",X"88",
		X"FF",X"80",X"18",X"30",X"60",X"C0",X"8F",X"80",X"18",X"16",X"08",X"08",X"00",X"00",X"00",X"00",
		X"70",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"04",X"08",X"10",X"20",X"40",X"00",
		X"00",X"38",X"20",X"20",X"00",X"00",X"00",X"00",X"FE",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"38",X"24",X"10",X"10",X"10",X"10",X"10",X"20",X"1C",X"30",X"20",X"20",X"20",X"20",X"24",X"10",
		X"FE",X"A0",X"80",X"98",X"10",X"00",X"38",X"A0",X"3E",X"44",X"A4",X"A4",X"A4",X"A5",X"A5",X"44",
		X"BE",X"68",X"28",X"28",X"10",X"28",X"28",X"10",X"7B",X"46",X"A5",X"A5",X"45",X"A5",X"A5",X"45",
		X"77",X"44",X"44",X"33",X"C4",X"88",X"88",X"88",X"38",X"20",X"20",X"18",X"60",X"40",X"40",X"40",
		X"00",X"62",X"44",X"28",X"10",X"28",X"44",X"00",X"00",X"00",X"38",X"20",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"60",X"50",X"40",X"40",X"00",X"2B",X"2B",X"2B",X"2B",X"2B",X"3F",X"16",
		X"00",X"93",X"93",X"93",X"9F",X"93",X"9F",X"8E",X"00",X"C9",X"C9",X"C9",X"C7",X"C9",X"CF",X"C7",
		X"00",X"38",X"4C",X"4C",X"4C",X"4C",X"7C",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"50",X"50",X"50",X"50",X"50",X"00",X"A0",X"EF",X"49",X"59",X"41",X"49",X"49",X"59",X"20",
		X"FB",X"92",X"92",X"96",X"88",X"92",X"96",X"88",X"0E",X"11",X"24",X"24",X"24",X"24",X"2C",X"10",
		X"00",X"00",X"F0",X"F0",X"F8",X"A0",X"00",X"00",X"00",X"00",X"07",X"07",X"07",X"03",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"24",X"24",X"42",X"42",X"24",X"24",X"18",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FC",X"80",X"10",X"10",X"10",X"10",X"10",X"10",X"8E",X"11",X"20",X"20",X"20",X"20",X"20",X"20",
		X"F3",X"0A",X"22",X"62",X"22",X"22",X"E2",X"02",X"1D",X"11",X"11",X"11",X"11",X"10",X"11",X"11",
		X"00",X"00",X"F0",X"F0",X"F8",X"A0",X"00",X"00",X"00",X"00",X"07",X"07",X"07",X"03",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"D3",X"D3",X"D3",X"8F",X"00",X"01",X"01",X"FE",X"AA",X"AA",X"AA",X"A9",X"00",X"80",X"80",X"7F",
		X"FE",X"01",X"01",X"00",X"81",X"C1",X"CF",X"D3",X"18",X"24",X"24",X"42",X"42",X"24",X"24",X"18",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E7",X"84",X"9C",X"80",X"84",X"8C",X"48",X"20",X"7F",X"C0",X"84",X"9C",X"40",X"84",X"9C",X"40",
		X"7C",X"C2",X"89",X"04",X"04",X"EC",X"98",X"00",X"3F",X"60",X"C4",X"84",X"84",X"94",X"4C",X"20",
		X"FF",X"80",X"04",X"7C",X"40",X"04",X"FC",X"80",X"07",X"04",X"04",X"7C",X"40",X"04",X"FC",X"80",
		X"FC",X"82",X"89",X"94",X"84",X"04",X"F8",X"80",X"E7",X"84",X"84",X"9C",X"80",X"84",X"84",X"84",
		X"FE",X"80",X"20",X"20",X"20",X"20",X"E6",X"80",X"7E",X"C1",X"84",X"84",X"80",X"80",X"80",X"80",
		X"F7",X"84",X"04",X"00",X"30",X"64",X"C4",X"84",X"FE",X"80",X"08",X"08",X"08",X"08",X"08",X"08",
		X"E7",X"84",X"9C",X"94",X"80",X"80",X"88",X"84",X"E7",X"84",X"84",X"84",X"80",X"90",X"88",X"84",
		X"3E",X"41",X"84",X"84",X"84",X"84",X"9C",X"40",X"07",X"04",X"7C",X"C0",X"84",X"84",X"9C",X"40",
		X"DE",X"A1",X"CC",X"84",X"84",X"84",X"9C",X"40",X"F7",X"84",X"04",X"E0",X"84",X"84",X"9C",X"40",
		X"7E",X"C1",X"84",X"9E",X"41",X"74",X"4C",X"20",X"38",X"20",X"20",X"20",X"20",X"20",X"E6",X"80",
		X"7E",X"C1",X"84",X"84",X"84",X"84",X"84",X"84",X"18",X"30",X"60",X"C0",X"88",X"84",X"84",X"84",
		X"E7",X"8C",X"88",X"80",X"80",X"94",X"84",X"84",X"E7",X"8C",X"88",X"00",X"60",X"C0",X"88",X"84",
		X"38",X"20",X"20",X"64",X"C2",X"88",X"88",X"88",X"FF",X"80",X"18",X"30",X"60",X"C0",X"8F",X"80",
		X"77",X"44",X"44",X"33",X"C4",X"88",X"88",X"88",X"00",X"0E",X"08",X"08",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"C0",X"C0",X"C0",X"C0",X"F0",X"00",X"00",X"E1",X"31",X"31",X"31",X"31",X"E7",X"00",
		X"00",X"E3",X"E6",X"E6",X"E6",X"E6",X"E3",X"00",X"00",X"00",X"00",X"0F",X"1C",X"1C",X"0F",X"00",
		X"00",X"E0",X"F0",X"00",X"06",X"F6",X"F0",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"07",X"0F",X"00",X"60",X"6F",X"0F",X"00",X"00",X"81",X"C3",X"C3",X"C3",X"FF",X"FF",X"00",
		X"00",X"81",X"C3",X"C3",X"C3",X"FF",X"FF",X"00",X"00",X"81",X"C3",X"C3",X"C3",X"FF",X"FF",X"00",
		X"00",X"EF",X"E7",X"E1",X"00",X"FE",X"7E",X"1E",X"2E",X"6E",X"6E",X"EE",X"1E",X"02",X"00",X"FF",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"1A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"C0",X"F8",X"F0",X"C0",X"F0",X"78",X"7C",X"7B",X"37",X"7F",X"65",X"46",X"46",X"04",X"00",X"00",
		X"00",X"EF",X"E7",X"E1",X"00",X"FE",X"7E",X"1E",X"2E",X"6E",X"6E",X"EE",X"1E",X"02",X"00",X"FF",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"1A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FE",X"BA",X"BB",X"77",X"FF",X"FF",X"FE",X"FF",X"FF",X"BB",X"BB",X"B7",X"7F",X"DD",X"EF",
		X"7F",X"7F",X"7B",X"77",X"FF",X"FF",X"FF",X"7F",X"80",X"C0",X"E0",X"F0",X"E8",X"DC",X"BE",X"80",
		X"80",X"C0",X"E0",X"F0",X"E8",X"DC",X"BE",X"80",X"80",X"C0",X"E0",X"F0",X"E8",X"DC",X"BE",X"80",
		X"00",X"E0",X"F0",X"00",X"06",X"F6",X"F0",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"07",X"0F",X"00",X"60",X"6F",X"0F",X"00",X"FF",X"01",X"01",X"01",X"01",X"03",X"06",X"FC",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"80",X"80",X"80",X"80",X"C0",X"60",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"83",X"C0",X"0C",X"5E",X"82",X"00",X"78",X"00",
		X"38",X"20",X"20",X"64",X"C2",X"88",X"88",X"88",X"3E",X"41",X"84",X"84",X"84",X"84",X"9C",X"40",
		X"7E",X"C1",X"84",X"84",X"84",X"84",X"84",X"84",X"3F",X"60",X"C4",X"84",X"84",X"94",X"4C",X"20",
		X"FE",X"80",X"20",X"20",X"20",X"20",X"E6",X"80",X"38",X"20",X"20",X"20",X"20",X"20",X"E6",X"80",
		X"F7",X"84",X"04",X"00",X"30",X"64",X"C4",X"84",X"FF",X"80",X"04",X"7C",X"40",X"04",X"FC",X"80",
		X"07",X"04",X"7C",X"C0",X"84",X"84",X"9C",X"40",X"FC",X"82",X"89",X"94",X"84",X"04",X"F8",X"80",
		X"E7",X"84",X"84",X"84",X"80",X"90",X"88",X"84",X"7E",X"C1",X"84",X"9E",X"41",X"74",X"4C",X"20",
		X"E7",X"84",X"84",X"9C",X"80",X"84",X"84",X"84",X"00",X"0E",X"08",X"08",X"00",X"00",X"00",X"00",
		X"77",X"44",X"44",X"33",X"C4",X"88",X"88",X"88",X"38",X"20",X"20",X"18",X"60",X"40",X"40",X"40",
		X"00",X"E0",X"F0",X"00",X"06",X"F6",X"F0",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"07",X"0F",X"00",X"60",X"6F",X"0F",X"00",X"77",X"77",X"00",X"88",X"88",X"00",X"77",X"77",
		X"77",X"77",X"00",X"88",X"88",X"00",X"77",X"77",X"77",X"77",X"00",X"08",X"08",X"00",X"77",X"77",
		X"07",X"04",X"7C",X"C0",X"84",X"84",X"9C",X"40",X"FF",X"80",X"04",X"7C",X"40",X"04",X"FC",X"80",
		X"F7",X"84",X"04",X"E0",X"84",X"84",X"9C",X"40",X"07",X"04",X"04",X"7C",X"40",X"04",X"FC",X"80",
		X"7C",X"C0",X"88",X"04",X"04",X"EC",X"98",X"00",X"38",X"20",X"20",X"20",X"20",X"20",X"E6",X"80",
		X"07",X"04",X"7C",X"C0",X"84",X"84",X"9C",X"40",X"38",X"20",X"20",X"20",X"20",X"20",X"E6",X"80",
		X"7E",X"C0",X"84",X"9E",X"40",X"74",X"4C",X"20",X"00",X"00",X"00",X"00",X"60",X"50",X"40",X"40",
		X"3C",X"62",X"C8",X"84",X"84",X"94",X"4C",X"20",X"FE",X"80",X"20",X"20",X"20",X"24",X"20",X"20",
		X"FF",X"80",X"38",X"60",X"C0",X"87",X"9C",X"40",X"7E",X"C0",X"84",X"9C",X"00",X"60",X"CE",X"80",
		X"70",X"40",X"CF",X"80",X"4C",X"48",X"40",X"40",X"7E",X"C0",X"80",X"80",X"9F",X"00",X"7C",X"40",
		X"7E",X"C0",X"84",X"9C",X"00",X"0C",X"78",X"40",X"1C",X"10",X"10",X"30",X"60",X"C7",X"9C",X"80",
		X"7E",X"C0",X"82",X"86",X"60",X"48",X"5C",X"20",X"3E",X"60",X"C0",X"9E",X"80",X"84",X"9C",X"40",
		X"07",X"04",X"04",X"7C",X"40",X"04",X"FC",X"80",X"E7",X"84",X"9C",X"80",X"84",X"8C",X"48",X"20",
		X"7C",X"C0",X"88",X"04",X"04",X"EC",X"98",X"00",X"FF",X"80",X"04",X"7C",X"40",X"04",X"FC",X"80",
		X"77",X"44",X"44",X"33",X"C4",X"88",X"88",X"88",X"38",X"20",X"20",X"18",X"60",X"40",X"40",X"40",
		X"3C",X"62",X"C8",X"84",X"84",X"94",X"4C",X"20",X"FE",X"80",X"20",X"20",X"20",X"24",X"20",X"20",
		X"FF",X"80",X"38",X"60",X"C0",X"87",X"9C",X"40",X"7E",X"C1",X"84",X"9C",X"00",X"60",X"CE",X"80",
		X"70",X"40",X"CF",X"80",X"4C",X"48",X"40",X"40",X"7E",X"C1",X"80",X"80",X"9F",X"00",X"7C",X"40",
		X"7E",X"C1",X"84",X"9C",X"00",X"0C",X"78",X"40",X"1C",X"10",X"10",X"30",X"60",X"C7",X"9C",X"80",
		X"7E",X"C1",X"82",X"86",X"61",X"48",X"5C",X"20",X"3E",X"60",X"C0",X"9E",X"81",X"84",X"9C",X"40",
		X"00",X"00",X"00",X"00",X"6C",X"5A",X"48",X"48",X"00",X"00",X"00",X"7E",X"40",X"00",X"00",X"00",
		X"78",X"40",X"20",X"10",X"18",X"30",X"60",X"40",X"00",X"00",X"7E",X"40",X"00",X"7E",X"40",X"00",
		X"1E",X"30",X"60",X"C0",X"80",X"40",X"20",X"10",X"38",X"20",X"38",X"60",X"C7",X"84",X"9C",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E7",X"84",X"9C",X"80",X"84",X"8C",X"48",X"20",
		X"7F",X"C0",X"84",X"9C",X"40",X"84",X"9C",X"40",X"7C",X"C2",X"89",X"04",X"04",X"EC",X"98",X"00",
		X"3F",X"60",X"C4",X"84",X"84",X"94",X"4C",X"20",X"FF",X"80",X"04",X"7C",X"40",X"04",X"FC",X"80",
		X"07",X"04",X"04",X"7C",X"40",X"04",X"FC",X"80",X"FC",X"82",X"89",X"94",X"84",X"04",X"F8",X"80",
		X"E7",X"84",X"84",X"9C",X"80",X"84",X"84",X"84",X"FE",X"80",X"20",X"20",X"20",X"20",X"E6",X"80",
		X"7E",X"C1",X"84",X"84",X"80",X"80",X"80",X"80",X"F7",X"84",X"04",X"00",X"30",X"64",X"C4",X"84",
		X"FE",X"80",X"08",X"08",X"08",X"08",X"08",X"08",X"E7",X"84",X"9C",X"94",X"80",X"80",X"88",X"84",
		X"E7",X"84",X"84",X"84",X"80",X"90",X"88",X"84",X"3E",X"41",X"84",X"84",X"84",X"84",X"9C",X"40",
		X"07",X"04",X"7C",X"C0",X"84",X"84",X"9C",X"40",X"DE",X"A1",X"CC",X"84",X"84",X"84",X"9C",X"40",
		X"F7",X"84",X"04",X"E0",X"84",X"84",X"9C",X"40",X"7E",X"C1",X"84",X"9E",X"41",X"74",X"4C",X"20",
		X"38",X"20",X"20",X"20",X"20",X"20",X"E6",X"80",X"7E",X"C1",X"84",X"84",X"84",X"84",X"84",X"84",
		X"18",X"30",X"60",X"C0",X"88",X"84",X"84",X"84",X"E7",X"8C",X"88",X"80",X"80",X"94",X"84",X"84",
		X"E7",X"8C",X"88",X"00",X"60",X"C0",X"88",X"84",X"38",X"20",X"20",X"64",X"C2",X"88",X"88",X"88",
		X"FF",X"80",X"18",X"30",X"60",X"C0",X"8F",X"80",X"18",X"16",X"08",X"08",X"00",X"00",X"00",X"00",
		X"70",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"04",X"08",X"10",X"20",X"40",X"00",
		X"00",X"38",X"20",X"20",X"00",X"00",X"00",X"00",X"FE",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"38",X"24",X"10",X"10",X"10",X"10",X"10",X"20",X"1C",X"30",X"20",X"20",X"20",X"20",X"24",X"10",
		X"FE",X"A0",X"80",X"98",X"10",X"00",X"38",X"A0",X"3E",X"44",X"A4",X"A4",X"A4",X"A5",X"A5",X"44",
		X"BE",X"68",X"28",X"28",X"10",X"28",X"28",X"10",X"7B",X"46",X"A5",X"A5",X"45",X"A5",X"A5",X"45",
		X"77",X"44",X"44",X"33",X"C4",X"88",X"88",X"88",X"38",X"20",X"20",X"18",X"60",X"40",X"40",X"40",
		X"00",X"62",X"44",X"28",X"10",X"28",X"44",X"00",X"00",X"00",X"38",X"20",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3C",X"62",X"C8",X"84",X"84",X"94",X"4C",X"20",X"FE",X"80",X"20",X"20",X"20",X"24",X"20",X"20",
		X"FF",X"80",X"38",X"60",X"C0",X"87",X"9C",X"40",X"7E",X"C1",X"84",X"9C",X"00",X"60",X"CE",X"80",
		X"70",X"40",X"CF",X"80",X"4C",X"48",X"40",X"40",X"7E",X"C1",X"80",X"80",X"9F",X"00",X"7C",X"40",
		X"7E",X"C1",X"84",X"9C",X"00",X"0C",X"78",X"40",X"1C",X"10",X"10",X"30",X"60",X"C7",X"9C",X"80",
		X"7E",X"C1",X"82",X"86",X"61",X"48",X"5C",X"20",X"3E",X"60",X"C0",X"9E",X"81",X"84",X"9C",X"40",
		X"00",X"00",X"00",X"00",X"6C",X"5A",X"48",X"48",X"00",X"00",X"00",X"7E",X"40",X"00",X"00",X"00",
		X"78",X"40",X"20",X"10",X"18",X"30",X"60",X"40",X"1E",X"30",X"60",X"C0",X"80",X"40",X"20",X"10",
		X"1E",X"30",X"60",X"C0",X"80",X"40",X"20",X"10",X"38",X"20",X"38",X"60",X"C7",X"84",X"9C",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E7",X"84",X"9C",X"80",X"84",X"8C",X"48",X"20",
		X"7F",X"C0",X"84",X"9C",X"40",X"84",X"9C",X"40",X"7C",X"C2",X"89",X"04",X"04",X"EC",X"98",X"00",
		X"3F",X"60",X"C4",X"84",X"84",X"94",X"4C",X"20",X"FF",X"80",X"04",X"7C",X"40",X"04",X"FC",X"80",
		X"07",X"04",X"04",X"7C",X"40",X"04",X"FC",X"80",X"FC",X"82",X"89",X"94",X"84",X"04",X"F8",X"80",
		X"E7",X"84",X"84",X"9C",X"80",X"84",X"84",X"84",X"FE",X"80",X"20",X"20",X"20",X"20",X"E6",X"80",
		X"7E",X"C1",X"84",X"84",X"80",X"80",X"80",X"80",X"F7",X"84",X"04",X"00",X"30",X"64",X"C4",X"84",
		X"FE",X"80",X"08",X"08",X"08",X"08",X"08",X"08",X"E7",X"84",X"9C",X"94",X"80",X"80",X"88",X"84",
		X"E7",X"84",X"84",X"84",X"80",X"90",X"88",X"84",X"3E",X"41",X"84",X"84",X"84",X"84",X"9C",X"40",
		X"07",X"04",X"7C",X"C0",X"84",X"84",X"9C",X"40",X"DE",X"A1",X"CC",X"84",X"84",X"84",X"9C",X"40",
		X"F7",X"84",X"04",X"E0",X"84",X"84",X"9C",X"40",X"7E",X"C1",X"84",X"9E",X"41",X"74",X"4C",X"20",
		X"38",X"20",X"20",X"20",X"20",X"20",X"E6",X"80",X"7E",X"C1",X"84",X"84",X"84",X"84",X"84",X"84",
		X"18",X"30",X"60",X"C0",X"88",X"84",X"84",X"84",X"E7",X"8C",X"88",X"80",X"80",X"94",X"84",X"84",
		X"E7",X"8C",X"88",X"00",X"60",X"C0",X"88",X"84",X"38",X"20",X"20",X"64",X"C2",X"88",X"88",X"88",
		X"FF",X"80",X"18",X"30",X"60",X"C0",X"8F",X"80",X"18",X"16",X"08",X"08",X"00",X"00",X"00",X"00",
		X"70",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"04",X"08",X"10",X"20",X"40",X"00",
		X"FE",X"48",X"48",X"48",X"49",X"48",X"78",X"48",X"FE",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"38",X"24",X"10",X"10",X"10",X"10",X"10",X"20",X"1C",X"30",X"20",X"20",X"20",X"20",X"24",X"10",
		X"FE",X"A0",X"80",X"98",X"10",X"00",X"38",X"A0",X"3E",X"44",X"A4",X"A4",X"A4",X"A5",X"A5",X"44",
		X"BE",X"68",X"28",X"28",X"10",X"28",X"28",X"10",X"7B",X"46",X"A5",X"A5",X"45",X"A5",X"A5",X"45",
		X"77",X"44",X"44",X"33",X"C4",X"88",X"88",X"88",X"38",X"20",X"20",X"18",X"60",X"40",X"40",X"40",
		X"00",X"62",X"44",X"28",X"10",X"28",X"44",X"00",X"00",X"00",X"38",X"20",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3C",X"62",X"C8",X"84",X"84",X"94",X"4C",X"20",X"FE",X"80",X"20",X"20",X"20",X"24",X"20",X"20",
		X"FF",X"80",X"38",X"60",X"C0",X"87",X"9C",X"40",X"7E",X"C1",X"84",X"9C",X"00",X"60",X"CE",X"80",
		X"70",X"40",X"CF",X"80",X"4C",X"48",X"40",X"40",X"7E",X"C1",X"80",X"80",X"9F",X"00",X"7C",X"40",
		X"7E",X"C1",X"84",X"9C",X"00",X"0C",X"78",X"40",X"1C",X"10",X"10",X"30",X"60",X"C7",X"9C",X"80",
		X"7E",X"C1",X"82",X"86",X"61",X"48",X"5C",X"20",X"3E",X"60",X"C0",X"9E",X"81",X"84",X"9C",X"40",
		X"00",X"00",X"00",X"00",X"6C",X"5A",X"48",X"48",X"00",X"00",X"00",X"7E",X"40",X"00",X"00",X"00",
		X"3E",X"41",X"BE",X"A2",X"BA",X"A2",X"BE",X"40",X"FE",X"08",X"08",X"F8",X"18",X"49",X"C8",X"08",
		X"F1",X"0A",X"24",X"64",X"0C",X"24",X"64",X"02",X"78",X"85",X"12",X"32",X"81",X"1E",X"33",X"81",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E7",X"84",X"9C",X"80",X"84",X"8C",X"48",X"20",
		X"7F",X"C0",X"84",X"9C",X"40",X"84",X"9C",X"40",X"7C",X"C2",X"89",X"04",X"04",X"EC",X"98",X"00",
		X"3F",X"60",X"C4",X"84",X"84",X"94",X"4C",X"20",X"FF",X"80",X"04",X"7C",X"40",X"04",X"FC",X"80",
		X"07",X"04",X"04",X"7C",X"40",X"04",X"FC",X"80",X"FC",X"82",X"89",X"94",X"84",X"04",X"F8",X"80",
		X"E7",X"84",X"84",X"9C",X"80",X"84",X"84",X"84",X"FE",X"80",X"20",X"20",X"20",X"20",X"E6",X"80",
		X"7E",X"C1",X"84",X"84",X"80",X"80",X"80",X"80",X"F7",X"84",X"04",X"00",X"30",X"64",X"C4",X"84",
		X"FE",X"80",X"08",X"08",X"08",X"08",X"08",X"08",X"E7",X"84",X"9C",X"94",X"80",X"80",X"88",X"84",
		X"E7",X"84",X"84",X"84",X"80",X"90",X"88",X"84",X"3E",X"41",X"84",X"84",X"84",X"84",X"9C",X"40",
		X"07",X"04",X"7C",X"C0",X"84",X"84",X"9C",X"40",X"DE",X"A1",X"CC",X"84",X"84",X"84",X"9C",X"40",
		X"F7",X"84",X"04",X"E0",X"84",X"84",X"9C",X"40",X"7E",X"C1",X"84",X"9E",X"41",X"74",X"4C",X"20",
		X"38",X"20",X"20",X"20",X"20",X"20",X"E6",X"80",X"7E",X"C1",X"84",X"84",X"84",X"84",X"84",X"84",
		X"18",X"30",X"60",X"C0",X"88",X"84",X"84",X"84",X"E7",X"8C",X"88",X"80",X"80",X"94",X"84",X"84",
		X"E7",X"8C",X"88",X"00",X"60",X"C0",X"88",X"84",X"38",X"20",X"20",X"64",X"C2",X"88",X"88",X"88",
		X"FF",X"80",X"18",X"30",X"60",X"C0",X"8F",X"80",X"18",X"16",X"08",X"08",X"00",X"00",X"00",X"00",
		X"70",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"70",X"40",X"41",X"41",X"40",X"01",X"81",X"40",
		X"FE",X"48",X"48",X"48",X"49",X"48",X"78",X"48",X"BB",X"22",X"22",X"22",X"66",X"10",X"00",X"00",
		X"F3",X"0A",X"E2",X"02",X"66",X"04",X"00",X"00",X"DF",X"12",X"13",X"12",X"32",X"80",X"00",X"00",
		X"FD",X"83",X"89",X"89",X"99",X"80",X"80",X"80",X"1E",X"21",X"44",X"44",X"4C",X"20",X"00",X"00",
		X"3C",X"42",X"88",X"88",X"98",X"40",X"00",X"00",X"8E",X"08",X"08",X"08",X"19",X"10",X"08",X"10",
		X"FB",X"26",X"20",X"20",X"22",X"26",X"10",X"08",X"BF",X"65",X"25",X"25",X"25",X"12",X"00",X"00",
		X"FF",X"90",X"9F",X"10",X"13",X"88",X"00",X"00",X"00",X"00",X"38",X"20",X"20",X"00",X"00",X"00",
		X"B8",X"60",X"20",X"27",X"24",X"24",X"38",X"20",X"EF",X"38",X"41",X"41",X"CF",X"08",X"00",X"00",
		X"CF",X"09",X"08",X"04",X"04",X"04",X"00",X"00",X"EF",X"89",X"89",X"89",X"99",X"41",X"01",X"01",
		X"FE",X"A1",X"04",X"04",X"3C",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3C",X"62",X"C8",X"84",X"84",X"94",X"4C",X"20",X"FE",X"80",X"20",X"20",X"20",X"24",X"20",X"20",
		X"FF",X"80",X"38",X"60",X"C0",X"87",X"9C",X"40",X"7E",X"C1",X"84",X"9C",X"00",X"60",X"CE",X"80",
		X"70",X"40",X"CF",X"80",X"4C",X"48",X"40",X"40",X"7E",X"C1",X"80",X"80",X"9F",X"00",X"7C",X"40",
		X"7E",X"C1",X"84",X"9C",X"00",X"0C",X"78",X"40",X"1C",X"10",X"10",X"30",X"60",X"C7",X"9C",X"80",
		X"7E",X"C1",X"82",X"86",X"61",X"48",X"5C",X"20",X"3E",X"60",X"C0",X"9E",X"81",X"84",X"9C",X"40",
		X"77",X"44",X"44",X"33",X"C4",X"88",X"88",X"88",X"00",X"00",X"00",X"7E",X"40",X"00",X"00",X"00",
		X"78",X"40",X"20",X"10",X"18",X"30",X"60",X"40",X"00",X"00",X"7E",X"40",X"00",X"7E",X"40",X"00",
		X"1E",X"30",X"60",X"C0",X"80",X"40",X"20",X"10",X"38",X"20",X"38",X"60",X"C7",X"84",X"9C",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E7",X"84",X"9C",X"80",X"84",X"8C",X"48",X"20",
		X"7F",X"C0",X"84",X"9C",X"40",X"84",X"9C",X"40",X"7C",X"C2",X"89",X"04",X"04",X"EC",X"98",X"00",
		X"3F",X"60",X"C4",X"84",X"84",X"94",X"4C",X"20",X"FF",X"80",X"04",X"7C",X"40",X"04",X"FC",X"80",
		X"07",X"04",X"04",X"7C",X"40",X"04",X"FC",X"80",X"FC",X"82",X"89",X"94",X"84",X"04",X"F8",X"80",
		X"E7",X"84",X"84",X"9C",X"80",X"84",X"84",X"84",X"FE",X"80",X"20",X"20",X"20",X"20",X"E6",X"80",
		X"7E",X"C1",X"84",X"84",X"80",X"80",X"80",X"80",X"F7",X"84",X"04",X"00",X"30",X"64",X"C4",X"84",
		X"FE",X"80",X"08",X"08",X"08",X"08",X"08",X"08",X"E7",X"84",X"9C",X"94",X"80",X"80",X"88",X"84",
		X"E7",X"84",X"84",X"84",X"80",X"90",X"88",X"84",X"3E",X"41",X"84",X"84",X"84",X"84",X"9C",X"40",
		X"07",X"04",X"7C",X"C0",X"84",X"84",X"9C",X"40",X"DE",X"A1",X"CC",X"84",X"84",X"84",X"9C",X"40",
		X"F7",X"84",X"04",X"E0",X"84",X"84",X"9C",X"40",X"7E",X"C1",X"84",X"9E",X"41",X"74",X"4C",X"20",
		X"38",X"20",X"20",X"20",X"20",X"20",X"E6",X"80",X"7E",X"C1",X"84",X"84",X"84",X"84",X"84",X"84",
		X"18",X"30",X"60",X"C0",X"88",X"84",X"84",X"84",X"E7",X"8C",X"88",X"80",X"80",X"94",X"84",X"84",
		X"E7",X"8C",X"88",X"00",X"60",X"C0",X"88",X"84",X"38",X"20",X"20",X"64",X"C2",X"88",X"88",X"88",
		X"FF",X"80",X"18",X"30",X"60",X"C0",X"8F",X"80",X"18",X"16",X"08",X"08",X"00",X"00",X"00",X"00",
		X"70",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"04",X"08",X"10",X"20",X"40",X"00",
		X"00",X"38",X"20",X"20",X"00",X"00",X"00",X"00",X"FE",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"38",X"24",X"10",X"10",X"10",X"10",X"10",X"20",X"1C",X"30",X"20",X"20",X"20",X"20",X"24",X"10",
		X"FE",X"A0",X"80",X"98",X"10",X"00",X"38",X"A0",X"3E",X"44",X"A4",X"A4",X"A4",X"A5",X"A5",X"44",
		X"BE",X"68",X"28",X"28",X"10",X"28",X"28",X"10",X"7B",X"46",X"A5",X"A5",X"45",X"A5",X"A5",X"45",
		X"77",X"44",X"44",X"33",X"C4",X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"20",X"20",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
