library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity bwidow_pgm_rom6 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of bwidow_pgm_rom6 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"F8",X"E5",X"CF",X"E5",X"00",X"E6",X"0E",X"E6",X"13",X"E6",X"1A",X"E6",X"1F",X"E6",X"2C",X"E6",
		X"49",X"E6",X"52",X"E6",X"62",X"E6",X"71",X"E6",X"8B",X"E6",X"A3",X"E6",X"B0",X"E6",X"BC",X"E6",
		X"C9",X"E6",X"E3",X"E6",X"02",X"E7",X"26",X"E7",X"61",X"0A",X"71",X"60",X"71",X"20",X"F1",X"56",
		X"71",X"38",X"41",X"A4",X"31",X"9C",X"61",X"94",X"21",X"60",X"21",X"08",X"E1",X"F8",X"21",X"F8",
		X"C1",X"98",X"21",X"92",X"71",X"E8",X"21",X"D8",X"C1",X"56",X"21",X"A1",X"21",X"A1",X"21",X"A1",
		X"21",X"A1",X"11",X"92",X"21",X"A0",X"21",X"89",X"21",X"B0",X"11",X"5A",X"C2",X"60",X"21",X"30",
		X"21",X"00",X"21",X"20",X"21",X"C0",X"21",X"C0",X"21",X"C0",X"21",X"C0",X"21",X"10",X"71",X"50",
		X"71",X"40",X"71",X"40",X"71",X"40",X"71",X"40",X"41",X"50",X"21",X"D0",X"21",X"F0",X"21",X"E0",
		X"71",X"40",X"71",X"30",X"71",X"20",X"71",X"40",X"E5",X"22",X"16",X"2E",X"1E",X"00",X"32",X"40",
		X"1E",X"B8",X"D9",X"20",X"26",X"30",X"00",X"1C",X"1E",X"00",X"34",X"16",X"38",X"3C",X"26",X"9E",
		X"E5",X"3A",X"34",X"26",X"1E",X"2C",X"1E",X"30",X"1C",X"9E",X"D3",X"28",X"3E",X"1E",X"22",X"32",
		X"00",X"3C",X"1E",X"38",X"2E",X"26",X"30",X"16",X"1C",X"B2",X"EB",X"34",X"2C",X"16",X"46",X"1E",
		X"38",X"80",X"EB",X"28",X"32",X"3E",X"1E",X"3E",X"38",X"80",X"E8",X"3A",X"34",X"26",X"1E",X"2C",
		X"1E",X"38",X"80",X"E8",X"28",X"3E",X"22",X"16",X"1C",X"32",X"38",X"80",X"DF",X"34",X"38",X"1E",
		X"3A",X"3A",X"00",X"3A",X"3C",X"16",X"38",X"BC",X"EE",X"20",X"38",X"1E",X"30",X"1A",X"A4",X"EE",
		X"22",X"1E",X"38",X"2E",X"16",X"B0",X"EB",X"3A",X"34",X"16",X"30",X"26",X"3A",X"A4",X"F4",X"34",
		X"2C",X"16",X"C6",X"F1",X"28",X"32",X"3E",X"1E",X"C8",X"F1",X"3A",X"34",X"26",X"1E",X"AC",X"EE",
		X"28",X"3E",X"1E",X"22",X"3E",X"9E",X"C7",X"1E",X"30",X"3C",X"1E",X"38",X"00",X"46",X"32",X"3E",
		X"38",X"00",X"26",X"30",X"26",X"3C",X"26",X"16",X"2C",X"BA",X"B8",X"3A",X"40",X"34",X"00",X"1E",
		X"30",X"3C",X"38",X"1E",X"48",X"00",X"40",X"32",X"3A",X"00",X"26",X"30",X"26",X"3C",X"26",X"16",
		X"2C",X"1E",X"BA",X"AC",X"22",X"1E",X"18",X"1E",X"30",X"00",X"3A",X"26",X"1E",X"00",X"26",X"24",
		X"38",X"1E",X"00",X"26",X"30",X"26",X"3C",X"26",X"16",X"2C",X"1E",X"30",X"00",X"1E",X"26",X"B0",
		X"C7",X"1E",X"30",X"3C",X"38",X"1E",X"00",X"3A",X"3E",X"3A",X"00",X"26",X"30",X"26",X"1A",X"26",
		X"16",X"2C",X"1E",X"BA",X"BE",X"1A",X"24",X"16",X"30",X"22",X"1E",X"00",X"42",X"26",X"3C",X"24",
		X"00",X"2C",X"1E",X"20",X"3C",X"00",X"3A",X"3C",X"26",X"1A",X"AA",X"A6",X"3C",X"32",X"3E",X"38",
		X"30",X"1E",X"48",X"00",X"2C",X"1E",X"00",X"18",X"32",X"3E",X"3C",X"32",X"30",X"00",X"34",X"32",
		X"3E",X"38",X"00",X"1A",X"24",X"16",X"30",X"22",X"1E",X"B8",X"B5",X"2A",X"30",X"32",X"34",X"20",
		X"00",X"1C",X"38",X"1E",X"24",X"1E",X"30",X"00",X"48",X"3E",X"2E",X"00",X"42",X"1E",X"1A",X"24",
		X"3A",X"1E",X"2C",X"B0",X"AC",X"22",X"26",X"38",X"1E",X"00",X"2C",X"16",X"00",X"34",X"1E",X"38",
		X"26",X"2C",X"2C",X"16",X"00",X"34",X"16",X"38",X"16",X"00",X"1A",X"16",X"2E",X"18",X"26",X"16",
		X"B8",X"B5",X"2E",X"32",X"40",X"1E",X"00",X"38",X"26",X"22",X"24",X"3C",X"00",X"3A",X"3C",X"26",
		X"1A",X"2A",X"00",X"3C",X"32",X"00",X"1E",X"30",X"3C",X"1E",X"B8",X"B2",X"34",X"32",X"3E",X"3A",
		X"3A",X"1E",X"48",X"00",X"20",X"1E",X"3E",X"00",X"36",X"3E",X"16",X"30",X"1C",X"00",X"1A",X"32",
		X"38",X"38",X"1E",X"1A",X"3C",X"9E",X"B2",X"20",X"26",X"38",X"1E",X"00",X"1C",X"38",X"3E",X"1E",
		X"1A",X"2A",X"1E",X"30",X"00",X"42",X"1E",X"30",X"30",X"00",X"38",X"26",X"1A",X"24",X"3C",X"26",
		X"A2",X"AC",X"32",X"34",X"38",X"26",X"2E",X"16",X"00",X"20",X"26",X"38",X"1E",X"00",X"34",X"16",
		X"38",X"16",X"00",X"3A",X"1E",X"2C",X"1E",X"1A",X"1A",X"26",X"32",X"30",X"16",X"B8",X"C0",X"18",
		X"2C",X"16",X"1A",X"2A",X"00",X"42",X"26",X"1C",X"32",X"42",X"00",X"24",X"16",X"2C",X"2C",X"00",
		X"32",X"20",X"00",X"20",X"16",X"2E",X"9E",X"EE",X"20",X"38",X"1E",X"30",X"1A",X"A4",X"EE",X"22",
		X"1E",X"38",X"2E",X"16",X"B0",X"EB",X"3A",X"34",X"16",X"30",X"26",X"3A",X"A4",X"9A",X"3A",X"1E",
		X"2C",X"1E",X"1A",X"3C",X"00",X"1C",X"26",X"20",X"20",X"26",X"1A",X"3E",X"2C",X"3C",X"46",X"00",
		X"42",X"26",X"3C",X"24",X"00",X"38",X"26",X"22",X"24",X"3C",X"00",X"3A",X"3C",X"26",X"1A",X"AA",
		X"EE",X"20",X"38",X"1E",X"30",X"1A",X"A4",X"EE",X"22",X"1E",X"38",X"2E",X"16",X"B0",X"EB",X"3A",
		X"34",X"16",X"30",X"26",X"3A",X"A4",X"90",X"34",X"3E",X"3A",X"24",X"00",X"2C",X"1E",X"20",X"3C",
		X"00",X"3A",X"3C",X"26",X"1A",X"2A",X"00",X"16",X"30",X"1C",X"00",X"34",X"38",X"1E",X"3A",X"3A",
		X"00",X"3A",X"3C",X"16",X"38",X"3C",X"00",X"3C",X"32",X"00",X"18",X"1E",X"22",X"26",X"B0",X"EE",
		X"20",X"38",X"1E",X"30",X"1A",X"A4",X"EE",X"22",X"1E",X"38",X"2E",X"16",X"B0",X"EB",X"3A",X"34",
		X"16",X"30",X"26",X"3A",X"A4",X"8B",X"18",X"32",X"30",X"3E",X"BA",X"E8",X"3C",X"26",X"2E",X"1E",
		X"80",X"E0",X"1C",X"3E",X"38",X"1E",X"1E",X"80",X"E8",X"48",X"1E",X"26",X"3C",X"80",X"E4",X"3C",
		X"26",X"1E",X"2E",X"34",X"32",X"80",X"E8",X"42",X"16",X"40",X"1E",X"80",X"DC",X"30",X"26",X"40",
		X"1E",X"16",X"3E",X"80",X"E8",X"22",X"38",X"16",X"1C",X"80",X"E2",X"30",X"26",X"40",X"1E",X"2C",
		X"80",X"B2",X"3A",X"24",X"32",X"32",X"3C",X"00",X"00",X"00",X"00",X"00",X"3C",X"32",X"00",X"1A",
		X"32",X"2C",X"2C",X"1E",X"1A",X"3C",X"00",X"18",X"32",X"30",X"3E",X"BA",X"EE",X"20",X"38",X"1E",
		X"30",X"1A",X"A4",X"EB",X"3A",X"34",X"16",X"30",X"26",X"3A",X"A4",X"EE",X"22",X"1E",X"38",X"2E",
		X"16",X"B0",X"BA",X"42",X"16",X"40",X"1E",X"00",X"00",X"18",X"32",X"30",X"3E",X"3A",X"00",X"00",
		X"00",X"00",X"00",X"1C",X"26",X"20",X"20",X"26",X"1A",X"3E",X"2C",X"3C",X"C6",X"EE",X"20",X"38",
		X"1E",X"30",X"1A",X"A4",X"EB",X"3A",X"34",X"16",X"30",X"26",X"3A",X"A4",X"EE",X"22",X"1E",X"38",
		X"2E",X"16",X"B0",X"DC",X"26",X"30",X"3A",X"1E",X"38",X"3C",X"00",X"1A",X"32",X"26",X"30",X"BA",
		X"C1",X"26",X"30",X"3C",X"38",X"32",X"1C",X"3E",X"26",X"38",X"1E",X"00",X"2C",X"1E",X"3A",X"00",
		X"34",X"26",X"1E",X"1A",X"1E",X"BA",X"D6",X"22",X"1E",X"2C",X"1C",X"00",X"1E",X"26",X"30",X"42",
		X"1E",X"38",X"20",X"1E",X"B0",X"D6",X"26",X"30",X"3A",X"1E",X"38",X"3C",X"1E",X"00",X"20",X"26",
		X"1A",X"24",X"16",X"BA",X"E5",X"20",X"38",X"1E",X"1E",X"00",X"34",X"2C",X"16",X"C6",X"D6",X"04",
		X"00",X"1A",X"32",X"26",X"30",X"00",X"06",X"00",X"34",X"2C",X"16",X"46",X"BA",X"CD",X"04",X"00",
		X"34",X"26",X"1E",X"1A",X"1E",X"00",X"06",X"00",X"28",X"32",X"3E",X"1E",X"3E",X"38",X"BA",X"D0",
		X"04",X"00",X"2E",X"3E",X"1E",X"30",X"48",X"00",X"06",X"00",X"3A",X"34",X"26",X"1E",X"2C",X"9E",
		X"CD",X"04",X"00",X"2E",X"32",X"30",X"1E",X"1C",X"16",X"00",X"06",X"00",X"28",X"3E",X"1E",X"22",
		X"32",X"BA",X"D9",X"04",X"00",X"1A",X"32",X"26",X"30",X"00",X"04",X"00",X"34",X"2C",X"16",X"C6",
		X"D0",X"04",X"00",X"34",X"26",X"1E",X"1A",X"1E",X"00",X"04",X"00",X"28",X"32",X"3E",X"1E",X"3E",
		X"B8",X"D0",X"04",X"00",X"2E",X"3E",X"1E",X"30",X"48",X"1E",X"00",X"04",X"00",X"3A",X"34",X"26",
		X"1E",X"AC",X"D0",X"04",X"00",X"2E",X"32",X"30",X"1E",X"1C",X"16",X"00",X"04",X"00",X"28",X"3E",
		X"1E",X"22",X"B2",X"D6",X"06",X"00",X"1A",X"32",X"26",X"30",X"3A",X"00",X"04",X"00",X"34",X"2C",
		X"16",X"C6",X"CD",X"06",X"00",X"34",X"26",X"1E",X"1A",X"1E",X"3A",X"00",X"04",X"00",X"28",X"32",
		X"3E",X"1E",X"3E",X"B8",X"CD",X"06",X"00",X"2E",X"3E",X"1E",X"30",X"48",X"1E",X"30",X"00",X"04",
		X"00",X"3A",X"34",X"26",X"1E",X"AC",X"CD",X"06",X"00",X"2E",X"32",X"30",X"1E",X"1C",X"16",X"3A",
		X"00",X"04",X"00",X"28",X"3E",X"1E",X"22",X"B2",X"CD",X"50",X"00",X"16",X"3C",X"16",X"38",X"26",
		X"00",X"2E",X"1A",X"2E",X"2C",X"44",X"44",X"44",X"26",X"A6",X"E6",X"1A",X"38",X"1E",X"1C",X"26",
		X"3C",X"3A",X"80",X"A0",X"2A",X"38",X"1E",X"1C",X"26",X"3C",X"1E",X"80",X"A0",X"1A",X"38",X"1E",
		X"1C",X"26",X"3C",X"32",X"3A",X"80",X"D0",X"06",X"00",X"1A",X"38",X"1E",X"1C",X"26",X"3C",X"00",
		X"2E",X"26",X"30",X"26",X"2E",X"3E",X"AE",X"D6",X"06",X"00",X"28",X"1E",X"3E",X"44",X"00",X"2E",
		X"26",X"30",X"26",X"2E",X"3E",X"AE",X"D0",X"06",X"00",X"3A",X"34",X"26",X"1E",X"2C",X"1E",X"00",
		X"2E",X"26",X"30",X"26",X"2E",X"3E",X"AE",X"D3",X"06",X"00",X"28",X"3E",X"1E",X"22",X"32",X"3A",
		X"00",X"2E",X"26",X"30",X"26",X"2E",X"B2",X"BC",X"18",X"32",X"30",X"3E",X"3A",X"00",X"3A",X"34",
		X"26",X"1C",X"1E",X"38",X"00",X"1E",X"40",X"1E",X"38",X"46",X"80",X"CE",X"18",X"32",X"30",X"3E",
		X"3A",X"00",X"1A",X"24",X"16",X"36",X"3E",X"1E",X"80",X"CE",X"18",X"32",X"30",X"3E",X"3A",X"00",
		X"28",X"1E",X"1C",X"1E",X"80",X"C8",X"18",X"32",X"30",X"3E",X"3A",X"00",X"1A",X"16",X"1C",X"16",
		X"80",X"E0",X"2C",X"1E",X"40",X"1E",X"AC",X"DA",X"30",X"26",X"40",X"1E",X"16",X"BE",X"E2",X"22",
		X"38",X"16",X"9C",X"E0",X"30",X"26",X"40",X"1E",X"AC",X"E4",X"30",X"1E",X"44",X"3C",X"00",X"18",
		X"32",X"30",X"3E",X"3A",X"80",X"E8",X"20",X"38",X"1E",X"30",X"1A",X"A4",X"E8",X"22",X"1E",X"38",
		X"2E",X"16",X"B0",X"E8",X"3A",X"34",X"16",X"30",X"26",X"3A",X"A4",X"C0",X"2C",X"26",X"40",X"1E",
		X"3A",X"00",X"34",X"1E",X"38",X"00",X"22",X"16",X"2E",X"1E",X"80",X"E8",X"20",X"38",X"1E",X"30",
		X"1A",X"A4",X"E8",X"22",X"1E",X"38",X"2E",X"16",X"B0",X"E8",X"3A",X"34",X"16",X"30",X"26",X"3A",
		X"A4",X"C0",X"2E",X"16",X"44",X"00",X"3A",X"3C",X"16",X"38",X"3C",X"00",X"42",X"16",X"40",X"1E",
		X"80",X"E8",X"20",X"38",X"1E",X"30",X"1A",X"A4",X"E8",X"22",X"1E",X"38",X"2E",X"16",X"B0",X"E8",
		X"3A",X"34",X"16",X"30",X"26",X"3A",X"A4",X"C0",X"16",X"40",X"1E",X"38",X"16",X"22",X"1E",X"00",
		X"22",X"16",X"2E",X"1E",X"00",X"3C",X"26",X"2E",X"1E",X"80",X"E8",X"20",X"38",X"1E",X"30",X"1A",
		X"A4",X"E8",X"22",X"1E",X"38",X"2E",X"16",X"B0",X"E8",X"3A",X"34",X"16",X"30",X"26",X"3A",X"A4",
		X"D9",X"1C",X"1E",X"2E",X"32",X"30",X"3A",X"3C",X"38",X"16",X"3C",X"26",X"32",X"B0",X"F4",X"1E",
		X"16",X"3A",X"C6",X"EE",X"2E",X"1E",X"1C",X"26",X"3E",X"AE",X"F4",X"24",X"16",X"38",X"9C",X"C0",
		X"22",X"16",X"2E",X"1E",X"3A",X"00",X"34",X"2C",X"16",X"46",X"1E",X"9C",X"AC",X"24",X"32",X"2C",
		X"1C",X"00",X"20",X"26",X"38",X"1E",X"00",X"3C",X"24",X"1E",X"30",X"00",X"34",X"38",X"1E",X"3A",
		X"3A",X"00",X"3A",X"3C",X"16",X"38",X"3C",X"00",X"84",X"E8",X"20",X"32",X"38",X"00",X"3C",X"1E",
		X"3A",X"BC",X"D3",X"3C",X"32",X"00",X"1A",X"2C",X"1E",X"16",X"38",X"00",X"3A",X"1A",X"32",X"38",
		X"1E",X"BA",X"D6",X"3C",X"32",X"00",X"1A",X"2C",X"1E",X"16",X"38",X"00",X"3C",X"26",X"2E",X"1E",
		X"BA",X"B5",X"3C",X"32",X"00",X"1A",X"2C",X"1E",X"16",X"38",X"00",X"3A",X"1A",X"32",X"38",X"1E",
		X"3A",X"00",X"16",X"30",X"1C",X"00",X"3C",X"26",X"2E",X"1E",X"BA",X"BB",X"1E",X"16",X"38",X"32",
		X"2E",X"00",X"18",X"3E",X"3A",X"46",X"00",X"00",X"34",X"2C",X"1E",X"16",X"3A",X"1E",X"00",X"42",
		X"16",X"26",X"BC",X"C0",X"18",X"32",X"30",X"3E",X"3A",X"00",X"16",X"1C",X"1C",X"1E",X"38",X"80",
		X"C0",X"2C",X"1E",X"20",X"3C",X"00",X"2E",X"1E",X"1A",X"24",X"00",X"C4",X"C0",X"38",X"26",X"22",
		X"24",X"3C",X"00",X"2E",X"1E",X"1A",X"24",X"00",X"C4",X"BA",X"3C",X"16",X"22",X"00",X"22",X"38",
		X"3E",X"18",X"3A",X"3C",X"1E",X"16",X"2A",X"3A",X"00",X"20",X"32",X"38",X"00",X"34",X"32",X"26",
		X"30",X"3C",X"BA",X"AB",X"3A",X"24",X"32",X"32",X"3C",X"00",X"18",X"3E",X"22",X"3A",X"00",X"3C",
		X"24",X"1E",X"30",X"00",X"3C",X"16",X"22",X"00",X"22",X"38",X"3E",X"18",X"3A",X"3C",X"1E",X"16",
		X"2A",X"BA",X"9C",X"34",X"3E",X"3A",X"24",X"00",X"1E",X"22",X"22",X"3A",X"00",X"32",X"20",X"20",
		X"00",X"42",X"1E",X"18",X"00",X"18",X"1E",X"20",X"32",X"38",X"1E",X"00",X"3C",X"24",X"1E",X"46",
		X"00",X"24",X"16",X"3C",X"1A",X"A4",X"A8",X"3A",X"24",X"32",X"32",X"3C",X"00",X"22",X"38",X"1E",
		X"30",X"16",X"1C",X"1E",X"00",X"18",X"3E",X"22",X"3A",X"00",X"42",X"26",X"3C",X"24",X"00",X"1A",
		X"16",X"3E",X"3C",X"26",X"32",X"B0",X"A8",X"DE",X"08",X"DF",X"68",X"DF",X"C8",X"DF",X"A9",X"00",
		X"0A",X"A8",X"B9",X"46",X"E7",X"85",X"9B",X"B9",X"47",X"E7",X"85",X"9C",X"60",X"F3",X"00",X"78",
		X"8D",X"80",X"89",X"8D",X"C0",X"88",X"8D",X"80",X"88",X"A2",X"FF",X"9A",X"AD",X"00",X"78",X"29",
		X"10",X"F0",X"03",X"4C",X"18",X"90",X"78",X"A9",X"C0",X"8D",X"00",X"88",X"A9",X"00",X"A2",X"00",
		X"95",X"00",X"9D",X"00",X"01",X"9D",X"00",X"02",X"9D",X"00",X"03",X"9D",X"00",X"04",X"9D",X"00",
		X"05",X"9D",X"00",X"06",X"9D",X"00",X"07",X"9D",X"00",X"20",X"9D",X"00",X"21",X"9D",X"00",X"22",
		X"9D",X"00",X"23",X"9D",X"00",X"24",X"9D",X"00",X"25",X"9D",X"00",X"26",X"9D",X"00",X"27",X"E8",
		X"D0",X"CE",X"A9",X"69",X"8D",X"FF",X"07",X"8D",X"80",X"88",X"4C",X"D3",X"E8",X"48",X"8A",X"48",
		X"98",X"48",X"D8",X"AD",X"FF",X"07",X"C9",X"69",X"D0",X"06",X"20",X"B3",X"D6",X"4C",X"CA",X"E8",
		X"8D",X"0B",X"60",X"AD",X"08",X"60",X"8D",X"2E",X"06",X"8D",X"0B",X"68",X"AD",X"08",X"68",X"8D",
		X"2F",X"06",X"24",X"EF",X"10",X"11",X"A5",X"8C",X"F0",X"14",X"AD",X"00",X"78",X"29",X"10",X"F0",
		X"0D",X"A5",X"8D",X"F0",X"1D",X"D0",X"07",X"AD",X"20",X"04",X"C9",X"07",X"D0",X"14",X"AD",X"00",
		X"88",X"49",X"FF",X"29",X"60",X"F0",X"08",X"4D",X"2D",X"06",X"F0",X"06",X"8D",X"2C",X"06",X"8D",
		X"2D",X"06",X"E6",X"94",X"A5",X"19",X"85",X"18",X"A5",X"94",X"29",X"0F",X"D0",X"03",X"20",X"B3",
		X"D6",X"A5",X"00",X"C9",X"55",X"D0",X"03",X"4C",X"6F",X"E8",X"20",X"83",X"BD",X"20",X"64",X"D5",
		X"A5",X"99",X"4A",X"4A",X"85",X"19",X"A5",X"8A",X"0A",X"26",X"19",X"A5",X"8B",X"0A",X"26",X"19",
		X"A5",X"19",X"85",X"99",X"8D",X"00",X"88",X"AD",X"20",X"01",X"D0",X"23",X"A5",X"00",X"C9",X"AA",
		X"F0",X"1D",X"AD",X"00",X"78",X"29",X"40",X"D0",X"0B",X"E6",X"81",X"A5",X"81",X"C9",X"0A",X"D0",
		X"0E",X"8D",X"80",X"88",X"A9",X"00",X"85",X"81",X"A9",X"AA",X"85",X"00",X"8D",X"40",X"88",X"A5",
		X"18",X"85",X"19",X"A5",X"FC",X"D0",X"50",X"CE",X"D0",X"03",X"D0",X"4B",X"A9",X"F6",X"8D",X"D0",
		X"03",X"CE",X"22",X"04",X"10",X"05",X"A9",X"00",X"8D",X"22",X"04",X"24",X"EF",X"10",X"1E",X"CE",
		X"24",X"04",X"10",X"19",X"A9",X"1E",X"8D",X"24",X"04",X"AD",X"2F",X"06",X"29",X"03",X"AA",X"AD",
		X"2B",X"06",X"DD",X"25",X"9C",X"90",X"06",X"38",X"E9",X"04",X"8D",X"2B",X"06",X"E6",X"79",X"E6",
		X"76",X"D0",X"06",X"E6",X"77",X"D0",X"02",X"E6",X"78",X"24",X"EF",X"30",X"0A",X"E6",X"7C",X"D0",
		X"06",X"E6",X"7D",X"D0",X"02",X"E6",X"7E",X"8D",X"80",X"89",X"8D",X"C0",X"88",X"68",X"A8",X"68",
		X"AA",X"68",X"40",X"A2",X"11",X"9A",X"8A",X"86",X"00",X"A0",X"00",X"A2",X"01",X"C8",X"B9",X"00",
		X"00",X"D0",X"21",X"E8",X"D0",X"F7",X"BA",X"8A",X"8D",X"80",X"89",X"C8",X"59",X"00",X"00",X"D0",
		X"13",X"8A",X"A2",X"00",X"96",X"00",X"C8",X"D0",X"05",X"0A",X"A2",X"00",X"B0",X"4B",X"AA",X"9A",
		X"96",X"00",X"D0",X"D7",X"AA",X"8A",X"A0",X"82",X"29",X"0F",X"F0",X"02",X"A0",X"12",X"8A",X"A2",
		X"82",X"29",X"F0",X"F0",X"02",X"A2",X"12",X"98",X"9A",X"AA",X"8E",X"00",X"60",X"A2",X"A8",X"8E",
		X"01",X"60",X"A0",X"0C",X"A2",X"64",X"2C",X"00",X"78",X"30",X"FB",X"2C",X"00",X"78",X"10",X"FB",
		X"8D",X"80",X"89",X"CA",X"D0",X"F0",X"C0",X"05",X"D0",X"03",X"8E",X"01",X"60",X"88",X"D0",X"E4",
		X"4A",X"B0",X"03",X"BA",X"D0",X"D4",X"4C",X"00",X"EA",X"A2",X"FF",X"9A",X"A2",X"00",X"8A",X"95",
		X"00",X"E8",X"D0",X"FB",X"A8",X"A9",X"01",X"85",X"01",X"A2",X"11",X"B1",X"00",X"D0",X"27",X"8A",
		X"91",X"00",X"51",X"00",X"D0",X"20",X"8A",X"0A",X"AA",X"90",X"F5",X"C8",X"D0",X"EB",X"8D",X"80",
		X"89",X"E6",X"01",X"A6",X"01",X"E0",X"04",X"90",X"E0",X"A9",X"20",X"E0",X"20",X"90",X"D8",X"E0",
		X"28",X"90",X"D6",X"4C",X"07",X"EA",X"A6",X"01",X"E0",X"20",X"85",X"02",X"90",X"03",X"8A",X"E9",
		X"1C",X"4A",X"4A",X"29",X"07",X"A8",X"A5",X"02",X"84",X"00",X"85",X"01",X"A9",X"01",X"85",X"02",
		X"A2",X"A8",X"A0",X"82",X"A5",X"00",X"D0",X"08",X"A5",X"01",X"29",X"0F",X"F0",X"02",X"A0",X"12",
		X"8E",X"01",X"60",X"8C",X"00",X"60",X"A9",X"09",X"C0",X"12",X"F0",X"02",X"A9",X"01",X"A8",X"A2",
		X"00",X"2C",X"00",X"78",X"30",X"FB",X"2C",X"00",X"78",X"10",X"FB",X"8D",X"80",X"89",X"CA",X"D0",
		X"F0",X"88",X"D0",X"ED",X"8E",X"01",X"60",X"A0",X"09",X"2C",X"00",X"78",X"30",X"FB",X"2C",X"00",
		X"78",X"10",X"FB",X"8D",X"80",X"89",X"CA",X"D0",X"F0",X"88",X"D0",X"ED",X"A5",X"00",X"D0",X"08",
		X"A5",X"01",X"4A",X"4A",X"4A",X"4A",X"85",X"01",X"C6",X"02",X"F0",X"A4",X"C6",X"00",X"10",X"9C",
		X"8D",X"80",X"89",X"A9",X"FF",X"85",X"D4",X"A9",X"00",X"AA",X"9D",X"00",X"01",X"9D",X"00",X"02",
		X"9D",X"00",X"03",X"CA",X"D0",X"F4",X"A8",X"85",X"C0",X"A9",X"30",X"85",X"C1",X"A9",X"10",X"85",
		X"C2",X"8A",X"51",X"C0",X"C8",X"D0",X"FB",X"E6",X"C1",X"8D",X"80",X"89",X"C6",X"C2",X"D0",X"F2",
		X"95",X"CB",X"E8",X"F0",X"18",X"A5",X"C1",X"C9",X"60",X"D0",X"04",X"A9",X"90",X"85",X"C1",X"C9",
		X"F0",X"90",X"D8",X"A2",X"FF",X"A9",X"28",X"85",X"C1",X"A9",X"08",X"D0",X"D2",X"A5",X"CA",X"05",
		X"CB",X"F0",X"0A",X"A9",X"F0",X"A2",X"A2",X"8D",X"04",X"60",X"8E",X"05",X"60",X"A2",X"05",X"AD",
		X"0A",X"68",X"CD",X"0A",X"68",X"D0",X"05",X"CA",X"10",X"F8",X"85",X"D5",X"A2",X"05",X"AD",X"0A",
		X"60",X"CD",X"0A",X"60",X"D0",X"05",X"CA",X"10",X"F8",X"85",X"D6",X"58",X"20",X"A9",X"D6",X"A0",
		X"02",X"AD",X"2D",X"01",X"F0",X"0A",X"85",X"D7",X"20",X"89",X"D6",X"A0",X"00",X"8C",X"2D",X"01",
		X"84",X"C9",X"4C",X"D8",X"EC",X"AD",X"2E",X"01",X"0D",X"2B",X"01",X"D0",X"0C",X"20",X"A9",X"D6",
		X"AD",X"2D",X"01",X"85",X"D7",X"A9",X"02",X"85",X"C9",X"60",X"A0",X"A7",X"A9",X"04",X"20",X"EF",
		X"D7",X"A2",X"20",X"A9",X"5E",X"20",X"E3",X"D7",X"A9",X"48",X"A2",X"40",X"A0",X"00",X"20",X"1B",
		X"D8",X"20",X"42",X"EC",X"A9",X"01",X"20",X"12",X"D8",X"A2",X"46",X"86",X"C2",X"A2",X"09",X"B5",
		X"CA",X"F0",X"1B",X"86",X"C1",X"20",X"F9",X"D7",X"A6",X"C2",X"8A",X"38",X"E9",X"08",X"85",X"C2",
		X"A9",X"F6",X"A0",X"00",X"20",X"1B",X"D8",X"A5",X"C1",X"20",X"C3",X"ED",X"A6",X"C1",X"CA",X"10",
		X"DE",X"20",X"F9",X"D7",X"A9",X"F6",X"A2",X"58",X"A0",X"00",X"20",X"1B",X"D8",X"A2",X"03",X"86",
		X"C1",X"A6",X"C1",X"A0",X"00",X"B5",X"D4",X"F0",X"03",X"BC",X"CA",X"EB",X"B9",X"C4",X"5D",X"BE",
		X"C5",X"5D",X"20",X"FD",X"D7",X"C6",X"C1",X"10",X"E8",X"20",X"A8",X"EC",X"60",X"A2",X"FE",X"A9",
		X"5E",X"4C",X"E3",X"D7",X"E6",X"C4",X"10",X"06",X"A9",X"00",X"85",X"C4",X"E6",X"C2",X"A5",X"C2",
		X"29",X"07",X"AA",X"BC",X"69",X"EB",X"A9",X"00",X"99",X"F1",X"67",X"BC",X"6A",X"EB",X"BD",X"73",
		X"EB",X"99",X"F0",X"67",X"A9",X"A8",X"99",X"F1",X"67",X"A2",X"04",X"A9",X"5F",X"20",X"E3",X"D7",
		X"20",X"F9",X"D7",X"A4",X"C4",X"A5",X"C2",X"29",X"07",X"D0",X"04",X"A9",X"01",X"85",X"C2",X"20",
		X"12",X"D8",X"A2",X"22",X"A9",X"5E",X"4C",X"E3",X"D7",X"16",X"00",X"10",X"02",X"12",X"04",X"14",
		X"06",X"16",X"00",X"10",X"10",X"40",X"40",X"90",X"90",X"FF",X"FF",X"A2",X"20",X"A9",X"5E",X"20",
		X"E3",X"D7",X"A0",X"06",X"84",X"C2",X"20",X"F9",X"D7",X"A4",X"C2",X"B9",X"BC",X"EB",X"BE",X"C3",
		X"EB",X"20",X"1B",X"D8",X"A5",X"C2",X"49",X"FF",X"29",X"07",X"A8",X"20",X"EF",X"D7",X"A5",X"C2",
		X"D0",X"07",X"A2",X"C0",X"A9",X"5E",X"4C",X"AD",X"EB",X"A2",X"BA",X"A9",X"5E",X"20",X"E3",X"D7",
		X"C6",X"C2",X"10",X"D2",X"A2",X"DE",X"A9",X"5E",X"20",X"E3",X"D7",X"60",X"DE",X"9D",X"1F",X"9D",
		X"DE",X"1F",X"DE",X"F4",X"D8",X"D8",X"10",X"D8",X"10",X"10",X"38",X"34",X"36",X"1E",X"20",X"F9",
		X"D7",X"A9",X"01",X"20",X"10",X"D8",X"A2",X"06",X"86",X"C1",X"A4",X"C1",X"A9",X"90",X"BE",X"1D",
		X"EC",X"20",X"1B",X"D8",X"A2",X"F6",X"A9",X"5E",X"20",X"E3",X"D7",X"C6",X"C1",X"10",X"EB",X"A2",
		X"06",X"86",X"C1",X"A4",X"C1",X"B9",X"24",X"EC",X"A2",X"6B",X"20",X"1B",X"D8",X"A2",X"EE",X"A9",
		X"5E",X"20",X"E3",X"D7",X"C6",X"C1",X"10",X"EB",X"AD",X"00",X"88",X"29",X"20",X"D0",X"09",X"06",
		X"C0",X"90",X"02",X"E6",X"C5",X"4C",X"1C",X"EC",X"A9",X"20",X"85",X"C0",X"60",X"B2",X"CC",X"E6",
		X"00",X"1A",X"34",X"4E",X"AC",X"C8",X"E4",X"00",X"1C",X"38",X"54",X"A2",X"46",X"A9",X"5F",X"20",
		X"E3",X"D7",X"A9",X"20",X"85",X"C0",X"A2",X"3A",X"A9",X"5F",X"20",X"E3",X"D7",X"C6",X"C0",X"10",
		X"F5",X"60",X"A2",X"0F",X"86",X"C1",X"8D",X"0B",X"60",X"EA",X"AD",X"08",X"60",X"85",X"C3",X"8D",
		X"0B",X"68",X"EA",X"AD",X"08",X"68",X"48",X"29",X"01",X"18",X"20",X"C3",X"ED",X"46",X"C3",X"68",
		X"6A",X"C6",X"C1",X"10",X"F1",X"A9",X"D0",X"A0",X"00",X"A2",X"F8",X"20",X"1B",X"D8",X"A2",X"07",
		X"86",X"C1",X"A9",X"78",X"85",X"C6",X"A9",X"07",X"85",X"C7",X"A9",X"00",X"85",X"C5",X"A8",X"B1",
		X"C5",X"49",X"FF",X"29",X"7F",X"48",X"29",X"01",X"18",X"20",X"C3",X"ED",X"68",X"6A",X"C8",X"C6",
		X"C7",X"10",X"F2",X"A9",X"D0",X"A0",X"00",X"A2",X"F8",X"20",X"1B",X"D8",X"A5",X"C6",X"18",X"69",
		X"08",X"85",X"C6",X"C9",X"90",X"90",X"CF",X"60",X"84",X"C3",X"AD",X"00",X"78",X"29",X"0F",X"85",
		X"C0",X"AD",X"00",X"80",X"29",X"1F",X"85",X"C1",X"AD",X"00",X"88",X"29",X"7F",X"85",X"C2",X"A5",
		X"C0",X"09",X"10",X"25",X"C1",X"09",X"60",X"25",X"C2",X"49",X"7F",X"F0",X"07",X"69",X"40",X"8D",
		X"00",X"60",X"A0",X"A4",X"8C",X"01",X"60",X"60",X"A2",X"18",X"2C",X"00",X"78",X"10",X"FB",X"2C",
		X"00",X"78",X"30",X"FB",X"CA",X"10",X"F3",X"E6",X"D9",X"2C",X"00",X"78",X"50",X"FB",X"A9",X"00",
		X"8D",X"11",X"00",X"A9",X"20",X"8D",X"12",X"00",X"AD",X"00",X"78",X"49",X"FF",X"29",X"24",X"F0",
		X"26",X"06",X"C8",X"90",X"1F",X"AD",X"00",X"88",X"29",X"40",X"D0",X"06",X"20",X"8E",X"ED",X"20",
		X"FF",X"ED",X"E6",X"C9",X"E6",X"C9",X"A9",X"00",X"A2",X"06",X"9D",X"00",X"60",X"9D",X"00",X"68",
		X"CA",X"CA",X"10",X"F6",X"4C",X"2B",X"ED",X"A9",X"20",X"85",X"C8",X"A5",X"C9",X"C9",X"0C",X"D0",
		X"0E",X"A5",X"C5",X"29",X"07",X"D0",X"02",X"A9",X"01",X"09",X"C0",X"A8",X"4C",X"41",X"ED",X"A0",
		X"A7",X"A9",X"04",X"20",X"EF",X"D7",X"A2",X"20",X"A9",X"5E",X"20",X"E3",X"D7",X"20",X"7B",X"ED",
		X"20",X"F9",X"D7",X"20",X"A6",X"D7",X"A9",X"C0",X"85",X"DA",X"8D",X"40",X"88",X"8D",X"80",X"89",
		X"AD",X"00",X"78",X"29",X"10",X"D0",X"03",X"4C",X"D8",X"EC",X"4C",X"6A",X"ED",X"94",X"EA",X"A9",
		X"EA",X"1C",X"EB",X"23",X"EB",X"2A",X"EC",X"7A",X"EB",X"CD",X"EB",X"A6",X"C9",X"E0",X"0E",X"90",
		X"04",X"A2",X"02",X"86",X"C9",X"BD",X"6E",X"ED",X"48",X"BD",X"6D",X"ED",X"48",X"60",X"A9",X"00",
		X"8D",X"0F",X"60",X"8D",X"0F",X"68",X"A9",X"07",X"8D",X"0F",X"60",X"8D",X"0F",X"68",X"A2",X"0F",
		X"A9",X"00",X"9D",X"00",X"60",X"9D",X"00",X"68",X"CA",X"10",X"F7",X"A9",X"00",X"8D",X"08",X"60",
		X"A2",X"00",X"8E",X"08",X"68",X"60",X"48",X"08",X"4A",X"4A",X"4A",X"4A",X"28",X"20",X"C3",X"ED",
		X"68",X"29",X"0F",X"90",X"05",X"29",X"0F",X"F0",X"08",X"18",X"0A",X"08",X"20",X"DD",X"ED",X"28",
		X"60",X"AE",X"C4",X"5D",X"AD",X"C5",X"5D",X"08",X"20",X"E8",X"ED",X"28",X"60",X"A8",X"BE",X"C6",
		X"5D",X"B9",X"C7",X"5D",X"20",X"E8",X"ED",X"60",X"A0",X"01",X"91",X"11",X"88",X"8A",X"91",X"11",
		X"AD",X"11",X"00",X"18",X"69",X"02",X"8D",X"11",X"00",X"90",X"03",X"EE",X"12",X"00",X"60",X"78",
		X"D8",X"A9",X"FF",X"85",X"02",X"D0",X"11",X"A5",X"00",X"F0",X"0D",X"AD",X"00",X"78",X"29",X"40",
		X"F0",X"06",X"8D",X"80",X"88",X"8D",X"40",X"88",X"8D",X"80",X"89",X"AD",X"00",X"78",X"29",X"10",
		X"D0",X"FE",X"AD",X"00",X"80",X"18",X"2A",X"2A",X"2A",X"2A",X"49",X"FF",X"29",X"07",X"85",X"00",
		X"A5",X"00",X"C5",X"02",X"F0",X"D1",X"85",X"02",X"AA",X"F0",X"21",X"A9",X"C7",X"8D",X"00",X"20",
		X"A9",X"60",X"8D",X"01",X"20",X"BC",X"B0",X"EE",X"BD",X"B8",X"EE",X"AA",X"B9",X"C0",X"EE",X"9D",
		X"02",X"20",X"88",X"CA",X"10",X"F6",X"8D",X"80",X"88",X"4C",X"07",X"EE",X"A9",X"20",X"85",X"04",
		X"A9",X"00",X"85",X"03",X"85",X"01",X"A8",X"A9",X"08",X"85",X"00",X"18",X"A5",X"01",X"91",X"03",
		X"69",X"05",X"85",X"01",X"C8",X"D0",X"F4",X"E6",X"04",X"C6",X"00",X"D0",X"EE",X"A0",X"07",X"A2",
		X"00",X"A9",X"11",X"9D",X"80",X"27",X"9D",X"80",X"26",X"48",X"8A",X"18",X"69",X"10",X"AA",X"68",
		X"88",X"10",X"F0",X"8D",X"B2",X"26",X"8D",X"B2",X"27",X"8D",X"DE",X"26",X"8D",X"EE",X"26",X"8D",
		X"DE",X"27",X"8D",X"EE",X"27",X"A9",X"80",X"8D",X"FE",X"26",X"8D",X"FE",X"27",X"4C",X"56",X"EE",
		X"01",X"01",X"15",X"2B",X"45",X"71",X"01",X"01",X"01",X"01",X"13",X"15",X"19",X"2B",X"01",X"01",
		X"00",X"20",X"40",X"80",X"00",X"71",X"80",X"01",X"00",X"22",X"40",X"80",X"00",X"60",X"80",X"1E",
		X"00",X"3E",X"40",X"80",X"00",X"20",X"40",X"80",X"00",X"71",X"80",X"01",X"00",X"22",X"07",X"E0",
		X"00",X"20",X"40",X"80",X"80",X"1E",X"00",X"3E",X"40",X"80",X"00",X"20",X"40",X"80",X"00",X"71",
		X"80",X"01",X"00",X"22",X"07",X"E0",X"00",X"20",X"40",X"80",X"80",X"1E",X"00",X"3E",X"40",X"80",
		X"2F",X"51",X"40",X"80",X"00",X"20",X"40",X"80",X"00",X"71",X"80",X"01",X"00",X"22",X"07",X"E0",
		X"00",X"20",X"40",X"80",X"80",X"1E",X"00",X"3E",X"40",X"80",X"2F",X"51",X"40",X"80",X"11",X"A0",
		X"20",X"51",X"40",X"80",X"00",X"20",X"13",X"A0",X"00",X"C0",X"15",X"A0",X"00",X"C0",X"2F",X"40",
		X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5F",X"E7",X"5F",X"E7",X"BD",X"E7");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
