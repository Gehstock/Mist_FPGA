`define BUILD_DATE "180913"
`define BUILD_TIME "214058"
