library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity cclimber_program is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of cclimber_program is
	type rom is array(0 to  20479) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"EA",X"AE",X"FF",X"EF",X"23",X"00",X"A0",X"33",X"01",X"A0",X"23",X"02",X"A0",X"33",X"07",X"A0",
		X"C2",X"AC",X"00",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",
		X"2B",X"7C",X"80",X"B2",X"93",X"B3",X"0B",X"3B",X"81",X"80",X"E7",X"93",X"B8",X"0B",X"C2",X"B3",
		X"0B",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",
		X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",
		X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",
		X"41",X"10",X"41",X"10",X"41",X"10",X"E1",X"3B",X"00",X"B8",X"EE",X"33",X"00",X"A0",X"A1",X"97",
		X"D9",X"00",X"2B",X"00",X"B8",X"EF",X"23",X"00",X"A0",X"70",X"FF",X"00",X"77",X"40",X"80",X"64",
		X"00",X"84",X"8D",X"43",X"01",X"EF",X"23",X"44",X"80",X"70",X"62",X"80",X"63",X"40",X"8D",X"CB",
		X"00",X"97",X"37",X"02",X"EE",X"33",X"00",X"A0",X"EE",X"33",X"44",X"80",X"74",X"5D",X"80",X"7E",
		X"04",X"76",X"00",X"77",X"7D",X"30",X"FA",X"76",X"20",X"97",X"37",X"02",X"74",X"00",X"80",X"44",
		X"00",X"04",X"63",X"00",X"72",X"4A",X"3B",X"F2",X"61",X"F8",X"30",X"00",X"84",X"7E",X"07",X"C2",
		X"08",X"7E",X"FF",X"C2",X"09",X"DD",X"A3",X"03",X"C2",X"72",X"00",X"70",X"5D",X"80",X"6B",X"04",
		X"63",X"20",X"72",X"2C",X"61",X"FA",X"63",X"40",X"9D",X"E5",X"85",X"C5",X"A5",X"CD",X"A5",X"ED",
		X"A5",X"DD",X"4A",X"01",X"2B",X"00",X"B8",X"64",X"00",X"84",X"2B",X"7A",X"80",X"AE",X"04",X"30",
		X"03",X"33",X"72",X"80",X"41",X"70",X"45",X"80",X"21",X"6B",X"E7",X"93",X"00",X"01",X"72",X"60",
		X"8D",X"63",X"01",X"DD",X"00",X"40",X"2B",X"75",X"80",X"E7",X"61",X"23",X"2B",X"00",X"B8",X"9F",
		X"22",X"30",X"07",X"7E",X"01",X"33",X"B4",X"82",X"0D",X"15",X"2B",X"B4",X"82",X"E7",X"69",X"0F",
		X"74",X"C0",X"4C",X"27",X"24",X"80",X"6B",X"84",X"23",X"27",X"80",X"EF",X"23",X"B4",X"82",X"DD",
		X"E3",X"01",X"2B",X"73",X"80",X"F3",X"01",X"93",X"85",X"00",X"8D",X"FC",X"01",X"DD",X"FC",X"01",
		X"C2",X"37",X"02",X"70",X"89",X"03",X"77",X"42",X"80",X"C8",X"E1",X"2F",X"40",X"80",X"6D",X"AE",
		X"FF",X"38",X"0E",X"44",X"49",X"80",X"7C",X"4C",X"EA",X"70",X"04",X"00",X"38",X"BF",X"36",X"77",
		X"33",X"B0",X"9D",X"3B",X"00",X"B8",X"F6",X"01",X"93",X"CD",X"01",X"3B",X"00",X"B8",X"F6",X"02",
		X"93",X"D8",X"01",X"3B",X"71",X"80",X"E7",X"9D",X"2B",X"77",X"80",X"B2",X"69",X"20",X"2B",X"72",
		X"80",X"AE",X"50",X"21",X"09",X"06",X"2B",X"7A",X"80",X"C4",X"32",X"33",X"72",X"80",X"EE",X"33",
		X"71",X"80",X"2B",X"75",X"80",X"B2",X"D4",X"EF",X"23",X"44",X"80",X"97",X"72",X"00",X"2B",X"79",
		X"80",X"68",X"23",X"79",X"80",X"06",X"EE",X"33",X"71",X"80",X"2B",X"78",X"80",X"E9",X"D4",X"7E",
		X"00",X"33",X"79",X"80",X"2B",X"72",X"80",X"AE",X"50",X"21",X"06",X"D3",X"01",X"72",X"23",X"72",
		X"80",X"3B",X"75",X"80",X"E7",X"95",X"EE",X"33",X"44",X"80",X"C2",X"72",X"00",X"7E",X"00",X"33",
		X"77",X"80",X"6B",X"01",X"23",X"71",X"80",X"C8",X"6B",X"01",X"23",X"77",X"80",X"7E",X"01",X"33",
		X"71",X"80",X"9D",X"02",X"0A",X"70",X"67",X"80",X"10",X"5D",X"80",X"EF",X"FB",X"38",X"03",X"24",
		X"61",X"04",X"0B",X"F3",X"EF",X"13",X"72",X"42",X"14",X"30",X"F0",X"C8",X"74",X"5D",X"80",X"3B",
		X"45",X"80",X"F6",X"00",X"FF",X"00",X"61",X"04",X"7B",X"A6",X"40",X"37",X"72",X"3B",X"45",X"80",
		X"F6",X"03",X"FF",X"03",X"61",X"04",X"7B",X"A6",X"40",X"37",X"72",X"3B",X"45",X"80",X"F6",X"00",
		X"FF",X"00",X"61",X"04",X"7B",X"A6",X"40",X"37",X"72",X"3B",X"45",X"80",X"F6",X"01",X"FF",X"00",
		X"61",X"04",X"7B",X"A6",X"40",X"37",X"9D",X"3B",X"00",X"B8",X"2B",X"44",X"80",X"B2",X"61",X"32",
		X"6B",X"FF",X"23",X"40",X"80",X"EF",X"23",X"00",X"A0",X"7E",X"01",X"33",X"00",X"A0",X"54",X"00",
		X"0A",X"70",X"5D",X"80",X"7B",X"F3",X"30",X"30",X"05",X"6B",X"F6",X"C0",X"61",X"07",X"72",X"5C",
		X"14",X"30",X"F1",X"09",X"E0",X"EF",X"23",X"00",X"A0",X"3D",X"23",X"40",X"80",X"6B",X"F6",X"80",
		X"69",X"20",X"7F",X"40",X"80",X"44",X"49",X"80",X"7C",X"4C",X"5B",X"77",X"53",X"BF",X"A9",X"ED",
		X"B5",X"CD",X"B5",X"E0",X"81",X"C0",X"EE",X"33",X"00",X"A0",X"6B",X"01",X"23",X"00",X"A0",X"B0",
		X"AD",X"41",X"63",X"80",X"7F",X"40",X"80",X"44",X"95",X"03",X"7C",X"4C",X"5B",X"77",X"53",X"BF",
		X"A9",X"2F",X"40",X"80",X"EA",X"2F",X"42",X"80",X"18",X"4C",X"5B",X"77",X"53",X"BF",X"EE",X"33",
		X"00",X"A0",X"6B",X"01",X"23",X"00",X"A0",X"E8",X"E1",X"EF",X"23",X"00",X"A0",X"B0",X"E1",X"D5",
		X"C1",X"F5",X"C9",X"F5",X"E9",X"F5",X"E1",X"3B",X"44",X"80",X"E7",X"09",X"1D",X"B0",X"8D",X"4A",
		X"01",X"64",X"00",X"84",X"7F",X"40",X"80",X"44",X"67",X"80",X"18",X"37",X"7F",X"40",X"80",X"44",
		X"5D",X"80",X"18",X"6B",X"F7",X"10",X"76",X"97",X"37",X"02",X"EE",X"33",X"00",X"A0",X"6B",X"01",
		X"23",X"00",X"A0",X"B0",X"D7",X"01",X"2D",X"0E",X"E1",X"70",X"00",X"01",X"A5",X"E0",X"7A",X"79",
		X"A4",X"30",X"F9",X"B0",X"0D",X"EE",X"E9",X"E0",X"C9",X"E0",X"B5",X"90",X"95",X"B0",X"9D",X"EF",
		X"23",X"00",X"A0",X"2F",X"40",X"80",X"10",X"5D",X"80",X"4C",X"7B",X"F3",X"7F",X"37",X"C2",X"37",
		X"02",X"E5",X"EE",X"33",X"00",X"A0",X"A1",X"E5",X"85",X"C5",X"A5",X"CD",X"A5",X"ED",X"A5",X"DD",
		X"4A",X"01",X"30",X"00",X"84",X"70",X"5D",X"80",X"43",X"00",X"5E",X"4C",X"7B",X"A6",X"20",X"37",
		X"C2",X"37",X"02",X"E5",X"EE",X"33",X"00",X"A0",X"A1",X"E5",X"85",X"C5",X"A5",X"CD",X"A5",X"ED",
		X"A5",X"DD",X"4A",X"01",X"30",X"00",X"84",X"70",X"5D",X"80",X"43",X"00",X"5E",X"4C",X"7B",X"A6",
		X"40",X"37",X"C2",X"37",X"02",X"E5",X"EE",X"33",X"00",X"A0",X"A1",X"E5",X"85",X"C5",X"A5",X"CD",
		X"A5",X"ED",X"A5",X"DD",X"4A",X"01",X"30",X"00",X"84",X"70",X"5D",X"80",X"43",X"00",X"5E",X"4C",
		X"7B",X"F3",X"DF",X"37",X"C2",X"37",X"02",X"C7",X"FB",X"20",X"10",X"90",X"13",X"40",X"1B",X"10",
		X"28",X"72",X"05",X"54",X"04",X"E0",X"83",X"A8",X"83",X"70",X"83",X"38",X"83",X"E0",X"83",X"00",
		X"83",X"C7",X"F3",X"10",X"2B",X"00",X"B0",X"F3",X"03",X"D3",X"03",X"33",X"7E",X"80",X"2B",X"00",
		X"B8",X"F3",X"10",X"30",X"07",X"7E",X"00",X"33",X"7C",X"80",X"0D",X"05",X"6B",X"01",X"23",X"7C",
		X"80",X"3B",X"00",X"B0",X"F6",X"04",X"61",X"07",X"6B",X"00",X"23",X"76",X"80",X"09",X"05",X"7E",
		X"01",X"33",X"76",X"80",X"2B",X"00",X"B0",X"F3",X"40",X"30",X"07",X"7E",X"03",X"33",X"7D",X"80",
		X"0D",X"05",X"6B",X"05",X"23",X"7D",X"80",X"3B",X"00",X"B0",X"1A",X"5A",X"1A",X"5A",X"F6",X"03",
		X"D6",X"01",X"23",X"78",X"80",X"3B",X"00",X"B0",X"1A",X"5A",X"1A",X"5A",X"1A",X"5A",X"F6",X"03",
		X"D6",X"01",X"23",X"7A",X"80",X"70",X"95",X"80",X"17",X"05",X"1F",X"0A",X"C9",X"70",X"3E",X"04",
		X"C9",X"6B",X"00",X"37",X"72",X"CD",X"72",X"5D",X"61",X"F6",X"72",X"77",X"72",X"77",X"14",X"30",
		X"E9",X"70",X"83",X"80",X"17",X"05",X"63",X"02",X"72",X"76",X"00",X"77",X"63",X"00",X"72",X"55",
		X"61",X"F4",X"2B",X"7A",X"80",X"AE",X"04",X"95",X"23",X"72",X"80",X"C8",X"C7",X"FB",X"30",X"31",
		X"32",X"33",X"34",X"35",X"36",X"37",X"52",X"52",X"C7",X"F3",X"7B",X"13",X"72",X"42",X"5A",X"3D",
		X"F1",X"30",X"F7",X"C8",X"41",X"E5",X"A5",X"70",X"22",X"81",X"7B",X"D3",X"01",X"37",X"B5",X"B0",
		X"41",X"09",X"F1",X"70",X"00",X"9C",X"54",X"00",X"04",X"76",X"0A",X"77",X"5A",X"6D",X"B4",X"30",
		X"F8",X"C8",X"41",X"ED",X"A5",X"CD",X"A5",X"E5",X"85",X"C5",X"A5",X"C5",X"C9",X"E0",X"74",X"00",
		X"90",X"ED",X"74",X"00",X"9C",X"50",X"20",X"00",X"C9",X"6B",X"01",X"B2",X"69",X"06",X"5C",X"ED",
		X"5C",X"2C",X"61",X"FA",X"C9",X"1A",X"02",X"02",X"00",X"58",X"E9",X"58",X"C9",X"12",X"00",X"CD",
		X"72",X"CD",X"72",X"CD",X"72",X"CD",X"7B",X"00",X"FF",X"FF",X"69",X"10",X"76",X"6D",X"FF",X"FF",
		X"69",X"03",X"E9",X"65",X"00",X"77",X"C9",X"77",X"E9",X"77",X"0D",X"E9",X"B5",X"90",X"95",X"B0",
		X"C9",X"E0",X"E9",X"E0",X"9D",X"10",X"E9",X"F5",X"C9",X"F5",X"E1",X"D5",X"C1",X"F5",X"C1",X"CD",
		X"B5",X"70",X"00",X"90",X"E9",X"70",X"00",X"9C",X"54",X"20",X"00",X"CD",X"7B",X"01",X"E7",X"38",
		X"06",X"58",X"E9",X"58",X"7D",X"30",X"FA",X"CD",X"0F",X"02",X"17",X"00",X"5C",X"ED",X"5C",X"CD",
		X"07",X"00",X"C9",X"1A",X"05",X"CD",X"53",X"04",X"C9",X"4B",X"03",X"9F",X"11",X"38",X"07",X"1B",
		X"F6",X"0F",X"76",X"42",X"0D",X"08",X"0B",X"5A",X"1A",X"5A",X"1A",X"F3",X"0F",X"37",X"3D",X"AE",
		X"FF",X"38",X"03",X"ED",X"35",X"00",X"E9",X"77",X"72",X"5D",X"61",X"DF",X"B5",X"90",X"95",X"B0",
		X"C9",X"E0",X"E9",X"E0",X"9D",X"10",X"74",X"00",X"90",X"50",X"00",X"04",X"63",X"52",X"72",X"5F",
		X"3D",X"F4",X"61",X"F8",X"41",X"70",X"00",X"98",X"54",X"A0",X"00",X"76",X"00",X"77",X"5A",X"6D",
		X"B4",X"30",X"F8",X"DD",X"47",X"05",X"9D",X"10",X"74",X"00",X"88",X"50",X"00",X"01",X"63",X"00",
		X"72",X"5F",X"3D",X"F4",X"61",X"F8",X"74",X"DC",X"98",X"02",X"04",X"76",X"00",X"77",X"14",X"30",
		X"FA",X"C8",X"41",X"70",X"30",X"81",X"54",X"C0",X"01",X"76",X"00",X"77",X"5A",X"6D",X"B4",X"30",
		X"F8",X"C8",X"41",X"7E",X"01",X"33",X"44",X"80",X"2B",X"73",X"80",X"B2",X"93",X"5F",X"06",X"02",
		X"00",X"3B",X"72",X"80",X"E7",X"38",X"01",X"54",X"3D",X"33",X"75",X"80",X"8D",X"D0",X"05",X"7E",
		X"01",X"33",X"74",X"80",X"6B",X"01",X"23",X"44",X"80",X"97",X"94",X"00",X"41",X"70",X"62",X"80",
		X"10",X"00",X"13",X"4C",X"10",X"C2",X"05",X"02",X"0C",X"1A",X"0B",X"D3",X"10",X"FC",X"61",X"06",
		X"72",X"42",X"14",X"30",X"F4",X"C8",X"2B",X"72",X"80",X"D3",X"05",X"72",X"23",X"72",X"80",X"C8",
		X"C7",X"FB",X"07",X"02",X"01",X"08",X"07",X"42",X"FB",X"0E",X"0C",X"0C",X"FA",X"07",X"C7",X"F3",
		X"41",X"7E",X"01",X"33",X"80",X"80",X"8D",X"25",X"05",X"3B",X"75",X"80",X"E7",X"30",X"19",X"DD",
		X"F4",X"07",X"8D",X"9C",X"05",X"DD",X"37",X"0E",X"6B",X"FF",X"8D",X"B8",X"02",X"7E",X"FF",X"DD",
		X"B8",X"02",X"EE",X"33",X"80",X"80",X"0D",X"51",X"8D",X"37",X"0E",X"3B",X"72",X"80",X"FF",X"01",
		X"61",X"08",X"8D",X"30",X"0A",X"DD",X"F8",X"09",X"0D",X"06",X"8D",X"6B",X"0A",X"DD",X"F8",X"09",
		X"41",X"3B",X"00",X"B8",X"F6",X"08",X"FF",X"08",X"69",X"0B",X"2B",X"00",X"B8",X"F3",X"04",X"AE",
		X"04",X"38",X"19",X"09",X"D6",X"3B",X"72",X"80",X"FF",X"02",X"2D",X"CF",X"6B",X"01",X"23",X"80",
		X"80",X"3B",X"72",X"80",X"D6",X"98",X"32",X"33",X"72",X"80",X"0D",X"0D",X"EE",X"33",X"80",X"80",
		X"2B",X"72",X"80",X"D3",X"99",X"72",X"23",X"72",X"80",X"DD",X"62",X"05",X"8D",X"36",X"07",X"EF",
		X"8D",X"F7",X"06",X"7E",X"01",X"DD",X"F7",X"06",X"2B",X"FC",X"80",X"33",X"82",X"80",X"9D",X"10",
		X"EE",X"33",X"73",X"80",X"8D",X"25",X"05",X"3B",X"D8",X"80",X"7D",X"33",X"D8",X"80",X"2B",X"81",
		X"80",X"DD",X"F7",X"06",X"2B",X"D8",X"80",X"B2",X"69",X"43",X"2B",X"80",X"80",X"B2",X"69",X"2C",
		X"2B",X"82",X"80",X"B2",X"69",X"26",X"2B",X"81",X"80",X"68",X"F6",X"01",X"23",X"81",X"80",X"3B",
		X"7C",X"80",X"E7",X"30",X"17",X"3B",X"81",X"80",X"E7",X"38",X"0A",X"7E",X"01",X"33",X"01",X"A0",
		X"23",X"02",X"A0",X"09",X"07",X"EF",X"23",X"01",X"A0",X"33",X"02",X"A0",X"8D",X"62",X"05",X"3B",
		X"81",X"80",X"8D",X"0D",X"07",X"7E",X"01",X"33",X"44",X"80",X"C2",X"94",X"00",X"3B",X"75",X"80",
		X"E7",X"9B",X"72",X"00",X"8D",X"A9",X"0A",X"DD",X"18",X"0B",X"2B",X"80",X"80",X"B2",X"69",X"06",
		X"2B",X"82",X"80",X"B2",X"61",X"B0",X"8D",X"F2",X"0A",X"EF",X"23",X"73",X"80",X"33",X"74",X"80",
		X"23",X"75",X"80",X"33",X"81",X"80",X"23",X"80",X"80",X"33",X"01",X"A0",X"23",X"02",X"A0",X"7E",
		X"01",X"33",X"44",X"80",X"C2",X"72",X"00",X"10",X"E7",X"30",X"05",X"44",X"EA",X"80",X"0D",X"03",
		X"10",X"FC",X"80",X"70",X"D8",X"80",X"54",X"12",X"00",X"DD",X"4A",X"04",X"9D",X"10",X"E7",X"30",
		X"0B",X"3B",X"FC",X"80",X"23",X"82",X"80",X"70",X"EA",X"80",X"0D",X"09",X"2B",X"EA",X"80",X"33",
		X"82",X"80",X"74",X"FC",X"80",X"44",X"D8",X"80",X"54",X"12",X"00",X"DD",X"4A",X"04",X"EE",X"33",
		X"20",X"81",X"23",X"21",X"81",X"C8",X"41",X"3B",X"7E",X"80",X"23",X"D8",X"80",X"EF",X"23",X"D9",
		X"80",X"33",X"DA",X"80",X"23",X"DB",X"80",X"7E",X"00",X"33",X"DC",X"80",X"23",X"DD",X"80",X"EF",
		X"23",X"DE",X"80",X"33",X"20",X"81",X"23",X"21",X"81",X"33",X"DF",X"80",X"23",X"E8",X"80",X"33",
		X"E9",X"80",X"9D",X"10",X"10",X"CD",X"07",X"DD",X"72",X"04",X"10",X"D7",X"07",X"DD",X"72",X"04",
		X"10",X"DF",X"07",X"DD",X"72",X"04",X"10",X"E8",X"07",X"DD",X"72",X"04",X"10",X"A7",X"07",X"DD",
		X"C5",X"04",X"10",X"AD",X"07",X"DD",X"C5",X"04",X"10",X"B3",X"07",X"DD",X"C5",X"04",X"2B",X"80",
		X"80",X"B2",X"D4",X"3B",X"75",X"80",X"E7",X"9D",X"10",X"B9",X"07",X"DD",X"72",X"04",X"10",X"C3",
		X"07",X"DD",X"72",X"04",X"9D",X"C7",X"FB",X"FF",X"09",X"02",X"EB",X"80",X"06",X"FF",X"05",X"02",
		X"83",X"80",X"06",X"FF",X"0D",X"02",X"FD",X"80",X"06",X"FF",X"0C",X"02",X"52",X"52",X"52",X"52",
		X"52",X"52",X"FF",X"FF",X"0D",X"02",X"52",X"52",X"52",X"52",X"52",X"52",X"FF",X"FF",X"08",X"02",
		X"1C",X"0C",X"18",X"1B",X"0E",X"01",X"FF",X"FF",X"03",X"02",X"11",X"12",X"10",X"11",X"FF",X"FF",
		X"04",X"02",X"1C",X"0C",X"18",X"1B",X"0E",X"FF",X"FF",X"0C",X"02",X"1C",X"0C",X"18",X"1B",X"0E",
		X"02",X"FF",X"C7",X"F3",X"41",X"DD",X"63",X"04",X"74",X"00",X"98",X"02",X"20",X"76",X"80",X"77",
		X"14",X"30",X"FA",X"97",X"00",X"10",X"41",X"02",X"08",X"6D",X"FF",X"01",X"69",X"1A",X"FF",X"07",
		X"61",X"0D",X"C9",X"4B",X"00",X"CD",X"53",X"01",X"8D",X"72",X"04",X"CD",X"72",X"CD",X"72",X"CD",
		X"5B",X"00",X"C9",X"43",X"01",X"DD",X"72",X"04",X"1F",X"10",X"C2",X"10",X"10",X"56",X"20",X"37",
		X"72",X"04",X"61",X"FB",X"8D",X"48",X"09",X"7E",X"08",X"DD",X"B8",X"02",X"1C",X"30",X"EB",X"CD",
		X"72",X"CD",X"72",X"55",X"61",X"C3",X"6B",X"FF",X"8D",X"B8",X"02",X"7E",X"FF",X"DD",X"B8",X"02",
		X"6B",X"FF",X"8D",X"B8",X"02",X"C8",X"C7",X"FB",X"68",X"08",X"7C",X"08",X"99",X"08",X"B6",X"08",
		X"CE",X"08",X"EE",X"08",X"0F",X"09",X"2D",X"09",X"0B",X"0E",X"02",X"0C",X"18",X"19",X"22",X"1B",
		X"12",X"10",X"11",X"1D",X"52",X"52",X"52",X"01",X"09",X"08",X"00",X"FF",X"1E",X"10",X"02",X"C0",
		X"C1",X"C4",X"C5",X"C8",X"C9",X"CC",X"CD",X"D0",X"D1",X"D4",X"D5",X"D8",X"D9",X"DC",X"DD",X"4F",
		X"E0",X"E1",X"E4",X"E5",X"E8",X"E9",X"EC",X"ED",X"FF",X"1E",X"11",X"02",X"C2",X"C3",X"C6",X"C7",
		X"CA",X"CB",X"CE",X"CF",X"D2",X"D3",X"D6",X"D7",X"DA",X"DB",X"DE",X"DF",X"4F",X"E2",X"E3",X"E6",
		X"E7",X"EA",X"EB",X"EE",X"EF",X"FF",X"0A",X"13",X"02",X"0A",X"15",X"15",X"52",X"1B",X"12",X"10",
		X"11",X"1D",X"1C",X"52",X"1B",X"0E",X"1C",X"0E",X"1B",X"1F",X"0E",X"0D",X"2C",X"FF",X"0A",X"15",
		X"02",X"17",X"18",X"52",X"19",X"0A",X"1B",X"1D",X"52",X"18",X"0F",X"52",X"1D",X"11",X"12",X"1C",
		X"52",X"1C",X"18",X"0F",X"1D",X"20",X"0A",X"1B",X"0E",X"52",X"16",X"0A",X"22",X"FF",X"0A",X"17",
		X"02",X"0B",X"0E",X"52",X"0C",X"18",X"19",X"12",X"0E",X"0D",X"52",X"18",X"1B",X"52",X"1E",X"1C",
		X"0E",X"0D",X"52",X"20",X"12",X"1D",X"11",X"18",X"1E",X"1D",X"52",X"1D",X"11",X"0E",X"FF",X"0A",
		X"19",X"02",X"0E",X"21",X"19",X"1B",X"0E",X"1C",X"1C",X"52",X"20",X"1B",X"12",X"1D",X"1D",X"0E",
		X"17",X"52",X"0C",X"18",X"17",X"1C",X"0E",X"17",X"1D",X"52",X"18",X"0F",X"FF",X"0A",X"1B",X"02",
		X"17",X"12",X"11",X"18",X"17",X"52",X"0B",X"1E",X"1C",X"1C",X"0A",X"17",X"52",X"0C",X"18",X"2F",
		X"52",X"15",X"1D",X"0D",X"2C",X"FF",X"C7",X"F3",X"E9",X"F5",X"A5",X"C5",X"85",X"ED",X"74",X"DC",
		X"98",X"3B",X"AF",X"82",X"E6",X"30",X"4D",X"3B",X"B1",X"82",X"E6",X"30",X"2F",X"ED",X"63",X"01",
		X"03",X"ED",X"63",X"02",X"F0",X"ED",X"63",X"03",X"40",X"ED",X"63",X"00",X"04",X"70",X"C4",X"09",
		X"10",X"F3",X"88",X"50",X"0A",X"00",X"8D",X"4A",X"04",X"50",X"E6",X"FF",X"EA",X"58",X"EA",X"ED",
		X"75",X"00",X"61",X"EF",X"6B",X"01",X"23",X"B1",X"82",X"97",X"BC",X"09",X"E9",X"6B",X"02",X"AE",
		X"E0",X"21",X"11",X"70",X"EC",X"09",X"10",X"B3",X"88",X"50",X"0A",X"00",X"8D",X"4A",X"04",X"7E",
		X"01",X"33",X"AF",X"82",X"FF",X"02",X"69",X"11",X"E9",X"24",X"02",X"ED",X"7B",X"02",X"FF",X"91",
		X"25",X"0A",X"6B",X"02",X"23",X"AF",X"82",X"09",X"03",X"ED",X"21",X"02",X"95",X"90",X"B5",X"ED",
		X"B5",X"C8",X"C7",X"FB",X"94",X"95",X"B4",X"B5",X"D4",X"D5",X"F4",X"F5",X"F5",X"CB",X"92",X"93",
		X"B2",X"B3",X"D2",X"D3",X"F2",X"F3",X"EA",X"EB",X"90",X"91",X"B0",X"B1",X"D0",X"D1",X"F0",X"F1",
		X"E8",X"E9",X"8E",X"8F",X"AE",X"AF",X"CE",X"CF",X"EE",X"EF",X"CA",X"C9",X"8C",X"8D",X"AC",X"AD",
		X"CC",X"CD",X"EC",X"ED",X"C8",X"C9",X"C7",X"F3",X"41",X"3B",X"7A",X"80",X"FF",X"04",X"69",X"0D",
		X"10",X"1E",X"0A",X"DD",X"72",X"04",X"10",X"28",X"0A",X"DD",X"C5",X"04",X"9D",X"44",X"16",X"0A",
		X"8D",X"72",X"04",X"C8",X"C7",X"FB",X"0A",X"1C",X"01",X"0F",X"1B",X"0E",X"0E",X"FF",X"0A",X"1C",
		X"01",X"0C",X"1B",X"0E",X"0D",X"12",X"1D",X"FF",X"0A",X"1D",X"04",X"72",X"80",X"02",X"C7",X"F3",
		X"41",X"44",X"46",X"0A",X"8D",X"72",X"04",X"44",X"4E",X"0A",X"8D",X"72",X"04",X"44",X"61",X"0A",
		X"8D",X"72",X"04",X"C8",X"C7",X"FB",X"0B",X"10",X"0C",X"19",X"1E",X"1C",X"11",X"FF",X"0B",X"12",
		X"07",X"01",X"52",X"19",X"15",X"0A",X"22",X"0E",X"1B",X"52",X"0B",X"1E",X"1D",X"1D",X"18",X"17",
		X"FF",X"0B",X"14",X"0C",X"18",X"17",X"15",X"22",X"FF",X"C7",X"F3",X"10",X"10",X"81",X"0A",X"DD",
		X"72",X"04",X"10",X"89",X"0A",X"DD",X"72",X"04",X"10",X"9D",X"0A",X"DD",X"72",X"04",X"9D",X"C7",
		X"FB",X"0B",X"10",X"0C",X"19",X"1E",X"1C",X"11",X"FF",X"0B",X"12",X"07",X"01",X"52",X"18",X"1B",
		X"52",X"02",X"52",X"19",X"15",X"0A",X"22",X"0E",X"1B",X"1C",X"52",X"52",X"FF",X"0B",X"14",X"0B",
		X"0B",X"1E",X"1D",X"1D",X"18",X"17",X"FF",X"C7",X"F3",X"10",X"8D",X"63",X"04",X"3B",X"81",X"80",
		X"E7",X"30",X"05",X"44",X"CE",X"0A",X"0D",X"03",X"10",X"DF",X"0A",X"DD",X"72",X"04",X"8D",X"63",
		X"07",X"7E",X"FF",X"DD",X"B8",X"02",X"6B",X"FF",X"8D",X"B8",X"02",X"C8",X"C7",X"FB",X"0B",X"0D",
		X"0A",X"19",X"15",X"0A",X"22",X"0E",X"1B",X"52",X"01",X"52",X"18",X"1F",X"0E",X"1B",X"FF",X"0B",
		X"0D",X"0A",X"19",X"15",X"0A",X"22",X"0E",X"1B",X"52",X"02",X"52",X"18",X"1F",X"0E",X"1B",X"FF",
		X"C7",X"F3",X"41",X"44",X"09",X"0B",X"8D",X"72",X"04",X"DD",X"63",X"07",X"6B",X"FF",X"8D",X"B8",
		X"02",X"7E",X"FF",X"DD",X"B8",X"02",X"9D",X"C7",X"FB",X"0B",X"11",X"0C",X"10",X"0A",X"16",X"0E",
		X"52",X"18",X"1F",X"0E",X"1B",X"FF",X"C7",X"F3",X"41",X"CD",X"74",X"D9",X"80",X"ED",X"74",X"83",
		X"80",X"22",X"05",X"2A",X"00",X"CD",X"7B",X"00",X"E9",X"D7",X"00",X"29",X"18",X"30",X"21",X"CD",
		X"7B",X"01",X"E9",X"D7",X"01",X"29",X"0E",X"30",X"17",X"CD",X"7B",X"02",X"E9",X"D7",X"02",X"29",
		X"04",X"38",X"02",X"09",X"0B",X"ED",X"72",X"ED",X"72",X"ED",X"72",X"7C",X"34",X"30",X"D6",X"C8",
		X"6D",X"33",X"1F",X"81",X"8D",X"79",X"0B",X"C8",X"41",X"E5",X"85",X"C5",X"A5",X"70",X"00",X"90",
		X"12",X"52",X"12",X"F3",X"F8",X"1F",X"43",X"00",X"18",X"4C",X"18",X"4C",X"17",X"20",X"63",X"52",
		X"72",X"55",X"61",X"FA",X"B5",X"90",X"95",X"B0",X"9D",X"10",X"8D",X"37",X"0E",X"DD",X"6A",X"0F",
		X"6B",X"59",X"23",X"B2",X"82",X"7E",X"10",X"33",X"B3",X"82",X"10",X"18",X"0E",X"DD",X"72",X"04",
		X"10",X"24",X"0E",X"DD",X"72",X"04",X"10",X"29",X"0E",X"DD",X"C5",X"04",X"10",X"2F",X"0E",X"DD",
		X"C5",X"04",X"EE",X"33",X"1C",X"81",X"EE",X"33",X"1D",X"81",X"C2",X"EF",X"0B",X"97",X"20",X"00",
		X"E7",X"30",X"05",X"3B",X"00",X"A0",X"0D",X"03",X"2B",X"00",X"A8",X"33",X"54",X"81",X"F6",X"04",
		X"61",X"12",X"2B",X"54",X"81",X"F3",X"08",X"30",X"18",X"3B",X"54",X"81",X"F6",X"F0",X"93",X"65",
		X"0C",X"97",X"DA",X"0C",X"2B",X"1C",X"81",X"B2",X"9B",X"DA",X"0C",X"2C",X"23",X"1C",X"81",X"09",
		X"0E",X"3B",X"1C",X"81",X"FF",X"1C",X"9B",X"DA",X"0C",X"68",X"23",X"1C",X"81",X"09",X"00",X"CD",
		X"74",X"80",X"98",X"70",X"29",X"0C",X"2B",X"1C",X"81",X"52",X"F6",X"FE",X"5E",X"56",X"00",X"4C",
		X"7B",X"02",X"12",X"C1",X"C9",X"37",X"03",X"77",X"07",X"7E",X"F2",X"C1",X"C9",X"37",X"02",X"CD",
		X"63",X"00",X"0E",X"CD",X"63",X"01",X"02",X"3B",X"81",X"80",X"E7",X"9B",X"C9",X"0B",X"C9",X"24",
		X"02",X"CD",X"75",X"02",X"C2",X"C9",X"0B",X"C7",X"FB",X"35",X"9C",X"45",X"9C",X"55",X"9C",X"65",
		X"9C",X"75",X"9C",X"85",X"9C",X"95",X"9C",X"A5",X"9C",X"B5",X"9C",X"35",X"AC",X"45",X"AC",X"55",
		X"AC",X"65",X"AC",X"75",X"AC",X"85",X"AC",X"95",X"AC",X"A5",X"AC",X"B5",X"AC",X"C9",X"AC",X"35",
		X"BC",X"45",X"BC",X"55",X"BC",X"65",X"BC",X"75",X"BC",X"85",X"BC",X"95",X"BC",X"A5",X"BC",X"B5",
		X"BC",X"C7",X"BC",X"C7",X"F3",X"3B",X"1C",X"81",X"FF",X"1C",X"9B",X"1A",X"0D",X"AE",X"12",X"38",
		X"30",X"AE",X"12",X"29",X"08",X"AE",X"1B",X"38",X"08",X"D3",X"09",X"09",X"06",X"D3",X"0A",X"09",
		X"02",X"7E",X"2C",X"33",X"1E",X"81",X"2B",X"1D",X"81",X"AE",X"03",X"21",X"4D",X"70",X"11",X"81",
		X"5E",X"56",X"00",X"4C",X"2B",X"1E",X"81",X"37",X"2B",X"1D",X"81",X"68",X"23",X"1D",X"81",X"09",
		X"1A",X"7E",X"52",X"33",X"1E",X"81",X"2B",X"1D",X"81",X"B2",X"69",X"2E",X"7D",X"33",X"1D",X"81",
		X"74",X"11",X"81",X"1F",X"43",X"00",X"18",X"3B",X"1E",X"81",X"76",X"CD",X"74",X"0E",X"81",X"CD",
		X"63",X"00",X"0B",X"CD",X"63",X"01",X"12",X"CD",X"63",X"02",X"0B",X"CD",X"63",X"0D",X"FF",X"44",
		X"0E",X"81",X"8D",X"72",X"04",X"7E",X"50",X"DD",X"B8",X"02",X"6B",X"30",X"8D",X"B8",X"02",X"70",
		X"B3",X"82",X"7B",X"86",X"01",X"72",X"76",X"30",X"08",X"76",X"10",X"7F",X"7B",X"86",X"01",X"72",
		X"76",X"70",X"B2",X"82",X"7B",X"AE",X"00",X"30",X"12",X"77",X"7B",X"AE",X"01",X"30",X"0C",X"EF",
		X"23",X"B3",X"82",X"44",X"2F",X"0E",X"8D",X"C5",X"04",X"09",X"0F",X"44",X"29",X"0E",X"8D",X"C5",
		X"04",X"44",X"2F",X"0E",X"8D",X"C5",X"04",X"97",X"AD",X"0B",X"2B",X"1F",X"81",X"06",X"6B",X"04",
		X"D1",X"06",X"E7",X"9B",X"70",X"0D",X"C9",X"70",X"8C",X"80",X"E9",X"70",X"8F",X"80",X"10",X"FA",
		X"FF",X"0A",X"03",X"CD",X"7B",X"00",X"E9",X"37",X"00",X"CD",X"72",X"ED",X"72",X"5D",X"61",X"F3",
		X"C9",X"4C",X"E9",X"4C",X"14",X"30",X"EA",X"3B",X"1F",X"81",X"02",X"7E",X"04",X"C1",X"02",X"CD",
		X"74",X"BF",X"80",X"ED",X"74",X"CD",X"80",X"0A",X"0A",X"CD",X"7B",X"00",X"E9",X"37",X"00",X"CD",
		X"72",X"ED",X"72",X"5D",X"61",X"F3",X"10",X"E8",X"FF",X"CD",X"18",X"ED",X"18",X"55",X"61",X"E7",
		X"2B",X"1F",X"81",X"06",X"0A",X"ED",X"74",X"83",X"80",X"B2",X"69",X"09",X"E9",X"77",X"E9",X"77",
		X"E9",X"77",X"14",X"30",X"F7",X"CD",X"74",X"D9",X"80",X"02",X"03",X"CD",X"7B",X"00",X"E9",X"37",
		X"00",X"CD",X"72",X"ED",X"72",X"55",X"61",X"F3",X"E9",X"70",X"95",X"80",X"68",X"B2",X"69",X"08",
		X"10",X"0E",X"00",X"ED",X"18",X"5D",X"61",X"FB",X"74",X"0E",X"0E",X"CD",X"74",X"11",X"81",X"02",
		X"0A",X"1A",X"C9",X"6B",X"00",X"FC",X"61",X"1F",X"72",X"CD",X"72",X"55",X"61",X"F3",X"2B",X"72",
		X"80",X"D3",X"02",X"72",X"23",X"72",X"80",X"CD",X"63",X"FF",X"52",X"CD",X"63",X"FE",X"52",X"CD",
		X"63",X"FD",X"52",X"CD",X"63",X"FC",X"52",X"CD",X"74",X"11",X"81",X"0A",X"0A",X"CD",X"7B",X"00",
		X"E9",X"37",X"00",X"CD",X"72",X"ED",X"72",X"5D",X"61",X"F3",X"8D",X"37",X"0E",X"EF",X"23",X"82",
		X"98",X"7E",X"FF",X"DD",X"B8",X"02",X"6B",X"FF",X"8D",X"B8",X"02",X"7E",X"FF",X"DD",X"B8",X"02",
		X"17",X"1C",X"6B",X"02",X"8D",X"58",X"0B",X"68",X"14",X"30",X"F9",X"C8",X"C7",X"FB",X"13",X"18",
		X"1B",X"0D",X"0A",X"17",X"2C",X"15",X"1D",X"0D",X"0A",X"1A",X"07",X"1B",X"0E",X"10",X"52",X"1D",
		X"12",X"16",X"0E",X"FF",X"0A",X"1C",X"0C",X"2D",X"FF",X"0A",X"1C",X"0A",X"B2",X"82",X"02",X"0A",
		X"1C",X"0D",X"B3",X"82",X"01",X"C7",X"F3",X"10",X"8D",X"47",X"05",X"DD",X"63",X"04",X"6B",X"02",
		X"17",X"34",X"8D",X"58",X"0B",X"68",X"14",X"30",X"F9",X"44",X"10",X"0F",X"8D",X"72",X"04",X"44",
		X"22",X"0F",X"8D",X"72",X"04",X"44",X"4A",X"0F",X"8D",X"C5",X"04",X"CD",X"74",X"92",X"80",X"CD",
		X"63",X"00",X"0A",X"CD",X"63",X"01",X"05",X"CD",X"63",X"02",X"11",X"CD",X"63",X"0D",X"FF",X"44",
		X"92",X"80",X"8D",X"72",X"04",X"44",X"2A",X"0F",X"8D",X"72",X"04",X"44",X"50",X"0F",X"8D",X"C5",
		X"04",X"CD",X"74",X"A0",X"80",X"CD",X"63",X"00",X"0A",X"CD",X"63",X"01",X"07",X"CD",X"63",X"02",
		X"11",X"CD",X"63",X"0D",X"FF",X"44",X"A0",X"80",X"8D",X"72",X"04",X"44",X"32",X"0F",X"8D",X"72",
		X"04",X"44",X"56",X"0F",X"8D",X"C5",X"04",X"CD",X"74",X"AE",X"80",X"CD",X"63",X"00",X"0A",X"CD",
		X"63",X"01",X"09",X"CD",X"63",X"02",X"11",X"CD",X"63",X"0D",X"FF",X"44",X"AE",X"80",X"8D",X"72",
		X"04",X"44",X"3A",X"0F",X"8D",X"72",X"04",X"44",X"5C",X"0F",X"8D",X"C5",X"04",X"CD",X"74",X"BC",
		X"80",X"CD",X"63",X"00",X"0A",X"CD",X"63",X"01",X"0B",X"CD",X"63",X"02",X"11",X"CD",X"63",X"0D",
		X"FF",X"44",X"BC",X"80",X"8D",X"72",X"04",X"44",X"42",X"0F",X"8D",X"72",X"04",X"44",X"62",X"0F",
		X"8D",X"C5",X"04",X"CD",X"74",X"CA",X"80",X"CD",X"63",X"00",X"0A",X"CD",X"63",X"01",X"0D",X"CD",
		X"63",X"02",X"11",X"CD",X"63",X"0D",X"FF",X"44",X"CA",X"80",X"8D",X"72",X"04",X"C8",X"C7",X"FB",
		X"0A",X"03",X"0A",X"1C",X"0C",X"18",X"1B",X"0E",X"52",X"52",X"52",X"52",X"52",X"17",X"0A",X"16",
		X"0E",X"FF",X"0A",X"05",X"04",X"17",X"18",X"01",X"2D",X"FF",X"0A",X"07",X"04",X"17",X"18",X"02",
		X"2D",X"FF",X"0A",X"09",X"04",X"17",X"18",X"03",X"2D",X"FF",X"0A",X"0B",X"04",X"17",X"18",X"04",
		X"2D",X"FF",X"0A",X"0D",X"04",X"17",X"18",X"05",X"2D",X"FF",X"0A",X"05",X"09",X"83",X"80",X"06",
		X"0A",X"07",X"09",X"86",X"80",X"06",X"0A",X"09",X"09",X"89",X"80",X"06",X"0A",X"0B",X"09",X"8C",
		X"80",X"06",X"0A",X"0D",X"09",X"8F",X"80",X"06",X"C7",X"F3",X"41",X"44",X"98",X"0F",X"8D",X"72",
		X"04",X"44",X"AD",X"0F",X"8D",X"72",X"04",X"44",X"B6",X"0F",X"8D",X"72",X"04",X"44",X"CC",X"0F",
		X"8D",X"72",X"04",X"44",X"E4",X"0F",X"8D",X"72",X"04",X"70",X"11",X"81",X"17",X"0A",X"63",X"52",
		X"72",X"55",X"93",X"8E",X"0F",X"C8",X"C7",X"FB",X"0A",X"10",X"06",X"17",X"0A",X"16",X"0E",X"52",
		X"1B",X"0E",X"10",X"12",X"1C",X"1D",X"1B",X"0A",X"1D",X"12",X"18",X"17",X"FF",X"0A",X"12",X"05",
		X"17",X"0A",X"16",X"0E",X"2D",X"FF",X"0A",X"14",X"05",X"0A",X"52",X"0B",X"52",X"0C",X"52",X"0D",
		X"52",X"0E",X"52",X"0F",X"52",X"10",X"52",X"11",X"52",X"12",X"52",X"FF",X"0A",X"16",X"05",X"13",
		X"52",X"14",X"52",X"15",X"52",X"16",X"52",X"17",X"52",X"18",X"52",X"19",X"52",X"1A",X"52",X"1B",
		X"52",X"3C",X"3D",X"FF",X"0A",X"18",X"05",X"1C",X"52",X"1D",X"52",X"1E",X"52",X"1F",X"52",X"20",
		X"52",X"21",X"52",X"22",X"52",X"23",X"52",X"2C",X"52",X"3E",X"3F",X"FF",X"C7",X"F3",X"41",X"10",
		X"C9",X"70",X"58",X"08",X"6B",X"80",X"23",X"31",X"81",X"97",X"07",X"08",X"41",X"10",X"41",X"10",
		X"74",X"00",X"98",X"3B",X"31",X"81",X"29",X"33",X"31",X"81",X"C2",X"2D",X"08",X"10",X"41",X"10",
		X"41",X"DD",X"27",X"10",X"8D",X"0F",X"03",X"CD",X"74",X"5C",X"81",X"44",X"08",X"00",X"37",X"04",
		X"C9",X"6B",X"00",X"AE",X"00",X"38",X"07",X"CD",X"7B",X"03",X"FF",X"07",X"25",X"0D",X"3F",X"08",
		X"C9",X"76",X"00",X"00",X"C9",X"77",X"3C",X"30",X"F7",X"09",X"02",X"CD",X"18",X"75",X"61",X"E0",
		X"C9",X"70",X"5C",X"81",X"E9",X"70",X"80",X"98",X"10",X"08",X"00",X"50",X"04",X"00",X"37",X"04",
		X"C9",X"6B",X"00",X"AE",X"F0",X"38",X"19",X"2A",X"04",X"CD",X"72",X"CD",X"7B",X"00",X"E9",X"37",
		X"00",X"CD",X"72",X"ED",X"72",X"7D",X"61",X"F3",X"C9",X"77",X"C9",X"77",X"C9",X"77",X"0D",X"04",
		X"C9",X"4C",X"E9",X"58",X"34",X"30",X"D9",X"CD",X"74",X"5C",X"81",X"ED",X"74",X"83",X"82",X"02",
		X"04",X"CD",X"7B",X"00",X"E6",X"30",X"14",X"ED",X"7B",X"06",X"FF",X"01",X"69",X"0D",X"1F",X"08",
		X"EE",X"ED",X"76",X"00",X"E9",X"77",X"1C",X"30",X"F8",X"09",X"02",X"ED",X"18",X"CD",X"18",X"55",
		X"61",X"DF",X"9D",X"7E",X"01",X"33",X"44",X"80",X"7F",X"00",X"80",X"6B",X"FF",X"FF",X"61",X"F8",
		X"2B",X"DF",X"80",X"D3",X"01",X"F3",X"03",X"33",X"DF",X"80",X"8D",X"62",X"05",X"EF",X"23",X"DC",
		X"80",X"33",X"DD",X"80",X"74",X"00",X"00",X"27",X"E8",X"80",X"6B",X"01",X"8D",X"65",X"03",X"7E",
		X"FF",X"DD",X"B8",X"02",X"6B",X"00",X"23",X"44",X"80",X"C8",X"6B",X"01",X"23",X"44",X"80",X"7E",
		X"FF",X"DD",X"B8",X"02",X"8D",X"62",X"05",X"EF",X"23",X"DC",X"80",X"33",X"DD",X"80",X"6B",X"01",
		X"23",X"73",X"80",X"7E",X"80",X"DD",X"B8",X"02",X"9D",X"3B",X"E6",X"80",X"0A",X"3B",X"E5",X"80",
		X"02",X"3B",X"E4",X"80",X"F1",X"F4",X"DC",X"3B",X"E3",X"80",X"0A",X"3B",X"E2",X"80",X"02",X"D5",
		X"8D",X"A5",X"27",X"DD",X"DD",X"27",X"95",X"DD",X"5D",X"11",X"6B",X"01",X"9D",X"70",X"30",X"00",
		X"77",X"E5",X"80",X"EF",X"23",X"E4",X"80",X"44",X"5F",X"1F",X"8D",X"C5",X"04",X"C8",X"2B",X"E4",
		X"80",X"B2",X"61",X"0D",X"2B",X"E6",X"80",X"2E",X"2B",X"E5",X"80",X"26",X"10",X"F0",X"CF",X"4C",
		X"C4",X"3B",X"E3",X"80",X"0A",X"3B",X"E2",X"80",X"02",X"DD",X"5D",X"11",X"9D",X"3B",X"75",X"80",
		X"E6",X"9D",X"2B",X"E6",X"80",X"D4",X"32",X"33",X"E6",X"80",X"2B",X"E5",X"80",X"C9",X"32",X"33",
		X"E5",X"80",X"2B",X"E4",X"80",X"02",X"00",X"C9",X"32",X"33",X"E4",X"80",X"10",X"5F",X"1F",X"DD",
		X"C5",X"04",X"9D",X"3B",X"7C",X"80",X"E6",X"30",X"08",X"3B",X"81",X"80",X"E6",X"38",X"02",X"EF",
		X"9D",X"7E",X"01",X"C8",X"2B",X"DF",X"80",X"52",X"5E",X"56",X"00",X"70",X"A9",X"11",X"18",X"4B",
		X"72",X"43",X"EA",X"27",X"20",X"81",X"9D",X"C7",X"FB",X"00",X"20",X"00",X"28",X"00",X"30",X"00",
		X"38",X"00",X"40",X"00",X"48",X"00",X"50",X"00",X"58",X"C7",X"F3",X"3B",X"75",X"80",X"E6",X"9D",
		X"C9",X"F5",X"A5",X"6D",X"17",X"00",X"FF",X"04",X"69",X"7A",X"FF",X"03",X"69",X"5B",X"FF",X"02",
		X"69",X"2C",X"68",X"52",X"12",X"52",X"0A",X"CD",X"74",X"6E",X"13",X"CD",X"5C",X"CD",X"27",X"00",
		X"C9",X"3A",X"01",X"27",X"0C",X"80",X"C9",X"6B",X"02",X"33",X"0F",X"80",X"C9",X"32",X"04",X"CD",
		X"2F",X"05",X"77",X"18",X"80",X"CD",X"7B",X"06",X"23",X"1B",X"80",X"97",X"8C",X"12",X"68",X"52",
		X"12",X"52",X"0A",X"CD",X"74",X"92",X"12",X"CD",X"5C",X"CD",X"27",X"00",X"C9",X"3A",X"01",X"27",
		X"00",X"80",X"C9",X"6B",X"02",X"33",X"03",X"80",X"C9",X"32",X"04",X"CD",X"2F",X"05",X"77",X"0C",
		X"80",X"CD",X"7B",X"06",X"23",X"0F",X"80",X"09",X"63",X"3D",X"12",X"52",X"0A",X"CD",X"74",X"AA",
		X"12",X"CD",X"5C",X"CD",X"27",X"00",X"C9",X"3A",X"01",X"27",X"24",X"80",X"C9",X"6B",X"02",X"33",
		X"27",X"80",X"0D",X"48",X"68",X"52",X"12",X"52",X"12",X"0E",X"C9",X"70",X"CE",X"12",X"C9",X"58",
		X"C9",X"32",X"00",X"CD",X"2F",X"01",X"77",X"00",X"80",X"CD",X"7B",X"02",X"23",X"03",X"80",X"CD",
		X"27",X"04",X"C9",X"3A",X"05",X"27",X"0C",X"80",X"C9",X"6B",X"06",X"33",X"0F",X"80",X"C9",X"32",
		X"08",X"CD",X"2F",X"09",X"77",X"18",X"80",X"CD",X"7B",X"0A",X"23",X"1B",X"80",X"CD",X"27",X"0C",
		X"C9",X"3A",X"0D",X"27",X"24",X"80",X"C9",X"6B",X"0E",X"33",X"27",X"80",X"B5",X"CD",X"B5",X"C8",
		X"C7",X"FB",X"4B",X"10",X"81",X"00",X"4B",X"10",X"81",X"00",X"4D",X"20",X"90",X"00",X"4D",X"50",
		X"90",X"00",X"46",X"E0",X"82",X"00",X"46",X"E0",X"82",X"00",X"48",X"A0",X"81",X"00",X"48",X"C0",
		X"81",X"00",X"48",X"E0",X"81",X"00",X"4D",X"10",X"84",X"00",X"4A",X"20",X"81",X"00",X"4A",X"F4",
		X"81",X"00",X"4E",X"80",X"80",X"00",X"4E",X"90",X"80",X"00",X"00",X"00",X"00",X"00",X"48",X"00",
		X"82",X"00",X"48",X"40",X"82",X"00",X"48",X"60",X"82",X"00",X"48",X"80",X"82",X"00",X"4A",X"40",
		X"84",X"00",X"4A",X"80",X"84",X"00",X"4A",X"C0",X"84",X"00",X"4A",X"F4",X"84",X"00",X"4B",X"30",
		X"82",X"00",X"4B",X"80",X"82",X"00",X"4B",X"C0",X"82",X"00",X"4B",X"E0",X"82",X"00",X"4C",X"00",
		X"83",X"00",X"4C",X"38",X"83",X"00",X"4C",X"68",X"83",X"00",X"4C",X"90",X"83",X"00",X"4E",X"A0",
		X"87",X"00",X"4E",X"E8",X"87",X"00",X"4F",X"48",X"87",X"00",X"4F",X"A8",X"87",X"00",X"45",X"00",
		X"80",X"00",X"45",X"80",X"80",X"00",X"45",X"E0",X"80",X"00",X"46",X"10",X"80",X"00",X"49",X"00",
		X"86",X"00",X"49",X"50",X"86",X"00",X"49",X"A0",X"86",X"00",X"4A",X"00",X"86",X"00",X"4C",X"A0",
		X"84",X"00",X"4C",X"C0",X"84",X"00",X"4C",X"E0",X"84",X"00",X"4D",X"00",X"84",X"00",X"4D",X"70",
		X"82",X"00",X"4D",X"E0",X"82",X"00",X"4E",X"38",X"82",X"00",X"4F",X"A8",X"82",X"00",X"4F",X"B8",
		X"80",X"00",X"4F",X"C0",X"80",X"00",X"4F",X"C8",X"80",X"00",X"4F",X"D0",X"80",X"00",X"4F",X"E0",
		X"80",X"00",X"4F",X"F0",X"80",X"00",X"46",X"40",X"83",X"00",X"46",X"90",X"83",X"00",X"C7",X"F3",
		X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",
		X"41",X"3B",X"5B",X"81",X"FF",X"00",X"98",X"0F",X"03",X"AE",X"01",X"D9",X"25",X"14",X"FF",X"02",
		X"90",X"0F",X"03",X"3B",X"4C",X"81",X"FF",X"00",X"90",X"0F",X"03",X"DD",X"44",X"15",X"2B",X"81",
		X"82",X"AE",X"FF",X"38",X"18",X"DD",X"77",X"1A",X"2B",X"82",X"82",X"E7",X"61",X"09",X"8D",X"52",
		X"15",X"DD",X"2D",X"16",X"8D",X"0F",X"03",X"DD",X"2E",X"18",X"8D",X"0F",X"03",X"7E",X"FB",X"DD",
		X"D1",X"18",X"2B",X"75",X"80",X"E5",X"E6",X"33",X"75",X"80",X"8D",X"52",X"15",X"B0",X"23",X"75",
		X"80",X"DD",X"F0",X"18",X"2B",X"34",X"81",X"AE",X"F0",X"89",X"0F",X"03",X"FF",X"F8",X"80",X"0F",
		X"03",X"7E",X"FF",X"33",X"AB",X"82",X"74",X"90",X"98",X"02",X"10",X"76",X"00",X"77",X"14",X"30",
		X"FA",X"DD",X"EA",X"10",X"8D",X"0F",X"03",X"3B",X"3D",X"81",X"23",X"E7",X"80",X"3B",X"31",X"81",
		X"23",X"E8",X"80",X"3B",X"30",X"81",X"23",X"E9",X"80",X"7E",X"FF",X"33",X"81",X"82",X"54",X"07",
		X"04",X"DD",X"BB",X"11",X"9D",X"7E",X"02",X"DD",X"21",X"03",X"6B",X"03",X"8D",X"21",X"03",X"70",
		X"AD",X"14",X"10",X"32",X"81",X"50",X"10",X"00",X"8D",X"4A",X"04",X"70",X"BD",X"14",X"10",X"46",
		X"81",X"50",X"06",X"00",X"8D",X"4A",X"04",X"DD",X"44",X"15",X"6B",X"20",X"8D",X"B8",X"02",X"50",
		X"00",X"04",X"8D",X"BB",X"11",X"10",X"8D",X"44",X"15",X"DD",X"77",X"1A",X"2B",X"AA",X"82",X"9F",
		X"76",X"38",X"10",X"7E",X"02",X"33",X"5B",X"81",X"6B",X"02",X"8D",X"65",X"03",X"7E",X"03",X"DD",
		X"65",X"03",X"9D",X"10",X"2B",X"55",X"81",X"1F",X"43",X"00",X"29",X"F3",X"0F",X"33",X"55",X"81",
		X"74",X"C3",X"14",X"4C",X"7B",X"33",X"54",X"81",X"8D",X"BA",X"15",X"DD",X"2D",X"16",X"2B",X"4C",
		X"81",X"7A",X"D6",X"01",X"8D",X"D1",X"18",X"EF",X"23",X"4C",X"81",X"7E",X"0A",X"DD",X"B8",X"02",
		X"2B",X"AA",X"82",X"D3",X"01",X"33",X"AA",X"82",X"C2",X"55",X"14",X"C7",X"FB",X"7B",X"06",X"12",
		X"A8",X"3B",X"06",X"12",X"B8",X"79",X"06",X"22",X"A8",X"39",X"06",X"22",X"B8",X"01",X"01",X"04",
		X"01",X"04",X"00",X"22",X"22",X"22",X"22",X"80",X"10",X"10",X"10",X"10",X"40",X"04",X"01",X"01",
		X"01",X"01",X"08",X"C7",X"F3",X"10",X"74",X"AD",X"14",X"44",X"32",X"81",X"54",X"10",X"00",X"DD",
		X"4A",X"04",X"74",X"32",X"81",X"02",X"04",X"77",X"72",X"6B",X"D6",X"40",X"76",X"77",X"72",X"55",
		X"61",X"F5",X"2B",X"E7",X"80",X"86",X"40",X"5A",X"1A",X"5A",X"F6",X"1F",X"74",X"30",X"15",X"1F",
		X"43",X"00",X"18",X"12",X"6B",X"10",X"D0",X"0E",X"C9",X"70",X"32",X"81",X"C9",X"65",X"03",X"CD",
		X"60",X"07",X"C9",X"65",X"0B",X"CD",X"60",X"0F",X"74",X"BD",X"14",X"44",X"46",X"81",X"54",X"06",
		X"00",X"DD",X"4A",X"04",X"8D",X"44",X"15",X"50",X"00",X"04",X"8D",X"BB",X"11",X"C8",X"C7",X"FB",
		X"48",X"48",X"48",X"60",X"60",X"60",X"78",X"78",X"78",X"90",X"90",X"90",X"A8",X"A8",X"A8",X"C0",
		X"C0",X"C0",X"C7",X"F3",X"41",X"70",X"32",X"81",X"10",X"90",X"98",X"50",X"10",X"00",X"8D",X"4A",
		X"04",X"C8",X"41",X"3B",X"75",X"80",X"E7",X"38",X"1D",X"3B",X"7C",X"80",X"E7",X"30",X"06",X"3B",
		X"81",X"80",X"E7",X"30",X"08",X"3B",X"00",X"A0",X"23",X"54",X"81",X"09",X"4D",X"10",X"2B",X"00",
		X"A8",X"33",X"54",X"81",X"0D",X"44",X"2B",X"45",X"80",X"F3",X"1F",X"30",X"06",X"EF",X"23",X"54",
		X"81",X"09",X"14",X"3B",X"55",X"81",X"29",X"F3",X"3F",X"33",X"55",X"81",X"5E",X"56",X"00",X"70",
		X"E3",X"15",X"18",X"6B",X"23",X"54",X"81",X"3B",X"00",X"B8",X"CA",X"26",X"61",X"07",X"6B",X"01",
		X"23",X"B4",X"82",X"09",X"15",X"3B",X"B4",X"82",X"E6",X"38",X"0F",X"70",X"C0",X"4C",X"77",X"24",
		X"80",X"7E",X"84",X"33",X"27",X"80",X"EE",X"33",X"B4",X"82",X"41",X"56",X"00",X"0A",X"04",X"CD",
		X"74",X"45",X"81",X"3B",X"54",X"81",X"02",X"F3",X"03",X"1F",X"74",X"DF",X"15",X"4C",X"7B",X"CD",
		X"76",X"00",X"1C",X"38",X"07",X"CD",X"7A",X"6D",X"1A",X"5A",X"0D",X"EA",X"9D",X"C7",X"FB",X"00",
		X"01",X"FF",X"00",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"15",X"12",X"12",X"12",X"12",X"12",
		X"12",X"12",X"12",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"44",X"44",X"44",X"44",X"44",
		X"44",X"00",X"00",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"88",X"88",X"88",X"88",X"88",
		X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C7",X"F3",X"3B",X"46",X"81",
		X"02",X"3B",X"47",X"81",X"D0",X"38",X"27",X"06",X"2B",X"43",X"81",X"E7",X"61",X"06",X"2B",X"45",
		X"81",X"E7",X"69",X"04",X"41",X"DD",X"63",X"16",X"41",X"3B",X"42",X"81",X"E6",X"30",X"06",X"3B",
		X"44",X"81",X"E6",X"38",X"04",X"10",X"8D",X"54",X"17",X"10",X"8D",X"F0",X"18",X"C8",X"41",X"DD",
		X"07",X"14",X"9D",X"10",X"3D",X"AE",X"02",X"30",X"5C",X"3B",X"4A",X"81",X"0A",X"3B",X"48",X"81",
		X"BC",X"93",X"29",X"17",X"2B",X"45",X"81",X"06",X"2B",X"43",X"81",X"C4",X"69",X"03",X"B2",X"96",
		X"16",X"10",X"EE",X"33",X"46",X"81",X"23",X"47",X"81",X"10",X"2B",X"4A",X"81",X"AE",X"00",X"9D",
		X"6B",X"FC",X"23",X"4C",X"81",X"C8",X"41",X"AE",X"02",X"38",X"0E",X"3B",X"4A",X"81",X"FF",X"04",
		X"DC",X"EF",X"23",X"46",X"81",X"33",X"47",X"81",X"9D",X"10",X"2B",X"AC",X"82",X"AE",X"00",X"38",
		X"08",X"EF",X"23",X"43",X"81",X"33",X"45",X"81",X"9D",X"3B",X"4A",X"81",X"FF",X"04",X"DC",X"7E",
		X"04",X"33",X"4C",X"81",X"9D",X"10",X"2B",X"47",X"81",X"E7",X"69",X"2E",X"2B",X"45",X"81",X"AE",
		X"00",X"9D",X"B2",X"E1",X"16",X"3B",X"4A",X"81",X"FF",X"00",X"DC",X"7E",X"FC",X"33",X"4C",X"81",
		X"9D",X"10",X"2B",X"AC",X"82",X"AE",X"00",X"38",X"05",X"EF",X"23",X"45",X"81",X"C8",X"2B",X"4A",
		X"81",X"AE",X"04",X"9D",X"6B",X"04",X"23",X"4C",X"81",X"C8",X"41",X"3B",X"43",X"81",X"FF",X"00",
		X"DC",X"E6",X"10",X"17",X"2B",X"48",X"81",X"AE",X"00",X"9D",X"6B",X"FC",X"23",X"4C",X"81",X"C8",
		X"41",X"3B",X"AC",X"82",X"FF",X"00",X"69",X"05",X"EE",X"33",X"43",X"81",X"9D",X"3B",X"48",X"81",
		X"FF",X"04",X"DC",X"7E",X"04",X"33",X"4C",X"81",X"9D",X"10",X"2B",X"4A",X"81",X"AE",X"04",X"30",
		X"0C",X"EF",X"23",X"46",X"81",X"3B",X"45",X"81",X"FF",X"FF",X"D4",X"09",X"11",X"10",X"2B",X"48",
		X"81",X"AE",X"04",X"95",X"EE",X"33",X"47",X"81",X"2B",X"43",X"81",X"AE",X"FF",X"95",X"6B",X"FC",
		X"23",X"4C",X"81",X"C8",X"41",X"3B",X"44",X"81",X"02",X"3B",X"42",X"81",X"D0",X"38",X"05",X"E6",
		X"82",X"17",X"0D",X"15",X"2B",X"47",X"81",X"E7",X"69",X"08",X"EE",X"33",X"44",X"81",X"8D",X"DD",
		X"17",X"C8",X"23",X"42",X"81",X"DD",X"8B",X"17",X"9D",X"DD",X"DD",X"17",X"E6",X"95",X"8D",X"8B",
		X"17",X"C8",X"8D",X"8B",X"17",X"E7",X"D4",X"DD",X"DD",X"17",X"9D",X"3B",X"44",X"81",X"E6",X"38",
		X"4A",X"10",X"2B",X"46",X"81",X"E7",X"61",X"06",X"EE",X"33",X"44",X"81",X"0D",X"3D",X"2B",X"44",
		X"81",X"AE",X"01",X"30",X"1A",X"3B",X"4B",X"81",X"FF",X"00",X"69",X"2F",X"2B",X"49",X"81",X"AE",
		X"00",X"38",X"28",X"7E",X"F8",X"DD",X"B2",X"18",X"6B",X"FF",X"23",X"42",X"81",X"09",X"19",X"10",
		X"2B",X"4B",X"81",X"AE",X"01",X"38",X"14",X"3B",X"49",X"81",X"FF",X"01",X"69",X"0D",X"6B",X"08",
		X"8D",X"B2",X"18",X"7E",X"01",X"33",X"42",X"81",X"6B",X"FF",X"9D",X"EF",X"9D",X"3B",X"42",X"81",
		X"E6",X"38",X"49",X"3B",X"47",X"81",X"E6",X"30",X"06",X"EF",X"23",X"42",X"81",X"09",X"3D",X"3B",
		X"42",X"81",X"FF",X"01",X"61",X"1A",X"2B",X"49",X"81",X"AE",X"00",X"38",X"2F",X"3B",X"4B",X"81",
		X"FF",X"00",X"69",X"28",X"6B",X"F8",X"8D",X"B2",X"18",X"7E",X"FF",X"33",X"44",X"81",X"0D",X"19",
		X"41",X"3B",X"49",X"81",X"FF",X"01",X"69",X"14",X"2B",X"4B",X"81",X"AE",X"01",X"38",X"0D",X"7E",
		X"08",X"DD",X"B2",X"18",X"6B",X"01",X"23",X"44",X"81",X"7E",X"FF",X"C8",X"EE",X"C8",X"41",X"3B",
		X"46",X"81",X"02",X"3B",X"47",X"81",X"D0",X"AE",X"02",X"21",X"04",X"DD",X"07",X"14",X"9D",X"10",
		X"2B",X"82",X"82",X"F3",X"80",X"30",X"22",X"EF",X"23",X"46",X"81",X"3B",X"48",X"81",X"FF",X"00",
		X"61",X"0B",X"2B",X"4A",X"81",X"AE",X"04",X"30",X"04",X"7E",X"01",X"09",X"02",X"7E",X"FF",X"33",
		X"43",X"81",X"6B",X"01",X"23",X"45",X"81",X"09",X"21",X"EF",X"23",X"47",X"81",X"3B",X"4A",X"81",
		X"FF",X"00",X"61",X"0C",X"2B",X"48",X"81",X"AE",X"04",X"30",X"05",X"7E",X"01",X"97",X"82",X"18",
		X"6B",X"FF",X"23",X"45",X"81",X"7E",X"01",X"33",X"43",X"81",X"41",X"DD",X"2D",X"16",X"8D",X"44",
		X"15",X"3B",X"82",X"82",X"D6",X"FF",X"0A",X"F3",X"0F",X"38",X"0F",X"3D",X"23",X"82",X"82",X"7E",
		X"05",X"DD",X"B8",X"02",X"8D",X"77",X"1A",X"97",X"3F",X"18",X"8D",X"3E",X"11",X"EF",X"23",X"82",
		X"82",X"C8",X"41",X"06",X"2B",X"41",X"81",X"C4",X"23",X"41",X"81",X"3B",X"39",X"81",X"D0",X"33",
		X"39",X"81",X"2B",X"3D",X"81",X"C4",X"23",X"3D",X"81",X"3B",X"35",X"81",X"D0",X"33",X"35",X"81",
		X"9D",X"10",X"02",X"3B",X"40",X"81",X"D0",X"33",X"40",X"81",X"2B",X"38",X"81",X"C4",X"23",X"38",
		X"81",X"3B",X"3C",X"81",X"D0",X"33",X"3C",X"81",X"2B",X"34",X"81",X"C4",X"23",X"34",X"81",X"C8",
		X"2B",X"48",X"81",X"06",X"2B",X"43",X"81",X"C4",X"02",X"EE",X"2F",X"19",X"D7",X"05",X"B2",X"2F",
		X"19",X"6D",X"FF",X"01",X"61",X"11",X"2B",X"48",X"81",X"AE",X"00",X"30",X"1E",X"3B",X"40",X"81",
		X"D6",X"04",X"23",X"40",X"81",X"09",X"14",X"6D",X"FF",X"00",X"61",X"0F",X"2B",X"48",X"81",X"AE",
		X"01",X"30",X"08",X"3B",X"40",X"81",X"D7",X"04",X"23",X"40",X"81",X"6D",X"23",X"48",X"81",X"10",
		X"2B",X"49",X"81",X"06",X"2B",X"42",X"81",X"C4",X"02",X"EE",X"45",X"19",X"D7",X"02",X"B2",X"45",
		X"19",X"6D",X"23",X"49",X"81",X"3B",X"4A",X"81",X"02",X"3B",X"45",X"81",X"D0",X"06",X"BA",X"84",
		X"19",X"86",X"05",X"E6",X"84",X"19",X"3D",X"AE",X"01",X"30",X"11",X"3B",X"4A",X"81",X"FF",X"00",
		X"61",X"1E",X"2B",X"3C",X"81",X"D3",X"04",X"33",X"3C",X"81",X"0D",X"14",X"3D",X"AE",X"00",X"30",
		X"0F",X"3B",X"4A",X"81",X"FF",X"01",X"61",X"08",X"2B",X"3C",X"81",X"86",X"04",X"33",X"3C",X"81",
		X"3D",X"33",X"4A",X"81",X"2B",X"4B",X"81",X"06",X"2B",X"44",X"81",X"C4",X"02",X"EE",X"99",X"19",
		X"D7",X"02",X"B2",X"99",X"19",X"6D",X"23",X"4B",X"81",X"10",X"2B",X"48",X"81",X"52",X"12",X"0E",
		X"2B",X"49",X"81",X"52",X"91",X"0E",X"17",X"00",X"74",X"D3",X"19",X"58",X"7B",X"33",X"3E",X"81",
		X"72",X"6B",X"23",X"36",X"81",X"3B",X"4A",X"81",X"12",X"52",X"0A",X"3B",X"4B",X"81",X"12",X"91",
		X"0A",X"02",X"00",X"70",X"E7",X"19",X"5C",X"6B",X"23",X"3A",X"81",X"77",X"7B",X"33",X"32",X"81",
		X"9D",X"C7",X"FB",X"30",X"3A",X"35",X"3B",X"31",X"3C",X"36",X"3D",X"32",X"3E",X"37",X"3F",X"33",
		X"3E",X"38",X"3D",X"34",X"3C",X"39",X"3B",X"75",X"7B",X"70",X"7A",X"76",X"7D",X"71",X"7C",X"77",
		X"7F",X"72",X"7E",X"78",X"7D",X"73",X"7E",X"79",X"7B",X"74",X"7C",X"C7",X"F3",X"10",X"2B",X"31",
		X"81",X"C1",X"02",X"F3",X"0F",X"30",X"42",X"3B",X"22",X"81",X"CA",X"06",X"69",X"0A",X"3D",X"5A",
		X"1A",X"5A",X"1A",X"F3",X"0F",X"33",X"D9",X"82",X"3D",X"5A",X"F6",X"F8",X"02",X"3D",X"1A",X"5A",
		X"1A",X"F3",X"1F",X"70",X"55",X"1A",X"5E",X"56",X"00",X"4C",X"7B",X"1A",X"FF",X"FF",X"69",X"19",
		X"74",X"81",X"81",X"6D",X"5E",X"56",X"00",X"4C",X"48",X"4C",X"7B",X"AE",X"FF",X"38",X"0A",X"AE",
		X"05",X"EE",X"4C",X"1A",X"FF",X"0C",X"B2",X"4C",X"1A",X"7E",X"00",X"C8",X"68",X"33",X"DA",X"82",
		X"6B",X"01",X"9D",X"C7",X"FB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",
		X"01",X"FF",X"02",X"02",X"FF",X"03",X"03",X"FF",X"04",X"04",X"FF",X"05",X"05",X"FF",X"06",X"06",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"C7",X"F3",X"10",X"C9",X"70",X"98",X"98",X"C9",X"6B",X"00",X"F3",
		X"0F",X"52",X"F6",X"1E",X"E9",X"70",X"E9",X"1A",X"5E",X"56",X"00",X"ED",X"18",X"CD",X"7B",X"02",
		X"E9",X"C3",X"00",X"06",X"C9",X"6B",X"03",X"ED",X"83",X"01",X"0A",X"DD",X"FD",X"19",X"23",X"47",
		X"81",X"3B",X"22",X"81",X"D6",X"01",X"23",X"22",X"81",X"CD",X"74",X"9C",X"98",X"CD",X"7B",X"00",
		X"F6",X"0F",X"12",X"F3",X"1E",X"ED",X"74",X"D5",X"1A",X"1F",X"43",X"00",X"E9",X"4C",X"C9",X"6B",
		X"02",X"ED",X"83",X"00",X"02",X"CD",X"7B",X"03",X"E9",X"C3",X"01",X"0E",X"8D",X"FD",X"19",X"33",
		X"46",X"81",X"9D",X"C7",X"FB",X"02",X"0B",X"02",X"0B",X"06",X"0B",X"0A",X"0B",X"0E",X"0B",X"02",
		X"03",X"02",X"03",X"06",X"03",X"0A",X"03",X"0E",X"03",X"02",X"04",X"02",X"04",X"06",X"04",X"0A",
		X"04",X"0E",X"04",X"02",X"0C",X"02",X"0C",X"06",X"0C",X"0A",X"0C",X"0E",X"0C",X"C7",X"F3",X"10",
		X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",
		X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",
		X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",
		X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",
		X"41",X"3B",X"5B",X"81",X"FF",X"01",X"69",X"2A",X"FF",X"02",X"9B",X"21",X"1C",X"7E",X"01",X"DD",
		X"21",X"03",X"6B",X"03",X"8D",X"21",X"03",X"DD",X"25",X"05",X"6B",X"10",X"23",X"AD",X"82",X"7E",
		X"F8",X"33",X"7E",X"81",X"8D",X"14",X"1D",X"DD",X"94",X"1C",X"6B",X"01",X"23",X"5B",X"81",X"DD",
		X"0F",X"03",X"7F",X"E8",X"80",X"44",X"00",X"FF",X"18",X"2D",X"F6",X"F0",X"2A",X"27",X"E8",X"80",
		X"6D",X"7A",X"E0",X"AE",X"FF",X"9B",X"14",X"1C",X"2B",X"E9",X"80",X"AE",X"F4",X"21",X"06",X"70",
		X"D0",X"F3",X"77",X"E8",X"80",X"7E",X"FF",X"33",X"4C",X"81",X"8D",X"DE",X"26",X"DD",X"D0",X"26",
		X"8D",X"FB",X"1C",X"7E",X"00",X"DD",X"B8",X"02",X"7F",X"E8",X"80",X"77",X"77",X"E8",X"80",X"79",
		X"A4",X"30",X"E2",X"DD",X"D5",X"14",X"8D",X"77",X"1A",X"3B",X"46",X"81",X"E6",X"30",X"12",X"02",
		X"10",X"D5",X"6B",X"01",X"23",X"4C",X"81",X"DD",X"DE",X"26",X"8D",X"D0",X"26",X"C0",X"14",X"30",
		X"F0",X"EF",X"23",X"4C",X"81",X"DD",X"77",X"1A",X"2B",X"46",X"81",X"E7",X"61",X"20",X"6B",X"48",
		X"23",X"E7",X"80",X"02",X"06",X"D5",X"8D",X"D5",X"14",X"DD",X"77",X"1A",X"2B",X"46",X"81",X"E7",
		X"61",X"0C",X"2B",X"E7",X"80",X"D3",X"18",X"33",X"E7",X"80",X"95",X"55",X"61",X"E7",X"6B",X"02",
		X"23",X"5B",X"81",X"3B",X"DC",X"80",X"1A",X"5A",X"F6",X"3F",X"D6",X"01",X"23",X"DB",X"82",X"7E",
		X"FF",X"33",X"AD",X"82",X"6B",X"01",X"8D",X"65",X"03",X"7E",X"03",X"DD",X"65",X"03",X"8D",X"0F",
		X"03",X"DD",X"FB",X"1C",X"2B",X"AD",X"82",X"2C",X"61",X"0A",X"8D",X"72",X"25",X"3B",X"DF",X"80",
		X"3A",X"F3",X"03",X"68",X"23",X"AD",X"82",X"7E",X"01",X"33",X"44",X"80",X"8D",X"DE",X"26",X"DD",
		X"D0",X"26",X"8D",X"A4",X"26",X"EF",X"23",X"44",X"80",X"3B",X"45",X"80",X"F6",X"1F",X"61",X"0F",
		X"2B",X"45",X"80",X"F3",X"20",X"30",X"05",X"DD",X"6C",X"1E",X"0D",X"03",X"8D",X"44",X"1E",X"3B",
		X"75",X"80",X"E7",X"38",X"19",X"3B",X"00",X"B0",X"F6",X"08",X"69",X"12",X"6B",X"01",X"23",X"44",
		X"80",X"02",X"03",X"DD",X"81",X"1C",X"6B",X"01",X"23",X"AB",X"82",X"DD",X"B3",X"10",X"8D",X"0F",
		X"03",X"10",X"74",X"02",X"04",X"3B",X"DF",X"80",X"F6",X"03",X"5E",X"56",X"00",X"4C",X"00",X"49",
		X"8D",X"BB",X"11",X"C8",X"E9",X"70",X"DC",X"98",X"E9",X"76",X"00",X"01",X"2B",X"DF",X"80",X"1F",
		X"43",X"00",X"74",X"E1",X"1C",X"4C",X"7B",X"ED",X"76",X"01",X"2B",X"DF",X"80",X"F3",X"03",X"52",
		X"12",X"1F",X"74",X"E9",X"1C",X"4C",X"10",X"F6",X"88",X"02",X"04",X"6B",X"03",X"77",X"06",X"55",
		X"61",X"F9",X"E9",X"76",X"02",X"36",X"8D",X"83",X"11",X"E7",X"61",X"0E",X"E9",X"6B",X"01",X"A6",
		X"10",X"ED",X"76",X"01",X"E9",X"76",X"03",X"5B",X"0D",X"04",X"E9",X"76",X"03",X"34",X"9D",X"C7",
		X"FB",X"07",X"06",X"05",X"04",X"04",X"05",X"06",X"07",X"C0",X"C1",X"E0",X"E1",X"C2",X"C3",X"E2",
		X"E3",X"C4",X"C5",X"E4",X"E5",X"C6",X"C7",X"E6",X"E7",X"C7",X"F3",X"3B",X"DC",X"80",X"FF",X"05",
		X"C4",X"ED",X"74",X"DC",X"98",X"ED",X"7B",X"02",X"FF",X"06",X"C4",X"ED",X"63",X"00",X"00",X"ED",
		X"63",X"02",X"F0",X"C8",X"41",X"EF",X"23",X"31",X"81",X"33",X"30",X"81",X"74",X"00",X"9C",X"50",
		X"00",X"04",X"2B",X"DF",X"80",X"52",X"12",X"52",X"F6",X"08",X"F7",X"07",X"76",X"77",X"5A",X"6D",
		X"B4",X"30",X"EF",X"DD",X"63",X"07",X"8D",X"DD",X"27",X"0A",X"20",X"3B",X"31",X"81",X"D7",X"08",
		X"23",X"31",X"81",X"D5",X"8D",X"FC",X"1F",X"C0",X"1C",X"30",X"F0",X"DD",X"AF",X"1F",X"8D",X"67",
		X"1F",X"DD",X"DD",X"1F",X"8D",X"2C",X"1E",X"3B",X"E9",X"80",X"E7",X"30",X"03",X"DD",X"B0",X"1E",
		X"8D",X"0F",X"1F",X"C8",X"41",X"D5",X"C9",X"70",X"A6",X"1D",X"2B",X"DF",X"80",X"52",X"12",X"F3",
		X"1F",X"1F",X"43",X"00",X"C9",X"4C",X"C9",X"3A",X"00",X"CD",X"27",X"01",X"C9",X"1A",X"02",X"CD",
		X"74",X"80",X"93",X"ED",X"74",X"80",X"9F",X"44",X"E0",X"FF",X"3D",X"B2",X"69",X"08",X"C9",X"4C",
		X"E9",X"4C",X"72",X"55",X"61",X"F8",X"7B",X"52",X"F6",X"06",X"D6",X"F8",X"C9",X"37",X"00",X"ED",
		X"60",X"00",X"95",X"C8",X"C7",X"FB",X"C6",X"1D",X"14",X"00",X"DF",X"1D",X"1C",X"00",X"F8",X"1D",
		X"14",X"00",X"11",X"1E",X"1C",X"00",X"C6",X"1D",X"14",X"00",X"DF",X"1D",X"1C",X"00",X"F8",X"1D",
		X"14",X"00",X"11",X"1E",X"1C",X"00",X"00",X"00",X"03",X"00",X"00",X"02",X"00",X"00",X"00",X"03",
		X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"02",X"02",X"00",X"00",X"03",X"00",X"00",X"00",X"00",
		X"01",X"02",X"02",X"02",X"02",X"01",X"00",X"03",X"03",X"03",X"03",X"01",X"01",X"01",X"01",X"03",
		X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"03",X"03",X"03",X"00",X"03",
		X"00",X"00",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"00",X"03",X"00",X"03",X"03",X"03",X"03",X"00",X"00",X"02",X"02",X"00",X"00",X"00",X"01",
		X"01",X"02",X"01",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"C7",X"F3",X"41",X"02",X"00",X"DD",
		X"64",X"1D",X"51",X"6D",X"FF",X"19",X"61",X"F7",X"6B",X"4E",X"23",X"40",X"90",X"33",X"60",X"90",
		X"23",X"A0",X"93",X"C8",X"41",X"3B",X"31",X"81",X"AD",X"00",X"2A",X"3B",X"30",X"81",X"AD",X"00",
		X"22",X"44",X"40",X"00",X"18",X"2D",X"12",X"F3",X"01",X"17",X"2C",X"52",X"F6",X"1E",X"96",X"06",
		X"E7",X"38",X"05",X"55",X"8D",X"64",X"1D",X"54",X"8D",X"64",X"1D",X"C8",X"41",X"DD",X"44",X"1E",
		X"2B",X"31",X"81",X"FD",X"00",X"D3",X"40",X"5A",X"1A",X"5A",X"1A",X"F3",X"06",X"1F",X"C9",X"6B",
		X"00",X"86",X"F8",X"52",X"12",X"F3",X"18",X"87",X"D6",X"60",X"C9",X"37",X"00",X"3B",X"41",X"81",
		X"FF",X"7C",X"CC",X"AE",X"94",X"29",X"15",X"AE",X"AC",X"29",X"09",X"ED",X"7B",X"00",X"F7",X"40",
		X"E9",X"37",X"00",X"C8",X"E9",X"6B",X"00",X"A6",X"40",X"ED",X"76",X"00",X"C9",X"60",X"00",X"C8",
		X"41",X"70",X"ED",X"1E",X"2B",X"DF",X"80",X"52",X"12",X"F3",X"FC",X"56",X"00",X"1F",X"18",X"6B",
		X"23",X"E0",X"80",X"77",X"7B",X"33",X"E1",X"80",X"72",X"6B",X"23",X"E4",X"80",X"EF",X"23",X"E5",
		X"80",X"33",X"E6",X"80",X"72",X"6B",X"23",X"E2",X"80",X"EF",X"23",X"E3",X"80",X"3B",X"DF",X"80",
		X"23",X"BA",X"82",X"EF",X"23",X"31",X"81",X"33",X"30",X"81",X"9D",X"C7",X"FB",X"01",X"00",X"01",
		X"01",X"01",X"50",X"02",X"01",X"02",X"00",X"03",X"02",X"02",X"50",X"04",X"02",X"03",X"00",X"05",
		X"02",X"03",X"00",X"05",X"02",X"03",X"00",X"05",X"02",X"03",X"00",X"05",X"02",X"C7",X"F3",X"10",
		X"10",X"37",X"1F",X"DD",X"72",X"04",X"10",X"3F",X"1F",X"DD",X"72",X"04",X"10",X"48",X"1F",X"DD",
		X"72",X"04",X"10",X"51",X"1F",X"DD",X"72",X"04",X"10",X"59",X"1F",X"DD",X"C5",X"04",X"10",X"5F",
		X"1F",X"DD",X"C5",X"04",X"9D",X"C7",X"FB",X"FF",X"12",X"02",X"1C",X"1D",X"0E",X"19",X"FF",X"FF",
		X"13",X"02",X"19",X"18",X"12",X"17",X"1D",X"FF",X"FF",X"16",X"02",X"0B",X"18",X"17",X"1E",X"1C",
		X"FF",X"FF",X"17",X"02",X"1B",X"0A",X"1D",X"0E",X"FF",X"FF",X"14",X"03",X"E0",X"80",X"03",X"FF",
		X"18",X"02",X"E4",X"80",X"05",X"C7",X"F3",X"10",X"2B",X"DF",X"80",X"68",X"C9",X"70",X"9E",X"93",
		X"E9",X"70",X"9E",X"9F",X"74",X"9D",X"1F",X"50",X"C0",X"FF",X"53",X"CD",X"33",X"00",X"01",X"CD",
		X"33",X"01",X"01",X"CD",X"33",X"20",X"01",X"CD",X"33",X"21",X"72",X"43",X"E9",X"66",X"00",X"ED",
		X"33",X"01",X"72",X"CD",X"5C",X"ED",X"5C",X"2C",X"61",X"E0",X"9D",X"C7",X"FB",X"80",X"03",X"84",
		X"00",X"88",X"00",X"8C",X"03",X"80",X"03",X"84",X"00",X"88",X"00",X"8C",X"03",X"C7",X"F3",X"10",
		X"C9",X"70",X"00",X"90",X"E9",X"70",X"00",X"9C",X"10",X"20",X"00",X"02",X"20",X"CD",X"63",X"01",
		X"7E",X"CD",X"63",X"1E",X"7C",X"CD",X"63",X"1F",X"7D",X"CD",X"18",X"ED",X"63",X"01",X"02",X"ED",
		X"63",X"1E",X"02",X"ED",X"63",X"1F",X"02",X"ED",X"18",X"55",X"61",X"E1",X"9D",X"10",X"2B",X"D8",
		X"80",X"2C",X"E7",X"9D",X"C9",X"70",X"82",X"93",X"E9",X"70",X"82",X"9F",X"C9",X"76",X"00",X"7F",
		X"E9",X"76",X"00",X"0D",X"C9",X"77",X"E9",X"77",X"7D",X"30",X"F1",X"C8",X"41",X"3B",X"DF",X"80",
		X"12",X"52",X"12",X"52",X"12",X"F3",X"60",X"1F",X"2B",X"DC",X"80",X"70",X"E6",X"20",X"C3",X"1F",
		X"43",X"00",X"18",X"6B",X"FF",X"FF",X"DC",X"33",X"4F",X"81",X"C9",X"70",X"66",X"21",X"2B",X"4F",
		X"81",X"52",X"F6",X"FE",X"5E",X"56",X"00",X"CD",X"18",X"CD",X"2F",X"00",X"C9",X"32",X"01",X"3B",
		X"DD",X"80",X"5E",X"56",X"00",X"4C",X"7B",X"33",X"51",X"81",X"C9",X"70",X"60",X"22",X"E7",X"38",
		X"08",X"44",X"15",X"00",X"C9",X"4C",X"7D",X"30",X"FB",X"ED",X"74",X"08",X"90",X"3B",X"31",X"81",
		X"5E",X"56",X"00",X"ED",X"18",X"ED",X"18",X"ED",X"18",X"ED",X"18",X"F5",X"74",X"DE",X"2B",X"3B",
		X"DF",X"80",X"5E",X"56",X"00",X"4C",X"0F",X"ED",X"A5",X"E0",X"10",X"00",X"0C",X"4C",X"17",X"15",
		X"C9",X"6B",X"00",X"ED",X"76",X"00",X"60",X"77",X"C9",X"77",X"E9",X"77",X"14",X"30",X"F1",X"E0",
		X"2B",X"51",X"81",X"CD",X"74",X"97",X"24",X"52",X"12",X"52",X"F6",X"F8",X"5E",X"56",X"00",X"CD",
		X"18",X"ED",X"74",X"81",X"81",X"3B",X"31",X"81",X"F6",X"F8",X"CA",X"1F",X"9B",X"A3",X"20",X"9F",
		X"CF",X"D3",X"10",X"5A",X"F6",X"7F",X"5E",X"56",X"00",X"ED",X"18",X"02",X"08",X"CD",X"7B",X"00",
		X"E9",X"37",X"00",X"CD",X"72",X"ED",X"72",X"55",X"61",X"F3",X"2B",X"31",X"81",X"50",X"00",X"03",
		X"CA",X"26",X"69",X"03",X"54",X"01",X"03",X"DD",X"BB",X"11",X"2B",X"DD",X"80",X"D3",X"01",X"33",
		X"DD",X"80",X"72",X"6B",X"FF",X"FF",X"D4",X"3B",X"DC",X"80",X"D6",X"01",X"23",X"DC",X"80",X"EF",
		X"23",X"DD",X"80",X"C8",X"C7",X"FB",X"00",X"01",X"02",X"01",X"01",X"05",X"01",X"01",X"01",X"02",
		X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"05",X"05",X"01",X"01",X"02",X"01",X"01",X"08",X"0B",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"00",X"03",X"05",X"05",X"05",X"05",X"03",X"01",X"02",X"02",
		X"02",X"02",X"03",X"04",X"04",X"04",X"02",X"02",X"03",X"04",X"04",X"04",X"04",X"04",X"09",X"0B",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"00",X"01",X"01",X"02",X"02",X"02",X"01",X"02",X"01",X"01",
		X"02",X"03",X"04",X"04",X"04",X"04",X"04",X"05",X"05",X"06",X"07",X"05",X"06",X"06",X"0A",X"0B",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"00",X"02",X"01",X"02",X"02",X"02",X"02",X"01",X"01",X"05",
		X"05",X"01",X"01",X"01",X"03",X"01",X"05",X"03",X"02",X"02",X"02",X"02",X"02",X"02",X"0C",X"0B",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"80",X"21",X"94",X"21",X"A5",X"21",X"B6",X"21",X"C7",X"21",
		X"D8",X"21",X"E9",X"21",X"FA",X"21",X"0B",X"22",X"1C",X"22",X"2D",X"22",X"3E",X"22",X"4F",X"22",
		X"0E",X"0E",X"00",X"01",X"02",X"01",X"03",X"0B",X"08",X"0B",X"08",X"0B",X"08",X"0B",X"08",X"0B",
		X"08",X"0B",X"08",X"FF",X"0B",X"08",X"0B",X"08",X"0B",X"08",X"0B",X"08",X"0B",X"08",X"0B",X"08",
		X"0B",X"08",X"0B",X"08",X"FF",X"04",X"0C",X"06",X"07",X"06",X"07",X"06",X"07",X"06",X"07",X"06",
		X"07",X"06",X"07",X"06",X"07",X"FF",X"10",X"11",X"12",X"13",X"12",X"13",X"12",X"13",X"12",X"13",
		X"12",X"13",X"12",X"13",X"12",X"13",X"FF",X"12",X"13",X"12",X"13",X"12",X"13",X"12",X"13",X"12",
		X"13",X"12",X"13",X"12",X"13",X"12",X"13",X"FF",X"05",X"0A",X"09",X"0A",X"09",X"0A",X"09",X"0A",
		X"09",X"0A",X"09",X"0A",X"09",X"0A",X"05",X"0D",X"FF",X"14",X"15",X"16",X"17",X"16",X"17",X"16",
		X"17",X"16",X"17",X"16",X"17",X"16",X"17",X"16",X"17",X"FF",X"16",X"17",X"16",X"17",X"16",X"17",
		X"16",X"17",X"16",X"17",X"16",X"17",X"16",X"17",X"16",X"17",X"FF",X"0B",X"08",X"0B",X"08",X"0B",
		X"08",X"0B",X"08",X"0B",X"08",X"0B",X"08",X"0B",X"08",X"0B",X"0E",X"FF",X"12",X"13",X"12",X"13",
		X"12",X"13",X"12",X"13",X"12",X"13",X"12",X"13",X"12",X"13",X"12",X"18",X"FF",X"16",X"17",X"16",
		X"17",X"16",X"17",X"16",X"17",X"16",X"17",X"16",X"17",X"16",X"17",X"16",X"19",X"FF",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"06",
		X"07",X"06",X"07",X"06",X"07",X"06",X"07",X"06",X"07",X"06",X"07",X"06",X"07",X"06",X"1A",X"FF",
		X"51",X"53",X"51",X"51",X"53",X"51",X"51",X"53",X"58",X"59",X"5E",X"59",X"5F",X"53",X"51",X"51",
		X"53",X"51",X"51",X"53",X"51",X"51",X"53",X"42",X"43",X"53",X"42",X"43",X"53",X"56",X"52",X"5C",
		X"52",X"5D",X"53",X"42",X"43",X"53",X"42",X"43",X"53",X"51",X"51",X"53",X"4E",X"4F",X"53",X"4E",
		X"4F",X"53",X"56",X"57",X"5C",X"57",X"5D",X"53",X"4E",X"4F",X"53",X"4E",X"4F",X"53",X"51",X"51",
		X"53",X"4E",X"4F",X"53",X"4E",X"4F",X"53",X"54",X"55",X"5A",X"55",X"5B",X"53",X"4E",X"4F",X"53",
		X"4E",X"4F",X"53",X"51",X"51",X"53",X"42",X"43",X"53",X"42",X"43",X"53",X"51",X"51",X"53",X"51",
		X"51",X"53",X"42",X"43",X"53",X"42",X"43",X"53",X"51",X"51",X"53",X"51",X"51",X"53",X"51",X"51",
		X"53",X"42",X"43",X"53",X"42",X"43",X"53",X"51",X"51",X"53",X"51",X"51",X"53",X"51",X"51",X"53",
		X"42",X"43",X"53",X"42",X"43",X"53",X"52",X"52",X"52",X"52",X"52",X"53",X"42",X"43",X"53",X"42",
		X"43",X"53",X"51",X"51",X"53",X"4E",X"4F",X"53",X"4E",X"4F",X"53",X"52",X"52",X"52",X"52",X"52",
		X"53",X"4E",X"4F",X"53",X"4E",X"4F",X"53",X"51",X"51",X"53",X"4E",X"4F",X"53",X"4E",X"4F",X"53",
		X"4E",X"4F",X"53",X"4E",X"4F",X"53",X"4E",X"4F",X"53",X"4E",X"4F",X"53",X"51",X"51",X"53",X"52",
		X"52",X"52",X"52",X"52",X"53",X"42",X"43",X"53",X"42",X"43",X"53",X"52",X"52",X"52",X"52",X"52",
		X"53",X"51",X"51",X"53",X"52",X"52",X"52",X"52",X"52",X"53",X"4E",X"4F",X"53",X"4E",X"4F",X"53",
		X"52",X"52",X"52",X"52",X"52",X"53",X"51",X"51",X"53",X"42",X"43",X"53",X"42",X"43",X"53",X"42",
		X"43",X"53",X"42",X"43",X"53",X"42",X"43",X"53",X"42",X"43",X"53",X"51",X"51",X"53",X"4E",X"4F",
		X"53",X"4E",X"4F",X"53",X"51",X"51",X"53",X"51",X"51",X"53",X"4E",X"4F",X"53",X"4E",X"4F",X"53",
		X"51",X"51",X"53",X"51",X"51",X"53",X"51",X"51",X"53",X"4E",X"4F",X"53",X"4E",X"4F",X"53",X"51",
		X"51",X"53",X"51",X"51",X"53",X"51",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"52",X"52",X"52",X"52",X"52",
		X"52",X"52",X"52",X"52",X"52",X"52",X"52",X"52",X"52",X"52",X"52",X"52",X"52",X"52",X"52",X"52",
		X"51",X"53",X"51",X"51",X"53",X"42",X"43",X"53",X"42",X"43",X"53",X"42",X"43",X"53",X"42",X"43",
		X"53",X"51",X"51",X"53",X"51",X"51",X"53",X"51",X"51",X"53",X"4E",X"4F",X"53",X"4E",X"4F",X"53",
		X"4E",X"4F",X"53",X"4E",X"4F",X"53",X"51",X"51",X"53",X"51",X"52",X"52",X"52",X"51",X"53",X"42",
		X"43",X"53",X"42",X"43",X"53",X"42",X"43",X"53",X"42",X"43",X"53",X"51",X"52",X"52",X"52",X"52",
		X"52",X"52",X"51",X"53",X"4E",X"4F",X"53",X"4E",X"4F",X"53",X"4E",X"4F",X"53",X"4E",X"4F",X"53",
		X"51",X"52",X"52",X"52",X"52",X"52",X"52",X"51",X"53",X"51",X"51",X"53",X"42",X"43",X"53",X"42",
		X"43",X"53",X"51",X"51",X"53",X"51",X"52",X"52",X"52",X"52",X"52",X"52",X"51",X"53",X"51",X"51",
		X"53",X"4E",X"4F",X"53",X"4E",X"4F",X"53",X"51",X"51",X"53",X"51",X"52",X"52",X"52",X"52",X"52",
		X"52",X"52",X"52",X"52",X"51",X"53",X"42",X"43",X"53",X"42",X"43",X"53",X"51",X"52",X"52",X"52",
		X"52",X"52",X"52",X"52",X"52",X"52",X"52",X"52",X"52",X"51",X"53",X"4E",X"4F",X"53",X"4E",X"4F",
		X"53",X"51",X"52",X"52",X"52",X"52",X"52",X"52",X"52",X"52",X"52",X"50",X"50",X"50",X"50",X"50",
		X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"52",X"52",X"52",X"52",X"52",X"52",
		X"52",X"52",X"52",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"52",X"52",X"52",X"52",
		X"52",X"52",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"52",X"52",X"52",X"52",X"52",X"50",
		X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"80",X"80",X"FF",X"FF",X"80",X"80",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"80",X"80",X"80",X"80",X"80",X"80",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",
		X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"80",X"80",X"80",X"80",X"FF",X"FF",X"FF",
		X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"80",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"80",X"80",X"80",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"80",X"80",X"FF",X"FF",X"FF",X"FF",X"80",X"80",X"FF",X"FF",X"80",X"80",X"FF",X"FF",
		X"C7",X"F3",X"2B",X"56",X"81",X"06",X"12",X"C4",X"5E",X"56",X"00",X"ED",X"74",X"01",X"82",X"ED",
		X"18",X"ED",X"7B",X"00",X"FF",X"00",X"69",X"18",X"E9",X"1A",X"01",X"ED",X"07",X"02",X"8D",X"3B",
		X"26",X"6B",X"FF",X"00",X"69",X"0A",X"FF",X"80",X"69",X"06",X"FF",X"FF",X"69",X"02",X"0D",X"56",
		X"2B",X"22",X"81",X"F3",X"01",X"30",X"1E",X"FD",X"4A",X"BB",X"82",X"ED",X"60",X"01",X"E9",X"65",
		X"02",X"F5",X"C1",X"D5",X"74",X"BD",X"82",X"44",X"BB",X"82",X"54",X"1E",X"00",X"DD",X"4A",X"04",
		X"95",X"90",X"B5",X"09",X"15",X"3B",X"22",X"81",X"02",X"3B",X"45",X"80",X"F8",X"F3",X"0F",X"0E",
		X"E9",X"35",X"01",X"6D",X"F6",X"07",X"02",X"ED",X"35",X"02",X"8D",X"3B",X"26",X"6B",X"FF",X"80",
		X"69",X"06",X"FF",X"FF",X"69",X"02",X"0D",X"0E",X"E9",X"76",X"00",X"00",X"E9",X"76",X"01",X"00",
		X"E9",X"76",X"02",X"00",X"0D",X"2B",X"29",X"F3",X"0F",X"37",X"E9",X"76",X"00",X"01",X"E9",X"70",
		X"62",X"26",X"12",X"52",X"5E",X"56",X"00",X"ED",X"18",X"ED",X"7B",X"00",X"C9",X"37",X"00",X"ED",
		X"7B",X"01",X"C9",X"37",X"01",X"ED",X"7B",X"02",X"C9",X"37",X"20",X"ED",X"7B",X"03",X"C9",X"37",
		X"21",X"02",X"14",X"3B",X"DC",X"80",X"1A",X"F3",X"0F",X"C4",X"02",X"3B",X"56",X"81",X"29",X"E9",
		X"69",X"04",X"FF",X"28",X"2D",X"01",X"EE",X"33",X"56",X"81",X"9D",X"70",X"81",X"81",X"C9",X"70",
		X"E7",X"93",X"68",X"B2",X"69",X"0C",X"10",X"08",X"00",X"4C",X"10",X"40",X"00",X"CD",X"18",X"2C",
		X"61",X"F4",X"3D",X"B2",X"69",X"09",X"10",X"03",X"00",X"77",X"C9",X"4C",X"7D",X"30",X"FA",X"C8",
		X"C7",X"FB",X"4E",X"4F",X"42",X"43",X"4C",X"4D",X"42",X"43",X"4A",X"4B",X"42",X"43",X"48",X"49",
		X"42",X"43",X"46",X"47",X"42",X"43",X"44",X"45",X"40",X"41",X"44",X"45",X"40",X"41",X"44",X"45",
		X"40",X"41",X"44",X"45",X"40",X"41",X"44",X"45",X"40",X"41",X"44",X"45",X"40",X"41",X"44",X"45",
		X"40",X"41",X"46",X"47",X"42",X"43",X"48",X"49",X"42",X"43",X"4A",X"4B",X"42",X"43",X"4C",X"4D",
		X"42",X"43",X"C7",X"F3",X"41",X"70",X"92",X"98",X"17",X"04",X"2B",X"4C",X"81",X"AE",X"00",X"9D",
		X"F6",X"80",X"69",X"03",X"75",X"09",X"01",X"60",X"72",X"77",X"72",X"77",X"14",X"30",X"EB",X"3B",
		X"4C",X"81",X"CA",X"3F",X"61",X"04",X"D7",X"01",X"0D",X"02",X"D6",X"01",X"23",X"4C",X"81",X"C8",
		X"74",X"08",X"98",X"0A",X"15",X"3B",X"31",X"81",X"76",X"77",X"1C",X"30",X"FB",X"C8",X"2B",X"30",
		X"81",X"AE",X"F5",X"21",X"07",X"7E",X"01",X"33",X"AC",X"82",X"0D",X"19",X"1F",X"19",X"2B",X"DC",
		X"80",X"AE",X"02",X"30",X"02",X"0A",X"08",X"3B",X"7E",X"81",X"02",X"3B",X"31",X"81",X"D1",X"FC",
		X"6B",X"01",X"25",X"01",X"EE",X"33",X"AC",X"82",X"2B",X"4C",X"81",X"AE",X"00",X"38",X"32",X"EE",
		X"16",X"27",X"17",X"01",X"0D",X"02",X"17",X"FF",X"8D",X"42",X"27",X"3B",X"31",X"81",X"D0",X"33",
		X"31",X"81",X"02",X"3B",X"7E",X"81",X"F9",X"30",X"18",X"86",X"08",X"33",X"7E",X"81",X"8D",X"FC",
		X"1F",X"DD",X"8A",X"27",X"2B",X"31",X"81",X"E7",X"61",X"07",X"2B",X"30",X"81",X"2C",X"23",X"30",
		X"81",X"C8",X"74",X"5C",X"81",X"44",X"80",X"98",X"C9",X"70",X"5F",X"81",X"1F",X"04",X"7B",X"AE",
		X"00",X"38",X"07",X"CD",X"7B",X"00",X"D0",X"CD",X"76",X"00",X"85",X"6B",X"FF",X"F0",X"72",X"30",
		X"09",X"50",X"04",X"00",X"5C",X"BF",X"5C",X"BF",X"0D",X"06",X"54",X"04",X"00",X"DD",X"4A",X"04",
		X"54",X"03",X"00",X"58",X"54",X"08",X"00",X"CD",X"5C",X"C0",X"1C",X"30",X"D1",X"3B",X"DC",X"98",
		X"E6",X"9D",X"2B",X"DE",X"98",X"C4",X"23",X"DE",X"98",X"C8",X"2B",X"5B",X"81",X"AE",X"01",X"9D",
		X"2B",X"7E",X"81",X"F3",X"0F",X"95",X"2B",X"E0",X"80",X"06",X"2B",X"E1",X"80",X"0E",X"8D",X"A5",
		X"27",X"DD",X"DD",X"27",X"9D",X"3B",X"75",X"80",X"E7",X"9D",X"74",X"DB",X"80",X"3D",X"83",X"72",
		X"76",X"7F",X"3D",X"CB",X"32",X"37",X"7A",X"7E",X"00",X"CB",X"32",X"37",X"2B",X"DE",X"80",X"B2",
		X"D4",X"3B",X"7D",X"80",X"02",X"3B",X"D9",X"80",X"F9",X"8D",X"74",X"D8",X"80",X"60",X"8D",X"DD",
		X"1F",X"50",X"00",X"01",X"8D",X"BB",X"11",X"7E",X"01",X"33",X"DE",X"80",X"9D",X"3B",X"81",X"80",
		X"E7",X"30",X"07",X"44",X"F3",X"27",X"8D",X"C5",X"04",X"C8",X"10",X"F9",X"27",X"DD",X"C5",X"04",
		X"9D",X"C7",X"FB",X"FF",X"09",X"02",X"D9",X"80",X"06",X"FF",X"0D",X"02",X"D9",X"80",X"06",X"C7",
		X"F3",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",
		X"2B",X"20",X"81",X"2C",X"23",X"20",X"81",X"30",X"1A",X"DD",X"3E",X"11",X"2B",X"21",X"81",X"2C",
		X"23",X"21",X"81",X"30",X"0E",X"DD",X"94",X"11",X"2B",X"BA",X"82",X"AE",X"07",X"38",X"04",X"68",
		X"23",X"BA",X"82",X"3B",X"B8",X"82",X"FF",X"00",X"9B",X"63",X"28",X"AE",X"FF",X"9B",X"98",X"28",
		X"8D",X"70",X"2A",X"3B",X"DC",X"80",X"1A",X"5A",X"F6",X"3F",X"02",X"3B",X"DB",X"82",X"FF",X"07",
		X"69",X"09",X"F9",X"38",X"06",X"DD",X"8B",X"33",X"C2",X"A3",X"28",X"2F",X"DC",X"82",X"10",X"A3",
		X"28",X"C5",X"BD",X"3B",X"DC",X"80",X"1A",X"5A",X"F6",X"3F",X"02",X"3B",X"DB",X"82",X"F9",X"21",
		X"04",X"6D",X"23",X"DB",X"82",X"1F",X"43",X"00",X"2B",X"DF",X"80",X"52",X"12",X"52",X"C3",X"1F",
		X"74",X"C0",X"28",X"4C",X"5B",X"70",X"A8",X"28",X"18",X"4B",X"72",X"43",X"EA",X"27",X"DC",X"82",
		X"6B",X"01",X"23",X"B8",X"82",X"97",X"A3",X"28",X"EE",X"33",X"B8",X"82",X"2B",X"DB",X"82",X"68",
		X"23",X"DB",X"82",X"DD",X"0F",X"03",X"C7",X"FB",X"02",X"29",X"08",X"29",X"0E",X"29",X"9A",X"33",
		X"EB",X"2E",X"30",X"37",X"30",X"37",X"DB",X"38",X"66",X"3B",X"04",X"3E",X"1A",X"2C",X"80",X"33",
		X"16",X"00",X"06",X"02",X"08",X"04",X"14",X"14",X"16",X"04",X"0A",X"06",X"10",X"0E",X"14",X"14",
		X"16",X"04",X"0C",X"12",X"08",X"0E",X"14",X"14",X"16",X"10",X"06",X"04",X"0C",X"12",X"14",X"14",
		X"16",X"0A",X"04",X"0C",X"08",X"12",X"14",X"14",X"16",X"04",X"06",X"12",X"10",X"0E",X"14",X"14",
		X"16",X"04",X"06",X"0C",X"12",X"0E",X"14",X"14",X"16",X"10",X"12",X"06",X"0C",X"10",X"14",X"14",
		X"C7",X"F3",X"6B",X"0A",X"17",X"01",X"0D",X"0A",X"6B",X"08",X"17",X"02",X"0D",X"04",X"6B",X"05",
		X"17",X"03",X"23",X"A3",X"82",X"3B",X"BA",X"82",X"F6",X"04",X"69",X"01",X"51",X"6D",X"23",X"A4",
		X"82",X"10",X"2B",X"DC",X"80",X"F3",X"03",X"AE",X"03",X"30",X"06",X"7E",X"FF",X"33",X"B8",X"82",
		X"9D",X"DD",X"35",X"29",X"9D",X"7E",X"01",X"33",X"44",X"80",X"2B",X"31",X"81",X"F3",X"0F",X"93",
		X"6B",X"2A",X"2B",X"A4",X"82",X"0E",X"C9",X"70",X"5C",X"81",X"E9",X"70",X"83",X"82",X"C9",X"6B",
		X"00",X"AE",X"00",X"30",X"07",X"ED",X"7B",X"06",X"FF",X"01",X"61",X"0D",X"1C",X"9B",X"6B",X"2A",
		X"10",X"08",X"00",X"CD",X"18",X"ED",X"18",X"09",X"E5",X"D5",X"74",X"81",X"81",X"3B",X"31",X"81",
		X"F6",X"F0",X"D6",X"10",X"1A",X"06",X"2B",X"22",X"81",X"F3",X"07",X"52",X"12",X"52",X"0A",X"C4",
		X"F6",X"7F",X"5E",X"56",X"00",X"4C",X"A5",X"3D",X"12",X"0E",X"6B",X"F0",X"94",X"CD",X"76",X"03",
		X"2B",X"31",X"81",X"91",X"5E",X"56",X"00",X"70",X"27",X"90",X"18",X"4C",X"18",X"4C",X"E9",X"25",
		X"01",X"ED",X"24",X"02",X"B5",X"C0",X"1C",X"93",X"BA",X"29",X"1F",X"01",X"2B",X"39",X"81",X"06",
		X"6B",X"60",X"F9",X"21",X"0E",X"D3",X"18",X"5C",X"0D",X"F8",X"2B",X"22",X"81",X"52",X"12",X"F3",
		X"03",X"68",X"0A",X"02",X"00",X"6B",X"FF",X"00",X"69",X"09",X"72",X"40",X"6B",X"07",X"AE",X"38",
		X"0C",X"09",X"F2",X"47",X"E9",X"25",X"03",X"ED",X"24",X"04",X"1C",X"30",X"ED",X"EF",X"F9",X"9B",
		X"6B",X"2A",X"E9",X"3A",X"03",X"ED",X"27",X"04",X"63",X"FF",X"3D",X"52",X"12",X"52",X"0A",X"52",
		X"91",X"D3",X"38",X"CD",X"76",X"04",X"3D",X"52",X"D0",X"ED",X"07",X"01",X"D0",X"ED",X"76",X"01",
		X"C9",X"76",X"00",X"F0",X"C9",X"76",X"06",X"05",X"C9",X"76",X"07",X"01",X"2B",X"A3",X"82",X"ED",
		X"76",X"00",X"E9",X"76",X"07",X"01",X"2B",X"22",X"81",X"F3",X"03",X"06",X"6B",X"20",X"D0",X"CD",
		X"76",X"01",X"51",X"9F",X"4C",X"02",X"03",X"38",X"02",X"02",X"00",X"3B",X"DF",X"80",X"CA",X"06",
		X"3D",X"38",X"02",X"D3",X"10",X"CD",X"76",X"02",X"E9",X"76",X"06",X"01",X"E9",X"76",X"05",X"00",
		X"2B",X"DF",X"80",X"1F",X"43",X"00",X"74",X"E6",X"2B",X"4C",X"0F",X"ED",X"2F",X"01",X"E9",X"32",
		X"02",X"F5",X"C9",X"E0",X"10",X"00",X"0C",X"4C",X"60",X"77",X"60",X"CD",X"63",X"00",X"90",X"CD",
		X"63",X"01",X"91",X"CD",X"63",X"20",X"92",X"CD",X"63",X"21",X"93",X"EF",X"23",X"44",X"80",X"C8",
		X"C9",X"70",X"5C",X"81",X"E9",X"70",X"83",X"82",X"17",X"04",X"85",X"CD",X"7B",X"00",X"FF",X"00",
		X"61",X"07",X"E9",X"6B",X"06",X"AE",X"01",X"30",X"1C",X"ED",X"7B",X"07",X"FF",X"01",X"61",X"05",
		X"8D",X"B1",X"2A",X"09",X"10",X"AE",X"02",X"30",X"05",X"DD",X"7C",X"35",X"0D",X"07",X"FF",X"03",
		X"61",X"03",X"8D",X"5E",X"37",X"C0",X"14",X"9D",X"10",X"08",X"00",X"CD",X"18",X"ED",X"18",X"09",
		X"C9",X"ED",X"7B",X"06",X"FF",X"01",X"93",X"34",X"2B",X"ED",X"7B",X"00",X"D7",X"01",X"E9",X"37",
		X"00",X"93",X"34",X"2B",X"2B",X"A3",X"82",X"ED",X"76",X"00",X"E9",X"3A",X"01",X"ED",X"27",X"02",
		X"C9",X"F5",X"A5",X"CD",X"B5",X"70",X"10",X"2C",X"E9",X"4B",X"05",X"56",X"00",X"4C",X"7B",X"CD",
		X"76",X"00",X"29",X"CD",X"76",X"01",X"29",X"AE",X"50",X"30",X"02",X"7E",X"42",X"CD",X"76",X"20",
		X"29",X"CD",X"76",X"21",X"C9",X"E0",X"E9",X"6B",X"05",X"68",X"E9",X"37",X"05",X"AE",X"04",X"38",
		X"2A",X"AE",X"08",X"30",X"2F",X"3B",X"DF",X"80",X"5E",X"56",X"00",X"70",X"DE",X"2B",X"18",X"1A",
		X"E9",X"3A",X"01",X"ED",X"27",X"02",X"10",X"00",X"0C",X"4C",X"60",X"77",X"60",X"ED",X"2F",X"03",
		X"E9",X"32",X"04",X"76",X"00",X"ED",X"63",X"06",X"00",X"09",X"09",X"CD",X"63",X"05",X"01",X"CD",
		X"63",X"00",X"01",X"C8",X"C9",X"6B",X"05",X"AE",X"02",X"9B",X"A1",X"2B",X"FF",X"01",X"D4",X"CD",
		X"07",X"03",X"C9",X"6B",X"04",X"D3",X"05",X"0E",X"8D",X"C0",X"32",X"E7",X"61",X"0A",X"68",X"D3",
		X"05",X"0E",X"8D",X"C0",X"32",X"E7",X"69",X"1D",X"F6",X"80",X"69",X"0A",X"C9",X"76",X"07",X"80",
		X"C9",X"76",X"05",X"02",X"0D",X"08",X"C9",X"76",X"07",X"00",X"C9",X"76",X"05",X"02",X"54",X"02",
		X"03",X"DD",X"BB",X"11",X"9D",X"CD",X"75",X"06",X"61",X"0E",X"C9",X"76",X"06",X"08",X"C9",X"6B",
		X"07",X"AE",X"04",X"21",X"03",X"CD",X"21",X"07",X"C9",X"6B",X"03",X"CD",X"D3",X"07",X"C9",X"37",
		X"03",X"CD",X"7B",X"06",X"F6",X"03",X"61",X"43",X"C9",X"6B",X"01",X"FB",X"40",X"CD",X"76",X"01",
		X"9D",X"CD",X"7B",X"07",X"CA",X"3F",X"74",X"EE",X"2B",X"9B",X"AF",X"2B",X"74",X"FF",X"2B",X"52",
		X"F6",X"FE",X"5E",X"56",X"00",X"4C",X"7B",X"AE",X"FF",X"38",X"14",X"CD",X"0F",X"03",X"91",X"CD",
		X"76",X"03",X"72",X"6B",X"C9",X"1A",X"04",X"91",X"C9",X"37",X"04",X"CD",X"21",X"07",X"9D",X"CD",
		X"63",X"05",X"01",X"CD",X"63",X"06",X"05",X"CD",X"63",X"07",X"03",X"C8",X"C7",X"FB",X"07",X"1F",
		X"17",X"0F",X"17",X"0F",X"07",X"1F",X"01",X"19",X"11",X"09",X"11",X"09",X"01",X"19",X"04",X"03",
		X"04",X"03",X"03",X"02",X"02",X"02",X"01",X"01",X"FE",X"02",X"FE",X"03",X"FE",X"04",X"FF",X"04",
		X"FD",X"04",X"FD",X"03",X"FE",X"02",X"FE",X"01",X"FF",X"FE",X"FE",X"FE",X"FD",X"FE",X"FC",X"FF",
		X"90",X"94",X"98",X"9C",X"98",X"94",X"90",X"4E",X"C7",X"F3",X"2B",X"A5",X"82",X"AE",X"02",X"C6",
		X"B8",X"2C",X"FF",X"00",X"61",X"17",X"74",X"00",X"03",X"27",X"B5",X"82",X"6B",X"01",X"23",X"A5",
		X"82",X"50",X"00",X"02",X"8D",X"BB",X"11",X"7E",X"F0",X"33",X"DE",X"98",X"9D",X"3B",X"DC",X"80",
		X"F6",X"03",X"FF",X"00",X"9B",X"D9",X"2C",X"AE",X"02",X"21",X"08",X"3B",X"DD",X"80",X"FF",X"0A",
		X"9A",X"D9",X"2C",X"ED",X"74",X"DC",X"98",X"ED",X"63",X"02",X"F0",X"ED",X"63",X"03",X"50",X"ED",
		X"63",X"00",X"01",X"3B",X"22",X"81",X"F6",X"01",X"61",X"06",X"E9",X"76",X"01",X"00",X"0D",X"04",
		X"E9",X"76",X"01",X"10",X"74",X"28",X"2E",X"CD",X"74",X"E6",X"88",X"DD",X"4F",X"35",X"72",X"CD",
		X"74",X"E8",X"88",X"DD",X"4F",X"35",X"72",X"CD",X"74",X"EA",X"88",X"DD",X"4F",X"35",X"72",X"CD",
		X"74",X"C6",X"88",X"DD",X"4F",X"35",X"72",X"CD",X"74",X"C8",X"88",X"DD",X"4F",X"35",X"72",X"CD",
		X"74",X"CA",X"88",X"DD",X"4F",X"35",X"6B",X"02",X"8D",X"B8",X"02",X"7E",X"02",X"33",X"A5",X"82",
		X"23",X"A8",X"82",X"33",X"A9",X"82",X"0D",X"21",X"8D",X"9E",X"2D",X"DD",X"F8",X"2C",X"2B",X"AB",
		X"82",X"AE",X"02",X"38",X"2C",X"7E",X"01",X"DD",X"21",X"03",X"8D",X"30",X"2E",X"3B",X"AB",X"82",
		X"FF",X"01",X"69",X"1D",X"6B",X"01",X"8D",X"65",X"03",X"2F",X"B5",X"82",X"7A",X"27",X"B5",X"82",
		X"6D",X"A4",X"D4",X"7E",X"02",X"33",X"AB",X"82",X"54",X"07",X"04",X"DD",X"BB",X"11",X"8D",X"2D",
		X"11",X"DD",X"70",X"2E",X"8D",X"B3",X"10",X"C8",X"E9",X"70",X"DC",X"98",X"E9",X"9F",X"01",X"66",
		X"E9",X"6B",X"03",X"30",X"06",X"AE",X"80",X"21",X"08",X"09",X"0E",X"AE",X"04",X"29",X"02",X"09",
		X"08",X"ED",X"7B",X"01",X"FE",X"10",X"E9",X"37",X"01",X"3B",X"A5",X"82",X"CA",X"06",X"61",X"49",
		X"2B",X"DD",X"80",X"AE",X"02",X"29",X"04",X"AE",X"04",X"29",X"09",X"ED",X"7B",X"02",X"FF",X"B0",
		X"25",X"12",X"0D",X"07",X"E9",X"6B",X"02",X"AE",X"70",X"21",X"09",X"3B",X"A5",X"82",X"CA",X"96",
		X"23",X"A5",X"82",X"C8",X"E9",X"6B",X"02",X"86",X"02",X"ED",X"76",X"02",X"2B",X"45",X"80",X"F3",
		X"03",X"30",X"15",X"ED",X"CA",X"01",X"66",X"ED",X"7B",X"03",X"61",X"07",X"D6",X"01",X"E9",X"37",
		X"03",X"09",X"05",X"86",X"01",X"ED",X"76",X"03",X"9D",X"ED",X"7B",X"02",X"FF",X"C0",X"2D",X"09",
		X"2B",X"A5",X"82",X"9F",X"C6",X"33",X"A5",X"82",X"9D",X"3B",X"45",X"80",X"F6",X"03",X"61",X"15",
		X"E9",X"9F",X"01",X"66",X"E9",X"6B",X"03",X"30",X"07",X"D3",X"01",X"ED",X"76",X"03",X"0D",X"05",
		X"D7",X"01",X"E9",X"37",X"03",X"ED",X"7B",X"02",X"D6",X"02",X"E9",X"37",X"02",X"C8",X"2B",X"A8",
		X"82",X"86",X"01",X"AE",X"00",X"30",X"25",X"3B",X"A6",X"82",X"12",X"1F",X"12",X"87",X"5E",X"56",
		X"00",X"70",X"FE",X"2D",X"18",X"44",X"C5",X"88",X"54",X"06",X"00",X"DD",X"4A",X"04",X"2B",X"A6",
		X"82",X"68",X"FF",X"06",X"2D",X"01",X"EE",X"33",X"A6",X"82",X"6B",X"01",X"23",X"A8",X"82",X"3B",
		X"A9",X"82",X"D7",X"01",X"FF",X"00",X"61",X"20",X"2B",X"A7",X"82",X"1F",X"43",X"00",X"74",X"22",
		X"2E",X"4C",X"C9",X"70",X"CC",X"88",X"8D",X"4F",X"35",X"3B",X"A7",X"82",X"29",X"AE",X"06",X"CE",
		X"F3",X"2D",X"EE",X"33",X"A7",X"82",X"6B",X"01",X"23",X"A9",X"82",X"C8",X"C7",X"FB",X"00",X"00",
		X"08",X"09",X"28",X"29",X"00",X"00",X"0A",X"0B",X"2A",X"2B",X"0C",X"0D",X"2C",X"2D",X"00",X"00",
		X"0E",X"0F",X"2E",X"2F",X"00",X"00",X"0C",X"0D",X"2C",X"2D",X"00",X"00",X"00",X"00",X"0A",X"0B",
		X"2A",X"2B",X"48",X"4C",X"60",X"64",X"68",X"6C",X"04",X"24",X"44",X"00",X"20",X"40",X"C7",X"F3",
		X"2B",X"DE",X"98",X"06",X"8D",X"83",X"11",X"E7",X"61",X"07",X"2B",X"DF",X"98",X"D3",X"40",X"09",
		X"07",X"3B",X"DF",X"98",X"AD",X"00",X"D7",X"31",X"0A",X"DD",X"C0",X"32",X"E6",X"30",X"13",X"3D",
		X"D7",X"08",X"0A",X"DD",X"C0",X"32",X"E6",X"30",X"09",X"3D",X"D7",X"08",X"0A",X"DD",X"C0",X"32",
		X"E6",X"9D",X"8D",X"44",X"15",X"7E",X"01",X"33",X"AB",X"82",X"17",X"00",X"8D",X"81",X"1C",X"C8",
		X"C9",X"70",X"DC",X"98",X"C9",X"76",X"00",X"00",X"C9",X"70",X"DC",X"98",X"2B",X"A5",X"82",X"AE",
		X"00",X"38",X"14",X"CD",X"7B",X"02",X"D6",X"01",X"C9",X"37",X"02",X"AE",X"EC",X"29",X"08",X"EF",
		X"23",X"A5",X"82",X"CD",X"63",X"02",X"F0",X"3B",X"AB",X"82",X"FF",X"01",X"69",X"0B",X"8D",X"09",
		X"11",X"3B",X"A5",X"82",X"E6",X"30",X"27",X"09",X"36",X"70",X"92",X"98",X"17",X"04",X"7B",X"AE",
		X"EC",X"29",X"0D",X"70",X"90",X"98",X"17",X"10",X"63",X"00",X"72",X"55",X"61",X"FA",X"0D",X"1F",
		X"7B",X"D3",X"01",X"37",X"72",X"77",X"72",X"77",X"14",X"30",X"F5",X"DD",X"09",X"11",X"17",X"04",
		X"85",X"7E",X"02",X"DD",X"B8",X"02",X"8D",X"9E",X"2D",X"C0",X"14",X"30",X"F3",X"09",X"99",X"7E",
		X"0A",X"DD",X"B8",X"02",X"8D",X"09",X"11",X"E7",X"61",X"F5",X"9D",X"3B",X"7F",X"81",X"E6",X"30",
		X"0C",X"3B",X"DC",X"80",X"F6",X"03",X"FF",X"01",X"D4",X"DD",X"01",X"2F",X"9D",X"DD",X"2C",X"30",
		X"9D",X"10",X"2B",X"DD",X"80",X"AE",X"03",X"CE",X"21",X"2F",X"FF",X"09",X"25",X"48",X"D7",X"03",
		X"02",X"7E",X"01",X"33",X"44",X"80",X"8D",X"60",X"2F",X"DD",X"D4",X"2F",X"EE",X"33",X"44",X"80",
		X"9D",X"10",X"2B",X"AF",X"82",X"E7",X"D4",X"3B",X"22",X"81",X"12",X"F3",X"01",X"33",X"58",X"81",
		X"EE",X"33",X"80",X"81",X"23",X"5A",X"81",X"33",X"59",X"81",X"74",X"5C",X"81",X"44",X"83",X"82",
		X"17",X"20",X"EE",X"37",X"03",X"77",X"06",X"55",X"61",X"F8",X"54",X"01",X"04",X"DD",X"BB",X"11",
		X"6B",X"01",X"23",X"AF",X"82",X"C8",X"6B",X"01",X"23",X"7F",X"81",X"EF",X"23",X"AF",X"82",X"C8",
		X"41",X"3B",X"80",X"81",X"F9",X"95",X"3D",X"52",X"F6",X"FE",X"0A",X"02",X"00",X"3B",X"31",X"81",
		X"F6",X"F8",X"5E",X"56",X"00",X"AE",X"F8",X"30",X"03",X"44",X"F8",X"FF",X"2B",X"58",X"81",X"E7",
		X"61",X"06",X"C9",X"70",X"2B",X"90",X"0D",X"04",X"C9",X"70",X"36",X"90",X"41",X"CD",X"18",X"CD",
		X"18",X"CD",X"18",X"CD",X"18",X"ED",X"74",X"EC",X"31",X"ED",X"5C",X"ED",X"2F",X"00",X"E9",X"32",
		X"01",X"CD",X"A5",X"ED",X"B5",X"44",X"00",X"0C",X"E9",X"4C",X"41",X"6B",X"FF",X"FF",X"69",X"0E",
		X"C9",X"37",X"00",X"ED",X"63",X"00",X"17",X"ED",X"72",X"77",X"C9",X"77",X"0D",X"EC",X"2B",X"80",
		X"81",X"D3",X"01",X"33",X"80",X"81",X"FF",X"06",X"61",X"09",X"6B",X"01",X"23",X"7F",X"81",X"EF",
		X"23",X"AF",X"82",X"C8",X"41",X"3B",X"80",X"81",X"FF",X"04",X"69",X"32",X"FF",X"02",X"69",X"06",
		X"FF",X"05",X"80",X"2C",X"30",X"C8",X"2B",X"5C",X"81",X"AE",X"01",X"9D",X"2B",X"58",X"81",X"E7",
		X"74",X"76",X"32",X"30",X"03",X"70",X"96",X"32",X"41",X"44",X"5C",X"81",X"54",X"10",X"00",X"DD",
		X"4A",X"04",X"54",X"08",X"00",X"58",X"10",X"74",X"81",X"DD",X"4A",X"04",X"0D",X"1C",X"41",X"3B",
		X"6C",X"81",X"FF",X"01",X"DC",X"3B",X"58",X"81",X"E6",X"70",X"86",X"32",X"61",X"03",X"74",X"A6",
		X"32",X"44",X"6C",X"81",X"54",X"08",X"00",X"DD",X"4A",X"04",X"41",X"C8",X"41",X"3B",X"6C",X"81",
		X"E6",X"30",X"0D",X"EF",X"23",X"7F",X"81",X"33",X"AF",X"82",X"6B",X"FF",X"23",X"B8",X"82",X"C8",
		X"41",X"3B",X"59",X"81",X"E6",X"38",X"05",X"2C",X"23",X"59",X"81",X"C8",X"41",X"3B",X"DF",X"80",
		X"5E",X"56",X"00",X"70",X"B6",X"32",X"18",X"6B",X"23",X"59",X"81",X"3B",X"5A",X"81",X"12",X"1F",
		X"43",X"00",X"2B",X"58",X"81",X"E7",X"C9",X"70",X"16",X"32",X"61",X"04",X"C9",X"70",X"46",X"32",
		X"41",X"CD",X"18",X"CD",X"2F",X"00",X"C9",X"32",X"01",X"6B",X"23",X"5D",X"81",X"77",X"7B",X"33",
		X"65",X"81",X"72",X"6B",X"23",X"6D",X"81",X"77",X"7B",X"33",X"75",X"81",X"2B",X"5A",X"81",X"D3",
		X"01",X"F3",X"07",X"33",X"5A",X"81",X"FF",X"03",X"61",X"40",X"54",X"05",X"03",X"DD",X"BB",X"11",
		X"2B",X"58",X"81",X"E7",X"61",X"18",X"2B",X"5F",X"81",X"D3",X"0A",X"06",X"2B",X"60",X"81",X"D3",
		X"0E",X"0E",X"8D",X"C0",X"32",X"3D",X"D7",X"04",X"0A",X"DD",X"C0",X"32",X"0D",X"16",X"2B",X"5F",
		X"81",X"D3",X"0A",X"06",X"2B",X"60",X"81",X"D3",X"02",X"0E",X"8D",X"C0",X"32",X"3D",X"D6",X"04",
		X"0A",X"DD",X"C0",X"32",X"6B",X"30",X"8D",X"B8",X"02",X"C8",X"2B",X"5F",X"81",X"06",X"6B",X"C0",
		X"F9",X"8D",X"2B",X"DF",X"80",X"F3",X"02",X"7E",X"4F",X"38",X"02",X"7E",X"3F",X"E9",X"C4",X"3B",
		X"5A",X"81",X"FF",X"05",X"D4",X"3B",X"31",X"81",X"F6",X"0F",X"D4",X"DD",X"FF",X"30",X"9D",X"7E",
		X"01",X"33",X"44",X"80",X"C9",X"70",X"5C",X"81",X"54",X"08",X"00",X"56",X"18",X"3B",X"58",X"81",
		X"FE",X"01",X"23",X"58",X"81",X"10",X"C9",X"6B",X"01",X"FB",X"40",X"CD",X"76",X"01",X"2B",X"58",
		X"81",X"AE",X"01",X"CD",X"7B",X"04",X"61",X"03",X"96",X"09",X"01",X"D6",X"41",X"CD",X"76",X"04",
		X"C9",X"58",X"6B",X"20",X"96",X"17",X"FF",X"98",X"61",X"DB",X"2B",X"5F",X"81",X"06",X"2B",X"79",
		X"32",X"D3",X"10",X"C1",X"F6",X"F8",X"02",X"3B",X"31",X"81",X"F6",X"F8",X"D0",X"1F",X"43",X"00",
		X"2B",X"58",X"81",X"E7",X"61",X"0A",X"C9",X"70",X"0B",X"94",X"E9",X"70",X"16",X"94",X"0D",X"08",
		X"C9",X"70",X"16",X"94",X"E9",X"70",X"0B",X"94",X"41",X"CD",X"18",X"CD",X"18",X"CD",X"18",X"CD",
		X"18",X"ED",X"18",X"ED",X"18",X"ED",X"18",X"ED",X"18",X"CD",X"A5",X"CD",X"A5",X"ED",X"A5",X"CD",
		X"B5",X"50",X"00",X"08",X"C9",X"58",X"74",X"DE",X"2B",X"3B",X"DF",X"80",X"5E",X"56",X"00",X"4C",
		X"07",X"0A",X"52",X"2A",X"06",X"44",X"E0",X"FF",X"E9",X"35",X"00",X"ED",X"60",X"01",X"E9",X"35",
		X"02",X"ED",X"60",X"03",X"E9",X"4C",X"C9",X"65",X"00",X"CD",X"35",X"01",X"C9",X"65",X"02",X"CD",
		X"35",X"03",X"C9",X"4C",X"3C",X"30",X"E1",X"CD",X"B5",X"ED",X"B5",X"50",X"00",X"08",X"E9",X"58",
		X"74",X"F8",X"31",X"02",X"06",X"44",X"DC",X"FF",X"1F",X"04",X"E9",X"76",X"00",X"17",X"7B",X"CD",
		X"76",X"00",X"72",X"ED",X"72",X"CD",X"72",X"5D",X"61",X"F0",X"14",X"38",X"07",X"77",X"C9",X"4C",
		X"E9",X"4C",X"0D",X"E4",X"41",X"EF",X"23",X"44",X"80",X"C8",X"C7",X"FB",X"F8",X"31",X"FD",X"31",
		X"02",X"32",X"07",X"32",X"0C",X"32",X"11",X"32",X"0A",X"0B",X"2A",X"2B",X"FF",X"08",X"09",X"28",
		X"29",X"FF",X"06",X"07",X"26",X"27",X"FF",X"04",X"05",X"24",X"25",X"FF",X"02",X"03",X"22",X"23",
		X"FF",X"00",X"01",X"20",X"21",X"FF",X"26",X"32",X"2A",X"32",X"2E",X"32",X"32",X"32",X"36",X"32",
		X"3A",X"32",X"3E",X"32",X"42",X"32",X"4B",X"43",X"06",X"04",X"4C",X"44",X"0F",X"03",X"4D",X"45",
		X"06",X"04",X"4C",X"44",X"07",X"03",X"4B",X"43",X"47",X"04",X"4C",X"44",X"0E",X"03",X"4B",X"43",
		X"07",X"04",X"4C",X"44",X"4E",X"03",X"56",X"32",X"5A",X"32",X"5E",X"32",X"62",X"32",X"66",X"32",
		X"6A",X"32",X"6E",X"32",X"72",X"32",X"0B",X"03",X"46",X"44",X"0C",X"04",X"4F",X"43",X"0D",X"05",
		X"46",X"44",X"0C",X"04",X"47",X"43",X"0B",X"03",X"07",X"44",X"0C",X"04",X"4E",X"43",X"0B",X"03",
		X"47",X"44",X"0C",X"04",X"0E",X"43",X"01",X"4B",X"15",X"F0",X"98",X"00",X"00",X"00",X"01",X"43",
		X"15",X"F0",X"A8",X"00",X"00",X"00",X"01",X"04",X"15",X"F0",X"B8",X"00",X"00",X"00",X"01",X"04",
		X"15",X"F0",X"C8",X"00",X"00",X"00",X"01",X"0B",X"15",X"F0",X"80",X"00",X"00",X"00",X"01",X"03",
		X"15",X"F0",X"70",X"00",X"00",X"00",X"01",X"46",X"15",X"F0",X"60",X"00",X"00",X"00",X"01",X"44",
		X"15",X"F0",X"50",X"00",X"00",X"00",X"04",X"04",X"03",X"03",X"02",X"02",X"01",X"01",X"C7",X"F3",
		X"C9",X"F5",X"A5",X"C5",X"C9",X"70",X"32",X"81",X"37",X"04",X"C9",X"43",X"02",X"6D",X"86",X"CE",
		X"2C",X"33",X"FF",X"10",X"92",X"2C",X"33",X"5A",X"1A",X"F3",X"3F",X"17",X"C9",X"4B",X"03",X"3D",
		X"D2",X"CE",X"2C",X"33",X"FF",X"10",X"92",X"2C",X"33",X"5A",X"1A",X"F3",X"3F",X"1F",X"74",X"3E",
		X"33",X"CD",X"7B",X"00",X"F6",X"0F",X"12",X"52",X"96",X"C5",X"5E",X"56",X"00",X"4C",X"81",X"CD",
		X"CA",X"00",X"76",X"38",X"05",X"2B",X"3A",X"F3",X"03",X"1F",X"7B",X"48",X"4E",X"0C",X"61",X"FC",
		X"25",X"16",X"C9",X"9F",X"00",X"76",X"69",X"04",X"4B",X"81",X"0D",X"02",X"4B",X"01",X"2B",X"82",
		X"82",X"87",X"23",X"82",X"82",X"2B",X"0D",X"0F",X"6B",X"00",X"0D",X"0B",X"34",X"38",X"F9",X"44",
		X"04",X"00",X"C9",X"4C",X"C2",X"CA",X"32",X"90",X"B5",X"CD",X"B5",X"C8",X"C7",X"FB",X"0F",X"07",
		X"01",X"01",X"0F",X"01",X"01",X"00",X"07",X"0D",X"01",X"00",X"07",X"05",X"0D",X"00",X"01",X"03",
		X"07",X"0C",X"03",X"03",X"01",X"01",X"03",X"01",X"01",X"00",X"07",X"03",X"01",X"00",X"03",X"03",
		X"03",X"00",X"03",X"03",X"03",X"03",X"04",X"06",X"03",X"01",X"02",X"02",X"01",X"01",X"03",X"01",
		X"03",X"01",X"00",X"03",X"03",X"01",X"00",X"01",X"02",X"03",X"00",X"00",X"07",X"03",X"C7",X"F3",
		X"6B",X"FF",X"8D",X"B8",X"02",X"7E",X"FF",X"33",X"B8",X"82",X"9D",X"3B",X"BA",X"82",X"F6",X"03",
		X"E6",X"9D",X"29",X"33",X"A4",X"82",X"8D",X"4E",X"38",X"C8",X"2B",X"AF",X"82",X"E7",X"61",X"1D",
		X"2B",X"DC",X"80",X"F3",X"03",X"AE",X"03",X"30",X"06",X"7E",X"FF",X"33",X"B8",X"82",X"9D",X"AE",
		X"00",X"30",X"06",X"50",X"06",X"04",X"8D",X"BB",X"11",X"DD",X"E0",X"33",X"9D",X"3B",X"DC",X"80",
		X"F6",X"03",X"FF",X"03",X"69",X"13",X"2B",X"AF",X"82",X"AE",X"09",X"21",X"0C",X"9F",X"02",X"D9",
		X"EA",X"35",X"8D",X"45",X"34",X"DD",X"04",X"35",X"9D",X"DD",X"04",X"35",X"8D",X"BA",X"34",X"C8",
		X"E9",X"70",X"DC",X"98",X"E9",X"76",X"00",X"00",X"E9",X"76",X"02",X"F0",X"2B",X"AE",X"82",X"FB",
		X"01",X"F3",X"01",X"33",X"AE",X"82",X"61",X"0A",X"E9",X"76",X"01",X"02",X"E9",X"76",X"03",X"F0",
		X"0D",X"08",X"E9",X"76",X"01",X"12",X"E9",X"76",X"03",X"90",X"8D",X"83",X"11",X"E7",X"61",X"08",
		X"E9",X"6B",X"03",X"D3",X"20",X"ED",X"76",X"03",X"C9",X"70",X"C6",X"88",X"74",X"62",X"35",X"DD",
		X"4F",X"35",X"C9",X"70",X"C8",X"88",X"72",X"DD",X"4F",X"35",X"C9",X"70",X"E6",X"88",X"72",X"DD",
		X"4F",X"35",X"C9",X"70",X"E8",X"88",X"72",X"DD",X"4F",X"35",X"6B",X"30",X"23",X"B0",X"82",X"7E",
		X"01",X"33",X"AF",X"82",X"9D",X"ED",X"74",X"DC",X"98",X"3B",X"AF",X"82",X"CA",X"06",X"69",X"35",
		X"E9",X"6B",X"02",X"AE",X"B0",X"21",X"09",X"3B",X"AF",X"82",X"D6",X"01",X"23",X"AF",X"82",X"C8",
		X"2B",X"45",X"80",X"F3",X"03",X"30",X"15",X"3B",X"AE",X"82",X"E6",X"ED",X"7B",X"03",X"61",X"07",
		X"D6",X"01",X"E9",X"37",X"03",X"09",X"05",X"86",X"01",X"ED",X"76",X"03",X"E9",X"6B",X"02",X"86",
		X"01",X"ED",X"76",X"02",X"9D",X"ED",X"7B",X"02",X"FF",X"D0",X"2D",X"09",X"2B",X"AF",X"82",X"D3",
		X"01",X"33",X"AF",X"82",X"9D",X"3B",X"45",X"80",X"F6",X"03",X"61",X"15",X"2B",X"AE",X"82",X"E7",
		X"E9",X"6B",X"03",X"30",X"07",X"D3",X"01",X"ED",X"76",X"03",X"0D",X"05",X"D7",X"01",X"E9",X"37",
		X"03",X"ED",X"7B",X"02",X"D6",X"01",X"E9",X"37",X"02",X"C8",X"E9",X"70",X"DC",X"98",X"E9",X"6B",
		X"02",X"AE",X"E8",X"29",X"1A",X"EF",X"23",X"B1",X"82",X"33",X"AF",X"82",X"E9",X"76",X"02",X"F0",
		X"E9",X"76",X"00",X"00",X"6B",X"C0",X"8D",X"1E",X"3F",X"7E",X"D0",X"DD",X"1E",X"3F",X"9D",X"3B",
		X"45",X"80",X"F6",X"03",X"61",X"15",X"2B",X"AE",X"82",X"E7",X"E9",X"6B",X"03",X"30",X"07",X"D3",
		X"01",X"ED",X"76",X"03",X"0D",X"05",X"D7",X"01",X"E9",X"37",X"03",X"ED",X"7B",X"02",X"D6",X"01",
		X"E9",X"37",X"02",X"C8",X"2B",X"B0",X"82",X"E7",X"69",X"05",X"7D",X"33",X"B0",X"82",X"9D",X"3B",
		X"B1",X"82",X"12",X"52",X"5E",X"56",X"00",X"70",X"62",X"35",X"18",X"CD",X"74",X"C6",X"88",X"DD",
		X"4F",X"35",X"72",X"CD",X"74",X"C8",X"88",X"DD",X"4F",X"35",X"72",X"CD",X"74",X"E6",X"88",X"DD",
		X"4F",X"35",X"72",X"CD",X"74",X"E8",X"88",X"DD",X"4F",X"35",X"2B",X"AF",X"82",X"F3",X"01",X"33",
		X"B0",X"82",X"2B",X"B1",X"82",X"68",X"FF",X"06",X"2D",X"01",X"EE",X"33",X"B1",X"82",X"9D",X"6B",
		X"C9",X"37",X"00",X"68",X"C9",X"37",X"01",X"68",X"C9",X"37",X"10",X"68",X"C9",X"37",X"11",X"C8",
		X"C7",X"FB",X"10",X"30",X"14",X"34",X"18",X"38",X"1C",X"3C",X"50",X"70",X"54",X"74",X"58",X"78",
		X"5C",X"7C",X"50",X"70",X"54",X"74",X"18",X"38",X"1C",X"3C",X"C7",X"F3",X"C9",X"6B",X"05",X"AE",
		X"01",X"38",X"1A",X"CD",X"75",X"06",X"D4",X"CD",X"7B",X"01",X"29",X"0E",X"F6",X"03",X"61",X"05",
		X"C9",X"76",X"00",X"00",X"9D",X"CD",X"60",X"01",X"C9",X"76",X"06",X"03",X"9D",X"CD",X"07",X"03",
		X"C9",X"6B",X"04",X"D3",X"08",X"0E",X"8D",X"C0",X"32",X"E7",X"69",X"0B",X"41",X"10",X"41",X"10",
		X"41",X"10",X"C9",X"76",X"05",X"02",X"9D",X"ED",X"75",X"02",X"61",X"10",X"E9",X"6B",X"05",X"ED",
		X"76",X"02",X"6B",X"05",X"E9",X"FF",X"03",X"29",X"03",X"ED",X"21",X"03",X"C9",X"6B",X"03",X"ED",
		X"D3",X"03",X"C9",X"37",X"03",X"ED",X"75",X"00",X"61",X"0F",X"C9",X"6B",X"04",X"ED",X"83",X"01",
		X"C9",X"37",X"04",X"ED",X"7B",X"04",X"E9",X"37",X"00",X"C8",X"2B",X"20",X"81",X"F3",X"07",X"95",
		X"2B",X"BA",X"82",X"F3",X"02",X"D3",X"02",X"06",X"C9",X"70",X"5C",X"81",X"E9",X"70",X"83",X"82",
		X"10",X"08",X"00",X"CD",X"7B",X"00",X"E6",X"30",X"07",X"ED",X"7B",X"06",X"FF",X"01",X"61",X"08",
		X"14",X"9D",X"C9",X"4C",X"E9",X"4C",X"0D",X"EB",X"54",X"04",X"03",X"DD",X"BB",X"11",X"2B",X"35",
		X"81",X"17",X"2B",X"DF",X"98",X"1F",X"2B",X"AE",X"82",X"E7",X"61",X"2D",X"2B",X"81",X"80",X"E7",
		X"3E",X"38",X"02",X"D3",X"80",X"FD",X"00",X"86",X"50",X"D6",X"4B",X"03",X"2D",X"0B",X"FF",X"18",
		X"2D",X"07",X"5D",X"38",X"04",X"86",X"10",X"09",X"F5",X"DD",X"83",X"11",X"E6",X"30",X"05",X"70",
		X"F4",X"36",X"0D",X"31",X"74",X"04",X"37",X"09",X"2C",X"DD",X"83",X"11",X"E6",X"2B",X"61",X"03",
		X"D7",X"80",X"5E",X"FD",X"00",X"86",X"30",X"D6",X"4B",X"03",X"25",X"0B",X"FF",X"D8",X"25",X"07",
		X"5D",X"38",X"04",X"D3",X"10",X"09",X"F5",X"DD",X"83",X"11",X"E6",X"30",X"05",X"70",X"04",X"37",
		X"0D",X"03",X"74",X"F4",X"36",X"2B",X"12",X"52",X"5E",X"56",X"00",X"4C",X"7B",X"ED",X"76",X"00",
		X"E9",X"37",X"04",X"77",X"7B",X"ED",X"76",X"01",X"72",X"6B",X"E9",X"37",X"02",X"ED",X"76",X"05",
		X"E9",X"76",X"03",X"01",X"E9",X"76",X"06",X"00",X"E9",X"76",X"07",X"02",X"C9",X"76",X"00",X"01",
		X"2B",X"22",X"81",X"9F",X"2A",X"38",X"0A",X"CD",X"63",X"01",X"28",X"CD",X"63",X"02",X"03",X"09",
		X"08",X"CD",X"63",X"01",X"2C",X"CD",X"63",X"02",X"05",X"CD",X"63",X"05",X"01",X"CD",X"63",X"06",
		X"03",X"CD",X"63",X"07",X"00",X"3B",X"DE",X"98",X"C9",X"37",X"03",X"DD",X"83",X"11",X"E6",X"3B",
		X"DF",X"98",X"69",X"08",X"AD",X"00",X"D7",X"40",X"C9",X"37",X"04",X"C8",X"D6",X"30",X"C9",X"37",
		X"04",X"C8",X"C7",X"FB",X"01",X"01",X"08",X"00",X"02",X"02",X"08",X"00",X"02",X"01",X"08",X"00",
		X"01",X"00",X"08",X"00",X"01",X"FF",X"08",X"00",X"02",X"FE",X"08",X"00",X"02",X"FF",X"08",X"00",
		X"01",X"00",X"08",X"00",X"C7",X"F3",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",
		X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",
		X"2B",X"DC",X"80",X"F3",X"03",X"AE",X"03",X"30",X"06",X"7E",X"FF",X"33",X"B8",X"82",X"9D",X"3B",
		X"BA",X"82",X"12",X"1F",X"43",X"00",X"74",X"32",X"3F",X"4C",X"7B",X"33",X"A3",X"82",X"02",X"3B",
		X"20",X"81",X"F0",X"30",X"08",X"77",X"7B",X"33",X"A4",X"82",X"8D",X"4E",X"38",X"C8",X"C9",X"6B",
		X"05",X"AE",X"01",X"95",X"C9",X"6B",X"03",X"AE",X"90",X"21",X"37",X"AE",X"50",X"29",X"47",X"CD",
		X"7B",X"01",X"F6",X"03",X"12",X"06",X"12",X"C4",X"5E",X"56",X"00",X"70",X"4A",X"3F",X"18",X"5E",
		X"03",X"CD",X"7B",X"03",X"83",X"06",X"72",X"CD",X"7B",X"04",X"83",X"0E",X"8D",X"C0",X"32",X"0C",
		X"72",X"30",X"EE",X"3B",X"82",X"82",X"F6",X"0E",X"69",X"1C",X"54",X"03",X"03",X"DD",X"BB",X"11",
		X"0D",X"14",X"E9",X"24",X"00",X"30",X"0F",X"CD",X"7B",X"04",X"E9",X"C3",X"01",X"CD",X"76",X"04",
		X"E9",X"6B",X"04",X"ED",X"76",X"00",X"C9",X"6B",X"03",X"ED",X"83",X"03",X"C9",X"37",X"03",X"ED",
		X"75",X"02",X"61",X"2C",X"E9",X"6B",X"05",X"ED",X"76",X"02",X"6B",X"FB",X"E9",X"24",X"03",X"ED",
		X"FB",X"03",X"2D",X"1C",X"54",X"01",X"01",X"DD",X"BB",X"11",X"C9",X"6B",X"03",X"AE",X"90",X"29",
		X"0B",X"CD",X"7B",X"04",X"FF",X"48",X"2D",X"04",X"FF",X"C8",X"2D",X"3A",X"E9",X"76",X"03",X"FC",
		X"C9",X"24",X"06",X"30",X"30",X"CD",X"5B",X"07",X"43",X"00",X"74",X"62",X"3F",X"4C",X"C9",X"6B",
		X"01",X"9F",X"56",X"6B",X"69",X"02",X"D6",X"04",X"C9",X"37",X"01",X"48",X"6B",X"06",X"FA",X"30",
		X"01",X"4E",X"C9",X"23",X"07",X"3B",X"22",X"81",X"F6",X"07",X"5E",X"56",X"00",X"70",X"68",X"3F",
		X"18",X"6B",X"C9",X"37",X"06",X"C8",X"2B",X"22",X"81",X"F3",X"07",X"52",X"12",X"1F",X"43",X"00",
		X"74",X"70",X"3F",X"4C",X"7B",X"ED",X"76",X"00",X"E9",X"37",X"04",X"77",X"7B",X"ED",X"76",X"01",
		X"72",X"6B",X"E9",X"37",X"02",X"ED",X"76",X"05",X"72",X"6B",X"E9",X"37",X"03",X"C8",X"2B",X"A4",
		X"82",X"06",X"C9",X"70",X"5C",X"81",X"E9",X"70",X"83",X"82",X"10",X"08",X"00",X"CD",X"7B",X"00",
		X"E6",X"30",X"07",X"ED",X"7B",X"06",X"FF",X"01",X"61",X"08",X"14",X"9D",X"C9",X"4C",X"E9",X"4C",
		X"0D",X"EB",X"54",X"01",X"01",X"DD",X"BB",X"11",X"6B",X"01",X"23",X"44",X"80",X"CD",X"63",X"00",
		X"01",X"CD",X"63",X"02",X"18",X"CD",X"63",X"03",X"F0",X"CD",X"63",X"05",X"01",X"3B",X"20",X"81",
		X"CA",X"06",X"61",X"06",X"C9",X"76",X"01",X"28",X"0D",X"04",X"C9",X"76",X"01",X"2C",X"2B",X"22",
		X"81",X"F3",X"07",X"1F",X"43",X"00",X"74",X"42",X"3F",X"4C",X"7B",X"CD",X"76",X"04",X"74",X"68",
		X"3F",X"4C",X"7B",X"CD",X"76",X"06",X"E9",X"76",X"02",X"08",X"E9",X"76",X"03",X"FF",X"E9",X"76",
		X"05",X"04",X"E9",X"76",X"07",X"03",X"EE",X"CD",X"76",X"07",X"E9",X"37",X"00",X"ED",X"76",X"01",
		X"E9",X"37",X"04",X"ED",X"76",X"06",X"EE",X"33",X"44",X"80",X"9D",X"ED",X"74",X"DC",X"98",X"3B",
		X"B8",X"82",X"FF",X"01",X"69",X"14",X"FF",X"02",X"69",X"08",X"FF",X"03",X"69",X"08",X"8D",X"14",
		X"3B",X"C8",X"8D",X"AA",X"39",X"C8",X"8D",X"CD",X"3A",X"C8",X"8D",X"FE",X"38",X"C8",X"6B",X"01",
		X"23",X"44",X"80",X"3B",X"B1",X"82",X"E6",X"38",X"07",X"2C",X"69",X"3A",X"7D",X"9B",X"61",X"39",
		X"54",X"01",X"02",X"DD",X"BB",X"11",X"E9",X"76",X"00",X"01",X"E9",X"76",X"01",X"01",X"E9",X"76",
		X"02",X"F0",X"2B",X"22",X"81",X"F3",X"3F",X"D3",X"40",X"ED",X"76",X"03",X"74",X"01",X"0C",X"27",
		X"B5",X"82",X"C9",X"70",X"E6",X"88",X"74",X"90",X"3F",X"DD",X"4F",X"35",X"C9",X"77",X"C9",X"77",
		X"72",X"DD",X"4F",X"35",X"0D",X"3F",X"E9",X"6B",X"02",X"AE",X"E6",X"21",X"3F",X"CD",X"74",X"C6",
		X"88",X"70",X"92",X"3F",X"8D",X"4F",X"35",X"CD",X"72",X"CD",X"72",X"77",X"8D",X"4F",X"35",X"09",
		X"24",X"ED",X"7B",X"02",X"FF",X"D6",X"25",X"24",X"C9",X"70",X"A6",X"88",X"74",X"94",X"3F",X"DD",
		X"4F",X"35",X"C9",X"77",X"C9",X"77",X"72",X"DD",X"4F",X"35",X"6B",X"02",X"23",X"B8",X"82",X"EF",
		X"23",X"B1",X"82",X"09",X"18",X"3B",X"B1",X"82",X"29",X"33",X"B1",X"82",X"17",X"02",X"8D",X"91",
		X"3A",X"02",X"01",X"DD",X"4B",X"3A",X"E9",X"76",X"00",X"00",X"C2",X"A5",X"39",X"ED",X"63",X"00",
		X"01",X"10",X"41",X"10",X"41",X"EF",X"23",X"44",X"80",X"C8",X"2B",X"DC",X"80",X"F3",X"03",X"AE",
		X"02",X"21",X"0B",X"2F",X"B5",X"82",X"7A",X"27",X"B5",X"82",X"6D",X"A4",X"61",X"08",X"6B",X"04",
		X"23",X"B8",X"82",X"97",X"46",X"3A",X"E9",X"12",X"02",X"DD",X"83",X"11",X"E6",X"30",X"09",X"56",
		X"00",X"ED",X"7B",X"03",X"D6",X"38",X"0D",X"09",X"43",X"01",X"E9",X"6B",X"03",X"FD",X"00",X"86",
		X"3A",X"0E",X"6B",X"01",X"8D",X"21",X"03",X"DD",X"C0",X"32",X"E6",X"38",X"46",X"9F",X"7E",X"30",
		X"12",X"3B",X"3E",X"81",X"F6",X"0F",X"FF",X"05",X"2B",X"41",X"81",X"21",X"02",X"D3",X"08",X"D3",
		X"04",X"09",X"10",X"3B",X"3A",X"81",X"F6",X"0F",X"FF",X"05",X"2B",X"3D",X"81",X"29",X"02",X"D3",
		X"08",X"D3",X"04",X"04",X"69",X"04",X"D7",X"38",X"0D",X"04",X"AD",X"00",X"D7",X"3A",X"E9",X"37",
		X"03",X"50",X"08",X"04",X"8D",X"BB",X"11",X"7E",X"03",X"33",X"B8",X"82",X"6B",X"80",X"23",X"B1",
		X"82",X"09",X"13",X"7E",X"01",X"DD",X"65",X"03",X"17",X"01",X"8D",X"4B",X"3A",X"02",X"01",X"DD",
		X"91",X"3A",X"8D",X"8B",X"33",X"C8",X"EE",X"33",X"DC",X"98",X"9D",X"3B",X"B5",X"82",X"CA",X"06",
		X"DC",X"3B",X"AF",X"82",X"CA",X"06",X"61",X"14",X"2B",X"B5",X"82",X"9F",X"76",X"30",X"1A",X"ED",
		X"7B",X"02",X"D1",X"ED",X"76",X"02",X"FF",X"6E",X"2D",X"0F",X"0D",X"14",X"E9",X"6B",X"02",X"AE",
		X"90",X"21",X"06",X"C4",X"E9",X"37",X"02",X"09",X"07",X"3B",X"AF",X"82",X"29",X"33",X"AF",X"82",
		X"E9",X"6B",X"02",X"AE",X"80",X"21",X"05",X"ED",X"63",X"00",X"00",X"C8",X"E9",X"76",X"00",X"01",
		X"9D",X"3B",X"B5",X"82",X"CA",X"06",X"D4",X"3B",X"AE",X"82",X"E6",X"30",X"20",X"ED",X"7B",X"03",
		X"D0",X"ED",X"76",X"03",X"8D",X"83",X"11",X"E7",X"61",X"04",X"1F",X"A0",X"0D",X"02",X"1F",X"80",
		X"E9",X"6B",X"03",X"FC",X"2D",X"16",X"6B",X"01",X"23",X"AE",X"82",X"09",X"0F",X"ED",X"7B",X"03",
		X"D1",X"ED",X"76",X"03",X"FF",X"F0",X"2D",X"04",X"EE",X"33",X"AE",X"82",X"9D",X"DD",X"44",X"15",
		X"2B",X"B1",X"82",X"E7",X"61",X"24",X"8D",X"77",X"1A",X"3B",X"46",X"81",X"02",X"3B",X"47",X"81",
		X"D0",X"38",X"29",X"EF",X"23",X"81",X"82",X"33",X"82",X"82",X"6B",X"04",X"23",X"B8",X"82",X"7E",
		X"80",X"33",X"81",X"81",X"6B",X"01",X"8D",X"65",X"03",X"C8",X"2B",X"4C",X"81",X"E7",X"61",X"0C",
		X"6B",X"FF",X"23",X"4C",X"81",X"3B",X"B1",X"82",X"7D",X"33",X"B1",X"82",X"6B",X"04",X"8D",X"B8",
		X"02",X"97",X"CD",X"3A",X"E9",X"6B",X"02",X"D3",X"02",X"ED",X"76",X"02",X"2B",X"B1",X"82",X"AE",
		X"00",X"ED",X"7B",X"02",X"61",X"15",X"FF",X"D8",X"2D",X"2E",X"6B",X"A0",X"8D",X"1E",X"3F",X"7E",
		X"B0",X"DD",X"1E",X"3F",X"6B",X"01",X"23",X"B1",X"82",X"09",X"1D",X"AE",X"EC",X"29",X"19",X"ED",
		X"63",X"02",X"F0",X"7E",X"FF",X"33",X"B8",X"82",X"EE",X"33",X"AF",X"82",X"6B",X"C0",X"8D",X"1E",
		X"3F",X"7E",X"D0",X"DD",X"1E",X"3F",X"0D",X"0D",X"17",X"02",X"8D",X"91",X"3A",X"3B",X"B5",X"82",
		X"FE",X"01",X"23",X"B5",X"82",X"C8",X"2B",X"B8",X"82",X"AE",X"01",X"30",X"04",X"DD",X"75",X"3B",
		X"9D",X"DD",X"65",X"3C",X"9D",X"ED",X"74",X"DC",X"98",X"3B",X"DC",X"80",X"F6",X"03",X"FF",X"01",
		X"D4",X"50",X"02",X"02",X"8D",X"BB",X"11",X"7E",X"01",X"33",X"44",X"80",X"23",X"B0",X"82",X"ED",
		X"63",X"00",X"01",X"DD",X"83",X"11",X"E6",X"ED",X"63",X"01",X"05",X"30",X"04",X"ED",X"63",X"01",
		X"15",X"ED",X"63",X"02",X"F0",X"3B",X"DF",X"80",X"F6",X"03",X"5E",X"56",X"00",X"DD",X"83",X"11",
		X"E6",X"30",X"07",X"70",X"B2",X"3F",X"1F",X"02",X"0D",X"05",X"74",X"B6",X"3F",X"0A",X"01",X"4C",
		X"7B",X"ED",X"76",X"03",X"C9",X"70",X"E4",X"88",X"74",X"AE",X"3F",X"02",X"04",X"DD",X"4F",X"35",
		X"72",X"CD",X"72",X"CD",X"72",X"55",X"61",X"F5",X"74",X"BA",X"3F",X"4C",X"07",X"DD",X"EA",X"3B",
		X"6B",X"02",X"23",X"B8",X"82",X"EF",X"23",X"44",X"80",X"C8",X"C9",X"70",X"5C",X"81",X"E9",X"70",
		X"83",X"82",X"C9",X"76",X"00",X"01",X"C9",X"76",X"01",X"18",X"C9",X"76",X"02",X"02",X"C9",X"76",
		X"03",X"F0",X"C9",X"76",X"06",X"03",X"E9",X"76",X"07",X"04",X"3D",X"F3",X"01",X"ED",X"76",X"00",
		X"CA",X"11",X"2B",X"DF",X"98",X"38",X"16",X"FD",X"00",X"9F",X"44",X"38",X"0C",X"86",X"19",X"CD",
		X"63",X"01",X"58",X"CD",X"63",X"07",X"0C",X"09",X"16",X"86",X"69",X"09",X"12",X"9F",X"44",X"30",
		X"04",X"D3",X"09",X"09",X"0A",X"D3",X"59",X"CD",X"63",X"01",X"58",X"CD",X"63",X"07",X"0C",X"CD",
		X"76",X"04",X"C9",X"76",X"08",X"01",X"C9",X"76",X"09",X"1D",X"C9",X"76",X"0A",X"03",X"C9",X"76",
		X"0B",X"F0",X"E9",X"76",X"0F",X"04",X"CA",X"6D",X"DC",X"02",X"01",X"44",X"10",X"00",X"C9",X"4C",
		X"E9",X"4C",X"C2",X"F2",X"3B",X"ED",X"74",X"DC",X"98",X"3B",X"B0",X"82",X"7D",X"33",X"B0",X"82",
		X"61",X"1A",X"6B",X"02",X"23",X"B0",X"82",X"ED",X"7B",X"01",X"02",X"F3",X"0F",X"68",X"FF",X"08",
		X"61",X"02",X"6B",X"04",X"0A",X"6D",X"F6",X"10",X"B4",X"ED",X"76",X"01",X"2B",X"B9",X"82",X"AE",
		X"0C",X"21",X"1A",X"ED",X"7B",X"02",X"FF",X"20",X"25",X"13",X"6B",X"80",X"23",X"B9",X"82",X"7E",
		X"06",X"33",X"33",X"81",X"23",X"37",X"81",X"33",X"3B",X"81",X"23",X"3F",X"81",X"ED",X"7B",X"02",
		X"FF",X"06",X"2D",X"06",X"FF",X"E4",X"88",X"D2",X"3C",X"C8",X"E9",X"76",X"00",X"00",X"E9",X"76",
		X"02",X"F0",X"6B",X"FF",X"23",X"B8",X"82",X"7E",X"E0",X"DD",X"1E",X"3F",X"6B",X"F0",X"8D",X"1E",
		X"3F",X"C8",X"C9",X"70",X"5C",X"81",X"E9",X"70",X"83",X"82",X"17",X"02",X"85",X"ED",X"7B",X"07",
		X"FF",X"04",X"69",X"0C",X"10",X"10",X"00",X"CD",X"18",X"ED",X"18",X"C0",X"14",X"30",X"ED",X"C8",
		X"2B",X"B9",X"82",X"9F",X"7E",X"30",X"25",X"7E",X"01",X"DD",X"21",X"03",X"C9",X"6B",X"0B",X"D3",
		X"08",X"06",X"C9",X"6B",X"0C",X"D3",X"08",X"0E",X"8D",X"C0",X"32",X"E7",X"69",X"09",X"54",X"07",
		X"03",X"DD",X"BB",X"11",X"8D",X"B7",X"3D",X"7E",X"01",X"DD",X"65",X"03",X"C9",X"24",X"06",X"93",
		X"93",X"3D",X"2B",X"22",X"81",X"F3",X"07",X"1F",X"43",X"00",X"74",X"BE",X"3F",X"4C",X"7B",X"CD",
		X"76",X"06",X"C9",X"6B",X"07",X"68",X"F6",X"0F",X"C9",X"37",X"07",X"1F",X"FF",X"05",X"61",X"0A",
		X"C9",X"6B",X"03",X"D3",X"10",X"CD",X"76",X"03",X"0D",X"0C",X"FF",X"0C",X"61",X"08",X"C9",X"6B",
		X"03",X"86",X"10",X"CD",X"76",X"03",X"74",X"C6",X"3F",X"4C",X"7B",X"CD",X"76",X"01",X"3E",X"52",
		X"5E",X"70",X"D6",X"3F",X"18",X"ED",X"CA",X"00",X"46",X"38",X"17",X"CD",X"CA",X"01",X"F6",X"CD",
		X"7B",X"04",X"07",X"C1",X"C9",X"37",X"0C",X"77",X"07",X"CD",X"7B",X"03",X"D0",X"CD",X"76",X"0B",
		X"0D",X"11",X"C9",X"6B",X"04",X"12",X"D0",X"CD",X"76",X"0C",X"72",X"CD",X"7B",X"03",X"07",X"C4",
		X"C9",X"37",X"0B",X"CD",X"21",X"0E",X"C9",X"9F",X"0E",X"56",X"C9",X"76",X"09",X"1D",X"61",X"0A",
		X"C9",X"76",X"09",X"1E",X"54",X"06",X"03",X"DD",X"BB",X"11",X"E9",X"9F",X"00",X"46",X"69",X"04",
		X"C9",X"9F",X"09",X"F6",X"C2",X"E4",X"3C",X"EF",X"23",X"82",X"82",X"3B",X"B9",X"82",X"FF",X"0D",
		X"25",X"1B",X"23",X"33",X"81",X"33",X"37",X"81",X"23",X"3B",X"81",X"33",X"3F",X"81",X"29",X"33",
		X"B9",X"82",X"6B",X"01",X"8D",X"65",X"03",X"7E",X"03",X"DD",X"B8",X"02",X"9D",X"0A",X"09",X"3D",
		X"23",X"33",X"81",X"33",X"37",X"81",X"23",X"3B",X"81",X"33",X"3F",X"81",X"6B",X"08",X"8D",X"B8",
		X"02",X"5D",X"61",X"EB",X"6B",X"80",X"23",X"B9",X"82",X"7E",X"03",X"33",X"82",X"82",X"6B",X"01",
		X"8D",X"65",X"03",X"C8",X"2B",X"B8",X"82",X"AE",X"01",X"30",X"18",X"3B",X"DC",X"80",X"F6",X"03",
		X"FF",X"03",X"61",X"06",X"6B",X"FF",X"23",X"B8",X"82",X"C8",X"8D",X"27",X"3E",X"7E",X"02",X"33",
		X"B8",X"82",X"9D",X"DD",X"44",X"3E",X"9D",X"ED",X"74",X"DC",X"98",X"DD",X"EB",X"3E",X"2B",X"22",
		X"81",X"F3",X"07",X"52",X"12",X"52",X"12",X"ED",X"76",X"03",X"6B",X"08",X"23",X"B0",X"82",X"EF",
		X"23",X"B7",X"82",X"C8",X"E9",X"70",X"DC",X"98",X"E9",X"12",X"02",X"6D",X"FF",X"90",X"25",X"47",
		X"FF",X"40",X"2D",X"43",X"8D",X"83",X"11",X"E7",X"69",X"09",X"E9",X"6B",X"03",X"FD",X"00",X"86",
		X"38",X"09",X"05",X"ED",X"7B",X"03",X"D6",X"40",X"0A",X"3B",X"41",X"81",X"BC",X"56",X"04",X"21",
		X"02",X"56",X"FC",X"5E",X"07",X"3D",X"96",X"0E",X"8D",X"C0",X"32",X"0C",X"61",X"F7",X"4B",X"05",
		X"3D",X"D3",X"04",X"06",X"8D",X"C0",X"32",X"0C",X"61",X"F6",X"2B",X"82",X"82",X"F3",X"0E",X"38",
		X"06",X"50",X"03",X"03",X"8D",X"BB",X"11",X"3B",X"B7",X"82",X"12",X"1F",X"43",X"00",X"74",X"9E",
		X"3F",X"4C",X"7B",X"ED",X"83",X"02",X"E9",X"37",X"02",X"AE",X"F1",X"29",X"1C",X"AE",X"F8",X"21",
		X"18",X"EF",X"E9",X"37",X"00",X"7E",X"01",X"33",X"B8",X"82",X"E9",X"76",X"02",X"F0",X"6B",X"C0",
		X"8D",X"1E",X"3F",X"D3",X"10",X"30",X"F9",X"09",X"21",X"3B",X"B0",X"82",X"7D",X"33",X"B0",X"82",
		X"61",X"18",X"2B",X"B7",X"82",X"68",X"F6",X"07",X"23",X"B7",X"82",X"AE",X"04",X"30",X"06",X"50",
		X"09",X"04",X"8D",X"BB",X"11",X"77",X"7B",X"33",X"B0",X"82",X"9D",X"ED",X"63",X"02",X"F0",X"ED",
		X"63",X"00",X"01",X"DD",X"83",X"11",X"E6",X"7E",X"06",X"30",X"02",X"7E",X"16",X"CD",X"74",X"E4",
		X"88",X"70",X"96",X"3F",X"54",X"04",X"02",X"DD",X"4F",X"35",X"72",X"CD",X"72",X"CD",X"72",X"5D",
		X"61",X"F5",X"14",X"38",X"08",X"CD",X"74",X"D4",X"88",X"0A",X"04",X"09",X"EA",X"C8",X"A5",X"E5",
		X"74",X"00",X"88",X"D0",X"2A",X"7E",X"10",X"76",X"00",X"7C",X"7D",X"30",X"FA",X"B0",X"B5",X"C8",
		X"C7",X"FB",X"00",X"01",X"00",X"01",X"0F",X"02",X"1F",X"02",X"00",X"03",X"1F",X"03",X"0F",X"04",
		X"00",X"04",X"50",X"80",X"C0",X"70",X"90",X"B0",X"60",X"A0",X"02",X"00",X"02",X"08",X"02",X"10",
		X"00",X"02",X"04",X"08",X"0C",X"0E",X"00",X"02",X"00",X"08",X"0C",X"08",X"00",X"04",X"00",X"0A",
		X"0C",X"08",X"28",X"29",X"2A",X"2B",X"6A",X"69",X"01",X"02",X"01",X"01",X"02",X"03",X"01",X"02",
		X"02",X"FE",X"08",X"FF",X"02",X"02",X"08",X"FF",X"01",X"00",X"08",X"FF",X"01",X"00",X"08",X"FF",
		X"01",X"00",X"02",X"01",X"01",X"00",X"02",X"01",X"02",X"FE",X"02",X"01",X"02",X"02",X"02",X"01",
		X"88",X"A8",X"84",X"A4",X"80",X"A0",X"9C",X"BC",X"DC",X"FC",X"9A",X"BA",X"DA",X"FA",X"FF",X"03",
		X"FE",X"05",X"FD",X"07",X"FC",X"01",X"03",X"02",X"02",X"02",X"01",X"02",X"00",X"04",X"96",X"B6",
		X"D6",X"F6",X"67",X"67",X"67",X"67",X"28",X"28",X"30",X"30",X"80",X"80",X"80",X"80",X"01",X"03",
		X"05",X"02",X"01",X"03",X"02",X"01",X"18",X"19",X"1A",X"1B",X"1C",X"9B",X"9A",X"99",X"98",X"99",
		X"9A",X"9B",X"1C",X"1B",X"1A",X"19",X"07",X"F8",X"00",X"F8",X"F8",X"F8",X"F8",X"00",X"F8",X"07",
		X"F8",X"00",X"F8",X"07",X"00",X"07",X"07",X"07",X"00",X"07",X"F8",X"07",X"F8",X"00",X"F8",X"07",
		X"F8",X"00",X"F8",X"F8",X"00",X"F8",X"C7",X"F3",X"41",X"10",X"41",X"10",X"41",X"10",X"41",X"10",
		X"C9",X"2F",X"00",X"80",X"E9",X"70",X"00",X"80",X"17",X"00",X"8D",X"35",X"40",X"CD",X"7F",X"0C",
		X"80",X"ED",X"74",X"0C",X"80",X"02",X"01",X"DD",X"35",X"40",X"C9",X"2F",X"18",X"80",X"E9",X"70",
		X"18",X"80",X"17",X"02",X"8D",X"35",X"40",X"CD",X"7F",X"24",X"80",X"ED",X"74",X"24",X"80",X"02",
		X"03",X"DD",X"35",X"40",X"9D",X"CD",X"7B",X"00",X"FF",X"80",X"9B",X"33",X"42",X"97",X"7E",X"42",
		X"C9",X"6B",X"00",X"AE",X"F8",X"C6",X"0B",X"41",X"3D",X"AE",X"03",X"9B",X"F5",X"41",X"C9",X"6B",
		X"00",X"AE",X"F0",X"30",X"08",X"7E",X"00",X"ED",X"76",X"02",X"C2",X"33",X"42",X"AE",X"F1",X"30",
		X"08",X"7E",X"01",X"ED",X"76",X"02",X"C2",X"33",X"42",X"AE",X"F2",X"30",X"0F",X"6D",X"F7",X"08",
		X"82",X"08",X"C9",X"6B",X"01",X"F3",X"0F",X"C2",X"09",X"97",X"3B",X"42",X"FF",X"F3",X"61",X"27",
		X"3D",X"A6",X"08",X"C2",X"08",X"7E",X"10",X"C2",X"09",X"7E",X"0D",X"C2",X"08",X"CD",X"7B",X"01",
		X"82",X"09",X"6B",X"0C",X"82",X"08",X"C9",X"6B",X"02",X"C2",X"09",X"7E",X"0B",X"C2",X"08",X"CD",
		X"7B",X"03",X"82",X"09",X"C2",X"4B",X"42",X"AE",X"F4",X"93",X"C5",X"43",X"6B",X"07",X"82",X"08",
		X"C9",X"6B",X"01",X"F3",X"80",X"30",X"25",X"6D",X"FF",X"00",X"61",X"08",X"8A",X"0C",X"F6",X"F7",
		X"82",X"09",X"0D",X"3B",X"FF",X"01",X"61",X"08",X"8A",X"0C",X"F6",X"EF",X"82",X"09",X"0D",X"2F",
		X"FF",X"02",X"61",X"21",X"8A",X"0C",X"F6",X"DF",X"82",X"09",X"0D",X"23",X"3D",X"AE",X"00",X"30",
		X"08",X"CA",X"0C",X"A6",X"08",X"C2",X"09",X"09",X"16",X"AE",X"01",X"30",X"08",X"CA",X"0C",X"A6",
		X"10",X"C2",X"09",X"09",X"0A",X"AE",X"02",X"30",X"FC",X"CA",X"0C",X"A6",X"20",X"C2",X"09",X"7E",
		X"06",X"C2",X"08",X"CD",X"7B",X"01",X"82",X"09",X"C2",X"3B",X"42",X"AE",X"F8",X"30",X"08",X"7E",
		X"01",X"33",X"04",X"A0",X"C2",X"33",X"42",X"AE",X"F9",X"30",X"22",X"6D",X"FF",X"03",X"61",X"09",
		X"C9",X"6B",X"01",X"ED",X"76",X"02",X"C2",X"3B",X"42",X"6D",X"F7",X"08",X"82",X"08",X"6B",X"10",
		X"82",X"09",X"6B",X"0D",X"82",X"08",X"6B",X"09",X"82",X"09",X"C2",X"33",X"42",X"AE",X"FA",X"30",
		X"17",X"ED",X"2F",X"00",X"E9",X"32",X"01",X"77",X"72",X"ED",X"65",X"06",X"E9",X"71",X"07",X"CD",
		X"7B",X"01",X"E9",X"37",X"08",X"97",X"3B",X"42",X"FF",X"FB",X"61",X"1B",X"E9",X"6B",X"08",X"2C",
		X"FF",X"FF",X"9B",X"33",X"42",X"ED",X"75",X"08",X"E9",X"3A",X"06",X"ED",X"27",X"07",X"E9",X"25",
		X"00",X"ED",X"24",X"01",X"C2",X"5D",X"42",X"AE",X"FC",X"30",X"17",X"ED",X"2F",X"00",X"E9",X"32",
		X"01",X"77",X"72",X"ED",X"65",X"09",X"E9",X"71",X"0A",X"CD",X"7B",X"01",X"E9",X"37",X"0B",X"97",
		X"3B",X"42",X"FF",X"FD",X"61",X"1B",X"E9",X"6B",X"0B",X"2C",X"FF",X"FF",X"9B",X"33",X"42",X"ED",
		X"75",X"0B",X"E9",X"3A",X"09",X"ED",X"27",X"0A",X"E9",X"25",X"00",X"ED",X"24",X"01",X"C2",X"5D",
		X"42",X"AE",X"FE",X"93",X"C5",X"43",X"6B",X"07",X"82",X"08",X"3D",X"AE",X"00",X"30",X"09",X"CA",
		X"0C",X"A6",X"01",X"C2",X"09",X"97",X"E5",X"41",X"FF",X"01",X"61",X"08",X"8A",X"0C",X"F7",X"02",
		X"82",X"09",X"0D",X"11",X"FF",X"02",X"61",X"08",X"8A",X"0C",X"F7",X"04",X"82",X"09",X"0D",X"05",
		X"6B",X"00",X"23",X"00",X"B0",X"ED",X"2F",X"00",X"E9",X"32",X"01",X"77",X"E9",X"25",X"00",X"ED",
		X"24",X"01",X"C2",X"C5",X"43",X"CD",X"7B",X"00",X"FF",X"F5",X"61",X"0D",X"C9",X"6B",X"01",X"A6",
		X"10",X"ED",X"76",X"0C",X"23",X"00",X"B0",X"09",X"32",X"AE",X"F6",X"30",X"08",X"CD",X"7B",X"01",
		X"23",X"00",X"A8",X"09",X"26",X"AE",X"F7",X"93",X"C5",X"43",X"6B",X"00",X"23",X"04",X"A0",X"7E",
		X"0E",X"C2",X"08",X"CD",X"7B",X"01",X"82",X"09",X"6B",X"0F",X"82",X"08",X"C9",X"6B",X"02",X"C2",
		X"09",X"09",X"10",X"ED",X"2F",X"00",X"E9",X"32",X"01",X"09",X"1B",X"ED",X"2F",X"00",X"E9",X"32",
		X"01",X"09",X"12",X"ED",X"2F",X"00",X"E9",X"32",X"01",X"09",X"09",X"ED",X"2F",X"00",X"E9",X"32",
		X"01",X"09",X"00",X"77",X"72",X"77",X"72",X"ED",X"65",X"00",X"E9",X"71",X"01",X"F5",X"C9",X"E0",
		X"6B",X"80",X"E9",X"37",X"04",X"ED",X"76",X"05",X"C2",X"35",X"40",X"ED",X"2F",X"00",X"E9",X"32",
		X"01",X"77",X"E9",X"25",X"00",X"ED",X"24",X"01",X"A5",X"CD",X"B5",X"97",X"35",X"40",X"F6",X"C0",
		X"FF",X"80",X"61",X"0C",X"C9",X"6B",X"00",X"F3",X"3F",X"A6",X"80",X"ED",X"76",X"05",X"0D",X"DB",
		X"E9",X"24",X"04",X"ED",X"7B",X"04",X"FF",X"80",X"92",X"C5",X"43",X"ED",X"7B",X"03",X"E9",X"37",
		X"04",X"ED",X"7B",X"05",X"FF",X"82",X"9A",X"C2",X"42",X"ED",X"75",X"05",X"3D",X"AE",X"03",X"93",
		X"C5",X"43",X"E9",X"6B",X"05",X"AE",X"82",X"C6",X"C5",X"43",X"6B",X"00",X"23",X"04",X"A0",X"97",
		X"C5",X"43",X"C9",X"6B",X"00",X"AE",X"F0",X"C6",X"40",X"40",X"E9",X"6B",X"02",X"AE",X"00",X"30",
		X"69",X"6D",X"FF",X"00",X"61",X"04",X"6B",X"01",X"0D",X"0E",X"FF",X"01",X"61",X"04",X"6B",X"03",
		X"0D",X"06",X"FF",X"02",X"61",X"2C",X"6B",X"05",X"82",X"08",X"C9",X"6B",X"00",X"C2",X"09",X"09",
		X"00",X"6D",X"FF",X"00",X"61",X"04",X"6B",X"00",X"0D",X"0E",X"FF",X"01",X"61",X"04",X"6B",X"02",
		X"0D",X"06",X"FF",X"02",X"61",X"34",X"6B",X"04",X"82",X"08",X"C9",X"6B",X"01",X"C2",X"09",X"97",
		X"29",X"43",X"6B",X"0E",X"82",X"08",X"C9",X"6B",X"00",X"C2",X"09",X"7E",X"0F",X"C2",X"08",X"7E",
		X"3F",X"C2",X"09",X"CD",X"7B",X"01",X"23",X"00",X"A8",X"ED",X"2F",X"00",X"E9",X"32",X"01",X"77",
		X"72",X"ED",X"65",X"00",X"E9",X"71",X"01",X"97",X"90",X"43",X"C9",X"3A",X"00",X"22",X"00",X"78",
		X"10",X"C8",X"43",X"4C",X"3D",X"AE",X"00",X"30",X"04",X"7E",X"00",X"09",X"0E",X"AE",X"01",X"30",
		X"04",X"7E",X"02",X"09",X"06",X"AE",X"02",X"30",X"27",X"7E",X"04",X"C2",X"08",X"6B",X"82",X"09",
		X"3D",X"AE",X"00",X"30",X"04",X"7E",X"01",X"09",X"0E",X"AE",X"01",X"30",X"04",X"7E",X"03",X"09",
		X"06",X"AE",X"02",X"30",X"0B",X"7E",X"05",X"C2",X"08",X"77",X"7B",X"C2",X"09",X"97",X"83",X"43",
		X"C2",X"12",X"43",X"ED",X"2F",X"00",X"E9",X"32",X"01",X"77",X"E9",X"25",X"00",X"ED",X"24",X"01",
		X"6B",X"07",X"82",X"08",X"3D",X"AE",X"00",X"30",X"06",X"CA",X"0C",X"F3",X"FE",X"09",X"12",X"AE",
		X"01",X"30",X"06",X"CA",X"0C",X"F3",X"FD",X"09",X"08",X"AE",X"02",X"30",X"08",X"CA",X"0C",X"F3",
		X"FB",X"C2",X"09",X"09",X"10",X"ED",X"7B",X"0C",X"F7",X"10",X"E9",X"37",X"0C",X"33",X"00",X"B0",
		X"6B",X"01",X"23",X"04",X"A0",X"C8",X"C7",X"FB",X"5D",X"0D",X"9C",X"0C",X"E7",X"0B",X"3C",X"0B",
		X"9B",X"0A",X"02",X"0A",X"73",X"09",X"EB",X"08",X"6B",X"08",X"F2",X"07",X"80",X"07",X"14",X"07",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AE",X"06",X"4E",X"06",X"F4",X"05",X"9E",X"05",
		X"4D",X"05",X"01",X"05",X"B9",X"04",X"75",X"04",X"35",X"04",X"F9",X"03",X"C0",X"03",X"8A",X"03",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"57",X"03",X"27",X"03",X"FA",X"02",X"CF",X"02",
		X"A7",X"02",X"81",X"02",X"5D",X"02",X"3B",X"02",X"1B",X"02",X"FC",X"01",X"E0",X"01",X"C5",X"01",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AC",X"01",X"94",X"01",X"7D",X"01",X"68",X"01",
		X"53",X"01",X"40",X"01",X"2E",X"01",X"1D",X"01",X"0D",X"01",X"FE",X"00",X"F0",X"00",X"E2",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"D6",X"00",X"CA",X"00",X"BE",X"00",X"B4",X"00",
		X"AA",X"00",X"A0",X"00",X"97",X"00",X"8F",X"00",X"87",X"00",X"7F",X"00",X"78",X"00",X"71",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"6B",X"00",X"65",X"00",X"5F",X"00",X"5A",X"00",
		X"55",X"00",X"50",X"00",X"4C",X"00",X"47",X"00",X"43",X"00",X"40",X"00",X"3C",X"00",X"39",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"35",X"00",X"32",X"00",X"30",X"00",X"2D",X"00",
		X"2A",X"00",X"28",X"00",X"26",X"00",X"24",X"00",X"22",X"00",X"20",X"00",X"1E",X"00",X"1C",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1B",X"00",X"19",X"00",X"18",X"00",X"16",X"00",
		X"15",X"00",X"14",X"00",X"13",X"00",X"12",X"00",X"11",X"00",X"10",X"00",X"0F",X"00",X"0E",X"00",
		X"08",X"08",X"00",X"02",X"05",X"10",X"01",X"00",X"18",X"04",X"00",X"00",X"00",X"00",X"01",X"01",
		X"09",X"06",X"02",X"00",X"80",X"84",X"00",X"01",X"00",X"00",X"18",X"08",X"01",X"05",X"05",X"00",
		X"09",X"00",X"00",X"02",X"00",X"0D",X"00",X"00",X"08",X"06",X"0C",X"00",X"01",X"04",X"08",X"00",
		X"48",X"00",X"04",X"00",X"02",X"84",X"25",X"00",X"04",X"00",X"00",X"05",X"0E",X"06",X"00",X"01",
		X"A0",X"F2",X"0D",X"FA",X"01",X"50",X"8A",X"FE",X"82",X"50",X"83",X"FE",X"81",X"50",X"8A",X"FE",
		X"82",X"4A",X"83",X"FE",X"81",X"50",X"8A",X"FE",X"82",X"50",X"83",X"FE",X"81",X"53",X"8A",X"FE",
		X"82",X"50",X"83",X"FE",X"81",X"50",X"8A",X"FE",X"82",X"4A",X"83",X"FE",X"81",X"47",X"8A",X"FE",
		X"82",X"45",X"83",X"FE",X"01",X"47",X"90",X"FE",X"90",X"45",X"8A",X"FE",X"82",X"43",X"83",X"FE",
		X"81",X"45",X"8A",X"FE",X"82",X"43",X"83",X"FE",X"81",X"45",X"8A",X"FE",X"82",X"43",X"83",X"FE",
		X"81",X"45",X"8A",X"FE",X"82",X"47",X"83",X"FE",X"81",X"4A",X"8A",X"FE",X"82",X"47",X"83",X"FE",
		X"81",X"4A",X"8A",X"FE",X"82",X"53",X"84",X"50",X"94",X"FE",X"88",X"4A",X"84",X"50",X"88",X"FE",
		X"84",X"4A",X"84",X"50",X"88",X"FE",X"84",X"4A",X"84",X"50",X"98",X"FE",X"98",X"FB",X"FE",X"FF",
		X"A0",X"FE",X"F3",X"09",X"20",X"00",X"FA",X"01",X"30",X"F9",X"9C",X"2A",X"F9",X"84",X"30",X"F9",
		X"A0",X"27",X"F9",X"9C",X"25",X"F9",X"84",X"27",X"F9",X"A0",X"25",X"F9",X"9C",X"23",X"F9",X"84",
		X"25",X"F9",X"A0",X"27",X"F9",X"9C",X"2A",X"F9",X"84",X"30",X"F9",X"A0",X"30",X"F9",X"90",X"30",
		X"F9",X"90",X"30",X"F9",X"B0",X"FB",X"FE",X"FF",X"A0",X"27",X"F3",X"09",X"20",X"00",X"9C",X"2A",
		X"F3",X"09",X"20",X"00",X"84",X"30",X"F3",X"09",X"20",X"00",X"A0",X"30",X"F3",X"09",X"20",X"00",
		X"90",X"30",X"F3",X"09",X"20",X"00",X"90",X"30",X"F3",X"09",X"20",X"00",X"B0",X"FB",X"FE",X"FF",
		X"FE",X"FF",X"F2",X"0C",X"FA",X"01",X"FE",X"82",X"2B",X"84",X"FE",X"84",X"27",X"84",X"FE",X"84",
		X"30",X"84",X"FE",X"84",X"30",X"84",X"FE",X"84",X"30",X"84",X"27",X"82",X"1B",X"84",X"22",X"82",
		X"1B",X"84",X"20",X"84",X"FE",X"84",X"FB",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"F5",X"0E",X"F6",X"80",X"F7",X"80",X"BF",X"82",X"F8",X"9E",X"FC",X"01",X"F5",X"0E",X"F6",
		X"C0",X"FA",X"06",X"8E",X"F7",X"70",X"7F",X"82",X"F8",X"94",X"FB",X"98",X"FA",X"02",X"F7",X"F8",
		X"FF",X"82",X"F8",X"92",X"FB",X"9E",X"FD",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"F1",X"F3",X"09",X"80",X"00",X"6B",X"6A",X"69",X"68",X"67",X"66",X"65",X"64",X"63",X"62",
		X"61",X"60",X"5B",X"5A",X"59",X"58",X"57",X"56",X"55",X"54",X"53",X"52",X"51",X"50",X"4B",X"4A",
		X"49",X"48",X"47",X"46",X"45",X"43",X"42",X"41",X"40",X"3B",X"3A",X"39",X"38",X"37",X"36",X"35",
		X"34",X"32",X"31",X"30",X"2B",X"2A",X"29",X"28",X"27",X"26",X"25",X"24",X"23",X"22",X"21",X"20",
		X"1B",X"1A",X"19",X"18",X"17",X"16",X"15",X"14",X"13",X"12",X"11",X"10",X"FE",X"FF",X"00",X"00",
		X"80",X"F1",X"F3",X"09",X"80",X"00",X"69",X"68",X"67",X"66",X"65",X"64",X"63",X"62",X"61",X"60",
		X"5B",X"5A",X"59",X"58",X"57",X"56",X"55",X"54",X"53",X"52",X"51",X"50",X"4B",X"4A",X"49",X"48",
		X"47",X"46",X"45",X"43",X"42",X"41",X"40",X"3B",X"3A",X"39",X"38",X"37",X"36",X"35",X"34",X"33",
		X"32",X"31",X"30",X"2B",X"2A",X"29",X"28",X"27",X"26",X"25",X"24",X"23",X"22",X"21",X"20",X"1B",
		X"1A",X"19",X"18",X"17",X"16",X"15",X"14",X"13",X"12",X"11",X"10",X"F2",X"00",X"FE",X"FF",X"00",
		X"80",X"F1",X"F2",X"0C",X"FC",X"01",X"FA",X"07",X"59",X"66",X"52",X"59",X"66",X"59",X"56",X"62",
		X"69",X"62",X"57",X"62",X"6B",X"62",X"5B",X"67",X"51",X"57",X"64",X"57",X"54",X"61",X"67",X"61",
		X"56",X"61",X"69",X"61",X"FB",X"F3",X"09",X"FF",X"FF",X"FD",X"FE",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"80",X"F4",X"FF",X"F1",X"F2",X"0C",X"FA",X"00",X"40",X"84",X"FE",X"81",X"44",X"81",X"FE",X"81",
		X"47",X"84",X"FE",X"81",X"50",X"83",X"53",X"81",X"54",X"83",X"FE",X"81",X"52",X"83",X"FE",X"81",
		X"50",X"83",X"FE",X"81",X"49",X"83",X"FE",X"81",X"46",X"90",X"47",X"82",X"FE",X"8E",X"FB",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"F4",X"FF",X"F1",X"F2",X"0C",X"FA",X"02",X"27",X"88",X"2A",X"84",X"2B",X"84",X"FB",X"FE",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"F4",X"FF",X"F1",X"FA",X"01",X"F3",X"09",X"30",X"00",X"22",X"90",X"F3",X"09",X"30",X"00",
		X"17",X"90",X"FB",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"F5",X"0E",X"F6",X"B0",X"FA",X"03",X"F7",X"F8",X"FF",X"82",X"F8",X"88",X"F7",X"70",X"7F",
		X"82",X"F8",X"88",X"FB",X"F6",X"50",X"FA",X"03",X"A0",X"F7",X"00",X"3F",X"82",X"F8",X"FB",X"FF",
		X"80",X"F5",X"0C",X"F6",X"90",X"F7",X"B8",X"BF",X"82",X"F8",X"B8",X"F5",X"0E",X"B0",X"F6",X"70",
		X"B0",X"F7",X"00",X"3F",X"82",X"F8",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"F5",X"0C",X"F6",X"70",X"F7",X"B8",X"BF",X"82",X"F8",X"B0",X"F5",X"0E",X"B0",X"F6",X"60",
		X"B0",X"F7",X"00",X"3F",X"82",X"F8",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"F5",X"0E",X"F6",X"90",X"F7",X"F8",X"FF",X"82",X"F8",X"88",X"F5",X"0F",X"F6",X"90",X"F7",
		X"40",X"7F",X"82",X"F8",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"82",X"FA",X"00",X"F1",X"F2",X"0C",X"45",X"83",X"FE",X"81",X"47",X"82",X"45",X"82",X"47",
		X"83",X"FE",X"81",X"48",X"83",X"FE",X"81",X"50",X"83",X"FE",X"81",X"51",X"82",X"50",X"82",X"48",
		X"83",X"FE",X"81",X"50",X"83",X"FE",X"81",X"51",X"81",X"FE",X"81",X"55",X"81",X"FE",X"81",X"55",
		X"82",X"58",X"82",X"57",X"82",X"55",X"82",X"51",X"83",X"FE",X"81",X"50",X"90",X"FB",X"FE",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"82",X"F1",X"F2",X"0C",X"FE",X"90",X"FA",X"00",X"55",X"83",X"FE",X"81",X"57",X"82",X"55",
		X"82",X"57",X"83",X"FE",X"81",X"58",X"83",X"FE",X"81",X"60",X"83",X"FE",X"81",X"61",X"82",X"60",
		X"82",X"58",X"83",X"FE",X"81",X"60",X"83",X"FE",X"81",X"61",X"81",X"FE",X"81",X"65",X"81",X"FE",
		X"81",X"65",X"82",X"68",X"82",X"67",X"82",X"65",X"82",X"61",X"83",X"FE",X"81",X"60",X"90",X"FB",
		X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"82",X"F1",X"F2",X"0C",X"FE",X"A0",X"FA",X"00",X"25",X"83",X"FE",X"81",X"27",X"82",X"25",
		X"82",X"27",X"83",X"FE",X"81",X"28",X"83",X"FE",X"81",X"30",X"83",X"FE",X"81",X"31",X"82",X"30",
		X"82",X"28",X"83",X"FE",X"81",X"30",X"83",X"FE",X"81",X"31",X"81",X"FE",X"81",X"35",X"81",X"FE",
		X"81",X"35",X"82",X"38",X"82",X"37",X"82",X"35",X"82",X"31",X"83",X"FE",X"81",X"30",X"87",X"FE",
		X"81",X"30",X"82",X"2A",X"82",X"28",X"82",X"27",X"82",X"FB",X"F3",X"09",X"20",X"00",X"25",X"90",
		X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"F5",X"0E",X"F6",X"B0",X"FA",X"0A",X"F7",X"30",X"3F",X"82",X"F8",X"84",X"F7",X"30",X"3F",
		X"82",X"F8",X"82",X"F7",X"30",X"3F",X"82",X"F8",X"88",X"FB",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"80",X"F5",X"0E",X"F6",X"B0",X"F7",X"30",X"3F",X"82",X"F8",X"88",X"F6",X"B4",X"F7",X"28",X"3F",
		X"82",X"F8",X"90",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"F1",X"F2",X"0C",X"FA",X"02",X"43",X"83",X"FE",X"81",X"F3",X"09",X"20",X"00",X"44",X"8C",
		X"F2",X"0C",X"46",X"83",X"FE",X"81",X"F3",X"09",X"20",X"00",X"47",X"8C",X"F2",X"0C",X"43",X"83",
		X"FE",X"81",X"44",X"83",X"FE",X"82",X"46",X"83",X"FE",X"81",X"47",X"83",X"FE",X"82",X"50",X"83",
		X"FE",X"81",X"4B",X"87",X"FE",X"81",X"4A",X"84",X"FE",X"81",X"FB",X"FF",X"00",X"00",X"00",X"00",
		X"80",X"F1",X"F3",X"09",X"20",X"00",X"FA",X"02",X"2A",X"F9",X"84",X"2B",X"F9",X"8C",X"21",X"F9",
		X"84",X"22",X"F9",X"8C",X"2A",X"F9",X"84",X"2B",X"F9",X"84",X"21",X"F9",X"84",X"22",X"F9",X"85",
		X"27",X"F9",X"84",X"26",X"F9",X"88",X"2A",X"F9",X"86",X"FB",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"F1",X"F2",X"0C",X"FA",X"02",X"33",X"83",X"FE",X"81",X"34",X"88",X"FE",X"84",X"36",X"83",
		X"FE",X"81",X"37",X"88",X"FE",X"84",X"33",X"83",X"FE",X"81",X"34",X"83",X"FE",X"81",X"36",X"83",
		X"FE",X"81",X"37",X"83",X"FE",X"82",X"40",X"83",X"FE",X"81",X"3B",X"87",X"FE",X"81",X"3A",X"84",
		X"FE",X"82",X"FB",X"FF",X"80",X"F5",X"0E",X"F6",X"60",X"F7",X"30",X"3F",X"82",X"F8",X"A0",X"FF",
		X"80",X"FE",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"F1",X"F2",X"0C",X"FE",X"80",X"FA",X"FF",X"21",X"82",X"1A",X"81",X"18",X"81",X"21",X"81",
		X"FE",X"81",X"1A",X"81",X"18",X"81",X"FB",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"8C",X"F1",X"F2",X"0C",X"FC",X"01",X"FA",X"01",X"45",X"83",X"FE",X"81",X"45",X"83",X"FE",
		X"81",X"45",X"83",X"FE",X"81",X"45",X"83",X"FE",X"81",X"45",X"82",X"44",X"82",X"45",X"83",X"FE",
		X"81",X"46",X"83",X"FE",X"81",X"45",X"83",X"FE",X"81",X"FB",X"FA",X"01",X"46",X"82",X"45",X"82",
		X"46",X"83",X"FE",X"81",X"47",X"83",X"FE",X"81",X"48",X"83",X"FE",X"81",X"FB",X"51",X"88",X"FE",
		X"88",X"FD",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"8C",X"F1",X"F2",X"0C",X"FC",X"01",X"FA",X"03",X"21",X"84",X"1A",X"82",X"18",X"82",X"21",
		X"83",X"FE",X"81",X"1A",X"82",X"18",X"82",X"FB",X"FA",X"01",X"26",X"82",X"25",X"82",X"26",X"83",
		X"FE",X"81",X"27",X"83",X"FE",X"81",X"28",X"83",X"FE",X"81",X"FB",X"31",X"88",X"FE",X"82",X"FE",
		X"82",X"FE",X"82",X"FE",X"82",X"FD",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"8C",X"F1",X"FC",X"01",X"FA",X"03",X"F3",X"09",X"20",X"00",X"21",X"90",X"FB",X"FA",X"03",
		X"FE",X"90",X"FB",X"FD",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"F5",X"0E",X"F6",X"80",X"F7",X"80",X"BF",X"82",X"F8",X"F8",X"92",X"F5",X"0E",X"F6",X"C0",
		X"FA",X"0D",X"F7",X"F8",X"FF",X"82",X"F8",X"88",X"F7",X"70",X"7F",X"82",X"F8",X"88",X"FB",X"FF",
		X"88",X"F1",X"F2",X"0E",X"FA",X"02",X"FE",X"82",X"42",X"82",X"43",X"82",X"44",X"82",X"50",X"84",
		X"44",X"82",X"50",X"84",X"44",X"82",X"50",X"87",X"FE",X"81",X"50",X"82",X"52",X"82",X"53",X"82",
		X"54",X"82",X"50",X"82",X"52",X"82",X"54",X"84",X"4B",X"82",X"52",X"84",X"50",X"84",X"FE",X"84",
		X"FB",X"FF",X"90",X"FB",X"FD",X"FF",X"00",X"00",X"88",X"F1",X"F1",X"F2",X"0E",X"FA",X"02",X"FE",
		X"82",X"27",X"84",X"30",X"84",X"34",X"84",X"30",X"84",X"37",X"84",X"35",X"84",X"39",X"84",X"30",
		X"84",X"34",X"84",X"37",X"82",X"2B",X"84",X"32",X"82",X"2B",X"84",X"30",X"84",X"FE",X"84",X"FB",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"F1",X"F2",X"08",X"FA",X"02",X"FE",X"82",
		X"2B",X"84",X"FE",X"84",X"27",X"84",X"FE",X"84",X"30",X"84",X"FE",X"84",X"30",X"84",X"FE",X"84",
		X"30",X"84",X"27",X"82",X"1B",X"84",X"22",X"82",X"1B",X"84",X"20",X"84",X"FE",X"84",X"FB",X"FF",
		X"80",X"F5",X"0E",X"F6",X"80",X"FA",X"00",X"F7",X"80",X"BF",X"82",X"F8",X"FB",X"FF",X"00",X"00",
		X"88",X"F1",X"F2",X"0C",X"FE",X"82",X"FA",X"01",X"40",X"82",X"3B",X"82",X"39",X"82",X"37",X"82",
		X"FB",X"F3",X"09",X"20",X"00",X"40",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"F1",X"F2",X"0C",X"FE",X"86",X"FA",X"01",X"39",X"82",X"37",X"82",X"35",X"82",X"34",X"82",
		X"FB",X"F3",X"09",X"20",X"00",X"39",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"F1",X"F2",X"0C",X"FE",X"8A",X"FA",X"01",X"35",X"82",X"34",X"82",X"32",X"82",X"30",X"82",
		X"FB",X"F3",X"09",X"20",X"00",X"35",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"84",X"F5",X"0E",X"F6",X"50",X"F7",X"C0",X"FF",X"82",X"F8",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"80",X"F5",X"0E",X"F6",X"00",X"F7",X"70",X"7F",X"82",X"F8",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"80",X"F1",X"F2",X"0C",X"FC",X"01",X"FA",X"01",X"34",X"38",X"3B",X"44",X"2B",X"33",X"36",X"3B",
		X"31",X"34",X"38",X"41",X"28",X"2B",X"33",X"38",X"29",X"31",X"34",X"39",X"21",X"24",X"28",X"34",
		X"26",X"29",X"34",X"39",X"2B",X"33",X"36",X"3B",X"FB",X"F3",X"09",X"FF",X"FF",X"FD",X"FE",X"FF",
		X"80",X"F1",X"F2",X"0C",X"FC",X"01",X"FA",X"01",X"21",X"84",X"18",X"84",X"19",X"84",X"14",X"84",
		X"16",X"84",X"11",X"84",X"16",X"84",X"18",X"84",X"FB",X"F3",X"09",X"FF",X"FF",X"FD",X"FE",X"FF",
		X"81",X"F1",X"F2",X"0C",X"FA",X"01",X"39",X"84",X"FE",X"82",X"42",X"FE",X"42",X"84",X"FE",X"82",
		X"46",X"FE",X"4B",X"84",X"FE",X"82",X"46",X"FE",X"49",X"84",X"FE",X"82",X"FE",X"82",X"49",X"84",
		X"FE",X"82",X"4B",X"FE",X"49",X"84",X"FE",X"82",X"46",X"FE",X"47",X"84",X"FE",X"82",X"46",X"FE",
		X"44",X"84",X"FE",X"82",X"FE",X"82",X"3B",X"84",X"FE",X"82",X"44",X"FE",X"44",X"84",X"FE",X"82",
		X"47",X"FE",X"51",X"84",X"FE",X"82",X"51",X"FE",X"4B",X"84",X"FE",X"82",X"49",X"FE",X"47",X"84",
		X"FE",X"82",X"47",X"FE",X"46",X"84",X"FE",X"82",X"44",X"FE",X"41",X"86",X"FE",X"82",X"44",X"86",
		X"FE",X"82",X"42",X"8E",X"FE",X"82",X"FB",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"81",X"F1",X"F2",X"0C",X"FA",X"01",X"39",X"84",X"FE",X"82",X"36",X"84",X"FE",X"84",X"32",X"84",
		X"FE",X"84",X"32",X"84",X"FE",X"84",X"36",X"FE",X"39",X"84",X"FE",X"82",X"36",X"84",X"FE",X"84",
		X"32",X"84",X"FE",X"84",X"31",X"84",X"FE",X"84",X"31",X"FE",X"37",X"84",X"FE",X"82",X"2B",X"84",
		X"FE",X"84",X"2B",X"84",X"FE",X"84",X"31",X"84",X"FE",X"84",X"31",X"84",X"FE",X"84",X"34",X"84",
		X"FE",X"84",X"28",X"84",X"FE",X"84",X"31",X"84",X"FE",X"84",X"31",X"FE",X"36",X"8E",X"FE",X"82",
		X"FB",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"F1",X"FE",X"F3",X"09",X"20",X"00",X"FA",
		X"01",X"1B",X"F9",X"88",X"19",X"F9",X"88",X"17",X"F9",X"88",X"16",X"F9",X"88",X"1B",X"F9",X"88",
		X"16",X"F9",X"88",X"21",X"F9",X"88",X"16",X"F9",X"88",X"21",X"F9",X"88",X"11",X"F9",X"88",X"16",
		X"F9",X"88",X"16",X"F9",X"88",X"21",X"F9",X"88",X"11",X"F9",X"88",X"16",X"F9",X"88",X"16",X"F9",
		X"88",X"1B",X"F9",X"88",X"0B",X"F9",X"88",X"FB",X"12",X"F9",X"88",X"FE",X"FF",X"00",X"00",X"00",
		X"80",X"F5",X"0F",X"F6",X"F0",X"FA",X"02",X"F7",X"70",X"7F",X"82",X"F8",X"84",X"FB",X"FF",X"00",
		X"80",X"F5",X"0F",X"F6",X"A0",X"F7",X"30",X"3F",X"82",X"F8",X"88",X"FE",X"FF",X"00",X"00",X"00",
		X"80",X"F1",X"F2",X"0C",X"FA",X"01",X"FE",X"32",X"36",X"3B",X"39",X"36",X"42",X"32",X"36",X"41",
		X"32",X"36",X"3B",X"32",X"36",X"39",X"32",X"36",X"39",X"2B",X"34",X"37",X"2B",X"36",X"37",X"2B",
		X"34",X"2B",X"34",X"37",X"FE",X"31",X"34",X"39",X"37",X"34",X"41",X"31",X"34",X"3B",X"31",X"34",
		X"39",X"31",X"34",X"37",X"31",X"34",X"37",X"29",X"32",X"36",X"29",X"35",X"36",X"29",X"32",X"29",
		X"FE",X"FE",X"FB",X"FF",X"00",X"00",X"00",X"00",X"80",X"F1",X"F2",X"0C",X"FA",X"01",X"FE",X"86",
		X"26",X"83",X"29",X"83",X"26",X"83",X"29",X"83",X"1B",X"83",X"27",X"83",X"17",X"86",X"21",X"84",
		X"FE",X"82",X"21",X"83",X"27",X"83",X"21",X"83",X"27",X"83",X"26",X"83",X"21",X"83",X"26",X"83",
		X"29",X"2B",X"31",X"FB",X"FE",X"FF",X"F9",X"82",X"32",X"F9",X"82",X"2B",X"F9",X"82",X"37",X"F9",
		X"84",X"21",X"F9",X"82",X"27",X"F9",X"82",X"34",X"F9",X"82",X"27",X"F9",X"82",X"24",X"F9",X"82",
		X"31",X"F9",X"82",X"37",X"F9",X"82",X"31",X"F9",X"82",X"26",X"F9",X"82",X"31",X"F9",X"82",X"39",
		X"F9",X"82",X"31",X"F9",X"82",X"FB",X"FF",X"00",X"80",X"F1",X"F2",X"08",X"FA",X"01",X"FE",X"8C",
		X"31",X"83",X"FE",X"83",X"31",X"83",X"FE",X"83",X"2B",X"83",X"FE",X"86",X"FE",X"86",X"2B",X"83",
		X"FE",X"83",X"2B",X"83",X"FE",X"8C",X"FB",X"FE",X"FF",X"39",X"F9",X"82",X"32",X"F9",X"82",X"27",
		X"F9",X"82",X"32",X"F9",X"82",X"3B",X"F9",X"82",X"32",X"F9",X"82",X"2B",X"F9",X"82",X"37",X"F9",
		X"84",X"21",X"F9",X"82",X"27",X"F9",X"82",X"34",X"F9",X"82",X"27",X"F9",X"82",X"24",X"F9",X"82",
		X"31",X"F9",X"82",X"37",X"F9",X"82",X"31",X"F9",X"82",X"26",X"F9",X"82",X"31",X"F9",X"82",X"39",
		X"F9",X"82",X"31",X"F9",X"82",X"FB",X"FF",X"00",X"80",X"F5",X"0E",X"F6",X"80",X"F7",X"80",X"BF",
		X"82",X"F8",X"FF",X"00",X"00",X"00",X"00",X"00",X"80",X"F1",X"F3",X"09",X"30",X"00",X"20",X"FF",
		X"80",X"F1",X"F3",X"09",X"30",X"00",X"22",X"FF",X"80",X"F1",X"F3",X"09",X"30",X"00",X"24",X"FF",
		X"80",X"F5",X"0E",X"F6",X"00",X"F7",X"70",X"7F",X"82",X"F8",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"80",X"F1",X"FA",X"07",X"F3",X"09",X"10",X"00",X"60",X"90",X"FB",X"FF",X"00",X"00",X"00",X"00",
		X"80",X"F1",X"FA",X"07",X"F3",X"09",X"10",X"00",X"62",X"90",X"FB",X"FF",X"00",X"00",X"C7",X"F3");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
