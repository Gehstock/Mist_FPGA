library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity spchip_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of spchip_rom is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"01",X"03",X"07",X"03",X"01",X"00",X"70",X"10",X"30",X"70",X"0F",X"70",X"30",
		X"00",X"B0",X"80",X"F0",X"FE",X"FF",X"F1",X"F1",X"00",X"C0",X"C0",X"C0",X"80",X"0E",X"C8",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"AA",X"AA",X"F0",X"30",X"00",X"00",X"00",
		X"FE",X"FF",X"FF",X"F0",X"F0",X"F0",X"E0",X"00",X"E0",X"E0",X"E0",X"E0",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"07",X"03",X"01",X"00",X"10",X"00",X"00",X"10",X"0F",X"10",X"30",
		X"00",X"E0",X"60",X"F0",X"FE",X"FF",X"F1",X"F1",X"00",X"00",X"00",X"80",X"C0",X"0E",X"C8",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"AA",X"AA",X"F0",X"30",X"00",X"00",X"00",
		X"FE",X"FF",X"FF",X"F0",X"F0",X"F0",X"E0",X"00",X"E0",X"E0",X"E0",X"E0",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"E6",X"91",X"F7",X"91",
		X"00",X"02",X"07",X"0F",X"02",X"52",X"D2",X"D2",X"00",X"00",X"00",X"08",X"00",X"20",X"A0",X"E0",
		X"70",X"70",X"70",X"30",X"30",X"10",X"00",X"00",X"F7",X"F7",X"F7",X"F6",X"F0",X"F0",X"F0",X"00",
		X"F3",X"F3",X"F3",X"FE",X"DE",X"42",X"02",X"00",X"E0",X"80",X"A0",X"A0",X"E0",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"E6",X"91",X"F7",X"91",
		X"00",X"02",X"07",X"0F",X"02",X"02",X"82",X"D2",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"20",
		X"70",X"70",X"70",X"30",X"30",X"10",X"00",X"00",X"F7",X"F7",X"F7",X"F6",X"F0",X"F0",X"F0",X"00",
		X"F3",X"F3",X"F3",X"FE",X"DE",X"52",X"02",X"00",X"A0",X"E0",X"E0",X"80",X"80",X"00",X"00",X"00",
		X"00",X"10",X"00",X"00",X"00",X"33",X"77",X"66",X"00",X"C0",X"E0",X"70",X"F0",X"F0",X"F0",X"70",
		X"00",X"00",X"30",X"F3",X"F3",X"F0",X"F1",X"F3",X"00",X"40",X"C0",X"C0",X"C8",X"CC",X"CC",X"88",
		X"00",X"11",X"11",X"10",X"00",X"00",X"00",X"00",X"FF",X"55",X"55",X"F0",X"70",X"10",X"10",X"00",
		X"FC",X"FE",X"FE",X"F0",X"F0",X"F0",X"C0",X"00",X"C0",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"30",X"00",X"30",X"F8",X"F8",X"F8",X"30",
		X"00",X"E0",X"E0",X"F0",X"FE",X"FF",X"FD",X"F1",X"00",X"00",X"00",X"80",X"C0",X"C0",X"C8",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"AA",X"AA",X"F0",X"30",X"00",X"00",X"00",
		X"FE",X"FF",X"FF",X"F0",X"F0",X"F0",X"E0",X"00",X"E0",X"E0",X"E0",X"E0",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"70",X"00",X"00",X"00",X"E6",X"91",X"F7",X"91",X"F7",
		X"00",X"CC",X"EE",X"66",X"70",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"20",X"60",X"E0",X"C0",X"80",
		X"70",X"70",X"30",X"30",X"10",X"00",X"00",X"00",X"F7",X"F7",X"F6",X"F0",X"F0",X"F0",X"00",X"00",
		X"F0",X"F0",X"F9",X"FD",X"FF",X"76",X"00",X"00",X"80",X"80",X"C8",X"C8",X"C0",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"E6",X"91",X"F7",X"91",
		X"00",X"00",X"00",X"22",X"77",X"70",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"A0",
		X"70",X"70",X"70",X"30",X"30",X"10",X"00",X"00",X"F7",X"F7",X"F7",X"F6",X"F0",X"F0",X"F0",X"00",
		X"F7",X"F7",X"F3",X"FE",X"FC",X"70",X"00",X"00",X"E0",X"E0",X"E0",X"80",X"80",X"00",X"00",X"00",
		X"00",X"01",X"03",X"06",X"0C",X"08",X"33",X"33",X"00",X"0F",X"0E",X"1E",X"34",X"34",X"0F",X"F8",
		X"00",X"30",X"10",X"F0",X"F0",X"FE",X"FF",X"F0",X"00",X"E0",X"C0",X"E0",X"E0",X"F0",X"FC",X"EC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"55",X"55",X"70",X"10",X"00",X"00",X"00",
		X"FF",X"77",X"77",X"F0",X"F0",X"70",X"70",X"00",X"F0",X"F8",X"F8",X"F0",X"E0",X"C0",X"00",X"00",
		X"00",X"01",X"03",X"16",X"3C",X"3B",X"33",X"00",X"00",X"0F",X"1E",X"1E",X"B4",X"0F",X"F0",X"FF",
		X"00",X"70",X"10",X"F0",X"FE",X"FF",X"F0",X"FC",X"00",X"80",X"C0",X"E0",X"E0",X"EC",X"EC",X"C0",
		X"11",X"11",X"10",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"F0",X"70",X"10",X"10",X"00",X"00",
		X"FE",X"FE",X"F0",X"F0",X"F0",X"C0",X"00",X"00",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"E6",X"91",X"F7",
		X"03",X"01",X"CC",X"CC",X"8C",X"87",X"B4",X"B4",X"00",X"08",X"0C",X"06",X"0E",X"0E",X"0E",X"82",
		X"10",X"70",X"70",X"70",X"30",X"30",X"10",X"00",X"91",X"F7",X"F7",X"F7",X"F6",X"F0",X"F0",X"F0",
		X"F6",X"F6",X"F6",X"F4",X"FC",X"FC",X"F0",X"60",X"80",X"80",X"A0",X"E0",X"E0",X"E0",X"A0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"73",X"40",X"F3",X"C0",X"F3",
		X"03",X"01",X"76",X"76",X"DA",X"CB",X"DA",X"DA",X"00",X"08",X"0C",X"86",X"0E",X"0E",X"0E",X"C2",
		X"30",X"30",X"10",X"10",X"00",X"00",X"00",X"00",X"F3",X"F3",X"F3",X"F0",X"F0",X"70",X"00",X"00",
		X"FB",X"FB",X"F3",X"F2",X"F6",X"F6",X"70",X"00",X"80",X"A0",X"A0",X"E0",X"E0",X"C0",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"00",X"00",X"00",X"00",X"11",X"77",X"00",X"E0",X"E0",X"70",X"10",X"74",X"FC",X"33",
		X"00",X"00",X"00",X"F0",X"F3",X"F3",X"F0",X"FF",X"00",X"30",X"70",X"F0",X"FC",X"EE",X"E6",X"F4",
		X"EE",X"FF",X"66",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"70",X"10",X"00",X"00",X"00",X"00",
		X"77",X"77",X"F0",X"F0",X"70",X"70",X"00",X"00",X"F8",X"F8",X"F0",X"E0",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"77",X"77",X"22",X"00",X"73",X"40",X"F3",
		X"00",X"88",X"88",X"CC",X"44",X"66",X"E8",X"F8",X"00",X"00",X"00",X"20",X"60",X"E0",X"E0",X"80",
		X"00",X"30",X"30",X"30",X"10",X"10",X"00",X"00",X"C0",X"F3",X"F3",X"F3",X"F3",X"F0",X"F0",X"70",
		X"F8",X"F8",X"FB",X"FB",X"F3",X"FF",X"F6",X"90",X"80",X"80",X"80",X"80",X"80",X"C0",X"E0",X"E0",
		X"00",X"00",X"00",X"03",X"07",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"0C",X"0E",X"0F",X"0F",X"0F",
		X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"03",X"03",X"03",X"03",
		X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"08",X"08",X"08",X"08",X"08",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"03",X"03",X"03",X"01",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0E",X"08",X"08",X"08",X"08",X"08",X"08",X"00",X"00",
		X"00",X"00",X"00",X"40",X"E0",X"B0",X"B0",X"10",X"10",X"70",X"00",X"30",X"F0",X"F0",X"F0",X"F0",
		X"C0",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F1",X"00",X"00",X"00",X"00",X"33",X"77",X"22",X"EE",
		X"10",X"11",X"11",X"55",X"FF",X"EE",X"00",X"00",X"F0",X"F0",X"55",X"00",X"55",X"70",X"00",X"00",
		X"F0",X"F0",X"DD",X"88",X"DD",X"F0",X"F0",X"30",X"EC",X"F0",X"F8",X"FC",X"FC",X"E0",X"C0",X"80",
		X"40",X"40",X"70",X"70",X"10",X"10",X"70",X"F0",X"00",X"00",X"80",X"C0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"11",X"00",X"F0",X"F1",X"F0",X"00",X"00",X"CC",X"EE",X"44",X"CC",X"CC",X"88",
		X"B0",X"B0",X"10",X"77",X"66",X"00",X"00",X"00",X"F0",X"F0",X"F3",X"66",X"44",X"33",X"30",X"00",
		X"F7",X"DD",X"99",X"DD",X"76",X"F8",X"F0",X"30",X"F0",X"F8",X"F8",X"F0",X"E0",X"E0",X"E0",X"C0",
		X"00",X"30",X"70",X"70",X"C0",X"80",X"30",X"30",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"30",
		X"C0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F3",X"DD",X"33",X"77",X"33",X"E6",X"CC",X"CC",X"F0",X"FC",
		X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"66",X"44",X"22",X"30",X"00",X"00",X"00",
		X"88",X"DD",X"77",X"FC",X"F0",X"70",X"00",X"00",X"FC",X"FC",X"E0",X"E0",X"E0",X"00",X"00",X"00",
		X"00",X"10",X"00",X"00",X"00",X"30",X"00",X"00",X"10",X"10",X"90",X"40",X"00",X"80",X"00",X"40",
		X"00",X"10",X"20",X"40",X"00",X"30",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",
		X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"10",X"10",X"00",X"00",X"00",X"00",X"00",
		X"20",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"11",X"00",X"31",X"20",X"31",X"00",X"88",X"00",X"FE",X"30",X"74",X"30",X"74",
		X"70",X"10",X"70",X"E0",X"F0",X"F0",X"F0",X"F0",X"00",X"80",X"00",X"00",X"00",X"20",X"A0",X"B0",
		X"71",X"71",X"E0",X"F1",X"F1",X"71",X"30",X"10",X"FC",X"74",X"30",X"74",X"FD",X"F9",X"F0",X"E0",
		X"F0",X"F0",X"F0",X"E8",X"88",X"AA",X"FF",X"33",X"F0",X"F0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"11",X"00",X"00",X"11",X"62",X"62",X"30",X"88",X"B8",X"F8",X"70",X"F8",X"FC",X"74",
		X"80",X"C0",X"C0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"F0",X"C0",X"C0",X"C0",X"80",X"00",X"00",
		X"62",X"71",X"F1",X"F0",X"F0",X"F0",X"70",X"00",X"FE",X"BB",X"11",X"FF",X"F6",X"F0",X"F0",X"F0",
		X"E0",X"E0",X"E0",X"E4",X"EE",X"77",X"00",X"00",X"00",X"00",X"00",X"88",X"CC",X"CC",X"88",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"10",X"00",X"00",X"66",X"BB",X"11",
		X"30",X"10",X"C0",X"C0",X"70",X"70",X"F0",X"F0",X"00",X"C0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",
		X"10",X"30",X"30",X"30",X"10",X"10",X"10",X"00",X"BB",X"EE",X"C4",X"E6",X"F3",X"F3",X"F0",X"30",
		X"F8",X"F8",X"74",X"FC",X"FB",X"FB",X"C0",X"C0",X"F0",X"F0",X"E0",X"C0",X"80",X"AA",X"FF",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"10",X"00",X"00",X"70",
		X"00",X"00",X"20",X"20",X"20",X"80",X"00",X"00",X"00",X"00",X"00",X"20",X"40",X"80",X"00",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"20",X"00",X"00",X"00",X"00",
		X"00",X"80",X"20",X"20",X"20",X"00",X"00",X"00",X"00",X"80",X"40",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"70",X"70",X"D5",X"88",X"DD",X"FF",X"F8",X"00",X"00",X"E0",X"E8",X"E8",X"E8",X"E0",X"E8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F6",X"F7",X"F3",X"F0",X"70",X"60",X"E0",X"00",X"EC",X"EC",X"E8",X"E0",X"60",X"60",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"73",X"51",X"51",X"F3",X"D1",X"00",X"20",X"60",X"E0",X"E0",X"C0",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"D1",X"D1",X"73",X"73",X"72",X"70",X"30",X"00",X"C0",X"C0",X"E0",X"E4",X"EC",X"E8",X"20",X"00",
		X"00",X"00",X"00",X"33",X"77",X"57",X"47",X"67",X"11",X"33",X"EF",X"EF",X"FF",X"F2",X"F8",X"3C",
		X"FF",X"F1",X"FF",X"7F",X"FF",X"F9",X"F0",X"F0",X"00",X"CC",X"E6",X"EE",X"EE",X"EE",X"EE",X"E6",
		X"33",X"00",X"00",X"11",X"11",X"11",X"00",X"00",X"BC",X"FF",X"F9",X"D2",X"3E",X"CF",X"77",X"00",
		X"FC",X"F4",X"F0",X"FD",X"F3",X"F4",X"8F",X"FF",X"EE",X"EE",X"CC",X"EE",X"EE",X"E6",X"E6",X"CC",
		X"00",X"00",X"00",X"33",X"77",X"FF",X"BE",X"9F",X"77",X"74",X"BF",X"9F",X"FF",X"FD",X"F0",X"F0",
		X"CC",X"F7",X"FD",X"FF",X"FF",X"F3",X"F1",X"F0",X"00",X"00",X"88",X"88",X"CC",X"CC",X"CC",X"CC",
		X"CF",X"77",X"11",X"11",X"32",X"11",X"11",X"00",X"79",X"7E",X"FE",X"D2",X"B4",X"4F",X"FF",X"00",
		X"F9",X"F9",X"F1",X"FB",X"F3",X"F4",X"8F",X"FF",X"CC",X"88",X"CC",X"EE",X"EE",X"E6",X"C4",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"00",X"00",X"70",X"F3",X"C4",X"F7",X"F7",X"C4",
		X"00",X"00",X"C2",X"E9",X"E9",X"C3",X"CB",X"E9",X"00",X"00",X"00",X"20",X"28",X"E0",X"28",X"08",
		X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"F7",X"F7",X"F3",X"78",X"3C",X"34",X"00",X"00",
		X"E9",X"E9",X"C3",X"87",X"1F",X"1D",X"77",X"00",X"28",X"28",X"E0",X"28",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"30",X"35",X"35",X"35",X"35",X"00",X"00",X"F0",X"FE",X"FE",X"30",X"FE",X"FE",
		X"00",X"00",X"28",X"96",X"96",X"1E",X"0E",X"A4",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",
		X"35",X"35",X"34",X"16",X"03",X"01",X"00",X"00",X"32",X"FE",X"FC",X"E1",X"C3",X"C3",X"00",X"00",
		X"B4",X"96",X"1E",X"0E",X"2E",X"2A",X"33",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"88",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"78",X"59",X"59",X"7A",X"7B",X"59",X"00",X"00",X"08",X"A4",X"A4",X"E0",X"A4",X"84",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"59",X"7A",X"78",X"2D",X"2D",X"25",X"00",X"00",X"A4",X"A4",X"68",X"2C",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"13",X"02",X"00",X"00",X"00",X"21",X"F0",X"BA",X"BB",X"33",
		X"30",X"00",X"10",X"2C",X"0F",X"87",X"C3",X"E9",X"00",X"80",X"00",X"00",X"00",X"28",X"1C",X"78",
		X"12",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"EE",X"E6",X"6A",X"3D",X"16",X"01",X"00",X"00",
		X"21",X"FC",X"ED",X"F8",X"F0",X"1E",X"00",X"00",X"1C",X"0C",X"0C",X"6E",X"91",X"22",X"00",X"00",
		X"00",X"00",X"10",X"10",X"30",X"30",X"30",X"30",X"00",X"00",X"11",X"88",X"11",X"88",X"91",X"90",
		X"00",X"00",X"80",X"C0",X"D0",X"E1",X"E1",X"F0",X"00",X"00",X"02",X"0E",X"86",X"C0",X"48",X"0C",
		X"30",X"30",X"11",X"11",X"00",X"00",X"00",X"00",X"90",X"FC",X"FE",X"99",X"99",X"77",X"00",X"00",
		X"F0",X"94",X"87",X"07",X"07",X"03",X"03",X"00",X"86",X"C2",X"C0",X"68",X"60",X"68",X"20",X"00",
		X"00",X"00",X"10",X"10",X"30",X"30",X"30",X"30",X"00",X"00",X"64",X"B8",X"74",X"B8",X"F4",X"90",
		X"00",X"00",X"01",X"00",X"10",X"90",X"B0",X"F0",X"00",X"00",X"08",X"06",X"C0",X"C0",X"C2",X"C2",
		X"30",X"30",X"11",X"11",X"00",X"00",X"00",X"00",X"D0",X"FC",X"32",X"11",X"BB",X"77",X"00",X"00",
		X"F0",X"B4",X"86",X"0C",X"0E",X"0C",X"06",X"00",X"0E",X"C2",X"C0",X"60",X"60",X"60",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"72",X"50",X"F2",X"D0",X"F2",X"D0",X"00",X"00",X"02",X"42",X"42",X"E0",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F4",X"BA",X"AB",X"AB",X"AB",X"45",X"00",X"C2",X"86",X"C2",X"60",X"28",X"20",X"68",X"00",
		X"00",X"00",X"00",X"00",X"10",X"10",X"30",X"30",X"00",X"00",X"00",X"20",X"A8",X"30",X"74",X"90",
		X"00",X"02",X"03",X"01",X"01",X"10",X"03",X"B0",X"00",X"00",X"00",X"08",X"00",X"80",X"08",X"0E",
		X"30",X"30",X"30",X"30",X"10",X"10",X"00",X"00",X"E2",X"E0",X"E0",X"F6",X"99",X"99",X"DD",X"66",
		X"F0",X"D2",X"94",X"87",X"84",X"86",X"04",X"00",X"48",X"C0",X"E0",X"A0",X"60",X"40",X"40",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"71",X"63",X"63",X"73",X"73",
		X"00",X"00",X"E0",X"FC",X"7C",X"7C",X"FC",X"E8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"73",X"73",X"63",X"63",X"71",X"30",X"00",X"00",
		X"E8",X"FC",X"7C",X"7C",X"FC",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"71",X"73",X"E3",X"E7",X"F7",
		X"00",X"00",X"E0",X"FE",X"7E",X"FC",X"FC",X"E8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F7",X"E7",X"E3",X"73",X"71",X"30",X"00",X"00",
		X"E8",X"FC",X"FC",X"7E",X"FE",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"11",X"11",X"00",X"00",X"00",X"66",X"BF",X"1F",X"1F",X"2E",X"CC",X"00",
		X"00",X"00",X"22",X"55",X"55",X"66",X"88",X"99",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"88",
		X"00",X"11",X"11",X"11",X"00",X"00",X"00",X"00",X"CC",X"2E",X"1F",X"1F",X"BF",X"66",X"00",X"00",
		X"88",X"66",X"55",X"55",X"22",X"00",X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"1F",X"8F",X"8F",X"9F",X"66",X"00",
		X"00",X"66",X"11",X"AA",X"AA",X"11",X"11",X"11",X"00",X"00",X"00",X"88",X"88",X"44",X"44",X"CC",
		X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"66",X"9F",X"8F",X"8F",X"1F",X"EE",X"00",X"00",
		X"11",X"11",X"AA",X"AA",X"11",X"66",X"00",X"00",X"44",X"44",X"88",X"88",X"00",X"00",X"00",X"00",
		X"01",X"02",X"03",X"01",X"00",X"00",X"01",X"01",X"01",X"00",X"0E",X"0D",X"06",X"01",X"03",X"0A",
		X"00",X"0C",X"06",X"0E",X"86",X"CA",X"C3",X"F5",X"00",X"00",X"02",X"04",X"0C",X"0C",X"08",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"10",X"10",X"10",X"30",X"31",X"32",X"44",
		X"7E",X"F6",X"ED",X"EC",X"C8",X"C0",X"00",X"00",X"0C",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",
		X"18",X"12",X"12",X"24",X"24",X"03",X"01",X"00",X"E1",X"7A",X"12",X"00",X"00",X"00",X"08",X"04",
		X"7E",X"3F",X"F2",X"F2",X"7E",X"3F",X"36",X"63",X"9A",X"BC",X"E8",X"C2",X"C2",X"8C",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"11",X"32",X"22",X"22",
		X"6A",X"68",X"CC",X"88",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"02",X"07",X"21",X"21",X"01",X"14",X"0B",X"00",X"00",X"01",X"00",X"00",X"08",X"0E",X"0F",
		X"00",X"08",X"24",X"12",X"03",X"01",X"00",X"01",X"04",X"80",X"08",X"08",X"08",X"0C",X"0E",X"0E",
		X"10",X"00",X"01",X"03",X"03",X"06",X"04",X"08",X"0F",X"E5",X"3E",X"69",X"3C",X"03",X"01",X"87",
		X"0B",X"1A",X"1F",X"B4",X"FA",X"E5",X"E3",X"7E",X"4A",X"84",X"48",X"80",X"82",X"02",X"01",X"92",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",
		X"71",X"71",X"3F",X"71",X"30",X"60",X"C0",X"80",X"CC",X"8E",X"E9",X"49",X"01",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"31",X"20",X"22",X"60",X"40",X"44",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"07",X"07",X"06",X"06",X"02",X"01",X"0F",X"4B",X"96",X"0B",X"01",X"00",X"01",X"03",
		X"7A",X"F4",X"F0",X"F0",X"3C",X"3C",X"3D",X"F6",X"CE",X"E3",X"C2",X"D3",X"E5",X"CE",X"FF",X"E2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"06",X"04",X"02",X"00",X"00",X"00",X"00",
		X"3C",X"1E",X"07",X"03",X"07",X"18",X"12",X"13",X"D2",X"AC",X"E1",X"E0",X"E2",X"F4",X"8E",X"84",
		X"00",X"03",X"06",X"06",X"0E",X"0F",X"2D",X"16",X"00",X"01",X"01",X"12",X"06",X"00",X"0C",X"86",
		X"06",X"0F",X"C7",X"6B",X"70",X"21",X"21",X"03",X"00",X"06",X"02",X"38",X"2C",X"6B",X"6A",X"D6",
		X"13",X"01",X"00",X"03",X"34",X"08",X"0A",X"04",X"58",X"C8",X"6C",X"1E",X"1E",X"87",X"43",X"01",
		X"07",X"3D",X"7B",X"F6",X"F0",X"F0",X"3D",X"7B",X"BD",X"E2",X"EE",X"E7",X"C6",X"E6",X"EE",X"E9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"06",X"1F",X"06",X"02",X"00",X"00",X"00",X"77",X"88",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"CC",X"22",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"22",X"CC",X"00",X"00",X"00",X"00",X"77",X"88",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"CC",X"22",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"07",X"0F",X"22",X"11",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"88",X"88",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"11",X"22",X"44",X"44",X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"44",X"22",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"11",X"22",X"44",X"44",X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"07",X"07",X"07",X"07",X"07",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"08",X"0C",X"0E",X"0E",X"0E",X"0E",X"0E",
		X"07",X"07",X"07",X"07",X"07",X"03",X"01",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"0E",X"0E",X"0E",X"0E",X"0E",X"0C",X"08",X"00",
		X"03",X"03",X"03",X"03",X"03",X"03",X"01",X"00",X"69",X"96",X"87",X"87",X"69",X"0F",X"0F",X"00",
		X"2D",X"2D",X"A5",X"69",X"2D",X"0F",X"0F",X"00",X"08",X"08",X"08",X"08",X"08",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"03",X"03",X"03",X"03",X"01",X"00",X"69",X"96",X"96",X"96",X"87",X"0F",X"0F",X"00",
		X"C3",X"2D",X"2D",X"2D",X"2D",X"0F",X"0F",X"00",X"08",X"08",X"08",X"08",X"08",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"03",X"03",X"03",X"03",X"01",X"00",X"0F",X"F0",X"4B",X"2D",X"1E",X"0F",X"0F",X"00",
		X"87",X"E1",X"87",X"87",X"87",X"0F",X"0F",X"00",X"08",X"08",X"08",X"08",X"08",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"03",X"03",X"03",X"03",X"01",X"00",X"96",X"A5",X"A5",X"A5",X"E1",X"0F",X"0F",X"00",
		X"C3",X"2D",X"2D",X"2D",X"4B",X"0F",X"0F",X"00",X"08",X"08",X"08",X"08",X"08",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"03",X"03",X"03",X"03",X"01",X"00",X"0F",X"96",X"96",X"5A",X"3C",X"0F",X"0F",X"00",
		X"C3",X"2D",X"2D",X"2D",X"C3",X"0F",X"0F",X"00",X"08",X"08",X"08",X"08",X"08",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"03",X"03",X"03",X"03",X"01",X"00",X"69",X"96",X"96",X"96",X"69",X"0F",X"0F",X"00",
		X"C3",X"2D",X"2D",X"2D",X"C3",X"0F",X"0F",X"00",X"08",X"08",X"08",X"08",X"08",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"78",X"87",X"87",X"78",X"0F",X"0F",X"F0",X"0F",
		X"C3",X"2D",X"2D",X"C3",X"0F",X"0F",X"E1",X"0F",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"96",X"A5",X"A5",X"E1",X"0F",X"69",X"96",X"87",
		X"C3",X"2D",X"2D",X"4B",X"0F",X"2D",X"2D",X"A5",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"87",X"4B",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"69",X"2D",X"0F",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"78",X"87",X"87",X"78",X"0F",X"0F",X"F0",X"4B",
		X"C3",X"2D",X"2D",X"C3",X"0F",X"87",X"E1",X"87",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"2D",X"1E",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"87",X"87",X"0F",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"78",X"87",X"87",X"78",X"0F",X"0F",X"96",X"96",
		X"C3",X"2D",X"2D",X"C3",X"0F",X"C3",X"2D",X"2D",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"5A",X"3C",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"2D",X"C3",X"0F",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"78",X"87",X"87",X"78",X"0F",X"69",X"96",X"96",
		X"C3",X"2D",X"2D",X"C3",X"0F",X"C3",X"2D",X"2D",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"96",X"69",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"2D",X"C3",X"0F",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"78",X"87",X"87",X"78",X"0F",X"78",X"87",X"87",
		X"C3",X"2D",X"2D",X"C3",X"0F",X"C3",X"2D",X"2D",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"78",X"0F",X"F0",X"4B",X"00",X"00",X"00",X"00",
		X"C3",X"0F",X"E1",X"0F",X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"78",X"87",X"87",X"78",X"0F",X"69",X"96",X"87",
		X"C3",X"2D",X"2D",X"C3",X"0F",X"2D",X"2D",X"A5",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"4B",X"0F",X"F0",X"4B",X"00",X"00",X"00",X"00",
		X"69",X"0F",X"E1",X"0F",X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"78",X"87",X"87",X"78",X"0F",X"96",X"A5",X"A5",
		X"C3",X"2D",X"2D",X"C3",X"0F",X"C3",X"2D",X"2D",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"E1",X"0F",X"F0",X"4B",X"00",X"00",X"00",X"00",
		X"4B",X"0F",X"E1",X"0F",X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"0F",X"78",X"87",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"C3",X"2D",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"87",X"78",X"0F",X"78",X"87",X"87",X"78",X"0F",
		X"2D",X"C3",X"0F",X"C3",X"2D",X"2D",X"C3",X"0F",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"FF",X"FF",X"CF",X"8F",X"9F",X"9F",X"9F",X"9F",
		X"FF",X"FF",X"0F",X"0F",X"FF",X"FF",X"FF",X"FF",X"EE",X"EE",X"6E",X"6E",X"EE",X"EE",X"EE",X"EE",
		X"11",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"8F",X"8F",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"6E",X"6E",X"EE",X"CC",X"00",X"00",X"00",X"00",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"8F",X"9F",X"9F",X"8F",X"8F",X"FF",X"FF",X"CF",
		X"0F",X"FF",X"FF",X"0F",X"0F",X"FF",X"FF",X"0F",X"6E",X"EE",X"EE",X"6E",X"6E",X"EE",X"EE",X"6E",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"8F",X"8F",X"9F",X"9F",X"9F",X"9F",X"9F",X"FF",
		X"0F",X"0F",X"2F",X"2F",X"2F",X"2F",X"0F",X"0F",X"6E",X"6E",X"6E",X"6E",X"6E",X"6E",X"6E",X"6E",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"FF",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"8F",
		X"FF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"0F",X"EE",X"6E",X"6E",X"6E",X"6E",X"6E",X"6E",X"6E",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"CF",X"FF",X"FF",X"CF",X"8F",X"9F",X"9F",X"8F",
		X"0F",X"FF",X"FF",X"0F",X"0F",X"FF",X"FF",X"0F",X"EE",X"EE",X"EE",X"6E",X"6E",X"EE",X"EE",X"6E",
		X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"00",X"00",X"00",X"00",X"FF",X"FF",X"CF",X"8F",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"0F",X"0F",X"00",X"00",X"00",X"00",X"CC",X"EE",X"EE",X"6E",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"9F",X"9F",X"9F",X"9F",X"9F",X"8F",X"CF",X"FF",
		X"EF",X"EF",X"EF",X"EF",X"EF",X"0F",X"0F",X"FF",X"6E",X"6E",X"6E",X"6E",X"6E",X"6E",X"EE",X"EE",
		X"00",X"10",X"00",X"00",X"10",X"10",X"10",X"33",X"00",X"E0",X"60",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"F0",X"30",X"F0",X"E0",X"E0",X"F1",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",
		X"66",X"DD",X"DD",X"DC",X"44",X"00",X"00",X"00",X"FF",X"22",X"AA",X"F0",X"70",X"10",X"10",X"00",
		X"FC",X"76",X"FE",X"F0",X"F0",X"F0",X"C0",X"00",X"CC",X"E6",X"E6",X"FF",X"E6",X"00",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"10",X"10",X"70",X"EE",X"FF",X"11",X"E6",X"D5",X"91",X"F7",X"91",
		X"00",X"00",X"88",X"F8",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"20",X"A0",X"E0",X"E0",X"80",
		X"70",X"70",X"30",X"30",X"10",X"11",X"11",X"00",X"D5",X"F7",X"F6",X"F0",X"F9",X"FF",X"EE",X"88",
		X"F0",X"F0",X"F0",X"C4",X"CC",X"00",X"00",X"00",X"A0",X"A0",X"E0",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"88",X"88",X"77",X"00",X"66",X"99",X"88",
		X"CC",X"22",X"22",X"CC",X"00",X"22",X"22",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"44",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"88",X"88",X"77",X"00",X"88",X"DD",X"BB",
		X"CC",X"22",X"22",X"CC",X"00",X"CC",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"88",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"88",X"88",X"77",X"00",X"99",X"AA",X"AA",
		X"CC",X"22",X"22",X"CC",X"00",X"CC",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"88",X"88",X"77",X"00",X"CC",X"AA",X"99",
		X"CC",X"22",X"22",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"74",X"16",X"07",X"05",X"07",X"07",X"07",X"07",
		X"00",X"C0",X"68",X"3C",X"16",X"0F",X"0D",X"0F",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"07",X"07",X"05",X"07",X"16",X"74",
		X"0F",X"0D",X"0F",X"16",X"3C",X"68",X"C0",X"00",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"20",X"10",X"00",X"70",X"11",X"01",X"01",X"40",X"40",X"40",X"C7",X"8F",X"0F",X"1F",X"6F",
		X"00",X"00",X"00",X"08",X"0C",X"0E",X"0F",X"2F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"07",X"03",X"00",X"00",X"00",X"00",X"00",
		X"4F",X"0F",X"1F",X"2F",X"07",X"01",X"00",X"00",X"08",X"08",X"0C",X"0C",X"0C",X"0C",X"00",X"00",
		X"00",X"30",X"70",X"11",X"00",X"00",X"00",X"00",X"00",X"F4",X"F0",X"F1",X"10",X"00",X"00",X"00",
		X"00",X"88",X"E0",X"F0",X"F2",X"F0",X"72",X"30",X"00",X"00",X"00",X"00",X"C0",X"C0",X"E0",X"E4",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"30",X"30",X"30",X"31",X"10",X"00",X"00",X"E0",X"E8",X"E0",X"C0",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"10",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"20",X"A0",X"60",X"F0",X"71",X"23",
		X"00",X"00",X"00",X"00",X"47",X"8F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"08",X"0C",X"0E",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"47",X"07",X"07",X"07",X"03",X"01",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"0E",X"0E",X"0E",X"0E",X"0E",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"10",X"10",X"10",X"00",X"30",X"00",X"F0",X"F0",X"F7",X"FF",X"D7",X"D7",X"F0",
		X"00",X"00",X"90",X"F9",X"FF",X"5F",X"6F",X"DF",X"00",X"00",X"80",X"C0",X"E8",X"FE",X"FC",X"E0",
		X"70",X"40",X"00",X"10",X"10",X"10",X"00",X"00",X"E1",X"E3",X"F3",X"F7",X"F7",X"F0",X"F0",X"00",
		X"AF",X"BF",X"FF",X"FF",X"F8",X"90",X"00",X"00",X"E8",X"FC",X"FC",X"E0",X"C0",X"80",X"00",X"00",
		X"00",X"11",X"77",X"33",X"33",X"00",X"00",X"00",X"00",X"CF",X"8F",X"EF",X"8F",X"8F",X"03",X"01",
		X"00",X"0C",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"08",X"0C",X"0C",X"0E",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"4B",X"69",X"3C",X"0F",X"07",X"03",X"00",X"0F",X"0F",X"0F",X"0F",X"0E",X"0E",X"0C",X"00",
		X"00",X"00",X"00",X"01",X"13",X"33",X"77",X"67",X"00",X"00",X"77",X"DF",X"9F",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"88",X"88",X"98",X"F8",X"F8",X"00",X"00",X"00",X"00",X"C0",X"68",X"2C",X"A4",
		X"47",X"77",X"33",X"33",X"11",X"00",X"00",X"00",X"CF",X"EF",X"FF",X"7F",X"3F",X"77",X"00",X"00",
		X"F8",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"84",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"22",X"11",X"11",X"01",X"77",X"00",X"01",X"07",X"0F",X"8F",X"CF",X"4F",X"AF",
		X"00",X"0C",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"08",X"0C",X"0C",X"0E",X"0E",
		X"11",X"11",X"10",X"11",X"00",X"00",X"00",X"00",X"E7",X"CF",X"CF",X"2D",X"1E",X"07",X"01",X"00",
		X"2D",X"69",X"C3",X"0F",X"87",X"0F",X"0C",X"00",X"0E",X"0E",X"0C",X"0C",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"10",X"30",X"30",X"61",X"D2",X"3C",
		X"00",X"F0",X"F0",X"F0",X"1E",X"E1",X"F0",X"F0",X"00",X"00",X"80",X"95",X"E6",X"84",X"7F",X"84",
		X"30",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F2",X"F1",X"70",X"31",X"10",X"00",X"00",
		X"F0",X"F1",X"FE",X"F0",X"F3",X"FC",X"F0",X"00",X"FF",X"84",X"F7",X"E2",X"D1",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"03",X"21",X"61",X"C3",
		X"00",X"00",X"00",X"88",X"CC",X"6E",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"C3",X"61",X"21",X"03",X"FF",X"00",X"00",
		X"0F",X"08",X"0C",X"6E",X"CC",X"88",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"50",X"50",X"20",X"93",X"70",X"00",X"00",X"00",X"00",X"13",X"A3",X"A7",X"D7",
		X"00",X"00",X"00",X"0D",X"8F",X"3F",X"CF",X"0F",X"00",X"00",X"00",X"08",X"CC",X"2E",X"0E",X"CE",
		X"61",X"B0",X"20",X"50",X"50",X"00",X"00",X"00",X"DF",X"A7",X"A3",X"13",X"00",X"00",X"00",X"00",
		X"3F",X"CF",X"0F",X"BF",X"0D",X"00",X"00",X"00",X"2E",X"0E",X"CE",X"0C",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"44",X"22",X"11",X"00",X"00",X"00",
		X"88",X"EE",X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"55",X"33",X"00",X"00",X"00",
		X"CC",X"22",X"22",X"22",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"99",X"99",X"99",X"66",X"00",X"00",X"00",
		X"CC",X"22",X"22",X"22",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"88",X"88",X"77",X"00",X"FF",X"44",X"00",
		X"CC",X"22",X"22",X"CC",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"88",X"88",X"77",X"00",X"00",X"FF",X"44",
		X"CC",X"22",X"22",X"CC",X"00",X"88",X"EE",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"11",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"88",X"88",X"77",X"00",X"00",X"99",X"99",
		X"CC",X"22",X"22",X"CC",X"00",X"CC",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"33",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"88",X"88",X"77",X"00",X"66",X"99",X"99",
		X"CC",X"22",X"22",X"CC",X"00",X"CC",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"66",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"77",X"00",X"77",X"88",X"88",X"77",X"00",
		X"22",X"CC",X"00",X"CC",X"22",X"22",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"40",X"40",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"20",X"40",X"40",X"40",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"22",X"22",X"22",X"22",X"EE",X"EE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"FF",X"88",X"88",X"88",X"FF",X"FF",X"00",X"00",X"88",X"88",X"88",X"88",X"EE",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"FF",X"11",X"11",X"FF",X"EE",X"00",X"00",X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"77",X"CC",X"88",X"CC",X"77",X"33",X"00",X"EE",X"EE",X"88",X"88",X"88",X"EE",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"FF",X"99",X"88",X"88",X"FF",X"FF",X"00",X"22",X"66",X"EE",X"CC",X"88",X"EE",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"99",X"99",X"99",X"99",X"FF",X"FF",X"00",X"22",X"22",X"22",X"22",X"22",X"EE",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"33",X"00",X"00",X"00",X"00",X"CC",X"EE",X"AE",X"1F",
		X"00",X"40",X"80",X"C0",X"70",X"70",X"30",X"00",X"00",X"00",X"20",X"40",X"40",X"A0",X"E0",X"60",
		X"33",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"1F",X"BF",X"EE",X"CC",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"30",X"70",X"40",X"20",X"10",X"00",X"E0",X"60",X"C0",X"20",X"20",X"40",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"44",X"00",X"00",X"00",X"22",X"22",X"EE",X"EE",X"22",X"22",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"FF",X"BB",X"99",X"99",X"CC",X"44",X"00",X"22",X"22",X"AA",X"AA",X"EE",X"EE",X"66",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"99",X"99",X"99",X"99",X"FF",X"FF",X"00",X"22",X"22",X"22",X"22",X"22",X"EE",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"FF",X"99",X"88",X"88",X"FF",X"FF",X"00",X"22",X"66",X"EE",X"CC",X"88",X"EE",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"77",X"CC",X"88",X"88",X"FF",X"FF",X"00",X"88",X"CC",X"66",X"22",X"22",X"EE",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"77",X"CC",X"88",X"CC",X"77",X"33",X"00",X"EE",X"EE",X"88",X"88",X"88",X"EE",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"FF",X"11",X"11",X"FF",X"EE",X"00",X"00",X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"77",X"CC",X"88",X"CC",X"77",X"33",X"00",X"EE",X"EE",X"88",X"88",X"88",X"EE",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"99",X"99",X"88",X"CC",X"77",X"33",X"00",X"EE",X"EE",X"22",X"22",X"66",X"CC",X"88",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"99",X"99",X"99",X"99",X"FF",X"FF",X"00",X"22",X"22",X"22",X"22",X"22",X"EE",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"77",X"33",X"77",X"FF",X"FF",X"00",X"EE",X"EE",X"00",X"88",X"00",X"EE",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"11",X"00",X"11",X"FF",X"FF",X"00",X"00",X"88",X"CC",X"EE",X"CC",X"88",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"FF",X"88",X"88",X"88",X"FF",X"77",X"00",X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"88",X"88",X"44",X"44",X"22",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"22",X"0F",X"07",X"02",X"88",X"88",X"88",X"00",X"00",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"88",X"88",X"44",X"44",X"22",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"11",X"22",X"44",X"44",X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",
		X"00",X"33",X"56",X"56",X"67",X"33",X"00",X"00",X"77",X"F8",X"F0",X"F0",X"F0",X"0F",X"FF",X"00",
		X"CC",X"7B",X"3F",X"BF",X"CF",X"F1",X"79",X"BC",X"00",X"62",X"62",X"88",X"EE",X"EE",X"EA",X"E2",
		X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"00",X"00",X"00",X"00",X"11",X"FE",X"3C",X"DE",X"33",
		X"76",X"11",X"33",X"FD",X"F8",X"F4",X"C3",X"FF",X"E6",X"CC",X"EE",X"EE",X"EA",X"E2",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"30",X"16",X"01",X"00",X"44",X"6A",X"26",X"00",X"C4",X"E2",X"6A",X"26",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"80",X"C4",X"48",X"08",X"44",X"6A",X"68",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"20",
		X"00",X"10",X"31",X"31",X"20",X"35",X"35",X"16",X"E1",X"ED",X"A9",X"30",X"31",X"FF",X"CC",X"CC",
		X"0F",X"0F",X"0F",X"87",X"C3",X"E9",X"65",X"ED",X"48",X"0C",X"0E",X"0E",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"16",X"07",X"03",X"03",X"01",X"01",X"00",X"00",X"D5",X"F3",X"79",X"3C",X"1E",X"0F",X"0F",X"03",
		X"ED",X"ED",X"E9",X"C3",X"4B",X"2D",X"3C",X"1E",X"0F",X"0F",X"0F",X"0F",X"0E",X"0E",X"2E",X"22",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"44",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"87",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",
		X"00",X"00",X"01",X"01",X"03",X"03",X"03",X"03",X"71",X"F3",X"80",X"80",X"D5",X"F7",X"F7",X"E6",
		X"CB",X"E9",X"E9",X"E9",X"C3",X"87",X"C3",X"E9",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"80",X"80",X"00",X"08",X"08",X"08",X"08",X"48",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"03",X"03",X"03",X"01",X"01",X"00",X"C4",X"C0",X"F3",X"7B",X"78",X"3C",X"1E",X"1E",
		X"74",X"74",X"FC",X"ED",X"E1",X"C3",X"0F",X"87",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C3",X"4B",X"43",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0E",X"48",X"C0",X"48",X"08",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"2E",X"2A",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"08",
		X"00",X"00",X"00",X"22",X"00",X"11",X"11",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"00",X"DD",X"66",X"26",X"06",X"0C",X"E1",X"FE",
		X"EE",X"88",X"01",X"00",X"08",X"04",X"06",X"0E",X"00",X"00",X"00",X"08",X"0C",X"0E",X"0E",X"07",
		X"00",X"00",X"00",X"00",X"00",X"88",X"99",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"26",X"03",X"01",X"09",X"09",X"0D",X"0F",X"00",X"00",X"00",X"00",X"08",X"08",X"48",X"48",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"31",X"31",X"30",X"10",X"01",X"01",X"00",X"00",X"DD",X"99",X"11",X"FF",X"F7",X"F3",X"79",X"3C",
		X"0F",X"F0",X"FE",X"11",X"33",X"77",X"FF",X"F6",X"0F",X"0F",X"87",X"87",X"C3",X"C3",X"C3",X"C3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"3C",X"0F",X"03",X"00",X"00",X"00",X"00",X"87",X"C3",X"4B",X"4B",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"C0",X"08",X"08",X"08",X"08",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"1F",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",
		X"00",X"31",X"20",X"60",X"60",X"F1",X"F0",X"F0",X"40",X"40",X"60",X"E8",X"70",X"70",X"74",X"30",
		X"00",X"71",X"73",X"F7",X"F7",X"F7",X"F3",X"F1",X"06",X"BE",X"FF",X"FF",X"EF",X"EF",X"EF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"C0",X"C0",X"48",X"48",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"71",X"71",X"31",X"00",X"90",X"D0",X"F0",X"FC",X"32",X"32",X"32",X"EC",
		X"F0",X"F0",X"F0",X"F0",X"E1",X"D2",X"43",X"03",X"F7",X"F0",X"F0",X"F0",X"F0",X"F0",X"78",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"84",X"C0",X"E0",X"E0",X"E0",X"60",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"D4",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"F3",
		X"00",X"10",X"10",X"10",X"30",X"30",X"30",X"30",X"90",X"B2",X"90",X"D4",X"90",X"D1",X"C0",X"E0",
		X"90",X"B1",X"F1",X"F1",X"F1",X"F1",X"F0",X"70",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C8",X"8C",X"CA",X"8E",X"8E",X"EC",X"EC",X"C8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"30",X"30",X"30",X"30",X"10",X"10",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F3",X"C4",X"C4",
		X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"F1",X"F0",X"F0",X"F0",X"E1",X"D2",X"C3",X"43",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"33",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"78",X"F0",X"86",X"86",X"84",X"C0",X"E0",X"E0",X"E0",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"68",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"00",X"99",X"55",X"00",X"00",X"00",X"22",X"33",X"FF",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"F0",X"00",X"22",X"00",X"70",X"74",X"30",X"10",X"99",
		X"77",X"22",X"62",X"71",X"F7",X"F0",X"F0",X"F0",X"00",X"00",X"11",X"11",X"88",X"D5",X"F6",X"F8",
		X"00",X"00",X"00",X"01",X"23",X"AA",X"77",X"33",X"00",X"00",X"00",X"00",X"08",X"0C",X"0C",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"DD",X"FF",X"FC",X"F4",X"F0",X"C8",X"C0",X"C8",X"E0",X"E0",X"2C",X"2C",X"86",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"70",X"70",X"30",X"30",X"10",X"10",X"00",X"80",X"D0",X"F0",X"F0",X"F3",X"C4",X"C4",X"C4",
		X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"74",X"74",X"F0",X"F0",X"F0",X"F0",X"F0",X"B4",X"87",X"B4",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"33",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"F8",X"E0",X"00",X"00",X"00",X"00",X"00",X"07",X"04",X"03",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"C2",X"86",X"E0",X"E0",X"E0",X"E0",X"60",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"77",X"33",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"77",X"77",X"33",X"11",X"11",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"77",X"77",X"33",X"33",X"11",X"11",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"77",X"33",X"11",X"11",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"74",X"76",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"F3",X"F1",X"F0",X"F8",X"F8",X"FC",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"F3",X"F3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"77",X"33",X"33",X"11",X"11",X"00",X"74",X"74",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",
		X"F1",X"F0",X"F8",X"FC",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"F3",X"F3",X"F1",X"F1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"F3",X"F1",X"F8",X"FC",X"FC",X"FE",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"F7",X"F3",X"F8",X"FC",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F1",X"F9",X"FC",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"F7",X"F3",X"F1",X"F9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"77",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"F8",X"F8",
		X"F8",X"F8",X"F1",X"F3",X"F3",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"76",X"32",X"00",X"00",X"00",X"11",X"11",X"F1",X"F3",X"F3",X"77",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"77",X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FC",X"FC",X"F8",X"F0",X"F0",X"F0",X"F0",
		X"33",X"33",X"11",X"11",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"77",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"F8",X"FC",X"FC",X"FE",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"FF",X"FE",X"FE",X"FC",X"F9",X"FB",X"F3",X"F7",X"F7",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"FF",X"FF",X"77",X"77",X"32",X"10",X"11",X"11",X"FC",X"F9",X"F9",X"F3",X"F7",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"F8",X"FC",X"F8",X"F8",X"F1",X"F1",X"F3",X"F7",X"F7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"77",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"F8",X"F0",
		X"F8",X"F1",X"F1",X"F3",X"F7",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"FF",X"FE",X"FC",X"FC",X"70",X"00",X"11",X"11",X"F1",X"F3",X"F3",X"F3",X"F7",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"FE",X"FC",X"F8",X"F1",X"F1",X"F3",X"F3",X"F7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"33",X"77",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",
		X"00",X"11",X"33",X"33",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"33",X"33",X"33",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"33",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"FD",X"FB",X"F3",
		X"0F",X"0F",X"87",X"87",X"C3",X"F0",X"F8",X"F8",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"E1",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"0F",
		X"FC",X"FE",X"EF",X"CF",X"8F",X"8F",X"0F",X"0F",X"87",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"C0",X"E0",X"3C",X"0F",X"0F",X"0F",X"0E",X"0C",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"1E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"08",X"0C",X"0C",X"0E",X"0E",X"0E",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"1E",X"3C",X"1E",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"F0",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"03",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"F0",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"E7",X"E3",X"E1",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0E",X"0C",
		X"CB",X"8F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"FE",X"7F",X"6F",X"6F",X"6F",X"6F",X"6F",X"6B",X"87",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"6B",X"69",X"69",X"78",X"78",X"3C",X"1E",X"0F",X"0F",X"0F",X"0F",X"0F",X"87",X"F0",X"F0",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"2C",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"1E",X"F0",X"F0",X"0F",X"0F",X"EF",X"EF",X"E7",X"E3",X"E3",X"C3",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"87",X"C3",X"E1",X"E1",X"F8",X"FC",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"87",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"FC",X"FE",X"FE",X"CF",X"8F",X"0F",X"0F",X"0F",X"E1",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0E",X"0C",X"08",
		X"0F",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"1E",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"80",X"C0",X"0C",X"0E",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"1E",X"3C",X"3C",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"8F",X"CB",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"C3",X"E3",X"E7",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0E",X"2C",X"C0",X"C0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F1",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"FC",X"FC",X"F6",X"F3",X"F3",X"F1",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"FC",X"FC",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"C0",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"C0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"E0",
		X"0F",X"0F",X"0F",X"8F",X"CB",X"F0",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"F0",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"F0",
		X"F0",X"87",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"4B",X"C7",X"E7",X"CF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"8F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"8F",X"CF",X"F8",X"F8",X"F0",X"F0",X"E1",X"0F",X"0F",X"0F",X"F0",X"F0",X"E1",X"C3",X"0F",
		X"0F",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"0F",
		X"C3",X"87",X"87",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"F0",X"F0",X"1E",X"0F",X"0F",X"0F",X"0E",X"2C",X"C0",X"80",X"80",X"08",X"0C",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0E",X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"03",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"08",X"09",X"2B",X"6F",X"6F",X"6F",X"6F",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"6F",X"6F",X"6F",X"7E",X"7C",X"3C",X"1E",X"0F",X"0F",X"0F",X"0F",X"0F",X"87",X"F0",X"F0",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0C",X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"1F",X"F3",X"F6",X"0F",X"0F",X"EF",X"ED",X"E9",X"E1",X"E1",X"C3",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"8F",X"CF",X"EF",X"FC",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"F8",X"F8",X"F0",X"87",X"0F",X"0F",X"0F",X"0F",X"87",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0E",
		X"0F",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0C",X"80",X"00",X"08",X"0C",X"0E",X"0F",X"0F",
		X"00",X"01",X"03",X"03",X"0F",X"69",X"69",X"69",X"3C",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"96",X"87",X"96",X"96",X"96",X"96",X"96",X"96",X"F0",X"C3",X"4B",X"F0",X"F0",X"F0",X"F0",X"B4",
		X"69",X"69",X"0F",X"69",X"2D",X"34",X"16",X"12",X"F0",X"F0",X"F0",X"F0",X"78",X"78",X"78",X"F0",
		X"96",X"87",X"96",X"D2",X"F0",X"E1",X"F0",X"F0",X"4B",X"C3",X"78",X"F0",X"F0",X"78",X"0F",X"C3",
		X"B4",X"78",X"78",X"F0",X"A5",X"69",X"B4",X"F0",X"86",X"C3",X"E1",X"3C",X"F0",X"78",X"3C",X"96",
		X"03",X"30",X"0F",X"0F",X"3C",X"3C",X"3C",X"3C",X"F6",X"F2",X"F3",X"F1",X"F1",X"F0",X"F0",X"F0",
		X"78",X"78",X"B4",X"78",X"F0",X"E1",X"0F",X"3C",X"F0",X"F0",X"F0",X"F0",X"1E",X"0F",X"E1",X"F0",
		X"3C",X"3C",X"3C",X"F0",X"F0",X"F0",X"78",X"78",X"F1",X"F1",X"F3",X"F2",X"F6",X"F4",X"FC",X"F9",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"78",X"3C",X"16",X"03",X"00",X"00",X"00",
		X"F0",X"F0",X"C3",X"87",X"3F",X"7F",X"37",X"03",X"F0",X"F0",X"0F",X"0F",X"FF",X"FF",X"FF",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"78",X"3C",X"BC",X"CE",X"8C",X"08",X"F0",X"F0",X"F0",X"C3",X"0F",X"0C",X"00",X"00",
		X"78",X"78",X"78",X"F0",X"16",X"12",X"03",X"01",X"F9",X"E1",X"F0",X"F0",X"F0",X"F0",X"F0",X"78",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"16",X"03",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"03",X"03",X"03",X"03",X"03",X"03",X"78",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",
		X"03",X"03",X"01",X"06",X"06",X"06",X"0E",X"1E",X"E1",X"E1",X"0F",X"0E",X"00",X"00",X"0F",X"F0",
		X"0D",X"87",X"E1",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"B4",X"B4",X"B4",X"D2",X"D2",X"D2",X"E1",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"1E",X"84",X"84",X"86",X"C2",X"C2",X"C3",X"E1",X"E1",
		X"C3",X"C2",X"0E",X"0E",X"00",X"00",X"0F",X"78",X"69",X"07",X"00",X"01",X"01",X"01",X"00",X"00",
		X"3C",X"34",X"78",X"78",X"78",X"78",X"78",X"16",X"E1",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"7F",X"7F",X"0F",X"00",X"0F",X"7F",X"7F",X"EF",X"FF",X"FF",X"7F",X"7F",X"7F",X"FF",X"FF",
		X"3C",X"9E",X"CF",X"FF",X"EF",X"DE",X"BC",X"78",X"F0",X"E1",X"69",X"2D",X"E1",X"E1",X"B4",X"5A",
		X"4F",X"0E",X"00",X"00",X"00",X"01",X"03",X"00",X"3F",X"33",X"11",X"17",X"3F",X"09",X"00",X"00",
		X"AD",X"DE",X"DE",X"FF",X"FF",X"7F",X"3F",X"17",X"E1",X"F0",X"F0",X"EF",X"FF",X"FF",X"EF",X"CF",
		X"A7",X"6F",X"EF",X"EF",X"EF",X"6F",X"A7",X"E7",X"0E",X"0E",X"0F",X"0E",X"0E",X"0E",X"0C",X"0C",
		X"01",X"01",X"09",X"13",X"13",X"13",X"13",X"37",X"EF",X"EF",X"EF",X"CF",X"DF",X"DF",X"DF",X"9F",
		X"E7",X"E7",X"7F",X"FF",X"DF",X"DF",X"57",X"77",X"0F",X"E1",X"69",X"0F",X"BF",X"DF",X"EF",X"EF",
		X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"EF",X"0E",X"BF",X"BF",X"3F",X"7F",X"0F",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"37",X"13",X"01",X"00",X"00",X"00",X"00",X"00",X"CE",X"8E",X"0C",X"08",X"00",X"00",X"00",X"00",
		X"02",X"02",X"02",X"02",X"02",X"03",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"4E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"4E",X"6F",X"37",X"13",X"3F",X"FF",X"3F",X"6F",X"7F",X"7D",X"F8",X"F0",X"E1",X"D3",X"B7",
		X"27",X"6F",X"EF",X"C6",X"4E",X"CF",X"EF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",
		X"00",X"00",X"00",X"02",X"07",X"2F",X"7F",X"FF",X"00",X"00",X"00",X"00",X"00",X"0B",X"3F",X"9F",
		X"0C",X"0E",X"4F",X"7F",X"7F",X"3F",X"07",X"01",X"17",X"37",X"3F",X"FF",X"EF",X"CF",X"BC",X"8F",
		X"FF",X"FF",X"FF",X"FF",X"78",X"F0",X"C3",X"C3",X"DF",X"FF",X"FF",X"FF",X"D3",X"E1",X"3C",X"3C",
		X"13",X"07",X"27",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"3F",X"8F",X"EF",X"EF",X"CF",X"CF",
		X"FF",X"FF",X"FF",X"CF",X"AF",X"7F",X"FF",X"FF",X"8E",X"CF",X"EF",X"EF",X"4F",X"5E",X"7E",X"7E",
		X"BF",X"BF",X"AF",X"AF",X"EF",X"EF",X"E7",X"E7",X"8F",X"2D",X"69",X"0F",X"0C",X"0C",X"0E",X"0E",
		X"7F",X"3F",X"37",X"37",X"13",X"13",X"13",X"13",X"3E",X"BE",X"BE",X"BE",X"9F",X"DF",X"DF",X"CF",
		X"F6",X"F6",X"F3",X"F3",X"F9",X"FD",X"F4",X"FD",X"87",X"B4",X"B4",X"B4",X"BC",X"BC",X"BC",X"BC",
		X"78",X"78",X"78",X"78",X"5A",X"0F",X"D2",X"D2",X"F0",X"F0",X"E1",X"C3",X"1E",X"78",X"69",X"69",
		X"F9",X"F3",X"F3",X"F6",X"F6",X"FC",X"8F",X"BC",X"BC",X"B4",X"B4",X"B4",X"B4",X"B4",X"0F",X"F0",
		X"D2",X"0F",X"5A",X"78",X"78",X"78",X"3C",X"B4",X"69",X"69",X"78",X"C3",X"E1",X"F0",X"F0",X"F0",
		X"87",X"3C",X"78",X"F0",X"F0",X"3C",X"D2",X"D2",X"0E",X"0F",X"E1",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"0C",X"0F",X"C3",X"F0",X"F0",X"F0",X"F0",X"00",X"03",X"0F",X"0F",X"C3",X"C3",X"C3",X"C3",
		X"D2",X"0F",X"F0",X"F0",X"78",X"3C",X"87",X"D2",X"F0",X"78",X"F0",X"F0",X"E1",X"0F",X"1E",X"F0",
		X"F0",X"F0",X"F0",X"C3",X"0F",X"0C",X"FF",X"FF",X"C3",X"C3",X"C3",X"0F",X"0F",X"03",X"CC",X"CF",
		X"BC",X"3C",X"B4",X"B4",X"D2",X"E1",X"D2",X"D2",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"3C",X"B4",
		X"B4",X"B4",X"B4",X"B4",X"D2",X"1E",X"84",X"C2",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"3C",X"16",
		X"F0",X"F0",X"F0",X"78",X"3C",X"16",X"03",X"00",X"87",X"F0",X"E1",X"E1",X"C3",X"C2",X"0E",X"00",
		X"0E",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E1",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"0F",X"0B",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"9D",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",
		X"C3",X"0E",X"0C",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"4F",X"4F",X"07",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"09",X"CF",X"EF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"0B",X"00",X"00",X"01",X"03",X"16",X"3C",X"78",X"F0",
		X"01",X"00",X"00",X"00",X"07",X"3F",X"17",X"03",X"7F",X"7F",X"7F",X"77",X"3F",X"FF",X"FF",X"FF",
		X"0E",X"8F",X"CF",X"EF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"08",X"0C",X"0E",X"8F",X"CE",X"0C",
		X"07",X"2D",X"78",X"F0",X"F0",X"F0",X"F0",X"D2",X"7F",X"7F",X"3F",X"B7",X"86",X"C2",X"C0",X"80",
		X"EF",X"CF",X"8E",X"0C",X"08",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"E9",X"CF",X"9F",X"3F",X"FF",X"FF",X"FF",X"6F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EF",X"CF",X"8F",X"FF",X"FF",X"EF",X"CF",X"EF",X"FF",X"FF",X"3F",X"9F",X"3F",X"7F",X"FF",X"7F",
		X"FF",X"FF",X"FF",X"FF",X"3F",X"0F",X"02",X"02",X"EF",X"CF",X"9F",X"3F",X"FF",X"7F",X"0F",X"00",
		X"3F",X"CF",X"FF",X"FF",X"FF",X"FF",X"0F",X"25",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",
		X"97",X"3F",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"0F",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"0F",X"0F",X"CE",X"CE",X"CE",X"EF",X"EF",X"EF",X"6F",X"2F",X"07",X"03",X"00",
		X"0E",X"0F",X"01",X"01",X"01",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"34",X"34",X"16",X"03",X"00",X"00",X"00",X"00",X"87",X"C3",X"0C",X"01",X"01",X"12",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"7F",X"3F",X"97",X"D3",X"C3",X"69",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"CE",X"CE",X"CE",X"CE",X"CE",X"8E",X"8C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"25",X"69",X"25",X"03",X"01",X"00",X"FF",X"EF",X"EF",X"CF",X"8E",X"8C",X"0C",X"00",
		X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"37",X"07",X"01",X"00",X"00",X"00",X"00",
		X"0F",X"FF",X"FF",X"7F",X"0F",X"00",X"00",X"00",X"0F",X"FF",X"FF",X"FF",X"3F",X"37",X"37",X"37",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0E",X"EF",X"EF",X"CF",X"8E",X"8C",X"8C",X"8C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"0F",X"B4",X"B4",X"B4",X"B4",X"96",X"0F",X"0F",X"D2",X"D2",X"C3",X"E1",X"E1",X"E1",
		X"0F",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"3F",X"1F",X"87",X"A5",X"B4",X"B4",X"3C",X"78",
		X"D2",X"D2",X"D2",X"F0",X"F0",X"F0",X"F0",X"F0",X"E1",X"E1",X"F0",X"F0",X"F0",X"1E",X"4F",X"6F",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"87",X"78",X"78",X"78",X"78",X"78",X"F0",X"F0",X"F0",
		X"FF",X"FF",X"3F",X"0F",X"A5",X"B4",X"B4",X"B4",X"FF",X"FF",X"FF",X"7F",X"3F",X"1F",X"C3",X"E1",
		X"8C",X"8C",X"8C",X"8C",X"8C",X"8C",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3C",X"78",X"78",X"78",X"F0",X"F0",X"E1",X"C3",X"F0",X"F0",X"F0",X"D2",X"97",X"3F",X"7F",X"FF",
		X"08",X"08",X"08",X"00",X"0D",X"8F",X"CF",X"EF",X"07",X"27",X"27",X"2F",X"6F",X"EF",X"EF",X"EF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"30",X"30",X"30",X"30",X"30",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"D0",X"00",X"00",X"00",X"00",X"10",X"70",X"60",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"30",X"30",X"30",X"30",X"30",X"30",X"00",X"0F",
		X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"60",X"60",X"30",X"00",X"00",X"00",X"00",X"00",
		X"00",X"30",X"70",X"F0",X"F0",X"30",X"D0",X"D0",X"00",X"00",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"C0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"C0",
		X"D0",X"00",X"F0",X"F0",X"70",X"30",X"00",X"00",X"F0",X"70",X"F0",X"F0",X"E0",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"C0",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"03",X"03",
		X"08",X"08",X"08",X"08",X"0C",X"00",X"08",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"13",X"37",X"7F",X"EF",
		X"00",X"00",X"00",X"0B",X"CE",X"CE",X"0F",X"00",X"00",X"00",X"00",X"0D",X"13",X"13",X"0F",X"00",
		X"13",X"37",X"7F",X"6F",X"6F",X"6F",X"6F",X"6F",X"CE",X"8C",X"08",X"01",X"12",X"12",X"12",X"12",
		X"00",X"07",X"78",X"F0",X"F0",X"0F",X"0F",X"F0",X"00",X"0C",X"C2",X"E1",X"E1",X"E1",X"E1",X"E1",
		X"00",X"00",X"00",X"0C",X"8F",X"EF",X"7F",X"7F",X"00",X"0E",X"69",X"34",X"12",X"3C",X"2D",X"8E",
		X"00",X"00",X"00",X"08",X"84",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"08",
		X"37",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"CF",X"EF",X"EF",X"EF",X"EE",X"8F",X"BC",X"BC",
		X"01",X"02",X"04",X"00",X"01",X"00",X"08",X"84",X"01",X"02",X"04",X"08",X"00",X"00",X"00",X"00",
		X"6F",X"6F",X"6F",X"6F",X"6F",X"6F",X"6F",X"6F",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"12",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"C3",X"A5",X"E1",X"C2",X"84",X"84",X"84",X"84",X"C2",X"E1",
		X"6F",X"27",X"03",X"01",X"00",X"00",X"00",X"00",X"12",X"01",X"00",X"08",X"0C",X"06",X"02",X"00",
		X"E1",X"F0",X"78",X"07",X"00",X"00",X"0F",X"0F",X"E1",X"E1",X"E1",X"0E",X"00",X"00",X"0F",X"0F",
		X"13",X"13",X"37",X"7F",X"7F",X"7F",X"37",X"13",X"DE",X"EF",X"DE",X"BC",X"DE",X"EF",X"0E",X"69",
		X"C2",X"E1",X"C2",X"84",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"13",X"13",X"13",X"13",X"17",X"3F",X"6F",X"02",X"78",X"BC",X"DE",X"BC",X"78",X"2D",X"02",X"00",
		X"08",X"84",X"C2",X"84",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"11",X"11",
		X"00",X"00",X"88",X"88",X"CC",X"CC",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"11",X"11",X"11",X"33",X"33",
		X"EE",X"EE",X"66",X"CC",X"CC",X"CC",X"CC",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"08",X"08",X"08",X"0C",X"0C",X"0C",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"06",X"00",X"06",X"02",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"07",X"00",X"00",X"07",X"0F",X"0F",X"17",X"1B",X"3F",
		X"00",X"00",X"0C",X"0E",X"1E",X"0D",X"0B",X"8F",X"00",X"00",X"00",X"00",X"C0",X"38",X"0C",X"0C",
		X"07",X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"FF",X"3F",X"1B",X"17",X"0F",X"0F",X"07",X"00",
		X"EF",X"8F",X"0B",X"0D",X"0E",X"0E",X"0C",X"00",X"0C",X"0C",X"0C",X"08",X"00",X"00",X"00",X"00",
		X"00",X"30",X"70",X"80",X"00",X"80",X"40",X"30",X"00",X"C0",X"E0",X"E0",X"60",X"20",X"10",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"30",X"30",X"70",X"40",X"00",X"E0",X"40",X"C0",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"33",X"77",X"77",X"00",X"00",X"77",X"FF",X"FF",X"67",X"AB",X"CF",
		X"00",X"00",X"CC",X"EE",X"FE",X"DD",X"BB",X"7F",X"00",X"00",X"00",X"00",X"E0",X"98",X"CC",X"CC",
		X"77",X"77",X"77",X"33",X"00",X"00",X"00",X"00",X"0F",X"CF",X"AB",X"67",X"FF",X"FF",X"77",X"00",
		X"1F",X"7F",X"BB",X"DD",X"EE",X"EE",X"CC",X"00",X"CC",X"CC",X"CC",X"88",X"00",X"00",X"00",X"00",
		X"00",X"30",X"70",X"F0",X"00",X"80",X"40",X"30",X"00",X"C0",X"E0",X"E0",X"E0",X"60",X"10",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"30",X"70",X"70",X"E0",X"00",X"F0",X"20",X"E0",X"C0",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
