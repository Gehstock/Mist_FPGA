library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ckong_tile_bit0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ckong_tile_bit0 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3C",X"7E",X"FF",X"FF",X"FF",X"FF",X"7E",X"3C",X"3C",X"7F",X"E7",X"C3",X"C3",X"E7",X"7E",X"3C",
		X"3C",X"42",X"81",X"81",X"81",X"81",X"42",X"3C",X"3C",X"42",X"99",X"BD",X"BD",X"99",X"42",X"3C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"3F",X"3F",X"3F",X"3C",X"30",X"00",X"00",X"30",X"30",X"30",X"30",X"30",X"30",X"00",X"00",
		X"0C",X"0C",X"0C",X"0C",X"0C",X"00",X"00",X"00",X"03",X"03",X"03",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"30",X"3C",X"3F",X"3F",X"3F",X"3F",X"00",X"00",X"30",X"30",X"30",X"30",X"30",X"30",
		X"00",X"00",X"00",X"0C",X"0C",X"0C",X"0C",X"0C",X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"03",
		X"00",X"00",X"3F",X"3F",X"1F",X"1F",X"0F",X"0F",X"00",X"00",X"3F",X"3F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"1F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",
		X"00",X"00",X"FC",X"FC",X"F8",X"F8",X"F0",X"F0",X"00",X"00",X"FC",X"FC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F8",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",
		X"00",X"00",X"0C",X"3C",X"FC",X"FC",X"FC",X"FC",X"00",X"00",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"00",X"00",X"00",X"30",X"30",X"30",X"30",X"30",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7B",X"7B",X"00",X"00",X"00",X"00",
		X"FC",X"FC",X"FC",X"FC",X"3C",X"0C",X"00",X"00",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"00",X"00",
		X"30",X"30",X"30",X"30",X"30",X"00",X"00",X"00",X"47",X"25",X"17",X"08",X"74",X"52",X"71",X"00",
		X"C0",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F8",X"F8",X"FC",X"FC",X"00",X"00",
		X"00",X"00",X"41",X"22",X"1C",X"00",X"00",X"00",X"00",X"00",X"3C",X"42",X"81",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FC",X"FC",X"00",X"00",X"00",X"00",X"08",X"1C",X"08",X"00",X"00",X"00",
		X"00",X"00",X"06",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"00",X"00",X"00",
		X"00",X"00",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"F8",X"00",X"00",X"00",X"00",
		X"1C",X"3E",X"61",X"41",X"43",X"3E",X"1C",X"00",X"01",X"01",X"7F",X"7F",X"21",X"01",X"00",X"00",
		X"31",X"79",X"5D",X"4D",X"4F",X"67",X"23",X"00",X"46",X"6F",X"79",X"59",X"49",X"43",X"02",X"00",
		X"04",X"7F",X"7F",X"64",X"34",X"1C",X"0C",X"00",X"0E",X"5F",X"51",X"51",X"51",X"73",X"72",X"00",
		X"06",X"4F",X"49",X"49",X"69",X"3F",X"1E",X"00",X"60",X"70",X"59",X"4F",X"47",X"61",X"60",X"00",
		X"06",X"37",X"4F",X"4D",X"5D",X"79",X"36",X"00",X"3C",X"7E",X"4B",X"49",X"49",X"79",X"30",X"00",
		X"00",X"00",X"33",X"33",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"1F",X"1F",X"3F",X"3F",X"00",X"00",X"00",X"00",X"14",X"14",X"14",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"3F",X"3F",X"00",X"00",X"00",X"00",X"1F",X"1F",X"00",X"00",X"00",X"00",
		X"3C",X"42",X"81",X"A5",X"A5",X"99",X"42",X"3C",X"1F",X"3F",X"64",X"44",X"64",X"3F",X"1F",X"00",
		X"36",X"7F",X"49",X"49",X"7F",X"7F",X"00",X"00",X"63",X"41",X"41",X"63",X"3E",X"1C",X"00",X"00",
		X"1C",X"3E",X"63",X"41",X"41",X"7F",X"7F",X"00",X"41",X"49",X"49",X"49",X"7F",X"7F",X"00",X"00",
		X"40",X"48",X"48",X"48",X"7F",X"7F",X"00",X"00",X"4F",X"4F",X"49",X"41",X"63",X"3E",X"1C",X"00",
		X"7F",X"7F",X"08",X"08",X"08",X"7F",X"7F",X"00",X"00",X"41",X"41",X"7F",X"7F",X"41",X"41",X"00",
		X"7E",X"7F",X"01",X"01",X"01",X"03",X"02",X"00",X"41",X"63",X"37",X"1E",X"0C",X"7F",X"7F",X"00",
		X"01",X"01",X"01",X"01",X"01",X"7F",X"7F",X"00",X"7F",X"7F",X"38",X"1C",X"38",X"7F",X"7F",X"00",
		X"7F",X"7F",X"0E",X"1C",X"38",X"7F",X"7F",X"00",X"3E",X"7F",X"41",X"41",X"41",X"7F",X"3E",X"00",
		X"38",X"7C",X"44",X"44",X"44",X"7F",X"7F",X"00",X"3D",X"7E",X"47",X"47",X"43",X"7F",X"3E",X"00",
		X"39",X"7B",X"5F",X"4E",X"4C",X"7F",X"7F",X"00",X"06",X"2F",X"69",X"49",X"49",X"7B",X"32",X"00",
		X"40",X"40",X"7F",X"7F",X"40",X"40",X"00",X"00",X"7E",X"7F",X"01",X"01",X"01",X"7F",X"7E",X"00",
		X"78",X"7C",X"0E",X"07",X"0E",X"7C",X"78",X"00",X"7C",X"7F",X"0E",X"1C",X"0E",X"7F",X"7C",X"00",
		X"63",X"77",X"3E",X"1C",X"3E",X"77",X"63",X"00",X"60",X"78",X"1F",X"1F",X"78",X"60",X"00",X"00",
		X"61",X"71",X"79",X"5D",X"4F",X"47",X"43",X"00",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"F0",X"C1",X"01",X"03",X"03",X"07",X"07",X"07",X"07",X"03",X"03",X"01",X"C1",X"F0",X"FC",
		X"E0",X"E0",X"C0",X"C0",X"80",X"83",X"0F",X"3F",X"3F",X"0F",X"83",X"80",X"C0",X"C0",X"E0",X"E0",
		X"C0",X"C0",X"C0",X"00",X"00",X"00",X"07",X"07",X"30",X"30",X"00",X"00",X"03",X"03",X"00",X"00",
		X"C0",X"C0",X"E0",X"60",X"70",X"3C",X"1F",X"07",X"07",X"1F",X"3C",X"70",X"60",X"E0",X"C0",X"C0",
		X"03",X"03",X"07",X"06",X"0E",X"3C",X"F8",X"E0",X"E0",X"F8",X"3C",X"0E",X"06",X"07",X"03",X"03",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"FF",X"FF",X"FF",X"FF",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"03",X"03",X"03",X"03",X"03",X"03",X"FF",X"FF",X"FF",X"FF",X"03",X"03",X"03",X"03",X"03",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",
		X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"00",X"00",X"18",X"3C",X"3C",X"18",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FC",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"7E",X"7C",X"78",X"70",X"70",X"70",X"70",X"70",
		X"1E",X"3C",X"38",X"30",X"30",X"30",X"30",X"30",X"06",X"0C",X"18",X"10",X"10",X"10",X"10",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"0F",X"1F",X"3F",X"7F",X"FF",
		X"00",X"00",X"01",X"03",X"07",X"0F",X"1F",X"3F",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"F2",X"FF",X"FF",X"E0",X"C0",X"80",X"00",X"00",X"FF",X"FF",X"FF",X"E0",X"C0",X"80",X"00",
		X"00",X"00",X"7F",X"FF",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"3F",X"60",X"C0",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"07",X"03",X"01",X"00",X"00",X"FF",X"FF",X"FF",X"07",X"03",X"01",X"00",
		X"00",X"00",X"FE",X"FF",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"DC",X"06",X"03",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"F0",X"F8",X"FC",X"FE",X"FF",
		X"00",X"00",X"80",X"C0",X"E0",X"F0",X"F8",X"FC",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"3F",X"1F",X"0F",X"0F",X"0F",X"0F",X"0F",X"7E",X"3E",X"1E",X"0E",X"0E",X"08",X"0E",X"0E",
		X"78",X"3C",X"1C",X"0C",X"0C",X"0C",X"0C",X"0C",X"60",X"30",X"18",X"08",X"08",X"08",X"08",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",X"3F",X"7F",X"0E",X"0E",X"0E",X"0E",X"0E",X"1E",X"3E",X"7E",
		X"0C",X"0C",X"0C",X"0C",X"0C",X"1C",X"3C",X"78",X"08",X"08",X"08",X"08",X"08",X"18",X"30",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FE",X"FC",X"F8",X"F0",X"E0",X"C0",X"80",
		X"FC",X"58",X"B0",X"E0",X"C0",X"80",X"00",X"00",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"07",X"FF",X"FF",X"FF",X"FF",X"00",X"01",X"03",X"07",X"FF",X"FF",X"FF",X"00",
		X"00",X"01",X"03",X"07",X"FF",X"FE",X"00",X"00",X"00",X"01",X"03",X"06",X"FC",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"C0",X"E0",X"FF",X"FF",X"FF",X"FF",X"00",X"80",X"C0",X"E0",X"FF",X"FF",X"FF",X"00",
		X"00",X"80",X"C0",X"E0",X"FF",X"7F",X"00",X"00",X"00",X"80",X"C0",X"60",X"3F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"7F",X"3F",X"1F",X"0F",X"07",X"03",X"01",
		X"3F",X"1F",X"0F",X"07",X"03",X"01",X"00",X"00",X"0F",X"07",X"03",X"01",X"00",X"00",X"00",X"00",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"FC",X"FE",X"70",X"70",X"70",X"70",X"70",X"78",X"7C",X"7E",
		X"30",X"30",X"30",X"30",X"30",X"38",X"3C",X"1E",X"10",X"10",X"10",X"10",X"10",X"18",X"0C",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"5A",X"3C",X"FF",X"FF",X"3C",X"5A",X"99",
		X"0C",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"07",X"07",X"00",X"00",X"00",X"C0",X"C0",X"C0",
		X"00",X"00",X"03",X"03",X"00",X"00",X"30",X"30",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"0C",
		X"E0",X"E0",X"00",X"00",X"00",X"03",X"03",X"03",X"00",X"00",X"C0",X"C0",X"00",X"00",X"0C",X"0C",
		X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"30",X"03",X"03",X"03",X"00",X"00",X"00",X"E0",X"E0",
		X"0C",X"0C",X"00",X"00",X"C0",X"C0",X"00",X"00",X"30",X"00",X"80",X"80",X"00",X"00",X"00",X"00",
		X"F9",X"E2",X"84",X"09",X"11",X"23",X"43",X"87",X"87",X"43",X"23",X"11",X"09",X"84",X"E2",X"F9",
		X"87",X"43",X"23",X"91",X"89",X"C4",X"C2",X"E1",X"E1",X"C2",X"C4",X"88",X"90",X"21",X"47",X"9F",
		X"F3",X"C7",X"8E",X"0C",X"11",X"21",X"43",X"87",X"87",X"43",X"21",X"11",X"0C",X"8E",X"C7",X"F3",
		X"CF",X"E3",X"71",X"30",X"88",X"84",X"C2",X"E1",X"E1",X"C2",X"84",X"88",X"30",X"71",X"E3",X"CF",
		X"E7",X"CF",X"8F",X"1E",X"38",X"31",X"43",X"87",X"87",X"43",X"31",X"38",X"1E",X"8F",X"CF",X"E7",
		X"E7",X"F3",X"F1",X"78",X"1C",X"8C",X"C2",X"E1",X"E1",X"C2",X"8C",X"1C",X"78",X"F1",X"F3",X"E7",
		X"EF",X"DF",X"9F",X"3F",X"3E",X"79",X"63",X"87",X"87",X"63",X"79",X"3E",X"3F",X"9F",X"DF",X"EF",
		X"F7",X"FB",X"F9",X"FC",X"7C",X"9E",X"C6",X"E1",X"E1",X"C6",X"9E",X"7C",X"FC",X"F9",X"FB",X"F7",
		X"DF",X"FF",X"BF",X"3F",X"7F",X"7E",X"73",X"87",X"87",X"73",X"7E",X"7F",X"3F",X"BF",X"FF",X"DF",
		X"FB",X"FF",X"FD",X"FC",X"FE",X"7E",X"CE",X"E1",X"E1",X"CE",X"7E",X"FE",X"FC",X"FD",X"FF",X"FB",
		X"BF",X"BF",X"3F",X"7F",X"7F",X"7F",X"78",X"83",X"83",X"78",X"7F",X"7F",X"7F",X"3F",X"BF",X"BF",
		X"FD",X"FD",X"FC",X"FE",X"FE",X"FE",X"1E",X"C1",X"C1",X"1E",X"FE",X"FE",X"FE",X"FC",X"FD",X"FD",
		X"18",X"18",X"0C",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0F",X"0C",X"18",X"18",
		X"18",X"18",X"30",X"F0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"F0",X"30",X"18",X"18",
		X"7F",X"1F",X"7F",X"0F",X"17",X"25",X"05",X"01",X"01",X"05",X"25",X"17",X"1F",X"7F",X"1F",X"FF",
		X"FF",X"F8",X"FE",X"F0",X"E8",X"A4",X"A0",X"80",X"80",X"A0",X"A4",X"E8",X"F0",X"FE",X"F8",X"FF",
		X"01",X"02",X"04",X"00",X"00",X"00",X"00",X"00",X"FF",X"01",X"0F",X"FF",X"01",X"07",X"1F",X"38",
		X"39",X"1F",X"07",X"01",X"FF",X"0F",X"01",X"FF",X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"01",
		X"7F",X"6D",X"6D",X"CD",X"C9",X"89",X"09",X"09",X"09",X"09",X"89",X"C9",X"CD",X"6D",X"6D",X"7F",
		X"FE",X"B6",X"B6",X"B3",X"93",X"91",X"90",X"90",X"90",X"90",X"91",X"93",X"B3",X"B6",X"B6",X"FE",
		X"80",X"40",X"20",X"00",X"00",X"00",X"00",X"00",X"FF",X"80",X"F0",X"FF",X"80",X"E0",X"F8",X"1C",
		X"1C",X"F8",X"E0",X"80",X"FF",X"F0",X"80",X"FF",X"00",X"00",X"00",X"00",X"00",X"20",X"40",X"80",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"01",X"02",X"02",X"01",X"00",X"00",
		X"00",X"03",X"04",X"08",X"08",X"04",X"03",X"00",X"00",X"0F",X"10",X"20",X"20",X"10",X"0F",X"00",
		X"00",X"3F",X"40",X"80",X"80",X"40",X"3F",X"00",X"99",X"95",X"B1",X"75",X"29",X"92",X"41",X"59",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C1",X"F1",X"7B",X"3B",X"3F",X"0F",X"3F",X"FF",X"83",X"8F",X"DE",X"DC",X"FC",X"F0",X"FC",X"FF",
		X"FF",X"3F",X"0F",X"3F",X"7B",X"7B",X"F1",X"C1",X"FF",X"FC",X"F0",X"FC",X"DE",X"DE",X"8F",X"83",
		X"07",X"1F",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"E0",X"F8",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",X"1F",X"07",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"F8",X"E0",
		X"E0",X"E0",X"E1",X"E7",X"EC",X"ED",X"FC",X"FF",X"00",X"00",X"E0",X"F8",X"FC",X"7C",X"FE",X"FE",
		X"FF",X"FC",X"ED",X"EC",X"E7",X"E1",X"E0",X"E0",X"FE",X"FE",X"7C",X"FC",X"F8",X"E0",X"00",X"00",
		X"E0",X"E0",X"E1",X"E7",X"EC",X"ED",X"FC",X"FF",X"00",X"00",X"E0",X"F8",X"FC",X"7C",X"FE",X"FE",
		X"FF",X"FC",X"ED",X"EC",X"E7",X"E1",X"E0",X"E0",X"FE",X"FE",X"7C",X"FC",X"F8",X"E0",X"00",X"00",
		X"E0",X"E0",X"E1",X"E7",X"EC",X"ED",X"FC",X"FF",X"00",X"00",X"E0",X"F8",X"FC",X"7C",X"FE",X"FE",
		X"FF",X"FC",X"ED",X"EC",X"E7",X"E1",X"E0",X"E0",X"FE",X"FE",X"7C",X"FC",X"F8",X"E0",X"00",X"00",
		X"E0",X"E0",X"E0",X"E0",X"E8",X"EC",X"FE",X"FF",X"00",X"00",X"00",X"00",X"04",X"0C",X"1E",X"3E",
		X"FF",X"FD",X"EC",X"EF",X"E7",X"E1",X"E0",X"E0",X"FE",X"7E",X"FC",X"FC",X"F8",X"E0",X"00",X"00",
		X"E0",X"E0",X"E0",X"E6",X"EE",X"EF",X"FF",X"FF",X"00",X"00",X"20",X"38",X"3C",X"3C",X"3E",X"BE",
		X"FF",X"FD",X"EC",X"EF",X"E7",X"E1",X"E0",X"E0",X"FE",X"7E",X"FC",X"FC",X"F8",X"E0",X"00",X"00",
		X"E0",X"E0",X"E1",X"E7",X"EC",X"ED",X"FC",X"FF",X"00",X"00",X"E0",X"F8",X"FC",X"7C",X"FE",X"FE",
		X"FF",X"FC",X"ED",X"EC",X"E7",X"E1",X"E0",X"E0",X"FE",X"FE",X"7C",X"FC",X"F8",X"E0",X"00",X"00",
		X"00",X"00",X"E1",X"E7",X"EC",X"ED",X"FC",X"FF",X"00",X"00",X"E0",X"F8",X"FC",X"7C",X"FE",X"FE",
		X"FF",X"FC",X"ED",X"EC",X"E7",X"E1",X"00",X"00",X"FE",X"FE",X"7C",X"FC",X"F8",X"E0",X"00",X"00",
		X"00",X"00",X"E1",X"E7",X"EC",X"ED",X"FC",X"FF",X"00",X"00",X"E0",X"F8",X"FC",X"7C",X"FE",X"FE",
		X"FF",X"FC",X"ED",X"EC",X"E7",X"E1",X"00",X"00",X"FE",X"FE",X"7C",X"FC",X"F8",X"E0",X"00",X"00",
		X"00",X"00",X"E1",X"E7",X"EC",X"ED",X"FC",X"FF",X"00",X"00",X"E0",X"F8",X"FC",X"7C",X"FE",X"FE",
		X"FF",X"FC",X"ED",X"EC",X"E7",X"E1",X"00",X"00",X"FE",X"FE",X"7C",X"FC",X"F8",X"E0",X"00",X"00",
		X"00",X"00",X"E0",X"E0",X"E8",X"EC",X"FE",X"FF",X"00",X"00",X"00",X"00",X"04",X"0C",X"1E",X"3E",
		X"FF",X"FD",X"EC",X"EF",X"E7",X"E1",X"00",X"00",X"FE",X"7E",X"FC",X"FC",X"F8",X"E0",X"00",X"00",
		X"00",X"00",X"E0",X"E6",X"EE",X"EF",X"FF",X"FF",X"00",X"00",X"20",X"38",X"3C",X"3C",X"3E",X"BE",
		X"FF",X"FD",X"EC",X"EF",X"E7",X"E1",X"00",X"00",X"FE",X"7E",X"FC",X"FC",X"F8",X"E0",X"00",X"00",
		X"00",X"00",X"E1",X"E7",X"EC",X"ED",X"FC",X"FF",X"00",X"00",X"E0",X"F8",X"FC",X"7C",X"FE",X"FE",
		X"FF",X"FC",X"ED",X"EC",X"E7",X"E1",X"00",X"00",X"FE",X"FE",X"7C",X"FC",X"F8",X"E0",X"00",X"00",
		X"00",X"00",X"01",X"07",X"EC",X"ED",X"FC",X"FF",X"00",X"00",X"E0",X"F8",X"FC",X"7C",X"FE",X"FE",
		X"FF",X"FC",X"ED",X"EC",X"07",X"01",X"00",X"00",X"FE",X"FE",X"7C",X"FC",X"F8",X"E0",X"00",X"00",
		X"00",X"00",X"01",X"07",X"EC",X"ED",X"FC",X"FF",X"00",X"00",X"E0",X"F8",X"FC",X"7C",X"FE",X"FE",
		X"FF",X"FC",X"ED",X"EC",X"07",X"01",X"00",X"00",X"FE",X"FE",X"7C",X"FC",X"F8",X"E0",X"00",X"00",
		X"00",X"00",X"01",X"07",X"EC",X"ED",X"FC",X"FF",X"00",X"00",X"E0",X"F8",X"FC",X"7C",X"FE",X"FE",
		X"FF",X"FC",X"ED",X"EC",X"07",X"01",X"00",X"00",X"FE",X"FE",X"7C",X"FC",X"F8",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"E8",X"EC",X"FE",X"FF",X"00",X"00",X"00",X"00",X"04",X"0C",X"1E",X"3E",
		X"FF",X"FD",X"EC",X"EF",X"07",X"01",X"00",X"00",X"FE",X"7E",X"FC",X"FC",X"F8",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"06",X"EE",X"EF",X"FF",X"FF",X"00",X"00",X"20",X"38",X"3C",X"3C",X"3E",X"BE",
		X"FF",X"FD",X"EC",X"EF",X"07",X"01",X"00",X"00",X"FE",X"7E",X"FC",X"FC",X"F8",X"E0",X"00",X"00",
		X"00",X"00",X"01",X"07",X"EC",X"ED",X"FC",X"FF",X"00",X"00",X"E0",X"F8",X"FC",X"7C",X"FE",X"FE",
		X"FF",X"FC",X"ED",X"EC",X"07",X"01",X"00",X"00",X"FE",X"FE",X"7C",X"FC",X"F8",X"E0",X"00",X"00",
		X"00",X"00",X"01",X"07",X"2C",X"0D",X"00",X"00",X"00",X"00",X"E0",X"F8",X"FC",X"7C",X"FE",X"FE",
		X"00",X"00",X"2D",X"0C",X"07",X"01",X"00",X"00",X"FE",X"FE",X"7C",X"FC",X"F8",X"E0",X"00",X"00",
		X"00",X"00",X"01",X"07",X"04",X"01",X"00",X"00",X"00",X"00",X"E0",X"F8",X"FC",X"7C",X"FE",X"FE",
		X"00",X"00",X"01",X"04",X"07",X"01",X"00",X"00",X"FE",X"FE",X"7C",X"FC",X"F8",X"E0",X"00",X"00",
		X"00",X"00",X"01",X"03",X"00",X"01",X"00",X"00",X"00",X"00",X"E0",X"F8",X"FC",X"7C",X"FE",X"FE",
		X"00",X"00",X"01",X"00",X"03",X"01",X"00",X"00",X"FE",X"FE",X"7C",X"FC",X"F8",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"F8",X"FC",X"7C",X"FE",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FE",X"7C",X"FC",X"F8",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"38",X"7C",X"7C",X"FE",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FE",X"7C",X"7C",X"38",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"1C",X"3C",X"7E",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"7E",X"3C",X"1C",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"3E",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"3E",X"0C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"12",X"08",X"00",X"30",X"00",X"00",X"80",X"90",X"20",X"08",X"10",X"00",
		X"00",X"08",X"10",X"04",X"09",X"01",X"00",X"00",X"0C",X"00",X"10",X"48",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"07",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",
		X"06",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",
		X"05",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"08",X"08",X"1D",X"1E",X"5F",X"7F",X"3F",X"EF",X"50",X"F0",X"E0",X"E0",X"C0",X"80",X"80",X"80",
		X"FF",X"7B",X"FF",X"7F",X"1E",X"19",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"C8",X"78",X"10",
		X"03",X"07",X"07",X"2E",X"1F",X"3F",X"5F",X"FB",X"08",X"98",X"B8",X"F8",X"F0",X"E0",X"C0",X"F0",
		X"57",X"07",X"3C",X"38",X"71",X"61",X"C3",X"01",X"F8",X"BC",X"F0",X"F8",X"FC",X"7E",X"37",X"12",
		X"00",X"03",X"0C",X"0C",X"03",X"00",X"03",X"0C",X"00",X"C0",X"30",X"30",X"C0",X"00",X"C0",X"30",
		X"0C",X"03",X"00",X"03",X"0C",X"0C",X"02",X"00",X"30",X"C0",X"00",X"30",X"B0",X"70",X"30",X"00",
		X"00",X"00",X"01",X"03",X"07",X"07",X"0F",X"0F",X"70",X"F0",X"E0",X"E0",X"FE",X"E2",X"E0",X"E0",
		X"1F",X"1B",X"15",X"11",X"1F",X"1F",X"0F",X"03",X"E0",X"E0",X"20",X"20",X"3E",X"22",X"20",X"20",
		X"00",X"00",X"01",X"03",X"07",X"07",X"0F",X"0F",X"70",X"F0",X"E0",X"E6",X"FA",X"E6",X"E2",X"E0",
		X"1F",X"1B",X"15",X"11",X"1F",X"1E",X"0E",X"04",X"E0",X"E0",X"20",X"26",X"3A",X"26",X"22",X"20",
		X"00",X"00",X"01",X"03",X"07",X"07",X"0F",X"0F",X"70",X"F0",X"E6",X"EA",X"F0",X"E8",X"E6",X"E2",
		X"1F",X"37",X"2A",X"22",X"3E",X"3C",X"18",X"08",X"E0",X"E0",X"26",X"2A",X"30",X"28",X"26",X"22",
		X"00",X"00",X"01",X"07",X"0F",X"3F",X"3F",X"77",X"70",X"F0",X"EC",X"E8",X"F0",X"E8",X"E6",X"E2",
		X"6B",X"63",X"6F",X"6E",X"28",X"00",X"00",X"00",X"E0",X"EC",X"28",X"28",X"30",X"28",X"26",X"22",
		X"00",X"0F",X"00",X"1F",X"50",X"50",X"50",X"50",X"00",X"F0",X"00",X"F8",X"0A",X"0A",X"0A",X"0A",
		X"50",X"50",X"50",X"50",X"1F",X"00",X"0F",X"00",X"0A",X"0A",X"0A",X"0A",X"F8",X"00",X"F0",X"00",
		X"4D",X"D6",X"B8",X"38",X"2A",X"44",X"77",X"DC",X"71",X"2D",X"E9",X"41",X"DE",X"EB",X"3A",X"2A",
		X"18",X"D5",X"6D",X"18",X"34",X"A1",X"40",X"69",X"3E",X"A4",X"45",X"DE",X"86",X"4D",X"D6",X"B1",
		X"AC",X"47",X"DE",X"EF",X"52",X"E4",X"37",X"22",X"56",X"77",X"A7",X"4D",X"72",X"28",X"D4",X"73",
		X"75",X"D1",X"86",X"F0",X"DF",X"3A",X"54",X"A7",X"9D",X"25",X"4B",X"7A",X"9C",X"E7",X"1A",X"24",
		X"17",X"F5",X"02",X"98",X"25",X"6E",X"70",X"D2",X"FC",X"77",X"22",X"04",X"77",X"DA",X"34",X"57",
		X"72",X"A4",X"47",X"7D",X"D1",X"E6",X"3D",X"34",X"7D",X"D3",X"95",X"5A",X"84",X"17",X"12",X"F3",
		X"40",X"70",X"8A",X"D3",X"D7",X"4D",X"7E",X"03",X"37",X"25",X"38",X"78",X"6E",X"F3",X"E6",X"0C",
		X"5A",X"8F",X"57",X"E1",X"E0",X"D7",X"35",X"5E",X"08",X"89",X"AE",X"1F",X"78",X"C5",X"5D",X"03",
		X"9F",X"27",X"6D",X"72",X"3F",X"A7",X"47",X"A8",X"34",X"5A",X"66",X"37",X"CD",X"4B",X"78",X"D5",
		X"8C",X"CB",X"1D",X"02",X"D1",X"77",X"5E",X"B8",X"24",X"F7",X"70",X"D0",X"30",X"50",X"D1",X"3D",
		X"37",X"DB",X"ED",X"3A",X"76",X"3D",X"24",X"47",X"05",X"0A",X"04",X"D7",X"9D",X"5E",X"A3",X"AF",
		X"D7",X"DD",X"B2",X"4A",X"7A",X"A4",X"63",X"72",X"14",X"71",X"9F",X"A7",X"15",X"70",X"BA",X"28",
		X"A7",X"40",X"70",X"D0",X"A9",X"6D",X"D1",X"45",X"81",X"37",X"AC",X"45",X"E9",X"4D",X"DE",X"65",
		X"8D",X"7B",X"D4",X"37",X"37",X"AD",X"62",X"73",X"31",X"3A",X"D4",X"A7",X"5D",X"E3",X"33",X"DA",
		X"AD",X"4B",X"D3",X"B5",X"3D",X"2D",X"46",X"7D",X"96",X"71",X"4D",X"19",X"A1",X"CE",X"7B",X"DA",
		X"6D",X"72",X"DA",X"BE",X"44",X"7A",X"3E",X"74",X"58",X"DF",X"BD",X"83",X"75",X"98",X"B6",X"2A",
		X"A9",X"8D",X"7B",X"76",X"D7",X"23",X"87",X"6D",X"2A",X"07",X"BB",X"D1",X"BD",X"AB",X"74",X"A7",
		X"8D",X"74",X"A3",X"4E",X"74",X"ED",X"56",X"51",X"86",X"D7",X"6E",X"14",X"98",X"D9",X"6D",X"1B",
		X"1E",X"D5",X"6A",X"14",X"37",X"7D",X"45",X"DB",X"AA",X"4D",X"76",X"A1",X"CB",X"7D",X"36",X"81",
		X"E3",X"37",X"6D",X"32",X"E8",X"39",X"67",X"33",X"DF",X"2D",X"FE",X"95",X"53",X"C0",X"D0",X"13",
		X"D8",X"A2",X"66",X"17",X"66",X"F0",X"E3",X"A3",X"56",X"71",X"6D",X"F5",X"5F",X"EF",X"0F",X"8F",
		X"75",X"0D",X"14",X"37",X"3C",X"50",X"11",X"8D",X"1D",X"6E",X"DB",X"40",X"79",X"ED",X"04",X"97",
		X"37",X"A1",X"7E",X"D3",X"A6",X"63",X"35",X"43",X"B1",X"2E",X"83",X"B6",X"B3",X"E5",X"DA",X"1F",
		X"9D",X"73",X"95",X"E1",X"38",X"75",X"8E",X"50",X"36",X"3D",X"54",X"17",X"68",X"3B",X"51",X"AD",
		X"89",X"73",X"74",X"D7",X"4F",X"70",X"00",X"B0",X"03",X"87",X"FF",X"F8",X"F1",X"FA",X"3F",X"87",
		X"0F",X"FF",X"FF",X"F0",X"F0",X"F1",X"F3",X"FF",X"F0",X"3F",X"FF",X"F0",X"00",X"00",X"0F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"85",X"1B",X"01",X"09",X"05",X"BF",X"16",X"EF",X"8F",X"7F",X"0F",X"2F",X"AF",X"99",X"55",X"21",
		X"1F",X"8F",X"0F",X"0F",X"7F",X"AF",X"FF",X"FF",X"F1",X"F2",X"F6",X"F1",X"F0",X"F0",X"F0",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
