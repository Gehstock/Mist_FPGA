library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity loc_chr_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of loc_chr_rom is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"0E",X"01",X"01",X"01",X"0F",X"0F",X"0E",X"00",X"07",X"08",X"08",X"08",X"0F",X"0F",X"07",
		X"00",X"00",X"00",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"07",X"04",X"00",
		X"00",X"01",X"09",X"0D",X"0F",X"07",X"03",X"01",X"00",X"07",X"0F",X"0F",X"08",X"08",X"08",X"06",
		X"00",X"0E",X"0F",X"0F",X"01",X"01",X"01",X"06",X"00",X"06",X"0F",X"0F",X"09",X"08",X"08",X"04",
		X"00",X"04",X"0F",X"0F",X"0F",X"04",X"04",X"0C",X"00",X"00",X"0F",X"0F",X"07",X"02",X"01",X"00",
		X"00",X"0E",X"0F",X"0F",X"01",X"01",X"02",X"02",X"00",X"08",X"09",X"09",X"09",X"09",X"09",X"0F",
		X"00",X"0E",X"01",X"01",X"01",X"0F",X"0F",X"0E",X"00",X"04",X"09",X"09",X"09",X"0F",X"0F",X"07",
		X"00",X"00",X"00",X"08",X"0F",X"0F",X"03",X"01",X"00",X"0C",X"0E",X"0F",X"0B",X"08",X"08",X"08",
		X"00",X"0E",X"0F",X"0D",X"09",X"01",X"01",X"0E",X"00",X"00",X"06",X"09",X"0B",X"0F",X"07",X"00",
		X"00",X"0E",X"0F",X"0F",X"09",X"09",X"09",X"02",X"00",X"07",X"0F",X"0F",X"08",X"08",X"08",X"07",
		X"0C",X"02",X"01",X"05",X"05",X"09",X"02",X"0C",X"03",X"04",X"08",X"0A",X"0A",X"09",X"04",X"03",
		X"0F",X"01",X"01",X"01",X"01",X"01",X"01",X"0F",X"0F",X"08",X"08",X"08",X"08",X"08",X"08",X"0F",
		X"00",X"00",X"00",X"0A",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"00",X"00",X"00",
		X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"0C",X"0E",X"0C",X"08",X"00",X"00",X"03",X"07",X"07",X"03",X"07",X"07",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"0F",X"0E",X"0A",X"02",X"0E",X"03",X"00",X"00",X"01",X"07",X"0F",X"03",X"00",X"00",
		X"00",X"0E",X"01",X"01",X"01",X"0F",X"0F",X"0F",X"00",X"06",X"09",X"09",X"09",X"0F",X"0F",X"0F",
		X"00",X"06",X"01",X"01",X"01",X"0F",X"0F",X"0E",X"00",X"04",X"08",X"08",X"08",X"0F",X"0F",X"07",
		X"00",X"0C",X"02",X"01",X"01",X"0F",X"0F",X"0F",X"00",X"03",X"04",X"08",X"08",X"0F",X"0F",X"0F",
		X"00",X"01",X"01",X"01",X"01",X"0F",X"0F",X"0F",X"00",X"09",X"09",X"09",X"09",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"00",X"09",X"09",X"09",X"09",X"0F",X"0F",X"0F",
		X"00",X"0E",X"01",X"01",X"01",X"0F",X"0F",X"0E",X"00",X"05",X"09",X"09",X"08",X"0F",X"0F",X"07",
		X"00",X"0F",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"00",X"0F",X"01",X"01",X"01",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"00",X"00",
		X"00",X"0E",X"0F",X"0F",X"01",X"01",X"01",X"02",X"00",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"03",X"0C",X"00",X"00",X"0F",X"0F",X"0F",X"00",X"08",X"04",X"03",X"02",X"0F",X"0F",X"0F",
		X"00",X"01",X"01",X"01",X"01",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",
		X"00",X"0F",X"08",X"0C",X"0E",X"0C",X"08",X"0F",X"00",X"0F",X"07",X"03",X"01",X"03",X"07",X"0F",
		X"00",X"0F",X"0F",X"0E",X"0C",X"08",X"00",X"0F",X"00",X"0F",X"00",X"01",X"03",X"07",X"0F",X"0F",
		X"00",X"0E",X"01",X"01",X"01",X"0F",X"0F",X"0E",X"00",X"07",X"08",X"08",X"08",X"0F",X"0F",X"07",
		X"00",X"08",X"04",X"04",X"04",X"0F",X"0F",X"0F",X"00",X"07",X"08",X"08",X"08",X"0F",X"0F",X"0F",
		X"00",X"0F",X"03",X"0D",X"01",X"0F",X"0F",X"0E",X"00",X"07",X"08",X"08",X"08",X"0F",X"0F",X"07",
		X"00",X"09",X"05",X"06",X"04",X"0F",X"0F",X"0F",X"00",X"07",X"08",X"08",X"08",X"0F",X"0F",X"0F",
		X"00",X"06",X"0F",X"0F",X"0F",X"09",X"01",X"02",X"00",X"04",X"08",X"09",X"0F",X"0F",X"0F",X"06",
		X"00",X"00",X"00",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"08",X"08",X"0F",X"0F",X"0F",X"08",X"08",
		X"00",X"0E",X"01",X"01",X"01",X"0F",X"0F",X"0E",X"00",X"0F",X"00",X"00",X"00",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"0C",X"0F",X"0E",X"08",X"00",X"00",X"0C",X"03",X"00",X"00",X"03",X"0F",X"0E",
		X"00",X"0F",X"0E",X"0C",X"08",X"0C",X"0E",X"0F",X"00",X"0F",X"01",X"03",X"07",X"03",X"01",X"0F",
		X"00",X"07",X"0E",X"0C",X"08",X"04",X"02",X"01",X"00",X"08",X"04",X"03",X"03",X"07",X"0E",X"0C",
		X"00",X"00",X"00",X"00",X"08",X"0C",X"02",X"01",X"00",X"0C",X"02",X"01",X"03",X"07",X"0F",X"0E",
		X"00",X"01",X"01",X"09",X"0F",X"0F",X"0F",X"03",X"00",X"08",X"0E",X"0F",X"0F",X"0B",X"08",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"03",X"03",X"00",
		X"0C",X"06",X"02",X"02",X"02",X"02",X"06",X"0C",X"07",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"07",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"01",X"07",X"03",X"03",X"03",X"03",X"03",X"03",
		X"0C",X"0E",X"0E",X"0E",X"0C",X"08",X"00",X"0E",X"07",X"08",X"08",X"00",X"01",X"03",X"07",X"0F",
		X"0C",X"0E",X"0E",X"0C",X"0E",X"0E",X"0E",X"0C",X"07",X"08",X"00",X"01",X"00",X"08",X"08",X"07",
		X"0C",X"0C",X"0C",X"0C",X"0C",X"0E",X"0C",X"0C",X"00",X"01",X"03",X"05",X"09",X"0F",X"01",X"01",
		X"0C",X"00",X"00",X"0C",X"0E",X"0E",X"0E",X"0C",X"0F",X"08",X"08",X"0F",X"00",X"00",X"0C",X"03",
		X"0C",X"02",X"00",X"0C",X"02",X"02",X"02",X"0C",X"07",X"0E",X"0E",X"0F",X"0E",X"0E",X"0E",X"07",
		X"0E",X"0E",X"0C",X"08",X"08",X"00",X"00",X"00",X"0F",X"00",X"01",X"01",X"03",X"03",X"07",X"0F",
		X"08",X"04",X"04",X"08",X"0E",X"0E",X"06",X"0C",X"03",X"06",X"07",X"07",X"09",X"08",X"08",X"07",
		X"0C",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0C",X"07",X"08",X"08",X"08",X"07",X"00",X"08",X"07",
		X"08",X"0E",X"00",X"02",X"0A",X"0A",X"0E",X"00",X"00",X"01",X"00",X"02",X"02",X"02",X"03",X"00",
		X"00",X"0C",X"02",X"02",X"0E",X"00",X"0E",X"04",X"00",X"00",X"01",X"01",X"01",X"00",X"01",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"74",X"BA",X"DD",X"EE",X"FF",X"33",X"CC",X"F3",X"BB",X"BB",X"D5",X"D5",X"E2",X"F1",X"F0",X"F0",
		X"F0",X"F0",X"F8",X"74",X"BA",X"BA",X"DD",X"DD",X"FC",X"33",X"CC",X"FF",X"77",X"BB",X"D5",X"E2",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"34",X"1A",X"0D",X"0E",X"0F",X"03",X"0C",X"C3",X"0B",X"0B",X"85",X"85",X"C2",X"E1",X"F0",X"F0",
		X"F0",X"F0",X"78",X"34",X"1A",X"1A",X"0D",X"0D",X"3C",X"03",X"0C",X"0F",X"07",X"0B",X"85",X"C2",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"D5",X"D5",X"D5",X"E2",X"E2",X"E2",X"F1",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"00",X"BA",X"BA",X"BA",X"DD",X"DD",X"EE",X"66",
		X"66",X"77",X"BB",X"BB",X"D5",X"D5",X"D5",X"D5",X"F1",X"F1",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"74",X"74",X"74",X"BA",X"BA",X"BA",X"BA",
		X"00",X"85",X"85",X"85",X"C2",X"C2",X"C2",X"E1",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"78",X"78",X"00",X"1A",X"1A",X"1A",X"0D",X"0D",X"0E",X"06",
		X"06",X"07",X"0B",X"0B",X"85",X"85",X"85",X"85",X"E1",X"E1",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"78",X"34",X"34",X"34",X"1A",X"1A",X"1A",X"1A",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FE",X"11",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"00",X"FF",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"EE",X"00",X"EE",X"F0",X"F0",X"F0",X"FC",X"33",X"CC",X"FF",X"77",
		X"EE",X"FF",X"33",X"CC",X"F3",X"F0",X"F0",X"F0",X"FF",X"00",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"EE",X"00",X"EE",X"E0",X"E0",X"E0",X"E0",X"E0",X"88",X"F7",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"1E",X"01",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"00",X"0F",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"0E",X"00",X"0E",X"F0",X"F0",X"F0",X"3C",X"03",X"0C",X"0F",X"07",
		X"0E",X"0F",X"03",X"0C",X"C3",X"F0",X"F0",X"F0",X"0F",X"00",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"0E",X"00",X"0E",X"E0",X"E0",X"E0",X"E0",X"E0",X"08",X"87",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"DD",X"DD",X"BA",X"BA",X"74",X"F8",X"F0",X"F0",X"E2",X"D5",X"BB",X"77",X"FF",X"CC",X"33",X"FC",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F3",X"CC",X"33",X"FF",X"EE",X"DD",X"BA",X"74",X"F0",X"F0",X"F1",X"E2",X"D5",X"D5",X"BB",X"BB",
		X"0D",X"0D",X"1A",X"1A",X"34",X"78",X"F0",X"F0",X"C2",X"85",X"0B",X"07",X"0F",X"0C",X"03",X"3C",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"C3",X"0C",X"03",X"0F",X"0E",X"0D",X"1A",X"34",X"F0",X"F0",X"E1",X"C2",X"85",X"85",X"0B",X"0B",
		X"00",X"D5",X"D5",X"D5",X"BB",X"BB",X"77",X"66",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F1",X"F1",
		X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"BA",X"BA",X"BA",X"74",X"74",X"74",X"F8",
		X"F1",X"E2",X"E2",X"E2",X"D5",X"D5",X"D5",X"D5",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"66",X"EE",X"DD",X"DD",X"BA",X"BA",X"BA",X"BA",
		X"00",X"85",X"85",X"85",X"0B",X"0B",X"07",X"06",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"E1",X"E1",
		X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"1A",X"1A",X"1A",X"34",X"34",X"34",X"78",
		X"E1",X"C2",X"C2",X"C2",X"85",X"85",X"85",X"85",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"78",X"78",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"06",X"0E",X"0D",X"0D",X"1A",X"1A",X"1A",X"1A",
		X"F0",X"F0",X"F0",X"F3",X"CC",X"33",X"FF",X"EE",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"00",X"FF",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"EE",X"00",X"EE",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F7",X"88",
		X"11",X"FE",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"00",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"EE",X"00",X"EE",X"E0",X"E0",X"E0",X"E0",X"E0",X"77",X"FF",X"CC",X"33",X"FC",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"C3",X"0C",X"03",X"0F",X"0E",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"00",X"0F",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"0E",X"00",X"0E",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"87",X"08",
		X"01",X"1E",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"00",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"0E",X"00",X"0E",X"E0",X"E0",X"E0",X"E0",X"E0",X"07",X"0F",X"0C",X"03",X"3C",X"F0",X"F0",X"F0",
		X"D5",X"D5",X"D5",X"D5",X"D5",X"DD",X"00",X"DD",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"00",X"FF",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"00",X"FF",X"BA",X"BA",X"BA",X"BA",X"BA",X"BB",X"00",X"BB",
		X"DD",X"00",X"DD",X"D5",X"D5",X"D5",X"D5",X"D5",X"FF",X"00",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"FF",X"00",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"BB",X"00",X"BB",X"BA",X"BA",X"BA",X"BA",X"BA",
		X"85",X"85",X"85",X"85",X"85",X"8D",X"00",X"8D",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"00",X"FF",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"00",X"FF",X"1A",X"1A",X"1A",X"1A",X"1A",X"1B",X"00",X"1B",
		X"8D",X"00",X"8D",X"85",X"85",X"85",X"85",X"85",X"FF",X"00",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"FF",X"00",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"1B",X"00",X"1B",X"1A",X"1A",X"1A",X"1A",X"1A",
		X"D5",X"D5",X"D5",X"D5",X"D5",X"0D",X"00",X"0D",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"00",X"0F",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"00",X"0F",X"BA",X"BA",X"BA",X"BA",X"BA",X"0B",X"00",X"0B",
		X"0D",X"00",X"0D",X"D5",X"D5",X"D5",X"D5",X"D5",X"0F",X"00",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"00",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"0B",X"00",X"0B",X"BA",X"BA",X"BA",X"BA",X"BA",
		X"85",X"85",X"85",X"85",X"85",X"0D",X"00",X"0D",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"00",X"0F",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"00",X"0F",X"1A",X"1A",X"1A",X"1A",X"1A",X"0B",X"00",X"0B",
		X"0D",X"00",X"0D",X"85",X"85",X"85",X"85",X"85",X"0F",X"00",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"00",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"0B",X"00",X"0B",X"1A",X"1A",X"1A",X"1A",X"1A",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"00",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"00",X"FF",
		X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"BA",X"BA",X"BA",X"BA",X"BA",X"BA",X"BA",
		X"FF",X"00",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"00",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"00",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"00",X"0F",
		X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",
		X"0F",X"00",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"00",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"85",X"85",X"85",X"85",X"85",X"85",X"85",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"95",X"4A",X"2D",X"1E",X"0F",X"C3",X"3C",X"8B",X"4B",X"4B",X"A5",X"A5",X"D6",X"A3",X"D5",X"A2",
		X"10",X"BA",X"54",X"BA",X"54",X"1E",X"F0",X"1E",X"00",X"AA",X"55",X"2E",X"C3",X"3C",X"0F",X"87",
		X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"D5",X"A2",X"D5",X"A2",X"D5",X"A2",X"D5",X"A2",
		X"1E",X"F0",X"1E",X"BA",X"54",X"BA",X"54",X"BA",X"78",X"8F",X"55",X"AA",X"55",X"AA",X"55",X"AA",
		X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"D5",X"A2",X"D5",X"A2",X"D5",X"A2",X"D5",X"A2",
		X"54",X"BA",X"54",X"BA",X"54",X"1E",X"F0",X"1E",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"07",X"78",
		X"47",X"3C",X"C3",X"0F",X"1E",X"2D",X"5B",X"A6",X"D5",X"A2",X"C5",X"92",X"A5",X"A5",X"4B",X"4B",
		X"1E",X"F0",X"1E",X"BA",X"54",X"BA",X"54",X"1C",X"87",X"0F",X"3C",X"C3",X"1D",X"AA",X"55",X"8B",
		X"11",X"AA",X"55",X"8B",X"3C",X"C3",X"0F",X"1E",X"80",X"A2",X"D5",X"A2",X"D5",X"0F",X"F0",X"0F",
		X"2D",X"2D",X"5A",X"5A",X"94",X"3A",X"54",X"BA",X"56",X"AD",X"4B",X"87",X"0F",X"3C",X"C3",X"2E",
		X"E1",X"0E",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"0F",X"F0",X"0F",X"A2",X"D5",X"A2",X"D5",X"A2",
		X"54",X"BA",X"54",X"BA",X"54",X"BA",X"54",X"BA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",
		X"55",X"AA",X"55",X"AA",X"55",X"AA",X"0F",X"E1",X"D5",X"A2",X"D5",X"A2",X"D5",X"0F",X"F0",X"0F",
		X"54",X"BA",X"54",X"BA",X"54",X"BA",X"54",X"BA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",
		X"1E",X"0F",X"C3",X"3C",X"47",X"AA",X"55",X"0C",X"0F",X"F0",X"0F",X"A2",X"D5",X"A2",X"D5",X"83",
		X"54",X"BA",X"5C",X"B6",X"5A",X"5A",X"2D",X"2D",X"1D",X"C3",X"3C",X"0F",X"87",X"4B",X"25",X"9A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"AA",X"45",X"AB",X"45",X"AB",X"4C",X"2A",X"5A",X"4A",X"5B",X"4A",X"2D",X"2D",X"1E",X"96",
		X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"F0",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"F0",
		X"95",X"4A",X"2D",X"1E",X"0F",X"C3",X"3C",X"C3",X"4B",X"4B",X"25",X"AD",X"56",X"AB",X"55",X"F0",
		X"F0",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"F0",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",
		X"C3",X"3C",X"C3",X"0F",X"1E",X"2D",X"5B",X"A6",X"F0",X"AA",X"45",X"9A",X"25",X"AD",X"4B",X"4B",
		X"45",X"9A",X"56",X"9A",X"25",X"AD",X"25",X"A5",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"F0",
		X"5D",X"2A",X"45",X"AB",X"45",X"AB",X"44",X"F0",X"96",X"1E",X"2D",X"2D",X"5B",X"4A",X"5B",X"5A",
		X"F0",X"AD",X"25",X"AD",X"4B",X"4B",X"87",X"96",X"F0",X"22",X"55",X"22",X"55",X"22",X"45",X"AB",
		X"F0",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"F0",X"4A",X"5B",X"4A",X"95",X"A6",X"95",X"2A",
		X"2D",X"2D",X"5B",X"4A",X"95",X"2A",X"55",X"F0",X"56",X"AD",X"4B",X"87",X"0F",X"3C",X"C3",X"3C",
		X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"F0",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"F0",
		X"F0",X"AA",X"5D",X"A6",X"5B",X"4A",X"2D",X"2D",X"3C",X"C3",X"3C",X"0F",X"87",X"4B",X"25",X"9A",
		X"F0",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"F0",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",
		X"96",X"87",X"4B",X"4B",X"25",X"AD",X"25",X"A5",X"45",X"23",X"55",X"22",X"55",X"22",X"55",X"F0",
		X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"F0",X"5D",X"A6",X"95",X"A6",X"5B",X"4A",X"5B",X"5A",
		X"C4",X"EA",X"FD",X"FE",X"FF",X"F3",X"FC",X"33",X"FB",X"FB",X"F5",X"F5",X"B2",X"91",X"80",X"80",
		X"10",X"10",X"10",X"10",X"10",X"FE",X"F0",X"FE",X"00",X"00",X"00",X"CC",X"F3",X"FC",X"FF",X"F7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"FE",X"F0",X"FE",X"10",X"10",X"10",X"10",X"10",X"F8",X"77",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"10",X"10",X"10",X"10",X"10",X"FE",X"F0",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"F8",
		X"33",X"FC",X"F3",X"FF",X"FE",X"FD",X"EA",X"C4",X"80",X"80",X"91",X"B2",X"F5",X"F5",X"FB",X"FB",
		X"FE",X"F0",X"FE",X"10",X"10",X"10",X"10",X"DC",X"F7",X"FF",X"FC",X"F3",X"CC",X"00",X"00",X"33",
		X"00",X"00",X"00",X"33",X"FC",X"F3",X"FF",X"FE",X"80",X"80",X"80",X"80",X"80",X"FF",X"F0",X"FF",
		X"FD",X"FD",X"FA",X"FA",X"D4",X"98",X"10",X"10",X"32",X"75",X"FB",X"F7",X"FF",X"FC",X"F3",X"CC",
		X"F1",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"F0",X"FF",X"80",X"80",X"80",X"80",X"80",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"F1",X"80",X"80",X"80",X"80",X"80",X"FF",X"F0",X"FF",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"FE",X"FF",X"F3",X"FC",X"33",X"00",X"00",X"CC",X"FF",X"F0",X"FF",X"80",X"80",X"80",X"80",X"B3",
		X"10",X"10",X"98",X"D4",X"FA",X"FA",X"FD",X"FD",X"CC",X"F3",X"FC",X"FF",X"F7",X"FB",X"75",X"32",
		X"F0",X"75",X"75",X"75",X"32",X"32",X"32",X"11",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"11",X"11",X"11",X"11",X"88",X"88",X"F0",X"EA",X"EA",X"EA",X"FD",X"FD",X"FE",X"F6",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",
		X"C4",X"EA",X"FD",X"FE",X"FF",X"F3",X"FC",X"F3",X"FB",X"FB",X"75",X"75",X"32",X"11",X"00",X"F0",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F3",X"FC",X"F3",X"FF",X"FE",X"FD",X"EA",X"C4",X"F0",X"00",X"11",X"32",X"75",X"75",X"FB",X"FB",
		X"11",X"32",X"32",X"32",X"75",X"75",X"75",X"F5",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",
		X"88",X"88",X"11",X"11",X"11",X"11",X"00",X"F0",X"F6",X"FE",X"FD",X"FD",X"EA",X"EA",X"EA",X"FA",
		X"F0",X"75",X"75",X"75",X"FB",X"FB",X"F7",X"F6",X"F0",X"00",X"00",X"00",X"00",X"00",X"11",X"11",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"EA",X"EA",X"EA",X"C4",X"C4",X"C4",X"88",
		X"FD",X"FD",X"EA",X"EA",X"C4",X"88",X"00",X"F0",X"32",X"75",X"FB",X"F7",X"FF",X"FC",X"F3",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",
		X"F0",X"00",X"88",X"C4",X"EA",X"EA",X"FD",X"FD",X"FC",X"F3",X"FC",X"FF",X"F7",X"FB",X"75",X"32",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F6",X"F7",X"FB",X"FB",X"75",X"75",X"75",X"F5",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"88",X"C4",X"C4",X"C4",X"EA",X"EA",X"EA",X"FA",
		X"81",X"40",X"20",X"10",X"00",X"C0",X"30",X"08",X"40",X"40",X"A0",X"A0",X"94",X"82",X"85",X"82",
		X"14",X"1A",X"14",X"1A",X"14",X"10",X"F0",X"10",X"05",X"0A",X"05",X"02",X"C0",X"30",X"00",X"80",
		X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"85",X"82",X"85",X"82",X"85",X"82",X"85",X"82",
		X"10",X"F0",X"10",X"1A",X"14",X"1A",X"14",X"1A",X"70",X"08",X"05",X"0A",X"05",X"0A",X"05",X"0A",
		X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"85",X"82",X"85",X"82",X"85",X"82",X"85",X"82",
		X"14",X"1A",X"14",X"1A",X"14",X"10",X"F0",X"10",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"00",X"70",
		X"04",X"30",X"C0",X"00",X"10",X"20",X"41",X"82",X"85",X"82",X"84",X"90",X"A0",X"A0",X"40",X"40",
		X"10",X"F0",X"10",X"1A",X"14",X"1A",X"14",X"1A",X"80",X"00",X"30",X"C0",X"01",X"0A",X"05",X"0A",
		X"05",X"0A",X"05",X"08",X"30",X"C0",X"00",X"10",X"85",X"82",X"85",X"82",X"85",X"00",X"F0",X"00",
		X"20",X"20",X"50",X"50",X"90",X"12",X"14",X"1A",X"20",X"40",X"80",X"00",X"00",X"30",X"C0",X"02",
		X"E0",X"00",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"00",X"F0",X"00",X"82",X"85",X"82",X"85",X"82",
		X"14",X"1A",X"14",X"1A",X"14",X"1A",X"14",X"1A",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"0A",
		X"05",X"0A",X"05",X"0A",X"05",X"0A",X"00",X"E0",X"85",X"82",X"85",X"82",X"85",X"00",X"F0",X"00",
		X"14",X"1A",X"14",X"1A",X"14",X"1A",X"14",X"1A",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"0A",
		X"10",X"00",X"C0",X"30",X"04",X"0A",X"05",X"0A",X"00",X"F0",X"00",X"82",X"85",X"82",X"85",X"82",
		X"14",X"1A",X"14",X"92",X"50",X"50",X"20",X"20",X"01",X"C0",X"30",X"00",X"80",X"40",X"20",X"18",
		X"F0",X"28",X"20",X"28",X"14",X"18",X"14",X"0A",X"F0",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"0A",
		X"F0",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"02",X"F0",X"40",X"41",X"40",X"20",X"20",X"10",X"90",
		X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"F0",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"F0",
		X"81",X"40",X"20",X"10",X"00",X"C0",X"30",X"C0",X"40",X"40",X"20",X"28",X"14",X"0A",X"05",X"F0",
		X"F0",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"F0",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"0A",
		X"C0",X"30",X"C0",X"00",X"10",X"20",X"41",X"82",X"F0",X"0A",X"04",X"18",X"20",X"28",X"40",X"40",
		X"04",X"18",X"14",X"18",X"20",X"28",X"20",X"A0",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"F0",
		X"05",X"02",X"05",X"0A",X"05",X"0A",X"05",X"F0",X"90",X"10",X"20",X"20",X"41",X"40",X"41",X"50",
		X"F0",X"28",X"20",X"28",X"40",X"40",X"80",X"90",X"F0",X"0A",X"05",X"0A",X"05",X"0A",X"04",X"0A",
		X"F0",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"F0",X"40",X"41",X"40",X"81",X"82",X"81",X"02",
		X"20",X"20",X"41",X"40",X"81",X"02",X"05",X"F0",X"14",X"28",X"40",X"80",X"00",X"30",X"C0",X"30",
		X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"F0",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"F0",
		X"F0",X"0A",X"05",X"82",X"41",X"40",X"20",X"20",X"30",X"C0",X"30",X"00",X"80",X"40",X"20",X"18",
		X"F0",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"F0",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"0A",
		X"90",X"80",X"40",X"40",X"20",X"28",X"20",X"A0",X"04",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"F0",
		X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"F0",X"05",X"82",X"81",X"82",X"41",X"40",X"41",X"50",
		X"84",X"A6",X"84",X"A6",X"84",X"A6",X"84",X"A6",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",
		X"00",X"AA",X"0F",X"F0",X"0F",X"0F",X"F0",X"0F",X"00",X"AA",X"0F",X"F0",X"0F",X"0F",X"F0",X"0F",
		X"81",X"82",X"81",X"82",X"81",X"82",X"81",X"82",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"05",X"0A",X"00",X"F0",X"00",X"00",X"F0",X"00",X"05",X"0A",X"00",X"F0",X"00",X"00",X"F0",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"0A",
		X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",
		X"00",X"00",X"FF",X"F0",X"FF",X"FF",X"F0",X"FF",X"00",X"00",X"FF",X"F0",X"FF",X"FF",X"F0",X"FF",
		X"08",X"0C",X"86",X"C2",X"C2",X"86",X"0C",X"08",X"07",X"1E",X"4B",X"0F",X"0F",X"4B",X"1E",X"07",
		X"0C",X"86",X"4B",X"69",X"69",X"4B",X"86",X"0C",X"03",X"07",X"2D",X"0F",X"0F",X"2D",X"07",X"03",
		X"88",X"CC",X"AE",X"2E",X"2E",X"AE",X"CC",X"88",X"77",X"FF",X"9F",X"FF",X"FF",X"9F",X"FF",X"77",
		X"CC",X"EE",X"DF",X"9F",X"9F",X"DF",X"EE",X"CC",X"33",X"77",X"CF",X"FF",X"FF",X"CF",X"77",X"33",
		X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"56",X"12",X"56",X"12",X"56",X"12",X"56",X"12",
		X"0F",X"F0",X"0F",X"0F",X"F0",X"0F",X"55",X"00",X"0F",X"F0",X"0F",X"0F",X"F0",X"0F",X"55",X"00",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"14",X"18",X"14",X"18",X"14",X"18",X"14",X"18",
		X"00",X"F0",X"00",X"00",X"F0",X"00",X"05",X"0A",X"00",X"F0",X"00",X"00",X"F0",X"00",X"05",X"0A",
		X"F0",X"AD",X"25",X"AD",X"16",X"9A",X"56",X"AB",X"F0",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",
		X"FF",X"F0",X"FF",X"FF",X"F0",X"FF",X"00",X"00",X"FF",X"F0",X"FF",X"FF",X"F0",X"FF",X"00",X"00",
		X"EE",X"DF",X"9F",X"9F",X"DF",X"EE",X"CC",X"00",X"77",X"CF",X"FF",X"FF",X"CF",X"77",X"33",X"00",
		X"86",X"4B",X"69",X"69",X"4B",X"86",X"0C",X"00",X"07",X"2D",X"0F",X"0F",X"2D",X"07",X"03",X"00",
		X"CC",X"EE",X"DF",X"9F",X"9F",X"DF",X"EE",X"CC",X"33",X"77",X"CF",X"FF",X"FF",X"CF",X"77",X"33",
		X"0C",X"86",X"4B",X"69",X"69",X"4B",X"86",X"0C",X"03",X"07",X"2D",X"0F",X"0F",X"2D",X"07",X"03",
		X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",
		X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"F0",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"F0",
		X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"0E",X"0F",X"0C",X"0C",X"0C",X"0C",
		X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"07",X"03",X"01",X"00",X"00",X"00",X"00",
		X"01",X"03",X"07",X"0F",X"03",X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DD",X"DD",X"99",X"99",X"55",X"DD",X"00",X"DD",X"E2",X"D5",X"BB",X"77",X"FF",X"CC",X"00",X"FF",
		X"74",X"BA",X"DD",X"EE",X"FF",X"33",X"00",X"FF",X"BB",X"BB",X"99",X"99",X"AA",X"BB",X"00",X"BB",
		X"DD",X"00",X"DD",X"55",X"99",X"99",X"DD",X"DD",X"FF",X"00",X"CC",X"FF",X"77",X"BB",X"D5",X"E2",
		X"FF",X"00",X"33",X"FF",X"EE",X"DD",X"BA",X"74",X"BB",X"00",X"BB",X"AA",X"99",X"99",X"BB",X"BB",
		X"F0",X"F1",X"F1",X"F3",X"F3",X"F3",X"F7",X"F7",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F1",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"F0",X"F0",X"F1",X"F1",X"F3",X"F7",X"FF",
		X"F7",X"F7",X"F3",X"F3",X"F3",X"F1",X"F1",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"F1",X"FF",X"F7",X"F3",X"F1",X"F1",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F7",X"FF",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F3",X"F7",
		X"F0",X"F0",X"F0",X"F7",X"FF",X"FF",X"FF",X"FF",X"F0",X"F0",X"F0",X"F0",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"F7",X"F0",X"F0",X"F0",X"F0",X"F0",X"F7",X"F3",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"F7",X"F0",X"F0",X"F0",X"FF",X"FF",X"FF",X"FF",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"0F",X"0D",X"0B",X"07",X"F0",X"F0",X"F0",X"F0",X"0F",X"0B",X"0D",X"0E",
		X"E0",X"E0",X"E0",X"E0",X"0E",X"0C",X"0A",X"06",X"F0",X"F0",X"F0",X"F0",X"0F",X"0B",X"0D",X"0E",
		X"07",X"0B",X"0D",X"0F",X"F0",X"F0",X"F0",X"F0",X"0E",X"0D",X"0B",X"0F",X"F0",X"F0",X"F0",X"F0",
		X"06",X"0A",X"0C",X"0E",X"E0",X"E0",X"E0",X"E0",X"0E",X"0D",X"0B",X"0F",X"F0",X"F0",X"F0",X"F0",
		X"00",X"0B",X"0D",X"0E",X"0E",X"0D",X"0B",X"0F",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"0D",X"0B",X"07",X"07",X"0B",X"0D",X"0F",
		X"0F",X"0B",X"0D",X"0E",X"0E",X"0D",X"0B",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"0D",X"0B",X"07",X"07",X"0B",X"0D",X"0F",
		X"00",X"01",X"03",X"0E",X"0C",X"00",X"00",X"00",X"00",X"08",X"0C",X"07",X"03",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"0E",X"03",X"01",X"00",X"00",X"00",X"00",X"03",X"07",X"0C",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"0F",X"0F",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0F",
		X"00",X"00",X"07",X"0F",X"0F",X"0F",X"0F",X"F0",X"00",X"00",X"00",X"03",X"0F",X"0F",X"0F",X"F0",
		X"0F",X"0F",X"01",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"07",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"03",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"01",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"03",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"01",X"00",
		X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"EE",X"00",X"EE",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"00",X"FF",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"BA",X"BA",X"BA",X"BA",X"BA",X"BA",X"BA",X"BA",
		X"EE",X"00",X"EE",X"E0",X"E0",X"E0",X"E0",X"E0",X"FF",X"00",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"0E",X"00",X"0E",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"00",X"0F",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",
		X"0E",X"00",X"0E",X"E0",X"E0",X"E0",X"E0",X"E0",X"0F",X"00",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"85",X"85",X"85",X"85",X"85",X"85",X"85",X"85",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F3",X"CC",X"33",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"00",X"FF",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"EE",X"00",X"EE",X"F0",X"F0",X"F0",X"FC",X"33",X"CC",X"00",X"00",
		X"00",X"00",X"33",X"CC",X"F3",X"F0",X"F0",X"F0",X"FF",X"00",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"EE",X"00",X"EE",X"E0",X"E0",X"E0",X"E0",X"E0",X"00",X"00",X"CC",X"33",X"FC",X"F0",X"F0",X"F0",
		X"00",X"D5",X"D5",X"D5",X"88",X"88",X"44",X"44",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F1",X"F1",
		X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"00",X"BA",X"BA",X"BA",X"11",X"11",X"22",X"22",
		X"44",X"44",X"88",X"88",X"D5",X"D5",X"D5",X"D5",X"F1",X"F1",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"22",X"22",X"11",X"11",X"BA",X"BA",X"BA",X"BA",
		X"00",X"04",X"E2",X"F3",X"FF",X"BB",X"EE",X"00",X"00",X"02",X"70",X"78",X"78",X"70",X"04",X"04",
		X"88",X"89",X"C1",X"E1",X"E1",X"E1",X"E1",X"C1",X"33",X"22",X"70",X"70",X"70",X"70",X"70",X"70",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"F0",
		X"0F",X"0F",X"0F",X"0F",X"78",X"F0",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"F0",
		X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"78",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"F0",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"11",X"11",X"30",X"70",X"F0",X"E1",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"CC",X"88",X"88",X"C0",X"E0",X"F0",X"78",
		X"E1",X"F0",X"70",X"30",X"11",X"11",X"33",X"33",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"78",X"F0",X"E0",X"C0",X"88",X"88",X"00",X"00",
		X"22",X"66",X"66",X"66",X"74",X"70",X"F0",X"E1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"EE",X"FF",X"00",X"00",X"00",X"00",X"00",X"C0",X"F1",X"F0",X"78",
		X"E1",X"F0",X"F8",X"30",X"00",X"00",X"00",X"00",X"00",X"FF",X"77",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"78",X"F0",X"E0",X"E2",X"66",X"66",X"66",X"44",
		X"00",X"00",X"00",X"00",X"30",X"70",X"F0",X"E1",X"00",X"00",X"00",X"66",X"66",X"33",X"33",X"00",
		X"00",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"77",X"66",X"C0",X"E0",X"F0",X"78",
		X"E1",X"F0",X"70",X"30",X"66",X"EE",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",
		X"00",X"CC",X"CC",X"66",X"66",X"00",X"00",X"00",X"78",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"C3",X"0C",X"03",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"00",X"0F",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"0E",X"00",X"0E",X"F0",X"F0",X"F0",X"3C",X"03",X"0C",X"00",X"00",
		X"00",X"00",X"03",X"0C",X"C3",X"F0",X"F0",X"F0",X"0F",X"00",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"0E",X"00",X"0E",X"E0",X"E0",X"E0",X"E0",X"E0",X"00",X"00",X"0C",X"03",X"3C",X"F0",X"F0",X"F0",
		X"00",X"85",X"85",X"85",X"08",X"08",X"04",X"04",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"E1",X"E1",
		X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"78",X"78",X"00",X"1A",X"1A",X"1A",X"01",X"01",X"02",X"02",
		X"04",X"04",X"08",X"08",X"85",X"85",X"85",X"85",X"E1",X"E1",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"78",X"78",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"02",X"02",X"01",X"01",X"1A",X"1A",X"1A",X"1A",
		X"00",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"00",X"11",X"33",X"77",X"77",X"77",X"77",X"77",
		X"00",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"33",
		X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"77",X"77",X"77",X"77",X"77",X"33",X"11",X"00",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"CC",X"88",X"00",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"EE",X"00",X"00",X"00",X"00",X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",
		X"33",X"33",X"00",X"33",X"33",X"33",X"33",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"33",X"11",X"00",X"33",X"33",X"33",X"33",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"00",X"00",X"00",X"EE",X"EE",X"EE",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"33",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",
		X"33",X"33",X"00",X"11",X"33",X"33",X"33",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"EE",X"CC",X"88",X"EE",X"EE",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"11",X"33",X"33",X"33",X"33",X"33",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"EE",X"EE",X"EE",X"EE",X"CC",X"EE",X"EE",X"00",X"FF",X"FF",X"FF",X"FF",X"99",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"BB",X"BB",X"BB",
		X"33",X"33",X"33",X"33",X"33",X"11",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"CC",X"00",X"EE",X"BB",X"88",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",
		X"33",X"33",X"33",X"33",X"33",X"33",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"EE",X"00",X"00",X"00",X"00",X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"CC",X"FF",X"FF",X"99",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"11",X"33",X"33",X"33",X"33",X"33",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"CC",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"00",X"FF",X"FF",X"FF",X"99",X"FF",X"FF",X"FF",
		X"33",X"11",X"00",X"33",X"33",X"33",X"33",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"CC",X"00",X"00",X"00",X"00",X"EE",X"EE",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"CF",X"C4",X"C6",X"CC",X"DD",X"FF",X"00",X"00",X"11",X"32",X"76",X"76",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",X"06",X"22",X"6E",X"66",X"EE",X"EE",
		X"FF",X"FF",X"DD",X"CC",X"C6",X"C4",X"CF",X"44",X"FF",X"FF",X"FF",X"76",X"76",X"32",X"11",X"00",
		X"00",X"00",X"00",X"C0",X"C0",X"00",X"00",X"00",X"EE",X"EE",X"EE",X"66",X"6E",X"22",X"06",X"00",
		X"00",X"01",X"02",X"19",X"13",X"19",X"BB",X"BB",X"00",X"00",X"00",X"23",X"77",X"75",X"FD",X"FD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"B8",X"88",X"CC",X"CC",X"EE",
		X"FF",X"FF",X"EE",X"EE",X"FF",X"F9",X"F8",X"77",X"FF",X"FF",X"FF",X"77",X"77",X"33",X"11",X"00",
		X"60",X"60",X"00",X"88",X"0C",X"00",X"00",X"00",X"EE",X"FF",X"FF",X"02",X"08",X"02",X"8C",X"88",
		X"00",X"00",X"0C",X"22",X"33",X"15",X"19",X"33",X"00",X"00",X"00",X"00",X"01",X"46",X"EE",X"F9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"00",X"00",X"C0",X"C0",X"00",X"88",X"CC",X"EE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FE",X"77",X"F9",X"FD",X"FF",X"77",X"77",X"33",X"11",X"00",
		X"00",X"88",X"04",X"04",X"00",X"00",X"00",X"00",X"FF",X"FF",X"89",X"00",X"8C",X"C5",X"E6",X"CC",
		X"00",X"30",X"30",X"CC",X"77",X"7F",X"33",X"33",X"00",X"00",X"00",X"01",X"00",X"02",X"04",X"CD",
		X"00",X"00",X"00",X"00",X"C0",X"C0",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"CC",X"FF",X"FF",
		X"33",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"FF",X"F9",X"F8",X"77",X"77",X"33",X"11",X"00",
		X"02",X"04",X"00",X"08",X"88",X"88",X"00",X"00",X"FF",X"CD",X"00",X"CE",X"FF",X"F1",X"FF",X"CC",
		X"00",X"00",X"80",X"80",X"00",X"FF",X"FF",X"77",X"00",X"00",X"10",X"10",X"00",X"37",X"15",X"01",
		X"00",X"00",X"00",X"00",X"00",X"8C",X"04",X"00",X"00",X"00",X"30",X"30",X"00",X"FF",X"FF",X"CD",
		X"77",X"33",X"FF",X"FF",X"F7",X"FF",X"FF",X"77",X"04",X"05",X"FF",X"74",X"74",X"33",X"11",X"00",
		X"04",X"04",X"EE",X"C4",X"C4",X"88",X"00",X"00",X"CC",X"89",X"FF",X"FE",X"FC",X"FF",X"FF",X"CC",
		X"00",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"11",X"33",X"77",X"77",X"F9",X"F9",
		X"00",X"00",X"00",X"88",X"08",X"08",X"00",X"04",X"00",X"CC",X"FF",X"F1",X"FF",X"CE",X"00",X"CD",
		X"33",X"77",X"77",X"7F",X"66",X"88",X"30",X"30",X"FB",X"CD",X"04",X"02",X"00",X"01",X"01",X"00",
		X"8A",X"88",X"00",X"C0",X"C0",X"00",X"00",X"00",X"FF",X"FF",X"EE",X"88",X"00",X"00",X"00",X"00",
		X"00",X"77",X"FE",X"FC",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"11",X"33",X"77",X"77",X"FF",X"FD",
		X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"88",X"00",X"CC",X"E6",X"C6",X"89",X"04",X"02",X"99",
		X"FF",X"77",X"33",X"33",X"37",X"22",X"0C",X"00",X"F9",X"F9",X"EF",X"44",X"02",X"00",X"00",X"00",
		X"00",X"60",X"60",X"00",X"00",X"00",X"00",X"00",X"FF",X"EE",X"CC",X"88",X"00",X"00",X"C0",X"C0",
		X"00",X"77",X"F9",X"F9",X"FB",X"EE",X"EE",X"FF",X"00",X"00",X"11",X"33",X"77",X"77",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"08",X"88",X"88",X"60",X"00",X"88",X"8C",X"02",X"08",X"02",X"33",X"FF",
		X"FF",X"BB",X"BB",X"19",X"13",X"08",X"02",X"01",X"FF",X"FD",X"FD",X"75",X"77",X"33",X"00",X"00",
		X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"EE",X"EE",X"CC",X"CC",X"B8",X"B8",X"00",
		X"00",X"00",X"00",X"00",X"01",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"0F",
		X"00",X"00",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"03",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"01",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"07",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"03",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"01",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"01",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"FF",X"FF",X"CC",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"EE",X"CC",X"CC",X"CC",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"CC",X"FF",X"FF",X"FF",X"CC",X"CC",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",
		X"EE",X"CC",X"88",X"88",X"88",X"88",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"EE",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"EE",X"88",X"00",X"00",
		X"00",X"88",X"88",X"88",X"88",X"CC",X"EE",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"EE",X"FF",X"FF",X"FF",X"00",X"88",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"88",X"88",X"88",X"88",X"00",X"00",X"00",
		X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"EE",X"EE",X"CC",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"88",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"CC",X"CC",X"EE",X"EE",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"EE",X"88",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"EE",X"CC",X"00",X"00",X"00",
		X"CC",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"88",X"EE",X"FF",X"00",X"00",X"00",X"CC",X"EE",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"FF",X"FF",
		X"EE",X"CC",X"CC",X"88",X"88",X"88",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"EE",X"CC",X"88",X"88",X"00",X"00",
		X"00",X"00",X"88",X"88",X"88",X"CC",X"CC",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"88",X"88",X"CC",X"EE",X"FF",X"FF",
		X"00",X"03",X"78",X"78",X"70",X"70",X"70",X"FF",X"00",X"00",X"03",X"03",X"00",X"00",X"00",X"33",
		X"00",X"00",X"00",X"00",X"0C",X"0C",X"00",X"00",X"00",X"0E",X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",
		X"11",X"11",X"11",X"11",X"FF",X"FF",X"FF",X"00",X"33",X"33",X"33",X"33",X"33",X"11",X"00",X"00",
		X"0C",X"0C",X"00",X"00",X"04",X"00",X"00",X"00",X"F8",X"F8",X"F8",X"FF",X"FF",X"EE",X"CC",X"00",
		X"00",X"34",X"78",X"F0",X"F0",X"F0",X"F0",X"F1",X"00",X"00",X"00",X"01",X"12",X"1E",X"0C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0C",X"00",X"80",X"C3",X"C3",X"E0",X"E0",X"F0",X"F8",
		X"77",X"88",X"88",X"88",X"CC",X"FF",X"FF",X"33",X"00",X"11",X"11",X"11",X"11",X"00",X"00",X"00",
		X"80",X"8A",X"CC",X"88",X"88",X"88",X"00",X"00",X"F8",X"FC",X"FF",X"77",X"FF",X"FF",X"EE",X"CC",
		X"00",X"24",X"78",X"F0",X"F0",X"F0",X"F0",X"F1",X"00",X"00",X"00",X"01",X"12",X"30",X"34",X"1E",
		X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"82",X"00",X"04",X"0C",X"84",X"C0",X"E1",X"F0",X"F8",
		X"F3",X"E6",X"CC",X"CC",X"EE",X"77",X"33",X"11",X"1C",X"00",X"00",X"11",X"00",X"00",X"00",X"00",
		X"CC",X"CC",X"CC",X"CC",X"88",X"00",X"00",X"00",X"FC",X"FF",X"77",X"33",X"77",X"FF",X"EE",X"CC",
		X"00",X"03",X"C3",X"F0",X"F0",X"F0",X"F0",X"F1",X"00",X"00",X"01",X"12",X"12",X"34",X"70",X"70",
		X"00",X"00",X"00",X"00",X"02",X"00",X"CC",X"CC",X"00",X"00",X"00",X"03",X"C3",X"F0",X"F0",X"F9",
		X"F3",X"E2",X"44",X"44",X"FF",X"77",X"11",X"00",X"34",X"0E",X"0C",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"EE",X"CC",X"CC",X"88",X"88",X"00",X"00",X"FF",X"FF",X"33",X"33",X"33",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"33",X"33",X"22",X"E2",X"E2",X"00",X"00",X"00",X"06",X"06",X"06",X"70",X"78",
		X"00",X"00",X"00",X"00",X"88",X"CC",X"CC",X"CC",X"00",X"00",X"00",X"FF",X"FF",X"11",X"11",X"11",
		X"F3",X"F3",X"F0",X"F0",X"F0",X"09",X"09",X"00",X"78",X"78",X"78",X"78",X"70",X"01",X"01",X"00",
		X"CC",X"CC",X"CC",X"88",X"00",X"00",X"00",X"00",X"FF",X"FF",X"F3",X"F3",X"F3",X"08",X"09",X"00",
		X"00",X"00",X"11",X"77",X"FF",X"44",X"44",X"E2",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0E",
		X"00",X"00",X"00",X"88",X"88",X"CC",X"CC",X"EE",X"00",X"00",X"FF",X"FF",X"33",X"33",X"33",X"FF",
		X"F3",X"F1",X"F0",X"F0",X"F0",X"F0",X"4B",X"03",X"34",X"70",X"70",X"70",X"12",X"03",X"01",X"00",
		X"CC",X"CC",X"CC",X"00",X"02",X"00",X"00",X"00",X"FF",X"F9",X"F0",X"F0",X"C3",X"03",X"00",X"00",
		X"00",X"11",X"33",X"77",X"EE",X"CC",X"CC",X"66",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"88",X"CC",X"CC",X"CC",X"00",X"CC",X"EE",X"FF",X"77",X"33",X"77",X"FF",
		X"F3",X"F1",X"F0",X"F0",X"F0",X"F0",X"78",X"24",X"0C",X"1E",X"34",X"30",X"12",X"01",X"00",X"00",
		X"CC",X"82",X"08",X"08",X"08",X"00",X"00",X"00",X"FC",X"F8",X"F0",X"E1",X"C0",X"84",X"0C",X"04",
		X"00",X"33",X"FF",X"FF",X"CC",X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"11",
		X"00",X"00",X"00",X"88",X"88",X"88",X"CC",X"8A",X"00",X"CC",X"EE",X"FF",X"FF",X"77",X"FF",X"FC",
		X"77",X"F1",X"F0",X"F0",X"F0",X"F0",X"78",X"07",X"00",X"00",X"0C",X"1E",X"12",X"10",X"00",X"00",
		X"80",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"F8",X"F8",X"F0",X"E0",X"E0",X"C3",X"C3",X"80",
		X"00",X"00",X"FF",X"FF",X"FF",X"11",X"11",X"11",X"00",X"00",X"00",X"11",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"0C",X"00",X"00",X"CC",X"EE",X"FF",X"FF",X"F8",X"F8",
		X"11",X"FF",X"70",X"70",X"70",X"78",X"78",X"03",X"33",X"33",X"00",X"00",X"00",X"03",X"03",X"00",
		X"0C",X"00",X"00",X"0C",X"0C",X"00",X"00",X"00",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"0E",
		X"00",X"22",X"FF",X"FF",X"FF",X"FF",X"33",X"33",X"00",X"00",X"00",X"33",X"77",X"77",X"66",X"66",
		X"00",X"00",X"00",X"00",X"08",X"08",X"00",X"00",X"00",X"01",X"CC",X"CC",X"E9",X"E1",X"F0",X"F8",
		X"11",X"33",X"FC",X"30",X"10",X"12",X"07",X"06",X"77",X"33",X"33",X"11",X"00",X"00",X"00",X"00",
		X"86",X"86",X"C0",X"C0",X"84",X"08",X"00",X"00",X"F8",X"F0",X"F0",X"F0",X"F0",X"E1",X"C2",X"00",
		X"00",X"00",X"FF",X"FF",X"FE",X"FE",X"77",X"33",X"00",X"00",X"00",X"11",X"33",X"77",X"FF",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"84",X"00",X"08",X"00",X"87",X"C2",X"E0",X"F0",X"F8",
		X"11",X"33",X"FE",X"DC",X"88",X"00",X"01",X"01",X"EE",X"77",X"33",X"11",X"00",X"00",X"00",X"00",
		X"C0",X"E0",X"C2",X"84",X"08",X"00",X"00",X"00",X"F8",X"F0",X"F0",X"F0",X"F0",X"69",X"0C",X"08",
		X"00",X"02",X"44",X"FE",X"FC",X"FC",X"FE",X"77",X"00",X"00",X"00",X"33",X"33",X"77",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"0C",X"0C",X"C0",X"C2",X"00",X"00",X"0C",X"0C",X"C0",X"F0",X"F0",X"F8",
		X"11",X"11",X"11",X"EE",X"EE",X"00",X"00",X"00",X"EE",X"EE",X"77",X"77",X"11",X"00",X"00",X"00",
		X"C2",X"C2",X"C2",X"84",X"80",X"00",X"00",X"00",X"F8",X"F0",X"F0",X"F0",X"34",X"07",X"0E",X"0C",
		X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"77",X"77",X"77",
		X"00",X"00",X"00",X"0C",X"0C",X"0C",X"C0",X"C2",X"00",X"00",X"00",X"88",X"88",X"88",X"F8",X"F8",
		X"FF",X"FF",X"F8",X"F8",X"F8",X"03",X"03",X"00",X"77",X"77",X"77",X"33",X"11",X"00",X"01",X"00",
		X"C2",X"C2",X"C2",X"C2",X"C0",X"00",X"00",X"00",X"F8",X"F8",X"F0",X"F0",X"F0",X"03",X"03",X"00",
		X"00",X"00",X"00",X"00",X"EE",X"EE",X"11",X"11",X"00",X"00",X"00",X"00",X"11",X"77",X"77",X"EE",
		X"00",X"00",X"00",X"00",X"08",X"84",X"C2",X"E0",X"00",X"06",X"06",X"03",X"30",X"F0",X"F0",X"F0",
		X"11",X"77",X"FE",X"FC",X"FC",X"FE",X"44",X"04",X"EE",X"FF",X"FF",X"77",X"33",X"33",X"00",X"00",
		X"E0",X"E0",X"C0",X"0C",X"0C",X"00",X"00",X"00",X"F8",X"F8",X"F0",X"F0",X"C0",X"0C",X"0C",X"00",
		X"00",X"01",X"01",X"00",X"88",X"DC",X"FE",X"33",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"77",
		X"00",X"00",X"00",X"00",X"08",X"84",X"C2",X"E0",X"00",X"08",X"0C",X"69",X"F0",X"F0",X"F0",X"F0",
		X"11",X"33",X"77",X"FE",X"FE",X"FF",X"FF",X"00",X"EE",X"EE",X"FF",X"77",X"33",X"11",X"00",X"00",
		X"C0",X"84",X"0E",X"00",X"00",X"00",X"00",X"00",X"F8",X"F8",X"F0",X"E0",X"C2",X"87",X"00",X"08",
		X"00",X"06",X"07",X"12",X"10",X"30",X"FC",X"33",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"33",
		X"00",X"00",X"00",X"08",X"84",X"C0",X"C0",X"86",X"00",X"00",X"C2",X"E1",X"F0",X"F0",X"F0",X"F0",
		X"11",X"33",X"33",X"FF",X"FF",X"FF",X"FF",X"22",X"77",X"66",X"66",X"77",X"77",X"33",X"00",X"00",
		X"86",X"00",X"00",X"08",X"08",X"00",X"00",X"00",X"F8",X"F8",X"F0",X"E1",X"E9",X"CC",X"CC",X"01");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
