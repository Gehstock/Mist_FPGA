library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity gfx1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of gfx1 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"11",X"11",X"1B",X"BA",X"BB",X"2B",X"FF",X"FF",X"44",X"44",X"44",X"44",X"FF",X"FF",X"33",X"33",
		X"12",X"22",X"22",X"22",X"FF",X"FF",X"F2",X"22",X"F2",X"B2",X"4F",X"FF",X"FF",X"FF",X"33",X"F2",
		X"33",X"33",X"FF",X"FF",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"33",X"FC",X"33",X"FC",X"33",X"CC",X"33",X"CF",X"33",X"C2",X"33",X"AC",X"33",X"BB",X"33",X"CC",
		X"33",X"DD",X"FF",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"77",X"88",X"77",X"18",X"FF",X"18",X"F2",X"1A",X"77",X"88",X"AA",X"77",X"7F",X"14",X"4F",
		X"DD",X"DF",X"11",X"1F",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"88",X"7F",X"87",X"4F",X"14",X"4F",X"17",X"4F",X"14",X"4F",X"11",X"4F",X"44",X"CF",X"14",X"CF",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FA",X"FF",X"12",X"11",X"11",X"12",X"A2",X"A2",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FA",X"AF",X"12",X"AF",X"11",X"AF",X"A2",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AF",X"AF",X"2F",X"2F",X"AF",X"2F",X"2A",X"2A",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AF",X"AA",X"2F",X"2F",X"2F",X"2F",X"2A",X"AA",X"AA",X"AA",
		X"22",X"11",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"22",X"11",X"22",X"22",
		X"22",X"12",X"22",X"12",X"22",X"12",X"22",X"12",X"22",X"12",X"22",X"12",X"22",X"12",X"22",X"22",
		X"22",X"11",X"21",X"21",X"22",X"21",X"22",X"11",X"21",X"22",X"21",X"22",X"21",X"11",X"22",X"22",
		X"22",X"11",X"21",X"21",X"22",X"21",X"22",X"11",X"22",X"21",X"21",X"21",X"22",X"11",X"22",X"22",
		X"22",X"11",X"22",X"11",X"22",X"11",X"21",X"11",X"21",X"11",X"21",X"11",X"22",X"11",X"22",X"22",
		X"21",X"11",X"21",X"22",X"21",X"11",X"22",X"21",X"22",X"21",X"21",X"21",X"22",X"11",X"22",X"22",
		X"22",X"11",X"21",X"21",X"21",X"22",X"21",X"11",X"21",X"21",X"21",X"21",X"22",X"11",X"22",X"22",
		X"21",X"11",X"22",X"21",X"22",X"11",X"22",X"12",X"22",X"12",X"22",X"12",X"22",X"12",X"22",X"22",
		X"22",X"11",X"21",X"21",X"21",X"21",X"22",X"11",X"21",X"21",X"21",X"21",X"22",X"11",X"22",X"22",
		X"22",X"11",X"21",X"21",X"21",X"21",X"22",X"11",X"22",X"21",X"21",X"21",X"22",X"11",X"22",X"22",
		X"33",X"33",X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00",
		X"33",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"00",X"1A",X"00",X"1A",X"00",X"AA",X"00",X"A0",X"01",X"00",X"01",X"00",X"00",X"00",
		X"2D",X"DD",X"21",X"11",X"21",X"11",X"21",X"11",X"21",X"11",X"21",X"11",X"21",X"11",X"21",X"11",
		X"DD",X"DD",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AF",X"AF",X"AF",X"AF",X"2F",X"2A",X"2A",X"2A",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"2A",X"AA",X"2A",X"FA",X"AA",X"22",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FF",X"FA",X"FF",X"F2",X"F2",X"F2",X"A2",X"A2",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FA",X"FA",X"22",X"22",X"2A",X"FA",X"2A",X"22",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FA",X"AA",X"F2",X"AA",X"22",X"AA",X"AA",X"AA",
		X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00",X"33",X"33",
		X"01",X"01",X"00",X"10",X"00",X"0A",X"00",X"10",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"33",
		X"FF",X"FF",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"FF",X"FF",X"AA",X"AA",X"AA",X"A2",X"AA",X"A2",
		X"FF",X"FF",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"FF",X"FF",X"22",X"AA",X"22",X"AA",X"22",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"A0",
		X"22",X"AA",X"22",X"2A",X"22",X"2A",X"22",X"22",X"22",X"22",X"FF",X"FF",X"EE",X"EE",X"EE",X"EE",
		X"01",X"11",X"11",X"33",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"01",X"11",X"00",X"33",
		X"01",X"10",X"00",X"13",X"00",X"13",X"00",X"13",X"00",X"13",X"00",X"13",X"00",X"13",X"00",X"33",
		X"01",X"11",X"10",X"11",X"03",X"11",X"01",X"11",X"11",X"33",X"11",X"00",X"11",X"11",X"03",X"33",
		X"01",X"11",X"10",X"11",X"03",X"11",X"00",X"11",X"00",X"11",X"10",X"11",X"01",X"11",X"00",X"33",
		X"00",X"11",X"00",X"11",X"01",X"11",X"10",X"11",X"13",X"11",X"11",X"11",X"03",X"11",X"00",X"33",
		X"11",X"11",X"11",X"33",X"11",X"11",X"11",X"11",X"03",X"11",X"10",X"11",X"01",X"11",X"00",X"33",
		X"01",X"11",X"11",X"33",X"11",X"00",X"11",X"11",X"11",X"33",X"11",X"00",X"01",X"11",X"00",X"33",
		X"11",X"11",X"03",X"11",X"00",X"11",X"00",X"11",X"00",X"13",X"00",X"13",X"00",X"13",X"00",X"33",
		X"01",X"11",X"11",X"33",X"11",X"00",X"01",X"11",X"11",X"33",X"11",X"00",X"01",X"11",X"00",X"33",
		X"01",X"11",X"10",X"11",X"13",X"11",X"01",X"11",X"00",X"11",X"10",X"11",X"01",X"11",X"00",X"33",
		X"AA",X"22",X"AA",X"22",X"AA",X"22",X"AA",X"22",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"22",X"AA",X"22",X"AA",X"22",X"2A",X"22",X"22",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"01",X"11",X"01",X"11",X"01",X"11",X"00",X"AA",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"11",X"00",X"AA",X"01",X"11",X"00",X"AA",X"00",X"00",X"00",X"00",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"01",X"11",X"11",X"11",X"0A",X"11",X"00",X"11",X"00",X"AA",X"00",X"A0",X"00",X"00",X"00",X"A0",
		X"AA",X"22",X"AA",X"22",X"AA",X"22",X"AA",X"22",X"A2",X"22",X"FF",X"FF",X"EE",X"EE",X"EE",X"EE",
		X"01",X"11",X"10",X"11",X"1A",X"11",X"1A",X"11",X"11",X"11",X"1A",X"11",X"1A",X"11",X"0A",X"0A",
		X"11",X"11",X"11",X"AA",X"11",X"00",X"11",X"11",X"11",X"AA",X"11",X"00",X"11",X"11",X"0A",X"AA",
		X"01",X"11",X"11",X"AA",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"01",X"11",X"00",X"AA",
		X"11",X"11",X"11",X"AA",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"11",X"0A",X"AA",
		X"11",X"11",X"11",X"AA",X"11",X"00",X"11",X"11",X"11",X"AA",X"11",X"00",X"11",X"11",X"0A",X"AA",
		X"11",X"11",X"11",X"AA",X"11",X"00",X"11",X"11",X"11",X"AA",X"11",X"00",X"11",X"00",X"0A",X"00",
		X"01",X"11",X"11",X"AA",X"11",X"00",X"11",X"11",X"11",X"0A",X"11",X"00",X"01",X"11",X"00",X"AA",
		X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"11",X"11",X"AA",X"11",X"00",X"11",X"00",X"0A",X"00",
		X"00",X"10",X"00",X"1A",X"00",X"1A",X"00",X"1A",X"00",X"1A",X"00",X"1A",X"00",X"1A",X"00",X"AA",
		X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"01",X"1A",X"00",X"AA",
		X"11",X"00",X"11",X"01",X"11",X"10",X"11",X"1A",X"11",X"11",X"11",X"01",X"11",X"01",X"0A",X"00",
		X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"11",X"0A",X"AA",
		X"11",X"01",X"11",X"11",X"11",X"11",X"11",X"1A",X"11",X"0A",X"11",X"00",X"11",X"00",X"0A",X"00",
		X"11",X"00",X"11",X"00",X"11",X"10",X"11",X"11",X"1A",X"11",X"1A",X"11",X"1A",X"11",X"0A",X"0A",
		X"01",X"11",X"11",X"AA",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"01",X"11",X"00",X"AA",
		X"11",X"11",X"11",X"AA",X"11",X"00",X"11",X"00",X"11",X"11",X"11",X"0A",X"11",X"00",X"0A",X"00",
		X"01",X"11",X"11",X"AA",X"11",X"00",X"11",X"00",X"11",X"10",X"11",X"1A",X"01",X"11",X"00",X"AA",
		X"11",X"11",X"11",X"AA",X"11",X"00",X"11",X"00",X"11",X"11",X"11",X"AA",X"11",X"00",X"0A",X"00",
		X"01",X"11",X"11",X"AA",X"11",X"00",X"01",X"11",X"00",X"11",X"10",X"11",X"01",X"11",X"00",X"AA",
		X"11",X"11",X"0A",X"1A",X"00",X"1A",X"00",X"1A",X"00",X"1A",X"00",X"1A",X"00",X"1A",X"00",X"AA",
		X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"01",X"11",X"00",X"AA",
		X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"01",X"01",X"00",X"10",X"00",X"AA",
		X"11",X"10",X"11",X"1A",X"11",X"1A",X"11",X"1A",X"11",X"1A",X"11",X"1A",X"01",X"01",X"00",X"A0",
		X"11",X"00",X"11",X"00",X"11",X"00",X"01",X"11",X"10",X"11",X"1A",X"11",X"1A",X"11",X"0A",X"0A",
		X"11",X"00",X"11",X"00",X"11",X"00",X"01",X"11",X"00",X"1A",X"00",X"1A",X"00",X"1A",X"00",X"AA",
		X"11",X"11",X"0A",X"11",X"00",X"11",X"00",X"1A",X"01",X"AA",X"11",X"A0",X"11",X"11",X"0A",X"AA",
		X"07",X"77",X"7F",X"77",X"79",X"77",X"77",X"77",X"07",X"77",X"00",X"70",X"00",X"00",X"00",X"00",
		X"00",X"33",X"08",X"22",X"8F",X"24",X"77",X"87",X"27",X"F7",X"02",X"77",X"00",X"77",X"00",X"22",
		X"00",X"00",X"00",X"03",X"0C",X"32",X"CF",X"20",X"CC",X"CC",X"2C",X"FC",X"02",X"CC",X"00",X"CB",
		X"00",X"00",X"00",X"C0",X"0C",X"CC",X"CF",X"CC",X"CC",X"CB",X"0B",X"BB",X"00",X"B0",X"00",X"00",
		X"00",X"04",X"08",X"47",X"8F",X"87",X"8F",X"87",X"88",X"77",X"07",X"77",X"00",X"70",X"00",X"00",
		X"22",X"22",X"2C",X"2C",X"2F",X"22",X"FF",X"FF",X"FF",X"EF",X"EE",X"21",X"FF",X"22",X"FF",X"F2",
		X"AA",X"BB",X"AA",X"BB",X"EA",X"AA",X"1E",X"BB",X"1E",X"B2",X"1A",X"2B",X"1A",X"BB",X"44",X"BB",
		X"FF",X"FF",X"CF",X"C4",X"CF",X"C4",X"CC",X"C4",X"CC",X"CC",X"FF",X"FC",X"FF",X"FC",X"F2",X"2C",
		X"44",X"4B",X"94",X"44",X"77",X"44",X"77",X"44",X"C4",X"44",X"CC",X"44",X"4C",X"44",X"44",X"11",
		X"BB",X"B1",X"BB",X"17",X"2F",X"17",X"F2",X"B7",X"FF",X"BB",X"FC",X"BB",X"CC",X"1B",X"FC",X"CC",
		X"77",X"7F",X"72",X"FF",X"27",X"22",X"77",X"22",X"77",X"18",X"77",X"89",X"C1",X"89",X"C1",X"99",
		X"CC",X"CC",X"CC",X"FC",X"CC",X"2C",X"AC",X"CC",X"AA",X"AC",X"1A",X"CC",X"AA",X"CC",X"2A",X"CC",
		X"C8",X"F9",X"C8",X"29",X"C8",X"29",X"B8",X"92",X"11",X"99",X"CC",X"99",X"B8",X"99",X"BB",X"88",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"2F",X"22",X"2F",X"22",X"F1",X"22",X"F1",
		X"F2",X"22",X"F2",X"22",X"1F",X"22",X"1F",X"22",X"11",X"22",X"11",X"22",X"11",X"22",X"11",X"22",
		X"22",X"11",X"22",X"11",X"22",X"11",X"22",X"11",X"2F",X"11",X"2F",X"11",X"F1",X"11",X"F1",X"11",
		X"11",X"F2",X"11",X"F2",X"11",X"1F",X"11",X"1F",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"22",X"22",X"22",X"22",X"22",X"2D",X"22",X"2E",X"22",X"DE",X"22",X"EE",X"22",X"EE",X"22",X"EE",
		X"ED",X"22",X"EE",X"22",X"EE",X"22",X"EE",X"22",X"EE",X"22",X"EE",X"22",X"EE",X"D2",X"EE",X"E2",
		X"22",X"EE",X"22",X"EE",X"2D",X"EE",X"2E",X"EE",X"2F",X"FF",X"2F",X"DD",X"2F",X"DD",X"2F",X"FF",
		X"EE",X"ED",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"FF",X"FF",X"DD",X"DD",X"DD",X"DD",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AF",X"AA",X"AF",X"AA",X"F1",X"AA",X"F1",
		X"FA",X"AA",X"FA",X"AA",X"1F",X"AA",X"1F",X"AA",X"11",X"AA",X"11",X"AA",X"11",X"AA",X"11",X"AA",
		X"AA",X"11",X"AA",X"11",X"AA",X"11",X"AA",X"11",X"AF",X"11",X"AF",X"11",X"F1",X"11",X"F1",X"11",
		X"11",X"FA",X"11",X"FA",X"11",X"1F",X"11",X"1F",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AD",X"AA",X"AE",X"AA",X"DE",X"AA",X"EE",
		X"DA",X"AA",X"EA",X"AA",X"ED",X"AA",X"EE",X"AA",X"EE",X"AA",X"EE",X"AA",X"EE",X"AA",X"EE",X"AA",
		X"AA",X"EE",X"AA",X"EE",X"AA",X"EE",X"AA",X"EE",X"AA",X"FF",X"AA",X"DD",X"AA",X"DD",X"AA",X"FF",
		X"EE",X"DA",X"EE",X"EA",X"EE",X"ED",X"EE",X"EE",X"FF",X"FF",X"DD",X"DF",X"DD",X"DF",X"FF",X"FF",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"FF",X"FF",X"EE",X"EE",X"EE",X"EE",
		X"FF",X"FF",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"FF",X"FF",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"D2",X"22",X"E2",X"22",
		X"01",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"01",X"11",X"01",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"01",X"11",X"01",X"11",
		X"11",X"01",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"01",X"11",X"00",X"00",
		X"11",X"01",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AF",
		X"AA",X"11",X"AF",X"11",X"EF",X"11",X"F1",X"11",X"E1",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"AA",X"EF",X"AA",X"F1",X"AA",X"E1",X"AA",X"11",X"AA",X"11",X"AF",X"11",X"EF",X"11",X"F1",X"11",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AF",X"AA",X"EF",X"AA",X"F1",X"AA",X"E1",X"AA",X"11",
		X"11",X"1F",X"11",X"1E",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FA",X"AA",X"FE",X"AA",X"1F",X"AA",X"1E",X"AA",
		X"FA",X"AA",X"FE",X"AA",X"1F",X"AA",X"1E",X"AA",X"11",X"AA",X"11",X"AA",X"11",X"FA",X"11",X"FE",
		X"11",X"AA",X"11",X"AA",X"11",X"FA",X"11",X"FE",X"11",X"1F",X"11",X"1E",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"FF",X"FF",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"FF",X"FF",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"FF",X"FF",X"EE",X"EE",X"EE",X"EE",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AE",X"AA",X"DE",X"AA",X"EE",
		X"AA",X"AA",X"AA",X"AA",X"EA",X"AA",X"ED",X"AA",X"EE",X"AA",X"EE",X"AA",X"EE",X"AA",X"EE",X"AA",
		X"AA",X"EE",X"AA",X"EE",X"AA",X"EE",X"AE",X"EE",X"AF",X"FF",X"AF",X"DD",X"AF",X"DD",X"AF",X"FF",
		X"EE",X"EA",X"EE",X"ED",X"EE",X"EE",X"EE",X"EE",X"FF",X"FF",X"DD",X"DD",X"DD",X"DD",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FF",X"AA",X"EE",X"AE",X"EE",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FF",X"FF",X"EE",X"EE",X"EE",X"EE",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"FF",X"FF",X"DD",X"DD",X"DD",X"DD",X"FF",X"FF",
		X"11",X"11",X"11",X"11",X"11",X"12",X"11",X"2A",X"11",X"AA",X"11",X"AA",X"12",X"AA",X"2A",X"AA",
		X"21",X"11",X"A2",X"11",X"AA",X"11",X"AA",X"11",X"AA",X"21",X"AA",X"A2",X"AA",X"AA",X"AA",X"AA",
		X"DD",X"DD",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"00",X"D1",X"00",X"11",X"DD",X"11",
		X"00",X"11",X"0D",X"11",X"D1",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",
		X"00",X"00",X"00",X"0D",X"00",X"D1",X"00",X"11",X"0D",X"11",X"D1",X"11",X"11",X"11",X"11",X"11",
		X"11",X"D0",X"11",X"1D",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"00",X"11",X"00",X"11",X"D0",X"11",X"1D",X"11",X"11",
		X"D0",X"00",X"1D",X"00",X"11",X"00",X"11",X"DD",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"1D",X"00",X"11",X"00",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"FF",X"FF",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"22",X"22",
		X"21",X"11",X"21",X"11",X"21",X"11",X"21",X"11",X"21",X"11",X"21",X"11",X"21",X"11",X"22",X"22",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"22",X"22",
		X"DD",X"DD",X"EE",X"EE",X"EE",X"EE",X"DD",X"DD",X"EE",X"EE",X"EE",X"EF",X"DD",X"DF",X"EE",X"EA",
		X"DD",X"88",X"E8",X"C8",X"28",X"CC",X"2A",X"AC",X"2A",X"AA",X"FF",X"CA",X"CA",X"CF",X"AA",X"FF",
		X"EE",X"A2",X"DD",X"DA",X"EE",X"22",X"EE",X"2A",X"DD",X"55",X"EE",X"5F",X"EE",X"C5",X"DD",X"CC",
		X"AB",X"FC",X"BB",X"FB",X"BB",X"CF",X"AA",X"FE",X"AC",X"FC",X"AB",X"FF",X"CC",X"EF",X"EE",X"EE",
		X"2A",X"AA",X"52",X"BA",X"5F",X"FF",X"5C",X"CF",X"5A",X"AA",X"52",X"AB",X"CA",X"AA",X"FF",X"BB",
		X"22",X"55",X"22",X"99",X"B2",X"99",X"BF",X"9F",X"2C",X"CF",X"B9",X"99",X"C2",X"99",X"28",X"98",
		X"FE",X"BB",X"FB",X"BC",X"EB",X"FB",X"2B",X"CB",X"CB",X"FB",X"C2",X"FF",X"BB",X"BB",X"CB",X"FB",
		X"48",X"9E",X"C2",X"9C",X"44",X"EE",X"4E",X"EE",X"4C",X"CE",X"2E",X"EE",X"44",X"EE",X"48",X"EE",
		X"22",X"FB",X"CC",X"FB",X"CC",X"BB",X"FC",X"B4",X"CF",X"AA",X"CF",X"BB",X"FF",X"BB",X"EE",X"FA",
		X"EE",X"EE",X"CC",X"EC",X"BE",X"EE",X"EE",X"EE",X"EE",X"EE",X"AA",X"EE",X"AB",X"EE",X"AA",X"E2",
		X"FF",X"FA",X"CC",X"FA",X"FF",X"CA",X"FF",X"AA",X"F1",X"2B",X"22",X"AA",X"22",X"1A",X"22",X"21",
		X"FA",X"B2",X"FA",X"B9",X"FA",X"99",X"AA",X"FF",X"AB",X"FC",X"BB",X"FF",X"BA",X"95",X"BA",X"29",
		X"12",X"12",X"22",X"12",X"1F",X"FF",X"FF",X"F2",X"FF",X"FB",X"11",X"2F",X"22",X"FF",X"12",X"2F",
		X"1F",X"BB",X"1B",X"BB",X"BB",X"B2",X"BB",X"2B",X"BB",X"F2",X"1B",X"AA",X"BA",X"FF",X"BA",X"FF",
		X"1C",X"FC",X"CA",X"FC",X"1C",X"CC",X"CC",X"FF",X"CC",X"F2",X"11",X"CB",X"CC",X"C1",X"11",X"CB",
		X"BE",X"FE",X"E2",X"FE",X"1E",X"EE",X"EE",X"EE",X"EE",X"2E",X"1E",X"2E",X"E1",X"EE",X"EE",X"EE",
		X"12",X"12",X"22",X"12",X"12",X"FF",X"FF",X"F2",X"FF",X"F2",X"FF",X"2F",X"22",X"FF",X"1C",X"2C",
		X"1F",X"BB",X"1B",X"B2",X"BB",X"2B",X"BB",X"F2",X"BB",X"AB",X"1B",X"AA",X"BA",X"FF",X"BE",X"FE",
		X"CA",X"FC",X"1C",X"CC",X"CC",X"FF",X"CC",X"F2",X"1C",X"CC",X"C1",X"2A",X"1C",X"CA",X"11",X"CA",
		X"E2",X"FE",X"1E",X"EE",X"1E",X"EE",X"EE",X"2E",X"EE",X"2E",X"1E",X"EE",X"11",X"EE",X"1E",X"2E",
		X"DE",X"AE",X"DE",X"EE",X"EF",X"EE",X"EE",X"E2",X"EE",X"2E",X"DE",X"2E",X"EE",X"EE",X"DE",X"EE",
		X"D4",X"55",X"43",X"FF",X"35",X"F2",X"35",X"75",X"DD",X"55",X"D3",X"55",X"35",X"55",X"32",X"22",
		X"DC",X"CC",X"CC",X"CC",X"C1",X"C1",X"1F",X"FF",X"12",X"2F",X"21",X"81",X"B2",X"11",X"11",X"11",
		X"32",X"22",X"DF",X"FF",X"FF",X"FF",X"F2",X"22",X"F2",X"A2",X"DF",X"FF",X"2D",X"F2",X"22",X"F2",
		X"AE",X"AE",X"AE",X"EE",X"EF",X"E2",X"EE",X"2E",X"EE",X"2E",X"DE",X"ED",X"EE",X"EE",X"EC",X"CC",
		X"DD",X"55",X"D3",X"FF",X"35",X"2F",X"35",X"75",X"DD",X"55",X"D3",X"55",X"35",X"55",X"D2",X"92",
		X"CC",X"CC",X"CC",X"1C",X"11",X"1F",X"11",X"1F",X"C1",X"77",X"C1",X"11",X"D1",X"11",X"B1",X"BB",
		X"D2",X"92",X"DF",X"FF",X"FF",X"FF",X"FF",X"F2",X"FF",X"FA",X"2D",X"2F",X"22",X"FF",X"D2",X"FF",
		X"DD",X"DD",X"EE",X"EE",X"EE",X"EE",X"DD",X"DD",X"EE",X"EE",X"EE",X"EE",X"DD",X"DF",X"EE",X"EF",
		X"DD",X"86",X"E2",X"85",X"22",X"CC",X"22",X"AA",X"2A",X"AA",X"2A",X"CA",X"FA",X"FF",X"CA",X"CF",
		X"EE",X"EA",X"DD",X"D2",X"EE",X"AA",X"EE",X"22",X"DD",X"55",X"EE",X"55",X"EE",X"5F",X"DD",X"CC",
		X"AA",X"CF",X"AB",X"FC",X"BB",X"EF",X"BB",X"CF",X"AB",X"FF",X"AB",X"FF",X"CC",X"EF",X"EE",X"EE",
		X"22",X"2A",X"82",X"BA",X"8F",X"AF",X"8F",X"AC",X"2A",X"CA",X"22",X"AB",X"CA",X"AA",X"FF",X"AA",
		X"22",X"BB",X"22",X"99",X"B2",X"99",X"BF",X"FF",X"2C",X"CF",X"29",X"99",X"B2",X"99",X"28",X"98",
		X"FE",X"BB",X"FE",X"BB",X"EB",X"BC",X"2B",X"FB",X"CB",X"CB",X"C2",X"FB",X"CC",X"FF",X"BB",X"BB",
		X"28",X"E9",X"42",X"E9",X"C4",X"EE",X"4E",X"EE",X"4E",X"EC",X"2E",X"EE",X"44",X"EE",X"28",X"EE",
		X"FF",X"77",X"FF",X"77",X"FF",X"17",X"2F",X"77",X"19",X"77",X"11",X"19",X"11",X"18",X"19",X"98",
		X"77",X"2B",X"77",X"BB",X"77",X"1F",X"27",X"B2",X"77",X"FF",X"CC",X"FC",X"CC",X"CC",X"CC",X"CC",
		X"9F",X"99",X"92",X"99",X"92",X"99",X"19",X"98",X"E9",X"88",X"E9",X"99",X"E9",X"98",X"18",X"88",
		X"FF",X"CC",X"FF",X"FF",X"2F",X"FF",X"AC",X"FF",X"C2",X"AA",X"CC",X"CC",X"CC",X"CC",X"1C",X"AA",
		X"2B",X"BB",X"BB",X"BA",X"BB",X"AA",X"BB",X"BA",X"FB",X"AA",X"FF",X"BA",X"FF",X"BA",X"FF",X"B4",
		X"1F",X"2F",X"F2",X"2F",X"F2",X"FF",X"1F",X"22",X"11",X"FE",X"11",X"FF",X"11",X"FF",X"44",X"FF",
		X"FF",X"44",X"FB",X"44",X"AB",X"44",X"A4",X"44",X"A4",X"44",X"14",X"44",X"C1",X"4C",X"1C",X"CC",
		X"44",X"FF",X"94",X"CC",X"94",X"AA",X"44",X"AC",X"44",X"CC",X"4C",X"FC",X"4C",X"FF",X"4C",X"FF",
		X"25",X"5E",X"11",X"5E",X"22",X"5C",X"22",X"15",X"22",X"21",X"22",X"22",X"22",X"22",X"22",X"22",
		X"EC",X"EE",X"EE",X"EC",X"EE",X"EC",X"EE",X"FF",X"EE",X"FC",X"EE",X"FC",X"1E",X"2F",X"21",X"CC",
		X"FF",X"FF",X"FD",X"DD",X"FD",X"DD",X"FD",X"DD",X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"22",X"2C",X"22",X"11",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"FF",X"CC",X"F4",X"CC",X"F4",X"FF",X"44",X"CC",X"EA",X"BC",X"AB",X"FF",X"AB",X"EE",X"FF",
		X"4E",X"EE",X"EE",X"EE",X"CC",X"EC",X"4E",X"EE",X"42",X"EE",X"2A",X"EE",X"2A",X"AE",X"AA",X"AE",
		X"FF",X"FF",X"FC",X"CF",X"FC",X"AC",X"CC",X"AA",X"11",X"2B",X"22",X"BA",X"22",X"1A",X"22",X"21",
		X"FF",X"BD",X"FF",X"B9",X"FF",X"99",X"AA",X"FF",X"AA",X"FF",X"BB",X"FC",X"AA",X"99",X"AA",X"25",
		X"22",X"BB",X"EB",X"BB",X"EC",X"CB",X"EF",X"BB",X"EC",X"BB",X"E2",X"44",X"BF",X"BB",X"2F",X"BC",
		X"2A",X"AA",X"4A",X"AA",X"CC",X"FF",X"4C",X"FF",X"FF",X"FF",X"FC",X"CC",X"FB",X"BC",X"FC",X"FC",
		X"2F",X"FB",X"99",X"FB",X"99",X"FB",X"FF",X"84",X"FF",X"E8",X"FF",X"CE",X"9E",X"EE",X"5E",X"EE",
		X"4F",X"FF",X"2C",X"FF",X"CC",X"FF",X"2C",X"FC",X"EE",X"FF",X"CE",X"FF",X"CC",X"FF",X"CC",X"AA",
		X"22",X"88",X"CC",X"AA",X"CC",X"A8",X"CC",X"88",X"CC",X"88",X"FF",X"FB",X"FF",X"BB",X"FF",X"BB",
		X"8A",X"CA",X"8C",X"AB",X"8C",X"AA",X"8A",X"AA",X"8A",X"AA",X"44",X"AA",X"B4",X"AA",X"BB",X"4B",
		X"F2",X"BB",X"FB",X"BB",X"2B",X"BB",X"2B",X"FB",X"2B",X"FC",X"22",X"CC",X"22",X"FF",X"2B",X"FF",
		X"BB",X"4B",X"BB",X"44",X"BB",X"44",X"BB",X"44",X"BB",X"44",X"BB",X"44",X"44",X"22",X"BB",X"42",
		X"22",X"BB",X"EC",X"BC",X"EF",X"BB",X"EC",X"BB",X"E2",X"BB",X"EF",X"4C",X"BF",X"BC",X"2F",X"FB",
		X"2A",X"AA",X"4A",X"AA",X"CC",X"FF",X"4C",X"FF",X"FF",X"FF",X"CC",X"CC",X"BC",X"CC",X"CF",X"CC",
		X"2F",X"FB",X"99",X"FB",X"99",X"FB",X"FF",X"84",X"FF",X"98",X"FF",X"EE",X"99",X"CE",X"59",X"EE",
		X"4F",X"FF",X"CC",X"FF",X"2C",X"EE",X"2C",X"FC",X"CF",X"FF",X"EE",X"FF",X"CC",X"FF",X"CE",X"BB",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"DC",X"C3",X"1D",X"33",X"11",X"32",X"11",X"DD",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"33",X"CC",X"33",X"CD",X"33",X"D1",X"32",X"11",X"3D",X"11",X"D1",X"11",X"11",X"11",X"11",X"11",
		X"1D",X"22",X"12",X"22",X"12",X"22",X"12",X"22",X"12",X"22",X"12",X"22",X"12",X"22",X"12",X"22",
		X"EE",X"EE",X"EE",X"EE",X"DE",X"CE",X"ED",X"CE",X"EE",X"EE",X"DE",X"EE",X"1D",X"EE",X"21",X"EE",
		X"EE",X"CB",X"EE",X"CC",X"EE",X"BB",X"EE",X"BA",X"ED",X"FF",X"DD",X"FF",X"ED",X"CA",X"DD",X"AC",
		X"22",X"EE",X"22",X"1E",X"22",X"21",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"D2",X"AA",X"ED",X"AB",X"DB",X"BA",X"DD",X"AA",X"11",X"AA",X"22",X"AA",X"22",X"1A",X"22",X"21",
		X"F2",X"AC",X"BB",X"C4",X"AA",X"C4",X"AA",X"BC",X"FF",X"AB",X"FF",X"AB",X"FF",X"AA",X"FF",X"AA",
		X"BB",X"B4",X"AB",X"44",X"A2",X"44",X"A2",X"44",X"2C",X"C2",X"CC",X"CF",X"CC",X"FF",X"CC",X"FF",
		X"FF",X"AA",X"AA",X"AB",X"AA",X"B2",X"BB",X"BB",X"AA",X"BB",X"AA",X"AB",X"CA",X"CB",X"CA",X"AB",
		X"FF",X"FF",X"FC",X"FC",X"CC",X"FC",X"CC",X"FC",X"FC",X"FF",X"FF",X"CF",X"2F",X"FF",X"A2",X"FE",
		X"AA",X"A8",X"C2",X"8A",X"C2",X"A8",X"CC",X"88",X"CC",X"88",X"FF",X"FB",X"FF",X"BB",X"FF",X"BB",
		X"8A",X"CC",X"8B",X"AA",X"8C",X"AA",X"88",X"AA",X"88",X"AA",X"44",X"AA",X"B4",X"AA",X"BB",X"4B",
		X"F2",X"BB",X"FB",X"BB",X"2B",X"FB",X"2B",X"FC",X"2B",X"CC",X"22",X"BB",X"22",X"FF",X"2B",X"FF",
		X"BB",X"4B",X"BB",X"C4",X"BB",X"44",X"BB",X"44",X"BB",X"44",X"BB",X"44",X"44",X"42",X"BB",X"42",
		X"EE",X"EE",X"EC",X"EC",X"EE",X"EE",X"EE",X"EE",X"DE",X"EE",X"ED",X"ED",X"1E",X"EE",X"21",X"EE",
		X"E2",X"CB",X"ED",X"CB",X"DD",X"BA",X"DD",X"AA",X"DE",X"FF",X"EE",X"FF",X"EE",X"FF",X"DD",X"CF",
		X"22",X"EE",X"22",X"1E",X"22",X"21",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"D2",X"AC",X"BA",X"AB",X"DB",X"BA",X"D2",X"AA",X"11",X"AA",X"22",X"AA",X"22",X"1A",X"22",X"21",
		X"22",X"CA",X"BB",X"44",X"AA",X"44",X"AA",X"B4",X"FF",X"BB",X"FF",X"AB",X"FF",X"AA",X"FF",X"AA",
		X"BB",X"B4",X"BB",X"44",X"22",X"C4",X"2C",X"CC",X"2C",X"CC",X"2C",X"FF",X"2C",X"FF",X"FF",X"FF",
		X"FA",X"AA",X"AA",X"AB",X"AA",X"B2",X"BB",X"BB",X"AA",X"BC",X"AA",X"CB",X"AB",X"AB",X"AA",X"AB",
		X"FC",X"FC",X"CC",X"FC",X"CB",X"FC",X"CC",X"FF",X"FF",X"CF",X"FF",X"FC",X"AF",X"FF",X"B2",X"FE",
		X"AC",X"AB",X"1A",X"AC",X"21",X"AB",X"22",X"AB",X"22",X"11",X"22",X"22",X"22",X"22",X"22",X"22",
		X"CC",X"FF",X"CC",X"FF",X"CC",X"FF",X"CC",X"FF",X"2F",X"FF",X"CC",X"FF",X"1C",X"FF",X"21",X"FF",
		X"FF",X"FF",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"22",X"FF",X"22",X"1F",X"22",X"21",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"33",X"00",X"33",X"03",X"33",X"03",X"33",X"3F",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"3F",X"33",X"3F",X"33",X"3F",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"33",X"00",X"33",X"2C",X"33",X"32",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"C0",X"00",X"C0",X"00",X"2C",X"00",X"2C",X"00",X"2C",X"00",X"22",X"00",X"22",X"00",X"22",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"33",X"03",X"33",X"3F",X"33",X"FF",X"33",X"FF",X"33",X"F3",X"33",X"F3",X"33",
		X"00",X"00",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"33",X"00",X"33",X"30",X"33",X"03",X"33",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"2C",X"00",X"33",X"00",X"33",X"C0",X"33",X"2C",X"33",X"2C",X"33",X"22",X"33",X"22",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"32",X"33",X"32",X"33",X"32",X"33",X"32",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"2C",X"00",
		X"00",X"33",X"00",X"33",X"00",X"3C",X"03",X"C0",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"0B",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"B3",X"33",X"BB",X"33",X"CC",X"33",X"00",X"33",X"00",X"CC",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"22",X"C0",X"22",X"2C",X"2C",X"22",X"22",X"C2",X"22",X"0C",X"22",X"00",X"22",X"00",X"2C",X"00",
		X"33",X"33",X"33",X"33",X"33",X"32",X"33",X"32",X"33",X"22",X"33",X"2C",X"23",X"C0",X"22",X"00",
		X"2B",X"00",X"2B",X"00",X"BB",X"00",X"BC",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"3C",X"00",X"C3",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"B3",X"00",X"B3",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"B3",X"00",X"BB",X"00",X"CB",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"C3",X"33",X"0C",X"33",X"00",X"22",X"00",X"CC",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"32",X"33",X"32",X"33",X"32",X"33",X"22",
		X"22",X"00",X"22",X"00",X"C2",X"00",X"CC",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",
		X"33",X"22",X"33",X"22",X"33",X"22",X"33",X"22",X"23",X"2B",X"22",X"CC",X"22",X"00",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"BC",X"00",X"BB",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"00",X"33",X"00",X"F3",X"03",X"33",X"03",X"33",X"3F",X"33",X"3F",X"33",X"3F",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"30",X"33",
		X"3F",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"33",X"00",X"33",X"2C",X"33",X"32",X"33",X"32",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"2C",X"00",X"2C",X"00",X"2C",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"3F",X"00",X"F3",X"00",X"33",X"03",X"33",X"03",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"33",X"C0",X"33",X"32",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"2C",X"00",X"2C",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"2C",X"00",X"22",X"00",X"22",X"00",X"32",X"00",X"32",X"00",X"32",X"00",X"32",X"00",X"32",X"C0",
		X"C3",X"33",X"0C",X"33",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"0B",X"00",X"0B",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"B3",X"33",X"BB",X"33",X"CC",X"33",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"22",X"22",X"2C",X"2C",X"22",X"C0",X"22",X"00",X"22",X"00",X"22",X"00",X"2C",X"00",X"2C",X"00",
		X"33",X"32",X"33",X"32",X"33",X"22",X"22",X"2C",X"22",X"C0",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"BB",X"00",X"BB",X"00",X"BB",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"00",X"33",X"00",X"33",X"00",X"3C",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"CC",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"B3",X"33",X"B3",X"33",X"BB",X"33",X"CC",X"22",X"00",X"CC",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"32",X"22",X"3C",X"22",X"32",X"CC",X"32",X"00",X"32",X"00",X"22",X"00",X"22",X"C0",X"22",X"BC",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"32",X"23",X"2C",X"22",X"C0",X"CC",X"00",
		X"22",X"C0",X"2B",X"00",X"BB",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"33",X"00",X"F3",X"03",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",
		X"33",X"33",X"3F",X"33",X"3F",X"33",X"3F",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"33",X"2C",X"33",X"22",X"33",X"32",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"C0",X"00",X"C0",X"00",X"2C",X"00",X"2C",X"00",X"2C",X"00",X"22",X"00",X"22",X"00",X"22",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"33",X"00",X"F3",X"03",X"33",X"03",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"33",X"3F",X"33",X"3F",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"33",X"00",X"33",X"2C",X"33",X"32",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"C0",X"00",X"C0",X"00",X"2C",X"00",X"2C",X"00",X"2C",X"02",X"22",X"22",X"22",X"22",X"22",X"2C",
		X"00",X"33",X"00",X"33",X"00",X"C3",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"0B",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"BF",X"33",X"CC",X"22",X"00",X"FF",X"00",X"CC",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"2C",X"C0",X"22",X"C0",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",
		X"33",X"33",X"33",X"33",X"33",X"32",X"33",X"22",X"23",X"22",X"C2",X"FC",X"FF",X"C0",X"CC",X"00",
		X"2C",X"00",X"2B",X"00",X"2B",X"00",X"BC",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"00",X"33",X"00",X"33",X"00",X"3C",X"03",X"C0",X"0C",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"0B",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"B3",X"33",X"BB",X"33",X"CC",X"33",X"00",X"33",X"00",X"CC",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"22",X"2C",X"22",X"C0",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"2C",X"00",
		X"33",X"33",X"33",X"33",X"33",X"32",X"33",X"32",X"33",X"22",X"33",X"2C",X"23",X"C0",X"22",X"00",
		X"2B",X"00",X"2B",X"00",X"BB",X"00",X"BC",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"33",X"00",X"F3",X"03",X"33",X"03",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"3F",X"33",X"3F",X"33",X"3F",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"33",X"2C",X"33",X"32",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"C0",X"00",X"C0",X"00",X"2C",X"00",X"2C",X"00",X"2C",X"00",X"22",X"20",X"22",X"2C",X"22",X"2C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"33",X"03",X"F3",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"33",X"3F",X"33",X"3F",X"33",X"3F",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"32",X"00",X"33",X"C0",X"33",X"2C",X"33",X"32",X"33",X"32",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"C0",X"00",X"C0",X"00",X"2C",X"00",X"2C",X"00",X"2C",X"00",X"22",X"00",X"22",X"00",X"2C",X"C0",
		X"00",X"00",X"00",X"03",X"00",X"33",X"00",X"33",X"00",X"3C",X"00",X"C0",X"00",X"00",X"00",X"0B",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"BB",X"00",X"CB",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"B3",X"33",X"CC",X"33",X"00",X"33",X"00",X"33",X"00",X"CC",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"2C",X"C0",X"22",X"C0",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"2C",X"00",
		X"33",X"33",X"33",X"33",X"33",X"32",X"33",X"32",X"33",X"22",X"33",X"2C",X"23",X"C0",X"22",X"00",
		X"2B",X"00",X"2B",X"00",X"BB",X"00",X"BC",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",X"00",X"33",X"00",X"3C",X"00",X"C0",X"00",X"00",
		X"33",X"33",X"33",X"33",X"23",X"33",X"C3",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"F3",X"33",X"BF",X"33",X"BB",X"33",X"CC",X"F3",X"00",X"CC",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"22",X"C0",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",
		X"33",X"33",X"33",X"33",X"33",X"32",X"33",X"32",X"33",X"22",X"33",X"22",X"22",X"22",X"C2",X"2C",
		X"2B",X"00",X"2B",X"00",X"2B",X"00",X"BC",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"00",X"33",X"03",X"F3",X"33",X"33",X"3F",X"33",X"33",X"33",X"33",X"F3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",
		X"33",X"FF",X"3F",X"FF",X"3F",X"CC",X"3F",X"CC",X"3F",X"FB",X"3F",X"BB",X"33",X"CC",X"33",X"FF",
		X"00",X"00",X"32",X"00",X"33",X"22",X"33",X"32",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"F3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"2C",X"00",X"2C",X"00",
		X"33",X"FF",X"33",X"FF",X"33",X"FF",X"33",X"FF",X"BB",X"FF",X"BB",X"BF",X"BB",X"FF",X"CC",X"33",
		X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"00",X"33",X"03",X"F3",X"33",X"33",X"3F",X"33",X"33",X"33",X"33",X"F3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",X"33",X"03",X"C3",X"03",X"0C",X"33",
		X"3F",X"FF",X"3F",X"CF",X"FF",X"CC",X"FF",X"FF",X"FF",X"FB",X"FF",X"BC",X"3F",X"BC",X"33",X"FB",
		X"00",X"00",X"32",X"00",X"33",X"22",X"33",X"32",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"2C",X"00",X"2C",X"00",
		X"33",X"FF",X"FF",X"CF",X"FF",X"CC",X"BF",X"FC",X"CB",X"FF",X"CC",X"BF",X"CC",X"CF",X"CC",X"F3",
		X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"22",X"22",X"22",
		X"00",X"03",X"00",X"33",X"00",X"33",X"00",X"22",X"03",X"CC",X"0C",X"00",X"00",X"00",X"00",X"00",
		X"33",X"FF",X"33",X"FF",X"33",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"FF",X"32",X"FF",X"32",X"FF",X"BB",X"FF",X"BB",X"FF",X"BB",X"CC",X"CC",X"C0",X"00",X"00",
		X"CF",X"F3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"22",X"00",X"22",X"00",X"22",X"20",X"2C",X"22",X"22",X"C2",X"22",X"0C",X"22",X"00",X"2C",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"FF",X"BB",X"CC",X"BB",X"00",X"CC",X"00",X"00",
		X"2C",X"00",X"2C",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"BC",X"00",X"C0",X"00",X"00",X"00",
		X"00",X"33",X"00",X"33",X"00",X"C3",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"FC",X"33",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",
		X"00",X"00",X"00",X"0B",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BC",X"FF",X"BB",X"FF",X"BB",X"FF",X"BB",X"FF",X"BB",X"FF",X"CC",X"22",X"00",X"CC",X"00",X"00",
		X"BB",X"FF",X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"22",X"2C",X"22",X"C0",X"22",X"00",X"2C",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"BC",X"00",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"CB",X"FF",X"CB",X"FF",X"FC",X"22",X"C0",X"C2",X"00",X"0C",X"00",
		X"BB",X"00",X"BB",X"00",X"BB",X"00",X"BC",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"33",X"03",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"3F",X"33",X"3F",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"C0",X"00",X"C0",X"00",X"2C",X"00",X"2C",X"00",X"22",X"00",X"22",X"00",X"22",X"03",X"22",X"22",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"0B",X"00",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"B0",X"0F",X"B0",X"FF",X"CF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",X"00",X"0C",X"03",X"00",X"33",
		X"3F",X"FF",X"3F",X"FF",X"33",X"FF",X"33",X"FC",X"33",X"BB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"FC",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"BC",X"00",
		X"FF",X"FF",X"FF",X"FF",X"BB",X"FF",X"CC",X"F3",X"BB",X"F3",X"BB",X"FF",X"3F",X"FF",X"3F",X"FF",
		X"C0",X"00",X"C0",X"00",X"3C",X"00",X"32",X"00",X"32",X"00",X"32",X"03",X"33",X"22",X"33",X"22",
		X"00",X"33",X"00",X"CC",X"00",X"0B",X"00",X"0B",X"00",X"0B",X"00",X"0C",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C3",X"33",X"0C",X"33",X"00",X"33",X"00",X"C2",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"32",
		X"22",X"C0",X"22",X"00",X"22",X"00",X"22",X"00",X"2B",X"00",X"2B",X"00",X"2C",X"00",X"C0",X"00",
		X"33",X"22",X"23",X"22",X"22",X"CC",X"22",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"33",X"00",X"33",X"00",X"C3",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"0C",X"00",X"00",
		X"FC",X"F3",X"FF",X"F3",X"FF",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"23",X"33",X"22",X"33",X"C2",X"33",X"0C",X"22",X"00",X"CC",X"00",X"00",X"0F",X"00",
		X"33",X"FC",X"33",X"FF",X"33",X"FF",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"32",X"2C",X"32",X"C0",X"32",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"0F",
		X"33",X"32",X"33",X"22",X"33",X"22",X"22",X"22",X"22",X"2C",X"22",X"C0",X"CC",X"00",X"00",X"0F",
		X"2C",X"00",X"2C",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0B",X"00",X"BB",X"00",X"BB",X"00",X"CB",X"00",X"0C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"B0",X"00",X"B0",X"00",X"BB",X"0F",X"BB",X"FF",X"BC",X"FF",X"CF",X"FF",X"3F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"33",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"FB",X"33",X"BC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"B0",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"CC",X"00",X"C0",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"FF",X"CB",X"FF",X"CC",X"FF",X"CC",X"BF",
		X"C0",X"00",X"3C",X"00",X"3C",X"00",X"F3",X"00",X"F3",X"00",X"33",X"00",X"33",X"00",X"33",X"2C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"BB",X"00",X"BB",X"0F",X"BB",X"FF",X"BC",X"FF",X"CF",X"FF",X"3F",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"C3",X"03",X"0C",X"33",X"00",X"33",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"FB",X"FF",X"FB",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"B0",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"CC",X"00",X"C0",X"00",X"C0",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"FF",X"BB",X"FF",X"CC",X"FF",X"CC",X"FF",
		X"3C",X"00",X"3C",X"00",X"F2",X"00",X"F2",X"00",X"F2",X"00",X"33",X"22",X"33",X"22",X"33",X"2C",
		X"00",X"33",X"03",X"C3",X"03",X"33",X"33",X"33",X"3C",X"C3",X"C0",X"03",X"00",X"03",X"00",X"0C",
		X"3F",X"BC",X"FF",X"FB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"F3",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"C2",X"33",X"0C",X"22",X"00",X"CC",X"00",X"00",
		X"CC",X"FF",X"BB",X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FF",X"FC",X"3F",X"FF",X"33",X"FF",
		X"33",X"22",X"F3",X"22",X"F3",X"C2",X"F2",X"CC",X"F2",X"00",X"F2",X"00",X"22",X"00",X"22",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"22",X"33",X"22",X"22",X"2C",X"22",X"C0",X"CC",X"00",
		X"22",X"00",X"2C",X"00",X"2C",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"C3",X"00",X"03",X"00",X"03",X"00",X"0C",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CC",X"FF",X"CC",X"FF",X"FF",X"FF",X"FF",X"F3",X"33",X"33",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"C2",X"33",X"0C",X"22",X"00",X"CC",X"00",X"00",X"00",X"00",
		X"BB",X"FF",X"FF",X"CF",X"FF",X"FF",X"FF",X"FF",X"33",X"FF",X"33",X"33",X"33",X"33",X"33",X"33",
		X"33",X"C0",X"33",X"C0",X"32",X"C0",X"32",X"00",X"32",X"00",X"22",X"00",X"22",X"00",X"22",X"00",
		X"33",X"33",X"33",X"33",X"33",X"22",X"33",X"22",X"22",X"2C",X"22",X"C0",X"CC",X"00",X"00",X"00",
		X"2C",X"00",X"2C",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"33",X"00",X"F3",X"03",X"33",X"03",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"3F",X"33",X"3F",X"33",X"3F",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"33",X"00",X"33",X"3C",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"C0",X"00",X"C0",X"00",X"2C",X"00",X"2C",X"00",X"2C",X"00",X"22",X"00",X"22",X"00",X"22",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"00",X"33",X"00",X"F3",X"03",X"33",X"03",X"33",X"33",X"33",X"3F",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"33",X"00",X"33",
		X"3F",X"33",X"3F",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"33",X"00",X"33",X"3C",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"C0",X"00",X"2C",X"00",X"2C",X"00",X"2C",X"00",X"22",X"00",X"22",X"02",X"22",X"22",X"22",X"2C",
		X"00",X"33",X"00",X"33",X"00",X"3C",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"0B",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"B3",X"33",X"BB",X"33",X"CC",X"33",X"00",X"CC",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"22",X"C0",X"22",X"2C",X"2C",X"2C",X"22",X"22",X"22",X"C2",X"22",X"0C",X"22",X"00",X"2C",X"00",
		X"33",X"33",X"33",X"32",X"33",X"22",X"33",X"22",X"23",X"22",X"C2",X"CC",X"C2",X"00",X"0C",X"00",
		X"2B",X"00",X"2B",X"00",X"BB",X"00",X"BC",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C3",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"BE",X"33",X"BB",X"33",X"BB",X"FF",X"CC",X"CC",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"22",X"00",X"2C",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"2C",X"00",X"2C",X"00",
		X"33",X"33",X"23",X"32",X"C2",X"22",X"F2",X"FF",X"FF",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"2C",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"11",X"11",X"BB",X"11",X"2B",X"A1",X"FF",X"FF",X"44",X"44",X"44",X"44",X"FF",X"FF",X"33",X"33",
		X"21",X"11",X"2F",X"21",X"FF",X"F1",X"2F",X"FF",X"BF",X"FF",X"F2",X"F1",X"FF",X"12",X"FF",X"21",
		X"33",X"33",X"FF",X"FF",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"FC",X"CC",X"FC",X"BC",X"FC",X"CC",X"FF",X"FC",X"F2",X"FC",X"FC",X"BB",X"FB",X"11",X"FC",X"CC",
		X"FD",X"DD",X"F1",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"88",X"11",X"87",X"71",X"FF",X"71",X"F2",X"71",X"87",X"AF",X"AA",X"F4",X"77",X"FF",X"44",X"33",
		X"DD",X"33",X"11",X"FF",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"77",X"33",X"44",X"33",X"44",X"33",X"74",X"33",X"94",X"33",X"44",X"33",X"CC",X"33",X"CC",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FA",X"FA",X"12",X"12",X"12",X"22",X"22",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FF",X"AA",X"22",X"1A",X"FF",X"22",X"22",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FF",X"FF",X"2F",X"FF",X"FF",X"2F",X"22",X"2A",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FF",X"FA",X"FF",X"FF",X"22",X"2F",X"2A",X"2A",X"AA",X"AA",
		X"11",X"22",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"11",X"22",X"22",X"22",
		X"21",X"22",X"11",X"22",X"21",X"22",X"21",X"22",X"21",X"22",X"21",X"22",X"21",X"22",X"22",X"22",
		X"11",X"22",X"22",X"12",X"22",X"12",X"11",X"22",X"12",X"22",X"12",X"22",X"11",X"12",X"22",X"22",
		X"11",X"22",X"12",X"12",X"22",X"12",X"22",X"22",X"22",X"12",X"12",X"12",X"11",X"22",X"22",X"22",
		X"22",X"22",X"21",X"22",X"12",X"22",X"22",X"22",X"22",X"22",X"11",X"12",X"22",X"22",X"22",X"22",
		X"11",X"12",X"12",X"22",X"11",X"22",X"22",X"12",X"22",X"12",X"12",X"12",X"11",X"22",X"22",X"22",
		X"11",X"22",X"12",X"12",X"12",X"22",X"11",X"22",X"12",X"12",X"12",X"12",X"11",X"22",X"22",X"22",
		X"11",X"12",X"22",X"12",X"22",X"22",X"21",X"22",X"21",X"22",X"21",X"22",X"21",X"22",X"22",X"22",
		X"11",X"22",X"12",X"12",X"12",X"12",X"11",X"22",X"12",X"12",X"12",X"12",X"11",X"22",X"22",X"22",
		X"11",X"22",X"12",X"12",X"12",X"12",X"11",X"12",X"22",X"12",X"12",X"12",X"11",X"22",X"22",X"22",
		X"33",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"0A",X"00",X"10",X"00",X"1A",X"00",X"AA",X"00",
		X"DD",X"DD",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"DD",X"D2",X"11",X"12",X"11",X"12",X"11",X"12",X"11",X"12",X"11",X"12",X"11",X"12",X"11",X"12",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FA",X"AF",X"2F",X"FF",X"2F",X"F2",X"2A",X"A2",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FA",X"FA",X"F2",X"F2",X"FF",X"F2",X"A2",X"A2",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FA",X"FF",X"F2",X"AF",X"F2",X"AF",X"A2",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FF",X"FF",X"FF",X"F2",X"FF",X"FF",X"A2",X"A2",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"33",
		X"00",X"00",X"10",X"A0",X"01",X"00",X"10",X"00",X"0A",X"00",X"A0",X"A0",X"00",X"00",X"00",X"00",
		X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"33",X"33",
		X"FF",X"FF",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"FF",X"FF",X"AA",X"22",X"AA",X"22",X"AA",X"22",
		X"FF",X"FF",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"FF",X"FF",X"AA",X"AA",X"2A",X"AA",X"2A",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"11",X"00",X"0A",X"00",
		X"22",X"AA",X"22",X"AA",X"22",X"AA",X"22",X"AA",X"22",X"2A",X"FF",X"FF",X"EE",X"EE",X"EE",X"EE",
		X"11",X"00",X"13",X"10",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"11",X"03",X"33",X"30",
		X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"03",X"00",
		X"11",X"00",X"33",X"10",X"00",X"13",X"11",X"33",X"13",X"30",X"13",X"00",X"11",X"10",X"33",X"33",
		X"11",X"00",X"33",X"10",X"00",X"13",X"01",X"33",X"00",X"10",X"00",X"13",X"11",X"33",X"33",X"30",
		X"01",X"00",X"11",X"30",X"01",X"30",X"31",X"30",X"01",X"30",X"11",X"10",X"31",X"33",X"00",X"30",
		X"11",X"10",X"13",X"33",X"11",X"00",X"33",X"10",X"30",X"13",X"00",X"13",X"11",X"33",X"33",X"30",
		X"11",X"00",X"13",X"10",X"13",X"03",X"11",X"00",X"13",X"10",X"13",X"13",X"11",X"03",X"33",X"30",
		X"11",X"10",X"33",X"13",X"01",X"33",X"01",X"30",X"11",X"30",X"11",X"00",X"11",X"00",X"03",X"00",
		X"11",X"00",X"13",X"10",X"13",X"13",X"11",X"03",X"13",X"10",X"13",X"13",X"11",X"03",X"33",X"30",
		X"11",X"00",X"33",X"10",X"00",X"13",X"11",X"13",X"33",X"13",X"00",X"13",X"11",X"33",X"33",X"30",
		X"AA",X"22",X"AA",X"22",X"A2",X"22",X"22",X"22",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"22",X"AA",X"22",X"AA",X"22",X"AA",X"22",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"11",X"10",X"11",X"1A",X"11",X"1A",X"AA",X"AA",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"00",X"AA",X"A0",X"11",X"00",X"AA",X"A0",X"00",X"00",X"00",X"00",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"11",X"00",X"AA",X"10",X"A0",X"1A",X"01",X"AA",X"11",X"A0",X"0A",X"00",X"11",X"00",X"0A",X"00",
		X"AA",X"22",X"A2",X"22",X"A2",X"22",X"22",X"22",X"22",X"22",X"FF",X"FF",X"EE",X"EE",X"EE",X"EE",
		X"11",X"00",X"AA",X"10",X"00",X"1A",X"00",X"1A",X"11",X"1A",X"AA",X"1A",X"00",X"1A",X"00",X"AA",
		X"11",X"00",X"1A",X"10",X"1A",X"1A",X"11",X"0A",X"1A",X"10",X"1A",X"1A",X"11",X"0A",X"AA",X"A0",
		X"11",X"00",X"1A",X"10",X"1A",X"0A",X"1A",X"00",X"1A",X"00",X"1A",X"10",X"11",X"0A",X"AA",X"A0",
		X"11",X"00",X"1A",X"10",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"11",X"0A",X"AA",X"A0",
		X"11",X"10",X"1A",X"AA",X"1A",X"00",X"11",X"10",X"1A",X"AA",X"1A",X"00",X"11",X"10",X"AA",X"AA",
		X"11",X"10",X"1A",X"AA",X"1A",X"00",X"11",X"10",X"1A",X"AA",X"1A",X"00",X"1A",X"00",X"AA",X"00",
		X"11",X"00",X"1A",X"10",X"1A",X"0A",X"1A",X"10",X"1A",X"1A",X"1A",X"1A",X"11",X"0A",X"AA",X"A0",
		X"10",X"10",X"1A",X"1A",X"1A",X"1A",X"11",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"AA",X"0A",
		X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"0A",X"00",
		X"01",X"00",X"01",X"A0",X"01",X"A0",X"01",X"A0",X"01",X"A0",X"01",X"A0",X"11",X"A0",X"AA",X"00",
		X"10",X"10",X"1A",X"0A",X"1A",X"A0",X"11",X"00",X"1A",X"00",X"1A",X"10",X"1A",X"1A",X"AA",X"AA",
		X"10",X"00",X"1A",X"00",X"1A",X"00",X"1A",X"00",X"1A",X"00",X"1A",X"00",X"11",X"10",X"AA",X"AA",
		X"11",X"10",X"11",X"1A",X"11",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"AA",X"0A",
		X"10",X"10",X"11",X"1A",X"11",X"1A",X"11",X"1A",X"11",X"1A",X"01",X"1A",X"00",X"1A",X"00",X"AA",
		X"11",X"00",X"1A",X"10",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"11",X"0A",X"AA",X"A0",
		X"11",X"00",X"1A",X"10",X"1A",X"1A",X"1A",X"1A",X"11",X"0A",X"1A",X"A0",X"1A",X"00",X"AA",X"00",
		X"11",X"00",X"1A",X"10",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"11",X"0A",X"AA",X"A0",
		X"11",X"00",X"1A",X"10",X"1A",X"1A",X"1A",X"1A",X"11",X"0A",X"1A",X"10",X"1A",X"1A",X"AA",X"0A",
		X"11",X"00",X"1A",X"10",X"1A",X"0A",X"11",X"00",X"AA",X"10",X"00",X"1A",X"11",X"AA",X"AA",X"A0",
		X"11",X"10",X"11",X"AA",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"0A",X"00",
		X"10",X"10",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"11",X"0A",X"AA",X"A0",
		X"10",X"10",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"0A",X"11",X"A0",X"0A",X"00",
		X"10",X"10",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"11",X"0A",X"AA",X"A0",
		X"10",X"10",X"1A",X"1A",X"1A",X"1A",X"11",X"0A",X"AA",X"10",X"00",X"1A",X"00",X"1A",X"00",X"AA",
		X"10",X"10",X"1A",X"1A",X"1A",X"1A",X"11",X"0A",X"11",X"A0",X"11",X"00",X"11",X"00",X"0A",X"00",
		X"11",X"10",X"AA",X"1A",X"01",X"AA",X"11",X"A0",X"11",X"00",X"1A",X"00",X"11",X"10",X"AA",X"AA",
		X"70",X"00",X"77",X"70",X"77",X"70",X"77",X"70",X"77",X"00",X"77",X"00",X"07",X"00",X"00",X"00",
		X"00",X"04",X"73",X"42",X"77",X"20",X"72",X"20",X"28",X"72",X"07",X"72",X"02",X"20",X"00",X"00",
		X"00",X"00",X"00",X"34",X"C0",X"24",X"CB",X"42",X"C2",X"20",X"2C",X"B0",X"2C",X"B0",X"02",X"20",
		X"00",X"00",X"CC",X"00",X"FC",X"00",X"CC",X"30",X"CC",X"B0",X"CC",X"00",X"BB",X"00",X"00",X"00",
		X"03",X"00",X"83",X"00",X"88",X"70",X"88",X"70",X"88",X"70",X"77",X"00",X"77",X"00",X"00",X"00",
		X"F2",X"F1",X"F2",X"2F",X"FF",X"2F",X"22",X"F1",X"EF",X"11",X"FF",X"11",X"FF",X"11",X"FF",X"44",
		X"BB",X"B2",X"AB",X"BB",X"AA",X"BB",X"AB",X"BB",X"AA",X"BF",X"AB",X"FF",X"AB",X"FF",X"4B",X"FF",
		X"FF",X"44",X"CC",X"49",X"AA",X"49",X"CA",X"44",X"CC",X"44",X"CF",X"C4",X"FF",X"C4",X"FF",X"C4",
		X"44",X"FF",X"44",X"BF",X"44",X"BA",X"44",X"4A",X"44",X"4A",X"44",X"41",X"C4",X"1C",X"CC",X"C1",
		X"B2",X"77",X"BB",X"77",X"F1",X"77",X"2B",X"72",X"FF",X"77",X"CF",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"77",X"FF",X"77",X"FF",X"71",X"FF",X"77",X"F2",X"77",X"91",X"91",X"11",X"81",X"11",X"89",X"91",
		X"CC",X"FF",X"FF",X"FF",X"FF",X"F2",X"FF",X"CA",X"AA",X"2C",X"CC",X"CC",X"CC",X"CC",X"AA",X"C1",
		X"99",X"F9",X"99",X"29",X"99",X"29",X"89",X"91",X"88",X"9E",X"99",X"9E",X"89",X"9E",X"88",X"81",
		X"22",X"2F",X"22",X"2F",X"22",X"F1",X"22",X"F1",X"22",X"11",X"22",X"11",X"22",X"11",X"22",X"11",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"F2",X"22",X"F2",X"22",X"1F",X"22",X"1F",X"22",
		X"2F",X"11",X"2F",X"11",X"F1",X"11",X"F1",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"22",X"11",X"22",X"11",X"22",X"11",X"22",X"11",X"F2",X"11",X"F2",X"11",X"1F",X"11",X"1F",
		X"22",X"DE",X"22",X"EE",X"22",X"EE",X"22",X"EE",X"22",X"EE",X"22",X"EE",X"2D",X"EE",X"2E",X"EE",
		X"22",X"22",X"22",X"22",X"D2",X"22",X"E2",X"22",X"ED",X"22",X"EE",X"22",X"EE",X"22",X"EE",X"22",
		X"DE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"FF",X"FF",X"DD",X"DD",X"DD",X"DD",X"FF",X"FF",
		X"EE",X"22",X"EE",X"22",X"EE",X"D2",X"EE",X"E2",X"FF",X"F2",X"DD",X"F2",X"DD",X"F2",X"FF",X"F2",
		X"AA",X"AF",X"AA",X"AF",X"AA",X"F1",X"AA",X"F1",X"AA",X"11",X"AA",X"11",X"AA",X"11",X"AA",X"11",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FA",X"AA",X"FA",X"AA",X"1F",X"AA",X"1F",X"AA",
		X"AF",X"11",X"AF",X"11",X"F1",X"11",X"F1",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"AA",X"11",X"AA",X"11",X"AA",X"11",X"AA",X"11",X"FA",X"11",X"FA",X"11",X"1F",X"11",X"1F",
		X"AA",X"AD",X"AA",X"AE",X"AA",X"DE",X"AA",X"EE",X"AA",X"EE",X"AA",X"EE",X"AA",X"EE",X"AA",X"EE",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"DA",X"AA",X"EA",X"AA",X"ED",X"AA",X"EE",X"AA",
		X"AD",X"EE",X"AE",X"EE",X"DE",X"EE",X"EE",X"EE",X"FF",X"FF",X"FD",X"DD",X"FD",X"DD",X"FF",X"FF",
		X"EE",X"AA",X"EE",X"AA",X"EE",X"AA",X"EE",X"AA",X"FF",X"AA",X"DD",X"AA",X"DD",X"AA",X"FF",X"AA",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"FF",X"FF",X"EE",X"EE",X"EE",X"EE",
		X"FF",X"FF",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"FF",X"FF",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"2D",X"22",X"2E",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"01",X"00",X"01",X"00",
		X"11",X"00",X"11",X"10",X"11",X"10",X"11",X"10",X"11",X"10",X"11",X"10",X"01",X"10",X"01",X"10",
		X"00",X"01",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"00",X"00",
		X"00",X"10",X"11",X"10",X"11",X"10",X"11",X"10",X"11",X"10",X"11",X"10",X"11",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AF",X"AA",X"EF",X"AA",X"F1",X"AA",X"E1",
		X"F1",X"11",X"E1",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"AA",X"11",X"AA",X"11",X"AF",X"11",X"EF",X"11",X"F1",X"11",X"E1",X"11",X"11",X"11",X"11",X"11",
		X"AA",X"AF",X"AA",X"EF",X"AA",X"F1",X"AA",X"E1",X"AA",X"11",X"AA",X"11",X"AF",X"11",X"EF",X"11",
		X"11",X"AA",X"11",X"FA",X"11",X"FE",X"11",X"1F",X"11",X"1E",X"11",X"11",X"11",X"11",X"11",X"11",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FA",X"AA",X"FE",X"AA",X"1F",X"AA",X"1E",X"AA",X"11",X"AA",
		X"FE",X"AA",X"1F",X"AA",X"1E",X"AA",X"11",X"AA",X"11",X"AA",X"11",X"FA",X"11",X"FE",X"11",X"1F",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"FF",X"FF",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"FF",X"FF",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"FF",X"FF",X"EE",X"EE",X"EE",X"EE",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AE",X"AA",X"DE",X"AA",X"EE",X"AA",X"EE",X"AA",X"EE",X"AA",X"EE",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"AA",X"ED",X"AA",X"EE",X"AA",
		X"AE",X"EE",X"DE",X"EE",X"EE",X"EE",X"EE",X"EE",X"FF",X"FF",X"DD",X"DD",X"DD",X"DD",X"FF",X"FF",
		X"EE",X"AA",X"EE",X"AA",X"EE",X"AA",X"EE",X"EA",X"FF",X"FA",X"DD",X"FA",X"DD",X"FA",X"FF",X"FA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FF",X"FF",X"EE",X"EE",X"EE",X"EE",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FF",X"AA",X"EE",X"AA",X"EE",X"EA",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"FF",X"FF",X"DD",X"DD",X"DD",X"DD",X"FF",X"FF",
		X"11",X"12",X"11",X"2A",X"11",X"AA",X"11",X"AA",X"12",X"AA",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"11",X"11",X"11",X"11",X"21",X"11",X"A2",X"11",X"AA",X"11",X"AA",X"11",X"AA",X"21",X"AA",X"A2",
		X"DD",X"DD",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"00",X"11",X"0D",X"11",X"D1",X"11",X"11",X"11",
		X"0D",X"11",X"D1",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"00",X"D1",X"00",X"11",
		X"00",X"0D",X"00",X"D1",X"00",X"11",X"DD",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"00",X"11",X"D0",X"11",X"1D",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"1D",X"00",X"11",X"00",X"11",X"DD",
		X"00",X"00",X"D0",X"00",X"1D",X"00",X"11",X"00",X"11",X"D0",X"11",X"1D",X"11",X"11",X"11",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"00",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"FF",X"FF",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"22",X"22",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"22",X"22",
		X"11",X"12",X"11",X"12",X"11",X"12",X"11",X"12",X"11",X"12",X"11",X"12",X"11",X"12",X"22",X"22",
		X"DD",X"DD",X"EE",X"EE",X"EE",X"EE",X"DD",X"AB",X"EE",X"AB",X"EE",X"FA",X"DD",X"CA",X"EE",X"AC",
		X"88",X"56",X"CC",X"56",X"CC",X"88",X"BA",X"88",X"BA",X"88",X"AC",X"CC",X"BC",X"CC",X"FF",X"FF",
		X"EE",X"AA",X"DD",X"AA",X"EE",X"AA",X"EE",X"AA",X"D5",X"A2",X"55",X"55",X"EC",X"EE",X"5C",X"EE",
		X"CC",X"CF",X"CB",X"CF",X"BF",X"FF",X"AE",X"EE",X"CC",X"CC",X"2C",X"FC",X"EE",X"FC",X"EE",X"CC",
		X"B2",X"B2",X"AA",X"AB",X"FA",X"FA",X"FA",X"FA",X"AA",X"AB",X"AC",X"BB",X"AA",X"AB",X"2B",X"44",
		X"55",X"52",X"29",X"82",X"99",X"98",X"99",X"99",X"F9",X"99",X"55",X"99",X"55",X"88",X"29",X"82",
		X"BB",X"44",X"CB",X"BC",X"BF",X"BB",X"BC",X"BB",X"BF",X"BB",X"FF",X"44",X"FF",X"BB",X"FF",X"BB",
		X"EE",X"E2",X"CE",X"E2",X"EE",X"E2",X"EE",X"EE",X"EE",X"EE",X"CE",X"EE",X"CE",X"EE",X"2E",X"E2",
		X"BF",X"BB",X"BF",X"44",X"CB",X"4B",X"CF",X"BB",X"FF",X"2E",X"FA",X"AE",X"FA",X"A2",X"EA",X"AA",
		X"EE",X"ED",X"EE",X"EC",X"EE",X"CC",X"EE",X"EE",X"EE",X"EE",X"AE",X"BB",X"AE",X"2B",X"BA",X"22",
		X"FF",X"FF",X"CC",X"CF",X"CA",X"AF",X"FF",X"AA",X"AA",X"AA",X"1A",X"BB",X"21",X"AA",X"22",X"AB",
		X"AA",X"22",X"AA",X"99",X"AB",X"99",X"A9",X"9F",X"BF",X"9C",X"AF",X"9F",X"A9",X"59",X"AA",X"99",
		X"21",X"21",X"21",X"22",X"FF",X"F1",X"22",X"2F",X"2B",X"2F",X"FF",X"F1",X"1F",X"12",X"F2",X"21",
		X"BB",X"22",X"BB",X"A2",X"2B",X"BA",X"B2",X"BA",X"2F",X"BA",X"BB",X"A2",X"FF",X"BA",X"FF",X"BA",
		X"CF",X"C1",X"CF",X"AC",X"CC",X"C1",X"FF",X"CB",X"F2",X"CB",X"CC",X"11",X"1C",X"BB",X"CC",X"11",
		X"EF",X"EA",X"EF",X"2E",X"EE",X"E1",X"2E",X"2E",X"EE",X"EE",X"EE",X"EE",X"EE",X"11",X"EE",X"EE",
		X"21",X"21",X"21",X"22",X"FF",X"21",X"22",X"2F",X"2B",X"BF",X"FF",X"FF",X"2F",X"22",X"C2",X"C1",
		X"BB",X"22",X"2B",X"A2",X"B2",X"BA",X"2F",X"BA",X"BA",X"BA",X"BB",X"A1",X"FF",X"BA",X"EF",X"EA",
		X"CF",X"AC",X"CC",X"C1",X"FF",X"CA",X"F2",X"CA",X"CC",X"C1",X"C2",X"1A",X"CC",X"A1",X"CC",X"11",
		X"EF",X"2E",X"EE",X"E2",X"2E",X"2E",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"11",X"EE",X"E1",
		X"DA",X"DA",X"FE",X"DA",X"EE",X"ED",X"2E",X"ED",X"E2",X"ED",X"E2",X"DD",X"EE",X"EE",X"EE",X"ED",
		X"35",X"4D",X"FF",X"54",X"F2",X"54",X"57",X"54",X"35",X"DD",X"55",X"4D",X"55",X"54",X"25",X"24",
		X"CC",X"BD",X"CC",X"CB",X"C1",X"CB",X"F1",X"11",X"F1",X"11",X"88",X"12",X"11",X"2B",X"11",X"11",
		X"25",X"24",X"FF",X"FD",X"FF",X"FF",X"2F",X"FF",X"AF",X"FF",X"F2",X"FD",X"2F",X"D2",X"2F",X"22",
		X"DA",X"DA",X"FE",X"DA",X"2E",X"ED",X"E2",X"ED",X"E2",X"ED",X"EE",X"DD",X"EE",X"EE",X"CC",X"BE",
		X"35",X"5D",X"FF",X"55",X"2F",X"55",X"57",X"55",X"35",X"DD",X"55",X"5D",X"55",X"55",X"22",X"25",
		X"CC",X"CB",X"1C",X"1B",X"FF",X"F1",X"F2",X"21",X"17",X"1C",X"11",X"1C",X"11",X"1D",X"BB",X"1B",
		X"22",X"2D",X"FF",X"FD",X"FF",X"FF",X"22",X"2F",X"2A",X"2F",X"FF",X"FD",X"2F",X"22",X"FF",X"2D",
		X"DD",X"DD",X"EE",X"EE",X"EE",X"EE",X"DD",X"DD",X"EE",X"AB",X"EE",X"AB",X"DD",X"FA",X"EE",X"CA",
		X"88",X"68",X"CC",X"58",X"AA",X"88",X"2A",X"88",X"B2",X"88",X"AC",X"CC",X"AC",X"FF",X"FC",X"CC",
		X"EE",X"AC",X"DD",X"AA",X"EE",X"AB",X"EE",X"AA",X"D5",X"AA",X"55",X"55",X"EC",X"EE",X"55",X"EE",
		X"FB",X"BC",X"FF",X"FF",X"BF",X"EF",X"CC",X"CC",X"FC",X"FC",X"2F",X"FF",X"EE",X"FC",X"EE",X"CC",
		X"AB",X"AB",X"AA",X"AB",X"FA",X"FA",X"CA",X"FA",X"AC",X"AB",X"2A",X"BB",X"AA",X"AB",X"2A",X"AB",
		X"BB",X"BB",X"B9",X"8B",X"99",X"98",X"F9",X"99",X"F9",X"99",X"55",X"99",X"99",X"88",X"29",X"82",
		X"2B",X"44",X"BB",X"B4",X"CB",X"BC",X"BF",X"BB",X"BC",X"BB",X"2F",X"44",X"FF",X"BB",X"FF",X"BB",
		X"EE",X"EE",X"EC",X"CE",X"EE",X"EE",X"EE",X"EE",X"CE",X"EE",X"EC",X"EE",X"EC",X"EE",X"2E",X"E2",
		X"F7",X"77",X"FF",X"27",X"22",X"72",X"22",X"77",X"81",X"77",X"98",X"77",X"98",X"1C",X"99",X"1C",
		X"1B",X"BB",X"71",X"BB",X"71",X"F2",X"7B",X"2F",X"BB",X"FF",X"BB",X"CF",X"B1",X"CC",X"CC",X"CF",
		X"9F",X"8C",X"92",X"8C",X"92",X"8C",X"29",X"8B",X"99",X"11",X"99",X"CC",X"99",X"8B",X"88",X"BB",
		X"CC",X"CC",X"CF",X"CC",X"C2",X"CC",X"CC",X"CA",X"CA",X"AA",X"CC",X"A1",X"CC",X"AA",X"CC",X"A2",
		X"BB",X"AA",X"BB",X"AA",X"AA",X"AE",X"BB",X"E1",X"2B",X"E1",X"B2",X"A1",X"BB",X"A1",X"BB",X"44",
		X"22",X"22",X"C2",X"C2",X"22",X"F2",X"FF",X"FF",X"FE",X"FF",X"12",X"EE",X"22",X"FF",X"2F",X"FF",
		X"B4",X"44",X"44",X"49",X"44",X"77",X"44",X"77",X"44",X"4C",X"44",X"CC",X"44",X"C4",X"11",X"44",
		X"FF",X"FF",X"4C",X"FC",X"4C",X"FC",X"4C",X"CC",X"CC",X"CC",X"CF",X"FF",X"CF",X"FF",X"C2",X"2F",
		X"55",X"CE",X"55",X"EC",X"15",X"EC",X"21",X"EE",X"22",X"EE",X"22",X"11",X"22",X"22",X"22",X"22",
		X"EE",X"C2",X"EE",X"C2",X"EE",X"CF",X"EC",X"FF",X"EE",X"CF",X"EE",X"BF",X"E2",X"FC",X"1C",X"CF",
		X"FF",X"FF",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"21",X"FF",X"22",X"FF",X"22",X"1F",X"22",X"21",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"BF",X"BB",X"CF",X"4B",X"CB",X"BB",X"CF",X"B4",X"FF",X"A4",X"FF",X"BA",X"FE",X"BA",X"EA",X"AA",
		X"EE",X"ED",X"EE",X"ED",X"EE",X"EC",X"EE",X"CC",X"EE",X"ED",X"AA",X"ED",X"BB",X"BB",X"BB",X"DB",
		X"FA",X"AF",X"CA",X"AC",X"CA",X"AA",X"FF",X"AA",X"FF",X"BA",X"1F",X"AB",X"21",X"AA",X"22",X"AA",
		X"AA",X"D2",X"AA",X"99",X"AB",X"99",X"A9",X"9F",X"BF",X"9F",X"BF",X"9C",X"A9",X"99",X"AA",X"55",
		X"BB",X"B4",X"BB",X"BB",X"BB",X"BC",X"FB",X"BB",X"CB",X"BB",X"B4",X"44",X"FB",X"BB",X"FF",X"BB",
		X"AA",X"B2",X"CC",X"B2",X"CC",X"CC",X"CF",X"CC",X"FF",X"FC",X"CF",X"CF",X"CF",X"CF",X"FC",X"CF",
		X"FF",X"CB",X"8F",X"B4",X"98",X"4C",X"99",X"42",X"FE",X"22",X"EC",X"2E",X"CC",X"EC",X"EE",X"EE",
		X"FF",X"FF",X"CF",X"EE",X"CF",X"FC",X"FF",X"CC",X"FF",X"FC",X"EF",X"CC",X"EF",X"CC",X"EA",X"C2",
		X"AA",X"88",X"AA",X"88",X"AA",X"88",X"2A",X"C8",X"2A",X"C8",X"22",X"BB",X"8F",X"BB",X"BB",X"BB",
		X"AA",X"AA",X"BB",X"AA",X"CC",X"BB",X"BA",X"CC",X"BA",X"AA",X"4B",X"AA",X"44",X"BB",X"44",X"CC",
		X"BB",X"BB",X"CB",X"CB",X"CB",X"CB",X"BF",X"BB",X"BF",X"BB",X"2C",X"BB",X"2F",X"FB",X"BF",X"FF",
		X"CC",X"AA",X"BB",X"AA",X"BB",X"4A",X"BB",X"4A",X"BB",X"42",X"B4",X"25",X"44",X"2C",X"44",X"55",
		X"BB",X"B4",X"BB",X"BB",X"FB",X"BC",X"CB",X"BB",X"4B",X"BB",X"F4",X"44",X"FF",X"BB",X"FF",X"CB",
		X"AA",X"B2",X"CC",X"B2",X"CC",X"CC",X"CF",X"CC",X"FF",X"FC",X"FC",X"FF",X"FB",X"FF",X"FF",X"FF",
		X"FF",X"BB",X"8F",X"BC",X"98",X"42",X"99",X"42",X"F9",X"2C",X"FE",X"2E",X"EC",X"2E",X"EC",X"EE",
		X"CF",X"FF",X"FF",X"EE",X"CF",X"FC",X"FF",X"CC",X"FF",X"FC",X"FF",X"CC",X"EF",X"CC",X"EB",X"C2",
		X"22",X"DD",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"CC",X"33",X"DC",X"33",X"1D",X"33",X"11",X"23",X"11",X"D3",X"11",X"1D",X"11",X"11",X"11",X"11",
		X"3C",X"CD",X"33",X"D1",X"23",X"11",X"DD",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"EE",X"EE",X"CE",X"CE",X"EC",X"EE",X"EC",X"EE",X"DE",X"EE",X"EE",X"DD",X"DE",X"EE",X"EE",X"EE",
		X"AB",X"A2",X"AB",X"AB",X"DA",X"AA",X"DA",X"AA",X"4F",X"AF",X"BF",X"AF",X"BF",X"AC",X"BA",X"AC",
		X"11",X"ED",X"22",X"EE",X"22",X"1D",X"22",X"21",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"BB",X"AA",X"2B",X"AA",X"BB",X"BB",X"BA",X"AA",X"BA",X"AA",X"1A",X"AA",X"21",X"AA",X"22",X"AA",
		X"2A",X"CA",X"BA",X"44",X"BB",X"44",X"AA",X"44",X"AA",X"BA",X"FA",X"BB",X"FA",X"AB",X"FA",X"AB",
		X"BB",X"45",X"BB",X"45",X"BB",X"25",X"CC",X"25",X"CC",X"2C",X"CC",X"FC",X"CF",X"FF",X"FF",X"FF",
		X"AA",X"BB",X"AA",X"BF",X"AB",X"2F",X"BB",X"2F",X"AA",X"2F",X"AA",X"22",X"AA",X"22",X"AC",X"2A",
		X"FF",X"FF",X"CC",X"CC",X"CC",X"CC",X"BC",X"BC",X"CF",X"CC",X"FC",X"FC",X"FF",X"FF",X"2F",X"FF",
		X"AA",X"88",X"AA",X"88",X"AA",X"88",X"AA",X"8C",X"AA",X"C8",X"28",X"BB",X"8F",X"BB",X"BB",X"BB",
		X"AA",X"AA",X"AA",X"AA",X"CC",X"AA",X"BA",X"CC",X"BA",X"AA",X"4B",X"AA",X"44",X"BB",X"44",X"AA",
		X"CC",X"CC",X"CB",X"CB",X"BF",X"BB",X"BF",X"BB",X"BC",X"BB",X"2B",X"BB",X"2F",X"FB",X"BF",X"FF",
		X"BB",X"AA",X"BC",X"AA",X"BB",X"4A",X"BB",X"4A",X"BB",X"45",X"B4",X"2C",X"44",X"2C",X"44",X"55",
		X"EE",X"EE",X"EE",X"EE",X"CC",X"EE",X"CC",X"EE",X"EE",X"ED",X"EE",X"DE",X"EE",X"EE",X"EE",X"EE",
		X"AB",X"A2",X"AB",X"BB",X"2A",X"AA",X"4A",X"AA",X"4F",X"AF",X"BF",X"AF",X"BF",X"AF",X"BF",X"AC",
		X"11",X"DD",X"22",X"EE",X"22",X"1E",X"22",X"21",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"4B",X"AA",X"A4",X"AA",X"AA",X"BB",X"BA",X"AA",X"BA",X"AA",X"1A",X"AA",X"21",X"AA",X"22",X"AA",
		X"AA",X"AF",X"AC",X"4A",X"BC",X"4A",X"AB",X"4A",X"AA",X"A2",X"FA",X"B2",X"FA",X"B2",X"AA",X"B2",
		X"BB",X"45",X"BB",X"45",X"CC",X"25",X"CC",X"25",X"CC",X"22",X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"B2",X"AA",X"2F",X"BB",X"2F",X"AB",X"2F",X"AB",X"2F",X"BB",X"22",X"BC",X"2A",X"AA",X"AB",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"BC",X"CF",X"CC",X"FC",X"FC",X"CF",X"FF",X"FF",X"FF",X"2F",X"FF",
		X"AC",X"B2",X"CA",X"CC",X"1A",X"CC",X"21",X"B2",X"22",X"22",X"22",X"12",X"22",X"21",X"22",X"22",
		X"CF",X"EE",X"CF",X"FF",X"CF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CF",X"FF",X"CC",X"FF",X"CC",X"FF",
		X"FF",X"FF",X"DD",X"DF",X"DD",X"DF",X"DD",X"DF",X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"11",X"CC",X"22",X"CC",X"22",X"1C",X"22",X"21",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"33",X"03",X"33",X"3F",X"33",X"F3",X"33",X"F3",X"33",X"F3",X"33",
		X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"33",X"00",X"33",X"00",X"33",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"2C",X"00",X"33",X"00",X"33",X"C0",X"33",X"2C",X"33",X"2C",X"33",X"22",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"32",X"33",X"32",X"33",X"32",X"33",X"32",X"33",X"32",X"33",X"32",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"2C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",X"00",X"3F",X"00",X"3F",
		X"00",X"00",X"03",X"33",X"33",X"33",X"F3",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"3F",X"00",X"3F",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"33",X"33",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"2C",X"00",X"32",X"00",X"32",X"00",X"33",X"00",X"33",X"C0",X"33",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"C0",X"33",X"2C",X"33",X"2C",X"33",X"2C",X"33",X"22",X"33",X"22",X"33",X"22",X"33",X"22",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"33",X"03",X"33",X"33",X"C3",X"3C",X"33",X"C0",X"33",X"00",X"33",X"00",X"33",X"00",X"C3",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"B3",X"00",X"B3",X"00",X"BB",X"00",X"CB",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"32",X"C3",X"32",X"0C",X"2C",X"00",X"20",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"32",X"33",X"32",X"33",X"32",X"33",X"32",
		X"22",X"00",X"22",X"00",X"C2",X"C0",X"CC",X"20",X"C0",X"C0",X"C0",X"00",X"C0",X"00",X"00",X"00",
		X"33",X"22",X"33",X"22",X"33",X"22",X"33",X"2B",X"33",X"BB",X"32",X"CC",X"22",X"00",X"CC",X"00",
		X"C0",X"00",X"B0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C3",X"33",X"0C",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"0B",X"33",X"BB",X"33",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"CB",X"33",X"0C",X"33",X"00",X"B3",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"32",X"33",X"32",X"C3",X"2C",X"0C",X"2C",X"00",X"C0",
		X"33",X"22",X"33",X"22",X"33",X"22",X"33",X"22",X"33",X"22",X"33",X"22",X"33",X"22",X"33",X"22",
		X"C0",X"00",X"C0",X"00",X"20",X"00",X"C2",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"2C",X"33",X"2C",X"32",X"BC",X"22",X"BB",X"22",X"BB",X"22",X"CC",X"CC",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"33",X"03",X"33",X"33",X"33",X"3F",X"33",X"FF",X"33",X"F3",X"33",X"F3",X"33",X"33",X"33",
		X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"03",X"33",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"2C",X"00",X"33",X"00",X"33",X"C0",X"33",X"2C",X"33",X"2C",X"33",X"22",X"33",X"32",X"33",X"32",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"32",X"33",X"32",X"33",X"32",X"33",X"32",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"2C",X"00",X"22",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"33",X"00",X"33",X"03",X"33",X"33",X"33",X"3F",X"33",X"3F",X"33",X"F3",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"33",
		X"F3",X"33",X"F3",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"32",X"00",X"33",X"C0",X"33",X"2C",X"33",X"22",X"33",X"32",X"33",X"32",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"2C",X"00",X"2C",X"00",X"2C",X"00",X"22",X"00",
		X"33",X"33",X"C3",X"C3",X"0C",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"C3",X"00",X"03",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"32",X"33",X"32",X"CC",X"2C",X"00",X"2C",X"00",X"C0",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"32",X"33",X"32",X"33",X"32",X"33",X"32",X"33",X"22",X"33",X"22",
		X"22",X"2C",X"22",X"C0",X"CC",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"33",X"22",X"33",X"2B",X"33",X"BB",X"22",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BC",X"00",X"BC",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C3",X"00",X"C3",X"00",X"C3",X"03",X"03",X"0C",X"03",X"00",X"03",X"00",X"03",X"00",X"0C",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"BB",X"00",X"CC",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"32",X"33",X"32",X"CC",X"2C",X"00",X"2C",X"00",X"CC",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"22",X"C0",X"C2",X"22",X"2C",X"CC",X"2C",X"00",X"2C",X"00",X"2C",X"00",X"BB",X"00",X"BB",X"00",
		X"33",X"32",X"33",X"32",X"33",X"22",X"33",X"2C",X"33",X"C0",X"32",X"00",X"2C",X"00",X"C0",X"00",
		X"BB",X"00",X"BC",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"03",X"33",X"3F",X"33",X"FF",X"33",
		X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"33",X"00",X"33",X"00",X"33",
		X"F3",X"33",X"F3",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2C",X"00",X"33",X"00",X"33",X"C0",X"33",X"2C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"22",X"33",X"22",X"33",X"22",X"33",X"32",X"33",X"32",X"33",X"32",X"33",X"32",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"C2",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"33",X"03",X"33",X"33",X"33",X"3F",X"33",X"F3",X"33",X"F3",X"33",
		X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"33",X"00",X"33",X"00",X"33",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"2C",X"00",X"33",X"00",X"33",X"C0",X"33",X"2C",X"33",X"2C",X"33",X"22",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"32",X"33",X"32",X"33",X"32",X"33",X"32",X"33",X"32",X"33",X"32",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"2C",X"C0",X"CC",X"C2",X"C0",X"22",X"00",
		X"00",X"C3",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"C3",X"00",X"B3",X"00",X"B3",X"00",X"CB",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"32",X"33",X"32",X"33",X"2C",X"F3",X"CF",X"CC",X"FF",X"00",X"CC",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"32",X"33",X"32",X"33",X"32",
		X"22",X"00",X"22",X"00",X"2C",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",
		X"33",X"22",X"33",X"22",X"33",X"22",X"33",X"22",X"22",X"FB",X"2F",X"CC",X"FC",X"00",X"C0",X"00",
		X"00",X"00",X"BC",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"33",X"00",X"33",X"03",X"33",X"33",X"C3",X"3C",X"33",X"C0",X"33",X"00",X"33",X"00",X"C3",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"B3",X"00",X"B3",X"00",X"BB",X"00",X"CB",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"32",X"C3",X"32",X"0C",X"2C",X"00",X"2C",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"32",X"33",X"32",X"33",X"32",X"33",X"32",
		X"22",X"00",X"22",X"00",X"2C",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",
		X"33",X"22",X"33",X"22",X"33",X"22",X"33",X"2B",X"33",X"BB",X"32",X"CC",X"22",X"00",X"CC",X"00",
		X"00",X"00",X"B0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"03",X"33",X"33",X"33",X"3F",X"33",X"FF",X"33",
		X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"33",X"00",X"33",X"00",X"33",
		X"F3",X"33",X"F3",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"2C",X"00",X"33",X"00",X"33",X"C0",X"33",X"2C",X"33",X"2C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"22",X"33",X"32",X"33",X"32",X"33",X"32",X"33",X"32",X"33",X"32",X"33",X"32",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"C2",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"33",X"3F",X"33",X"FF",X"33",X"FF",X"33",
		X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",
		X"F3",X"33",X"F3",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"32",X"00",X"33",X"00",X"33",X"C0",X"33",X"2C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"22",X"33",X"22",X"33",X"32",X"33",X"32",X"33",X"32",X"33",X"32",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"C2",X"00",X"22",X"00",
		X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"CC",X"03",X"33",X"03",X"33",X"0C",X"33",X"00",X"C3",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"B3",X"00",X"B3",X"00",X"BB",X"00",X"CB",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"32",X"C3",X"32",X"0C",X"2C",X"00",X"2C",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"32",X"33",X"32",X"33",X"32",X"33",X"32",
		X"22",X"00",X"22",X"00",X"2C",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",
		X"33",X"22",X"33",X"22",X"33",X"22",X"33",X"2B",X"33",X"BB",X"32",X"CC",X"22",X"00",X"CC",X"00",
		X"00",X"00",X"B0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"23",X"00",X"33",X"00",X"33",X"00",X"3C",X"00",X"C3",X"00",X"33",X"00",X"33",X"00",X"C3",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"0F",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"CB",X"00",X"0C",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"F3",X"33",X"CF",X"33",X"0C",X"33",X"00",X"CC",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"32",X"33",X"32",X"33",X"32",X"33",X"32",
		X"22",X"00",X"2C",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",
		X"33",X"22",X"33",X"22",X"33",X"22",X"33",X"22",X"33",X"2B",X"22",X"2C",X"C2",X"C0",X"2C",X"00",
		X"C0",X"00",X"B0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",
		X"00",X"00",X"00",X"33",X"33",X"33",X"3F",X"33",X"F3",X"33",X"33",X"33",X"33",X"33",X"3F",X"33",
		X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",
		X"FF",X"33",X"FF",X"33",X"FF",X"33",X"FF",X"33",X"FF",X"BB",X"FB",X"BB",X"FF",X"BB",X"33",X"CB",
		X"00",X"00",X"2C",X"00",X"32",X"C0",X"33",X"2C",X"33",X"22",X"33",X"22",X"33",X"32",X"3F",X"32",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"32",X"FF",X"F2",X"CC",X"F2",X"CC",X"F2",X"BF",X"F3",X"BB",X"F3",X"CC",X"33",X"CF",X"33",
		X"C0",X"00",X"C0",X"00",X"C0",X"00",X"2C",X"00",X"2C",X"00",X"2C",X"00",X"2C",X"00",X"2C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",
		X"00",X"00",X"00",X"33",X"33",X"33",X"3F",X"33",X"F3",X"33",X"33",X"33",X"33",X"33",X"FF",X"33",
		X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"33",X"33",X"33",X"33",
		X"FF",X"33",X"FC",X"FF",X"CC",X"FF",X"CF",X"FB",X"FF",X"BC",X"FB",X"CC",X"FF",X"CC",X"3F",X"CC",
		X"00",X"00",X"2C",X"00",X"32",X"C0",X"33",X"2C",X"33",X"22",X"33",X"22",X"33",X"32",X"3F",X"32",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"F2",X"FC",X"F2",X"CC",X"FF",X"FF",X"FF",X"BF",X"FF",X"CB",X"FF",X"CB",X"F3",X"BC",X"33",
		X"C0",X"00",X"C0",X"00",X"C0",X"00",X"2C",X"00",X"2C",X"00",X"2C",X"22",X"2C",X"2C",X"22",X"C0",
		X"00",X"33",X"00",X"33",X"03",X"23",X"33",X"C3",X"32",X"33",X"CC",X"33",X"00",X"33",X"00",X"C3",
		X"3F",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"0C",X"00",X"0B",X"00",X"BB",X"00",X"0C",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"FF",X"BB",X"FF",X"BB",X"CC",X"CC",X"00",X"00",X"00",
		X"FF",X"33",X"FF",X"33",X"FF",X"33",X"FF",X"F3",X"FF",X"F3",X"FF",X"F3",X"FF",X"F3",X"FF",X"F2",
		X"20",X"00",X"22",X"00",X"22",X"00",X"22",X"00",X"CC",X"20",X"C0",X"C0",X"C0",X"00",X"00",X"00",
		X"FF",X"F2",X"FF",X"22",X"FF",X"22",X"FF",X"BC",X"FF",X"BB",X"CC",X"BB",X"00",X"CC",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C3",X"33",X"0C",X"33",X"00",X"33",X"00",X"23",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"CB",
		X"FF",X"BB",X"FF",X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"CB",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"CF",X"FF",X"BC",X"FF",X"BC",X"FF",X"CF",X"FF",X"CC",X"22",X"00",X"22",X"00",X"CC",
		X"CF",X"33",X"FF",X"33",X"FF",X"F3",X"FF",X"F3",X"FF",X"F3",X"FF",X"F3",X"FF",X"F3",X"FF",X"FC",
		X"22",X"00",X"22",X"00",X"CC",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",
		X"FF",X"CB",X"FF",X"BB",X"FF",X"BB",X"FF",X"BB",X"FF",X"BB",X"22",X"CC",X"CC",X"00",X"00",X"00",
		X"C0",X"00",X"BC",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"03",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",X"00",X"33",X"00",X"33",X"30",X"33",X"33",X"33",
		X"3F",X"33",X"F3",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"00",X"33",X"C0",X"33",X"2C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"32",X"33",X"32",X"33",X"32",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"3C",X"C0",X"2C",X"C3",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"CB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"0F",X"FF",X"FF",X"FF",
		X"00",X"0C",X"00",X"00",X"00",X"03",X"00",X"33",X"00",X"33",X"30",X"33",X"33",X"3F",X"33",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"BB",X"3F",X"CC",X"FF",X"BB",X"FF",X"BB",X"FF",X"33",X"FF",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"FC",X"0B",X"FF",X"0B",X"FF",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"BC",X"00",X"BC",X"00",X"C0",X"00",X"00",X"00",
		X"FF",X"F3",X"FF",X"F3",X"FF",X"33",X"CF",X"33",X"BB",X"33",X"FF",X"F3",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"3C",X"C0",X"3C",X"2C",X"C0",X"22",X"C0",
		X"0C",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"B3",X"00",X"B3",X"00",X"C3",X"00",X"0C",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"32",X"C3",X"2C",X"0C",X"2C",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"32",X"33",X"32",X"33",X"32",X"33",X"22",X"33",X"22",X"33",X"22",
		X"22",X"00",X"CC",X"00",X"BC",X"00",X"BC",X"00",X"BC",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"33",X"2C",X"22",X"C0",X"22",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C3",X"3F",X"0C",X"3F",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"23",X"00",X"23",
		X"FF",X"33",X"FF",X"33",X"FF",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"C2",X"00",X"02",X"00",X"0C",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"22",X"32",X"C2",X"22",X"0C",X"22",X"00",X"CC",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"3F",X"F3",X"33",X"33",X"33",X"33",X"33",X"32",X"33",X"32",X"33",X"22",
		X"22",X"00",X"22",X"00",X"2C",X"00",X"2C",X"00",X"2C",X"00",X"2C",X"00",X"C0",X"00",X"C0",X"00",
		X"33",X"22",X"32",X"22",X"22",X"22",X"22",X"2C",X"22",X"C0",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0B",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"CC",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"03",X"00",X"03",X"00",X"3F",X"00",X"3F",X"00",X"33",X"00",X"33",X"03",X"33",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"FF",X"BC",X"FF",X"CC",X"FB",X"CC",
		X"00",X"00",X"00",X"0B",X"00",X"0B",X"F0",X"BB",X"FF",X"BB",X"FF",X"CB",X"FF",X"FC",X"FF",X"F3",
		X"00",X"00",X"B0",X"00",X"BB",X"00",X"BB",X"00",X"BC",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"F3",X"CB",X"F3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"2C",X"00",X"22",X"00",
		X"00",X"00",X"00",X"0B",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"CC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"03",X"00",X"03",X"00",X"3F",X"00",X"3F",X"00",X"33",X"33",X"33",X"33",X"33",X"C3",X"33",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"FF",X"BB",X"FF",X"CC",X"FF",X"CC",
		X"00",X"00",X"00",X"BB",X"F0",X"BB",X"FF",X"BB",X"FF",X"CB",X"FF",X"FC",X"FF",X"F3",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"F3",X"BF",X"FF",
		X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"22",X"2C",X"2C",X"22",X"C0",X"22",X"00",
		X"33",X"33",X"33",X"33",X"3C",X"33",X"C0",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",
		X"FF",X"CC",X"FF",X"BB",X"FF",X"FB",X"CF",X"FF",X"FF",X"33",X"FF",X"33",X"33",X"33",X"33",X"33",
		X"00",X"33",X"00",X"C3",X"00",X"03",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"23",X"33",X"C2",X"22",X"0C",X"22",X"00",X"CC",
		X"BB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CF",X"FF",X"CF",X"FF",X"FF",X"FF",X"F3",
		X"22",X"00",X"2C",X"20",X"22",X"2C",X"22",X"22",X"2C",X"C2",X"2C",X"0C",X"2C",X"00",X"C0",X"00",
		X"33",X"32",X"33",X"22",X"33",X"22",X"33",X"22",X"22",X"2C",X"22",X"C0",X"CC",X"00",X"00",X"00",
		X"C0",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"F0",X"00",
		X"0C",X"3F",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"3F",X"00",X"33",X"00",X"33",
		X"FF",X"BB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"FF",X"33",X"33",X"33",
		X"00",X"C3",X"00",X"03",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"23",X"33",X"C2",X"22",X"0C",X"22",X"00",X"CC",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"FF",X"33",X"33",X"33",X"33",X"33",X"33",X"32",
		X"22",X"00",X"22",X"00",X"22",X"00",X"2C",X"00",X"2C",X"00",X"2C",X"00",X"C0",X"00",X"C0",X"00",
		X"33",X"22",X"33",X"22",X"33",X"22",X"22",X"2C",X"22",X"C0",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"33",X"03",X"33",X"33",X"33",X"3F",X"33",X"FF",X"33",X"F3",X"33",
		X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"33",X"00",X"33",X"00",X"33",
		X"F3",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"3C",X"00",X"33",X"00",X"33",X"C0",X"33",X"2C",X"33",X"2C",X"33",X"32",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"32",X"33",X"32",X"33",X"32",X"33",X"32",X"33",X"32",X"33",X"32",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"2C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"33",X"03",X"33",X"33",X"33",X"3F",X"33",X"F3",X"33",X"F3",X"33",X"33",X"33",
		X"00",X"00",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"33",X"30",X"33",X"33",X"33",X"03",X"33",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"3C",X"00",X"33",X"00",X"33",X"C0",X"33",X"2C",X"33",X"2C",X"33",X"32",X"33",X"32",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"32",X"33",X"32",X"33",X"32",X"33",X"32",X"33",X"32",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"2C",X"22",X"C0",X"22",X"00",
		X"00",X"33",X"03",X"33",X"03",X"C3",X"33",X"33",X"3C",X"33",X"C0",X"33",X"00",X"33",X"00",X"C3",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"B3",X"00",X"B3",X"00",X"BB",X"00",X"CB",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"CC",X"32",X"00",X"C2",X"00",X"0C",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"32",X"33",X"32",X"33",X"32",X"33",X"22",
		X"22",X"00",X"22",X"00",X"C2",X"00",X"CC",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",
		X"33",X"22",X"33",X"22",X"33",X"22",X"32",X"2B",X"22",X"BB",X"22",X"CC",X"CC",X"00",X"00",X"00",
		X"C0",X"00",X"B0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"33",X"00",X"C3",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"C3",X"00",X"03",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"03",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"32",X"FF",X"32",X"CC",X"FF",X"00",X"CC",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"32",X"33",X"32",X"33",X"32",X"33",X"32",X"33",X"22",
		X"2C",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"33",X"22",X"33",X"22",X"32",X"EB",X"2E",X"BB",X"FF",X"BB",X"CC",X"CC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"00",X"BC",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
