library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity snd1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of snd1 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"55",X"04",X"52",X"C5",X"A5",X"8A",X"40",X"8A",X"80",X"B9",X"02",X"BA",X"40",X"BB",X"40",X"FA",
		X"77",X"77",X"53",X"3F",X"6A",X"AA",X"AB",X"34",X"00",X"FB",X"97",X"67",X"6B",X"AB",X"34",X"00",
		X"E9",X"0F",X"FA",X"47",X"00",X"53",X"0F",X"37",X"17",X"6A",X"07",X"AA",X"AB",X"03",X"D8",X"E6",
		X"3C",X"34",X"00",X"FB",X"97",X"67",X"6B",X"AB",X"34",X"00",X"04",X"22",X"D5",X"23",X"2B",X"34",
		X"81",X"14",X"45",X"04",X"52",X"80",X"37",X"B4",X"33",X"C6",X"51",X"53",X"F0",X"96",X"51",X"04",
		X"45",X"83",X"05",X"85",X"A5",X"B8",X"20",X"B0",X"00",X"D5",X"27",X"AE",X"AF",X"C5",X"8A",X"80",
		X"14",X"73",X"26",X"74",X"A5",X"0A",X"37",X"B2",X"A8",X"27",X"AE",X"AF",X"A9",X"B4",X"35",X"14",
		X"73",X"04",X"62",X"93",X"B8",X"20",X"F0",X"03",X"05",X"C6",X"69",X"F0",X"03",X"09",X"C6",X"69",
		X"B8",X"08",X"A5",X"B5",X"D4",X"1A",X"D4",X"38",X"8A",X"80",X"C6",X"62",X"B9",X"03",X"34",X"3F",
		X"B4",X"35",X"E9",X"8E",X"B9",X"04",X"B4",X"35",X"E9",X"96",X"FA",X"03",X"F9",X"A9",X"C6",X"86",
		X"9A",X"7F",X"B4",X"35",X"E9",X"A2",X"04",X"86",X"BB",X"20",X"34",X"15",X"FB",X"77",X"77",X"53",
		X"3F",X"6B",X"AB",X"26",X"74",X"E6",X"AA",X"34",X"15",X"FB",X"77",X"77",X"53",X"3F",X"6B",X"AB",
		X"26",X"74",X"E6",X"B7",X"04",X"62",X"BA",X"08",X"B9",X"FF",X"8A",X"80",X"A5",X"B5",X"FA",X"AB",
		X"34",X"31",X"34",X"31",X"FA",X"97",X"67",X"6A",X"F6",X"62",X"AB",X"34",X"31",X"34",X"31",X"34",
		X"31",X"FA",X"AB",X"34",X"31",X"34",X"31",X"FA",X"97",X"67",X"97",X"67",X"6A",X"AA",X"04",X"CE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"B8",X"03",X"34",X"23",X"E8",X"02",X"B8",X"03",X"34",X"0D",X"E8",X"08",X"83",X"27",X"AE",X"AF",
		X"D5",X"AE",X"AF",X"C4",X"7B",X"FB",X"47",X"E7",X"53",X"1F",X"AF",X"FB",X"47",X"E7",X"53",X"E0",
		X"AE",X"A4",X"35",X"FB",X"77",X"77",X"AE",X"53",X"3F",X"AF",X"FE",X"53",X"C0",X"AE",X"D5",X"C4",
		X"7B",X"FB",X"77",X"77",X"AE",X"53",X"3F",X"AF",X"FE",X"53",X"C0",X"AE",X"D5",X"A4",X"35",X"FE",
		X"6F",X"E6",X"44",X"1F",X"6F",X"E6",X"48",X"1F",X"AE",X"83",X"AB",X"D5",X"FB",X"1B",X"C5",X"B4",
		X"33",X"C6",X"9E",X"F2",X"9F",X"A8",X"D4",X"1A",X"D4",X"38",X"D4",X"4B",X"C6",X"4B",X"B9",X"03",
		X"8A",X"80",X"34",X"3F",X"D5",X"34",X"3F",X"D4",X"7B",X"E9",X"62",X"B9",X"04",X"D5",X"D4",X"7B",
		X"E9",X"6D",X"FA",X"03",X"F9",X"A9",X"C6",X"58",X"9A",X"7F",X"D5",X"D4",X"7B",X"E9",X"7A",X"24",
		X"58",X"AB",X"D5",X"FB",X"1B",X"C5",X"B4",X"33",X"C6",X"9E",X"F2",X"9F",X"A8",X"D4",X"1A",X"D4",
		X"38",X"D4",X"4B",X"C6",X"82",X"FA",X"A9",X"D5",X"D4",X"7B",X"E9",X"97",X"24",X"8F",X"83",X"BE",
		X"80",X"A4",X"A2",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"03",X"06",X"09",X"0C",X"0F",X"12",X"15",X"18",X"1B",X"1E",X"21",X"24",X"27",X"2A",X"2D",
		X"30",X"33",X"36",X"39",X"3C",X"3F",X"42",X"45",X"48",X"4B",X"4E",X"51",X"54",X"57",X"5A",X"5D",
		X"60",X"5D",X"5A",X"57",X"54",X"51",X"4E",X"4B",X"48",X"45",X"42",X"3F",X"3C",X"39",X"36",X"33",
		X"30",X"2D",X"2A",X"27",X"24",X"21",X"1E",X"1B",X"18",X"15",X"12",X"0F",X"0C",X"09",X"06",X"03",
		X"FC",X"6E",X"AC",X"FD",X"7F",X"AD",X"77",X"77",X"53",X"3F",X"A3",X"A8",X"C5",X"FC",X"6E",X"AC",
		X"FD",X"7F",X"AD",X"77",X"77",X"43",X"C0",X"A3",X"D5",X"68",X"39",X"16",X"5F",X"44",X"40",X"C5",
		X"83",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"05",X"0A",X"0F",X"14",X"19",X"1E",X"23",X"28",X"2D",X"32",X"37",X"3C",X"41",X"46",X"4B",
		X"50",X"55",X"5A",X"5F",X"64",X"69",X"6E",X"73",X"78",X"7D",X"82",X"87",X"8C",X"91",X"96",X"9B",
		X"9F",X"9B",X"96",X"91",X"8C",X"87",X"82",X"7D",X"78",X"73",X"6E",X"69",X"64",X"5F",X"5A",X"55",
		X"50",X"4B",X"46",X"41",X"3C",X"37",X"32",X"2D",X"28",X"23",X"1E",X"19",X"14",X"0F",X"0A",X"05",
		X"00",X"2A",X"80",X"1C",X"84",X"0E",X"88",X"8A",X"88",X"00",X"16",X"84",X"0B",X"84",X"84",X"00",
		X"00",X"18",X"84",X"0C",X"80",X"80",X"00",X"10",X"B8",X"B4",X"B0",X"00",X"12",X"90",X"09",X"90",
		X"90",X"12",X"90",X"90",X"94",X"90",X"94",X"90",X"94",X"09",X"94",X"94",X"12",X"94",X"94",X"98",
		X"94",X"98",X"94",X"00",X"00",X"09",X"B0",X"B2",X"B4",X"12",X"BA",X"B6",X"00",X"0E",X"A4",X"1C",
		X"E8",X"90",X"D8",X"88",X"38",X"E0",X"80",X"00",X"60",X"CA",X"82",X"20",X"CC",X"84",X"40",X"D0",
		X"86",X"CA",X"82",X"08",X"DA",X"89",X"D9",X"89",X"DA",X"89",X"D9",X"89",X"DA",X"89",X"D9",X"89",
		X"DA",X"89",X"D9",X"89",X"08",X"DA",X"89",X"D9",X"89",X"DA",X"89",X"D9",X"89",X"DA",X"89",X"D9",
		X"89",X"DA",X"89",X"D9",X"89",X"7F",X"DA",X"8A",X"00",X"00",X"24",X"88",X"82",X"88",X"82",X"12",
		X"D8",X"88",X"D6",X"88",X"D8",X"82",X"D6",X"82",X"D6",X"88",X"88",X"D6",X"82",X"82",X"24",X"DA",
		X"87",X"D9",X"83",X"DA",X"87",X"D7",X"83",X"09",X"D8",X"88",X"D7",X"88",X"D8",X"88",X"D7",X"88",
		X"D8",X"82",X"D7",X"82",X"D8",X"82",X"D7",X"82",X"48",X"D8",X"88",X"00",X"00",X"00",X"20",X"E8",
		X"88",X"82",X"E2",X"88",X"10",X"82",X"A4",X"20",X"DC",X"88",X"82",X"84",X"18",X"E0",X"87",X"08",
		X"A2",X"20",X"E4",X"88",X"E7",X"82",X"E8",X"88",X"EA",X"82",X"20",X"EA",X"88",X"EC",X"82",X"88",
		X"82",X"EC",X"88",X"82",X"F0",X"90",X"88",X"EC",X"88",X"82",X"10",X"84",X"AA",X"E8",X"8C",X"AA",
		X"20",X"E7",X"92",X"8A",X"10",X"84",X"A4",X"E2",X"8C",X"A4",X"00",X"1B",X"E2",X"88",X"09",X"A4",
		X"12",X"82",X"A8",X"12",X"88",X"A4",X"E2",X"82",X"A4",X"12",X"E0",X"80",X"09",X"82",X"83",X"86",
		X"88",X"8A",X"8C",X"24",X"D0",X"88",X"00",X"20",X"80",X"DC",X"98",X"E0",X"9A",X"E2",X"9C",X"20",
		X"90",X"E4",X"88",X"10",X"E3",X"90",X"A4",X"20",X"88",X"DA",X"8A",X"EA",X"84",X"10",X"E8",X"8A",
		X"A4",X"20",X"84",X"E2",X"82",X"E2",X"87",X"16",X"E8",X"88",X"0A",X"A3",X"10",X"E4",X"82",X"A0",
		X"15",X"C8",X"80",X"2B",X"CA",X"83",X"40",X"CB",X"80",X"00",X"10",X"E8",X"A4",X"E8",X"A4",X"E6",
		X"A2",X"E6",X"A2",X"E4",X"A0",X"E4",X"A0",X"E2",X"9C",X"E2",X"9C",X"10",X"E0",X"90",X"A0",X"E4",
		X"88",X"A0",X"E4",X"80",X"A0",X"E4",X"88",X"A8",X"20",X"EA",X"96",X"E8",X"90",X"40",X"F0",X"80",
		X"00",X"10",X"E8",X"A4",X"E8",X"A4",X"E6",X"A2",X"E6",X"A2",X"E4",X"A0",X"E4",X"A0",X"E2",X"9C",
		X"E2",X"9C",X"20",X"E0",X"90",X"10",X"88",X"08",X"A0",X"A2",X"20",X"E4",X"90",X"E0",X"88",X"20",
		X"E2",X"92",X"10",X"8A",X"08",X"A2",X"A4",X"20",X"E6",X"92",X"E2",X"8A",X"20",X"E8",X"88",X"10",
		X"82",X"A8",X"EA",X"88",X"A8",X"E6",X"82",X"A4",X"E8",X"80",X"2B",X"83",X"40",X"80",X"00",X"0A",
		X"E8",X"A4",X"EA",X"A6",X"14",X"EC",X"A8",X"28",X"E8",X"A4",X"0A",X"E8",X"A4",X"EA",X"A6",X"14",
		X"EC",X"A8",X"28",X"E8",X"A4",X"00",X"0A",X"E0",X"98",X"E0",X"98",X"3C",X"E0",X"98",X"12",X"88",
		X"84",X"88",X"84",X"88",X"84",X"88",X"84",X"88",X"84",X"88",X"84",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"A3",X"83",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"20",X"10",X"05",X"06",X"12",X"40",X"16",X"01",X"02",X"00",X"04",X"14",X"FA",X"1E",X"2D",
		X"10",X"00",X"13",X"00",X"11",X"00",X"14",X"83",X"FE",X"85",X"FE",X"85",X"FE",X"00",X"15",X"00",
		X"0A",X"00",X"95",X"FE",X"85",X"FE",X"85",X"FE",X"00",X"00",X"00",X"09",X"00",X"FE",X"84",X"FE",
		X"83",X"FE",X"00",X"A3",X"83",X"D5",X"B8",X"20",X"80",X"37",X"53",X"0F",X"20",X"37",X"17",X"60",
		X"96",X"64",X"B6",X"BD",X"46",X"BA",X"F0",X"A3",X"C6",X"5D",X"F2",X"5F",X"34",X"3F",X"E9",X"5D",
		X"FF",X"96",X"56",X"FE",X"C6",X"75",X"FA",X"03",X"F8",X"A9",X"27",X"AE",X"AF",X"C4",X"7B",X"27",
		X"AE",X"AF",X"C4",X"7B",X"F0",X"A3",X"C6",X"5F",X"F2",X"8C",X"92",X"7D",X"B2",X"81",X"D2",X"E5",
		X"8A",X"80",X"A8",X"D4",X"1A",X"D4",X"38",X"C6",X"64",X"B9",X"08",X"C4",X"7B",X"34",X"4A",X"04",
		X"52",X"34",X"81",X"04",X"52",X"C5",X"BE",X"80",X"F4",X"06",X"04",X"52",X"76",X"91",X"C5",X"04",
		X"74",X"B0",X"08",X"A4",X"46",X"D5",X"FB",X"1B",X"C5",X"A3",X"C6",X"9E",X"96",X"A2",X"14",X"45",
		X"04",X"52",X"D2",X"B6",X"97",X"F7",X"97",X"F7",X"A9",X"23",X"80",X"62",X"16",X"AE",X"16",X"B2",
		X"A4",X"AE",X"E9",X"A9",X"A4",X"95",X"F4",X"06",X"A4",X"95",X"95",X"BB",X"F0",X"FB",X"E7",X"E7",
		X"47",X"53",X"03",X"96",X"C6",X"17",X"37",X"17",X"6B",X"AB",X"03",X"E0",X"F6",X"D7",X"85",X"27",
		X"AE",X"AF",X"B8",X"20",X"A0",X"C4",X"7B",X"FB",X"47",X"E7",X"53",X"1F",X"AF",X"FB",X"47",X"E7",
		X"53",X"E0",X"AE",X"C4",X"7B",X"B0",X"04",X"C5",X"F9",X"F2",X"ED",X"04",X"C6",X"D5",X"A4",X"46",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"28",X"00",X"2A",X"61",X"2C",X"E6",X"2F",X"91",X"32",X"66",X"FF",X"FF",X"35",X"65",X"38",X"92",
		X"3B",X"EF",X"3F",X"75",X"43",X"46",X"47",X"46",X"4B",X"83",X"BB",X"00",X"B9",X"30",X"B1",X"FF",
		X"D4",X"27",X"96",X"20",X"E8",X"20",X"83",X"B9",X"30",X"FB",X"96",X"2D",X"11",X"F1",X"96",X"34",
		X"FB",X"1B",X"E3",X"83",X"FB",X"1B",X"84",X"F8",X"D4",X"27",X"C6",X"5C",X"F2",X"46",X"AA",X"D4",
		X"27",X"F2",X"46",X"A9",X"D4",X"27",X"A8",X"D4",X"5D",X"F8",X"83",X"D2",X"54",X"D5",X"BE",X"00",
		X"BF",X"00",X"C5",X"83",X"D4",X"27",X"D5",X"A8",X"D4",X"5D",X"C5",X"F8",X"83",X"F8",X"53",X"0F",
		X"E7",X"AC",X"A3",X"AF",X"FC",X"17",X"A3",X"AE",X"F8",X"53",X"30",X"47",X"AC",X"FF",X"97",X"67",
		X"AF",X"FE",X"67",X"AE",X"1C",X"FC",X"03",X"FC",X"96",X"6D",X"83",X"42",X"03",X"80",X"62",X"76",
		X"A2",X"FC",X"6E",X"AC",X"FD",X"7F",X"AD",X"77",X"77",X"43",X"C0",X"A3",X"A8",X"C5",X"FC",X"6E",
		X"AC",X"FD",X"7F",X"AD",X"77",X"77",X"43",X"C0",X"A3",X"D5",X"68",X"39",X"16",X"A0",X"C4",X"81",
		X"C5",X"83",X"44",X"40",X"A3",X"83",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"03",X"06",X"09",X"0C",X"0F",X"12",X"15",X"18",X"1B",X"1E",X"21",X"24",X"27",X"2A",X"2D",
		X"30",X"33",X"36",X"39",X"3C",X"3F",X"42",X"45",X"48",X"4B",X"4E",X"51",X"54",X"57",X"5A",X"5D",
		X"60",X"5D",X"5A",X"57",X"54",X"51",X"4E",X"4B",X"48",X"45",X"42",X"3F",X"3C",X"39",X"36",X"33",
		X"30",X"2D",X"2A",X"27",X"24",X"21",X"1E",X"1B",X"18",X"15",X"12",X"0F",X"0C",X"09",X"06",X"03",
		X"02",X"04",X"06",X"0C",X"14",X"FF",X"A8",X"A3",X"28",X"17",X"A3",X"A9",X"12",X"24",X"C9",X"F4",
		X"24",X"9A",X"7F",X"B8",X"00",X"B9",X"FF",X"F4",X"24",X"9A",X"7F",X"B8",X"00",X"B9",X"FF",X"F4",
		X"24",X"8A",X"80",X"83",X"BF",X"00",X"9A",X"BF",X"A5",X"23",X"B0",X"48",X"3A",X"BA",X"08",X"81",
		X"E9",X"3B",X"AB",X"C8",X"F8",X"F2",X"BA",X"43",X"B0",X"3A",X"FB",X"77",X"AB",X"F2",X"78",X"76",
		X"5B",X"1F",X"FF",X"A3",X"F2",X"4A",X"37",X"17",X"E4",X"4E",X"CF",X"00",X"23",X"EC",X"6E",X"AE",
		X"F6",X"59",X"27",X"AE",X"39",X"EA",X"AC",X"E4",X"2D",X"E4",X"54",X"A5",X"CF",X"FF",X"F2",X"62",
		X"E4",X"64",X"27",X"AF",X"A3",X"37",X"17",X"6E",X"F6",X"71",X"27",X"AE",X"39",X"EA",X"AC",X"E4",
		X"2D",X"00",X"AE",X"39",X"EA",X"AC",X"E4",X"2D",X"76",X"93",X"B5",X"CF",X"FF",X"F2",X"81",X"E4",
		X"83",X"27",X"AF",X"A3",X"6E",X"AE",X"E6",X"90",X"23",X"FF",X"AE",X"39",X"EA",X"AC",X"E4",X"2D",
		X"00",X"E4",X"8B",X"1F",X"FF",X"A3",X"F2",X"9C",X"00",X"00",X"E4",X"9F",X"CF",X"FF",X"A3",X"6E",
		X"E6",X"AA",X"23",X"FF",X"AE",X"39",X"EA",X"AC",X"E4",X"2D",X"E4",X"A4",X"FB",X"C6",X"B4",X"00",
		X"00",X"00",X"E4",X"3B",X"81",X"C6",X"BA",X"FB",X"E4",X"3B",X"8A",X"40",X"A5",X"83",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"FF",X"05",X"FF",X"02",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
