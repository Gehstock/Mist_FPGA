library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ckong_big_sprite_tile_bit0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ckong_big_sprite_tile_bit0 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"1E",X"3F",X"3F",X"3F",X"7D",X"7F",X"3E",X"CC",X"E6",X"EF",X"C3",X"E7",X"E7",X"E7",X"C3",
		X"1E",X"3F",X"7D",X"3F",X"1F",X"0C",X"00",X"0F",X"F7",X"F7",X"E7",X"C3",X"E7",X"F6",X"E6",X"FC",
		X"00",X"1E",X"3F",X"3F",X"3F",X"6F",X"7F",X"3E",X"CC",X"E6",X"EF",X"C3",X"E7",X"E7",X"E7",X"C3",
		X"1E",X"3F",X"7F",X"3F",X"1B",X"0C",X"00",X"0F",X"F7",X"F7",X"E7",X"C3",X"E7",X"F6",X"E6",X"FC",
		X"00",X"1E",X"3B",X"3F",X"3F",X"7F",X"7F",X"3E",X"CC",X"E6",X"EF",X"C3",X"E7",X"E7",X"E7",X"C3",
		X"1E",X"3F",X"77",X"3F",X"1F",X"0C",X"00",X"0F",X"F7",X"F7",X"E7",X"C3",X"E7",X"F6",X"E6",X"FC",
		X"0F",X"01",X"09",X"1F",X"3F",X"3F",X"1A",X"0E",X"E0",X"D8",X"B8",X"BC",X"BC",X"BC",X"BC",X"BC",
		X"1A",X"3F",X"3F",X"1F",X"09",X"01",X"01",X"0F",X"BC",X"BC",X"BC",X"BC",X"B8",X"D8",X"E0",X"E0",
		X"0F",X"01",X"09",X"1F",X"3F",X"3F",X"1A",X"0E",X"D0",X"F8",X"D8",X"8C",X"DC",X"FC",X"DC",X"8C",
		X"1A",X"3F",X"3F",X"1F",X"09",X"01",X"01",X"0F",X"DC",X"FC",X"DC",X"8C",X"D8",X"F8",X"D8",X"F0",
		X"38",X"FC",X"FF",X"EF",X"FF",X"FF",X"FF",X"7F",X"00",X"00",X"40",X"80",X"80",X"C0",X"00",X"80",
		X"7F",X"FF",X"FF",X"FF",X"EF",X"FF",X"FC",X"38",X"C0",X"80",X"C0",X"80",X"80",X"40",X"00",X"00",
		X"00",X"00",X"09",X"00",X"00",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"04",
		X"08",X"04",X"04",X"03",X"00",X"00",X"00",X"00",X"04",X"08",X"0C",X"0C",X"14",X"1C",X"1C",X"0C",
		X"00",X"00",X"00",X"00",X"01",X"02",X"04",X"08",X"01",X"03",X"07",X"E3",X"07",X"05",X"03",X"03",
		X"00",X"00",X"48",X"B4",X"00",X"00",X"00",X"00",X"03",X"07",X"05",X"03",X"06",X"00",X"00",X"00",
		X"00",X"00",X"38",X"3C",X"7C",X"7F",X"FF",X"FC",X"00",X"00",X"00",X"00",X"40",X"80",X"00",X"00",
		X"FC",X"FC",X"78",X"20",X"00",X"00",X"06",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"EE",X"60",X"00",X"0E",X"1A",X"1D",X"18",X"00",X"10",X"30",X"30",
		X"10",X"08",X"08",X"04",X"02",X"02",X"01",X"00",X"60",X"40",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"3C",X"60",X"C0",
		X"01",X"03",X"06",X"04",X"04",X"01",X"06",X"0E",X"80",X"00",X"00",X"00",X"00",X"01",X"03",X"E0",
		X"00",X"00",X"00",X"00",X"C0",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"17",X"E7",X"87",X"06",X"06",X"00",X"40",X"E0",X"70",X"B0",X"F8",X"18",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"78",X"FE",X"33",
		X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"40",X"07",X"81",X"83",X"03",X"03",X"01",X"00",X"00",
		X"0F",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"03",X"03",X"05",X"07",X"07",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0E",X"5E",X"FF",X"FF",X"CF",X"C6",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"E0",X"E0",
		X"01",X"01",X"03",X"03",X"87",X"C7",X"7F",X"3F",X"E0",X"E0",X"C0",X"C1",X"83",X"87",X"07",X"03",
		X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"04",X"00",X"01",X"07",X"3C",X"C0",X"00",X"00",X"00",
		X"04",X"08",X"09",X"09",X"08",X"10",X"10",X"10",X"00",X"00",X"FC",X"07",X"01",X"00",X"00",X"00",
		X"03",X"07",X"07",X"03",X"08",X"1C",X"1E",X"3F",X"00",X"00",X"C0",X"60",X"30",X"1C",X"3E",X"7E",
		X"3F",X"3B",X"1F",X"03",X"03",X"03",X"01",X"00",X"F6",X"EE",X"DC",X"DC",X"DC",X"D8",X"D0",X"60",
		X"00",X"00",X"01",X"01",X"02",X"02",X"02",X"04",X"40",X"80",X"00",X"00",X"00",X"42",X"33",X"07",
		X"04",X"04",X"08",X"08",X"08",X"08",X"08",X"08",X"07",X"07",X"07",X"07",X"00",X"00",X"00",X"00",
		X"00",X"80",X"C0",X"40",X"61",X"3A",X"0E",X"07",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"0A",X"32",X"41",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",
		X"60",X"F0",X"A0",X"80",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"60",X"20",X"20",
		X"00",X"08",X"08",X"04",X"0E",X"08",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"0C",X"06",X"06",X"06",X"04",X"08",X"10",X"00",X"00",X"0C",X"0E",X"0F",X"0F",X"0F",X"07",
		X"20",X"00",X"80",X"60",X"18",X"0C",X"00",X"00",X"07",X"03",X"03",X"01",X"00",X"00",X"00",X"00",
		X"00",X"18",X"20",X"40",X"80",X"00",X"00",X"21",X"00",X"00",X"10",X"70",X"70",X"F0",X"F0",X"F0",
		X"11",X"09",X"04",X"04",X"06",X"06",X"06",X"06",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"01",X"03",X"06",X"0C",X"15",X"00",X"00",X"80",X"40",X"E0",X"30",X"18",X"54",
		X"15",X"0C",X"06",X"03",X"01",X"00",X"00",X"00",X"54",X"18",X"30",X"E0",X"40",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"20",X"50",X"70",X"50",X"D8",X"88",X"88",X"04",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"88",X"88",X"D8",X"50",X"70",X"50",X"20",
		X"00",X"44",X"02",X"01",X"05",X"43",X"0F",X"16",X"00",X"00",X"00",X"78",X"FE",X"86",X"03",X"73",
		X"03",X"0E",X"5B",X"21",X"00",X"00",X"00",X"00",X"7B",X"3B",X"33",X"86",X"FE",X"3C",X"00",X"00",
		X"00",X"00",X"28",X"87",X"33",X"1E",X"0C",X"44",X"00",X"80",X"78",X"FC",X"86",X"03",X"71",X"F9",
		X"32",X"1E",X"0D",X"03",X"01",X"00",X"00",X"00",X"F9",X"79",X"7B",X"32",X"86",X"FC",X"38",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"19",X"3C",X"7F",X"00",X"00",X"00",X"00",X"04",X"08",X"10",X"50",
		X"EF",X"F2",X"DC",X"6C",X"30",X"18",X"03",X"07",X"E0",X"00",X"00",X"00",X"00",X"00",X"CC",X"9E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"08",X"10",X"20",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"05",X"07",X"87",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"07",X"03",X"07",X"05",X"03",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"07",X"07",X"1F",X"1F",X"0C",X"07",X"3A",X"3B",X"FB",X"C1",X"FB",X"FB",X"E1",X"BB",
		X"07",X"0C",X"1F",X"1F",X"07",X"07",X"03",X"00",X"BB",X"E1",X"FB",X"FB",X"C1",X"FB",X"3B",X"3A",
		X"0F",X"0C",X"1F",X"1F",X"1F",X"1B",X"0F",X"80",X"C0",X"60",X"70",X"8C",X"E7",X"E8",X"EA",X"0A",
		X"83",X"87",X"0F",X"1F",X"1F",X"1F",X"1F",X"0C",X"1C",X"1C",X"DE",X"CE",X"E8",X"E9",X"5F",X"26",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"80",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"9E",X"CC",X"80",X"20",X"10",X"08",X"04",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"01",X"00",X"00",X"00",X"00",X"00",
		X"08",X"18",X"30",X"30",X"20",X"40",X"40",X"80",X"5C",X"B0",X"C0",X"00",X"C0",X"40",X"40",X"40",
		X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"40",X"40",X"20",X"38",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"0C",X"0C",X"0C",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"18",X"3C",X"3C",X"2C",X"2C",X"3C",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
