library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity prom_palette_ic41 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(6 downto 0);
	data : out std_logic_vector(2 downto 0)
);
end entity;

architecture prom of prom_palette_ic41 is
	type rom is array(0 to  127) of std_logic_vector(2 downto 0);
	signal rom_data: rom := (
		"000","000","000","000","000","000","000","000","010","110","101","011","101","110","110","110",
		"001","011","011","110","010","011","011","011","111","101","101","011","111","101","101","101",
		"000","000","000","000","000","000","000","000","110","001","001","011","011","011","001","100",
		"110","101","101","111","111","111","111","011","110","111","111","101","101","101","011","111",
		"000","000","000","000","000","000","000","000","010","010","101","011","011","011","011","011",
		"001","011","011","110","110","110","110","110","101","101","101","011","101","101","101","101",
		"000","000","000","000","000","000","000","000","110","001","001","100","100","100","011","100",
		"110","101","101","101","101","101","111","011","101","111","111","111","111","111","101","111");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
