library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity exerion_01 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of exerion_01 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"48",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"84",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"68",X"00",X"00",X"CC",X"33",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"C3",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"CC",X"77",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"0C",X"F0",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"78",X"00",X"00",X"EE",X"77",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"0F",X"0F",X"07",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"C3",X"F0",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"78",X"00",X"00",X"EE",X"FF",X"00",X"00",X"00",X"00",
		X"08",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"E1",X"00",X"00",X"00",X"00",X"0C",X"F0",X"F0",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"F0",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"0C",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"87",X"00",X"00",X"00",X"0C",X"C3",X"F0",X"F0",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"78",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"3C",X"0F",X"00",X"00",X"08",X"C3",X"F0",X"F0",X"F0",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"80",X"F0",X"78",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"0E",X"0F",X"0F",X"8F",X"FF",X"1F",X"E1",X"0F",X"00",X"08",X"87",X"F0",X"F0",X"F0",X"F0",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"F0",X"F0",X"00",X"88",X"FF",X"B3",X"00",X"00",X"00",X"00",
		X"0F",X"FF",X"87",X"EF",X"FF",X"7F",X"C3",X"1E",X"00",X"00",X"86",X"F0",X"F0",X"F0",X"F0",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"F0",X"F8",X"00",X"88",X"FF",X"D9",X"30",X"00",X"00",X"00",
		X"CF",X"FF",X"97",X"EF",X"FF",X"FF",X"87",X"3C",X"00",X"00",X"08",X"69",X"F0",X"F0",X"F0",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"FF",X"00",X"88",X"FF",X"EC",X"73",X"00",X"00",X"00",
		X"CF",X"FF",X"B7",X"FF",X"FF",X"FF",X"97",X"F0",X"00",X"00",X"00",X"86",X"F0",X"F0",X"F0",X"FC",
		X"00",X"00",X"00",X"00",X"80",X"F0",X"FE",X"FF",X"00",X"88",X"7F",X"CF",X"F7",X"00",X"00",X"00",
		X"EF",X"FF",X"F7",X"FE",X"FF",X"FF",X"B7",X"F8",X"00",X"00",X"08",X"E1",X"F0",X"F0",X"F0",X"FC",
		X"00",X"00",X"00",X"00",X"C0",X"FC",X"FF",X"FF",X"00",X"88",X"BF",X"BF",X"D7",X"00",X"00",X"00",
		X"FF",X"FF",X"F7",X"FC",X"FF",X"FF",X"F7",X"FC",X"00",X"00",X"87",X"F0",X"F0",X"F0",X"F0",X"FC",
		X"00",X"00",X"00",X"00",X"E8",X"FF",X"9F",X"FF",X"00",X"88",X"DF",X"FF",X"B7",X"00",X"00",X"00",
		X"FF",X"FF",X"F7",X"F8",X"FF",X"FF",X"F7",X"FC",X"00",X"0C",X"F0",X"F0",X"F8",X"F3",X"F0",X"FE",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"9F",X"FF",X"00",X"88",X"EF",X"FF",X"7F",X"10",X"00",X"00",
		X"FF",X"FF",X"F7",X"F0",X"FC",X"FF",X"F7",X"FE",X"0E",X"C3",X"78",X"E1",X"F8",X"F7",X"F0",X"FE",
		X"00",X"00",X"00",X"00",X"EE",X"FF",X"FF",X"FF",X"00",X"00",X"EF",X"FF",X"FF",X"01",X"00",X"00",
		X"FF",X"FF",X"FF",X"F1",X"F0",X"FF",X"F7",X"FE",X"00",X"86",X"96",X"F2",X"FE",X"F6",X"F0",X"FE",
		X"00",X"00",X"80",X"F0",X"CC",X"FF",X"9F",X"33",X"00",X"00",X"EF",X"FF",X"FF",X"01",X"00",X"00",
		X"FF",X"FF",X"FF",X"F7",X"F0",X"FE",X"F7",X"FF",X"00",X"08",X"E1",X"F2",X"FE",X"FC",X"F0",X"F7",
		X"00",X"00",X"C0",X"F0",X"98",X"00",X"9F",X"C0",X"00",X"00",X"EF",X"FF",X"FF",X"01",X"00",X"00",
		X"FF",X"FF",X"F7",X"FE",X"F3",X"FC",X"F7",X"FF",X"00",X"86",X"F8",X"F7",X"F6",X"FC",X"F9",X"F7",
		X"00",X"00",X"68",X"87",X"30",X"F0",X"00",X"F0",X"00",X"00",X"CE",X"FF",X"FF",X"01",X"00",X"00",
		X"EE",X"FF",X"F7",X"F8",X"F7",X"FE",X"F7",X"FF",X"08",X"E1",X"FC",X"FD",X"F6",X"F8",X"F9",X"F7",
		X"00",X"00",X"3E",X"0F",X"3D",X"F0",X"0F",X"F0",X"00",X"00",X"CE",X"FF",X"FF",X"01",X"00",X"00",
		X"88",X"FF",X"F7",X"FF",X"F7",X"FF",X"F7",X"F7",X"87",X"F0",X"F6",X"FD",X"F7",X"F8",X"FB",X"F7",
		X"00",X"08",X"FF",X"FF",X"3F",X"F0",X"F0",X"FC",X"00",X"00",X"8C",X"FF",X"FF",X"01",X"00",X"00",
		X"04",X"EE",X"F7",X"FF",X"FF",X"FF",X"77",X"F0",X"08",X"C3",X"F2",X"F8",X"F5",X"F0",X"F3",X"F7",
		X"00",X"68",X"7F",X"8F",X"3F",X"FF",X"0F",X"FF",X"00",X"00",X"4C",X"EF",X"7F",X"00",X"00",X"00",
		X"0C",X"89",X"77",X"EE",X"FF",X"FF",X"7F",X"87",X"00",X"0C",X"E1",X"F0",X"F1",X"F0",X"F3",X"F3",
		X"88",X"7F",X"3F",X"0F",X"3F",X"FF",X"0F",X"FF",X"00",X"00",X"EE",X"FF",X"3F",X"00",X"00",X"00",
		X"0C",X"07",X"08",X"01",X"EE",X"FF",X"3B",X"87",X"00",X"00",X"0E",X"E1",X"F0",X"F0",X"FE",X"F3",
		X"00",X"6E",X"7F",X"8F",X"3F",X"FF",X"F0",X"FF",X"00",X"00",X"FF",X"FF",X"53",X"00",X"00",X"00",
		X"CC",X"3F",X"87",X"0F",X"01",X"00",X"48",X"87",X"00",X"08",X"E1",X"1E",X"F0",X"F0",X"FE",X"F3",
		X"00",X"08",X"FF",X"FF",X"3F",X"FF",X"0F",X"FF",X"00",X"00",X"FF",X"FF",X"F7",X"00",X"00",X"00",
		X"CC",X"FF",X"B7",X"7F",X"0F",X"0F",X"CB",X"97",X"00",X"86",X"F0",X"F0",X"F0",X"F0",X"FC",X"F3",
		X"00",X"00",X"3F",X"0F",X"33",X"FF",X"00",X"FF",X"00",X"88",X"FF",X"FF",X"7F",X"10",X"00",X"00",
		X"CC",X"FF",X"F7",X"FE",X"FF",X"FF",X"DB",X"B7",X"0C",X"E1",X"F0",X"F0",X"F0",X"F0",X"F8",X"F1",
		X"00",X"00",X"6E",X"8F",X"D1",X"00",X"1E",X"CC",X"00",X"88",X"FF",X"FF",X"7F",X"10",X"00",X"00",
		X"CC",X"FF",X"F7",X"FC",X"FF",X"FF",X"FB",X"F7",X"00",X"86",X"F0",X"F0",X"F0",X"F0",X"F8",X"F1",
		X"00",X"00",X"DC",X"FF",X"E0",X"D2",X"5A",X"30",X"00",X"88",X"FF",X"FF",X"7F",X"10",X"00",X"00",
		X"CC",X"FF",X"F7",X"F0",X"FB",X"FF",X"FB",X"F7",X"00",X"08",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"B8",X"77",X"E1",X"D2",X"5A",X"F0",X"00",X"88",X"FF",X"FF",X"7F",X"10",X"00",X"00",
		X"CC",X"FF",X"FF",X"F3",X"F0",X"FF",X"FB",X"F7",X"00",X"00",X"00",X"87",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"70",X"80",X"E1",X"D2",X"1E",X"F0",X"00",X"00",X"FF",X"DF",X"B7",X"10",X"00",X"00",
		X"88",X"FF",X"FF",X"FF",X"F0",X"FF",X"FB",X"F7",X"00",X"00",X"00",X"08",X"87",X"F0",X"F0",X"F0",
		X"00",X"00",X"F0",X"F0",X"E1",X"D2",X"5A",X"F0",X"00",X"00",X"EF",X"EF",X"B7",X"00",X"00",X"00",
		X"00",X"FF",X"F7",X"FC",X"F3",X"FF",X"FB",X"F3",X"00",X"00",X"08",X"87",X"F0",X"F0",X"B4",X"F0",
		X"00",X"00",X"F0",X"F0",X"E1",X"D2",X"5A",X"F0",X"00",X"00",X"0E",X"FF",X"D3",X"00",X"00",X"00",
		X"00",X"CC",X"F7",X"FF",X"FB",X"FF",X"33",X"F0",X"00",X"00",X"87",X"F0",X"F0",X"F0",X"B4",X"F0",
		X"00",X"00",X"F0",X"F0",X"E1",X"D2",X"1E",X"F0",X"00",X"00",X"EE",X"FF",X"53",X"00",X"00",X"00",
		X"00",X"00",X"77",X"EE",X"FF",X"FF",X"33",X"F0",X"00",X"00",X"08",X"C3",X"F0",X"F0",X"B4",X"F0",
		X"00",X"00",X"F3",X"F0",X"EF",X"D3",X"5A",X"FF",X"00",X"00",X"CC",X"FF",X"61",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"EE",X"FF",X"11",X"F0",X"00",X"00",X"00",X"0C",X"E1",X"F0",X"B4",X"F0",
		X"00",X"00",X"EE",X"FF",X"EF",X"DF",X"59",X"FF",X"00",X"00",X"88",X"FF",X"21",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"0E",X"F0",X"D2",X"F0",
		X"00",X"00",X"CC",X"FF",X"00",X"CC",X"11",X"FF",X"00",X"00",X"00",X"6E",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"87",X"D2",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",
		X"00",X"00",X"0E",X"09",X"0F",X"0F",X"01",X"F0",X"00",X"00",X"00",X"00",X"00",X"08",X"C3",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"53",X"00",
		X"00",X"08",X"0F",X"2D",X"CF",X"3F",X"1E",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"C2",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"B7",X"00",
		X"00",X"0E",X"0F",X"2D",X"FF",X"7F",X"2D",X"E1",X"00",X"00",X"00",X"00",X"00",X"84",X"E1",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"B7",X"00",
		X"00",X"0F",X"EF",X"E9",X"FF",X"FF",X"4B",X"E1",X"00",X"00",X"00",X"00",X"00",X"4B",X"E1",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"7F",X"10",
		X"00",X"CF",X"FF",X"F1",X"FF",X"FE",X"DB",X"F1",X"00",X"00",X"00",X"00",X"0C",X"F0",X"E1",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"7F",X"10",
		X"00",X"FF",X"FF",X"F1",X"FC",X"FC",X"FB",X"F1",X"00",X"00",X"00",X"00",X"C2",X"78",X"F0",X"F0",
		X"80",X"F0",X"F0",X"F0",X"F0",X"34",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"7F",X"10",
		X"00",X"FF",X"FF",X"F1",X"F0",X"FC",X"FB",X"F1",X"00",X"00",X"00",X"00",X"0C",X"78",X"F0",X"F0",
		X"E0",X"F0",X"F0",X"F0",X"F0",X"78",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"6F",X"10",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FC",X"FB",X"F1",X"00",X"00",X"00",X"00",X"00",X"4B",X"F0",X"F0",
		X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"6E",X"7F",X"10",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FC",X"FB",X"F1",X"00",X"00",X"00",X"00",X"00",X"84",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"8C",X"7F",X"10",
		X"00",X"FF",X"FF",X"F1",X"FF",X"FC",X"FB",X"F1",X"00",X"00",X"00",X"00",X"00",X"8C",X"F1",X"F0",
		X"F0",X"78",X"0F",X"0F",X"0F",X"F1",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"7F",X"10",
		X"00",X"FF",X"FF",X"F9",X"FF",X"FE",X"FB",X"F1",X"00",X"00",X"00",X"00",X"00",X"8C",X"F7",X"F0",
		X"F0",X"1E",X"0F",X"0F",X"0F",X"E3",X"47",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"37",X"00",
		X"00",X"FF",X"FF",X"FD",X"FF",X"FF",X"FB",X"F1",X"00",X"00",X"00",X"00",X"00",X"CE",X"F3",X"F0",
		X"F0",X"1E",X"0F",X"0F",X"0F",X"E3",X"47",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"7F",X"00",
		X"00",X"FF",X"FF",X"FD",X"FF",X"FF",X"FB",X"F1",X"00",X"00",X"00",X"00",X"00",X"CE",X"F0",X"F0",
		X"F0",X"0F",X"F1",X"F0",X"3C",X"C7",X"CF",X"11",X"00",X"26",X"00",X"00",X"00",X"88",X"7F",X"00",
		X"00",X"EE",X"FF",X"FD",X"FF",X"FF",X"FD",X"F1",X"00",X"00",X"00",X"00",X"00",X"EF",X"F0",X"F0",
		X"F0",X"8F",X"F0",X"F0",X"78",X"C7",X"CF",X"FF",X"00",X"7F",X"10",X"00",X"40",X"00",X"7F",X"00",
		X"00",X"88",X"FF",X"FD",X"FF",X"FF",X"FE",X"F0",X"00",X"00",X"00",X"00",X"08",X"FF",X"F0",X"F0",
		X"F0",X"0F",X"F1",X"F0",X"3C",X"C7",X"CF",X"FF",X"00",X"FF",X"21",X"00",X"73",X"00",X"6F",X"00",
		X"00",X"00",X"EE",X"99",X"FF",X"FF",X"11",X"F0",X"00",X"00",X"00",X"00",X"8C",X"F7",X"F2",X"F0",
		X"F0",X"1E",X"0F",X"0F",X"0F",X"E3",X"CF",X"FF",X"00",X"BF",X"21",X"00",X"F7",X"00",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"CE",X"D3",X"F2",X"F0",
		X"F0",X"1E",X"0F",X"0F",X"0F",X"E3",X"CF",X"FF",X"00",X"DF",X"21",X"88",X"FF",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"EF",X"D3",X"F7",X"F0",
		X"F0",X"78",X"0F",X"0F",X"8F",X"F0",X"CF",X"11",X"00",X"EE",X"21",X"88",X"FF",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"CC",X"FF",X"00",X"F0",X"00",X"00",X"00",X"00",X"CE",X"E1",X"F7",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"47",X"00",X"00",X"EE",X"21",X"CC",X"FF",X"31",X"00",X"00",
		X"00",X"00",X"00",X"88",X"FF",X"FF",X"11",X"F0",X"00",X"00",X"00",X"00",X"8C",X"EF",X"F2",X"F0",
		X"F0",X"78",X"8F",X"78",X"8F",X"F0",X"47",X"00",X"00",X"6E",X"10",X"CC",X"FF",X"31",X"00",X"00",
		X"00",X"88",X"33",X"FF",X"FB",X"FF",X"31",X"F0",X"00",X"00",X"00",X"00",X"08",X"FE",X"F2",X"F0",
		X"F0",X"1E",X"8F",X"78",X"0F",X"E3",X"03",X"00",X"00",X"4C",X"10",X"CC",X"FF",X"31",X"00",X"00",
		X"00",X"EE",X"FB",X"FF",X"F3",X"FF",X"FD",X"F0",X"00",X"00",X"00",X"00",X"08",X"F7",X"F0",X"F0",
		X"F0",X"1E",X"8F",X"78",X"0F",X"E3",X"03",X"00",X"00",X"84",X"00",X"CE",X"FF",X"73",X"00",X"00",
		X"88",X"FF",X"FB",X"FE",X"F3",X"FE",X"FD",X"F1",X"00",X"00",X"00",X"00",X"8C",X"F3",X"F0",X"F0",
		X"F0",X"0F",X"F1",X"F0",X"3C",X"C7",X"03",X"00",X"00",X"00",X"00",X"CE",X"FF",X"73",X"00",X"00",
		X"CC",X"FF",X"F3",X"FF",X"F0",X"FE",X"FD",X"F1",X"00",X"00",X"00",X"00",X"CE",X"F1",X"F0",X"F0",
		X"F0",X"8F",X"F0",X"F0",X"78",X"C7",X"03",X"00",X"00",X"00",X"00",X"CE",X"FF",X"73",X"00",X"00",
		X"CC",X"FF",X"FF",X"F3",X"F0",X"FF",X"FD",X"F1",X"00",X"00",X"00",X"00",X"EB",X"F0",X"F0",X"F0",
		X"F0",X"0F",X"F1",X"F0",X"3C",X"C7",X"03",X"00",X"00",X"00",X"00",X"CE",X"FF",X"73",X"00",X"00",
		X"CC",X"FF",X"FF",X"F0",X"FF",X"FF",X"ED",X"F1",X"00",X"00",X"00",X"00",X"FE",X"F6",X"F1",X"F3",
		X"F0",X"1E",X"0F",X"0F",X"0F",X"E3",X"03",X"00",X"00",X"00",X"00",X"CE",X"FF",X"03",X"00",X"00",
		X"CC",X"FF",X"F3",X"F8",X"FF",X"7F",X"ED",X"F1",X"00",X"00",X"00",X"08",X"FF",X"F6",X"F1",X"F3",
		X"F0",X"1E",X"0F",X"0F",X"0F",X"E3",X"03",X"00",X"00",X"00",X"00",X"8C",X"FF",X"37",X"00",X"00",
		X"CC",X"FF",X"F3",X"FC",X"FF",X"3F",X"FC",X"E1",X"00",X"00",X"00",X"8C",X"FB",X"F6",X"F9",X"F3",
		X"F0",X"78",X"0F",X"0F",X"8F",X"F0",X"03",X"00",X"00",X"00",X"00",X"8C",X"FF",X"7F",X"00",X"00",
		X"8C",X"FF",X"F3",X"FF",X"FF",X"0F",X"9E",X"E1",X"00",X"00",X"00",X"CE",X"FD",X"F6",X"F8",X"F7",
		X"F0",X"8F",X"F0",X"1E",X"78",X"C7",X"03",X"00",X"00",X"00",X"00",X"08",X"FF",X"FF",X"01",X"00",
		X"0C",X"EF",X"4B",X"0F",X"0F",X"87",X"0F",X"E1",X"00",X"00",X"08",X"EF",X"F4",X"F1",X"F8",X"F7",
		X"F0",X"8F",X"F0",X"1E",X"78",X"C7",X"03",X"00",X"00",X"00",X"00",X"EE",X"FF",X"FF",X"01",X"00",
		X"0C",X"03",X"00",X"00",X"00",X"00",X"0F",X"F0",X"00",X"00",X"00",X"CC",X"F5",X"F1",X"FA",X"F4",
		X"F0",X"8F",X"F0",X"1E",X"78",X"C7",X"03",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"01",X"00",
		X"0C",X"0C",X"0F",X"0F",X"0F",X"0F",X"00",X"F0",X"00",X"00",X"CC",X"FF",X"F1",X"F1",X"FE",X"F4",
		X"F0",X"8F",X"F0",X"1E",X"78",X"C7",X"03",X"00",X"00",X"00",X"00",X"FF",X"FF",X"7F",X"00",X"00",
		X"00",X"0F",X"0F",X"0F",X"0F",X"4B",X"0F",X"E1",X"00",X"0C",X"EF",X"FE",X"F3",X"F0",X"F6",X"F0",
		X"F0",X"8F",X"F0",X"1E",X"78",X"C7",X"47",X"00",X"00",X"00",X"88",X"FF",X"FF",X"7F",X"00",X"00",
		X"0C",X"0F",X"0F",X"0F",X"0F",X"87",X"0F",X"C3",X"00",X"00",X"88",X"FD",X"F2",X"F8",X"F6",X"F0",
		X"F0",X"0F",X"F1",X"1E",X"3C",X"C7",X"47",X"00",X"00",X"00",X"88",X"FF",X"FF",X"6F",X"00",X"00",
		X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"1E",X"C3",X"00",X"00",X"00",X"CC",X"F2",X"F8",X"F4",X"F0",
		X"F0",X"1E",X"0F",X"0F",X"0F",X"E3",X"CF",X"11",X"00",X"00",X"88",X"FF",X"FF",X"1F",X"00",X"00",
		X"0E",X"0F",X"87",X"0F",X"EF",X"7F",X"2D",X"C3",X"00",X"0C",X"EF",X"F7",X"F0",X"FB",X"F0",X"F0",
		X"F0",X"1E",X"0F",X"0F",X"0F",X"E3",X"CF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"53",X"00",X"00",
		X"0E",X"0F",X"87",X"EF",X"FF",X"FF",X"4B",X"C3",X"08",X"8F",X"FF",X"F7",X"FA",X"FB",X"F1",X"F0",
		X"F0",X"78",X"0F",X"0F",X"8F",X"F0",X"CF",X"FF",X"00",X"00",X"00",X"F7",X"FF",X"53",X"00",X"00",
		X"0E",X"FF",X"B7",X"FE",X"FF",X"FF",X"DB",X"D3",X"00",X"0C",X"F0",X"F1",X"FE",X"FF",X"F1",X"F0",
		X"F0",X"F0",X"F0",X"1E",X"78",X"C7",X"CF",X"FF",X"00",X"00",X"00",X"E8",X"FF",X"53",X"00",X"00",
		X"8E",X"FF",X"F7",X"FE",X"FF",X"FF",X"FB",X"F3",X"00",X"00",X"C3",X"F0",X"FF",X"FF",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"1E",X"78",X"C7",X"CF",X"FF",X"00",X"00",X"00",X"CC",X"FF",X"53",X"00",X"00",
		X"CE",X"FF",X"F7",X"FC",X"FF",X"FF",X"FB",X"F3",X"00",X"00",X"08",X"3C",X"8F",X"F5",X"F2",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"78",X"C7",X"CF",X"11",X"00",X"00",X"00",X"CC",X"FF",X"43",X"00",X"00",
		X"EE",X"FF",X"F7",X"F0",X"FF",X"FD",X"FB",X"F3",X"00",X"00",X"00",X"C0",X"7F",X"CF",X"F2",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"78",X"C7",X"47",X"00",X"00",X"00",X"00",X"88",X"7F",X"30",X"00",X"00",
		X"EE",X"FF",X"F7",X"F0",X"FC",X"FC",X"FB",X"F3",X"00",X"00",X"0E",X"FB",X"FF",X"FD",X"FC",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"78",X"C7",X"47",X"00",X"00",X"00",X"00",X"88",X"3F",X"10",X"00",X"00",
		X"EE",X"FF",X"FF",X"F3",X"F1",X"FC",X"FB",X"F3",X"00",X"0E",X"EF",X"FD",X"F7",X"FF",X"F7",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"78",X"C7",X"03",X"00",X"00",X"00",X"00",X"08",X"C3",X"10",X"00",X"00",
		X"EE",X"FF",X"FF",X"FF",X"FF",X"FC",X"FB",X"F3",X"00",X"88",X"FF",X"FD",X"FC",X"F9",X"F1",X"F0",
		X"F0",X"0F",X"0F",X"0F",X"0F",X"C7",X"03",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",
		X"EE",X"FF",X"F7",X"FC",X"FF",X"FC",X"FB",X"F3",X"88",X"FF",X"FB",X"F4",X"FC",X"F1",X"F1",X"F0",
		X"F0",X"0F",X"0F",X"0F",X"0F",X"C7",X"03",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",
		X"CC",X"FF",X"F7",X"F2",X"FF",X"FD",X"FB",X"F3",X"EF",X"FD",X"FB",X"F2",X"FB",X"F0",X"F1",X"F0",
		X"F0",X"0F",X"0F",X"0F",X"0F",X"C7",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"FF",X"F7",X"FF",X"FF",X"FF",X"FB",X"F1",X"00",X"EE",X"F1",X"F7",X"F2",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"1E",X"F0",X"F0",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"EE",X"F7",X"FF",X"FF",X"FF",X"75",X"F0",X"00",X"80",X"FA",X"F7",X"B4",X"F4",X"F0",X"F0",
		X"F0",X"78",X"0F",X"0F",X"0F",X"C7",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"88",X"77",X"EE",X"FF",X"FF",X"11",X"F0",X"00",X"00",X"EE",X"F7",X"F0",X"F4",X"F4",X"F0",
		X"F0",X"1E",X"0F",X"0F",X"0F",X"C7",X"03",X"00",X"00",X"00",X"00",X"13",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"EE",X"FF",X"F9",X"F0",X"F4",X"F0",X"F0",
		X"F0",X"1E",X"0F",X"0F",X"0F",X"C7",X"03",X"00",X"00",X"00",X"88",X"37",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"CF",X"FF",X"F5",X"F9",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"0F",X"E3",X"1E",X"F0",X"F0",X"03",X"00",X"00",X"00",X"CC",X"7F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"0C",X"FF",X"F3",X"F8",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"0F",X"F1",X"1E",X"F0",X"F0",X"03",X"00",X"00",X"00",X"CC",X"7F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"CC",X"F0",X"F8",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"0F",X"E3",X"F0",X"F0",X"F0",X"03",X"00",X"00",X"00",X"EE",X"7F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"0E",X"E1",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"1E",X"0F",X"0F",X"0F",X"C7",X"03",X"00",X"00",X"00",X"EE",X"7F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"1E",X"0F",X"0F",X"0F",X"C7",X"47",X"00",X"00",X"00",X"FF",X"7F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"8E",X"F3",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"78",X"0F",X"0F",X"0F",X"C7",X"47",X"00",X"00",X"00",X"FF",X"7F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"08",X"EF",X"F5",X"F0",X"F2",X"F1",X"F1",
		X"F0",X"F0",X"F0",X"1E",X"F0",X"F0",X"CF",X"11",X"00",X"00",X"EE",X"7F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"0C",X"E1",X"F0",X"F0",X"F8",X"FE",X"F0",
		X"F0",X"0F",X"0F",X"0F",X"8F",X"F0",X"CF",X"FF",X"00",X"00",X"EE",X"7F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"0E",X"F0",X"F0",X"F8",X"FE",X"F1",
		X"F0",X"0F",X"0F",X"0F",X"0F",X"E3",X"CF",X"FF",X"00",X"00",X"CC",X"36",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"0F",X"E1",X"F0",X"F5",X"F1",
		X"F0",X"0F",X"0F",X"0F",X"0F",X"C7",X"CF",X"FF",X"00",X"00",X"CE",X"71",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"0E",X"E1",X"F5",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"3C",X"C7",X"CF",X"FF",X"00",X"00",X"FF",X"73",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"9F",X"E3",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"78",X"C7",X"CF",X"11",X"00",X"00",X"FF",X"73",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"8E",X"FF",X"F3",X"F0",
		X"E1",X"F0",X"F0",X"1E",X"3C",X"C7",X"47",X"00",X"00",X"00",X"FF",X"B7",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"0C",X"EF",X"FF",X"F2",X"FC",
		X"E1",X"F0",X"F0",X"1E",X"0F",X"C7",X"47",X"00",X"00",X"00",X"FF",X"B7",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"CF",X"FF",X"F2",X"F0",X"ED",
		X"C3",X"F0",X"F0",X"1E",X"0F",X"E3",X"03",X"00",X"00",X"00",X"FF",X"B7",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"0C",X"FF",X"FB",X"F0",X"F0",X"EF",
		X"C3",X"F0",X"F0",X"1E",X"8F",X"78",X"03",X"00",X"00",X"00",X"EE",X"B7",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"CF",X"F0",X"F0",X"78",X"FA",
		X"86",X"F0",X"F0",X"F0",X"F0",X"3C",X"01",X"00",X"00",X"00",X"EE",X"B7",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"0C",X"E1",X"F0",X"78",X"FB",
		X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"01",X"00",X"00",X"00",X"CC",X"B7",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"86",X"F0",X"BC",X"FB",
		X"08",X"0F",X"0F",X"0F",X"0F",X"07",X"00",X"00",X"00",X"00",X"0C",X"53",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"08",X"E1",X"DE",X"F1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"43",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"86",X"EF",X"F1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"08",X"FF",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"8C",X"F7",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"CF",X"FF",X"F1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"0C",X"CF",X"F3",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"0C",X"F0",X"F4",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"E1",X"F7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"CE",X"F3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"08",X"EF",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"0E",X"FD",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0E",X"09",X"0F",X"0F",X"01",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"C3",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"0F",X"2D",X"CF",X"3F",X"1E",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"84",X"F0",
		X"00",X"00",X"E0",X"30",X"F0",X"90",X"F0",X"70",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"0F",X"2D",X"FF",X"7F",X"2D",X"E1",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"F0",
		X"00",X"00",X"E0",X"B4",X"F0",X"96",X"F0",X"78",X"FF",X"13",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"EF",X"E9",X"FF",X"FF",X"4B",X"E1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E1",
		X"00",X"30",X"E1",X"B4",X"F0",X"96",X"F0",X"78",X"FF",X"13",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"CF",X"FF",X"F1",X"FF",X"FE",X"DB",X"F1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E1",
		X"80",X"B4",X"E1",X"B4",X"F0",X"F0",X"F0",X"78",X"EE",X"37",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"F1",X"FC",X"FC",X"FB",X"F1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C2",
		X"C0",X"3C",X"E1",X"B4",X"F0",X"96",X"F0",X"78",X"EE",X"37",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"F1",X"F0",X"FC",X"FB",X"F1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C2",
		X"C0",X"B4",X"E1",X"B4",X"F0",X"96",X"F0",X"78",X"CC",X"37",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FC",X"FB",X"F1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"84",
		X"C0",X"3C",X"E1",X"B4",X"F0",X"F0",X"F0",X"78",X"EE",X"37",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FC",X"FB",X"F1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"84",
		X"C0",X"B4",X"E1",X"B4",X"F0",X"96",X"F0",X"78",X"FF",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"F1",X"FF",X"FC",X"FB",X"F1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"8C",
		X"C4",X"3C",X"E1",X"BC",X"FF",X"97",X"F0",X"78",X"FF",X"37",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"F9",X"FF",X"FE",X"FB",X"F1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CE",
		X"CC",X"B4",X"E1",X"BC",X"FF",X"F9",X"FF",X"7F",X"FF",X"37",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"FD",X"FF",X"FF",X"FB",X"F1",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"E3",
		X"CC",X"3F",X"EF",X"BF",X"FF",X"9F",X"FF",X"7F",X"EE",X"17",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"FD",X"FF",X"FF",X"FB",X"F1",X"00",X"00",X"00",X"00",X"00",X"00",X"8F",X"F3",
		X"88",X"B7",X"EF",X"BF",X"FF",X"9F",X"FF",X"7F",X"EE",X"13",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"EE",X"FF",X"FD",X"FF",X"FF",X"FD",X"F1",X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"F1",
		X"00",X"33",X"EF",X"BF",X"FF",X"F9",X"FF",X"7F",X"CC",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"88",X"FF",X"FD",X"FF",X"FF",X"FE",X"F0",X"00",X"00",X"00",X"00",X"0E",X"FF",X"F7",X"F8",
		X"00",X"00",X"EE",X"BF",X"FF",X"9F",X"FF",X"7F",X"08",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"EE",X"99",X"FF",X"FF",X"11",X"F0",X"00",X"00",X"00",X"00",X"00",X"CF",X"F1",X"F8",
		X"00",X"00",X"EE",X"33",X"FF",X"99",X"FF",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"0C",X"F4",X"F5",
		X"00",X"00",X"00",X"00",X"AE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"13",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"CF",X"F5",
		X"00",X"00",X"00",X"00",X"AE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"37",
		X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"0E",X"FF",X"F5",
		X"00",X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"7F",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"11",X"F0",X"00",X"00",X"00",X"00",X"08",X"EF",X"FF",X"F1",
		X"00",X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"7F",
		X"00",X"88",X"77",X"EE",X"FB",X"FF",X"31",X"F0",X"00",X"00",X"00",X"0E",X"8F",X"FF",X"F7",X"F3",
		X"00",X"00",X"00",X"00",X"AE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"7F",
		X"00",X"EE",X"F7",X"FF",X"F3",X"FF",X"FD",X"F0",X"00",X"00",X"0E",X"EF",X"F7",X"FF",X"F4",X"F3",
		X"00",X"00",X"C0",X"F0",X"AE",X"C0",X"10",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"7F",
		X"00",X"FF",X"F7",X"FE",X"F3",X"FE",X"FD",X"F1",X"00",X"00",X"00",X"0E",X"FE",X"F0",X"FF",X"F2",
		X"00",X"00",X"E0",X"F0",X"E1",X"D2",X"5A",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"7F",
		X"88",X"FF",X"F7",X"FF",X"F0",X"FE",X"FD",X"F1",X"00",X"00",X"00",X"00",X"C3",X"F1",X"F3",X"FA",
		X"00",X"00",X"F0",X"F0",X"E1",X"D2",X"5A",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"7F",
		X"88",X"FF",X"FF",X"F3",X"F0",X"FF",X"FD",X"F1",X"00",X"00",X"00",X"00",X"84",X"F1",X"F0",X"F8",
		X"00",X"00",X"F0",X"F0",X"E1",X"D2",X"1E",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"7F",
		X"88",X"FF",X"FF",X"F0",X"FF",X"FF",X"ED",X"F1",X"00",X"00",X"00",X"00",X"0C",X"EB",X"F0",X"F1",
		X"00",X"00",X"F0",X"F0",X"E1",X"D2",X"5A",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"37",
		X"88",X"FF",X"F7",X"F8",X"FF",X"FF",X"AD",X"F1",X"00",X"00",X"00",X"0C",X"CF",X"F7",X"F7",X"F1",
		X"00",X"00",X"F0",X"F0",X"E1",X"D2",X"5A",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"EF",X"12",
		X"88",X"FF",X"F7",X"FC",X"FF",X"7F",X"3C",X"E1",X"00",X"00",X"08",X"CF",X"F7",X"F4",X"F2",X"F4",
		X"00",X"00",X"F0",X"F0",X"E1",X"D2",X"1E",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"DF",X"71",
		X"88",X"FF",X"F7",X"FF",X"FF",X"3F",X"1E",X"E1",X"00",X"00",X"8E",X"F7",X"F7",X"F9",X"F5",X"F6",
		X"00",X"00",X"F3",X"F0",X"EF",X"D3",X"5A",X"FF",X"00",X"00",X"00",X"00",X"00",X"88",X"FF",X"73",
		X"08",X"EF",X"B7",X"EF",X"FF",X"97",X"0F",X"E1",X"00",X"00",X"08",X"6B",X"F7",X"FB",X"FD",X"F2",
		X"00",X"00",X"EE",X"FF",X"EF",X"DF",X"5B",X"FF",X"00",X"00",X"00",X"00",X"00",X"88",X"FF",X"73",
		X"08",X"0F",X"87",X"CF",X"7F",X"0F",X"0F",X"E1",X"00",X"00",X"00",X"86",X"F9",X"FA",X"FD",X"F2",
		X"00",X"00",X"CC",X"FF",X"AE",X"CC",X"11",X"FF",X"00",X"00",X"00",X"00",X"00",X"88",X"FF",X"B7",
		X"08",X"0F",X"87",X"0F",X"0F",X"0F",X"0F",X"E1",X"00",X"00",X"08",X"CF",X"F9",X"F4",X"F6",X"F7",
		X"00",X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"FF",X"B7",
		X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"E1",X"00",X"00",X"8F",X"FF",X"F2",X"F0",X"F6",X"F5",
		X"00",X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F7",X"B7",
		X"00",X"0C",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"00",X"00",X"08",X"C7",X"F4",X"F1",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"AE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E8",X"B7",
		X"00",X"00",X"0F",X"0F",X"03",X"00",X"00",X"F0",X"00",X"00",X"00",X"0C",X"F0",X"F9",X"E9",X"F2",
		X"00",X"00",X"00",X"E0",X"F0",X"30",X"F0",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"B7",
		X"00",X"00",X"00",X"00",X"CC",X"FF",X"11",X"F0",X"00",X"00",X"00",X"00",X"C0",X"CF",X"E5",X"F2",
		X"00",X"00",X"80",X"E1",X"B4",X"3C",X"F0",X"2E",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"B7",
		X"00",X"88",X"FF",X"CC",X"FF",X"FF",X"33",X"F0",X"00",X"00",X"00",X"00",X"00",X"FE",X"E7",X"F3",
		X"00",X"00",X"E0",X"E1",X"B4",X"3C",X"F0",X"2F",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"53",
		X"00",X"EE",X"FF",X"FE",X"FF",X"FF",X"73",X"F0",X"00",X"00",X"00",X"00",X"C3",X"7A",X"F6",X"F5",
		X"00",X"C0",X"E1",X"E1",X"F0",X"3C",X"F0",X"2F",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"43",
		X"88",X"FF",X"FF",X"F8",X"FF",X"FE",X"FB",X"F1",X"00",X"00",X"00",X"00",X"0C",X"69",X"FF",X"F4",
		X"00",X"D2",X"E1",X"E1",X"B4",X"3C",X"F0",X"2F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",
		X"CC",X"FF",X"FF",X"FC",X"FF",X"FC",X"FB",X"F3",X"00",X"00",X"00",X"00",X"00",X"86",X"F9",X"F4",
		X"80",X"D2",X"E1",X"E1",X"B4",X"3C",X"F0",X"2F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"FF",X"FF",X"FF",X"F3",X"FC",X"FB",X"F3",X"00",X"00",X"00",X"00",X"00",X"08",X"F1",X"F4",
		X"84",X"D2",X"E1",X"E1",X"F0",X"3C",X"F0",X"2F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"FF",X"FF",X"F3",X"F0",X"FC",X"FB",X"F3",X"00",X"00",X"00",X"00",X"00",X"84",X"F4",X"FC",
		X"84",X"D2",X"E1",X"E1",X"B4",X"3C",X"F0",X"2F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"FF",X"FF",X"F0",X"FE",X"FE",X"FB",X"F3",X"00",X"00",X"00",X"00",X"0F",X"8F",X"F4",X"FD",
		X"84",X"D2",X"E1",X"E1",X"B4",X"3C",X"F0",X"2F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"8C",X"FF",X"FF",X"F8",X"FF",X"FF",X"DB",X"F3",X"00",X"00",X"00",X"00",X"00",X"0F",X"F8",X"FB",
		X"88",X"D3",X"E1",X"E1",X"F0",X"3C",X"F0",X"2F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"FF",X"7F",X"BC",X"EF",X"FF",X"4B",X"D3",X"00",X"00",X"00",X"00",X"00",X"00",X"CB",X"FF",
		X"00",X"DF",X"E1",X"E1",X"B4",X"3C",X"F0",X"2F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"0F",X"0F",X"3C",X"0F",X"3F",X"4B",X"C3",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"F7",
		X"00",X"CC",X"EF",X"EF",X"BF",X"3F",X"FF",X"2F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"0F",X"0F",X"1E",X"0F",X"0F",X"69",X"C3",X"00",X"00",X"00",X"00",X"00",X"08",X"E9",X"F6",
		X"00",X"00",X"EE",X"EF",X"FF",X"3F",X"FF",X"2F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"00",X"00",X"00",X"08",X"0F",X"2D",X"C3",X"00",X"00",X"00",X"00",X"00",X"8E",X"F9",X"F4",
		X"00",X"E0",X"98",X"EF",X"BF",X"3F",X"FF",X"2E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"0F",X"0F",X"0F",X"07",X"00",X"0C",X"C3",X"00",X"00",X"00",X"00",X"8E",X"E9",X"F4",X"F2",
		X"00",X"F0",X"70",X"EE",X"BF",X"33",X"FF",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"0F",X"0F",X"0F",X"0F",X"0F",X"03",X"F0",X"00",X"00",X"00",X"08",X"EB",X"F0",X"F6",X"F1",
		X"00",X"F0",X"F0",X"01",X"00",X"C0",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"87",X"00",X"00",X"00",X"87",X"FE",X"F0",X"F2",X"F5",
		X"00",X"F0",X"F0",X"87",X"F0",X"D2",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"0F",X"87",X"8F",X"FF",X"D3",X"0F",X"0F",X"00",X"00",X"00",X"08",X"E5",X"F4",X"FF",X"F4",
		X"00",X"F0",X"F0",X"A5",X"F0",X"D2",X"87",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"FF",X"87",X"EF",X"FF",X"B7",X"3C",X"0F",X"00",X"00",X"00",X"00",X"86",X"C7",X"F9",X"F5",
		X"00",X"F0",X"F0",X"87",X"F0",X"D2",X"87",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CF",X"FF",X"97",X"FE",X"FF",X"7F",X"F0",X"0F",X"00",X"00",X"00",X"00",X"00",X"3F",X"F1",X"FD",
		X"00",X"F0",X"F0",X"A5",X"F0",X"D2",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CF",X"FF",X"B7",X"FE",X"FF",X"FF",X"D3",X"3C",X"00",X"00",X"00",X"00",X"00",X"84",X"F1",X"FF",
		X"00",X"F0",X"F0",X"87",X"F0",X"D2",X"87",X"F0",X"00",X"00",X"00",X"17",X"00",X"00",X"00",X"00",
		X"EF",X"FF",X"F7",X"FE",X"FF",X"FF",X"B7",X"F0",X"00",X"00",X"00",X"00",X"0C",X"87",X"F2",X"FA",
		X"00",X"F1",X"F0",X"A5",X"F0",X"D2",X"87",X"F0",X"00",X"00",X"88",X"7F",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"F7",X"F8",X"FF",X"FF",X"7F",X"F0",X"00",X"00",X"00",X"00",X"CF",X"F4",X"F2",X"FA",
		X"00",X"F3",X"F0",X"8F",X"FF",X"D3",X"F8",X"FF",X"00",X"00",X"CC",X"7F",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"F7",X"F0",X"FF",X"FF",X"FF",X"78",X"00",X"00",X"00",X"0E",X"EF",X"F0",X"F8",X"F5",
		X"00",X"EE",X"FF",X"AF",X"FF",X"DF",X"8F",X"FF",X"00",X"00",X"8C",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"F7",X"F0",X"F4",X"FF",X"FF",X"3C",X"00",X"00",X"0C",X"CF",X"F3",X"F1",X"F0",X"F0",
		X"00",X"CC",X"FF",X"8F",X"FF",X"DF",X"8F",X"FF",X"00",X"00",X"6E",X"FF",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"F1",X"F0",X"FC",X"FF",X"3C",X"00",X"00",X"00",X"86",X"FD",X"F0",X"E1",X"F0",
		X"00",X"88",X"FF",X"01",X"00",X"CC",X"88",X"FF",X"00",X"00",X"FF",X"CF",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"F7",X"F0",X"FC",X"FF",X"1E",X"00",X"00",X"00",X"08",X"F8",X"F0",X"E5",X"F1",
		X"00",X"00",X"00",X"E0",X"F0",X"30",X"00",X"00",X"00",X"88",X"FF",X"FF",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"F7",X"FE",X"F3",X"FC",X"FF",X"9E",X"00",X"00",X"08",X"8F",X"F0",X"78",X"F5",X"F5",
		X"00",X"00",X"00",X"E1",X"F0",X"3C",X"00",X"0E",X"00",X"88",X"FF",X"FF",X"13",X"00",X"00",X"00",
		X"EE",X"FF",X"F7",X"F8",X"F7",X"FE",X"FF",X"9E",X"00",X"00",X"8E",X"F7",X"F0",X"B4",X"F7",X"F7",
		X"00",X"00",X"80",X"E1",X"F0",X"3C",X"10",X"0F",X"00",X"88",X"FF",X"FF",X"13",X"00",X"00",X"00",
		X"88",X"FF",X"F7",X"FF",X"F7",X"FF",X"FF",X"DE",X"00",X"0C",X"ED",X"F1",X"F0",X"D6",X"F6",X"F6",
		X"00",X"00",X"C0",X"E1",X"F0",X"3C",X"38",X"01",X"00",X"88",X"FF",X"FF",X"13",X"00",X"00",X"00",
		X"00",X"EE",X"F7",X"FF",X"FF",X"FF",X"FF",X"E7",X"00",X"00",X"0E",X"F2",X"F4",X"E9",X"F2",X"F2",
		X"00",X"00",X"C2",X"E1",X"F0",X"3C",X"3C",X"00",X"00",X"00",X"FF",X"FF",X"13",X"00",X"00",X"00",
		X"00",X"88",X"77",X"EE",X"FF",X"FF",X"FF",X"F0",X"00",X"00",X"00",X"87",X"3C",X"FB",X"F2",X"F1",
		X"00",X"00",X"D2",X"E1",X"F0",X"3C",X"34",X"00",X"00",X"00",X"FF",X"FF",X"13",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"EE",X"FF",X"FF",X"F0",X"00",X"00",X"00",X"08",X"CF",X"F3",X"F0",X"F1",
		X"00",X"80",X"D2",X"E1",X"F0",X"3C",X"34",X"00",X"00",X"00",X"EE",X"FF",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"88",X"FF",X"77",X"F0",X"00",X"00",X"00",X"0E",X"F3",X"F5",X"F0",X"F1",
		X"00",X"84",X"D2",X"E1",X"F0",X"3C",X"34",X"00",X"00",X"00",X"EE",X"FF",X"13",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"0C",X"EF",X"FD",X"78",X"F8",X"F8",
		X"00",X"A4",X"D2",X"E1",X"F0",X"00",X"24",X"08",X"00",X"00",X"0E",X"FF",X"37",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"0E",X"CF",X"F7",X"F0",X"B4",X"F8",X"FC",
		X"00",X"B4",X"D2",X"E1",X"70",X"F0",X"14",X"0E",X"00",X"00",X"EF",X"EF",X"37",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"0E",X"FB",X"F0",X"C7",X"F8",X"FC",
		X"00",X"A6",X"D2",X"E1",X"38",X"F0",X"12",X"07",X"00",X"08",X"FF",X"FF",X"37",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"87",X"3C",X"F6",X"F0",X"FD",
		X"00",X"8C",X"D3",X"E1",X"58",X"F0",X"5A",X"00",X"00",X"08",X"FF",X"FF",X"37",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"08",X"C7",X"F0",X"F0",X"FB",
		X"00",X"88",X"DF",X"E1",X"4A",X"F0",X"D2",X"00",X"00",X"88",X"FF",X"FF",X"37",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"8E",X"F6",X"F4",X"F2",X"F2",
		X"00",X"00",X"DF",X"67",X"5A",X"F0",X"D2",X"0C",X"00",X"88",X"FF",X"FF",X"13",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"08",X"EF",X"FF",X"F0",X"F0",X"F2",
		X"00",X"00",X"CE",X"A3",X"5B",X"F0",X"DA",X"0F",X"00",X"88",X"FF",X"7F",X"63",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"8E",X"F7",X"F6",X"F1",X"F0",X"F2",
		X"00",X"00",X"CC",X"67",X"5F",X"F0",X"DE",X"0C",X"00",X"00",X"FF",X"FF",X"73",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"08",X"EF",X"FB",X"FD",X"F1",X"F0",X"F2",
		X"00",X"00",X"88",X"EF",X"4E",X"FF",X"DF",X"00",X"00",X"00",X"FF",X"FF",X"73",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"8F",X"FF",X"F4",X"F9",X"F1",X"F7",X"F3",
		X"00",X"00",X"00",X"EF",X"5D",X"FF",X"5F",X"00",X"00",X"00",X"EE",X"FF",X"31",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"0F",X"FF",X"F7",X"F1",X"F0",X"F9",X"F9",X"F3",
		X"00",X"00",X"00",X"EE",X"3B",X"FF",X"13",X"07",X"00",X"00",X"CC",X"FF",X"31",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"08",X"CF",X"F1",X"FA",X"F0",X"FD",X"F8",X"F3",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"11",X"0E",X"00",X"00",X"CC",X"FF",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"0C",X"F0",X"F0",X"F4",X"FD",X"F0",X"F1",
		X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"08",X"00",X"00",X"80",X"F7",X"00",X"00",X"00",X"00",
		X"00",X"08",X"0F",X"0C",X"0F",X"0F",X"03",X"F0",X"00",X"00",X"C3",X"F0",X"F6",X"FC",X"F4",X"F1",
		X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"80",X"F3",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"0F",X"1E",X"0F",X"0F",X"2D",X"E1",X"00",X"00",X"0C",X"F0",X"FA",X"F2",X"F8",X"F1",
		X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"22",X"00",
		X"00",X"0F",X"0F",X"1E",X"FF",X"3F",X"4B",X"C3",X"00",X"00",X"00",X"CF",X"F9",X"F3",X"F0",X"F5",
		X"00",X"00",X"C2",X"78",X"F0",X"06",X"78",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"E6",X"00",
		X"08",X"EF",X"3F",X"BC",X"FF",X"FF",X"4B",X"C3",X"00",X"00",X"0C",X"FF",X"FD",X"F8",X"F2",X"F1",
		X"00",X"00",X"D2",X"78",X"F0",X"0F",X"78",X"78",X"00",X"00",X"00",X"00",X"00",X"88",X"FF",X"10",
		X"0C",X"FF",X"7F",X"F8",X"FF",X"FF",X"DB",X"D3",X"00",X"08",X"8F",X"FD",X"F6",X"F8",X"FB",X"F0",
		X"00",X"80",X"D2",X"78",X"F0",X"0F",X"78",X"78",X"00",X"00",X"00",X"00",X"00",X"88",X"FF",X"10",
		X"8C",X"FF",X"FF",X"F0",X"FE",X"FD",X"FB",X"F3",X"00",X"00",X"08",X"C3",X"F0",X"F0",X"FA",X"F0",
		X"00",X"80",X"D2",X"78",X"FF",X"0F",X"78",X"78",X"00",X"00",X"00",X"00",X"00",X"80",X"FE",X"10",
		X"CC",X"FF",X"FF",X"F0",X"F0",X"FC",X"FB",X"F3",X"00",X"00",X"00",X"0C",X"E1",X"F0",X"FA",X"F0",
		X"00",X"80",X"DF",X"7F",X"FF",X"0F",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",X"C8",X"FF",X"10",
		X"CC",X"FF",X"FF",X"FF",X"FF",X"FC",X"FB",X"F3",X"00",X"00",X"00",X"00",X"86",X"F4",X"F4",X"F0",
		X"00",X"88",X"DF",X"7F",X"FF",X"0F",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",X"CC",X"FF",X"10",
		X"CC",X"FF",X"FF",X"FF",X"FF",X"FC",X"FB",X"F3",X"00",X"00",X"00",X"00",X"08",X"E9",X"F0",X"F6",
		X"00",X"00",X"DF",X"7F",X"FF",X"00",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",X"CC",X"F7",X"00",
		X"CC",X"FF",X"FF",X"F0",X"FE",X"FD",X"FB",X"F3",X"00",X"00",X"00",X"00",X"00",X"86",X"F4",X"F7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"37",X"00",
		X"CC",X"FF",X"FF",X"FC",X"FF",X"FD",X"FB",X"F3",X"00",X"00",X"00",X"00",X"00",X"08",X"7F",X"F5",
		X"00",X"00",X"80",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"7F",X"00",
		X"CC",X"FF",X"FF",X"FC",X"FF",X"FF",X"FB",X"F3",X"00",X"00",X"00",X"00",X"00",X"8E",X"7B",X"F7",
		X"00",X"00",X"C0",X"F0",X"10",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"88",X"7F",X"00",
		X"88",X"FF",X"FF",X"FC",X"FF",X"FF",X"FB",X"F3",X"00",X"00",X"00",X"00",X"0C",X"EF",X"BD",X"F7",
		X"00",X"00",X"68",X"87",X"30",X"F0",X"00",X"F0",X"00",X"00",X"00",X"00",X"40",X"00",X"7F",X"00",
		X"00",X"FF",X"FF",X"FC",X"FF",X"FF",X"FB",X"F3",X"00",X"00",X"00",X"00",X"00",X"86",X"BC",X"F3",
		X"00",X"00",X"3E",X"0F",X"3D",X"F0",X"0F",X"F0",X"00",X"00",X"00",X"00",X"70",X"00",X"6F",X"00",
		X"00",X"EE",X"FF",X"FE",X"FF",X"FF",X"FD",X"F1",X"00",X"00",X"00",X"00",X"00",X"08",X"DE",X"FB",
		X"00",X"00",X"FF",X"FF",X"3F",X"F0",X"F0",X"FC",X"00",X"00",X"00",X"00",X"F3",X"00",X"06",X"00",
		X"00",X"88",X"FF",X"44",X"FF",X"FF",X"33",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"ED",X"FF",
		X"00",X"00",X"7F",X"8F",X"3F",X"FF",X"0F",X"FF",X"00",X"00",X"00",X"88",X"F7",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"0C",X"F7",X"FC",
		X"00",X"00",X"3F",X"0F",X"3F",X"FF",X"0F",X"FF",X"00",X"00",X"00",X"88",X"FF",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"CF",X"F7",X"F4",
		X"00",X"00",X"7F",X"8F",X"3F",X"FF",X"F0",X"FF",X"00",X"00",X"00",X"CC",X"FF",X"31",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"11",X"F0",X"00",X"00",X"00",X"00",X"00",X"0C",X"F0",X"F4",
		X"00",X"00",X"FF",X"FF",X"3F",X"FF",X"0F",X"FF",X"00",X"00",X"00",X"CC",X"FF",X"31",X"00",X"00",
		X"00",X"88",X"77",X"EE",X"FB",X"FF",X"31",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"CB",X"F4",
		X"00",X"00",X"3F",X"0F",X"33",X"FF",X"00",X"FF",X"00",X"00",X"00",X"CC",X"FF",X"31",X"00",X"00",
		X"00",X"EE",X"F7",X"FF",X"F3",X"FF",X"FD",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"84",X"F3",
		X"00",X"00",X"6E",X"8F",X"11",X"00",X"00",X"CC",X"00",X"00",X"00",X"CE",X"FF",X"73",X"00",X"00",
		X"00",X"FF",X"F7",X"FE",X"F3",X"FE",X"FD",X"F1",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"F3",
		X"00",X"00",X"CC",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CE",X"FF",X"73",X"00",X"00",
		X"88",X"FF",X"F7",X"FF",X"F0",X"FE",X"FD",X"F1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E3",
		X"00",X"00",X"88",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CE",X"FF",X"73",X"00",X"00",
		X"88",X"FF",X"FF",X"F3",X"F0",X"FD",X"FD",X"F1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CE",X"FF",X"73",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"E8",X"F1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E9",
		X"00",X"00",X"E0",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CE",X"FF",X"03",X"00",X"00",
		X"00",X"00",X"00",X"80",X"F0",X"FC",X"AD",X"F1",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"F8",
		X"00",X"00",X"E0",X"B4",X"90",X"1E",X"F0",X"30",X"00",X"00",X"00",X"8C",X"FF",X"37",X"00",X"00",
		X"00",X"00",X"80",X"F0",X"F8",X"7F",X"3C",X"E1",X"00",X"00",X"00",X"00",X"00",X"0C",X"E3",X"F8",
		X"00",X"30",X"E1",X"B4",X"96",X"F0",X"F0",X"3C",X"00",X"00",X"00",X"8C",X"FF",X"7F",X"00",X"00",
		X"00",X"00",X"C0",X"F8",X"FF",X"3F",X"1E",X"E1",X"00",X"00",X"00",X"00",X"08",X"CF",X"F3",X"FD",
		X"80",X"3C",X"E1",X"B4",X"96",X"1E",X"F0",X"3C",X"00",X"00",X"00",X"08",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"00",X"C0",X"F0",X"16",X"0F",X"E1",X"00",X"00",X"00",X"08",X"8F",X"FF",X"F5",X"FD",
		X"C0",X"B4",X"E1",X"B4",X"96",X"1E",X"F0",X"3C",X"00",X"00",X"00",X"EE",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"00",X"00",X"70",X"00",X"0F",X"E1",X"00",X"00",X"0C",X"8F",X"FF",X"F3",X"F5",X"FF",
		X"C0",X"3C",X"E1",X"B4",X"96",X"F0",X"F0",X"3C",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E1",X"00",X"00",X"00",X"08",X"F5",X"F0",X"FF",X"FF",
		X"C0",X"B4",X"E1",X"BC",X"9F",X"1F",X"FF",X"3F",X"00",X"00",X"00",X"FF",X"FF",X"7F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"87",X"F9",X"F0",X"FF",X"FE",
		X"CC",X"3C",X"EF",X"BF",X"9F",X"1F",X"FF",X"3F",X"00",X"00",X"88",X"FF",X"FF",X"7F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"0E",X"F7",X"F9",X"F3",X"FF",X"FE",
		X"CC",X"3F",X"EF",X"BF",X"9F",X"FF",X"FF",X"3F",X"00",X"00",X"88",X"FF",X"FF",X"6F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"0E",X"EF",X"F7",X"FB",X"FB",X"FF",X"FE",
		X"CC",X"B7",X"EF",X"BF",X"9F",X"1F",X"FF",X"37",X"00",X"00",X"88",X"FF",X"FF",X"1F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"CE",X"FF",X"FB",X"FF",X"FF",X"FE",
		X"CC",X"3F",X"EF",X"BF",X"9F",X"1F",X"FF",X"B3",X"00",X"00",X"00",X"FF",X"FF",X"53",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"0C",X"EF",X"FF",X"FB",X"FF",X"FF",X"FE",
		X"CC",X"B7",X"EF",X"BF",X"9F",X"FF",X"FF",X"D1",X"00",X"00",X"00",X"F7",X"FF",X"53",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"0E",X"CF",X"FF",X"FF",X"F9",X"FF",X"FC",X"FE",
		X"88",X"3F",X"EF",X"BF",X"9F",X"1F",X"FF",X"E0",X"00",X"00",X"00",X"E8",X"FF",X"53",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"0C",X"CF",X"FD",X"FD",X"FE",X"F0",X"F7",
		X"00",X"33",X"EF",X"BF",X"9F",X"1F",X"77",X"F0",X"00",X"00",X"00",X"CC",X"FF",X"53",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"0C",X"E9",X"FD",X"FE",X"F0",X"F0",
		X"00",X"00",X"EE",X"BF",X"99",X"FF",X"B3",X"F0",X"00",X"00",X"00",X"CC",X"FF",X"43",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"CA",X"FD",X"F4",X"F0",X"F0",
		X"00",X"00",X"EE",X"33",X"00",X"00",X"C0",X"F0",X"00",X"00",X"00",X"88",X"7F",X"30",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"0C",X"CB",X"F2",X"F0",X"F0",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"F0",X"00",X"00",X"00",X"88",X"3F",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"08",X"CF",X"3D",X"F7",X"F0",X"F0",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"FE",X"00",X"00",X"00",X"08",X"C3",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"8F",X"FF",X"FE",X"F7",X"FA",X"F1",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"80",X"78",X"FF",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"F1",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"7E",X"7F",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"0F",X"FA",X"F9",X"FE",X"FD",X"F3",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"E8",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"87",X"F0",X"F9",X"FD",X"F7",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"EE",X"7F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"08",X"C3",X"F3",X"FD",X"F7",X"F7",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"0C",X"F7",X"FB",X"F6",X"F7",
		X"00",X"00",X"00",X"00",X"00",X"88",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"8F",X"FB",X"F5",X"F7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"08",X"CF",X"FF",X"F7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"6E",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"0C",X"ED",X"F7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"4C",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"CE",X"F3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"0C",X"EF",X"FB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"8E",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"6E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
