library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity jng_prg_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of jng_prg_rom is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"AF",X"32",X"81",X"A1",X"C3",X"24",X"14",X"FF",X"85",X"6F",X"D0",X"24",X"C9",X"FF",X"FF",X"FF",
		X"7B",X"C6",X"20",X"5F",X"D0",X"14",X"C9",X"FF",X"87",X"CF",X"5E",X"23",X"56",X"C9",X"FF",X"FF",
		X"7D",X"D6",X"20",X"6F",X"D0",X"25",X"C9",X"FF",X"7B",X"D6",X"20",X"5F",X"D0",X"15",X"C9",X"FF",
		X"E1",X"DF",X"EB",X"E9",X"FF",X"FF",X"FF",X"FF",X"7E",X"FE",X"40",X"C8",X"12",X"23",X"D7",X"18",
		X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AF",X"32",X"81",X"A1",X"32",X"80",X"A0",X"3A",X"2C",X"99",
		X"32",X"30",X"A1",X"3A",X"2D",X"99",X"32",X"40",X"A1",X"21",X"00",X"9C",X"11",X"14",X"80",X"01",
		X"0C",X"00",X"ED",X"B0",X"21",X"10",X"9C",X"11",X"14",X"88",X"01",X"0C",X"00",X"ED",X"B0",X"21",
		X"24",X"9C",X"11",X"34",X"80",X"01",X"08",X"00",X"ED",X"B0",X"21",X"34",X"9C",X"11",X"34",X"88",
		X"01",X"08",X"00",X"ED",X"B0",X"21",X"44",X"9C",X"11",X"34",X"A0",X"01",X"08",X"00",X"ED",X"B0",
		X"CD",X"5E",X"2D",X"CD",X"84",X"2D",X"3A",X"00",X"A0",X"2F",X"32",X"03",X"98",X"3A",X"80",X"A0",
		X"2F",X"32",X"04",X"98",X"3A",X"00",X"A1",X"2F",X"32",X"05",X"98",X"CD",X"C2",X"2F",X"CD",X"0E",
		X"30",X"CD",X"DB",X"2F",X"21",X"E8",X"00",X"E5",X"3A",X"20",X"99",X"F7",X"D4",X"01",X"01",X"04",
		X"D0",X"07",X"35",X"0A",X"D0",X"0C",X"6B",X"0E",X"CD",X"69",X"30",X"CD",X"8D",X"30",X"CD",X"5F",
		X"33",X"21",X"02",X"98",X"34",X"21",X"00",X"98",X"7E",X"A7",X"28",X"01",X"35",X"2A",X"06",X"98",
		X"7C",X"B5",X"28",X"04",X"2B",X"22",X"06",X"98",X"3E",X"01",X"32",X"81",X"A1",X"C9",X"4A",X"55",
		X"4E",X"47",X"4C",X"45",X"52",X"40",X"43",X"52",X"45",X"44",X"49",X"54",X"40",X"4C",X"4F",X"4F",
		X"50",X"20",X"40",X"42",X"4F",X"4D",X"42",X"20",X"54",X"49",X"4D",X"45",X"52",X"20",X"40",X"48",
		X"49",X"20",X"53",X"43",X"4F",X"52",X"45",X"40",X"50",X"55",X"53",X"48",X"20",X"53",X"54",X"41",
		X"52",X"54",X"20",X"42",X"55",X"54",X"54",X"4F",X"4E",X"40",X"4F",X"4E",X"45",X"20",X"50",X"4C",
		X"41",X"59",X"45",X"52",X"20",X"4F",X"4E",X"4C",X"59",X"20",X"20",X"20",X"40",X"4F",X"4E",X"45",
		X"20",X"4F",X"52",X"20",X"54",X"57",X"4F",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"53",X"40",
		X"4F",X"4E",X"45",X"40",X"54",X"57",X"4F",X"40",X"01",X"55",X"50",X"40",X"02",X"55",X"50",X"40",
		X"47",X"41",X"4D",X"45",X"20",X"4F",X"56",X"45",X"52",X"40",X"53",X"43",X"4F",X"52",X"45",X"20",
		X"52",X"41",X"4E",X"4B",X"49",X"4E",X"47",X"40",X"50",X"4C",X"41",X"59",X"45",X"52",X"40",X"45",
		X"4E",X"44",X"40",X"45",X"4E",X"45",X"4D",X"59",X"40",X"50",X"4F",X"49",X"4E",X"54",X"53",X"40",
		X"5C",X"20",X"4B",X"4F",X"4E",X"41",X"4D",X"49",X"20",X"01",X"09",X"08",X"01",X"40",X"50",X"4C",
		X"41",X"59",X"45",X"52",X"20",X"4F",X"4E",X"45",X"40",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",
		X"54",X"57",X"4F",X"40",X"21",X"F0",X"01",X"E5",X"3A",X"21",X"99",X"F7",X"F1",X"01",X"1B",X"02",
		X"27",X"02",X"34",X"02",X"44",X"02",X"56",X"02",X"67",X"02",X"6E",X"02",X"97",X"02",X"F8",X"02",
		X"C9",X"3E",X"01",X"32",X"83",X"A1",X"32",X"2F",X"99",X"CD",X"0A",X"02",X"CD",X"05",X"1B",X"3E",
		X"1E",X"32",X"00",X"98",X"CD",X"1B",X"03",X"C3",X"FC",X"03",X"CD",X"84",X"1A",X"21",X"0E",X"01",
		X"11",X"85",X"81",X"0E",X"BA",X"CD",X"DA",X"16",X"C3",X"48",X"30",X"3A",X"00",X"98",X"A7",X"C0",
		X"CD",X"D1",X"1A",X"C0",X"C3",X"FC",X"03",X"3A",X"23",X"99",X"A7",X"CA",X"FC",X"03",X"3E",X"07",
		X"32",X"21",X"99",X"C9",X"3A",X"23",X"99",X"A7",X"20",X"F4",X"AF",X"32",X"21",X"99",X"3E",X"05",
		X"32",X"20",X"99",X"C9",X"3A",X"23",X"99",X"A7",X"20",X"E4",X"CD",X"B9",X"19",X"D8",X"3E",X"FF",
		X"32",X"00",X"98",X"C3",X"FC",X"03",X"3A",X"23",X"99",X"A7",X"20",X"05",X"3A",X"00",X"98",X"A7",
		X"C0",X"CD",X"1B",X"03",X"C3",X"FC",X"03",X"CD",X"D1",X"1A",X"C0",X"C3",X"FC",X"03",X"3A",X"23",
		X"99",X"A7",X"20",X"0A",X"AF",X"32",X"21",X"99",X"3E",X"04",X"32",X"20",X"99",X"C9",X"3E",X"01",
		X"32",X"83",X"A1",X"32",X"2F",X"99",X"21",X"38",X"01",X"11",X"16",X"85",X"0E",X"A3",X"CD",X"DA",
		X"16",X"CD",X"17",X"0F",X"C3",X"FC",X"03",X"CD",X"75",X"03",X"11",X"15",X"85",X"3A",X"23",X"99",
		X"FE",X"01",X"20",X"05",X"21",X"4A",X"01",X"18",X"03",X"21",X"5D",X"01",X"0E",X"A3",X"CD",X"DA",
		X"16",X"3A",X"04",X"98",X"E6",X"C0",X"C8",X"21",X"23",X"99",X"E6",X"80",X"28",X"0C",X"7E",X"D6",
		X"01",X"27",X"77",X"3E",X"00",X"32",X"10",X"99",X"18",X"13",X"7E",X"FE",X"02",X"D8",X"D6",X"01",
		X"27",X"D6",X"01",X"27",X"77",X"CD",X"4E",X"03",X"3E",X"01",X"32",X"10",X"99",X"AF",X"32",X"11",
		X"99",X"CD",X"27",X"03",X"CD",X"48",X"30",X"CD",X"AD",X"1A",X"CD",X"FB",X"33",X"3E",X"1E",X"32",
		X"00",X"98",X"CD",X"1B",X"03",X"C3",X"FC",X"03",X"3A",X"00",X"98",X"A7",X"C0",X"CD",X"D1",X"1A",
		X"C0",X"21",X"A2",X"88",X"11",X"20",X"00",X"06",X"03",X"36",X"8E",X"19",X"10",X"FB",X"21",X"62",
		X"8B",X"06",X"03",X"36",X"8E",X"19",X"10",X"FB",X"C3",X"F4",X"03",X"3E",X"20",X"32",X"01",X"98",
		X"21",X"00",X"84",X"22",X"52",X"98",X"C9",X"3E",X"03",X"32",X"00",X"9F",X"AF",X"32",X"01",X"9F",
		X"32",X"02",X"9F",X"32",X"0A",X"9F",X"3A",X"34",X"99",X"A7",X"28",X"05",X"3E",X"FF",X"32",X"00",
		X"9F",X"21",X"01",X"9F",X"34",X"CD",X"94",X"03",X"3E",X"0A",X"32",X"03",X"9F",X"C9",X"3E",X"03",
		X"32",X"40",X"9F",X"AF",X"32",X"41",X"9F",X"32",X"42",X"9F",X"32",X"4A",X"9F",X"3A",X"34",X"99",
		X"A7",X"28",X"05",X"3E",X"FF",X"32",X"40",X"9F",X"21",X"41",X"9F",X"34",X"CD",X"AB",X"03",X"3E",
		X"0A",X"32",X"43",X"9F",X"C9",X"21",X"00",X"99",X"06",X"10",X"36",X"00",X"23",X"10",X"FB",X"21",
		X"00",X"9F",X"06",X"10",X"36",X"00",X"23",X"10",X"FB",X"21",X"40",X"9F",X"06",X"10",X"36",X"00",
		X"23",X"10",X"FB",X"C9",X"7E",X"FE",X"19",X"38",X"02",X"3E",X"17",X"21",X"C2",X"03",X"CF",X"7E",
		X"32",X"08",X"9F",X"3E",X"19",X"CF",X"7E",X"32",X"09",X"9F",X"C9",X"7E",X"FE",X"19",X"38",X"02",
		X"3E",X"17",X"21",X"C2",X"03",X"CF",X"7E",X"32",X"48",X"9F",X"3E",X"19",X"CF",X"7E",X"32",X"49",
		X"9F",X"C9",X"00",X"03",X"04",X"05",X"04",X"05",X"06",X"07",X"04",X"07",X"07",X"07",X"05",X"07",
		X"07",X"07",X"05",X"08",X"08",X"08",X"06",X"08",X"08",X"08",X"07",X"00",X"02",X"03",X"04",X"03",
		X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"05",X"05",X"05",X"04",X"06",X"06",X"06",X"04",
		X"07",X"07",X"07",X"04",X"21",X"20",X"99",X"34",X"23",X"36",X"00",X"C9",X"21",X"21",X"99",X"34",
		X"C9",X"21",X"1F",X"04",X"E5",X"3A",X"21",X"99",X"F7",X"20",X"04",X"42",X"04",X"52",X"04",X"8F",
		X"04",X"F3",X"04",X"3F",X"05",X"16",X"06",X"8B",X"06",X"A6",X"06",X"B6",X"06",X"D2",X"06",X"C9",
		X"AF",X"32",X"08",X"98",X"3C",X"32",X"83",X"A1",X"32",X"2F",X"99",X"21",X"00",X"9F",X"7E",X"A7",
		X"28",X"04",X"35",X"C3",X"FC",X"03",X"21",X"0A",X"9F",X"7E",X"36",X"00",X"32",X"04",X"9F",X"C3",
		X"FC",X"03",X"3A",X"01",X"9F",X"32",X"01",X"99",X"CD",X"84",X"32",X"C0",X"CD",X"C3",X"1A",X"C3",
		X"FC",X"03",X"CD",X"B8",X"1A",X"CD",X"0A",X"02",X"CD",X"8F",X"31",X"3A",X"10",X"99",X"A7",X"20",
		X"29",X"21",X"2F",X"01",X"11",X"C2",X"82",X"CD",X"E7",X"30",X"21",X"2F",X"01",X"11",X"C1",X"82",
		X"CD",X"E7",X"30",X"CD",X"DD",X"04",X"21",X"00",X"9F",X"11",X"00",X"99",X"01",X"10",X"00",X"ED",
		X"B0",X"CD",X"06",X"19",X"CD",X"57",X"19",X"C3",X"FC",X"03",X"CD",X"B3",X"31",X"18",X"E4",X"CD",
		X"1D",X"17",X"CD",X"72",X"17",X"CD",X"FB",X"17",X"CD",X"84",X"18",X"3A",X"03",X"99",X"32",X"0F",
		X"99",X"CD",X"B8",X"3F",X"3E",X"78",X"32",X"00",X"98",X"21",X"20",X"1C",X"22",X"06",X"98",X"CD",
		X"65",X"2E",X"CD",X"25",X"2E",X"CD",X"E5",X"2D",X"CD",X"A0",X"2D",X"CD",X"63",X"1F",X"CD",X"BA",
		X"1F",X"CD",X"09",X"20",X"CD",X"58",X"20",X"CD",X"AD",X"23",X"06",X"0A",X"11",X"71",X"85",X"CD",
		X"18",X"05",X"06",X"09",X"11",X"8E",X"85",X"CD",X"13",X"05",X"C3",X"FC",X"03",X"21",X"98",X"01",
		X"11",X"46",X"80",X"0E",X"A3",X"CD",X"DA",X"16",X"21",X"70",X"01",X"11",X"A5",X"80",X"0E",X"A3",
		X"C3",X"DA",X"16",X"3A",X"00",X"98",X"A7",X"20",X"0E",X"06",X"0A",X"11",X"71",X"85",X"CD",X"2E",
		X"05",X"CD",X"BB",X"33",X"C3",X"FC",X"03",X"21",X"BE",X"01",X"11",X"71",X"85",X"01",X"20",X"00",
		X"C3",X"5B",X"06",X"21",X"EC",X"98",X"18",X"03",X"21",X"D4",X"98",X"1A",X"77",X"CB",X"DA",X"23",
		X"1A",X"77",X"23",X"CB",X"9A",X"D7",X"10",X"F3",X"C9",X"21",X"EC",X"98",X"18",X"03",X"21",X"D4",
		X"98",X"7E",X"12",X"CB",X"DA",X"23",X"7E",X"12",X"CB",X"9A",X"23",X"D7",X"10",X"F3",X"C9",X"2A",
		X"06",X"98",X"7D",X"A7",X"CC",X"12",X"07",X"CD",X"47",X"2A",X"CD",X"65",X"2E",X"CD",X"A8",X"28",
		X"CD",X"25",X"2E",X"CD",X"F5",X"26",X"CD",X"E5",X"2D",X"CD",X"DE",X"25",X"CD",X"A0",X"2D",X"CD",
		X"63",X"1F",X"CD",X"BA",X"1F",X"CD",X"09",X"20",X"CD",X"58",X"20",X"CD",X"AD",X"23",X"CD",X"A7",
		X"20",X"CD",X"59",X"1B",X"CD",X"C6",X"1B",X"CD",X"E5",X"1C",X"CD",X"54",X"1E",X"CD",X"3A",X"25",
		X"CD",X"7C",X"21",X"CD",X"E5",X"21",X"CD",X"7D",X"22",X"CD",X"15",X"23",X"CD",X"3C",X"3F",X"CD",
		X"3C",X"3E",X"CD",X"33",X"39",X"CD",X"D4",X"31",X"3A",X"04",X"99",X"A7",X"CA",X"05",X"06",X"FD",
		X"21",X"80",X"98",X"DD",X"21",X"04",X"99",X"DD",X"7E",X"01",X"FD",X"B6",X"01",X"CC",X"6B",X"17",
		X"DD",X"7E",X"02",X"FD",X"B6",X"02",X"CC",X"F4",X"17",X"DD",X"7E",X"03",X"FD",X"B6",X"03",X"CC",
		X"7D",X"18",X"DD",X"7E",X"01",X"DD",X"B6",X"02",X"DD",X"B6",X"03",X"C0",X"FD",X"7E",X"01",X"FD",
		X"B6",X"02",X"FD",X"B6",X"03",X"C0",X"CD",X"C0",X"33",X"CD",X"0A",X"34",X"3E",X"78",X"32",X"00",
		X"98",X"CD",X"1B",X"03",X"3E",X"0A",X"32",X"21",X"99",X"C9",X"CD",X"C0",X"33",X"3E",X"78",X"32",
		X"00",X"98",X"CD",X"1B",X"03",X"3A",X"00",X"99",X"21",X"0A",X"99",X"B6",X"C2",X"FC",X"03",X"CD",
		X"20",X"34",X"C3",X"FC",X"03",X"CD",X"0B",X"06",X"C0",X"18",X"DF",X"21",X"80",X"98",X"7E",X"23",
		X"B6",X"23",X"B6",X"23",X"B6",X"C9",X"3A",X"00",X"98",X"FE",X"01",X"38",X"08",X"28",X"59",X"CD",
		X"4A",X"06",X"C3",X"E2",X"1E",X"CD",X"D1",X"1A",X"C0",X"3A",X"00",X"99",X"21",X"0A",X"99",X"B6",
		X"28",X"15",X"3A",X"10",X"99",X"A7",X"28",X"0C",X"3A",X"40",X"9F",X"21",X"4A",X"9F",X"B6",X"28",
		X"03",X"CD",X"FC",X"03",X"CD",X"FC",X"03",X"C3",X"FC",X"03",X"3A",X"00",X"99",X"21",X"0A",X"99",
		X"B6",X"C0",X"21",X"80",X"01",X"11",X"8E",X"85",X"01",X"20",X"00",X"7E",X"FE",X"40",X"C8",X"D5",
		X"E5",X"CD",X"72",X"2D",X"3A",X"02",X"98",X"0F",X"0F",X"E6",X"07",X"21",X"83",X"06",X"CF",X"7E",
		X"12",X"D1",X"E1",X"13",X"09",X"EB",X"18",X"E3",X"CD",X"05",X"1B",X"11",X"8E",X"85",X"06",X"09",
		X"C3",X"29",X"05",X"87",X"8E",X"95",X"A3",X"87",X"9C",X"95",X"BE",X"3A",X"10",X"99",X"A7",X"20",
		X"0A",X"3E",X"03",X"32",X"20",X"99",X"AF",X"32",X"21",X"99",X"C9",X"3A",X"40",X"9F",X"21",X"4A",
		X"9F",X"B6",X"28",X"ED",X"18",X"10",X"AF",X"32",X"21",X"99",X"21",X"00",X"99",X"11",X"00",X"9F",
		X"01",X"10",X"00",X"ED",X"B0",X"C9",X"3A",X"2E",X"99",X"32",X"83",X"A1",X"32",X"2F",X"99",X"3E",
		X"01",X"32",X"11",X"99",X"21",X"00",X"99",X"11",X"00",X"9F",X"01",X"10",X"00",X"ED",X"B0",X"C3",
		X"F4",X"03",X"3A",X"00",X"98",X"FE",X"01",X"38",X"06",X"CA",X"05",X"1B",X"C3",X"E2",X"1E",X"CD",
		X"D1",X"1A",X"C0",X"3A",X"04",X"99",X"FE",X"09",X"38",X"14",X"3E",X"08",X"32",X"04",X"99",X"21",
		X"0A",X"99",X"34",X"7E",X"FE",X"08",X"38",X"06",X"36",X"00",X"21",X"00",X"99",X"34",X"3E",X"01",
		X"32",X"21",X"99",X"21",X"00",X"99",X"11",X"00",X"9F",X"01",X"10",X"00",X"ED",X"B0",X"CD",X"41",
		X"03",X"C9",X"7C",X"FE",X"10",X"30",X"28",X"E6",X"03",X"20",X"24",X"3A",X"65",X"98",X"FE",X"38",
		X"30",X"05",X"C6",X"08",X"32",X"65",X"98",X"3A",X"68",X"98",X"FE",X"38",X"30",X"05",X"C6",X"08",
		X"32",X"68",X"98",X"3A",X"6B",X"98",X"FE",X"38",X"D0",X"C6",X"08",X"32",X"6B",X"98",X"C9",X"7C",
		X"FE",X"17",X"28",X"10",X"FE",X"13",X"28",X"41",X"FE",X"0B",X"28",X"38",X"FE",X"11",X"C0",X"AF",
		X"32",X"18",X"9C",X"C9",X"CD",X"A5",X"2F",X"E6",X"03",X"32",X"1A",X"98",X"4F",X"3A",X"2F",X"99",
		X"A7",X"28",X"05",X"21",X"BC",X"07",X"18",X"03",X"21",X"C6",X"07",X"7E",X"32",X"08",X"9C",X"23",
		X"7E",X"32",X"19",X"9C",X"23",X"79",X"87",X"CF",X"7E",X"32",X"18",X"9C",X"23",X"7E",X"32",X"09",
		X"9C",X"C3",X"2F",X"34",X"AF",X"32",X"1A",X"9C",X"C9",X"CD",X"A5",X"2F",X"E6",X"03",X"21",X"1A",
		X"98",X"BE",X"28",X"F5",X"4F",X"3A",X"2F",X"99",X"A7",X"28",X"05",X"21",X"BC",X"07",X"18",X"03",
		X"21",X"C6",X"07",X"7E",X"32",X"0A",X"9C",X"23",X"7E",X"32",X"1B",X"9C",X"23",X"79",X"87",X"CF",
		X"7E",X"32",X"1A",X"9C",X"23",X"7E",X"32",X"0B",X"9C",X"C3",X"2F",X"34",X"7C",X"0F",X"94",X"8C",
		X"94",X"BC",X"5C",X"BC",X"5C",X"8C",X"7F",X"0F",X"5C",X"84",X"5C",X"54",X"94",X"54",X"94",X"84",
		X"21",X"EE",X"07",X"E5",X"3A",X"21",X"99",X"F7",X"EF",X"07",X"06",X"08",X"16",X"08",X"39",X"08",
		X"96",X"08",X"B6",X"08",X"82",X"09",X"B1",X"09",X"C4",X"09",X"D4",X"09",X"F5",X"09",X"C9",X"21",
		X"40",X"9F",X"7E",X"A7",X"28",X"04",X"35",X"C3",X"FC",X"03",X"21",X"4A",X"9F",X"7E",X"36",X"00",
		X"32",X"44",X"9F",X"C3",X"FC",X"03",X"3A",X"41",X"9F",X"32",X"01",X"99",X"CD",X"84",X"32",X"C0",
		X"CD",X"C3",X"1A",X"C3",X"FC",X"03",X"CD",X"B8",X"1A",X"CD",X"0A",X"02",X"CD",X"8F",X"31",X"CD",
		X"B3",X"31",X"CD",X"87",X"08",X"21",X"40",X"9F",X"11",X"00",X"99",X"01",X"10",X"00",X"ED",X"B0",
		X"CD",X"06",X"19",X"CD",X"57",X"19",X"C3",X"FC",X"03",X"CD",X"1D",X"17",X"CD",X"72",X"17",X"CD",
		X"FB",X"17",X"CD",X"84",X"18",X"3A",X"03",X"99",X"32",X"0F",X"99",X"CD",X"B8",X"3F",X"3E",X"78",
		X"32",X"00",X"98",X"21",X"20",X"1C",X"22",X"06",X"98",X"CD",X"65",X"2E",X"CD",X"25",X"2E",X"CD",
		X"E5",X"2D",X"CD",X"A0",X"2D",X"CD",X"63",X"1F",X"CD",X"BA",X"1F",X"CD",X"09",X"20",X"CD",X"58",
		X"20",X"CD",X"AD",X"23",X"06",X"0A",X"11",X"71",X"85",X"CD",X"18",X"05",X"06",X"09",X"11",X"8E",
		X"85",X"CD",X"13",X"05",X"C3",X"FC",X"03",X"21",X"98",X"01",X"11",X"46",X"80",X"FF",X"21",X"74",
		X"01",X"11",X"A5",X"80",X"FF",X"C9",X"3A",X"00",X"98",X"A7",X"20",X"0E",X"06",X"0A",X"11",X"71",
		X"85",X"CD",X"2E",X"05",X"CD",X"BB",X"33",X"C3",X"FC",X"03",X"21",X"C9",X"01",X"11",X"71",X"85",
		X"01",X"20",X"00",X"C3",X"5B",X"06",X"2A",X"06",X"98",X"7D",X"A7",X"CC",X"12",X"07",X"CD",X"47",
		X"2A",X"CD",X"65",X"2E",X"CD",X"A8",X"28",X"CD",X"25",X"2E",X"CD",X"F5",X"26",X"CD",X"E5",X"2D",
		X"CD",X"DE",X"25",X"CD",X"A0",X"2D",X"CD",X"63",X"1F",X"CD",X"BA",X"1F",X"CD",X"09",X"20",X"CD",
		X"58",X"20",X"CD",X"AD",X"23",X"CD",X"A7",X"20",X"CD",X"59",X"1B",X"CD",X"C6",X"1B",X"CD",X"E5",
		X"1C",X"CD",X"54",X"1E",X"CD",X"3A",X"25",X"CD",X"7C",X"21",X"CD",X"E5",X"21",X"CD",X"7D",X"22",
		X"CD",X"15",X"23",X"CD",X"3C",X"3F",X"CD",X"3C",X"3E",X"CD",X"33",X"39",X"CD",X"D4",X"31",X"3A",
		X"04",X"99",X"A7",X"CA",X"7C",X"09",X"FD",X"21",X"80",X"98",X"DD",X"21",X"04",X"99",X"DD",X"7E",
		X"01",X"FD",X"B6",X"01",X"CC",X"6B",X"17",X"DD",X"7E",X"02",X"FD",X"B6",X"02",X"CC",X"F4",X"17",
		X"DD",X"7E",X"03",X"FD",X"B6",X"03",X"CC",X"7D",X"18",X"DD",X"7E",X"01",X"DD",X"B6",X"02",X"DD",
		X"B6",X"03",X"C0",X"FD",X"7E",X"01",X"FD",X"B6",X"02",X"FD",X"B6",X"03",X"C0",X"CD",X"C0",X"33",
		X"CD",X"0A",X"34",X"3E",X"78",X"32",X"00",X"98",X"CD",X"1B",X"03",X"3E",X"0A",X"32",X"21",X"99",
		X"C9",X"CD",X"C0",X"33",X"3E",X"78",X"32",X"00",X"98",X"CD",X"1B",X"03",X"3A",X"00",X"99",X"21",
		X"0A",X"99",X"B6",X"C2",X"FC",X"03",X"CD",X"20",X"34",X"C3",X"FC",X"03",X"CD",X"0B",X"06",X"C0",
		X"18",X"DF",X"3A",X"00",X"98",X"FE",X"01",X"38",X"09",X"CA",X"78",X"06",X"CD",X"4A",X"06",X"C3",
		X"E2",X"1E",X"CD",X"D1",X"1A",X"C0",X"3A",X"00",X"99",X"21",X"0A",X"99",X"B6",X"28",X"0F",X"3A",
		X"00",X"9F",X"21",X"0A",X"9F",X"B6",X"28",X"03",X"CD",X"FC",X"03",X"CD",X"FC",X"03",X"C3",X"FC",
		X"03",X"3A",X"00",X"9F",X"21",X"0A",X"9F",X"B6",X"20",X"1A",X"3E",X"03",X"32",X"20",X"99",X"AF",
		X"32",X"21",X"99",X"C9",X"AF",X"32",X"21",X"99",X"21",X"00",X"99",X"11",X"40",X"9F",X"01",X"10",
		X"00",X"ED",X"B0",X"C9",X"3E",X"01",X"32",X"83",X"A1",X"32",X"2F",X"99",X"3E",X"00",X"32",X"11",
		X"99",X"21",X"00",X"99",X"11",X"40",X"9F",X"01",X"10",X"00",X"ED",X"B0",X"AF",X"32",X"21",X"99",
		X"3C",X"32",X"20",X"99",X"C9",X"3A",X"00",X"98",X"FE",X"01",X"38",X"06",X"CA",X"05",X"1B",X"C3",
		X"E2",X"1E",X"CD",X"D1",X"1A",X"C0",X"3A",X"04",X"99",X"FE",X"09",X"38",X"14",X"3E",X"08",X"32",
		X"04",X"99",X"21",X"0A",X"99",X"34",X"7E",X"FE",X"08",X"38",X"06",X"36",X"00",X"21",X"00",X"99",
		X"34",X"3E",X"01",X"32",X"21",X"99",X"21",X"00",X"99",X"11",X"40",X"9F",X"01",X"10",X"00",X"ED",
		X"B0",X"CD",X"68",X"03",X"C9",X"21",X"57",X"0A",X"E5",X"3A",X"21",X"99",X"F7",X"77",X"0A",X"29",
		X"0B",X"2F",X"0B",X"79",X"0B",X"45",X"0C",X"70",X"0C",X"91",X"0C",X"AA",X"0C",X"AD",X"0C",X"B0",
		X"0C",X"B3",X"0C",X"B6",X"0C",X"BF",X"0C",X"3A",X"23",X"99",X"A7",X"C8",X"4F",X"3A",X"04",X"98",
		X"E6",X"C0",X"C8",X"E6",X"80",X"28",X"0A",X"AF",X"32",X"20",X"99",X"3E",X"05",X"32",X"21",X"99",
		X"C9",X"79",X"FE",X"02",X"D8",X"18",X"F0",X"AF",X"32",X"11",X"99",X"FD",X"21",X"12",X"99",X"DD",
		X"21",X"40",X"98",X"DD",X"36",X"00",X"00",X"21",X"42",X"99",X"06",X"0A",X"E5",X"22",X"52",X"98",
		X"FD",X"7E",X"02",X"BE",X"38",X"48",X"28",X"02",X"18",X"12",X"FD",X"7E",X"01",X"2B",X"BE",X"38",
		X"3D",X"28",X"02",X"18",X"07",X"FD",X"7E",X"00",X"2B",X"BE",X"38",X"32",X"E1",X"2B",X"2B",X"E5",
		X"05",X"78",X"32",X"47",X"98",X"28",X"0F",X"87",X"87",X"87",X"87",X"4F",X"06",X"00",X"21",X"CF",
		X"99",X"11",X"DF",X"99",X"ED",X"B8",X"E1",X"FD",X"7E",X"00",X"77",X"23",X"FD",X"7E",X"01",X"77",
		X"23",X"FD",X"7E",X"02",X"77",X"06",X"0C",X"23",X"36",X"5B",X"10",X"FB",X"18",X"1C",X"DD",X"34",
		X"00",X"E1",X"11",X"10",X"00",X"19",X"10",X"A4",X"CD",X"FC",X"03",X"CD",X"FC",X"03",X"CD",X"FC",
		X"03",X"CD",X"FC",X"03",X"CD",X"FC",X"03",X"C3",X"FC",X"03",X"AF",X"32",X"41",X"98",X"32",X"42",
		X"98",X"21",X"E0",X"99",X"06",X"0C",X"36",X"5B",X"23",X"10",X"FB",X"3A",X"21",X"99",X"FE",X"06",
		X"30",X"0B",X"3E",X"01",X"32",X"83",X"A1",X"32",X"2F",X"99",X"C3",X"FC",X"03",X"3A",X"2E",X"99",
		X"32",X"83",X"A1",X"32",X"2F",X"99",X"C3",X"FC",X"03",X"CD",X"88",X"19",X"C3",X"FC",X"03",X"CD",
		X"B9",X"19",X"D8",X"CD",X"23",X"0C",X"CD",X"5B",X"1A",X"3A",X"47",X"98",X"87",X"21",X"98",X"01",
		X"11",X"06",X"8D",X"83",X"5F",X"0E",X"87",X"CD",X"F2",X"30",X"3A",X"42",X"98",X"06",X"95",X"CD",
		X"5F",X"0C",X"3A",X"41",X"98",X"0E",X"95",X"CD",X"54",X"0C",X"3A",X"21",X"99",X"FE",X"06",X"30",
		X"0C",X"CD",X"DD",X"04",X"21",X"08",X"07",X"22",X"06",X"98",X"C3",X"FC",X"03",X"CD",X"DD",X"04",
		X"21",X"08",X"07",X"22",X"06",X"98",X"C3",X"FC",X"03",X"3A",X"02",X"98",X"E6",X"07",X"C0",X"2A",
		X"06",X"98",X"7C",X"B5",X"CA",X"32",X"0C",X"CD",X"06",X"2D",X"28",X"5F",X"3A",X"16",X"98",X"CB",
		X"47",X"28",X"2E",X"21",X"42",X"98",X"CB",X"4F",X"7E",X"32",X"43",X"98",X"28",X"0A",X"34",X"7E",
		X"FE",X"1B",X"38",X"0B",X"36",X"00",X"18",X"07",X"7E",X"A7",X"20",X"02",X"36",X"1B",X"35",X"3A",
		X"43",X"98",X"06",X"8E",X"CD",X"5F",X"0C",X"3A",X"42",X"98",X"06",X"95",X"CD",X"5F",X"0C",X"18",
		X"2A",X"21",X"41",X"98",X"CB",X"4F",X"7E",X"32",X"44",X"98",X"28",X"0A",X"34",X"7E",X"FE",X"0C",
		X"38",X"09",X"36",X"0B",X"18",X"05",X"7E",X"A7",X"28",X"01",X"35",X"3A",X"44",X"98",X"0E",X"8E",
		X"CD",X"54",X"0C",X"3A",X"41",X"98",X"0E",X"95",X"CD",X"54",X"0C",X"CD",X"AB",X"1B",X"20",X"33",
		X"3A",X"42",X"98",X"FE",X"1A",X"28",X"3B",X"21",X"E0",X"99",X"3A",X"41",X"98",X"CF",X"3A",X"42",
		X"98",X"C6",X"41",X"77",X"21",X"41",X"98",X"7E",X"32",X"44",X"98",X"34",X"7E",X"FE",X"0C",X"38",
		X"02",X"36",X"0B",X"3A",X"44",X"98",X"0E",X"8E",X"CD",X"54",X"0C",X"3A",X"41",X"98",X"0E",X"95",
		X"CD",X"54",X"0C",X"21",X"E0",X"99",X"11",X"E4",X"85",X"06",X"0C",X"7E",X"12",X"23",X"D7",X"10",
		X"FA",X"C9",X"ED",X"5B",X"52",X"98",X"13",X"21",X"E0",X"99",X"01",X"0C",X"00",X"ED",X"B0",X"CD",
		X"88",X"19",X"C3",X"FC",X"03",X"CD",X"B9",X"19",X"D8",X"3E",X"1E",X"32",X"00",X"98",X"CD",X"1B",
		X"03",X"C3",X"FC",X"03",X"11",X"C4",X"8D",X"3C",X"47",X"D7",X"10",X"FD",X"79",X"12",X"C9",X"21",
		X"61",X"8F",X"4F",X"3E",X"1A",X"91",X"CF",X"70",X"EB",X"D7",X"78",X"12",X"D7",X"78",X"12",X"C9",
		X"3A",X"00",X"98",X"A7",X"C0",X"CD",X"D1",X"1A",X"C0",X"3A",X"10",X"99",X"A7",X"C2",X"FC",X"03",
		X"AF",X"32",X"20",X"99",X"3C",X"32",X"83",X"A1",X"32",X"2F",X"99",X"3E",X"03",X"32",X"21",X"99",
		X"C9",X"3E",X"01",X"32",X"11",X"99",X"FD",X"21",X"17",X"99",X"DD",X"21",X"40",X"98",X"DD",X"36",
		X"00",X"00",X"21",X"42",X"99",X"06",X"0A",X"C3",X"8C",X"0A",X"C3",X"29",X"0B",X"C3",X"2F",X"0B",
		X"C3",X"79",X"0B",X"C3",X"45",X"0C",X"3A",X"00",X"98",X"A7",X"C0",X"CD",X"D1",X"1A",X"C0",X"AF",
		X"32",X"20",X"99",X"3C",X"32",X"83",X"A1",X"32",X"2F",X"99",X"3E",X"03",X"32",X"21",X"99",X"C9",
		X"21",X"EA",X"0C",X"E5",X"3A",X"21",X"99",X"F7",X"F7",X"0C",X"07",X"0D",X"17",X"0D",X"31",X"0D",
		X"6F",X"0D",X"77",X"0D",X"21",X"0E",X"2C",X"0E",X"50",X"0E",X"3A",X"23",X"99",X"A7",X"C8",X"AF",
		X"32",X"20",X"99",X"32",X"21",X"99",X"C9",X"AF",X"32",X"10",X"99",X"32",X"11",X"99",X"CD",X"75",
		X"03",X"CD",X"27",X"03",X"C3",X"FC",X"03",X"3A",X"01",X"9F",X"32",X"01",X"99",X"CD",X"84",X"32",
		X"C0",X"CD",X"C3",X"1A",X"C3",X"FC",X"03",X"CD",X"B8",X"1A",X"CD",X"0A",X"02",X"CD",X"DD",X"04",
		X"21",X"00",X"9F",X"11",X"00",X"99",X"01",X"10",X"00",X"ED",X"B0",X"CD",X"06",X"19",X"C3",X"FC",
		X"03",X"CD",X"1D",X"17",X"CD",X"72",X"17",X"CD",X"FB",X"17",X"CD",X"84",X"18",X"3A",X"03",X"99",
		X"32",X"0F",X"99",X"CD",X"B8",X"3F",X"3E",X"3C",X"32",X"00",X"98",X"21",X"20",X"1C",X"22",X"06",
		X"98",X"CD",X"65",X"2E",X"CD",X"25",X"2E",X"CD",X"E5",X"2D",X"CD",X"A0",X"2D",X"CD",X"63",X"1F",
		X"CD",X"BA",X"1F",X"CD",X"09",X"20",X"CD",X"58",X"20",X"CD",X"AD",X"23",X"C3",X"FC",X"03",X"3A",
		X"00",X"98",X"A7",X"C0",X"C3",X"FC",X"03",X"2A",X"06",X"98",X"7D",X"A7",X"CC",X"12",X"07",X"CD",
		X"B0",X"3E",X"CD",X"47",X"2A",X"CD",X"65",X"2E",X"CD",X"A8",X"28",X"CD",X"25",X"2E",X"CD",X"F5",
		X"26",X"CD",X"E5",X"2D",X"CD",X"E6",X"2B",X"CD",X"A0",X"2D",X"CD",X"63",X"1F",X"CD",X"BA",X"1F",
		X"CD",X"09",X"20",X"CD",X"58",X"20",X"CD",X"AD",X"23",X"CD",X"A7",X"20",X"CD",X"A3",X"1C",X"CD",
		X"C6",X"1B",X"CD",X"E5",X"1C",X"CD",X"54",X"1E",X"CD",X"3A",X"25",X"CD",X"7C",X"21",X"CD",X"E5",
		X"21",X"CD",X"7D",X"22",X"CD",X"15",X"23",X"CD",X"3C",X"3F",X"CD",X"3C",X"3E",X"CD",X"D4",X"31",
		X"3A",X"04",X"99",X"A7",X"28",X"3A",X"FD",X"21",X"80",X"98",X"DD",X"21",X"04",X"99",X"DD",X"7E",
		X"01",X"FD",X"B6",X"01",X"CC",X"6B",X"17",X"DD",X"7E",X"02",X"FD",X"B6",X"02",X"CC",X"F4",X"17",
		X"DD",X"7E",X"03",X"FD",X"B6",X"03",X"CC",X"7D",X"18",X"DD",X"7E",X"01",X"DD",X"B6",X"02",X"DD",
		X"B6",X"03",X"C0",X"FD",X"7E",X"01",X"FD",X"B6",X"02",X"FD",X"B6",X"03",X"C0",X"C3",X"FC",X"03",
		X"CD",X"0B",X"06",X"C0",X"3E",X"08",X"32",X"21",X"99",X"3E",X"78",X"32",X"00",X"98",X"C3",X"1B",
		X"03",X"3E",X"78",X"32",X"00",X"98",X"CD",X"1B",X"03",X"C3",X"FC",X"03",X"3A",X"00",X"98",X"FE",
		X"01",X"38",X"06",X"CA",X"05",X"1B",X"C3",X"E2",X"1E",X"CD",X"D1",X"1A",X"C0",X"21",X"00",X"99",
		X"11",X"00",X"9F",X"01",X"10",X"00",X"ED",X"B0",X"3E",X"01",X"32",X"21",X"99",X"C3",X"41",X"03",
		X"3A",X"00",X"98",X"FE",X"01",X"38",X"06",X"CA",X"05",X"1B",X"C3",X"E2",X"1E",X"CD",X"D1",X"1A",
		X"C0",X"AF",X"32",X"20",X"99",X"3E",X"03",X"32",X"21",X"99",X"C9",X"21",X"95",X"0E",X"E5",X"3A",
		X"21",X"99",X"F7",X"A2",X"0E",X"A5",X"0E",X"22",X"0F",X"84",X"0F",X"AE",X"0F",X"E1",X"0F",X"44",
		X"10",X"60",X"10",X"6E",X"10",X"B4",X"10",X"D8",X"10",X"E0",X"10",X"36",X"11",X"52",X"11",X"66",
		X"11",X"F3",X"11",X"FE",X"11",X"3A",X"23",X"99",X"A7",X"C8",X"AF",X"32",X"20",X"99",X"32",X"21",
		X"99",X"C9",X"C3",X"FC",X"03",X"21",X"23",X"01",X"11",X"B0",X"84",X"0E",X"A3",X"CD",X"F2",X"30",
		X"21",X"23",X"01",X"11",X"AA",X"84",X"0E",X"A3",X"CD",X"F2",X"30",X"21",X"98",X"01",X"11",X"7A",
		X"86",X"0E",X"BA",X"CD",X"DA",X"16",X"21",X"A3",X"01",X"11",X"1A",X"85",X"0E",X"8E",X"CD",X"DA",
		X"16",X"21",X"A9",X"01",X"11",X"B0",X"84",X"FF",X"21",X"A9",X"01",X"11",X"AA",X"84",X"FF",X"CD",
		X"17",X"0F",X"DD",X"21",X"A0",X"13",X"21",X"78",X"86",X"CD",X"13",X"12",X"DD",X"21",X"A0",X"13",
		X"21",X"76",X"86",X"CD",X"13",X"12",X"DD",X"21",X"A0",X"13",X"21",X"74",X"86",X"CD",X"13",X"12",
		X"DD",X"21",X"8F",X"13",X"21",X"6E",X"86",X"CD",X"13",X"12",X"DD",X"21",X"A0",X"13",X"21",X"68",
		X"86",X"CD",X"13",X"12",X"C3",X"FC",X"03",X"21",X"B0",X"01",X"11",X"42",X"85",X"0E",X"BA",X"C3",
		X"DA",X"16",X"DD",X"21",X"CB",X"13",X"21",X"98",X"85",X"CD",X"18",X"12",X"DD",X"21",X"BE",X"13",
		X"21",X"96",X"85",X"CD",X"18",X"12",X"DD",X"21",X"AD",X"13",X"21",X"94",X"85",X"CD",X"18",X"12",
		X"DD",X"21",X"D4",X"13",X"21",X"8E",X"85",X"CD",X"18",X"12",X"DD",X"21",X"AD",X"13",X"21",X"88",
		X"85",X"CD",X"18",X"12",X"3E",X"0A",X"32",X"F4",X"85",X"3C",X"32",X"14",X"86",X"3C",X"32",X"F6",
		X"85",X"3C",X"32",X"16",X"86",X"3C",X"32",X"F8",X"85",X"3C",X"32",X"18",X"86",X"3E",X"BA",X"32",
		X"F4",X"8D",X"32",X"14",X"8E",X"32",X"F6",X"8D",X"32",X"16",X"8E",X"32",X"F8",X"8D",X"32",X"18",
		X"8E",X"C3",X"FC",X"03",X"AF",X"32",X"10",X"99",X"32",X"11",X"99",X"CD",X"75",X"03",X"CD",X"27",
		X"03",X"CD",X"B8",X"1A",X"CD",X"C3",X"1A",X"21",X"00",X"9F",X"11",X"00",X"99",X"01",X"10",X"00",
		X"ED",X"B0",X"AF",X"32",X"45",X"98",X"3E",X"3C",X"32",X"00",X"98",X"C3",X"FC",X"03",X"3A",X"00",
		X"98",X"A7",X"C0",X"3A",X"45",X"98",X"21",X"57",X"12",X"87",X"4F",X"87",X"81",X"CF",X"7E",X"23",
		X"5E",X"23",X"56",X"23",X"E5",X"EB",X"CD",X"E3",X"16",X"E1",X"7E",X"32",X"46",X"98",X"23",X"5E",
		X"23",X"56",X"EB",X"CD",X"00",X"17",X"3E",X"20",X"32",X"62",X"98",X"32",X"65",X"98",X"C3",X"FC",
		X"03",X"CD",X"89",X"3F",X"CD",X"E5",X"2D",X"CD",X"C9",X"3E",X"CD",X"A0",X"2D",X"CD",X"63",X"1F",
		X"CD",X"BA",X"1F",X"CD",X"AD",X"23",X"CD",X"A7",X"20",X"CD",X"E5",X"1C",X"CD",X"3A",X"25",X"CD",
		X"7C",X"21",X"CD",X"E5",X"21",X"FD",X"21",X"80",X"98",X"DD",X"21",X"04",X"99",X"DD",X"7E",X"00",
		X"A7",X"28",X"16",X"DD",X"7E",X"01",X"FD",X"B6",X"01",X"C0",X"ED",X"5B",X"02",X"9B",X"3E",X"77",
		X"CD",X"72",X"2D",X"3E",X"AB",X"12",X"C3",X"FC",X"03",X"FD",X"7E",X"00",X"A7",X"C0",X"3E",X"4A",
		X"ED",X"5B",X"42",X"9B",X"CB",X"DA",X"12",X"CB",X"9A",X"3E",X"76",X"CD",X"72",X"2D",X"3E",X"4A",
		X"12",X"C3",X"FC",X"03",X"21",X"45",X"98",X"34",X"7E",X"FE",X"03",X"30",X"0B",X"3E",X"04",X"32",
		X"21",X"99",X"3E",X"3C",X"32",X"00",X"98",X"C9",X"3E",X"3C",X"32",X"00",X"98",X"C3",X"FC",X"03",
		X"3A",X"00",X"98",X"A7",X"C0",X"CD",X"FC",X"03",X"AF",X"32",X"12",X"9C",X"18",X"18",X"3A",X"00",
		X"98",X"A7",X"C0",X"AF",X"32",X"10",X"9C",X"32",X"12",X"9C",X"21",X"00",X"9B",X"CD",X"47",X"1B",
		X"21",X"40",X"9B",X"CD",X"47",X"1B",X"3A",X"45",X"98",X"21",X"57",X"12",X"87",X"4F",X"87",X"81",
		X"CF",X"7E",X"23",X"5E",X"23",X"56",X"23",X"E5",X"EB",X"CD",X"E3",X"16",X"E1",X"7E",X"32",X"46",
		X"98",X"23",X"5E",X"23",X"56",X"EB",X"CD",X"00",X"17",X"3E",X"20",X"32",X"62",X"98",X"32",X"65",
		X"98",X"C3",X"FC",X"03",X"21",X"70",X"85",X"11",X"20",X"00",X"06",X"04",X"36",X"20",X"19",X"10",
		X"FB",X"CD",X"E5",X"2D",X"CD",X"A0",X"2D",X"CD",X"BA",X"1F",X"CD",X"63",X"1F",X"CD",X"AD",X"23",
		X"3E",X"3C",X"32",X"00",X"98",X"C3",X"FC",X"03",X"3A",X"00",X"98",X"A7",X"C0",X"C3",X"FC",X"03",
		X"CD",X"89",X"3F",X"CD",X"E5",X"2D",X"CD",X"C9",X"3E",X"CD",X"A0",X"2D",X"CD",X"63",X"1F",X"CD",
		X"BA",X"1F",X"CD",X"AD",X"23",X"CD",X"A7",X"20",X"CD",X"E5",X"1C",X"CD",X"3A",X"25",X"CD",X"7C",
		X"21",X"CD",X"E5",X"21",X"FD",X"21",X"80",X"98",X"DD",X"21",X"04",X"99",X"DD",X"7E",X"00",X"FD",
		X"B6",X"00",X"CA",X"FC",X"03",X"DD",X"7E",X"01",X"FD",X"B6",X"01",X"CA",X"FC",X"03",X"3A",X"46",
		X"98",X"21",X"68",X"21",X"DF",X"7B",X"32",X"42",X"98",X"7A",X"11",X"70",X"85",X"CD",X"B1",X"30",
		X"3A",X"42",X"98",X"C3",X"B6",X"30",X"21",X"45",X"98",X"34",X"7E",X"FE",X"0B",X"30",X"0B",X"3E",
		X"08",X"32",X"21",X"99",X"3E",X"3C",X"32",X"00",X"98",X"C9",X"3E",X"3C",X"32",X"00",X"98",X"C3",
		X"FC",X"03",X"3A",X"00",X"98",X"A7",X"C0",X"ED",X"5B",X"02",X"9B",X"3E",X"77",X"CD",X"72",X"2D",
		X"3E",X"AB",X"12",X"C3",X"AE",X"0F",X"AF",X"32",X"62",X"98",X"32",X"65",X"98",X"CD",X"C1",X"11",
		X"3A",X"05",X"99",X"A7",X"28",X"0F",X"3A",X"02",X"98",X"E6",X"3F",X"20",X"08",X"3E",X"FF",X"32",
		X"70",X"98",X"CD",X"E5",X"11",X"CD",X"E5",X"2D",X"CD",X"A0",X"2D",X"CD",X"63",X"1F",X"CD",X"BA",
		X"1F",X"CD",X"AD",X"23",X"CD",X"A3",X"1C",X"CD",X"E5",X"1C",X"CD",X"3A",X"25",X"CD",X"7C",X"21",
		X"CD",X"E5",X"21",X"FD",X"21",X"80",X"98",X"DD",X"21",X"04",X"99",X"DD",X"7E",X"01",X"FD",X"B6",
		X"01",X"C0",X"ED",X"5B",X"02",X"9B",X"3E",X"77",X"CD",X"72",X"2D",X"3E",X"AB",X"12",X"C3",X"FC",
		X"03",X"3A",X"47",X"98",X"A7",X"C8",X"AF",X"32",X"47",X"98",X"3A",X"05",X"99",X"A7",X"28",X"08",
		X"11",X"AA",X"85",X"3E",X"60",X"C3",X"B6",X"30",X"3E",X"05",X"11",X"6A",X"85",X"CD",X"B1",X"30",
		X"3E",X"00",X"C3",X"B6",X"30",X"21",X"6A",X"85",X"11",X"20",X"00",X"06",X"04",X"36",X"20",X"19",
		X"10",X"FB",X"C9",X"3E",X"3C",X"32",X"00",X"98",X"CD",X"1B",X"03",X"C3",X"FC",X"03",X"3A",X"00",
		X"98",X"A7",X"C0",X"CD",X"D1",X"1A",X"C0",X"CD",X"88",X"19",X"32",X"20",X"99",X"3E",X"04",X"32",
		X"21",X"99",X"C9",X"11",X"20",X"00",X"18",X"03",X"11",X"E0",X"FF",X"DD",X"46",X"00",X"DD",X"23",
		X"DD",X"7E",X"00",X"77",X"DD",X"23",X"DD",X"7E",X"00",X"CB",X"DC",X"77",X"CB",X"9C",X"19",X"10",
		X"01",X"C9",X"05",X"28",X"13",X"DD",X"23",X"DD",X"7E",X"00",X"77",X"DD",X"23",X"DD",X"7E",X"00",
		X"CB",X"DC",X"77",X"CB",X"9C",X"19",X"10",X"ED",X"DD",X"23",X"DD",X"7E",X"00",X"77",X"DD",X"23",
		X"DD",X"7E",X"00",X"CB",X"DC",X"77",X"C9",X"06",X"9F",X"12",X"04",X"17",X"13",X"06",X"B7",X"12",
		X"06",X"2F",X"13",X"06",X"CF",X"12",X"08",X"47",X"13",X"08",X"E7",X"12",X"08",X"5F",X"13",X"08",
		X"E7",X"12",X"07",X"5F",X"13",X"08",X"E7",X"12",X"06",X"5F",X"13",X"08",X"E7",X"12",X"05",X"5F",
		X"13",X"08",X"E7",X"12",X"04",X"5F",X"13",X"08",X"E7",X"12",X"03",X"5F",X"13",X"08",X"E7",X"12",
		X"02",X"5F",X"13",X"08",X"E7",X"12",X"01",X"5F",X"13",X"06",X"FF",X"12",X"08",X"77",X"13",X"58",
		X"86",X"78",X"86",X"98",X"86",X"B8",X"86",X"D8",X"86",X"F8",X"86",X"18",X"87",X"38",X"87",X"58",
		X"87",X"78",X"87",X"98",X"87",X"B8",X"87",X"56",X"86",X"76",X"86",X"96",X"86",X"B6",X"86",X"D6",
		X"86",X"F6",X"86",X"16",X"87",X"36",X"87",X"56",X"87",X"76",X"87",X"96",X"87",X"B6",X"87",X"54",
		X"86",X"74",X"86",X"94",X"86",X"B4",X"86",X"D4",X"86",X"F4",X"86",X"14",X"87",X"34",X"87",X"54",
		X"87",X"74",X"87",X"94",X"87",X"B4",X"87",X"4E",X"86",X"6E",X"86",X"8E",X"86",X"AE",X"86",X"CE",
		X"86",X"EE",X"86",X"0E",X"87",X"2E",X"87",X"4E",X"87",X"6E",X"87",X"8E",X"87",X"AE",X"87",X"48",
		X"86",X"68",X"86",X"88",X"86",X"A8",X"86",X"C8",X"86",X"E8",X"86",X"08",X"87",X"28",X"87",X"48",
		X"87",X"68",X"87",X"88",X"87",X"A8",X"87",X"B8",X"85",X"98",X"85",X"78",X"85",X"58",X"85",X"38",
		X"85",X"18",X"85",X"F8",X"84",X"D8",X"84",X"B8",X"84",X"98",X"84",X"78",X"84",X"58",X"84",X"B6",
		X"85",X"96",X"85",X"76",X"85",X"56",X"85",X"36",X"85",X"16",X"85",X"F6",X"84",X"D6",X"84",X"B6",
		X"84",X"96",X"84",X"76",X"84",X"56",X"84",X"B4",X"85",X"94",X"85",X"74",X"85",X"54",X"85",X"34",
		X"85",X"14",X"85",X"F4",X"84",X"D4",X"84",X"B4",X"84",X"94",X"84",X"74",X"84",X"54",X"84",X"AE",
		X"85",X"8E",X"85",X"6E",X"85",X"4E",X"85",X"2E",X"85",X"0E",X"85",X"EE",X"84",X"CE",X"84",X"AE",
		X"84",X"8E",X"84",X"6E",X"84",X"5E",X"84",X"A8",X"85",X"88",X"85",X"68",X"85",X"48",X"85",X"28",
		X"85",X"08",X"85",X"E8",X"84",X"C8",X"84",X"A8",X"84",X"88",X"84",X"68",X"84",X"58",X"84",X"08",
		X"77",X"AB",X"80",X"B0",X"80",X"B0",X"80",X"B0",X"80",X"B0",X"80",X"B0",X"A0",X"B0",X"C0",X"6A",
		X"06",X"77",X"AB",X"80",X"B0",X"80",X"B0",X"80",X"B0",X"80",X"B0",X"C0",X"6A",X"08",X"76",X"4A",
		X"80",X"88",X"80",X"88",X"80",X"88",X"80",X"88",X"80",X"88",X"A0",X"88",X"C0",X"88",X"06",X"76",
		X"56",X"80",X"98",X"80",X"98",X"80",X"98",X"80",X"98",X"C0",X"98",X"04",X"76",X"4F",X"80",X"90",
		X"80",X"90",X"C0",X"90",X"08",X"76",X"56",X"80",X"98",X"80",X"98",X"80",X"98",X"80",X"98",X"80",
		X"98",X"A0",X"98",X"C0",X"98",X"07",X"76",X"4F",X"80",X"90",X"80",X"90",X"80",X"90",X"80",X"90",
		X"A0",X"90",X"C0",X"90",X"06",X"76",X"4F",X"80",X"90",X"80",X"90",X"80",X"90",X"A0",X"90",X"C0",
		X"90",X"05",X"76",X"4F",X"80",X"90",X"80",X"90",X"A0",X"90",X"C0",X"90",X"04",X"76",X"4F",X"80",
		X"90",X"A0",X"90",X"C0",X"90",X"03",X"76",X"4F",X"A0",X"90",X"C0",X"90",X"02",X"76",X"4F",X"C0",
		X"90",X"01",X"76",X"4F",X"3A",X"00",X"40",X"FE",X"55",X"CA",X"00",X"40",X"31",X"00",X"A0",X"ED",
		X"46",X"F3",X"32",X"80",X"A0",X"21",X"00",X"98",X"11",X"01",X"98",X"01",X"00",X"08",X"36",X"00",
		X"ED",X"B0",X"21",X"00",X"80",X"06",X"40",X"36",X"00",X"23",X"10",X"FB",X"01",X"C0",X"07",X"11",
		X"41",X"80",X"36",X"20",X"ED",X"B0",X"32",X"80",X"A0",X"21",X"00",X"88",X"06",X"08",X"36",X"BA",
		X"23",X"10",X"FB",X"06",X"18",X"36",X"20",X"23",X"10",X"FB",X"21",X"00",X"88",X"11",X"20",X"88",
		X"01",X"E0",X"03",X"ED",X"B0",X"21",X"00",X"88",X"06",X"40",X"36",X"00",X"23",X"10",X"FB",X"21",
		X"42",X"88",X"11",X"20",X"00",X"06",X"1C",X"36",X"8E",X"19",X"10",X"FB",X"21",X"00",X"8C",X"11",
		X"01",X"8C",X"01",X"00",X"04",X"36",X"48",X"ED",X"B0",X"21",X"3F",X"A0",X"06",X"10",X"36",X"00",
		X"23",X"10",X"FB",X"21",X"80",X"A1",X"06",X"08",X"36",X"00",X"23",X"10",X"FB",X"21",X"21",X"15",
		X"11",X"00",X"9E",X"01",X"11",X"00",X"ED",X"B0",X"21",X"32",X"15",X"11",X"40",X"99",X"01",X"A0",
		X"00",X"ED",X"B0",X"3E",X"02",X"32",X"1E",X"99",X"3A",X"80",X"A1",X"2F",X"4F",X"07",X"E6",X"01",
		X"32",X"34",X"99",X"79",X"07",X"07",X"E6",X"01",X"32",X"2E",X"99",X"79",X"E6",X"07",X"21",X"19",
		X"15",X"CF",X"7E",X"32",X"26",X"99",X"79",X"0F",X"0F",X"0F",X"E6",X"07",X"21",X"19",X"15",X"CF",
		X"7E",X"32",X"29",X"99",X"AF",X"CD",X"78",X"33",X"3E",X"00",X"32",X"2D",X"99",X"3E",X"01",X"32",
		X"83",X"A1",X"32",X"2F",X"99",X"3A",X"34",X"99",X"A7",X"C2",X"DF",X"15",X"C3",X"D2",X"15",X"3E",
		X"01",X"32",X"81",X"A1",X"32",X"80",X"A0",X"18",X"FE",X"01",X"02",X"03",X"04",X"11",X"21",X"31",
		X"33",X"FF",X"05",X"F6",X"80",X"32",X"17",X"9C",X"C9",X"DD",X"21",X"74",X"98",X"FD",X"BF",X"24",
		X"AE",X"46",X"00",X"00",X"02",X"48",X"49",X"52",X"4F",X"53",X"48",X"49",X"54",X"41",X"5B",X"5B",
		X"5B",X"5B",X"80",X"99",X"01",X"49",X"4E",X"4F",X"55",X"45",X"5B",X"5B",X"5B",X"5B",X"5B",X"5B",
		X"5B",X"5B",X"50",X"88",X"01",X"4E",X"55",X"4D",X"41",X"5B",X"5B",X"5B",X"5B",X"5B",X"5B",X"5B",
		X"5B",X"5B",X"00",X"64",X"01",X"46",X"55",X"4A",X"49",X"4E",X"41",X"4B",X"41",X"5B",X"5B",X"5B",
		X"5B",X"5B",X"10",X"13",X"01",X"46",X"55",X"4B",X"55",X"54",X"41",X"4B",X"45",X"5B",X"5B",X"5B",
		X"5B",X"5B",X"60",X"05",X"01",X"54",X"41",X"4D",X"4F",X"54",X"53",X"55",X"5B",X"5B",X"5B",X"5B",
		X"5B",X"5B",X"90",X"90",X"00",X"4F",X"53",X"48",X"49",X"54",X"41",X"5B",X"5B",X"5B",X"5B",X"5B",
		X"5B",X"5B",X"30",X"90",X"00",X"54",X"53",X"55",X"44",X"41",X"5B",X"5B",X"5B",X"5B",X"5B",X"5B",
		X"5B",X"5B",X"90",X"86",X"00",X"4D",X"49",X"59",X"4F",X"53",X"48",X"49",X"5B",X"5B",X"5B",X"5B",
		X"5B",X"5B",X"10",X"82",X"00",X"48",X"41",X"52",X"41",X"5B",X"54",X"5B",X"5B",X"5B",X"5B",X"5B",
		X"5B",X"5B",X"11",X"BA",X"84",X"21",X"D3",X"16",X"0E",X"8E",X"CD",X"DA",X"16",X"18",X"16",X"11",
		X"44",X"80",X"21",X"BF",X"16",X"0E",X"87",X"CD",X"DA",X"16",X"11",X"BA",X"84",X"21",X"BF",X"16",
		X"0E",X"87",X"CD",X"DA",X"16",X"11",X"B8",X"84",X"21",X"A3",X"16",X"0E",X"BA",X"CD",X"DA",X"16",
		X"11",X"F8",X"85",X"21",X"B3",X"16",X"0E",X"BA",X"CD",X"DA",X"16",X"11",X"D8",X"86",X"21",X"B9",
		X"16",X"0E",X"BA",X"CD",X"DA",X"16",X"11",X"98",X"85",X"3A",X"26",X"99",X"0F",X"0F",X"0F",X"0F",
		X"E6",X"07",X"3C",X"CD",X"B1",X"30",X"11",X"78",X"86",X"3A",X"26",X"99",X"E6",X"07",X"CD",X"B1",
		X"30",X"11",X"B6",X"84",X"21",X"AB",X"16",X"0E",X"BA",X"CD",X"DA",X"16",X"11",X"F6",X"85",X"21",
		X"B3",X"16",X"0E",X"BA",X"CD",X"DA",X"16",X"11",X"D6",X"86",X"21",X"B9",X"16",X"0E",X"BA",X"CD",
		X"DA",X"16",X"11",X"96",X"85",X"3A",X"29",X"99",X"0F",X"0F",X"0F",X"0F",X"E6",X"07",X"3C",X"CD",
		X"B1",X"30",X"11",X"76",X"86",X"3A",X"29",X"99",X"E6",X"07",X"CD",X"B1",X"30",X"11",X"B4",X"84",
		X"0E",X"BA",X"21",X"CD",X"16",X"3A",X"2E",X"99",X"A7",X"28",X"03",X"21",X"C4",X"16",X"CD",X"DA",
		X"16",X"06",X"06",X"C5",X"06",X"00",X"C5",X"32",X"80",X"A0",X"3E",X"87",X"32",X"B8",X"8D",X"32",
		X"98",X"8E",X"32",X"B6",X"8D",X"32",X"96",X"8E",X"10",X"F0",X"C1",X"10",X"E9",X"C1",X"10",X"E3",
		X"C3",X"0F",X"15",X"43",X"4F",X"49",X"4E",X"01",X"20",X"20",X"40",X"43",X"4F",X"49",X"4E",X"02",
		X"20",X"20",X"40",X"43",X"4F",X"49",X"4E",X"20",X"40",X"50",X"4C",X"41",X"59",X"20",X"40",X"54",
		X"45",X"53",X"54",X"40",X"55",X"50",X"20",X"52",X"49",X"47",X"48",X"54",X"40",X"54",X"41",X"42",
		X"4C",X"45",X"40",X"4E",X"4F",X"52",X"4D",X"41",X"4C",X"40",X"E5",X"D5",X"CD",X"F2",X"30",X"D1",
		X"E1",X"FF",X"C9",X"11",X"00",X"9B",X"01",X"18",X"00",X"ED",X"B0",X"32",X"04",X"99",X"21",X"80",
		X"9A",X"11",X"81",X"9A",X"01",X"0C",X"00",X"36",X"00",X"ED",X"B0",X"AF",X"32",X"60",X"98",X"C9",
		X"11",X"40",X"9B",X"01",X"18",X"00",X"ED",X"B0",X"32",X"05",X"99",X"21",X"A0",X"9A",X"11",X"A1",
		X"9A",X"01",X"0C",X"00",X"36",X"02",X"ED",X"B0",X"AF",X"32",X"63",X"98",X"C9",X"21",X"04",X"99",
		X"7E",X"A7",X"20",X"03",X"3E",X"08",X"77",X"CD",X"4F",X"1E",X"32",X"62",X"98",X"21",X"48",X"17",
		X"11",X"80",X"9A",X"01",X"0C",X"00",X"ED",X"B0",X"21",X"53",X"17",X"11",X"00",X"9B",X"01",X"18",
		X"00",X"ED",X"B0",X"AF",X"32",X"60",X"98",X"C9",X"01",X"01",X"05",X"10",X"0F",X"0A",X"05",X"00",
		X"02",X"10",X"07",X"EF",X"85",X"EE",X"85",X"ED",X"85",X"0D",X"86",X"0E",X"86",X"EE",X"85",X"ED",
		X"85",X"0D",X"86",X"ED",X"85",X"0D",X"86",X"0E",X"86",X"EE",X"85",X"3A",X"03",X"99",X"E6",X"03",
		X"28",X"44",X"21",X"79",X"84",X"22",X"40",X"9B",X"21",X"7A",X"84",X"22",X"42",X"9B",X"21",X"42",
		X"9B",X"11",X"44",X"9B",X"01",X"16",X"00",X"ED",X"B0",X"3A",X"05",X"99",X"A7",X"20",X"0F",X"21",
		X"03",X"99",X"7E",X"A7",X"C8",X"35",X"CD",X"B8",X"3F",X"3E",X"09",X"32",X"05",X"99",X"CD",X"40",
		X"1E",X"32",X"65",X"98",X"21",X"A0",X"9A",X"11",X"A1",X"9A",X"01",X"0C",X"00",X"36",X"03",X"ED",
		X"B0",X"AF",X"32",X"63",X"98",X"C9",X"21",X"7A",X"87",X"22",X"40",X"9B",X"21",X"9A",X"87",X"22",
		X"42",X"9B",X"21",X"42",X"9B",X"11",X"44",X"9B",X"01",X"16",X"00",X"ED",X"B0",X"21",X"03",X"99",
		X"7E",X"A7",X"C8",X"35",X"CD",X"B8",X"3F",X"3E",X"09",X"32",X"05",X"99",X"CD",X"40",X"1E",X"32",
		X"65",X"98",X"21",X"A0",X"9A",X"11",X"A1",X"9A",X"01",X"0C",X"00",X"36",X"00",X"ED",X"B0",X"AF",
		X"32",X"63",X"98",X"C9",X"3A",X"03",X"99",X"E6",X"03",X"28",X"44",X"21",X"82",X"84",X"22",X"80",
		X"9B",X"21",X"62",X"84",X"22",X"82",X"9B",X"21",X"82",X"9B",X"11",X"84",X"9B",X"01",X"16",X"00",
		X"ED",X"B0",X"3A",X"06",X"99",X"A7",X"20",X"0F",X"21",X"03",X"99",X"7E",X"A7",X"C8",X"35",X"CD",
		X"B8",X"3F",X"3E",X"09",X"32",X"06",X"99",X"CD",X"40",X"1E",X"32",X"68",X"98",X"21",X"C0",X"9A",
		X"11",X"C1",X"9A",X"01",X"0C",X"00",X"36",X"02",X"ED",X"B0",X"AF",X"32",X"66",X"98",X"C9",X"21",
		X"7A",X"87",X"22",X"80",X"9B",X"21",X"9A",X"87",X"22",X"82",X"9B",X"21",X"82",X"9B",X"11",X"84",
		X"9B",X"01",X"16",X"00",X"ED",X"B0",X"21",X"03",X"99",X"7E",X"A7",X"C8",X"35",X"CD",X"B8",X"3F",
		X"3E",X"09",X"32",X"06",X"99",X"CD",X"40",X"1E",X"32",X"68",X"98",X"21",X"C0",X"9A",X"11",X"C1",
		X"9A",X"01",X"0C",X"00",X"36",X"00",X"ED",X"B0",X"AF",X"32",X"66",X"98",X"C9",X"3A",X"03",X"99",
		X"E6",X"03",X"28",X"44",X"21",X"83",X"87",X"22",X"C0",X"9B",X"21",X"82",X"87",X"22",X"C2",X"9B",
		X"21",X"C2",X"9B",X"11",X"C4",X"9B",X"01",X"16",X"00",X"ED",X"B0",X"3A",X"07",X"99",X"A7",X"20",
		X"0F",X"21",X"03",X"99",X"7E",X"A7",X"C8",X"35",X"CD",X"B8",X"3F",X"3E",X"09",X"32",X"07",X"99",
		X"CD",X"40",X"1E",X"32",X"6B",X"98",X"21",X"E0",X"9A",X"11",X"E1",X"9A",X"01",X"0C",X"00",X"36",
		X"01",X"ED",X"B0",X"AF",X"32",X"69",X"98",X"C9",X"21",X"7A",X"87",X"22",X"C0",X"9B",X"21",X"9A",
		X"87",X"22",X"C2",X"9B",X"21",X"C2",X"9B",X"11",X"C4",X"9B",X"01",X"16",X"00",X"ED",X"B0",X"21",
		X"03",X"99",X"7E",X"A7",X"C8",X"35",X"CD",X"B8",X"3F",X"3E",X"09",X"32",X"07",X"99",X"CD",X"40",
		X"1E",X"32",X"6B",X"98",X"21",X"E0",X"9A",X"11",X"E1",X"9A",X"01",X"0C",X"00",X"36",X"00",X"ED",
		X"B0",X"AF",X"32",X"69",X"98",X"C9",X"21",X"A7",X"80",X"11",X"E0",X"FF",X"3A",X"00",X"99",X"FE",
		X"05",X"30",X"1C",X"4F",X"3E",X"04",X"91",X"28",X"06",X"47",X"36",X"20",X"19",X"10",X"FB",X"79",
		X"A7",X"28",X"0C",X"47",X"36",X"5E",X"CB",X"DC",X"36",X"AB",X"CB",X"9C",X"19",X"10",X"F5",X"21",
		X"24",X"81",X"11",X"E0",X"FF",X"3A",X"0A",X"99",X"FE",X"09",X"D0",X"4F",X"3E",X"08",X"91",X"28",
		X"06",X"47",X"36",X"20",X"19",X"10",X"FB",X"79",X"A7",X"C8",X"47",X"36",X"5F",X"CB",X"DC",X"36",
		X"AB",X"CB",X"9C",X"19",X"10",X"F5",X"C9",X"3A",X"01",X"99",X"FE",X"19",X"D0",X"4F",X"21",X"A7",
		X"8B",X"11",X"E0",X"FF",X"06",X"06",X"36",X"89",X"19",X"36",X"89",X"19",X"36",X"89",X"19",X"36",
		X"95",X"19",X"10",X"F2",X"21",X"A7",X"83",X"41",X"36",X"5D",X"19",X"10",X"FB",X"3E",X"18",X"91",
		X"C8",X"47",X"36",X"20",X"19",X"10",X"FB",X"C9",X"11",X"78",X"8C",X"01",X"18",X"04",X"3E",X"8E",
		X"CD",X"6D",X"1A",X"11",X"18",X"8D",X"01",X"18",X"06",X"3E",X"BA",X"CD",X"6D",X"1A",X"11",X"F8",
		X"8D",X"01",X"13",X"0C",X"3E",X"95",X"CD",X"6D",X"1A",X"21",X"8A",X"01",X"11",X"3A",X"85",X"0E",
		X"BE",X"CD",X"DA",X"16",X"AF",X"32",X"40",X"98",X"C9",X"3A",X"02",X"98",X"E6",X"01",X"FE",X"01",
		X"D8",X"11",X"D8",X"84",X"21",X"47",X"1A",X"3A",X"40",X"98",X"47",X"A7",X"28",X"05",X"23",X"1B",
		X"1B",X"10",X"FB",X"7E",X"12",X"11",X"B8",X"84",X"21",X"51",X"1A",X"3A",X"40",X"98",X"47",X"A7",
		X"28",X"05",X"23",X"1B",X"1B",X"10",X"FB",X"7E",X"12",X"11",X"78",X"84",X"3A",X"40",X"98",X"47",
		X"A7",X"28",X"04",X"1B",X"1B",X"10",X"FC",X"C6",X"01",X"27",X"CD",X"B1",X"30",X"11",X"18",X"85",
		X"21",X"42",X"99",X"01",X"10",X"00",X"3A",X"40",X"98",X"A7",X"28",X"06",X"1B",X"1B",X"09",X"3D",
		X"20",X"FA",X"06",X"00",X"7E",X"CD",X"C9",X"30",X"2B",X"7E",X"CD",X"C9",X"30",X"2B",X"7E",X"CD",
		X"B6",X"30",X"11",X"F8",X"85",X"21",X"43",X"99",X"01",X"10",X"00",X"3A",X"40",X"98",X"A7",X"28",
		X"06",X"1B",X"1B",X"09",X"3D",X"20",X"FA",X"06",X"0C",X"7E",X"12",X"23",X"D7",X"10",X"FA",X"21",
		X"40",X"98",X"34",X"7E",X"FE",X"0A",X"C9",X"54",X"44",X"44",X"48",X"48",X"48",X"48",X"48",X"48",
		X"48",X"53",X"4E",X"52",X"54",X"54",X"54",X"54",X"54",X"54",X"54",X"11",X"9B",X"87",X"06",X"1A",
		X"3E",X"41",X"12",X"1B",X"3C",X"10",X"FB",X"EF",X"21",X"9F",X"01",X"FF",X"C9",X"C5",X"41",X"D5",
		X"12",X"1B",X"10",X"FC",X"D1",X"F5",X"D7",X"F1",X"C1",X"10",X"F2",X"C9",X"21",X"40",X"98",X"7E",
		X"C6",X"01",X"27",X"77",X"21",X"2F",X"01",X"11",X"82",X"81",X"D5",X"E5",X"FF",X"21",X"1F",X"FF",
		X"19",X"EB",X"3A",X"1E",X"99",X"06",X"00",X"CD",X"C9",X"30",X"3A",X"1D",X"99",X"CD",X"C9",X"30",
		X"3A",X"1C",X"99",X"CD",X"B6",X"30",X"E1",X"D1",X"0E",X"87",X"C3",X"F2",X"30",X"21",X"12",X"99",
		X"06",X"0A",X"36",X"00",X"23",X"10",X"FB",X"C9",X"21",X"00",X"98",X"06",X"00",X"36",X"00",X"23",
		X"10",X"FB",X"C9",X"21",X"00",X"9A",X"11",X"01",X"9A",X"01",X"FF",X"03",X"36",X"00",X"ED",X"B0",
		X"C9",X"AF",X"21",X"34",X"9C",X"06",X"08",X"77",X"23",X"10",X"FC",X"32",X"10",X"9C",X"32",X"12",
		X"9C",X"32",X"14",X"9C",X"32",X"16",X"9C",X"32",X"18",X"9C",X"32",X"1A",X"9C",X"2A",X"52",X"98",
		X"06",X"20",X"36",X"20",X"CB",X"DC",X"36",X"BF",X"CB",X"9C",X"23",X"10",X"F5",X"22",X"52",X"98",
		X"21",X"01",X"98",X"35",X"C9",X"21",X"A4",X"83",X"11",X"E0",X"FF",X"06",X"08",X"36",X"20",X"19",
		X"10",X"FB",X"AF",X"21",X"34",X"9C",X"06",X"08",X"77",X"23",X"10",X"FC",X"32",X"00",X"9D",X"21",
		X"00",X"9B",X"CD",X"47",X"1B",X"21",X"40",X"9B",X"CD",X"47",X"1B",X"21",X"80",X"9B",X"CD",X"47",
		X"1B",X"21",X"C0",X"9B",X"AF",X"32",X"10",X"9C",X"32",X"12",X"9C",X"32",X"14",X"9C",X"32",X"16",
		X"9C",X"32",X"18",X"9C",X"32",X"1A",X"9C",X"06",X"0A",X"3E",X"20",X"5E",X"23",X"56",X"23",X"7B",
		X"B2",X"28",X"03",X"3E",X"20",X"12",X"10",X"F3",X"C9",X"CD",X"AB",X"1B",X"C0",X"3A",X"04",X"99",
		X"A7",X"C8",X"DD",X"21",X"74",X"98",X"DD",X"7E",X"00",X"A7",X"28",X"07",X"DD",X"23",X"DD",X"7E",
		X"00",X"A7",X"C0",X"CD",X"A5",X"33",X"3A",X"61",X"98",X"DD",X"77",X"10",X"3A",X"6C",X"98",X"DD",
		X"77",X"20",X"3A",X"80",X"9A",X"E6",X"03",X"87",X"21",X"A3",X"1B",X"CF",X"7E",X"DD",X"77",X"30",
		X"23",X"7E",X"DD",X"77",X"40",X"3E",X"FF",X"DD",X"77",X"00",X"C9",X"02",X"00",X"00",X"02",X"FE",
		X"00",X"00",X"FE",X"03",X"00",X"00",X"03",X"FD",X"00",X"00",X"FD",X"21",X"15",X"98",X"3A",X"2F",
		X"99",X"A7",X"3A",X"04",X"98",X"28",X"03",X"3A",X"03",X"98",X"0F",X"0F",X"0F",X"0F",X"CB",X"16",
		X"7E",X"E6",X"07",X"FE",X"01",X"C9",X"3A",X"71",X"98",X"A7",X"28",X"07",X"DD",X"21",X"76",X"98",
		X"CD",X"27",X"1C",X"3A",X"72",X"98",X"A7",X"28",X"07",X"DD",X"21",X"78",X"98",X"CD",X"65",X"1C",
		X"3A",X"73",X"98",X"A7",X"C8",X"DD",X"21",X"7A",X"98",X"DD",X"7E",X"00",X"A7",X"28",X"07",X"DD",
		X"23",X"DD",X"7E",X"00",X"A7",X"C0",X"3A",X"02",X"98",X"E6",X"0F",X"C0",X"32",X"73",X"98",X"CD",
		X"A9",X"33",X"3A",X"6A",X"98",X"DD",X"77",X"10",X"3A",X"6F",X"98",X"DD",X"77",X"20",X"3A",X"E0",
		X"9A",X"E6",X"03",X"87",X"21",X"9B",X"1B",X"CF",X"7E",X"DD",X"77",X"30",X"23",X"7E",X"DD",X"77",
		X"40",X"3E",X"FF",X"DD",X"77",X"00",X"C9",X"DD",X"7E",X"00",X"A7",X"28",X"07",X"DD",X"23",X"DD",
		X"7E",X"00",X"A7",X"C0",X"3A",X"02",X"98",X"E6",X"0F",X"C0",X"32",X"71",X"98",X"CD",X"A9",X"33",
		X"3A",X"64",X"98",X"DD",X"77",X"10",X"3A",X"6D",X"98",X"DD",X"77",X"20",X"3A",X"A0",X"9A",X"E6",
		X"03",X"87",X"21",X"9B",X"1B",X"CF",X"7E",X"DD",X"77",X"30",X"23",X"7E",X"DD",X"77",X"40",X"3E",
		X"FF",X"DD",X"77",X"00",X"C9",X"DD",X"7E",X"00",X"A7",X"28",X"07",X"DD",X"23",X"DD",X"7E",X"00",
		X"A7",X"C0",X"3A",X"02",X"98",X"E6",X"0F",X"C0",X"32",X"72",X"98",X"CD",X"A9",X"33",X"3A",X"67",
		X"98",X"DD",X"77",X"10",X"3A",X"6E",X"98",X"DD",X"77",X"20",X"3A",X"C0",X"9A",X"E6",X"03",X"87",
		X"21",X"9B",X"1B",X"CF",X"7E",X"DD",X"77",X"30",X"23",X"7E",X"DD",X"77",X"40",X"3E",X"FF",X"DD",
		X"77",X"00",X"C9",X"3A",X"70",X"98",X"A7",X"C8",X"AF",X"32",X"70",X"98",X"DD",X"21",X"74",X"98",
		X"DD",X"7E",X"00",X"A7",X"28",X"07",X"DD",X"23",X"DD",X"7E",X"00",X"A7",X"C0",X"CD",X"A5",X"33",
		X"3A",X"61",X"98",X"DD",X"77",X"10",X"3A",X"6C",X"98",X"DD",X"77",X"20",X"3A",X"80",X"9A",X"E6",
		X"03",X"87",X"21",X"A3",X"1B",X"CF",X"7E",X"DD",X"77",X"30",X"23",X"7E",X"DD",X"77",X"40",X"3E",
		X"FF",X"DD",X"77",X"00",X"C9",X"FD",X"21",X"74",X"98",X"CD",X"EE",X"1C",X"FD",X"23",X"FD",X"7E",
		X"00",X"A7",X"C8",X"FD",X"7E",X"20",X"FD",X"86",X"40",X"FD",X"77",X"20",X"4F",X"FD",X"7E",X"10",
		X"FD",X"86",X"30",X"FD",X"77",X"10",X"2F",X"E6",X"F8",X"26",X"00",X"6F",X"29",X"29",X"79",X"E6",
		X"F8",X"0F",X"0F",X"0F",X"CF",X"11",X"00",X"84",X"19",X"7E",X"FE",X"E8",X"D2",X"DF",X"1D",X"EB",
		X"3A",X"05",X"99",X"A7",X"28",X"3B",X"DD",X"21",X"C4",X"98",X"CD",X"E4",X"1D",X"20",X"32",X"21",
		X"05",X"99",X"35",X"20",X"1E",X"AF",X"32",X"71",X"98",X"3E",X"40",X"32",X"81",X"98",X"CD",X"BF",
		X"31",X"28",X"03",X"32",X"B1",X"98",X"3E",X"01",X"32",X"91",X"98",X"32",X"A1",X"98",X"CD",X"11",
		X"1E",X"18",X"03",X"CD",X"F8",X"1D",X"3A",X"05",X"99",X"CD",X"40",X"1E",X"32",X"65",X"98",X"18",
		X"7E",X"3A",X"06",X"99",X"A7",X"28",X"3B",X"DD",X"21",X"C8",X"98",X"CD",X"E4",X"1D",X"20",X"32",
		X"21",X"06",X"99",X"35",X"20",X"1E",X"AF",X"32",X"72",X"98",X"3E",X"40",X"32",X"82",X"98",X"CD",
		X"BF",X"31",X"28",X"03",X"32",X"B2",X"98",X"3E",X"01",X"32",X"92",X"98",X"32",X"A2",X"98",X"CD",
		X"11",X"1E",X"18",X"03",X"CD",X"F8",X"1D",X"3A",X"06",X"99",X"CD",X"40",X"1E",X"32",X"68",X"98",
		X"18",X"3D",X"3A",X"07",X"99",X"A7",X"C8",X"DD",X"21",X"CC",X"98",X"CD",X"E4",X"1D",X"C0",X"21",
		X"07",X"99",X"35",X"20",X"1E",X"AF",X"32",X"73",X"98",X"3E",X"40",X"32",X"83",X"98",X"CD",X"BF",
		X"31",X"28",X"03",X"32",X"B3",X"98",X"3E",X"01",X"32",X"93",X"98",X"32",X"A3",X"98",X"CD",X"11",
		X"1E",X"18",X"03",X"CD",X"F8",X"1D",X"3A",X"07",X"99",X"CD",X"40",X"1E",X"32",X"6B",X"98",X"AF",
		X"FD",X"77",X"00",X"C9",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"AF",X"ED",X"52",X"C8",X"DD",X"6E",
		X"02",X"DD",X"66",X"03",X"AF",X"ED",X"52",X"C9",X"FD",X"E5",X"21",X"60",X"00",X"3E",X"FF",X"32",
		X"47",X"98",X"22",X"15",X"99",X"22",X"1A",X"99",X"CD",X"FE",X"30",X"CD",X"EB",X"33",X"FD",X"E1",
		X"C9",X"FD",X"E5",X"21",X"00",X"05",X"3E",X"FF",X"32",X"47",X"98",X"22",X"15",X"99",X"22",X"1A",
		X"99",X"CD",X"FE",X"30",X"CD",X"EF",X"33",X"FD",X"E1",X"C9",X"00",X"2A",X"28",X"26",X"24",X"22",
		X"20",X"1E",X"1C",X"1A",X"16",X"00",X"2C",X"2A",X"28",X"26",X"24",X"22",X"20",X"1E",X"1C",X"1A",
		X"21",X"2A",X"1E",X"CF",X"3A",X"01",X"99",X"3D",X"86",X"FE",X"39",X"D8",X"3E",X"38",X"C9",X"21",
		X"35",X"1E",X"18",X"EF",X"DD",X"21",X"76",X"98",X"CD",X"71",X"1E",X"DD",X"23",X"CD",X"71",X"1E",
		X"DD",X"23",X"CD",X"71",X"1E",X"DD",X"23",X"CD",X"71",X"1E",X"DD",X"23",X"CD",X"71",X"1E",X"DD",
		X"23",X"DD",X"7E",X"00",X"A7",X"C8",X"DD",X"7E",X"20",X"DD",X"86",X"40",X"DD",X"77",X"20",X"4F",
		X"DD",X"7E",X"10",X"DD",X"86",X"30",X"DD",X"77",X"10",X"2F",X"E6",X"F8",X"26",X"00",X"6F",X"29",
		X"29",X"79",X"E6",X"F8",X"0F",X"0F",X"0F",X"CF",X"11",X"00",X"84",X"19",X"7E",X"FE",X"E8",X"30",
		X"3C",X"3A",X"04",X"99",X"A7",X"C8",X"EB",X"2A",X"C0",X"98",X"A7",X"ED",X"52",X"20",X"07",X"3A",
		X"60",X"98",X"FE",X"A0",X"38",X"0D",X"2A",X"C2",X"98",X"A7",X"ED",X"52",X"C0",X"3A",X"60",X"98",
		X"FE",X"80",X"D8",X"CD",X"E7",X"33",X"21",X"04",X"99",X"35",X"20",X"0A",X"3E",X"40",X"32",X"80",
		X"98",X"3E",X"01",X"32",X"90",X"98",X"7E",X"CD",X"4F",X"1E",X"32",X"62",X"98",X"AF",X"DD",X"77",
		X"00",X"C9",X"FD",X"21",X"74",X"98",X"06",X"08",X"CD",X"2B",X"1F",X"FD",X"23",X"10",X"F9",X"CD",
		X"3A",X"25",X"3A",X"D3",X"98",X"A7",X"20",X"03",X"CD",X"47",X"2A",X"CD",X"65",X"2E",X"3A",X"D2",
		X"98",X"A7",X"20",X"03",X"CD",X"A8",X"28",X"CD",X"25",X"2E",X"3A",X"D1",X"98",X"A7",X"20",X"03",
		X"CD",X"F5",X"26",X"CD",X"E5",X"2D",X"CD",X"DE",X"25",X"CD",X"A0",X"2D",X"CD",X"63",X"1F",X"CD",
		X"BA",X"1F",X"CD",X"09",X"20",X"CD",X"58",X"20",X"C3",X"AD",X"23",X"FD",X"7E",X"00",X"A7",X"C8",
		X"FD",X"7E",X"20",X"FD",X"86",X"40",X"FD",X"77",X"20",X"4F",X"FD",X"7E",X"10",X"FD",X"86",X"30",
		X"FD",X"77",X"10",X"2F",X"E6",X"F8",X"26",X"00",X"6F",X"29",X"29",X"79",X"E6",X"F8",X"0F",X"0F",
		X"0F",X"CF",X"11",X"00",X"84",X"19",X"7E",X"FE",X"E8",X"D8",X"FD",X"36",X"00",X"00",X"FD",X"36",
		X"10",X"00",X"C9",X"2A",X"02",X"9B",X"11",X"00",X"84",X"A7",X"ED",X"52",X"7D",X"E6",X"1F",X"87",
		X"87",X"87",X"C6",X"04",X"32",X"6C",X"98",X"CB",X"3C",X"CB",X"1D",X"CB",X"3C",X"CB",X"1D",X"7D",
		X"E6",X"F8",X"C6",X"04",X"2F",X"32",X"61",X"98",X"3A",X"60",X"98",X"07",X"07",X"07",X"E6",X"07",
		X"C8",X"47",X"4F",X"3A",X"80",X"9A",X"E6",X"03",X"21",X"B2",X"1F",X"87",X"CF",X"3A",X"61",X"98",
		X"86",X"10",X"FD",X"32",X"61",X"98",X"23",X"3A",X"6C",X"98",X"41",X"86",X"10",X"FD",X"32",X"6C",
		X"98",X"C9",X"01",X"00",X"00",X"01",X"FF",X"00",X"00",X"FF",X"2A",X"42",X"9B",X"11",X"00",X"84",
		X"A7",X"ED",X"52",X"7D",X"E6",X"1F",X"87",X"87",X"87",X"C6",X"04",X"32",X"6D",X"98",X"CB",X"3C",
		X"CB",X"1D",X"CB",X"3C",X"CB",X"1D",X"7D",X"E6",X"F8",X"C6",X"04",X"2F",X"32",X"64",X"98",X"3A",
		X"63",X"98",X"07",X"07",X"07",X"E6",X"07",X"C8",X"47",X"4F",X"3A",X"A1",X"9A",X"E6",X"03",X"21",
		X"B2",X"1F",X"87",X"CF",X"3A",X"64",X"98",X"86",X"10",X"FD",X"32",X"64",X"98",X"23",X"3A",X"6D",
		X"98",X"41",X"86",X"10",X"FD",X"32",X"6D",X"98",X"C9",X"2A",X"82",X"9B",X"11",X"00",X"84",X"A7",
		X"ED",X"52",X"7D",X"E6",X"1F",X"87",X"87",X"87",X"C6",X"04",X"32",X"6E",X"98",X"CB",X"3C",X"CB",
		X"1D",X"CB",X"3C",X"CB",X"1D",X"7D",X"E6",X"F8",X"C6",X"04",X"2F",X"32",X"67",X"98",X"3A",X"66",
		X"98",X"07",X"07",X"07",X"E6",X"07",X"C8",X"47",X"4F",X"3A",X"C1",X"9A",X"E6",X"03",X"21",X"B2",
		X"1F",X"87",X"CF",X"3A",X"67",X"98",X"86",X"10",X"FD",X"32",X"67",X"98",X"23",X"3A",X"6E",X"98",
		X"41",X"86",X"10",X"FD",X"32",X"6E",X"98",X"C9",X"2A",X"C2",X"9B",X"11",X"00",X"84",X"A7",X"ED",
		X"52",X"7D",X"E6",X"1F",X"87",X"87",X"87",X"C6",X"04",X"32",X"6F",X"98",X"CB",X"3C",X"CB",X"1D",
		X"CB",X"3C",X"CB",X"1D",X"7D",X"E6",X"F8",X"C6",X"04",X"2F",X"32",X"6A",X"98",X"3A",X"69",X"98",
		X"07",X"07",X"07",X"E6",X"07",X"C8",X"47",X"4F",X"3A",X"E1",X"9A",X"E6",X"03",X"21",X"B2",X"1F",
		X"87",X"CF",X"3A",X"6A",X"98",X"86",X"10",X"FD",X"32",X"6A",X"98",X"23",X"3A",X"6F",X"98",X"41",
		X"86",X"10",X"FD",X"32",X"6F",X"98",X"C9",X"3A",X"05",X"99",X"32",X"40",X"98",X"21",X"64",X"98",
		X"11",X"6D",X"98",X"DD",X"21",X"81",X"98",X"CD",X"04",X"21",X"3A",X"40",X"98",X"32",X"05",X"99",
		X"A7",X"20",X"03",X"32",X"71",X"98",X"3A",X"06",X"99",X"32",X"40",X"98",X"21",X"67",X"98",X"11",
		X"6E",X"98",X"DD",X"21",X"82",X"98",X"CD",X"04",X"21",X"3A",X"40",X"98",X"32",X"06",X"99",X"A7",
		X"20",X"03",X"32",X"72",X"98",X"3A",X"07",X"99",X"32",X"40",X"98",X"21",X"6A",X"98",X"11",X"6F",
		X"98",X"DD",X"21",X"83",X"98",X"CD",X"04",X"21",X"3A",X"40",X"98",X"32",X"07",X"99",X"A7",X"C0",
		X"32",X"73",X"98",X"C9",X"3A",X"04",X"99",X"A7",X"C8",X"3A",X"40",X"98",X"A7",X"C8",X"3A",X"61",
		X"98",X"96",X"30",X"02",X"ED",X"44",X"FE",X"08",X"D0",X"47",X"EB",X"3A",X"6C",X"98",X"96",X"30",
		X"02",X"ED",X"44",X"FE",X"08",X"D0",X"A7",X"28",X"03",X"78",X"A7",X"C0",X"21",X"40",X"98",X"3A",
		X"04",X"99",X"BE",X"38",X"24",X"3E",X"40",X"DD",X"77",X"00",X"CD",X"BF",X"31",X"28",X"03",X"DD",
		X"77",X"30",X"21",X"40",X"98",X"7E",X"36",X"00",X"DD",X"77",X"10",X"21",X"68",X"21",X"DF",X"EB",
		X"22",X"15",X"99",X"22",X"1A",X"99",X"C3",X"FE",X"30",X"3E",X"40",X"32",X"80",X"98",X"21",X"04",
		X"99",X"7E",X"36",X"00",X"32",X"90",X"98",X"C9",X"00",X"00",X"80",X"00",X"60",X"01",X"40",X"02",
		X"20",X"03",X"00",X"04",X"80",X"04",X"60",X"05",X"40",X"06",X"00",X"08",X"21",X"80",X"98",X"7E",
		X"A7",X"C8",X"35",X"28",X"2F",X"7E",X"FE",X"2A",X"28",X"4F",X"FE",X"15",X"28",X"51",X"FE",X"3E",
		X"C0",X"CD",X"AD",X"33",X"21",X"02",X"9B",X"3A",X"90",X"98",X"3D",X"28",X"0B",X"47",X"04",X"3E",
		X"74",X"5E",X"2C",X"56",X"2C",X"12",X"10",X"F9",X"5E",X"2C",X"56",X"3E",X"20",X"12",X"3E",X"64",
		X"32",X"00",X"9C",X"C9",X"3A",X"90",X"98",X"3D",X"28",X"19",X"4F",X"0C",X"11",X"02",X"9B",X"21",
		X"50",X"9C",X"7E",X"3C",X"87",X"47",X"7E",X"81",X"77",X"78",X"85",X"6F",X"EB",X"CB",X"21",X"06",
		X"00",X"ED",X"B0",X"3E",X"20",X"32",X"00",X"9C",X"C9",X"3E",X"68",X"32",X"00",X"9C",X"C9",X"3E",
		X"6C",X"32",X"00",X"9C",X"C9",X"21",X"81",X"98",X"7E",X"A7",X"C8",X"35",X"28",X"35",X"3A",X"A1",
		X"98",X"A7",X"20",X"67",X"7E",X"FE",X"2A",X"28",X"56",X"FE",X"15",X"28",X"58",X"FE",X"3E",X"C0",
		X"CD",X"C5",X"33",X"21",X"42",X"9B",X"3A",X"91",X"98",X"3D",X"28",X"0B",X"47",X"04",X"3E",X"74",
		X"5E",X"2C",X"56",X"2C",X"12",X"10",X"F9",X"5E",X"2C",X"56",X"3E",X"20",X"12",X"3E",X"64",X"32",
		X"02",X"9C",X"C9",X"3A",X"91",X"98",X"3D",X"28",X"19",X"4F",X"0C",X"11",X"42",X"9B",X"21",X"50",
		X"9C",X"7E",X"3C",X"87",X"47",X"7E",X"81",X"77",X"78",X"85",X"6F",X"EB",X"CB",X"21",X"06",X"00",
		X"ED",X"B0",X"3E",X"20",X"32",X"02",X"9C",X"AF",X"32",X"A1",X"98",X"32",X"D1",X"98",X"C9",X"3E",
		X"68",X"32",X"02",X"9C",X"C9",X"3E",X"6C",X"32",X"02",X"9C",X"C9",X"7E",X"FE",X"3E",X"C0",X"3A",
		X"2F",X"99",X"A7",X"28",X"04",X"3E",X"34",X"18",X"02",X"3E",X"37",X"32",X"02",X"9C",X"21",X"42",
		X"9B",X"5E",X"2C",X"56",X"3E",X"20",X"12",X"2C",X"5E",X"2C",X"56",X"12",X"C9",X"21",X"82",X"98",
		X"7E",X"A7",X"C8",X"35",X"28",X"35",X"3A",X"A2",X"98",X"A7",X"20",X"67",X"7E",X"FE",X"2A",X"28",
		X"56",X"FE",X"15",X"28",X"58",X"FE",X"3E",X"C0",X"CD",X"C5",X"33",X"21",X"82",X"9B",X"3A",X"92",
		X"98",X"3D",X"28",X"0B",X"47",X"04",X"3E",X"74",X"5E",X"2C",X"56",X"2C",X"12",X"10",X"F9",X"5E",
		X"2C",X"56",X"3E",X"20",X"12",X"3E",X"64",X"32",X"04",X"9C",X"C9",X"3A",X"92",X"98",X"3D",X"28",
		X"19",X"4F",X"0C",X"11",X"82",X"9B",X"21",X"50",X"9C",X"7E",X"3C",X"87",X"47",X"7E",X"81",X"77",
		X"78",X"85",X"6F",X"EB",X"CB",X"21",X"06",X"00",X"ED",X"B0",X"3E",X"20",X"32",X"04",X"9C",X"AF",
		X"32",X"A2",X"98",X"32",X"D2",X"98",X"C9",X"3E",X"68",X"32",X"04",X"9C",X"C9",X"3E",X"6C",X"32",
		X"04",X"9C",X"C9",X"7E",X"FE",X"3E",X"C0",X"3A",X"2F",X"99",X"A7",X"28",X"04",X"3E",X"34",X"18",
		X"02",X"3E",X"37",X"32",X"04",X"9C",X"21",X"82",X"9B",X"5E",X"2C",X"56",X"3E",X"20",X"12",X"2C",
		X"5E",X"2C",X"56",X"12",X"C9",X"21",X"83",X"98",X"7E",X"A7",X"C8",X"35",X"28",X"35",X"3A",X"A3",
		X"98",X"A7",X"20",X"67",X"7E",X"FE",X"2A",X"28",X"56",X"FE",X"15",X"28",X"58",X"FE",X"3E",X"C0",
		X"CD",X"C5",X"33",X"21",X"C2",X"9B",X"3A",X"93",X"98",X"3D",X"28",X"0B",X"47",X"04",X"3E",X"74",
		X"5E",X"2C",X"56",X"2C",X"12",X"10",X"F9",X"5E",X"2C",X"56",X"3E",X"20",X"12",X"3E",X"64",X"32",
		X"06",X"9C",X"C9",X"3A",X"93",X"98",X"3D",X"28",X"19",X"4F",X"0C",X"11",X"C2",X"9B",X"21",X"50",
		X"9C",X"7E",X"3C",X"87",X"47",X"7E",X"81",X"77",X"78",X"85",X"6F",X"EB",X"CB",X"21",X"06",X"00",
		X"ED",X"B0",X"3E",X"20",X"32",X"06",X"9C",X"AF",X"32",X"A3",X"98",X"32",X"D3",X"98",X"C9",X"3E",
		X"68",X"32",X"06",X"9C",X"C9",X"3E",X"6C",X"32",X"06",X"9C",X"C9",X"7E",X"FE",X"3E",X"C0",X"3A",
		X"2F",X"99",X"A7",X"28",X"04",X"3E",X"34",X"18",X"02",X"3E",X"37",X"32",X"06",X"9C",X"21",X"C2",
		X"9B",X"5E",X"2C",X"56",X"3E",X"20",X"12",X"2C",X"5E",X"2C",X"56",X"12",X"C9",X"3A",X"2F",X"99",
		X"A7",X"C2",X"65",X"24",X"3A",X"04",X"99",X"A7",X"28",X"0E",X"3A",X"80",X"9A",X"C6",X"02",X"E6",
		X"03",X"87",X"87",X"C6",X"10",X"32",X"00",X"9C",X"3A",X"05",X"99",X"A7",X"28",X"0E",X"3A",X"A1",
		X"9A",X"C6",X"02",X"E6",X"03",X"87",X"87",X"C6",X"24",X"32",X"02",X"9C",X"3A",X"06",X"99",X"A7",
		X"28",X"0E",X"3A",X"C1",X"9A",X"C6",X"02",X"E6",X"03",X"87",X"87",X"C6",X"24",X"32",X"04",X"9C",
		X"3A",X"07",X"99",X"A7",X"28",X"0E",X"3A",X"E1",X"9A",X"C6",X"02",X"E6",X"03",X"87",X"87",X"C6",
		X"24",X"32",X"06",X"9C",X"3A",X"61",X"98",X"C6",X"FA",X"32",X"10",X"9C",X"3A",X"6C",X"98",X"C6",
		X"F8",X"32",X"01",X"9C",X"3A",X"11",X"9C",X"E6",X"7F",X"32",X"11",X"9C",X"3A",X"64",X"98",X"C6",
		X"FA",X"32",X"12",X"9C",X"3A",X"6D",X"98",X"C6",X"F8",X"32",X"03",X"9C",X"3A",X"13",X"9C",X"E6",
		X"7F",X"32",X"13",X"9C",X"3A",X"67",X"98",X"C6",X"FA",X"32",X"14",X"9C",X"3A",X"6E",X"98",X"C6",
		X"F8",X"32",X"05",X"9C",X"3A",X"15",X"9C",X"E6",X"7F",X"32",X"15",X"9C",X"3A",X"6A",X"98",X"C6",
		X"FA",X"32",X"16",X"9C",X"3A",X"6F",X"98",X"C6",X"F8",X"32",X"07",X"9C",X"3A",X"17",X"9C",X"E6",
		X"7F",X"32",X"17",X"9C",X"C9",X"3A",X"04",X"99",X"A7",X"28",X"0C",X"3A",X"80",X"9A",X"E6",X"03",
		X"87",X"87",X"C6",X"10",X"32",X"00",X"9C",X"3A",X"05",X"99",X"A7",X"28",X"0C",X"3A",X"A1",X"9A",
		X"E6",X"03",X"87",X"87",X"C6",X"24",X"32",X"02",X"9C",X"3A",X"06",X"99",X"A7",X"28",X"0C",X"3A",
		X"C1",X"9A",X"E6",X"03",X"87",X"87",X"C6",X"24",X"32",X"04",X"9C",X"3A",X"07",X"99",X"A7",X"28",
		X"0C",X"3A",X"E1",X"9A",X"E6",X"03",X"87",X"87",X"C6",X"24",X"32",X"06",X"9C",X"3A",X"61",X"98",
		X"2F",X"C6",X"F9",X"32",X"10",X"9C",X"3A",X"6C",X"98",X"2F",X"C6",X"19",X"32",X"01",X"9C",X"3A",
		X"11",X"9C",X"38",X"07",X"E6",X"7F",X"32",X"11",X"9C",X"18",X"05",X"F6",X"80",X"32",X"11",X"9C",
		X"3A",X"64",X"98",X"2F",X"C6",X"F9",X"32",X"12",X"9C",X"3A",X"6D",X"98",X"2F",X"C6",X"19",X"32",
		X"03",X"9C",X"3A",X"13",X"9C",X"38",X"07",X"E6",X"7F",X"32",X"13",X"9C",X"18",X"05",X"F6",X"80",
		X"32",X"13",X"9C",X"3A",X"67",X"98",X"2F",X"C6",X"F9",X"32",X"14",X"9C",X"3A",X"6E",X"98",X"2F",
		X"C6",X"19",X"32",X"05",X"9C",X"3A",X"15",X"9C",X"38",X"07",X"E6",X"7F",X"32",X"15",X"9C",X"18",
		X"05",X"F6",X"80",X"32",X"15",X"9C",X"3A",X"6A",X"98",X"2F",X"C6",X"F9",X"32",X"16",X"9C",X"3A",
		X"6F",X"98",X"2F",X"C6",X"19",X"32",X"07",X"9C",X"3A",X"17",X"9C",X"38",X"07",X"E6",X"7F",X"32",
		X"17",X"9C",X"18",X"05",X"F6",X"80",X"32",X"17",X"9C",X"C9",X"DD",X"21",X"74",X"98",X"FD",X"21",
		X"24",X"9C",X"06",X"06",X"CD",X"5C",X"25",X"FD",X"23",X"DD",X"23",X"CD",X"5C",X"25",X"FD",X"23",
		X"DD",X"23",X"CD",X"9D",X"25",X"FD",X"23",X"DD",X"23",X"10",X"F7",X"C9",X"DD",X"7E",X"00",X"A7",
		X"28",X"37",X"3A",X"2F",X"99",X"A7",X"28",X"19",X"DD",X"7E",X"10",X"2F",X"C6",X"FF",X"FD",X"77",
		X"10",X"DD",X"7E",X"20",X"2F",X"C6",X"1F",X"FD",X"77",X"00",X"38",X"18",X"FD",X"36",X"20",X"0C",
		X"C9",X"DD",X"7E",X"10",X"FD",X"77",X"10",X"DD",X"7E",X"20",X"C6",X"FE",X"FD",X"77",X"00",X"FD",
		X"36",X"20",X"0C",X"C9",X"FD",X"36",X"20",X"04",X"C9",X"FD",X"77",X"10",X"C9",X"DD",X"7E",X"00",
		X"A7",X"28",X"37",X"3A",X"2F",X"99",X"A7",X"28",X"19",X"DD",X"7E",X"10",X"2F",X"C6",X"FF",X"FD",
		X"77",X"10",X"DD",X"7E",X"20",X"2F",X"C6",X"1F",X"FD",X"77",X"00",X"38",X"18",X"FD",X"36",X"20",
		X"08",X"C9",X"DD",X"7E",X"10",X"FD",X"77",X"10",X"DD",X"7E",X"20",X"C6",X"FE",X"FD",X"77",X"00",
		X"FD",X"36",X"20",X"08",X"C9",X"FD",X"36",X"20",X"00",X"C9",X"FD",X"77",X"10",X"C9",X"3A",X"04",
		X"99",X"A7",X"C8",X"CD",X"06",X"2D",X"3A",X"17",X"98",X"A7",X"C2",X"6D",X"26",X"3A",X"62",X"98",
		X"21",X"60",X"98",X"86",X"77",X"D0",X"21",X"8A",X"9A",X"11",X"8B",X"9A",X"01",X"0B",X"00",X"ED",
		X"B8",X"21",X"15",X"9B",X"11",X"17",X"9B",X"01",X"16",X"00",X"ED",X"B8",X"3A",X"16",X"98",X"4F",
		X"21",X"80",X"9A",X"96",X"E6",X"03",X"28",X"06",X"FE",X"02",X"28",X"73",X"18",X"29",X"79",X"21",
		X"DD",X"26",X"DF",X"2A",X"00",X"9B",X"19",X"7E",X"FE",X"EC",X"30",X"10",X"FE",X"E8",X"30",X"7A",
		X"22",X"00",X"9B",X"3A",X"80",X"9A",X"E6",X"03",X"32",X"80",X"9A",X"C9",X"3E",X"00",X"32",X"60",
		X"98",X"3E",X"FF",X"32",X"17",X"98",X"C9",X"79",X"21",X"DD",X"26",X"DF",X"2A",X"00",X"9B",X"19",
		X"7E",X"FE",X"E8",X"3A",X"80",X"9A",X"30",X"C7",X"22",X"00",X"9B",X"3A",X"80",X"9A",X"E6",X"03",
		X"87",X"87",X"81",X"C6",X"04",X"32",X"81",X"9A",X"79",X"32",X"80",X"9A",X"C9",X"3A",X"16",X"98",
		X"4F",X"21",X"80",X"9A",X"96",X"E6",X"03",X"C8",X"E6",X"01",X"28",X"13",X"79",X"21",X"DD",X"26",
		X"DF",X"2A",X"00",X"9B",X"19",X"7E",X"FE",X"E8",X"D0",X"AF",X"32",X"17",X"98",X"18",X"C9",X"AF",
		X"32",X"60",X"98",X"32",X"17",X"98",X"2A",X"04",X"9B",X"22",X"00",X"9B",X"3A",X"80",X"9A",X"C6",
		X"02",X"E6",X"03",X"32",X"80",X"9A",X"32",X"81",X"9A",X"C9",X"D6",X"EC",X"E6",X"03",X"4F",X"3A",
		X"80",X"9A",X"E6",X"03",X"87",X"87",X"81",X"21",X"E5",X"26",X"CF",X"7E",X"4F",X"21",X"DD",X"26",
		X"DF",X"2A",X"00",X"9B",X"19",X"7E",X"FE",X"E8",X"30",X"02",X"18",X"8C",X"79",X"C6",X"02",X"E6",
		X"03",X"4F",X"21",X"DD",X"26",X"DF",X"2A",X"00",X"9B",X"19",X"C3",X"58",X"26",X"E0",X"FF",X"01",
		X"00",X"20",X"00",X"FF",X"FF",X"01",X"01",X"03",X"03",X"00",X"02",X"00",X"02",X"01",X"01",X"03",
		X"03",X"00",X"02",X"00",X"02",X"3A",X"05",X"99",X"A7",X"C8",X"3A",X"D1",X"98",X"A7",X"C2",X"77",
		X"28",X"3A",X"65",X"98",X"21",X"63",X"98",X"86",X"77",X"D0",X"21",X"AA",X"9A",X"11",X"AB",X"9A",
		X"01",X"0B",X"00",X"ED",X"B8",X"21",X"55",X"9B",X"11",X"57",X"9B",X"01",X"16",X"00",X"ED",X"B8",
		X"3A",X"C0",X"98",X"E6",X"1F",X"47",X"3A",X"40",X"9B",X"E6",X"1F",X"90",X"32",X"41",X"98",X"3E",
		X"03",X"30",X"02",X"3E",X"01",X"32",X"42",X"98",X"2A",X"C0",X"98",X"29",X"29",X"29",X"7C",X"E6",
		X"1F",X"47",X"2A",X"40",X"9B",X"29",X"29",X"29",X"7C",X"E6",X"1F",X"90",X"32",X"43",X"98",X"3E",
		X"00",X"30",X"02",X"3E",X"02",X"32",X"44",X"98",X"3A",X"A0",X"9A",X"E6",X"03",X"4F",X"21",X"DD",
		X"26",X"DF",X"2A",X"40",X"9B",X"19",X"22",X"50",X"98",X"7E",X"FE",X"E8",X"30",X"3C",X"CD",X"A5",
		X"2F",X"E6",X"07",X"28",X"4A",X"21",X"08",X"99",X"BE",X"D2",X"13",X"28",X"3A",X"41",X"98",X"A7",
		X"20",X"05",X"3A",X"44",X"98",X"18",X"0A",X"3A",X"43",X"98",X"A7",X"C2",X"42",X"28",X"3A",X"42",
		X"98",X"47",X"CD",X"A5",X"2F",X"E6",X"0F",X"FE",X"02",X"38",X"78",X"79",X"90",X"E6",X"03",X"28",
		X"7B",X"E6",X"01",X"28",X"1A",X"48",X"79",X"C3",X"4E",X"28",X"CD",X"A5",X"2F",X"E6",X"01",X"28",
		X"0E",X"79",X"E6",X"01",X"3A",X"42",X"98",X"28",X"03",X"3A",X"44",X"98",X"4F",X"18",X"09",X"CD",
		X"A5",X"2F",X"F6",X"01",X"81",X"E6",X"03",X"4F",X"21",X"DD",X"26",X"DF",X"2A",X"40",X"9B",X"19",
		X"7E",X"FE",X"E8",X"30",X"18",X"79",X"32",X"A0",X"9A",X"22",X"40",X"9B",X"21",X"A1",X"9A",X"7E",
		X"E6",X"03",X"87",X"87",X"81",X"C6",X"04",X"77",X"AF",X"32",X"71",X"98",X"C9",X"79",X"C6",X"02",
		X"E6",X"03",X"4F",X"21",X"DD",X"26",X"DF",X"2A",X"40",X"9B",X"19",X"7E",X"FE",X"E8",X"38",X"D5",
		X"3A",X"A0",X"9A",X"E6",X"03",X"4F",X"21",X"DD",X"26",X"DF",X"2A",X"40",X"9B",X"19",X"7E",X"FE",
		X"E8",X"30",X"4B",X"CD",X"A5",X"2F",X"E6",X"1F",X"28",X"10",X"18",X"13",X"CD",X"39",X"34",X"CD",
		X"A5",X"2F",X"E6",X"07",X"21",X"09",X"99",X"BE",X"30",X"05",X"3E",X"FF",X"32",X"71",X"98",X"2A",
		X"50",X"98",X"22",X"40",X"9B",X"C9",X"79",X"E6",X"01",X"78",X"20",X"03",X"3A",X"41",X"98",X"4F",
		X"18",X"86",X"79",X"E6",X"01",X"3A",X"42",X"98",X"28",X"03",X"3A",X"44",X"98",X"4F",X"21",X"DD",
		X"26",X"DF",X"2A",X"40",X"9B",X"19",X"7E",X"FE",X"E8",X"DA",X"D5",X"27",X"18",X"B5",X"3E",X"80",
		X"32",X"63",X"98",X"3E",X"F0",X"32",X"D1",X"98",X"21",X"00",X"03",X"22",X"15",X"99",X"22",X"1A",
		X"99",X"CD",X"F3",X"33",X"C3",X"FE",X"30",X"21",X"D1",X"98",X"35",X"20",X"16",X"21",X"05",X"99",
		X"7E",X"32",X"91",X"98",X"36",X"00",X"3E",X"40",X"32",X"81",X"98",X"CD",X"BF",X"31",X"C8",X"32",
		X"B1",X"98",X"C9",X"7E",X"0F",X"E6",X"07",X"21",X"A0",X"28",X"CF",X"7E",X"32",X"63",X"98",X"C9",
		X"C0",X"C0",X"A0",X"A0",X"80",X"80",X"60",X"60",X"3A",X"06",X"99",X"A7",X"C8",X"3A",X"D2",X"98",
		X"A7",X"C2",X"1E",X"2A",X"3A",X"68",X"98",X"21",X"66",X"98",X"86",X"77",X"D0",X"21",X"CA",X"9A",
		X"11",X"CB",X"9A",X"01",X"0B",X"00",X"ED",X"B8",X"21",X"95",X"9B",X"11",X"97",X"9B",X"01",X"16",
		X"00",X"ED",X"B8",X"3A",X"C0",X"98",X"E6",X"1F",X"47",X"3A",X"80",X"9B",X"E6",X"1F",X"90",X"32",
		X"41",X"98",X"3E",X"03",X"30",X"02",X"3E",X"01",X"32",X"42",X"98",X"2A",X"C0",X"98",X"29",X"29",
		X"29",X"7C",X"E6",X"1F",X"47",X"2A",X"80",X"9B",X"29",X"29",X"29",X"7C",X"E6",X"1F",X"90",X"32",
		X"43",X"98",X"3E",X"00",X"30",X"02",X"3E",X"02",X"32",X"44",X"98",X"3A",X"C0",X"9A",X"E6",X"03",
		X"4F",X"21",X"DD",X"26",X"DF",X"2A",X"80",X"9B",X"19",X"22",X"50",X"98",X"7E",X"FE",X"E8",X"30",
		X"3C",X"CD",X"A5",X"2F",X"E6",X"07",X"28",X"4A",X"21",X"08",X"99",X"BE",X"D2",X"C6",X"29",X"3A",
		X"41",X"98",X"A7",X"20",X"05",X"3A",X"44",X"98",X"18",X"0A",X"3A",X"43",X"98",X"A7",X"C2",X"F5",
		X"29",X"3A",X"42",X"98",X"47",X"CD",X"A5",X"2F",X"E6",X"0F",X"FE",X"08",X"38",X"78",X"79",X"90",
		X"E6",X"03",X"28",X"7B",X"E6",X"01",X"28",X"1A",X"48",X"79",X"C3",X"01",X"2A",X"CD",X"A5",X"2F",
		X"E6",X"01",X"28",X"0E",X"79",X"E6",X"01",X"3A",X"42",X"98",X"28",X"03",X"3A",X"44",X"98",X"4F",
		X"18",X"09",X"CD",X"A5",X"2F",X"F6",X"01",X"81",X"E6",X"03",X"4F",X"21",X"DD",X"26",X"DF",X"2A",
		X"80",X"9B",X"19",X"7E",X"FE",X"E8",X"30",X"18",X"79",X"32",X"C0",X"9A",X"22",X"80",X"9B",X"21",
		X"C1",X"9A",X"7E",X"E6",X"03",X"87",X"87",X"81",X"C6",X"04",X"77",X"AF",X"32",X"72",X"98",X"C9",
		X"79",X"C6",X"02",X"E6",X"03",X"4F",X"21",X"DD",X"26",X"DF",X"2A",X"80",X"9B",X"19",X"7E",X"FE",
		X"E8",X"38",X"D5",X"3A",X"C0",X"9A",X"E6",X"03",X"4F",X"21",X"DD",X"26",X"DF",X"2A",X"80",X"9B",
		X"19",X"7E",X"FE",X"E8",X"30",X"4B",X"CD",X"A5",X"2F",X"E6",X"1F",X"28",X"10",X"18",X"13",X"CD",
		X"39",X"34",X"CD",X"A5",X"2F",X"E6",X"07",X"21",X"09",X"99",X"BE",X"30",X"05",X"3E",X"FF",X"32",
		X"72",X"98",X"2A",X"50",X"98",X"22",X"80",X"9B",X"C9",X"79",X"E6",X"01",X"78",X"20",X"03",X"3A",
		X"41",X"98",X"4F",X"18",X"86",X"79",X"E6",X"01",X"3A",X"42",X"98",X"28",X"03",X"3A",X"44",X"98",
		X"4F",X"21",X"DD",X"26",X"DF",X"2A",X"80",X"9B",X"19",X"7E",X"FE",X"E8",X"DA",X"88",X"29",X"18",
		X"B5",X"3E",X"80",X"32",X"66",X"98",X"3E",X"F0",X"32",X"D2",X"98",X"C3",X"68",X"28",X"21",X"D2",
		X"98",X"35",X"20",X"16",X"21",X"06",X"99",X"7E",X"32",X"92",X"98",X"36",X"00",X"3E",X"40",X"32",
		X"82",X"98",X"CD",X"BF",X"31",X"C8",X"32",X"B2",X"98",X"C9",X"7E",X"0F",X"E6",X"07",X"21",X"A0",
		X"28",X"CF",X"7E",X"32",X"66",X"98",X"C9",X"3A",X"07",X"99",X"A7",X"C8",X"3A",X"D3",X"98",X"A7",
		X"C2",X"BD",X"2B",X"3A",X"6B",X"98",X"21",X"69",X"98",X"86",X"77",X"D0",X"21",X"EA",X"9A",X"11",
		X"EB",X"9A",X"01",X"0B",X"00",X"ED",X"B8",X"21",X"D5",X"9B",X"11",X"D7",X"9B",X"01",X"16",X"00",
		X"ED",X"B8",X"3A",X"C0",X"98",X"E6",X"1F",X"47",X"3A",X"C0",X"9B",X"E6",X"1F",X"90",X"32",X"41",
		X"98",X"3E",X"03",X"30",X"02",X"3E",X"01",X"32",X"42",X"98",X"2A",X"C0",X"98",X"29",X"29",X"29",
		X"7C",X"E6",X"1F",X"47",X"2A",X"C0",X"9B",X"29",X"29",X"29",X"7C",X"E6",X"1F",X"90",X"32",X"43",
		X"98",X"3E",X"00",X"30",X"02",X"3E",X"02",X"32",X"44",X"98",X"3A",X"E0",X"9A",X"E6",X"03",X"4F",
		X"21",X"DD",X"26",X"DF",X"2A",X"C0",X"9B",X"19",X"22",X"50",X"98",X"7E",X"FE",X"E8",X"30",X"3C",
		X"CD",X"A5",X"2F",X"E6",X"07",X"28",X"4A",X"21",X"08",X"99",X"BE",X"D2",X"65",X"2B",X"3A",X"41",
		X"98",X"A7",X"20",X"05",X"3A",X"44",X"98",X"18",X"0A",X"3A",X"43",X"98",X"A7",X"C2",X"94",X"2B",
		X"3A",X"42",X"98",X"47",X"CD",X"A5",X"2F",X"E6",X"0F",X"FE",X"0C",X"38",X"78",X"79",X"90",X"E6",
		X"03",X"28",X"7B",X"E6",X"01",X"28",X"1A",X"48",X"79",X"C3",X"A0",X"2B",X"CD",X"A5",X"2F",X"E6",
		X"01",X"28",X"0E",X"79",X"E6",X"01",X"3A",X"42",X"98",X"28",X"03",X"3A",X"44",X"98",X"4F",X"18",
		X"09",X"CD",X"A5",X"2F",X"F6",X"01",X"81",X"E6",X"03",X"4F",X"21",X"DD",X"26",X"DF",X"2A",X"C0",
		X"9B",X"19",X"7E",X"FE",X"E8",X"30",X"18",X"79",X"32",X"E0",X"9A",X"22",X"C0",X"9B",X"21",X"E1",
		X"9A",X"7E",X"E6",X"03",X"87",X"87",X"81",X"C6",X"04",X"77",X"AF",X"32",X"73",X"98",X"C9",X"79",
		X"C6",X"02",X"E6",X"03",X"4F",X"21",X"DD",X"26",X"DF",X"2A",X"C0",X"9B",X"19",X"7E",X"FE",X"E8",
		X"38",X"D5",X"3A",X"E0",X"9A",X"E6",X"03",X"4F",X"21",X"DD",X"26",X"DF",X"2A",X"C0",X"9B",X"19",
		X"7E",X"FE",X"E8",X"30",X"4B",X"CD",X"A5",X"2F",X"E6",X"1F",X"28",X"10",X"18",X"13",X"CD",X"39",
		X"34",X"CD",X"A5",X"2F",X"E6",X"07",X"21",X"09",X"99",X"BE",X"30",X"05",X"3E",X"FF",X"32",X"73",
		X"98",X"2A",X"50",X"98",X"22",X"C0",X"9B",X"C9",X"79",X"E6",X"01",X"78",X"20",X"03",X"3A",X"41",
		X"98",X"4F",X"18",X"86",X"79",X"E6",X"01",X"3A",X"42",X"98",X"28",X"03",X"3A",X"44",X"98",X"4F",
		X"21",X"DD",X"26",X"DF",X"2A",X"C0",X"9B",X"19",X"7E",X"FE",X"E8",X"DA",X"27",X"2B",X"18",X"B5",
		X"3E",X"80",X"32",X"69",X"98",X"3E",X"F0",X"32",X"D3",X"98",X"C3",X"68",X"28",X"21",X"D3",X"98",
		X"35",X"20",X"16",X"21",X"07",X"99",X"7E",X"32",X"93",X"98",X"36",X"00",X"3E",X"40",X"32",X"83",
		X"98",X"CD",X"BF",X"31",X"C8",X"32",X"B3",X"98",X"C9",X"7E",X"0F",X"E6",X"07",X"21",X"A0",X"28",
		X"CF",X"7E",X"32",X"69",X"98",X"C9",X"3A",X"04",X"99",X"A7",X"C8",X"3A",X"62",X"98",X"21",X"60",
		X"98",X"86",X"77",X"D0",X"21",X"8A",X"9A",X"11",X"8B",X"9A",X"01",X"0B",X"00",X"ED",X"B8",X"21",
		X"15",X"9B",X"11",X"17",X"9B",X"01",X"16",X"00",X"ED",X"B8",X"3A",X"80",X"9A",X"E6",X"03",X"4F",
		X"21",X"DD",X"26",X"DF",X"2A",X"00",X"9B",X"19",X"22",X"50",X"98",X"7E",X"FE",X"E8",X"30",X"79",
		X"CD",X"A5",X"2F",X"E6",X"07",X"FE",X"01",X"38",X"70",X"3A",X"05",X"99",X"A7",X"28",X"05",X"2A",
		X"C6",X"98",X"18",X"0E",X"3A",X"06",X"99",X"A7",X"28",X"05",X"2A",X"CA",X"98",X"18",X"03",X"2A",
		X"CE",X"98",X"22",X"58",X"98",X"3A",X"58",X"98",X"E6",X"1F",X"47",X"3A",X"00",X"9B",X"E6",X"1F",
		X"90",X"28",X"1C",X"06",X"03",X"30",X"02",X"06",X"01",X"2A",X"58",X"98",X"7D",X"E6",X"E0",X"6F",
		X"ED",X"5B",X"00",X"9B",X"7B",X"E6",X"E0",X"5F",X"ED",X"52",X"C2",X"EE",X"2C",X"18",X"17",X"2A",
		X"58",X"98",X"7D",X"E6",X"E0",X"6F",X"ED",X"5B",X"00",X"9B",X"7B",X"E6",X"E0",X"5F",X"ED",X"52",
		X"06",X"02",X"30",X"02",X"06",X"00",X"3E",X"FF",X"32",X"70",X"98",X"79",X"90",X"E6",X"03",X"28",
		X"5D",X"E6",X"01",X"28",X"04",X"48",X"79",X"18",X"0D",X"AF",X"32",X"70",X"98",X"CD",X"A5",X"2F",
		X"F6",X"01",X"81",X"E6",X"03",X"4F",X"21",X"DD",X"26",X"DF",X"2A",X"00",X"9B",X"19",X"7E",X"FE",
		X"E8",X"30",X"14",X"79",X"32",X"80",X"9A",X"22",X"00",X"9B",X"21",X"81",X"9A",X"7E",X"E6",X"03",
		X"87",X"87",X"81",X"C6",X"04",X"77",X"C9",X"79",X"C6",X"02",X"E6",X"03",X"4F",X"21",X"DD",X"26",
		X"DF",X"2A",X"00",X"9B",X"19",X"7E",X"FE",X"E8",X"38",X"D9",X"3A",X"80",X"9A",X"E6",X"03",X"4F",
		X"21",X"DD",X"26",X"DF",X"2A",X"00",X"9B",X"19",X"7E",X"FE",X"E8",X"D2",X"8F",X"26",X"2A",X"50",
		X"98",X"22",X"00",X"9B",X"C9",X"CD",X"A5",X"2F",X"E6",X"0F",X"20",X"08",X"CD",X"A5",X"2F",X"E6",
		X"03",X"3C",X"4F",X"C9",X"AF",X"C9",X"3A",X"2F",X"99",X"A7",X"28",X"29",X"0E",X"04",X"3A",X"05",
		X"98",X"CB",X"7F",X"20",X"17",X"0D",X"3A",X"03",X"98",X"CB",X"6F",X"20",X"0F",X"0D",X"3A",X"04",
		X"98",X"CB",X"47",X"20",X"07",X"0D",X"3A",X"03",X"98",X"CB",X"67",X"C8",X"79",X"3D",X"32",X"16",
		X"98",X"3E",X"FF",X"A7",X"C9",X"0E",X"04",X"3A",X"04",X"98",X"CB",X"4F",X"20",X"17",X"0D",X"3A",
		X"04",X"98",X"CB",X"67",X"20",X"0F",X"0D",X"3A",X"03",X"98",X"CB",X"47",X"20",X"07",X"0D",X"3A",
		X"04",X"98",X"CB",X"6F",X"C8",X"79",X"3D",X"32",X"16",X"98",X"3E",X"FF",X"A7",X"C9",X"21",X"50",
		X"9C",X"7E",X"A7",X"C8",X"47",X"36",X"00",X"3E",X"20",X"2C",X"2C",X"5E",X"2C",X"56",X"12",X"10",
		X"F9",X"C9",X"21",X"00",X"9D",X"34",X"08",X"7E",X"87",X"87",X"6F",X"73",X"2C",X"72",X"2C",X"08",
		X"77",X"2C",X"EB",X"C9",X"3A",X"00",X"9D",X"A7",X"C8",X"47",X"21",X"04",X"9D",X"AF",X"32",X"00",
		X"9D",X"5E",X"2C",X"56",X"2C",X"7E",X"12",X"2C",X"CB",X"DA",X"7E",X"12",X"2C",X"10",X"F2",X"C9",
		X"3A",X"04",X"99",X"A7",X"C8",X"32",X"40",X"98",X"21",X"99",X"2F",X"11",X"48",X"98",X"01",X"03",
		X"00",X"ED",X"B0",X"21",X"05",X"9B",X"87",X"CF",X"E5",X"DD",X"E1",X"3A",X"40",X"98",X"21",X"80",
		X"9A",X"CF",X"E5",X"FD",X"E1",X"3A",X"60",X"98",X"07",X"07",X"07",X"E6",X"07",X"32",X"41",X"98",
		X"21",X"11",X"9C",X"22",X"54",X"98",X"CD",X"A5",X"2E",X"21",X"56",X"98",X"11",X"C0",X"98",X"01",
		X"04",X"00",X"ED",X"B0",X"C9",X"3A",X"05",X"99",X"A7",X"C8",X"32",X"40",X"98",X"CD",X"7B",X"2F",
		X"3A",X"40",X"98",X"21",X"45",X"9B",X"87",X"CF",X"E5",X"DD",X"E1",X"3A",X"40",X"98",X"21",X"A0",
		X"9A",X"CF",X"E5",X"FD",X"E1",X"3A",X"63",X"98",X"07",X"07",X"07",X"E6",X"07",X"32",X"41",X"98",
		X"21",X"13",X"9C",X"22",X"54",X"98",X"CD",X"A5",X"2E",X"21",X"56",X"98",X"11",X"C4",X"98",X"01",
		X"04",X"00",X"ED",X"B0",X"C9",X"3A",X"06",X"99",X"A7",X"C8",X"32",X"40",X"98",X"CD",X"7B",X"2F",
		X"3A",X"40",X"98",X"21",X"85",X"9B",X"87",X"CF",X"E5",X"DD",X"E1",X"3A",X"40",X"98",X"21",X"C0",
		X"9A",X"CF",X"E5",X"FD",X"E1",X"3A",X"66",X"98",X"07",X"07",X"07",X"E6",X"07",X"32",X"41",X"98",
		X"21",X"15",X"9C",X"22",X"54",X"98",X"CD",X"A5",X"2E",X"21",X"56",X"98",X"11",X"C8",X"98",X"01",
		X"04",X"00",X"ED",X"B0",X"C9",X"3A",X"07",X"99",X"A7",X"C8",X"32",X"40",X"98",X"CD",X"7B",X"2F",
		X"3A",X"40",X"98",X"21",X"C5",X"9B",X"87",X"CF",X"E5",X"DD",X"E1",X"3A",X"40",X"98",X"21",X"E0",
		X"9A",X"CF",X"E5",X"FD",X"E1",X"3A",X"69",X"98",X"07",X"07",X"07",X"E6",X"07",X"32",X"41",X"98",
		X"21",X"17",X"9C",X"22",X"54",X"98",X"CD",X"A5",X"2E",X"21",X"56",X"98",X"11",X"CC",X"98",X"01",
		X"04",X"00",X"ED",X"B0",X"C9",X"3A",X"48",X"98",X"2A",X"54",X"98",X"CB",X"7E",X"77",X"28",X"02",
		X"CB",X"FE",X"DD",X"56",X"00",X"DD",X"2B",X"DD",X"5E",X"00",X"DD",X"2B",X"21",X"50",X"9C",X"34",
		X"7E",X"87",X"85",X"6F",X"73",X"2C",X"72",X"DD",X"56",X"00",X"DD",X"2B",X"DD",X"5E",X"00",X"DD",
		X"2B",X"21",X"50",X"9C",X"34",X"7E",X"87",X"85",X"6F",X"73",X"2C",X"72",X"21",X"40",X"98",X"35",
		X"20",X"13",X"DD",X"66",X"00",X"DD",X"6E",X"FF",X"22",X"56",X"98",X"DD",X"66",X"FE",X"DD",X"6E",
		X"FD",X"22",X"58",X"98",X"C9",X"DD",X"56",X"00",X"DD",X"2B",X"DD",X"5E",X"00",X"DD",X"2B",X"FD",
		X"7E",X"00",X"FD",X"2B",X"ED",X"53",X"56",X"98",X"21",X"28",X"3F",X"85",X"6F",X"46",X"25",X"3A",
		X"41",X"98",X"86",X"CD",X"72",X"2D",X"3A",X"4A",X"98",X"B0",X"12",X"DD",X"66",X"00",X"DD",X"6E",
		X"FF",X"22",X"58",X"98",X"DD",X"56",X"00",X"DD",X"2B",X"DD",X"5E",X"00",X"DD",X"2B",X"FD",X"7E",
		X"00",X"FD",X"2B",X"21",X"14",X"3F",X"85",X"6F",X"46",X"25",X"3A",X"41",X"98",X"86",X"CD",X"72",
		X"2D",X"3A",X"4A",X"98",X"B0",X"12",X"3A",X"40",X"98",X"3D",X"28",X"29",X"47",X"C5",X"DD",X"56",
		X"00",X"DD",X"2B",X"DD",X"5E",X"00",X"DD",X"2B",X"FD",X"7E",X"00",X"FD",X"2B",X"21",X"00",X"3F",
		X"85",X"6F",X"46",X"25",X"3A",X"41",X"98",X"86",X"CD",X"72",X"2D",X"3A",X"4A",X"98",X"B0",X"12",
		X"78",X"C1",X"10",X"D9",X"47",X"3A",X"49",X"98",X"B0",X"12",X"C9",X"21",X"04",X"99",X"BE",X"28",
		X"07",X"30",X"0A",X"21",X"9C",X"2F",X"18",X"08",X"21",X"9F",X"2F",X"18",X"03",X"21",X"A2",X"2F",
		X"11",X"48",X"98",X"01",X"03",X"00",X"ED",X"B0",X"C9",X"2B",X"06",X"30",X"0F",X"02",X"10",X"16",
		X"03",X"18",X"0A",X"01",X"08",X"D9",X"21",X"0F",X"9E",X"11",X"10",X"9E",X"01",X"10",X"00",X"ED",
		X"B8",X"21",X"10",X"9E",X"3A",X"07",X"9E",X"AE",X"32",X"00",X"9E",X"21",X"02",X"98",X"86",X"D9",
		X"C9",X"D9",X"3A",X"03",X"98",X"0F",X"0F",X"0F",X"21",X"22",X"99",X"CB",X"16",X"7E",X"E6",X"07",
		X"FE",X"01",X"C0",X"CD",X"A1",X"33",X"3E",X"01",X"C3",X"3E",X"30",X"3A",X"03",X"98",X"21",X"27",
		X"99",X"07",X"07",X"CB",X"16",X"7E",X"E6",X"07",X"FE",X"01",X"C0",X"EB",X"CD",X"A1",X"33",X"21",
		X"30",X"99",X"34",X"EB",X"23",X"7E",X"C6",X"10",X"77",X"47",X"23",X"7E",X"90",X"D0",X"7E",X"4F",
		X"E6",X"F0",X"C6",X"10",X"2B",X"ED",X"44",X"86",X"77",X"79",X"E6",X"0F",X"18",X"30",X"3A",X"03",
		X"98",X"21",X"24",X"99",X"07",X"CB",X"16",X"7E",X"E6",X"07",X"FE",X"01",X"C0",X"EB",X"CD",X"A1",
		X"33",X"21",X"2A",X"99",X"34",X"EB",X"23",X"7E",X"C6",X"10",X"77",X"47",X"23",X"7E",X"90",X"D0",
		X"7E",X"4F",X"E6",X"F0",X"C6",X"10",X"2B",X"ED",X"44",X"86",X"77",X"79",X"E6",X"0F",X"21",X"23",
		X"99",X"86",X"27",X"77",X"30",X"02",X"36",X"99",X"11",X"06",X"83",X"21",X"16",X"01",X"FF",X"21",
		X"BF",X"FF",X"19",X"EB",X"3A",X"23",X"99",X"CD",X"B1",X"30",X"21",X"06",X"8B",X"11",X"20",X"00",
		X"3E",X"A3",X"06",X"06",X"77",X"19",X"10",X"FC",X"C9",X"3A",X"2A",X"99",X"A7",X"C8",X"21",X"2B",
		X"99",X"7E",X"A7",X"20",X"07",X"36",X"30",X"3C",X"32",X"84",X"A1",X"C9",X"35",X"28",X"09",X"7E",
		X"FE",X"18",X"C0",X"AF",X"32",X"84",X"A1",X"C9",X"21",X"2A",X"99",X"35",X"C9",X"3A",X"30",X"99",
		X"A7",X"C8",X"21",X"31",X"99",X"7E",X"A7",X"20",X"07",X"36",X"30",X"3C",X"32",X"86",X"A1",X"C9",
		X"35",X"28",X"09",X"7E",X"FE",X"18",X"C0",X"AF",X"32",X"86",X"A1",X"C9",X"21",X"30",X"99",X"35",
		X"C9",X"FE",X"0A",X"4F",X"38",X"0F",X"4F",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"12",X"D7",X"79",
		X"E6",X"0F",X"12",X"D7",X"C9",X"3E",X"20",X"18",X"F4",X"4F",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",
		X"CD",X"D6",X"30",X"79",X"E6",X"0F",X"28",X"04",X"04",X"12",X"D7",X"C9",X"78",X"A7",X"28",X"03",
		X"AF",X"18",X"F6",X"3E",X"20",X"18",X"F2",X"7E",X"FE",X"40",X"C8",X"3E",X"20",X"12",X"23",X"D7",
		X"18",X"F5",X"CB",X"DA",X"7E",X"FE",X"40",X"C8",X"79",X"12",X"23",X"D7",X"18",X"F6",X"3A",X"20",
		X"99",X"FE",X"04",X"D0",X"3A",X"11",X"99",X"A7",X"20",X"79",X"FD",X"21",X"12",X"99",X"11",X"A2",
		X"80",X"21",X"78",X"01",X"FD",X"7E",X"03",X"FD",X"86",X"00",X"27",X"FD",X"77",X"00",X"FD",X"7E",
		X"04",X"FD",X"8E",X"01",X"27",X"FD",X"77",X"01",X"3E",X"00",X"FD",X"8E",X"02",X"27",X"FD",X"77",
		X"02",X"E6",X"0F",X"FE",X"02",X"28",X"0A",X"FE",X"07",X"28",X"06",X"AF",X"32",X"02",X"99",X"18",
		X"03",X"CD",X"9A",X"3E",X"DD",X"21",X"1C",X"99",X"FD",X"7E",X"02",X"DD",X"BE",X"02",X"38",X"49",
		X"28",X"02",X"18",X"14",X"FD",X"7E",X"01",X"DD",X"BE",X"01",X"38",X"3D",X"28",X"02",X"18",X"08",
		X"DD",X"7E",X"00",X"FD",X"BE",X"00",X"30",X"31",X"FD",X"7E",X"00",X"DD",X"77",X"00",X"FD",X"7E",
		X"01",X"DD",X"77",X"01",X"FD",X"7E",X"02",X"DD",X"77",X"02",X"D5",X"E5",X"CD",X"84",X"1A",X"E1",
		X"D1",X"18",X"16",X"FD",X"21",X"17",X"99",X"11",X"62",X"83",X"21",X"7C",X"01",X"18",X"85",X"FD",
		X"21",X"12",X"99",X"11",X"A2",X"80",X"21",X"78",X"01",X"FF",X"21",X"3F",X"FF",X"19",X"EB",X"FD",
		X"7E",X"02",X"06",X"00",X"CD",X"C9",X"30",X"FD",X"7E",X"01",X"CD",X"C9",X"30",X"FD",X"7E",X"00",
		X"C3",X"B6",X"30",X"FD",X"21",X"17",X"99",X"11",X"62",X"83",X"21",X"7C",X"01",X"18",X"DA",X"21",
		X"0F",X"99",X"7E",X"A7",X"C8",X"35",X"7E",X"FE",X"03",X"28",X"03",X"3E",X"40",X"C9",X"3E",X"40",
		X"32",X"B0",X"98",X"C9",X"3A",X"01",X"99",X"E6",X"03",X"06",X"9C",X"20",X"02",X"06",X"8E",X"21",
		X"B0",X"98",X"11",X"BB",X"8F",X"CD",X"FA",X"31",X"23",X"11",X"5B",X"8C",X"CD",X"FA",X"31",X"23",
		X"11",X"41",X"8C",X"CD",X"FA",X"31",X"23",X"11",X"A1",X"8F",X"7E",X"A7",X"C8",X"35",X"28",X"11",
		X"CB",X"56",X"3E",X"00",X"28",X"02",X"3E",X"87",X"E6",X"3F",X"4F",X"1A",X"E6",X"C0",X"B1",X"12",
		X"C9",X"78",X"18",X"F4",X"3A",X"04",X"99",X"A7",X"C8",X"3A",X"02",X"98",X"E6",X"3F",X"C0",X"CD",
		X"A5",X"2F",X"E6",X"07",X"FE",X"03",X"D0",X"FE",X"01",X"38",X"3C",X"28",X"1D",X"3A",X"07",X"99",
		X"A7",X"28",X"04",X"32",X"73",X"98",X"C9",X"3A",X"05",X"99",X"A7",X"28",X"04",X"32",X"71",X"98",
		X"C9",X"3A",X"06",X"99",X"A7",X"C8",X"32",X"72",X"98",X"C9",X"3A",X"06",X"99",X"A7",X"28",X"04",
		X"32",X"72",X"98",X"C9",X"3A",X"07",X"99",X"A7",X"28",X"04",X"32",X"73",X"98",X"C9",X"3A",X"05",
		X"99",X"A7",X"C8",X"32",X"71",X"98",X"C9",X"3A",X"05",X"99",X"A7",X"28",X"04",X"32",X"71",X"98",
		X"C9",X"3A",X"06",X"99",X"A7",X"28",X"04",X"32",X"72",X"98",X"C9",X"3A",X"07",X"99",X"A7",X"C8",
		X"32",X"73",X"98",X"C9",X"3A",X"01",X"99",X"E6",X"03",X"0E",X"1D",X"20",X"02",X"0E",X"0F",X"21",
		X"08",X"98",X"7E",X"47",X"34",X"87",X"87",X"87",X"6F",X"26",X"00",X"29",X"29",X"11",X"41",X"84",
		X"19",X"78",X"A7",X"CA",X"1D",X"33",X"FE",X"1B",X"CA",X"3E",X"33",X"E5",X"3A",X"01",X"99",X"3D",
		X"E6",X"07",X"21",X"43",X"34",X"DF",X"EB",X"11",X"0C",X"00",X"05",X"28",X"03",X"19",X"10",X"FD",
		X"EB",X"E1",X"36",X"F8",X"CB",X"DC",X"CB",X"F1",X"71",X"CB",X"9C",X"23",X"36",X"20",X"23",X"06",
		X"0C",X"CB",X"F9",X"CB",X"B1",X"1A",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"FE",X"0F",X"28",X"2D",
		X"C6",X"E8",X"77",X"CB",X"DC",X"FE",X"F5",X"28",X"2C",X"71",X"CB",X"9C",X"23",X"1A",X"E6",X"0F",
		X"FE",X"0F",X"28",X"1D",X"C6",X"E8",X"77",X"CB",X"DC",X"FE",X"F5",X"28",X"1C",X"71",X"CB",X"9C",
		X"23",X"13",X"10",X"D1",X"36",X"F8",X"CB",X"DC",X"71",X"3E",X"FF",X"A7",X"C9",X"3E",X"20",X"18",
		X"D1",X"3E",X"20",X"18",X"E1",X"36",X"BE",X"18",X"D1",X"36",X"BE",X"18",X"E1",X"CB",X"F1",X"36",
		X"FA",X"CB",X"DC",X"71",X"CB",X"9C",X"23",X"CB",X"B1",X"06",X"19",X"36",X"F9",X"CB",X"DC",X"71",
		X"CB",X"9C",X"23",X"10",X"F6",X"36",X"FA",X"CB",X"DC",X"71",X"3E",X"FF",X"A7",X"C9",X"36",X"FA",
		X"CB",X"DC",X"CB",X"F9",X"CB",X"F1",X"71",X"CB",X"9C",X"23",X"06",X"19",X"36",X"F9",X"CB",X"DC",
		X"71",X"CB",X"9C",X"23",X"10",X"F6",X"36",X"FA",X"CB",X"DC",X"CB",X"B1",X"71",X"AF",X"C9",X"21",
		X"F0",X"99",X"7E",X"A7",X"C8",X"35",X"F5",X"23",X"7E",X"CD",X"78",X"33",X"F1",X"C8",X"3D",X"06",
		X"00",X"4F",X"5D",X"54",X"23",X"ED",X"B0",X"C9",X"32",X"00",X"A1",X"3E",X"00",X"32",X"80",X"A1",
		X"00",X"00",X"00",X"00",X"3E",X"01",X"32",X"80",X"A1",X"C9",X"F5",X"FE",X"05",X"28",X"07",X"3A",
		X"20",X"99",X"FE",X"04",X"30",X"09",X"21",X"F0",X"99",X"34",X"7E",X"CF",X"F1",X"77",X"C9",X"F1",
		X"C9",X"3E",X"05",X"18",X"E5",X"3E",X"07",X"18",X"E1",X"3E",X"06",X"18",X"DD",X"AF",X"CD",X"8A",
		X"33",X"3E",X"02",X"CD",X"8A",X"33",X"3E",X"0F",X"C3",X"8A",X"33",X"3E",X"01",X"C3",X"8A",X"33",
		X"3E",X"81",X"C3",X"8A",X"33",X"3E",X"03",X"CD",X"8A",X"33",X"3E",X"08",X"CD",X"8A",X"33",X"3A",
		X"01",X"99",X"E6",X"03",X"C0",X"21",X"04",X"99",X"7E",X"A7",X"C8",X"FE",X"09",X"D0",X"34",X"7E",
		X"CD",X"4F",X"1E",X"32",X"62",X"98",X"C9",X"3E",X"09",X"18",X"9F",X"3E",X"0B",X"18",X"9B",X"3E",
		X"04",X"18",X"D9",X"3E",X"19",X"18",X"93",X"3E",X"0A",X"18",X"8F",X"3E",X"10",X"CD",X"8A",X"33",
		X"3E",X"11",X"CD",X"8A",X"33",X"3E",X"12",X"C3",X"8A",X"33",X"AF",X"32",X"18",X"9C",X"CD",X"8A",
		X"33",X"3E",X"13",X"CD",X"8A",X"33",X"3E",X"14",X"CD",X"8A",X"33",X"3E",X"15",X"C3",X"8A",X"33",
		X"3E",X"16",X"CD",X"8A",X"33",X"3E",X"17",X"CD",X"8A",X"33",X"3E",X"18",X"C3",X"8A",X"33",X"3E",
		X"0D",X"C3",X"8A",X"33",X"3E",X"0C",X"C3",X"8A",X"33",X"3A",X"04",X"99",X"A7",X"C8",X"3E",X"0E",
		X"C3",X"8A",X"33",X"53",X"34",X"53",X"34",X"8B",X"35",X"8B",X"35",X"C3",X"36",X"C3",X"36",X"FB",
		X"37",X"FB",X"37",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"24",
		X"44",X"0F",X"24",X"44",X"0F",X"20",X"F2",X"0F",X"24",X"44",X"0F",X"35",X"55",X"1F",X"35",X"55",
		X"1F",X"76",X"F3",X"1F",X"35",X"5B",X"6F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"76",X"FF",X"FF",
		X"FF",X"F7",X"6F",X"24",X"44",X"44",X"40",X"F2",X"44",X"A6",X"F2",X"0F",X"20",X"F7",X"6F",X"35",
		X"55",X"55",X"51",X"F3",X"55",X"51",X"F3",X"1F",X"31",X"F7",X"6F",X"DF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"6F",X"24",X"44",X"44",X"44",X"44",X"0F",X"24",X"44",X"44",
		X"40",X"F7",X"6F",X"35",X"55",X"55",X"55",X"5B",X"6F",X"35",X"55",X"55",X"B6",X"F3",X"1F",X"FF",
		X"FF",X"FF",X"FF",X"F7",X"6F",X"FF",X"FF",X"FF",X"76",X"FF",X"FF",X"24",X"44",X"0F",X"20",X"F7",
		X"6F",X"24",X"44",X"0F",X"76",X"F2",X"0F",X"35",X"55",X"1F",X"31",X"F3",X"1F",X"35",X"55",X"1F",
		X"31",X"F3",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"24",X"44",X"44",X"40",X"F2",
		X"0F",X"24",X"44",X"44",X"40",X"F2",X"0F",X"35",X"55",X"55",X"51",X"F7",X"6F",X"35",X"55",X"55",
		X"51",X"F7",X"6F",X"FF",X"FF",X"FF",X"FF",X"F7",X"6F",X"FF",X"FF",X"FF",X"FF",X"F7",X"6F",X"20",
		X"F2",X"0F",X"20",X"F7",X"6F",X"20",X"F2",X"0F",X"24",X"4A",X"6F",X"31",X"F3",X"1F",X"76",X"F3",
		X"1F",X"31",X"F7",X"6F",X"35",X"5B",X"6F",X"FF",X"FF",X"FF",X"76",X"FF",X"FF",X"FF",X"F7",X"6F",
		X"FF",X"F7",X"6F",X"24",X"44",X"0F",X"76",X"F2",X"44",X"40",X"F7",X"84",X"40",X"F7",X"6F",X"35",
		X"55",X"1F",X"76",X"F3",X"55",X"B6",X"F3",X"55",X"51",X"F3",X"1F",X"FF",X"FF",X"FF",X"76",X"FF",
		X"FF",X"76",X"FF",X"FF",X"FF",X"FF",X"FF",X"20",X"F2",X"44",X"A6",X"F2",X"0F",X"78",X"44",X"44",
		X"44",X"44",X"0F",X"31",X"F3",X"55",X"51",X"F3",X"1F",X"35",X"55",X"55",X"55",X"55",X"1F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"20",X"F2",X"44",X"44",X"44",X"0F",X"20",X"F2",X"44",
		X"40",X"F2",X"0F",X"76",X"F7",X"95",X"55",X"5B",X"6F",X"76",X"F3",X"55",X"51",X"F7",X"6F",X"76",
		X"F7",X"6F",X"FF",X"F7",X"6F",X"76",X"FF",X"FF",X"FF",X"F7",X"6F",X"76",X"F7",X"6F",X"20",X"F7",
		X"6F",X"76",X"F2",X"44",X"44",X"4A",X"6F",X"76",X"F7",X"6F",X"76",X"F7",X"6F",X"76",X"F7",X"95",
		X"55",X"55",X"1F",X"76",X"F7",X"6F",X"76",X"F7",X"6F",X"76",X"F7",X"6F",X"FF",X"FF",X"FF",X"76",
		X"F7",X"6F",X"76",X"F7",X"6F",X"76",X"F7",X"6F",X"24",X"44",X"0F",X"76",X"F3",X"1F",X"76",X"F7",
		X"6F",X"31",X"F7",X"6F",X"35",X"55",X"1F",X"76",X"FF",X"FF",X"76",X"F7",X"6F",X"FF",X"F7",X"6F",
		X"DF",X"FF",X"FF",X"78",X"44",X"44",X"A6",X"F7",X"6F",X"24",X"4A",X"6F",X"24",X"44",X"0F",X"35",
		X"55",X"55",X"51",X"F3",X"1F",X"35",X"55",X"1F",X"35",X"55",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"20",X"F2",X"0F",X"20",X"F2",X"0F",X"24",X"44",X"44",X"40",X"F2",X"0F",X"76",
		X"F7",X"6F",X"76",X"F7",X"6F",X"79",X"55",X"55",X"B6",X"F7",X"6F",X"76",X"F7",X"6F",X"76",X"F7",
		X"6F",X"76",X"FF",X"FF",X"76",X"F7",X"6F",X"76",X"F7",X"6F",X"76",X"F7",X"6F",X"76",X"F2",X"0F",
		X"76",X"F7",X"6F",X"76",X"F7",X"6F",X"76",X"F7",X"6F",X"31",X"F7",X"6F",X"31",X"F3",X"1F",X"76",
		X"F7",X"6F",X"76",X"F7",X"6F",X"FF",X"F7",X"6F",X"FF",X"FF",X"FF",X"76",X"F7",X"6F",X"76",X"F7",
		X"6F",X"24",X"4A",X"84",X"44",X"44",X"0F",X"31",X"F7",X"6F",X"31",X"F7",X"6F",X"35",X"55",X"55",
		X"55",X"55",X"1F",X"FF",X"F7",X"6F",X"FF",X"F7",X"6F",X"FF",X"FF",X"DF",X"FF",X"FF",X"FF",X"20",
		X"F7",X"84",X"44",X"4A",X"6F",X"24",X"44",X"0F",X"24",X"44",X"0F",X"31",X"F3",X"55",X"55",X"55",
		X"1F",X"35",X"55",X"1F",X"35",X"55",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"24",
		X"44",X"44",X"40",X"F2",X"0F",X"24",X"44",X"0F",X"20",X"F2",X"0F",X"79",X"55",X"55",X"51",X"F7",
		X"6F",X"35",X"55",X"1F",X"76",X"F3",X"1F",X"76",X"DF",X"FF",X"FF",X"F7",X"6F",X"FF",X"FF",X"FF",
		X"76",X"FF",X"FF",X"76",X"F2",X"0F",X"20",X"F7",X"6F",X"20",X"F2",X"44",X"A6",X"F2",X"0F",X"76",
		X"F3",X"1F",X"76",X"F7",X"6F",X"76",X"F3",X"55",X"51",X"F7",X"6F",X"76",X"FF",X"FF",X"76",X"F7",
		X"6F",X"76",X"FF",X"FF",X"FF",X"F7",X"6F",X"76",X"F2",X"44",X"A6",X"F7",X"6F",X"78",X"44",X"0F",
		X"20",X"F7",X"6F",X"76",X"F3",X"55",X"51",X"F7",X"6F",X"79",X"55",X"1F",X"76",X"F7",X"6F",X"76",
		X"FF",X"FF",X"FF",X"F7",X"6F",X"76",X"FF",X"FF",X"76",X"F7",X"6F",X"76",X"F2",X"44",X"44",X"4A",
		X"6F",X"76",X"F2",X"44",X"A6",X"F7",X"6F",X"31",X"F3",X"55",X"55",X"55",X"1F",X"31",X"F3",X"55",
		X"51",X"F3",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"20",X"F2",X"44",X"40",X"F2",
		X"0F",X"24",X"44",X"0F",X"24",X"44",X"0F",X"76",X"F3",X"55",X"B6",X"F7",X"6F",X"35",X"55",X"1F",
		X"35",X"5B",X"6F",X"76",X"FF",X"FF",X"76",X"F7",X"6F",X"FF",X"FF",X"FF",X"FF",X"F7",X"6F",X"76",
		X"F2",X"0F",X"76",X"F7",X"6F",X"20",X"F2",X"44",X"40",X"F7",X"6F",X"31",X"F7",X"6F",X"31",X"F3",
		X"1F",X"76",X"F3",X"55",X"51",X"F7",X"6F",X"FF",X"F7",X"6F",X"FF",X"FF",X"FF",X"76",X"FF",X"FF",
		X"FF",X"F7",X"6F",X"20",X"F7",X"84",X"44",X"44",X"0F",X"76",X"F2",X"44",X"40",X"F7",X"6F",X"31",
		X"F3",X"55",X"55",X"5B",X"6F",X"76",X"F3",X"55",X"51",X"F3",X"1F",X"FF",X"FF",X"FF",X"FF",X"F7",
		X"6F",X"76",X"FF",X"FF",X"FF",X"FF",X"FF",X"24",X"44",X"44",X"40",X"F7",X"6F",X"78",X"44",X"0F",
		X"24",X"44",X"0F",X"35",X"55",X"55",X"51",X"F3",X"1F",X"35",X"55",X"1F",X"35",X"55",X"1F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"20",X"F2",X"0F",X"20",X"F2",X"0F",X"20",X"F2",X"0F",
		X"20",X"F2",X"0F",X"31",X"F3",X"1F",X"31",X"F3",X"1F",X"31",X"F3",X"1F",X"31",X"F3",X"1F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"20",X"F2",X"0F",X"20",X"F2",
		X"0F",X"20",X"F2",X"0F",X"20",X"F2",X"0F",X"31",X"F3",X"1F",X"31",X"F3",X"1F",X"31",X"F3",X"1F",
		X"31",X"F3",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"20",
		X"F2",X"0F",X"20",X"F2",X"0F",X"20",X"F2",X"0F",X"20",X"F2",X"0F",X"31",X"F3",X"1F",X"31",X"F3",
		X"1F",X"31",X"F3",X"1F",X"31",X"F3",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"20",X"F2",X"0F",X"20",X"F2",X"0F",X"20",X"F2",X"0F",X"20",X"F2",X"0F",X"31",
		X"F3",X"1F",X"31",X"F3",X"1F",X"31",X"F3",X"1F",X"31",X"F3",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"20",X"F2",X"0F",X"20",X"F2",X"0F",X"20",X"F2",X"0F",X"20",X"F2",X"0F",X"31",
		X"F3",X"1F",X"31",X"F3",X"1F",X"31",X"F3",X"1F",X"31",X"F3",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"20",X"F2",X"0F",X"20",X"F2",X"0F",X"20",X"F2",X"0F",
		X"20",X"F2",X"0F",X"31",X"F3",X"1F",X"31",X"F3",X"1F",X"31",X"F3",X"1F",X"31",X"F3",X"1F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",X"FF",X"20",X"F2",X"0F",X"20",X"F2",
		X"0F",X"20",X"F2",X"0F",X"20",X"F2",X"0F",X"31",X"F3",X"1F",X"31",X"F3",X"1F",X"31",X"F3",X"1F",
		X"31",X"F3",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"20",
		X"F2",X"0F",X"20",X"F2",X"0F",X"20",X"F2",X"0F",X"20",X"F2",X"0F",X"31",X"F3",X"1F",X"31",X"F3",
		X"1F",X"31",X"F3",X"1F",X"31",X"F3",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"3A",X"1A",X"9C",X"A7",X"C8",X"3A",X"04",X"99",X"A7",X"C8",X"3A",X"19",X"98",
		X"A7",X"20",X"44",X"21",X"1A",X"9C",X"11",X"0B",X"9C",X"3A",X"10",X"9C",X"96",X"30",X"02",X"ED",
		X"44",X"FE",X"08",X"D0",X"47",X"EB",X"3A",X"01",X"9C",X"96",X"30",X"02",X"ED",X"44",X"FE",X"08",
		X"D0",X"CD",X"34",X"34",X"CD",X"D5",X"33",X"3E",X"40",X"32",X"19",X"98",X"3A",X"2F",X"99",X"A7",
		X"28",X"04",X"3E",X"34",X"18",X"02",X"3E",X"37",X"32",X"0A",X"9C",X"21",X"00",X"05",X"22",X"15",
		X"99",X"22",X"1A",X"99",X"C3",X"FE",X"30",X"3D",X"32",X"19",X"98",X"C0",X"AF",X"32",X"1A",X"9C",
		X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"80",X"88",X"80",X"88",X"FF",X"98",X"FF",X"98",X"90",X"FF",X"90",X"FF",X"FF",X"98",X"FF",X"98",
		X"90",X"FF",X"90",X"FF",X"A0",X"A8",X"A0",X"A8",X"FF",X"B8",X"FF",X"B8",X"B0",X"FF",X"B0",X"FF",
		X"FF",X"B8",X"FF",X"B8",X"B0",X"FF",X"B0",X"FF",X"C0",X"C8",X"C0",X"C8",X"FF",X"D8",X"FF",X"D8",
		X"D0",X"FF",X"D0",X"FF",X"FF",X"D8",X"FF",X"D8",X"D0",X"FF",X"D0",X"FF",X"3A",X"18",X"9C",X"A7",
		X"C8",X"3A",X"04",X"99",X"A7",X"C8",X"3A",X"18",X"98",X"A7",X"20",X"44",X"21",X"18",X"9C",X"11",
		X"09",X"9C",X"3A",X"10",X"9C",X"96",X"30",X"02",X"ED",X"44",X"FE",X"08",X"D0",X"47",X"EB",X"3A",
		X"01",X"9C",X"96",X"30",X"02",X"ED",X"44",X"FE",X"08",X"D0",X"CD",X"34",X"34",X"CD",X"D5",X"33",
		X"3E",X"40",X"32",X"18",X"98",X"3A",X"2F",X"99",X"A7",X"28",X"04",X"3E",X"34",X"18",X"02",X"3E",
		X"37",X"32",X"08",X"9C",X"21",X"00",X"05",X"22",X"15",X"99",X"22",X"1A",X"99",X"C3",X"FE",X"30",
		X"3D",X"32",X"18",X"98",X"C0",X"AF",X"32",X"18",X"9C",X"C9",X"3A",X"02",X"99",X"A7",X"C0",X"2F",
		X"32",X"02",X"99",X"D9",X"21",X"00",X"99",X"34",X"CD",X"06",X"19",X"CD",X"F7",X"33",X"D9",X"C9",
		X"3A",X"04",X"99",X"A7",X"C8",X"3A",X"02",X"98",X"E6",X"1F",X"C0",X"CD",X"A5",X"2F",X"E6",X"07",
		X"FE",X"03",X"D0",X"3E",X"FF",X"32",X"70",X"98",X"C9",X"3A",X"04",X"99",X"A7",X"C8",X"3A",X"62",
		X"98",X"21",X"60",X"98",X"86",X"77",X"D0",X"21",X"8A",X"9A",X"11",X"8B",X"9A",X"01",X"0B",X"00",
		X"ED",X"B8",X"21",X"15",X"9B",X"11",X"17",X"9B",X"01",X"16",X"00",X"ED",X"B8",X"2A",X"00",X"9B",
		X"11",X"E0",X"FF",X"19",X"22",X"00",X"9B",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"40",X"80",X"80",X"40",X"FF",X"C0",X"FF",X"80",X"00",X"FF",X"80",X"FF",X"FF",X"40",X"FF",X"00",
		X"40",X"FF",X"C0",X"FF",X"40",X"80",X"80",X"40",X"FF",X"C0",X"FF",X"80",X"00",X"FF",X"80",X"FF",
		X"FF",X"40",X"FF",X"00",X"40",X"FF",X"C0",X"FF",X"40",X"80",X"80",X"40",X"FF",X"C0",X"FF",X"80",
		X"00",X"FF",X"80",X"FF",X"FF",X"40",X"FF",X"00",X"40",X"FF",X"C0",X"FF",X"DD",X"21",X"74",X"98",
		X"DD",X"7E",X"00",X"A7",X"C4",X"4E",X"3F",X"DD",X"23",X"DD",X"7E",X"00",X"A7",X"C8",X"FD",X"21",
		X"86",X"98",X"06",X"06",X"FD",X"7E",X"F0",X"A7",X"28",X"2A",X"FD",X"7E",X"00",X"DD",X"96",X"10",
		X"30",X"02",X"ED",X"44",X"FE",X"04",X"30",X"1C",X"FD",X"7E",X"10",X"DD",X"96",X"20",X"30",X"02",
		X"ED",X"44",X"FE",X"04",X"30",X"0E",X"AF",X"DD",X"77",X"00",X"DD",X"77",X"10",X"FD",X"77",X"F0",
		X"FD",X"77",X"00",X"C9",X"FD",X"23",X"10",X"CC",X"C9",X"3A",X"05",X"99",X"A7",X"C8",X"3A",X"65",
		X"98",X"21",X"63",X"98",X"86",X"77",X"D0",X"21",X"AA",X"9A",X"11",X"AB",X"9A",X"01",X"0B",X"00",
		X"ED",X"B8",X"21",X"55",X"9B",X"11",X"57",X"9B",X"01",X"16",X"00",X"ED",X"B8",X"2A",X"40",X"9B",
		X"11",X"20",X"00",X"19",X"22",X"40",X"9B",X"C9",X"3A",X"03",X"99",X"A7",X"28",X"2A",X"FE",X"08",
		X"D0",X"21",X"A4",X"8B",X"11",X"E0",X"FF",X"47",X"4F",X"36",X"96",X"19",X"10",X"FB",X"21",X"44",
		X"8B",X"36",X"A4",X"21",X"A4",X"83",X"47",X"36",X"38",X"19",X"10",X"FB",X"3E",X"07",X"91",X"D8",
		X"C8",X"47",X"36",X"20",X"19",X"10",X"FB",X"C9",X"21",X"A4",X"83",X"11",X"E0",X"FF",X"06",X"08",
		X"36",X"20",X"19",X"10",X"FB",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
