library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity kick_sp_bits_3 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of kick_sp_bits_3 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"00",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"E0",X"00",X"0E",
		X"00",X"00",X"00",X"0E",X"00",X"00",X"E0",X"0E",X"00",X"00",X"0E",X"0E",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"0E",X"00",X"00",X"E0",X"E0",X"00",X"00",X"E0",
		X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",X"00",X"00",X"EE",X"E0",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",
		X"D0",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",
		X"E0",X"00",X"00",X"E0",X"0E",X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"EE",X"00",X"00",X"0E",X"0E",X"00",X"00",X"E0",X"0E",X"00",X"00",X"00",X"0E",
		X"00",X"E0",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"EE",X"00",X"00",X"0E",X"EE",X"EE",X"00",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",
		X"E0",X"00",X"00",X"E0",X"0E",X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"0D",X"00",X"00",X"EE",
		X"0D",X"00",X"00",X"EE",X"0D",X"00",X"0E",X"0E",X"5D",X"00",X"E0",X"0E",X"DD",X"00",X"00",X"0E",
		X"DD",X"E0",X"00",X"0E",X"DD",X"0E",X"00",X"0E",X"BD",X"11",X"00",X"0E",X"BD",X"EE",X"EE",X"EE",
		X"44",X"44",X"77",X"77",X"44",X"44",X"77",X"77",X"44",X"44",X"77",X"77",X"44",X"44",X"77",X"77",
		X"44",X"44",X"77",X"77",X"44",X"44",X"77",X"77",X"44",X"44",X"77",X"77",X"44",X"44",X"77",X"70",
		X"44",X"44",X"77",X"70",X"00",X"44",X"77",X"00",X"00",X"44",X"00",X"00",X"00",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"77",X"22",X"44",X"33",X"77",X"22",X"44",X"33",X"77",X"33",X"44",X"33",X"77",X"33",
		X"44",X"33",X"77",X"33",X"44",X"33",X"77",X"33",X"44",X"33",X"77",X"30",X"44",X"33",X"77",X"00",
		X"44",X"00",X"70",X"00",X"44",X"00",X"7B",X"00",X"44",X"44",X"BB",X"00",X"44",X"44",X"B0",X"00",
		X"44",X"44",X"BB",X"00",X"44",X"44",X"BB",X"00",X"04",X"44",X"B0",X"00",X"04",X"00",X"BB",X"00",
		X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"77",X"77",X"33",X"33",X"77",X"77",X"44",X"33",X"77",X"77",X"44",X"33",X"77",X"77",
		X"44",X"35",X"77",X"77",X"44",X"5F",X"77",X"00",X"44",X"55",X"77",X"00",X"44",X"55",X"77",X"00",
		X"44",X"5F",X"77",X"00",X"44",X"F5",X"77",X"00",X"44",X"40",X"00",X"00",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BA",X"00",X"00",X"04",X"BA",X"00",X"00",X"04",X"BA",
		X"00",X"00",X"44",X"BB",X"00",X"00",X"44",X"BB",X"00",X"00",X"44",X"BB",X"00",X"00",X"44",X"BB",
		X"00",X"00",X"44",X"BB",X"00",X"00",X"44",X"AB",X"00",X"00",X"44",X"AA",X"00",X"00",X"04",X"A0",
		X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0A",X"00",X"00",X"04",X"0A",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"BB",X"00",X"00",X"44",X"BB",X"00",X"00",X"44",X"BB",X"00",X"00",X"44",X"BA",
		X"00",X"00",X"44",X"AA",X"00",X"00",X"44",X"AA",X"00",X"00",X"44",X"AA",X"00",X"00",X"04",X"AA",
		X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"04",X"BB",X"00",X"00",X"44",X"AA",X"00",X"00",X"44",X"BB",
		X"00",X"00",X"44",X"BB",X"00",X"00",X"44",X"BB",X"00",X"00",X"44",X"AB",X"00",X"00",X"44",X"AA",
		X"00",X"00",X"44",X"A0",X"00",X"00",X"44",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"01",X"11",
		X"00",X"00",X"01",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",
		X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"77",X"11",
		X"00",X"00",X"77",X"11",X"00",X"00",X"77",X"01",X"00",X"33",X"77",X"77",X"00",X"33",X"77",X"77",
		X"40",X"33",X"77",X"77",X"45",X"33",X"77",X"77",X"33",X"33",X"77",X"77",X"33",X"33",X"77",X"77",
		X"00",X"00",X"DD",X"D0",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"D0",
		X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"B0",X"B0",X"00",X"00",
		X"BB",X"00",X"00",X"70",X"0B",X"00",X"00",X"70",X"0B",X"00",X"00",X"77",X"00",X"0B",X"00",X"77",
		X"00",X"B0",X"00",X"77",X"00",X"B0",X"00",X"77",X"0B",X"00",X"00",X"77",X"BB",X"00",X"00",X"77",
		X"B0",X"00",X"00",X"77",X"00",X"F0",X"00",X"77",X"00",X"F0",X"07",X"77",X"00",X"F0",X"07",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"00",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"E0",X"00",X"0E",
		X"00",X"00",X"00",X"0E",X"00",X"00",X"E0",X"0E",X"00",X"00",X"0E",X"0E",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"0E",X"00",X"00",X"E0",X"E0",X"00",X"00",X"E0",
		X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",X"00",X"00",X"EE",X"E0",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BD",X"EE",X"D0",X"0E",X"DD",X"55",X"DD",X"0E",X"DD",X"7E",X"DD",X"0E",X"77",X"E5",X"00",X"0E",
		X"00",X"00",X"E0",X"0E",X"00",X"00",X"0E",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"0E",X"00",X"00",X"E0",X"E0",X"00",X"00",X"E0",
		X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"EE",X"EE",X"EE",X"77",X"88",X"00",X"0E",X"77",X"88",X"00",X"0E",X"00",X"88",X"00",X"0E",
		X"00",X"88",X"00",X"0E",X"00",X"88",X"00",X"0E",X"00",X"0E",X"E0",X"0E",X"00",X"0E",X"E0",X"EE",
		X"0E",X"E0",X"0E",X"EE",X"E0",X"E0",X"0E",X"EE",X"00",X"E0",X"00",X"E0",X"00",X"E0",X"00",X"E0",
		X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",
		X"00",X"00",X"07",X"70",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",
		X"00",X"50",X"77",X"77",X"00",X"55",X"77",X"77",X"00",X"F5",X"77",X"77",X"00",X"45",X"77",X"77",
		X"00",X"40",X"77",X"77",X"05",X"43",X"77",X"07",X"03",X"43",X"77",X"11",X"33",X"44",X"77",X"11",
		X"33",X"44",X"77",X"11",X"33",X"44",X"77",X"11",X"33",X"44",X"77",X"22",X"33",X"44",X"77",X"22",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",
		X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"11",X"00",X"04",X"00",X"11",X"00",X"04",X"77",X"11",X"00",X"B4",X"77",X"11",
		X"00",X"BB",X"77",X"11",X"05",X"BB",X"77",X"11",X"03",X"BB",X"77",X"11",X"33",X"BB",X"77",X"11",
		X"33",X"F5",X"77",X"77",X"33",X"F5",X"77",X"77",X"33",X"F5",X"77",X"77",X"33",X"44",X"77",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"B0",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"0B",X"00",X"01",X"10",X"00",X"00",X"01",X"11",
		X"0B",X"00",X"11",X"11",X"BB",X"00",X"11",X"11",X"B0",X"00",X"11",X"11",X"00",X"00",X"11",X"11",
		X"00",X"40",X"11",X"11",X"00",X"44",X"11",X"11",X"00",X"44",X"77",X"11",X"00",X"44",X"77",X"11",
		X"00",X"54",X"77",X"01",X"05",X"33",X"77",X"77",X"03",X"33",X"77",X"77",X"33",X"33",X"77",X"77",
		X"33",X"33",X"77",X"77",X"33",X"33",X"77",X"77",X"33",X"33",X"77",X"77",X"33",X"33",X"77",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"5F",X"00",X"00",X"00",X"5F",X"00",X"00",X"00",X"5F",X"00",X"00",X"00",X"44",X"00",X"07",
		X"00",X"44",X"00",X"77",X"00",X"44",X"00",X"77",X"00",X"44",X"00",X"77",X"00",X"44",X"00",X"77",
		X"00",X"44",X"00",X"77",X"00",X"44",X"00",X"77",X"00",X"54",X"77",X"77",X"00",X"33",X"77",X"77",
		X"00",X"33",X"77",X"77",X"05",X"33",X"77",X"77",X"03",X"33",X"77",X"77",X"33",X"33",X"77",X"77",
		X"33",X"33",X"77",X"77",X"33",X"33",X"77",X"77",X"33",X"33",X"77",X"72",X"33",X"33",X"77",X"22",
		X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",
		X"00",X"00",X"DD",X"DD",X"00",X"0D",X"DD",X"D0",X"00",X"0D",X"DD",X"00",X"00",X"0D",X"DD",X"00",
		X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"07",X"00",X"00",X"BB",X"07",
		X"00",X"00",X"B0",X"77",X"00",X"00",X"00",X"77",X"00",X"04",X"00",X"77",X"00",X"44",X"00",X"77",
		X"00",X"44",X"00",X"77",X"00",X"44",X"00",X"77",X"44",X"44",X"00",X"77",X"44",X"44",X"00",X"77",
		X"44",X"40",X"00",X"77",X"44",X"00",X"07",X"77",X"44",X"00",X"77",X"77",X"44",X"00",X"77",X"77",
		X"44",X"00",X"77",X"70",X"33",X"33",X"77",X"70",X"33",X"33",X"77",X"20",X"35",X"53",X"77",X"2E",
		X"35",X"53",X"77",X"EE",X"33",X"33",X"77",X"11",X"33",X"33",X"77",X"11",X"44",X"03",X"77",X"11",
		X"44",X"00",X"77",X"11",X"44",X"00",X"77",X"11",X"44",X"00",X"77",X"11",X"44",X"40",X"00",X"11",
		X"44",X"44",X"00",X"11",X"44",X"44",X"00",X"11",X"00",X"44",X"00",X"11",X"00",X"44",X"00",X"11",
		X"00",X"44",X"00",X"01",X"00",X"44",X"00",X"00",X"B0",X"44",X"00",X"00",X"BB",X"44",X"00",X"11",
		X"BB",X"44",X"00",X"11",X"BB",X"44",X"00",X"11",X"BB",X"40",X"00",X"11",X"BB",X"00",X"00",X"11",
		X"0B",X"00",X"01",X"11",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"DD",
		X"00",X"00",X"F5",X"DD",X"00",X"00",X"5F",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",
		X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"0D",X"DD",X"00",X"00",X"00",X"DD",
		X"77",X"75",X"D2",X"0E",X"77",X"7F",X"D2",X"0E",X"77",X"05",X"DD",X"0E",X"77",X"0E",X"DD",X"0E",
		X"00",X"E0",X"DD",X"EE",X"EE",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"E0",X"E0",X"00",X"00",X"E0",X"E0",
		X"E0",X"00",X"0E",X"00",X"E0",X"00",X"0E",X"00",X"EE",X"00",X"0E",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3E",X"DD",X"00",X"0E",X"E3",X"DD",X"00",X"0E",X"33",X"DD",X"00",X"0E",X"33",X"D2",X"00",X"0E",
		X"30",X"D2",X"EE",X"0E",X"00",X"D2",X"00",X"0E",X"00",X"02",X"00",X"0E",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"0E",X"00",X"00",X"E0",X"E0",X"00",X"00",X"E0",
		X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"EE",X"88",X"00",X"00",X"E0",X"88",X"00",X"00",X"E0",X"88",X"00",X"00",
		X"E0",X"88",X"00",X"E0",X"7E",X"88",X"20",X"E0",X"77",X"00",X"20",X"EE",X"77",X"00",X"20",X"EE",
		X"77",X"00",X"20",X"EE",X"77",X"00",X"80",X"0E",X"77",X"00",X"80",X"0E",X"77",X"00",X"EE",X"0E",
		X"77",X"30",X"00",X"0E",X"77",X"33",X"00",X"0E",X"77",X"33",X"00",X"0E",X"77",X"5D",X"00",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"DD",X"00",X"00",
		X"00",X"DD",X"00",X"E0",X"00",X"DD",X"00",X"E0",X"E0",X"DD",X"0E",X"EE",X"7E",X"DD",X"0E",X"EE",
		X"77",X"0E",X"E0",X"EE",X"77",X"0E",X"E0",X"0E",X"77",X"0E",X"00",X"0E",X"77",X"0E",X"00",X"0E",
		X"77",X"0E",X"00",X"0E",X"77",X"75",X"00",X"0E",X"77",X"77",X"00",X"0E",X"77",X"77",X"00",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"EE",X"00",X"0E",X"00",X"E0",X"00",X"0E",X"00",X"E0",X"00",X"0E",X"00",
		X"00",X"00",X"E0",X"E0",X"00",X"00",X"E0",X"E0",X"00",X"00",X"D0",X"EE",X"00",X"00",X"DD",X"EE",
		X"00",X"00",X"DD",X"EE",X"00",X"00",X"DD",X"0E",X"EE",X"00",X"DD",X"0E",X"00",X"E0",X"DD",X"EE",
		X"77",X"0E",X"DD",X"0E",X"77",X"05",X"DD",X"0E",X"77",X"7F",X"D2",X"0E",X"77",X"75",X"D2",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"55",
		X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",
		X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",
		X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",
		X"00",X"00",X"00",X"44",X"00",X"00",X"05",X"44",X"00",X"00",X"B5",X"44",X"00",X"00",X"BF",X"04",
		X"00",X"00",X"B5",X"04",X"00",X"0B",X"05",X"00",X"00",X"0B",X"00",X"00",X"00",X"B0",X"00",X"00",
		X"00",X"00",X"44",X"BB",X"00",X"00",X"44",X"BA",X"00",X"00",X"44",X"AB",X"00",X"00",X"44",X"BB",
		X"00",X"00",X"04",X"B0",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"B0",
		X"00",X"00",X"44",X"BB",X"00",X"00",X"44",X"AB",X"00",X"00",X"44",X"BA",X"00",X"00",X"44",X"BB",
		X"33",X"55",X"77",X"77",X"33",X"53",X"77",X"77",X"33",X"33",X"77",X"77",X"33",X"33",X"77",X"77",
		X"44",X"33",X"77",X"77",X"44",X"03",X"77",X"00",X"44",X"00",X"77",X"00",X"44",X"00",X"77",X"00",
		X"44",X"00",X"77",X"00",X"44",X"00",X"77",X"00",X"44",X"00",X"00",X"00",X"04",X"00",X"00",X"00",
		X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"5F",X"00",X"00",X"00",
		X"BF",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",
		X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",
		X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",
		X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",
		X"5F",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"02",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",
		X"04",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"70",X"00",
		X"44",X"00",X"77",X"00",X"44",X"00",X"77",X"00",X"44",X"03",X"77",X"00",X"44",X"33",X"77",X"77",
		X"33",X"33",X"77",X"77",X"33",X"33",X"77",X"77",X"33",X"53",X"77",X"77",X"33",X"55",X"77",X"77",
		X"33",X"44",X"77",X"22",X"44",X"44",X"77",X"22",X"44",X"43",X"77",X"11",X"44",X"33",X"77",X"11",
		X"44",X"33",X"77",X"11",X"44",X"33",X"77",X"10",X"44",X"33",X"77",X"00",X"44",X"33",X"77",X"00",
		X"44",X"44",X"77",X"00",X"00",X"44",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"04",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"04",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"77",X"00",X"00",X"3F",X"77",X"00",X"00",X"3F",X"77",X"00",X"00",X"3F",X"77",
		X"00",X"00",X"3F",X"77",X"00",X"00",X"33",X"77",X"00",X"00",X"33",X"77",X"00",X"00",X"33",X"77",
		X"00",X"00",X"33",X"00",X"00",X"03",X"33",X"00",X"00",X"33",X"33",X"00",X"00",X"33",X"33",X"00",
		X"00",X"33",X"33",X"00",X"00",X"33",X"33",X"00",X"00",X"33",X"33",X"00",X"00",X"33",X"33",X"00",
		X"00",X"35",X"30",X"00",X"00",X"33",X"00",X"00",X"04",X"33",X"00",X"00",X"04",X"B3",X"00",X"00",
		X"AA",X"B3",X"00",X"00",X"AA",X"B3",X"44",X"44",X"BB",X"B3",X"44",X"44",X"6B",X"B3",X"44",X"44",
		X"B6",X"B3",X"44",X"44",X"6B",X"B3",X"44",X"00",X"BB",X"A4",X"44",X"00",X"4A",X"A0",X"00",X"00",
		X"44",X"A0",X"00",X"00",X"44",X"A0",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"0D",X"D0",X"E0",X"77",X"00",X"D0",X"00",X"77",X"00",X"D0",X"00",X"77",X"00",X"D0",X"00",
		X"77",X"00",X"D0",X"00",X"77",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",X"00",X"00",X"00",
		X"00",X"0E",X"0E",X"00",X"00",X"E0",X"EE",X"00",X"00",X"E0",X"EE",X"00",X"EE",X"00",X"E0",X"00",
		X"EE",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0B",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"B0",X"00",X"00",X"BB",X"00",X"00",X"00",
		X"BB",X"BB",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",
		X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",
		X"0E",X"00",X"00",X"EE",X"0E",X"00",X"00",X"EE",X"EE",X"00",X"00",X"EE",X"EE",X"00",X"00",X"0E",
		X"E0",X"00",X"00",X"0E",X"E0",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",
		X"00",X"00",X"0E",X"0E",X"00",X"0D",X"E0",X"0E",X"00",X"DD",X"E0",X"0E",X"00",X"DD",X"00",X"0E",
		X"00",X"DD",X"00",X"0E",X"07",X"DD",X"00",X"EE",X"77",X"DD",X"00",X"EE",X"77",X"DD",X"DE",X"EE",
		X"33",X"34",X"00",X"BE",X"33",X"44",X"00",X"EE",X"33",X"44",X"44",X"BB",X"33",X"44",X"44",X"EE",
		X"33",X"44",X"44",X"BB",X"33",X"44",X"44",X"EB",X"33",X"44",X"00",X"EE",X"33",X"43",X"00",X"EE",
		X"33",X"33",X"00",X"EE",X"03",X"55",X"E0",X"EE",X"03",X"5F",X"0E",X"E0",X"AA",X"F5",X"00",X"E0",
		X"AA",X"B5",X"00",X"00",X"BB",X"B0",X"00",X"00",X"BA",X"B4",X"00",X"00",X"AB",X"A4",X"00",X"00",
		X"AB",X"B4",X"00",X"00",X"BB",X"44",X"EE",X"00",X"BB",X"44",X"44",X"00",X"BB",X"44",X"44",X"0B",
		X"BB",X"04",X"45",X"BB",X"BB",X"00",X"45",X"00",X"BB",X"00",X"45",X"00",X"00",X"00",X"45",X"00",
		X"00",X"40",X"05",X"BB",X"00",X"40",X"00",X"0B",X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"B0",
		X"00",X"40",X"00",X"BB",X"00",X"40",X"00",X"0B",X"00",X"40",X"00",X"00",X"00",X"04",X"00",X"00",
		X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",
		X"DB",X"DD",X"00",X"00",X"DB",X"0D",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"70",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"70",X"00",
		X"00",X"EE",X"77",X"00",X"00",X"EE",X"77",X"00",X"00",X"00",X"E7",X"00",X"00",X"00",X"E7",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"77",X"EE",X"00",X"0E",X"77",X"7E",X"00",X"0E",X"77",X"7E",X"00",
		X"0E",X"77",X"77",X"00",X"77",X"77",X"77",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",
		X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"33",X"77",X"00",X"00",
		X"33",X"7E",X"00",X"00",X"33",X"70",X"EE",X"B0",X"33",X"30",X"00",X"00",X"33",X"3E",X"00",X"0B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"04",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"04",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"4F",X"40",X"00",X"00",X"FF",X"44",X"00",
		X"00",X"44",X"44",X"00",X"04",X"44",X"45",X"00",X"04",X"44",X"45",X"00",X"04",X"44",X"45",X"00",
		X"04",X"44",X"55",X"00",X"04",X"44",X"55",X"00",X"04",X"44",X"55",X"00",X"04",X"44",X"55",X"E0",
		X"00",X"44",X"55",X"E0",X"00",X"44",X"54",X"E0",X"00",X"45",X"50",X"0E",X"00",X"55",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"60",X"00",X"00",X"F6",X"66",X"00",
		X"00",X"FF",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"00",
		X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"66",X"6D",X"00",X"00",X"66",X"DD",X"E0",
		X"00",X"66",X"DD",X"E0",X"00",X"66",X"D6",X"E0",X"00",X"DD",X"60",X"0E",X"00",X"DD",X"00",X"00",
		X"00",X"DD",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"00",
		X"00",X"CC",X"AA",X"00",X"0C",X"FF",X"AA",X"00",X"0C",X"FF",X"AA",X"00",X"CC",X"FF",X"AA",X"00",
		X"CA",X"CC",X"AA",X"00",X"CA",X"CC",X"AA",X"00",X"CA",X"CC",X"AA",X"00",X"CA",X"CC",X"AA",X"00",
		X"CA",X"FF",X"AA",X"00",X"CA",X"FF",X"AA",X"00",X"CA",X"FF",X"AA",X"00",X"CA",X"CC",X"AA",X"00",
		X"CC",X"CC",X"AA",X"00",X"0C",X"CC",X"AA",X"00",X"0C",X"CC",X"AA",X"00",X"00",X"AA",X"AA",X"00",
		X"00",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"00",
		X"00",X"CC",X"66",X"00",X"0C",X"FF",X"66",X"00",X"0C",X"FF",X"66",X"00",X"CC",X"FF",X"66",X"00",
		X"C6",X"CC",X"66",X"00",X"C6",X"CC",X"66",X"00",X"C6",X"CC",X"66",X"00",X"C6",X"CC",X"66",X"00",
		X"C6",X"FF",X"66",X"00",X"C6",X"FF",X"66",X"00",X"C6",X"FF",X"66",X"00",X"C6",X"CC",X"66",X"00",
		X"CC",X"CC",X"66",X"00",X"0C",X"CC",X"66",X"00",X"0C",X"CC",X"66",X"00",X"00",X"66",X"66",X"00",
		X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",
		X"00",X"CC",X"BB",X"00",X"0C",X"FF",X"BB",X"00",X"0C",X"FF",X"BB",X"00",X"CC",X"FF",X"BB",X"00",
		X"CB",X"CC",X"BB",X"00",X"CB",X"CC",X"BB",X"00",X"CB",X"CC",X"BB",X"00",X"CB",X"CC",X"BB",X"00",
		X"CB",X"FF",X"BB",X"00",X"CB",X"FF",X"BB",X"00",X"CB",X"FF",X"BB",X"00",X"CB",X"CC",X"BB",X"00",
		X"CC",X"CC",X"BB",X"00",X"0C",X"CC",X"BB",X"00",X"0C",X"CC",X"BB",X"00",X"00",X"BB",X"BB",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",
		X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AF",X"A0",X"00",X"00",X"FF",X"AA",X"00",
		X"00",X"FF",X"AA",X"00",X"0A",X"AA",X"AA",X"00",X"0A",X"AA",X"AA",X"00",X"0A",X"AA",X"AA",X"00",
		X"0A",X"AA",X"A9",X"00",X"0A",X"AA",X"99",X"00",X"0A",X"AA",X"99",X"00",X"0A",X"AA",X"99",X"E0",
		X"00",X"AA",X"99",X"E0",X"00",X"A9",X"9A",X"E0",X"00",X"99",X"A0",X"0E",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"A9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"70",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"50",X"00",
		X"00",X"40",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"0F",X"05",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"04",X"00",
		X"00",X"00",X"40",X"00",X"00",X"0A",X"00",X"00",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"A0",X"00",X"00",X"AA",X"05",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"05",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",
		X"00",X"A0",X"00",X"00",X"00",X"0A",X"A0",X"00",X"00",X"0A",X"AA",X"00",X"00",X"50",X"A0",X"00",
		X"00",X"45",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",
		X"04",X"44",X"04",X"00",X"00",X"54",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"A0",X"40",X"05",X"00",X"0A",X"00",
		X"45",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"04",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"04",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"04",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"04",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"44",X"00",X"00",X"40",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"09",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"A9",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"A9",X"00",X"BB",X"99",X"99",X"00",
		X"00",X"99",X"A9",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"A9",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"99",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"40",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",
		X"00",X"60",X"AA",X"00",X"00",X"60",X"AA",X"00",X"00",X"60",X"66",X"00",X"00",X"60",X"00",X"00",
		X"00",X"60",X"00",X"00",X"00",X"66",X"06",X"00",X"00",X"AA",X"06",X"00",X"00",X"AA",X"06",X"00",
		X"00",X"66",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"60",X"A6",X"00",
		X"00",X"60",X"AA",X"00",X"00",X"60",X"AA",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",
		X"00",X"60",X"AA",X"00",X"00",X"60",X"AA",X"00",X"00",X"60",X"66",X"00",X"00",X"60",X"00",X"00",
		X"00",X"60",X"00",X"00",X"00",X"66",X"06",X"00",X"00",X"AA",X"06",X"00",X"00",X"AA",X"06",X"00",
		X"00",X"66",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"AA",X"AA",X"00",
		X"00",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"00",X"00",X"66",X"66",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"AA",X"AA",X"00",
		X"00",X"AA",X"AA",X"00",X"00",X"AA",X"66",X"00",X"00",X"AA",X"00",X"00",X"00",X"6A",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"60",X"AA",X"00",
		X"00",X"60",X"AA",X"00",X"00",X"60",X"66",X"00",X"00",X"60",X"00",X"00",X"00",X"60",X"00",X"00",
		X"00",X"66",X"06",X"00",X"00",X"AA",X"06",X"00",X"00",X"AA",X"06",X"00",X"00",X"66",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"AA",X"AA",X"00",
		X"00",X"AA",X"AA",X"00",X"00",X"AA",X"66",X"00",X"00",X"AA",X"00",X"00",X"00",X"6A",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"66",X"60",X"00",X"00",X"60",X"66",X"00",
		X"00",X"60",X"A6",X"00",X"00",X"66",X"AA",X"00",X"00",X"A6",X"AA",X"00",X"00",X"A6",X"6A",X"00",
		X"00",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"00",X"00",X"06",X"6A",X"00",
		X"00",X"06",X"AA",X"00",X"00",X"06",X"A6",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"66",X"00",X"00",X"06",X"A6",X"00",X"00",X"06",X"AA",X"00",X"00",X"06",X"6A",X"00",
		X"00",X"06",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",
		X"00",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"00",X"00",X"66",X"66",X"00",X"00",X"60",X"00",X"00",
		X"00",X"60",X"00",X"00",X"00",X"66",X"06",X"00",X"00",X"A6",X"06",X"00",X"00",X"A6",X"06",X"00",
		X"00",X"66",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"00",X"00",X"06",X"6A",X"00",
		X"00",X"06",X"AA",X"00",X"00",X"06",X"A6",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"66",X"00",X"00",X"06",X"A6",X"00",X"00",X"06",X"AA",X"00",X"00",X"06",X"6A",X"00",
		X"00",X"06",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"00",
		X"00",X"00",X"66",X"00",X"00",X"A0",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"6A",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"00",X"00",X"06",X"6A",X"00",
		X"00",X"06",X"AA",X"00",X"00",X"06",X"A6",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"66",X"00",X"00",X"06",X"A6",X"00",X"00",X"06",X"AA",X"00",X"00",X"06",X"6A",X"00",
		X"00",X"06",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",
		X"00",X"60",X"AA",X"00",X"00",X"60",X"AA",X"00",X"00",X"60",X"66",X"00",X"00",X"60",X"00",X"00",
		X"00",X"60",X"00",X"00",X"00",X"66",X"06",X"00",X"00",X"AA",X"06",X"00",X"00",X"AA",X"06",X"00",
		X"00",X"66",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"00",X"00",X"06",X"6A",X"00",
		X"00",X"06",X"AA",X"00",X"00",X"06",X"A6",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"66",X"00",X"00",X"06",X"A6",X"00",X"00",X"06",X"AA",X"00",X"00",X"06",X"6A",X"00",
		X"00",X"06",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"55",X"55",X"00",X"00",X"55",X"55",X"00",
		X"00",X"CC",X"55",X"00",X"0C",X"FF",X"55",X"00",X"0C",X"FF",X"55",X"00",X"CC",X"FF",X"55",X"00",
		X"C5",X"CC",X"55",X"00",X"C5",X"CC",X"55",X"00",X"C5",X"CC",X"55",X"00",X"C5",X"CC",X"55",X"00",
		X"C5",X"FF",X"55",X"00",X"C5",X"FF",X"55",X"00",X"C5",X"FF",X"55",X"00",X"C5",X"CC",X"55",X"00",
		X"CC",X"CC",X"55",X"00",X"0C",X"CC",X"55",X"00",X"0C",X"CC",X"55",X"00",X"00",X"55",X"55",X"00",
		X"00",X"55",X"55",X"00",X"00",X"55",X"55",X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
