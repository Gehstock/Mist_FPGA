library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity GALAXIAN_1H is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of GALAXIAN_1H is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",X"00",X"02",X"02",X"FE",X"FE",X"42",X"02",X"00",X"00",
		X"62",X"F2",X"BA",X"9A",X"9E",X"CE",X"46",X"00",X"8C",X"DE",X"F2",X"B2",X"92",X"86",X"04",X"00",
		X"08",X"FE",X"FE",X"C8",X"68",X"38",X"18",X"00",X"1C",X"BE",X"A2",X"A2",X"A2",X"E6",X"E4",X"00",
		X"0C",X"9E",X"92",X"92",X"D2",X"7E",X"3C",X"00",X"C0",X"E0",X"B0",X"9E",X"8E",X"C0",X"C0",X"00",
		X"0C",X"6E",X"9A",X"9A",X"B2",X"F2",X"6C",X"00",X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",X"00",
		X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",
		X"44",X"C6",X"82",X"82",X"C6",X"7C",X"38",X"00",X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",
		X"82",X"92",X"92",X"92",X"FE",X"FE",X"00",X"00",X"80",X"90",X"90",X"90",X"90",X"FE",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",
		X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",X"44",X"C6",X"82",X"82",X"C6",X"7C",X"38",X"00",
		X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",X"82",X"92",X"92",X"92",X"FE",X"FE",X"00",X"00",
		X"80",X"90",X"90",X"90",X"90",X"FE",X"FE",X"00",X"9E",X"9E",X"92",X"82",X"C6",X"7C",X"38",X"00",
		X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",X"82",X"82",X"FE",X"FE",X"82",X"82",X"00",X"00",
		X"FC",X"FE",X"02",X"02",X"02",X"06",X"04",X"00",X"82",X"C6",X"6E",X"3C",X"18",X"FE",X"FE",X"00",
		X"02",X"02",X"02",X"02",X"FE",X"FE",X"00",X"00",X"FE",X"FE",X"70",X"38",X"70",X"FE",X"FE",X"00",
		X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",X"00",
		X"70",X"F8",X"88",X"88",X"88",X"FE",X"FE",X"00",X"7A",X"FC",X"8E",X"8A",X"82",X"FE",X"7C",X"00",
		X"72",X"F6",X"9E",X"8C",X"88",X"FE",X"FE",X"00",X"0C",X"5E",X"D2",X"92",X"92",X"F6",X"64",X"00",
		X"80",X"80",X"FE",X"FE",X"80",X"80",X"00",X"00",X"FC",X"FE",X"02",X"02",X"02",X"FE",X"FC",X"00",
		X"F0",X"F8",X"1C",X"0E",X"1C",X"F8",X"F0",X"00",X"F8",X"FE",X"1C",X"38",X"1C",X"FE",X"F8",X"00",
		X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",X"C0",X"F0",X"1E",X"1E",X"F0",X"C0",X"00",X"00",
		X"C2",X"E2",X"F2",X"BA",X"9E",X"8E",X"86",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"C0",X"20",X"20",X"70",X"FC",X"7E",X"FC",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"70",X"20",X"20",X"C0",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",X"00",X"00",X"00",X"60",X"20",X"20",X"3C",X"FE",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",X"3F",X"FE",X"3C",X"20",X"20",X"60",X"00",X"00",
		X"00",X"00",X"00",X"06",X"02",X"02",X"03",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",
		X"03",X"0F",X"03",X"02",X"02",X"06",X"00",X"00",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"02",X"02",X"07",X"0F",X"07",X"0F",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"C0",
		X"07",X"02",X"02",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"10",X"10",X"38",X"FE",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"38",X"10",X"10",X"30",X"00",X"00",X"00",
		X"00",X"00",X"03",X"01",X"01",X"03",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"F0",
		X"0F",X"03",X"01",X"01",X"03",X"00",X"00",X"00",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"01",X"01",X"0F",X"07",X"1F",X"00",X"00",X"80",X"00",X"00",X"80",X"C0",X"E0",
		X"07",X"07",X"02",X"04",X"0C",X"00",X"00",X"00",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"0A",X"07",X"1F",X"0F",X"00",X"00",X"80",X"80",X"80",X"80",X"C0",X"C0",
		X"07",X"0F",X"08",X"10",X"00",X"00",X"00",X"00",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"07",X"1B",X"0F",X"0F",X"00",X"00",X"40",X"60",X"C0",X"80",X"C0",X"C0",
		X"0F",X"3B",X"10",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"05",X"07",X"27",X"3F",X"00",X"00",X"00",X"00",X"08",X"D8",X"E0",X"C0",
		X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"05",X"02",X"07",X"2F",X"3B",X"00",X"00",X"00",X"88",X"C8",X"F0",X"C0",X"C0",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"13",X"1F",X"00",X"00",X"00",X"00",X"40",X"40",X"E4",X"FC",
		X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"E0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"38",X"70",X"F7",X"FF",X"00",X"00",X"FC",X"20",X"70",X"E0",X"FC",X"F0",
		X"F7",X"70",X"38",X"00",X"00",X"00",X"00",X"00",X"FC",X"E0",X"70",X"20",X"FC",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"0C",X"7F",X"00",X"00",X"00",X"18",X"08",X"1C",X"FE",X"F8",
		X"0C",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"1C",X"08",X"18",X"00",X"00",X"00",X"00",
		X"02",X"07",X"07",X"0F",X"0F",X"0F",X"1F",X"18",X"00",X"00",X"00",X"80",X"80",X"80",X"C0",X"C0",
		X"17",X"37",X"38",X"3F",X"70",X"7F",X"7F",X"00",X"40",X"60",X"E0",X"E0",X"70",X"F0",X"F0",X"00",
		X"02",X"02",X"07",X"07",X"0F",X"0F",X"1F",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"00",
		X"C3",X"FF",X"FF",X"7E",X"00",X"00",X"C3",X"C3",X"00",X"00",X"7E",X"FF",X"FF",X"C3",X"C3",X"C3",
		X"00",X"01",X"03",X"07",X"03",X"07",X"0F",X"3F",X"80",X"80",X"D8",X"F8",X"F8",X"F0",X"F0",X"F0",
		X"1F",X"1F",X"1F",X"0F",X"03",X"07",X"07",X"01",X"F8",X"F8",X"F0",X"E0",X"F8",X"FC",X"78",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"90",
		X"07",X"02",X"02",X"08",X"00",X"00",X"00",X"00",X"C0",X"80",X"A0",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"24",X"04",X"4E",X"27",X"00",X"00",X"20",X"40",X"11",X"80",X"A4",X"C8",
		X"07",X"03",X"25",X"00",X"08",X"00",X"00",X"00",X"C0",X"20",X"90",X"A0",X"20",X"50",X"00",X"00",
		X"00",X"00",X"42",X"20",X"04",X"0F",X"E7",X"3F",X"00",X"20",X"44",X"C8",X"80",X"80",X"D0",X"EC",
		X"07",X"07",X"0D",X"1D",X"29",X"42",X"01",X"00",X"C0",X"A0",X"B0",X"88",X"44",X"20",X"10",X"08",
		X"07",X"08",X"08",X"08",X"07",X"00",X"09",X"0A",X"C0",X"20",X"20",X"20",X"C0",X"00",X"C0",X"20",
		X"0A",X"0A",X"0E",X"00",X"00",X"0F",X"04",X"00",X"20",X"20",X"40",X"00",X"20",X"E0",X"20",X"00",
		X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"C0",X"20",X"20",X"C0",X"00",X"C0",X"20",X"20",
		X"07",X"00",X"06",X"09",X"08",X"08",X"04",X"00",X"C0",X"00",X"20",X"20",X"A0",X"60",X"20",X"00",
		X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"C0",X"20",X"20",X"C0",X"00",X"C0",X"20",X"20",
		X"07",X"00",X"08",X"0D",X"0B",X"09",X"08",X"00",X"C0",X"00",X"C0",X"20",X"20",X"20",X"20",X"00",
		X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"C0",X"20",X"20",X"C0",X"00",X"C0",X"20",X"20",
		X"07",X"00",X"06",X"09",X"09",X"09",X"06",X"00",X"C0",X"00",X"C0",X"20",X"20",X"20",X"C0",X"00",
		X"1C",X"3E",X"61",X"41",X"43",X"3E",X"1C",X"00",X"01",X"01",X"7F",X"7F",X"21",X"01",X"00",X"00",
		X"31",X"79",X"5D",X"4D",X"4F",X"67",X"23",X"00",X"46",X"6F",X"79",X"59",X"49",X"43",X"02",X"00",
		X"04",X"7F",X"7F",X"64",X"34",X"1C",X"0C",X"00",X"0E",X"5F",X"51",X"51",X"51",X"73",X"72",X"00",
		X"06",X"4F",X"49",X"49",X"69",X"3F",X"1E",X"00",X"60",X"70",X"58",X"4F",X"47",X"60",X"60",X"00",
		X"06",X"37",X"4D",X"4D",X"59",X"79",X"36",X"00",X"3C",X"7E",X"4B",X"49",X"49",X"79",X"30",X"00",
		X"C0",X"C0",X"C0",X"FF",X"FF",X"FF",X"00",X"00",X"DF",X"1F",X"00",X"00",X"7F",X"FF",X"FF",X"C0",
		X"7F",X"FF",X"FF",X"DB",X"DB",X"DB",X"DB",X"DF",X"FF",X"C0",X"C0",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"7F",X"FF",X"FF",X"C0",X"C0",X"FF",X"FF",X"C3",X"C3",X"C3",X"C3",X"FF",X"FF",X"7E",X"00",
		X"20",X"20",X"00",X"10",X"28",X"28",X"28",X"3E",X"2A",X"2A",X"2A",X"12",X"00",X"20",X"20",X"3E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"03",X"01",X"01",X"03",X"00",X"00",X"00",X"80",X"C0",X"E0",X"F0",X"80",X"FC",
		X"03",X"01",X"01",X"03",X"0F",X"00",X"00",X"00",X"80",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"00",
		X"00",X"00",X"06",X"03",X"01",X"01",X"01",X"03",X"00",X"00",X"00",X"C0",X"C0",X"E0",X"F0",X"C0",
		X"00",X"03",X"03",X"07",X"1F",X"07",X"00",X"00",X"F0",X"9C",X"C0",X"E0",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"80",X"E0",X"70",X"F0",X"F0",X"F8",
		X"02",X"03",X"27",X"1F",X"0F",X"02",X"00",X"00",X"48",X"E0",X"98",X"CC",X"E0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"00",X"00",X"60",X"30",X"38",X"78",X"F8",X"F8",
		X"03",X"27",X"3F",X"1F",X"0F",X"00",X"00",X"00",X"78",X"C8",X"A0",X"90",X"C8",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"23",X"00",X"00",X"20",X"10",X"18",X"38",X"FC",X"78",
		X"33",X"1F",X"1F",X"0F",X"01",X"00",X"00",X"00",X"78",X"D8",X"48",X"20",X"B0",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"31",X"1F",X"00",X"00",X"00",X"08",X"08",X"1C",X"7C",X"7C",
		X"1F",X"1F",X"06",X"02",X"00",X"00",X"00",X"00",X"F8",X"B8",X"90",X"C0",X"40",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"10",X"19",X"1F",X"00",X"00",X"00",X"00",X"04",X"04",X"4C",X"7C",
		X"1F",X"0E",X"06",X"02",X"00",X"00",X"00",X"00",X"FC",X"B8",X"B0",X"A0",X"80",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"04",X"00",X"03",X"04",X"08",X"10",X"21",X"20",X"80",
		X"08",X"10",X"10",X"20",X"1C",X"08",X"04",X"08",X"C0",X"A1",X"07",X"01",X"38",X"70",X"F7",X"FF",
		X"00",X"00",X"C3",X"2C",X"10",X"11",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"20",X"10",X"10",
		X"00",X"FE",X"FF",X"FE",X"70",X"E0",X"FC",X"F0",X"08",X"08",X"14",X"14",X"28",X"48",X"10",X"20",
		X"08",X"10",X"10",X"09",X"04",X"03",X"00",X"00",X"F7",X"70",X"38",X"81",X"67",X"11",X"D0",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"03",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"E0",X"70",X"FE",X"FF",X"FE",X"00",X"00",X"40",X"40",X"00",X"00",X"00",X"40",X"40",X"80",
		X"00",X"21",X"19",X"C2",X"24",X"18",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"0D",X"02",X"04",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"02",X"62",X"27",X"10",X"E6",X"92",X"0C",X"68",X"20",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"61",X"13",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"12",X"04",X"F1",X"52",X"31",X"36",X"05",X"04",X"C0",X"20",X"A0",X"20",X"20",X"40",X"40",X"80",
		X"05",X"04",X"02",X"01",X"00",X"01",X"01",X"01",X"C0",X"40",X"40",X"40",X"C0",X"C0",X"FC",X"8A",
		X"01",X"06",X"08",X"00",X"00",X"00",X"00",X"00",X"72",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"02",X"00",X"78",X"20",X"20",X"10",X"10",X"20",X"20",
		X"13",X"0F",X"E3",X"00",X"00",X"00",X"00",X"00",X"70",X"D0",X"10",X"0C",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"00",X"00",X"00",X"10",X"7C",X"FF",X"FF",X"DF",
		X"03",X"07",X"07",X"09",X"0F",X"0F",X"05",X"0D",X"37",X"8F",X"C7",X"82",X"01",X"87",X"E1",X"F9",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"9F",X"FF",X"00",X"00",X"00",X"00",X"00",X"40",X"B8",X"78",
		X"9C",X"2F",X"74",X"F8",X"F1",X"A7",X"0F",X"CF",X"70",X"60",X"F0",X"E0",X"E0",X"C0",X"C0",X"E0",
		X"0E",X"07",X"07",X"0B",X"07",X"03",X"01",X"01",X"FF",X"7F",X"EF",X"F6",X"74",X"8F",X"8B",X"8E",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DF",X"77",X"23",X"03",X"03",X"03",X"00",X"00",
		X"EF",X"EF",X"7F",X"2F",X"8F",X"9F",X"3F",X"7E",X"E0",X"D0",X"F0",X"F0",X"E0",X"E0",X"80",X"10",
		X"6E",X"3E",X"DC",X"F8",X"F8",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"94",X"F7",X"33",
		X"00",X"01",X"00",X"00",X"00",X"03",X"02",X"00",X"1A",X"8E",X"C8",X"FA",X"D6",X"33",X"7D",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"02",X"14",X"35",X"00",X"00",X"00",X"00",X"00",X"40",X"80",X"00",
		X"24",X"28",X"49",X"DF",X"D7",X"77",X"CE",X"F8",X"00",X"00",X"00",X"00",X"80",X"80",X"20",X"00",
		X"01",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"87",X"FB",X"8E",X"19",X"F7",X"63",X"42",X"9C",
		X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"82",X"01",X"01",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"F8",X"EA",X"AE",X"79",X"DC",X"4A",X"C0",X"80",X"40",X"00",X"00",X"00",X"80",X"00",
		X"40",X"70",X"58",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
