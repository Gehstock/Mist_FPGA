library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity gravitar_vec_rom2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of gravitar_vec_rom2 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"FF",X"00",X"01",X"9F",X"FF",X"00",X"FF",X"80",X"00",X"C0",X"01",X"1F",X"FF",X"80",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"01",X"9F",X"FF",X"00",X"00",X"00",X"FF",X"00",X"FF",X"80",
		X"FF",X"01",X"00",X"00",X"01",X"1F",X"01",X"9F",X"FF",X"01",X"00",X"00",X"FF",X"00",X"FF",X"80",
		X"00",X"C0",X"00",X"00",X"FF",X"80",X"FF",X"00",X"00",X"00",X"00",X"00",X"01",X"9F",X"FF",X"01",
		X"00",X"00",X"FF",X"00",X"FF",X"80",X"FF",X"00",X"00",X"00",X"00",X"00",X"01",X"9F",X"FF",X"01",
		X"00",X"00",X"00",X"00",X"FF",X"80",X"00",X"C0",X"00",X"00",X"FF",X"80",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"01",X"9F",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"01",X"9F",X"FF",X"00",X"FF",X"80",
		X"00",X"00",X"01",X"9F",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"80",X"B2",X"00",X"00",X"00",
		X"6E",X"01",X"01",X"9F",X"00",X"C0",X"FF",X"00",X"FF",X"80",X"00",X"00",X"01",X"1F",X"FF",X"00",
		X"FF",X"80",X"00",X"00",X"01",X"9F",X"FF",X"00",X"FF",X"00",X"00",X"00",X"01",X"9F",X"FF",X"00",
		X"FF",X"80",X"FF",X"00",X"01",X"9F",X"B2",X"00",X"00",X"00",X"B0",X"1E",X"FF",X"80",X"00",X"C0",
		X"FF",X"00",X"FF",X"80",X"FF",X"00",X"01",X"9F",X"60",X"01",X"00",X"00",X"B0",X"1E",X"FF",X"80",
		X"D4",X"1E",X"FF",X"80",X"00",X"C0",X"C0",X"01",X"FF",X"80",X"00",X"00",X"01",X"9F",X"FF",X"00",
		X"FF",X"80",X"00",X"C0",X"00",X"00",X"80",X"80",X"C0",X"00",X"80",X"80",X"00",X"C0",X"FF",X"01",
		X"FF",X"80",X"00",X"C0",X"00",X"00",X"FF",X"80",X"80",X"1D",X"00",X"00",X"00",X"00",X"01",X"9F",
		X"40",X"1E",X"FF",X"80",X"00",X"C0",X"00",X"00",X"FF",X"80",X"C0",X"01",X"01",X"1F",X"C0",X"01",
		X"FF",X"80",X"C0",X"00",X"01",X"9F",X"00",X"C0",X"40",X"1E",X"FF",X"80",X"00",X"C0",X"FF",X"00",
		X"FF",X"80",X"C0",X"00",X"00",X"00",X"FF",X"00",X"01",X"9F",X"00",X"00",X"FF",X"80",X"FF",X"00",
		X"01",X"9F",X"00",X"00",X"FF",X"80",X"00",X"C0",X"00",X"00",X"FF",X"80",X"C0",X"00",X"01",X"1F",
		X"00",X"00",X"FF",X"80",X"60",X"00",X"00",X"00",X"00",X"00",X"60",X"9F",X"A0",X"00",X"A0",X"80",
		X"FF",X"00",X"01",X"1F",X"00",X"00",X"FF",X"80",X"C0",X"01",X"01",X"9F",X"80",X"00",X"80",X"80",
		X"00",X"00",X"80",X"80",X"00",X"C0",X"00",X"00",X"FF",X"80",X"C0",X"00",X"01",X"1F",X"00",X"00",
		X"FF",X"80",X"60",X"00",X"00",X"00",X"00",X"00",X"01",X"9F",X"A0",X"00",X"00",X"00",X"FF",X"00",
		X"FF",X"80",X"80",X"00",X"00",X"00",X"C0",X"01",X"01",X"9F",X"00",X"C0",X"00",X"00",X"FF",X"80",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"01",X"9F",X"60",X"00",X"00",X"00",X"00",X"00",X"FF",X"80",
		X"80",X"00",X"00",X"00",X"20",X"01",X"01",X"9F",X"80",X"00",X"00",X"00",X"01",X"1F",X"FF",X"80",
		X"00",X"C0",X"00",X"00",X"FF",X"80",X"C0",X"00",X"01",X"1F",X"00",X"00",X"60",X"80",X"60",X"00",
		X"A0",X"9F",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"1F",X"80",X"80",X"A0",X"1F",
		X"A0",X"9F",X"00",X"00",X"60",X"80",X"80",X"01",X"00",X"00",X"00",X"00",X"01",X"9F",X"00",X"C0",
		X"00",X"00",X"FF",X"80",X"C0",X"00",X"01",X"1F",X"00",X"00",X"FF",X"80",X"80",X"01",X"01",X"9F",
		X"00",X"C0",X"00",X"00",X"80",X"80",X"80",X"1F",X"80",X"80",X"00",X"C0",X"01",X"1F",X"FF",X"80",
		X"00",X"02",X"01",X"1F",X"00",X"00",X"FF",X"80",X"01",X"1F",X"01",X"9F",X"00",X"C0",X"00",X"00",
		X"FF",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"9F",X"80",X"1F",X"80",X"9F",X"FF",X"00",
		X"00",X"00",X"60",X"00",X"FF",X"80",X"20",X"01",X"00",X"00",X"80",X"1F",X"80",X"9F",X"00",X"00",
		X"80",X"9F",X"FF",X"00",X"FF",X"80",X"00",X"C0",X"00",X"00",X"FF",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"01",X"9F",X"E0",X"00",X"00",X"00",X"A0",X"1F",X"FF",X"80",X"80",X"00",X"00",X"00",
		X"FF",X"00",X"01",X"9F",X"80",X"00",X"00",X"00",X"00",X"00",X"FF",X"80",X"00",X"C0",X"00",X"00",
		X"FF",X"80",X"80",X"00",X"01",X"1F",X"E0",X"00",X"FF",X"80",X"40",X"00",X"C0",X"9F",X"60",X"1F",
		X"40",X"9F",X"80",X"00",X"00",X"00",X"FF",X"00",X"FF",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"01",X"9F",X"00",X"C0",X"00",X"00",X"FF",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"01",X"9F",
		X"FF",X"00",X"FF",X"80",X"FF",X"00",X"01",X"9F",X"80",X"00",X"00",X"00",X"00",X"00",X"FF",X"80",
		X"00",X"C0",X"C0",X"00",X"FF",X"80",X"C0",X"00",X"00",X"00",X"01",X"1F",X"01",X"9F",X"80",X"02",
		X"00",X"00",X"00",X"00",X"FF",X"80",X"00",X"C0",X"00",X"00",X"FF",X"80",X"C0",X"00",X"00",X"00",
		X"80",X"00",X"80",X"9F",X"80",X"1F",X"80",X"9F",X"80",X"01",X"00",X"00",X"00",X"00",X"FF",X"80",
		X"00",X"C0",X"00",X"00",X"40",X"80",X"C0",X"00",X"C0",X"80",X"C0",X"00",X"00",X"00",X"40",X"1F",
		X"40",X"9F",X"00",X"00",X"C0",X"9F",X"80",X"01",X"00",X"00",X"00",X"00",X"FF",X"80",X"00",X"C0",
		X"00",X"00",X"FF",X"80",X"C0",X"00",X"00",X"00",X"00",X"00",X"01",X"9F",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"80",X"00",X"C0",X"01",X"1F",X"FF",X"80",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"9F",X"C0",X"00",X"40",X"9F",X"C0",X"00",X"00",X"00",X"00",X"00",X"FF",X"80",X"00",X"C0",
		X"00",X"00",X"FF",X"80",X"FF",X"00",X"01",X"1F",X"C0",X"00",X"C0",X"80",X"00",X"00",X"40",X"80",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"01",X"9F",X"00",X"C0",X"00",X"00",X"FF",X"80",X"FF",X"00",
		X"00",X"00",X"C0",X"00",X"40",X"9F",X"00",X"00",X"C0",X"9F",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"80",X"00",X"C0",X"FF",X"00",X"FF",X"80",X"40",X"00",X"00",X"00",X"80",X"1F",X"80",X"9F",
		X"80",X"00",X"80",X"9F",X"FF",X"00",X"00",X"00",X"80",X"1F",X"80",X"80",X"80",X"00",X"80",X"80",
		X"80",X"01",X"00",X"00",X"00",X"00",X"01",X"9F",X"00",X"C0",X"FF",X"00",X"FF",X"80",X"80",X"1F",
		X"01",X"1F",X"40",X"00",X"40",X"80",X"00",X"00",X"C0",X"9F",X"FF",X"00",X"00",X"00",X"80",X"00",
		X"80",X"80",X"80",X"1F",X"80",X"80",X"80",X"01",X"00",X"00",X"00",X"00",X"01",X"9F",X"00",X"C0",
		X"E0",X"00",X"E0",X"80",X"60",X"00",X"A0",X"9F",X"80",X"1F",X"80",X"9F",X"80",X"01",X"00",X"00",
		X"00",X"00",X"FF",X"80",X"00",X"C0",X"01",X"1F",X"FF",X"80",X"00",X"03",X"00",X"00",X"00",X"1E",
		X"01",X"9F",X"00",X"03",X"FF",X"00",X"FF",X"00",X"01",X"9F",X"FF",X"00",X"FF",X"80",X"00",X"C0",
		X"01",X"1F",X"FF",X"80",X"00",X"02",X"00",X"00",X"00",X"02",X"01",X"9F",X"FF",X"00",X"00",X"00",
		X"80",X"1F",X"FF",X"80",X"80",X"02",X"01",X"1F",X"FF",X"00",X"FF",X"80",X"00",X"C0",X"00",X"00",
		X"FF",X"80",X"FF",X"00",X"80",X"9F",X"00",X"00",X"80",X"80",X"FF",X"00",X"01",X"1F",X"00",X"02",
		X"FF",X"80",X"80",X"00",X"01",X"9F",X"80",X"01",X"FF",X"00",X"00",X"00",X"01",X"9F",X"FF",X"00",
		X"FF",X"80",X"FF",X"00",X"00",X"00",X"00",X"00",X"01",X"9F",X"00",X"C0",X"00",X"00",X"FF",X"80",
		X"00",X"05",X"01",X"1F",X"FF",X"00",X"FF",X"80",X"00",X"00",X"01",X"1F",X"FF",X"00",X"FF",X"80",
		X"00",X"00",X"01",X"9F",X"00",X"C0",X"01",X"1F",X"FF",X"80",X"00",X"03",X"00",X"00",X"00",X"02",
		X"00",X"80",X"01",X"1F",X"01",X"9F",X"01",X"1F",X"FF",X"80",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"01",X"9F",X"00",X"03",X"00",X"00",X"FF",X"00",X"80",X"80",X"FF",X"00",X"80",X"9F",X"00",X"C0",
		X"FF",X"00",X"FF",X"80",X"00",X"02",X"01",X"1F",X"FF",X"00",X"FF",X"80",X"00",X"00",X"01",X"9F",
		X"FF",X"00",X"00",X"00",X"01",X"1F",X"FF",X"80",X"00",X"03",X"00",X"00",X"FF",X"00",X"80",X"9F",
		X"FF",X"00",X"80",X"80",X"00",X"C0",X"00",X"00",X"FF",X"80",X"00",X"05",X"00",X"00",X"FF",X"00",
		X"01",X"9F",X"00",X"00",X"FF",X"00",X"FF",X"00",X"01",X"9F",X"00",X"00",X"FF",X"80",X"00",X"C0",
		X"00",X"00",X"80",X"80",X"01",X"1F",X"80",X"9F",X"00",X"00",X"FF",X"80",X"00",X"02",X"00",X"00",
		X"00",X"02",X"01",X"9F",X"80",X"00",X"FF",X"80",X"80",X"01",X"01",X"1F",X"00",X"00",X"FF",X"80",
		X"FF",X"00",X"01",X"9F",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"80",X"00",X"C0",X"FF",X"00",
		X"FF",X"80",X"FF",X"00",X"01",X"1F",X"00",X"02",X"FF",X"80",X"80",X"00",X"01",X"1F",X"80",X"00",
		X"FF",X"80",X"00",X"02",X"00",X"00",X"FF",X"00",X"01",X"9F",X"00",X"C0",X"FF",X"00",X"FF",X"80",
		X"00",X"02",X"01",X"9F",X"FF",X"00",X"00",X"00",X"FF",X"00",X"FF",X"80",X"FF",X"00",X"01",X"9F",
		X"00",X"C0",X"00",X"00",X"FF",X"80",X"80",X"00",X"01",X"1F",X"00",X"00",X"FF",X"80",X"80",X"00",
		X"80",X"9F",X"00",X"00",X"80",X"9F",X"FF",X"00",X"00",X"00",X"FF",X"00",X"FF",X"80",X"80",X"00",
		X"01",X"1F",X"FF",X"00",X"FF",X"80",X"00",X"C0",X"00",X"00",X"FF",X"80",X"80",X"00",X"00",X"00",
		X"FF",X"00",X"01",X"9F",X"00",X"00",X"FF",X"80",X"80",X"00",X"00",X"00",X"FF",X"00",X"01",X"9F",
		X"80",X"01",X"00",X"00",X"01",X"1F",X"FF",X"80",X"00",X"C0",X"00",X"00",X"FF",X"80",X"80",X"00",
		X"00",X"00",X"00",X"00",X"01",X"9F",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"80",X"80",X"00",
		X"01",X"1F",X"FF",X"00",X"FF",X"80",X"80",X"00",X"01",X"1F",X"FF",X"00",X"FF",X"80",X"00",X"C0",
		X"00",X"00",X"FF",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"01",X"9F",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"80",X"80",X"00",X"00",X"00",X"FF",X"00",X"01",X"9F",X"80",X"01",X"00",X"00",
		X"01",X"1F",X"FF",X"80",X"00",X"C0",X"00",X"00",X"FF",X"80",X"80",X"00",X"01",X"1F",X"FF",X"00",
		X"FF",X"80",X"00",X"00",X"01",X"1F",X"FF",X"00",X"FF",X"80",X"80",X"00",X"00",X"00",X"01",X"1F",
		X"01",X"9F",X"80",X"01",X"00",X"00",X"FF",X"00",X"FF",X"80",X"00",X"C0",X"00",X"00",X"FF",X"80",
		X"80",X"02",X"00",X"00",X"01",X"1F",X"01",X"9F",X"FF",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"80",X"00",X"80",X"9F",X"80",X"01",X"00",X"00",X"01",X"1F",X"FF",X"80",X"00",X"C0",X"00",X"00",
		X"FF",X"80",X"FF",X"00",X"00",X"00",X"00",X"00",X"01",X"9F",X"FF",X"00",X"FF",X"80",X"80",X"00",
		X"01",X"1F",X"FF",X"00",X"FF",X"80",X"00",X"00",X"01",X"9F",X"00",X"C0",X"00",X"00",X"FF",X"80",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"01",X"9F",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"80",
		X"00",X"C0",X"00",X"00",X"FF",X"80",X"FF",X"00",X"01",X"1F",X"00",X"00",X"FF",X"80",X"FF",X"00",
		X"01",X"9F",X"80",X"00",X"FF",X"00",X"FF",X"00",X"01",X"9F",X"FF",X"00",X"FF",X"80",X"00",X"C0",
		X"00",X"00",X"FF",X"80",X"80",X"01",X"00",X"00",X"FF",X"00",X"01",X"9F",X"00",X"02",X"00",X"00",
		X"01",X"1F",X"FF",X"80",X"00",X"C0",X"00",X"00",X"FF",X"80",X"80",X"00",X"00",X"00",X"FF",X"00",
		X"01",X"9F",X"00",X"00",X"FF",X"00",X"80",X"00",X"01",X"9F",X"00",X"00",X"FF",X"80",X"80",X"01",
		X"01",X"1F",X"FF",X"00",X"FF",X"80",X"00",X"C0",X"00",X"00",X"FF",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"01",X"9F",X"80",X"00",X"FF",X"00",X"80",X"00",X"01",X"9F",X"80",X"00",X"00",X"00",
		X"FF",X"00",X"FF",X"80",X"80",X"00",X"00",X"00",X"FF",X"00",X"01",X"9F",X"00",X"C0",X"00",X"00",
		X"FF",X"80",X"80",X"00",X"01",X"1F",X"00",X"00",X"FF",X"80",X"80",X"00",X"01",X"9F",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"01",X"9F",X"80",X"00",X"00",X"00",X"FF",X"00",X"FF",X"80",X"00",X"C0",
		X"00",X"00",X"FF",X"80",X"80",X"00",X"00",X"00",X"80",X"00",X"01",X"9F",X"FF",X"00",X"FF",X"80",
		X"00",X"00",X"01",X"1F",X"FF",X"00",X"FF",X"80",X"80",X"00",X"00",X"00",X"FF",X"00",X"01",X"9F",
		X"00",X"C0",X"00",X"00",X"FF",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"01",X"9F",X"80",X"00",
		X"FF",X"00",X"FF",X"00",X"01",X"9F",X"00",X"00",X"FF",X"00",X"FF",X"00",X"01",X"9F",X"80",X"00",
		X"00",X"00",X"FF",X"00",X"FF",X"80",X"00",X"C0",X"00",X"00",X"FF",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"01",X"9F",X"80",X"00",X"00",X"00",X"00",X"00",X"FF",X"80",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"01",X"9F",X"80",X"01",X"FF",X"00",X"FF",X"00",X"01",X"9F",X"00",X"C0",X"00",X"00",
		X"FF",X"80",X"C0",X"00",X"A0",X"9F",X"A0",X"00",X"60",X"9F",X"00",X"00",X"FF",X"80",X"00",X"C0",
		X"00",X"00",X"FF",X"80",X"60",X"01",X"01",X"1F",X"00",X"00",X"FF",X"80",X"60",X"1F",X"60",X"9F",
		X"40",X"1F",X"A0",X"9F",X"00",X"C0",X"00",X"00",X"FF",X"80",X"00",X"02",X"01",X"1F",X"00",X"00",
		X"FF",X"80",X"A0",X"1F",X"A0",X"9F",X"C0",X"1F",X"E0",X"9F",X"40",X"00",X"E0",X"9F",X"60",X"00",
		X"A0",X"9F",X"00",X"C0",X"00",X"00",X"FF",X"80",X"40",X"00",X"E0",X"9F",X"60",X"00",X"A0",X"9F",
		X"00",X"00",X"80",X"80",X"60",X"02",X"01",X"1F",X"00",X"00",X"FF",X"80",X"A0",X"1F",X"A0",X"9F",
		X"C0",X"1F",X"E0",X"9F",X"40",X"00",X"E0",X"9F",X"60",X"00",X"A0",X"9F",X"00",X"C0",X"00",X"00",
		X"FF",X"80",X"A0",X"00",X"01",X"1F",X"00",X"00",X"80",X"80",X"A0",X"1F",X"A0",X"9F",X"C0",X"1F",
		X"E0",X"9F",X"00",X"C0",X"00",X"00",X"FF",X"80",X"A0",X"00",X"00",X"00",X"00",X"00",X"01",X"9F",
		X"A0",X"1F",X"60",X"80",X"C0",X"1F",X"20",X"80",X"40",X"00",X"20",X"80",X"60",X"00",X"60",X"80",
		X"80",X"01",X"00",X"00",X"C0",X"00",X"A0",X"9F",X"A0",X"00",X"60",X"9F",X"00",X"00",X"FF",X"80",
		X"00",X"C0",X"00",X"00",X"FF",X"80",X"20",X"02",X"01",X"1F",X"C0",X"00",X"60",X"80",X"A0",X"00",
		X"A0",X"80",X"00",X"00",X"01",X"9F",X"00",X"C0",X"00",X"00",X"FF",X"80",X"00",X"03",X"00",X"00",
		X"00",X"00",X"01",X"9F",X"A0",X"1F",X"60",X"80",X"C0",X"1F",X"20",X"80",X"40",X"00",X"20",X"80",
		X"60",X"00",X"60",X"80",X"00",X"C0",X"00",X"00",X"FF",X"80",X"A0",X"00",X"00",X"00",X"00",X"00",
		X"01",X"9F",X"A0",X"1F",X"60",X"80",X"C0",X"1F",X"20",X"80",X"40",X"00",X"20",X"80",X"60",X"00",
		X"60",X"80",X"00",X"C0",X"00",X"00",X"FF",X"80",X"FF",X"00",X"00",X"00",X"C0",X"00",X"A0",X"9F",
		X"A0",X"00",X"60",X"9F",X"00",X"00",X"FF",X"80",X"00",X"C0",X"00",X"00",X"FF",X"80",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"01",X"9F",X"A0",X"1F",X"60",X"80",X"C0",X"1F",X"20",X"80",X"40",X"00",
		X"20",X"80",X"60",X"00",X"60",X"80",X"20",X"00",X"01",X"1F",X"C0",X"00",X"60",X"80",X"A0",X"00",
		X"A0",X"80",X"00",X"00",X"01",X"9F",X"00",X"C0",X"00",X"00",X"C0",X"1F",X"00",X"00",X"20",X"80",
		X"E0",X"1F",X"10",X"80",X"E0",X"1F",X"F0",X"9F",X"00",X"C0",X"2C",X"AC",X"38",X"00",X"04",X"00",
		X"8C",X"48",X"84",X"58",X"94",X"58",X"00",X"C0",X"D8",X"1F",X"10",X"00",X"9C",X"4C",X"88",X"4C",
		X"8C",X"44",X"00",X"C0",X"3C",X"AC",X"12",X"5A",X"98",X"42",X"9E",X"5C",X"86",X"5A",X"00",X"C0",
		X"EC",X"1F",X"CC",X"1F",X"8C",X"44",X"88",X"4C",X"9C",X"4C",X"00",X"C0",X"48",X"AC",X"02",X"52",
		X"88",X"5C",X"9C",X"58",X"98",X"44",X"00",X"C0",X"00",X"00",X"C0",X"1F",X"8C",X"40",X"E0",X"1F",
		X"10",X"80",X"9C",X"54",X"00",X"C0",X"54",X"AC",X"20",X"00",X"04",X"80",X"8A",X"46",X"9C",X"46",
		X"96",X"5E",X"00",X"C0",X"40",X"00",X"E0",X"1F",X"E0",X"1F",X"10",X"80",X"E0",X"1F",X"F0",X"9F",
		X"00",X"00",X"E0",X"9F",X"00",X"C0",X"62",X"AC",X"08",X"00",X"24",X"00",X"8C",X"5A",X"84",X"48",
		X"94",X"48",X"00",X"C0",X"C0",X"1F",X"00",X"00",X"28",X"00",X"00",X"80",X"8C",X"4A",X"F4",X"1F",
		X"28",X"80",X"00",X"C0",X"72",X"AC",X"08",X"00",X"D4",X"1F",X"9A",X"48",X"98",X"5A",X"86",X"58",
		X"00",X"C0",X"F0",X"1F",X"C8",X"1F",X"08",X"00",X"20",X"80",X"E8",X"1F",X"20",X"80",X"E0",X"1F",
		X"08",X"80",X"00",X"C0",X"81",X"AC",X"28",X"00",X"F0",X"1F",X"84",X"4A",X"9C",X"42",X"98",X"5A",
		X"00",X"C0",X"C0",X"1F",X"20",X"00",X"20",X"00",X"F0",X"9F",X"20",X"00",X"10",X"80",X"00",X"00",
		X"20",X"80",X"00",X"C0",X"91",X"AC",X"F8",X"1F",X"DC",X"1F",X"94",X"46",X"9C",X"5C",X"8C",X"56",
		X"00",X"C0",X"40",X"00",X"E0",X"1F",X"D0",X"1F",X"10",X"80",X"00",X"00",X"20",X"80",X"30",X"00",
		X"10",X"80",X"00",X"C0",X"A1",X"AC",X"D0",X"1F",X"E8",X"1F",X"80",X"58",X"98",X"40",X"80",X"48",
		X"00",X"C0",X"C0",X"1F",X"E0",X"1F",X"30",X"00",X"10",X"80",X"00",X"00",X"20",X"80",X"D0",X"1F",
		X"10",X"80",X"00",X"C0",X"B1",X"AC",X"30",X"00",X"E8",X"1F",X"80",X"48",X"98",X"40",X"80",X"58",
		X"00",X"C0",X"00",X"00",X"C0",X"1F",X"00",X"00",X"20",X"80",X"20",X"00",X"20",X"80",X"20",X"00",
		X"00",X"80",X"00",X"C0",X"C1",X"AC",X"D8",X"1F",X"F8",X"1F",X"88",X"58",X"98",X"58",X"98",X"48",
		X"00",X"C0",X"C0",X"1F",X"00",X"00",X"20",X"00",X"00",X"80",X"20",X"00",X"20",X"80",X"00",X"00",
		X"20",X"80",X"00",X"C0",X"D1",X"AC",X"F8",X"1F",X"D8",X"1F",X"98",X"48",X"98",X"58",X"88",X"58",
		X"00",X"C0",X"00",X"00",X"C0",X"1F",X"00",X"00",X"20",X"80",X"E0",X"1F",X"20",X"80",X"E0",X"1F",
		X"00",X"80",X"00",X"C0",X"E1",X"AC",X"28",X"00",X"F8",X"1F",X"88",X"48",X"98",X"48",X"98",X"58",
		X"00",X"C0",X"40",X"00",X"F8",X"1F",X"E0",X"1F",X"00",X"80",X"E0",X"1F",X"20",X"80",X"00",X"00",
		X"20",X"80",X"00",X"C0",X"F1",X"AC",X"08",X"00",X"D8",X"1F",X"98",X"58",X"98",X"48",X"88",X"48",
		X"00",X"C0",X"20",X"00",X"20",X"00",X"98",X"58",X"E0",X"1F",X"10",X"80",X"F0",X"1F",X"20",X"80",
		X"00",X"C0",X"01",X"AD",X"18",X"00",X"DC",X"1F",X"96",X"5E",X"9C",X"46",X"8A",X"46",X"00",X"C0",
		X"00",X"00",X"40",X"00",X"94",X"40",X"98",X"54",X"84",X"54",X"00",X"C0",X"10",X"AD",X"1E",X"4E",
		X"98",X"46",X"82",X"44",X"8A",X"5E",X"00",X"C0",X"E8",X"1F",X"C8",X"1F",X"8C",X"46",X"EC",X"1F",
		X"30",X"80",X"84",X"54",X"00",X"C0",X"1C",X"AD",X"18",X"4E",X"80",X"4C",X"98",X"44",X"98",X"56",
		X"00",X"C0",X"F8",X"1F",X"50",X"00",X"04",X"00",X"DC",X"9F",X"28",X"00",X"E0",X"9F",X"24",X"00",
		X"04",X"80",X"00",X"C0",X"29",X"AD",X"D4",X"1F",X"04",X"00",X"98",X"54",X"84",X"5C",X"8C",X"44",
		X"00",X"C0",X"F8",X"1F",X"38",X"00",X"92",X"42",X"20",X"00",X"E8",X"9F",X"82",X"4E",X"00",X"C0",
		X"39",X"AD",X"24",X"00",X"04",X"00",X"98",X"58",X"84",X"5C",X"88",X"44",X"00",X"C0",X"E0",X"1F",
		X"00",X"E0",X"00",X"00",X"20",X"E0",X"20",X"00",X"00",X"E0",X"00",X"C0",X"20",X"00",X"00",X"E0",
		X"00",X"00",X"20",X"E0",X"E0",X"1F",X"00",X"E0",X"00",X"C0",X"8E",X"3A",X"9C",X"3A",X"D0",X"00",
		X"E0",X"1F",X"FC",X"1F",X"FB",X"1F",X"04",X"C0",X"05",X"00",X"04",X"C0",X"F7",X"1F",X"F3",X"1F",
		X"00",X"C0",X"E1",X"1F",X"F5",X"1F",X"FA",X"1F",X"03",X"C0",X"05",X"00",X"05",X"C0",X"0C",X"00",
		X"F5",X"1F",X"00",X"C0",X"18",X"52",X"F9",X"1F",X"02",X"C0",X"04",X"00",X"05",X"C0",X"1A",X"47",
		X"00",X"C0",X"E8",X"1F",X"EB",X"1F",X"F9",X"1F",X"00",X"C0",X"02",X"00",X"07",X"C0",X"11",X"00",
		X"F7",X"1F",X"00",X"C0",X"13",X"56",X"F9",X"1F",X"00",X"C0",X"01",X"00",X"06",X"C0",X"13",X"00",
		X"FA",X"1F",X"00",X"C0",X"F1",X"1F",X"E3",X"1F",X"DF",X"5D",X"00",X"00",X"07",X"C0",X"ED",X"1F",
		X"FE",X"1F",X"00",X"C0",X"F7",X"1F",X"E1",X"1F",X"FD",X"1F",X"FA",X"DF",X"FF",X"1F",X"07",X"C0",
		X"13",X"00",X"01",X"00",X"00",X"C0",X"FD",X"1F",X"E0",X"1F",X"FB",X"1F",X"FB",X"DF",X"FD",X"1F",
		X"06",X"C0",X"13",X"00",X"05",X"00",X"00",X"C0",X"04",X"00",X"E0",X"1F",X"FC",X"1F",X"FB",X"DF",
		X"FC",X"1F",X"05",X"C0",X"0D",X"00",X"09",X"00",X"00",X"C0",X"0B",X"00",X"E1",X"1F",X"FD",X"1F",
		X"FA",X"DF",X"FB",X"1F",X"05",X"C0",X"0B",X"00",X"0C",X"00",X"00",X"C0",X"12",X"48",X"FE",X"1F",
		X"F9",X"DF",X"FB",X"1F",X"04",X"C0",X"07",X"46",X"00",X"C0",X"15",X"00",X"E8",X"1F",X"00",X"00",
		X"F9",X"DF",X"F9",X"1F",X"02",X"C0",X"09",X"00",X"11",X"00",X"00",X"C0",X"16",X"4D",X"00",X"00",
		X"F9",X"DF",X"FA",X"1F",X"01",X"C0",X"06",X"00",X"13",X"00",X"00",X"C0",X"1D",X"00",X"F1",X"1F",
		X"DD",X"41",X"F9",X"1F",X"00",X"C0",X"02",X"00",X"ED",X"1F",X"00",X"C0",X"1F",X"00",X"F7",X"1F",
		X"06",X"00",X"FD",X"DF",X"F9",X"1F",X"FF",X"DF",X"FF",X"1F",X"13",X"00",X"00",X"C0",X"20",X"00",
		X"FD",X"1F",X"05",X"00",X"FB",X"DF",X"FA",X"1F",X"FD",X"DF",X"FB",X"1F",X"13",X"00",X"00",X"C0",
		X"20",X"00",X"04",X"00",X"05",X"00",X"FC",X"DF",X"FB",X"1F",X"FC",X"DF",X"F7",X"1F",X"0D",X"00",
		X"00",X"C0",X"1F",X"00",X"0B",X"00",X"06",X"00",X"FD",X"DF",X"FB",X"1F",X"FB",X"DF",X"F4",X"1F",
		X"0B",X"00",X"00",X"C0",X"08",X"4E",X"07",X"00",X"FE",X"DF",X"FC",X"1F",X"FB",X"DF",X"06",X"59",
		X"00",X"C0",X"18",X"00",X"15",X"00",X"07",X"00",X"00",X"C0",X"FE",X"1F",X"F9",X"DF",X"EF",X"1F",
		X"09",X"00",X"00",X"C0",X"0D",X"4A",X"07",X"00",X"00",X"C0",X"FF",X"1F",X"FA",X"DF",X"ED",X"1F",
		X"06",X"00",X"00",X"C0",X"0F",X"00",X"1D",X"00",X"C1",X"43",X"00",X"00",X"F9",X"DF",X"13",X"00",
		X"02",X"00",X"00",X"C0",X"09",X"00",X"1F",X"00",X"03",X"00",X"06",X"C0",X"01",X"00",X"F9",X"DF",
		X"ED",X"1F",X"FF",X"1F",X"00",X"C0",X"03",X"00",X"20",X"00",X"05",X"00",X"05",X"C0",X"03",X"00",
		X"FA",X"DF",X"ED",X"1F",X"FB",X"1F",X"00",X"C0",X"FC",X"1F",X"20",X"00",X"04",X"00",X"05",X"C0",
		X"04",X"00",X"FB",X"DF",X"F3",X"1F",X"F7",X"1F",X"00",X"C0",X"F5",X"1F",X"1F",X"00",X"03",X"00",
		X"06",X"C0",X"05",X"00",X"FB",X"DF",X"F5",X"1F",X"F4",X"1F",X"00",X"C0",X"0E",X"58",X"02",X"00",
		X"07",X"C0",X"05",X"00",X"FC",X"DF",X"1A",X"54",X"00",X"C0",X"EB",X"1F",X"18",X"00",X"00",X"00",
		X"07",X"C0",X"07",X"00",X"FE",X"DF",X"F7",X"1F",X"EF",X"1F",X"00",X"C0",X"0A",X"53",X"00",X"00",
		X"07",X"C0",X"06",X"00",X"FF",X"DF",X"FA",X"1F",X"ED",X"1F",X"00",X"C0",X"E3",X"1F",X"0F",X"00",
		X"C3",X"5F",X"07",X"00",X"00",X"C0",X"FE",X"1F",X"13",X"00",X"00",X"C0",X"E1",X"1F",X"09",X"00",
		X"FA",X"1F",X"03",X"C0",X"07",X"00",X"01",X"C0",X"01",X"00",X"ED",X"1F",X"00",X"C0",X"E0",X"1F",
		X"03",X"00",X"FB",X"1F",X"05",X"C0",X"06",X"00",X"03",X"C0",X"05",X"00",X"ED",X"1F",X"00",X"C0",
		X"80",X"1F",X"CC",X"BF",X"80",X"00",X"4C",X"00",X"80",X"1F",X"34",X"A0",X"00",X"C0",X"80",X"00",
		X"34",X"A0",X"80",X"1F",X"B4",X"1F",X"80",X"00",X"CC",X"BF",X"00",X"C0",X"40",X"80",X"00",X"1F",
		X"00",X"02",X"E0",X"1F",X"60",X"E0",X"E0",X"1F",X"A0",X"FF",X"00",X"00",X"40",X"E0",X"20",X"00",
		X"A0",X"FF",X"20",X"00",X"60",X"E0",X"E0",X"1F",X"20",X"E0",X"E0",X"1F",X"E0",X"FF",X"00",X"00",
		X"C0",X"FF",X"20",X"00",X"E0",X"FF",X"20",X"00",X"20",X"E0",X"00",X"C0",X"A7",X"64",X"38",X"1F",
		X"CC",X"1F",X"28",X"00",X"0E",X"20",X"0E",X"00",X"28",X"20",X"F2",X"1F",X"28",X"20",X"D8",X"1F",
		X"0E",X"20",X"D8",X"1F",X"F2",X"3F",X"F2",X"1F",X"D8",X"3F",X"0E",X"00",X"D8",X"3F",X"28",X"00",
		X"F2",X"3F",X"00",X"C0",X"08",X"40",X"25",X"4E",X"2E",X"45",X"2E",X"5B",X"25",X"52",X"3B",X"52",
		X"32",X"5B",X"32",X"45",X"3B",X"4E",X"00",X"C0",X"40",X"80",X"8E",X"EE",X"40",X"80",X"8E",X"AE",
		X"A4",X"64",X"A2",X"EE",X"40",X"80",X"8E",X"AE",X"A1",X"64",X"A2",X"EE",X"40",X"80",X"8E",X"AE",
		X"95",X"64",X"A2",X"EE",X"40",X"80",X"8E",X"AE",X"B2",X"64",X"A2",X"EE",X"40",X"80",X"8E",X"AE",
		X"A6",X"64",X"A2",X"EE",X"40",X"80",X"8E",X"AE",X"A3",X"64",X"A2",X"EE",X"C6",X"64",X"C8",X"00",
		X"7C",X"00",X"2A",X"43",X"23",X"4A",X"23",X"56",X"2A",X"5D",X"36",X"5D",X"3D",X"56",X"3D",X"4A",
		X"36",X"43",X"00",X"C0",X"A4",X"64",X"33",X"40",X"1A",X"00",X"34",X"00",X"20",X"4D",X"CC",X"1F",
		X"1A",X"00",X"2D",X"40",X"E6",X"1F",X"CC",X"1F",X"20",X"53",X"34",X"00",X"E6",X"1F",X"00",X"C0",
		X"A4",X"64",X"0A",X"43",X"20",X"00",X"E0",X"3F",X"E0",X"1F",X"2C",X"00",X"20",X"00",X"20",X"20",
		X"D4",X"1F",X"E0",X"1F",X"E0",X"1F",X"20",X"20",X"20",X"00",X"D4",X"1F",X"E0",X"1F",X"E0",X"3F",
		X"00",X"C0",X"40",X"80",X"C6",X"AE",X"D2",X"EE",X"40",X"80",X"C6",X"AE",X"E0",X"EE",X"40",X"80",
		X"C6",X"AE",X"D2",X"AE",X"E0",X"EE",X"40",X"80",X"C6",X"64",X"C8",X"00",X"06",X"1F",X"C9",X"AE",
		X"D2",X"EE",X"40",X"80",X"C6",X"64",X"C8",X"00",X"06",X"1F",X"C9",X"AE",X"E0",X"EE",X"40",X"80",
		X"C6",X"64",X"C8",X"00",X"06",X"1F",X"C9",X"AE",X"D2",X"AE",X"E0",X"EE",X"40",X"80",X"70",X"1E",
		X"40",X"02",X"D6",X"64",X"98",X"EF",X"91",X"64",X"03",X"5A",X"0C",X"00",X"E0",X"3F",X"0C",X"00",
		X"20",X"20",X"00",X"00",X"40",X"20",X"F4",X"1F",X"20",X"20",X"F4",X"1F",X"E0",X"3F",X"0C",X"00",
		X"BA",X"1F",X"00",X"C0",X"91",X"64",X"03",X"46",X"F4",X"1F",X"E0",X"3F",X"F4",X"1F",X"20",X"20",
		X"00",X"00",X"40",X"20",X"0C",X"00",X"20",X"20",X"0C",X"00",X"E0",X"3F",X"00",X"C0",X"0E",X"AF",
		X"13",X"EF",X"0E",X"AF",X"22",X"EF",X"40",X"80",X"84",X"64",X"BC",X"1D",X"8E",X"1D",X"34",X"F2",
		X"62",X"64",X"06",X"49",X"3A",X"43",X"D0",X"1F",X"30",X"20",X"3D",X"45",X"0C",X"00",X"D6",X"1F",
		X"00",X"C0",X"62",X"64",X"0E",X"4B",X"3E",X"46",X"BC",X"1F",X"00",X"20",X"22",X"46",X"12",X"4B",
		X"00",X"C0",X"62",X"64",X"0C",X"00",X"2A",X"00",X"23",X"46",X"D0",X"1F",X"D0",X"3F",X"26",X"43",
		X"1A",X"49",X"00",X"C0",X"62",X"64",X"01",X"5E",X"3A",X"42",X"00",X"00",X"44",X"20",X"3A",X"5E",
		X"00",X"C0",X"33",X"AF",X"41",X"EF",X"33",X"AF",X"49",X"EF",X"33",X"AF",X"52",X"EF",X"33",X"AF",
		X"38",X"EF",X"40",X"80",X"A4",X"64",X"C2",X"01",X"4C",X"1E",X"98",X"EF",X"C7",X"64",X"03",X"5E",
		X"F8",X"1F",X"E0",X"3F",X"2F",X"42",X"22",X"44",X"3E",X"44",X"31",X"42",X"FA",X"1F",X"20",X"20",
		X"1D",X"5E",X"00",X"C0",X"C7",X"64",X"00",X"00",X"22",X"00",X"24",X"40",X"3E",X"46",X"3E",X"5A",
		X"22",X"5A",X"22",X"46",X"1F",X"43",X"23",X"5D",X"3D",X"5D",X"3E",X"40",X"3D",X"43",X"23",X"43",
		X"FA",X"1F",X"DC",X"1F",X"00",X"C0",X"C7",X"64",X"FC",X"1F",X"46",X"00",X"F8",X"1F",X"20",X"20",
		X"31",X"42",X"3E",X"44",X"22",X"44",X"2F",X"42",X"F8",X"1F",X"E0",X"3F",X"00",X"C0",X"61",X"AF",
		X"66",X"AF",X"83",X"EF",X"61",X"AF",X"72",X"EF",X"40",X"80",X"85",X"64",X"F4",X"01",X"1A",X"02",
		X"26",X"4D",X"2D",X"46",X"2D",X"5A",X"26",X"53",X"3A",X"53",X"33",X"5A",X"33",X"46",X"3A",X"4D",
		X"00",X"C0",X"C6",X"64",X"02",X"5C",X"22",X"44",X"3E",X"44",X"01",X"5E",X"39",X"5E",X"27",X"5E",
		X"1D",X"42",X"00",X"C0",X"C4",X"64",X"22",X"00",X"1E",X"00",X"24",X"5E",X"24",X"42",X"1E",X"41",
		X"3E",X"4F",X"3E",X"51",X"E0",X"1F",X"DE",X"1F",X"00",X"C0",X"C1",X"64",X"08",X"00",X"48",X"00",
		X"3E",X"5C",X"22",X"5C",X"1F",X"42",X"27",X"42",X"39",X"42",X"FC",X"1F",X"BA",X"1F",X"00",X"C0",
		X"C7",X"64",X"DE",X"1F",X"1E",X"00",X"24",X"42",X"24",X"5E",X"1E",X"41",X"3E",X"51",X"3E",X"4F",
		X"20",X"00",X"DE",X"1F",X"00",X"C0",X"C6",X"64",X"02",X"5C",X"22",X"44",X"3E",X"44",X"01",X"5E",
		X"31",X"5E",X"2F",X"5E",X"1D",X"42",X"00",X"C0",X"C4",X"64",X"22",X"00",X"1E",X"00",X"24",X"5E",
		X"24",X"42",X"1E",X"41",X"3E",X"47",X"3E",X"59",X"E0",X"1F",X"DE",X"1F",X"00",X"C0",X"C1",X"64",
		X"08",X"00",X"48",X"00",X"3E",X"5C",X"22",X"5C",X"1F",X"42",X"04",X"00",X"22",X"20",X"04",X"00",
		X"DE",X"3F",X"FC",X"1F",X"BA",X"1F",X"00",X"C0",X"C7",X"64",X"DE",X"1F",X"1E",X"00",X"24",X"42",
		X"24",X"5E",X"1E",X"41",X"3E",X"59",X"3E",X"47",X"20",X"00",X"DE",X"1F",X"00",X"C0",X"94",X"AF",
		X"A1",X"AF",X"AA",X"AF",X"B5",X"AF",X"C0",X"EF",X"94",X"AF",X"CB",X"AF",X"D4",X"AF",X"DF",X"AF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
