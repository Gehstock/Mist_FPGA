library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity sol_bg_bits_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of sol_bg_bits_1 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"02",X"20",X"02",X"AA",X"AA",X"AA",X"AA",X"00",X"02",X"00",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"20",X"02",X"AA",X"AA",X"AA",X"AA",X"00",X"02",X"00",X"02",X"00",X"00",
		X"0A",X"88",X"08",X"88",X"08",X"A8",X"00",X"00",X"08",X"00",X"0A",X"A8",X"08",X"00",X"00",X"00",
		X"00",X"00",X"20",X"2A",X"A0",X"AA",X"80",X"A2",X"82",X"82",X"AA",X"82",X"2A",X"02",X"00",X"00",
		X"0A",X"A8",X"02",X"80",X"00",X"A0",X"0A",X"A8",X"00",X"00",X"0A",X"A8",X"08",X"08",X"02",X"A0",
		X"09",X"00",X"29",X"68",X"0A",X"50",X"0A",X"93",X"0A",X"93",X"0A",X"50",X"29",X"68",X"09",X"00",
		X"F3",X"00",X"FC",X"7C",X"35",X"DF",X"04",X"F4",X"04",X"F4",X"35",X"DF",X"FC",X"7C",X"F3",X"00",
		X"43",X"C0",X"3E",X"F4",X"39",X"B5",X"E8",X"6D",X"E8",X"6D",X"39",X"B5",X"3E",X"F4",X"43",X"C0",
		X"00",X"00",X"15",X"42",X"1A",X"D2",X"1E",X"E2",X"06",X"6A",X"1E",X"E2",X"1A",X"D2",X"15",X"42",
		X"00",X"00",X"15",X"42",X"1A",X"D2",X"1E",X"E2",X"06",X"6A",X"1E",X"E2",X"1A",X"D2",X"15",X"42",
		X"05",X"01",X"0C",X"05",X"00",X"75",X"33",X"F0",X"3C",X"30",X"00",X"75",X"0C",X"05",X"05",X"01",
		X"FF",X"0C",X"C3",X"F3",X"CF",X"FF",X"FF",X"3F",X"FF",X"3F",X"CF",X"FF",X"C3",X"F3",X"FF",X"0C",
		X"00",X"FF",X"03",X"FC",X"1D",X"70",X"55",X"C0",X"55",X"C0",X"1D",X"70",X"03",X"FC",X"00",X"FF",
		X"55",X"25",X"05",X"A0",X"00",X"00",X"01",X"43",X"01",X"43",X"00",X"00",X"05",X"A0",X"55",X"25",
		X"00",X"00",X"2A",X"A8",X"A0",X"2A",X"E2",X"A0",X"8A",X"B0",X"E2",X"A0",X"A0",X"2A",X"2A",X"A8",
		X"00",X"00",X"00",X"40",X"4F",X"28",X"9F",X"03",X"5C",X"C0",X"9F",X"03",X"4F",X"28",X"00",X"40",
		X"F0",X"0F",X"C0",X"03",X"CF",X"F3",X"CC",X"33",X"CC",X"33",X"CF",X"F3",X"C0",X"03",X"F0",X"0F",
		X"0E",X"B0",X"3A",X"AC",X"EB",X"EB",X"AD",X"7A",X"AD",X"7A",X"EB",X"EB",X"3A",X"AC",X"0E",X"B0",
		X"2A",X"A2",X"0A",X"A8",X"02",X"00",X"0A",X"08",X"0A",X"08",X"02",X"00",X"0A",X"A8",X"2A",X"A2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"31",X"00",X"05",X"42",X"04",X"87",X"56",X"54",X"56",X"54",X"04",X"84",X"05",X"42",X"31",X"00",
		X"C0",X"F1",X"F3",X"D4",X"0F",X"D1",X"FF",X"55",X"0F",X"D1",X"F3",X"D4",X"C0",X"F1",X"00",X"00",
		X"03",X"3F",X"3F",X"FF",X"3F",X"FC",X"FD",X"FC",X"FD",X"FC",X"3F",X"FC",X"3F",X"FF",X"03",X"3F",
		X"03",X"F0",X"F3",X"D6",X"33",X"58",X"3D",X"E0",X"3D",X"E0",X"33",X"58",X"F3",X"D6",X"03",X"F0",
		X"05",X"48",X"14",X"21",X"DB",X"11",X"E2",X"0C",X"DB",X"11",X"14",X"21",X"05",X"48",X"00",X"00",
		X"F4",X"50",X"5E",X"D0",X"1C",X"F0",X"02",X"5F",X"02",X"5F",X"1C",X"F0",X"5E",X"D0",X"F4",X"50",
		X"FC",X"3F",X"FD",X"7E",X"7D",X"79",X"17",X"D4",X"17",X"D4",X"7D",X"79",X"FD",X"7E",X"FC",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"15",X"50",X"55",X"54",X"40",X"04",X"40",X"04",X"55",X"54",X"15",X"50",X"00",X"00",
		X"00",X"00",X"00",X"04",X"10",X"04",X"55",X"54",X"55",X"54",X"00",X"04",X"00",X"04",X"00",X"00",
		X"00",X"00",X"10",X"54",X"51",X"54",X"51",X"04",X"51",X"04",X"55",X"14",X"14",X"14",X"00",X"00",
		X"00",X"00",X"50",X"50",X"40",X"54",X"44",X"04",X"44",X"04",X"51",X"54",X"51",X"50",X"00",X"00",
		X"00",X"00",X"05",X"40",X"15",X"40",X"00",X"40",X"00",X"40",X"55",X"54",X"55",X"54",X"00",X"00",
		X"00",X"00",X"55",X"10",X"55",X"14",X"44",X"04",X"44",X"04",X"45",X"54",X"45",X"50",X"00",X"00",
		X"00",X"00",X"15",X"50",X"55",X"54",X"41",X"04",X"41",X"04",X"51",X"54",X"10",X"50",X"00",X"00",
		X"00",X"00",X"50",X"00",X"50",X"00",X"40",X"54",X"41",X"54",X"55",X"00",X"54",X"00",X"00",X"00",
		X"00",X"00",X"11",X"50",X"55",X"54",X"45",X"04",X"45",X"04",X"55",X"54",X"11",X"50",X"00",X"00",
		X"00",X"00",X"14",X"10",X"55",X"14",X"41",X"04",X"41",X"04",X"55",X"54",X"15",X"50",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"55",X"54",X"55",X"54",X"50",X"40",X"50",X"40",X"55",X"54",X"15",X"54",X"00",X"00",
		X"00",X"00",X"55",X"54",X"55",X"54",X"44",X"14",X"54",X"14",X"55",X"54",X"11",X"50",X"00",X"00",
		X"00",X"00",X"15",X"50",X"55",X"54",X"40",X"04",X"40",X"04",X"54",X"54",X"14",X"50",X"00",X"00",
		X"00",X"00",X"55",X"54",X"55",X"54",X"40",X"04",X"40",X"04",X"55",X"54",X"15",X"50",X"00",X"00",
		X"00",X"00",X"55",X"54",X"55",X"54",X"41",X"04",X"41",X"04",X"40",X"04",X"50",X"14",X"00",X"00",
		X"00",X"00",X"55",X"54",X"55",X"54",X"41",X"00",X"41",X"00",X"40",X"00",X"50",X"00",X"00",X"00",
		X"00",X"00",X"15",X"50",X"55",X"54",X"40",X"04",X"41",X"04",X"51",X"54",X"11",X"50",X"00",X"00",
		X"00",X"00",X"55",X"54",X"55",X"54",X"01",X"00",X"01",X"00",X"55",X"54",X"55",X"54",X"00",X"00",
		X"00",X"00",X"40",X"04",X"40",X"04",X"55",X"54",X"55",X"54",X"40",X"04",X"40",X"04",X"00",X"00",
		X"00",X"00",X"00",X"50",X"40",X"54",X"40",X"04",X"55",X"54",X"55",X"50",X"40",X"00",X"00",X"00",
		X"00",X"00",X"55",X"54",X"55",X"54",X"05",X"40",X"14",X"50",X"50",X"14",X"40",X"04",X"00",X"00",
		X"00",X"00",X"55",X"54",X"55",X"54",X"00",X"04",X"00",X"04",X"00",X"14",X"00",X"14",X"00",X"00",
		X"00",X"00",X"55",X"54",X"55",X"54",X"40",X"00",X"55",X"54",X"40",X"00",X"15",X"54",X"00",X"00",
		X"00",X"00",X"55",X"54",X"55",X"54",X"15",X"00",X"01",X"50",X"55",X"54",X"55",X"54",X"00",X"00",
		X"00",X"00",X"15",X"50",X"55",X"54",X"40",X"04",X"40",X"04",X"55",X"54",X"15",X"50",X"00",X"00",
		X"00",X"00",X"55",X"54",X"55",X"54",X"41",X"00",X"41",X"00",X"55",X"00",X"14",X"00",X"00",X"00",
		X"00",X"00",X"15",X"50",X"55",X"54",X"40",X"04",X"40",X"44",X"55",X"50",X"15",X"44",X"00",X"00",
		X"00",X"00",X"55",X"54",X"55",X"54",X"41",X"00",X"41",X"40",X"54",X"54",X"10",X"04",X"00",X"00",
		X"00",X"00",X"14",X"10",X"55",X"14",X"41",X"04",X"41",X"04",X"51",X"54",X"10",X"50",X"00",X"00",
		X"00",X"00",X"54",X"00",X"40",X"00",X"55",X"54",X"55",X"54",X"40",X"00",X"54",X"00",X"00",X"00",
		X"00",X"00",X"55",X"50",X"55",X"54",X"00",X"04",X"00",X"04",X"55",X"54",X"55",X"50",X"00",X"00",
		X"00",X"00",X"54",X"00",X"15",X"50",X"00",X"14",X"01",X"54",X"55",X"40",X"40",X"00",X"00",X"00",
		X"00",X"00",X"55",X"50",X"55",X"54",X"00",X"04",X"15",X"50",X"00",X"04",X"55",X"50",X"00",X"00",
		X"00",X"00",X"40",X"04",X"54",X"54",X"15",X"50",X"05",X"40",X"54",X"54",X"40",X"04",X"00",X"00",
		X"00",X"00",X"50",X"00",X"54",X"00",X"05",X"54",X"01",X"54",X"55",X"00",X"50",X"00",X"00",X"00",
		X"00",X"00",X"50",X"14",X"40",X"54",X"41",X"44",X"45",X"04",X"54",X"04",X"50",X"14",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AF",X"FA",X"BF",X"FA",X"AA",X"BA",X"FF",X"FF",X"FF",X"FF",X"AA",X"BA",X"AA",X"AA",
		X"AE",X"AA",X"AF",X"FE",X"AE",X"AA",X"AA",X"AA",X"AF",X"FE",X"AA",X"EA",X"AA",X"EA",X"AF",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"50",X"01",X"10",X"01",X"50",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"2A",X"A0",X"AA",X"A8",X"80",X"08",X"80",X"08",X"AA",X"A8",X"2A",X"A0",X"00",X"00",
		X"00",X"00",X"00",X"08",X"20",X"08",X"AA",X"A8",X"AA",X"A8",X"00",X"08",X"00",X"08",X"00",X"00",
		X"00",X"00",X"20",X"A8",X"A2",X"A8",X"82",X"08",X"82",X"08",X"AA",X"28",X"28",X"28",X"00",X"00",
		X"00",X"00",X"A0",X"A0",X"80",X"A8",X"88",X"08",X"88",X"08",X"A2",X"A8",X"A0",X"A0",X"00",X"00",
		X"00",X"00",X"0A",X"80",X"2A",X"80",X"00",X"80",X"00",X"80",X"AA",X"A8",X"AA",X"A8",X"00",X"00",
		X"00",X"00",X"AA",X"20",X"AA",X"28",X"88",X"08",X"88",X"08",X"8A",X"A8",X"82",X"A0",X"00",X"00",
		X"00",X"00",X"2A",X"A0",X"AA",X"A8",X"82",X"08",X"82",X"08",X"A2",X"A8",X"20",X"A0",X"00",X"00",
		X"00",X"00",X"A0",X"00",X"A0",X"00",X"80",X"A8",X"82",X"A8",X"AA",X"00",X"A8",X"00",X"00",X"00",
		X"00",X"00",X"22",X"A0",X"AA",X"A8",X"8A",X"08",X"8A",X"08",X"AA",X"A8",X"22",X"A0",X"00",X"00",
		X"00",X"00",X"28",X"20",X"AA",X"28",X"82",X"08",X"82",X"08",X"AA",X"A8",X"2A",X"A0",X"00",X"00",
		X"00",X"00",X"AA",X"A8",X"AA",X"A8",X"A0",X"80",X"A0",X"80",X"AA",X"A8",X"2A",X"A8",X"00",X"00",
		X"00",X"00",X"AA",X"A8",X"AA",X"A8",X"82",X"08",X"82",X"08",X"AA",X"A8",X"28",X"A0",X"00",X"00",
		X"00",X"00",X"2A",X"A0",X"AA",X"A8",X"80",X"08",X"80",X"08",X"A8",X"A8",X"28",X"A0",X"00",X"00",
		X"00",X"00",X"AA",X"A8",X"AA",X"A8",X"80",X"08",X"A0",X"28",X"AA",X"A8",X"2A",X"A0",X"00",X"00",
		X"00",X"00",X"AA",X"A8",X"AA",X"A8",X"82",X"08",X"82",X"08",X"80",X"08",X"A0",X"28",X"00",X"00",
		X"00",X"00",X"AA",X"A8",X"AA",X"A8",X"82",X"00",X"82",X"00",X"80",X"00",X"A0",X"00",X"00",X"00",
		X"00",X"00",X"2A",X"A0",X"AA",X"A8",X"80",X"08",X"82",X"08",X"A2",X"A8",X"22",X"A0",X"00",X"00",
		X"00",X"00",X"AA",X"A8",X"AA",X"A8",X"02",X"00",X"02",X"00",X"AA",X"A8",X"AA",X"A8",X"00",X"00",
		X"00",X"00",X"80",X"08",X"80",X"08",X"AA",X"A8",X"AA",X"A8",X"80",X"08",X"80",X"08",X"00",X"00",
		X"00",X"00",X"00",X"A0",X"80",X"A8",X"80",X"08",X"AA",X"A8",X"AA",X"A0",X"80",X"00",X"00",X"00",
		X"00",X"00",X"AA",X"A8",X"AA",X"A8",X"0A",X"80",X"28",X"A0",X"A0",X"28",X"80",X"08",X"00",X"00",
		X"00",X"00",X"AA",X"A8",X"AA",X"A8",X"00",X"08",X"00",X"08",X"00",X"28",X"00",X"28",X"00",X"00",
		X"00",X"00",X"AA",X"A8",X"AA",X"A8",X"80",X"00",X"AA",X"A8",X"80",X"00",X"2A",X"A8",X"00",X"00",
		X"00",X"00",X"AA",X"A8",X"AA",X"A8",X"2A",X"00",X"02",X"A0",X"AA",X"A8",X"AA",X"A8",X"00",X"00",
		X"00",X"00",X"2A",X"A0",X"AA",X"A8",X"80",X"08",X"80",X"08",X"AA",X"A8",X"2A",X"A0",X"00",X"00",
		X"00",X"00",X"AA",X"A8",X"AA",X"A8",X"82",X"00",X"82",X"00",X"AA",X"00",X"28",X"00",X"00",X"00",
		X"00",X"00",X"2A",X"A0",X"AA",X"A8",X"80",X"08",X"80",X"88",X"AA",X"A0",X"2A",X"88",X"00",X"00",
		X"00",X"00",X"AA",X"A8",X"AA",X"A8",X"82",X"00",X"82",X"80",X"A8",X"A8",X"20",X"08",X"00",X"00",
		X"00",X"00",X"28",X"20",X"AA",X"28",X"82",X"08",X"82",X"08",X"A2",X"A8",X"20",X"A0",X"00",X"00",
		X"00",X"00",X"A8",X"00",X"80",X"00",X"AA",X"A8",X"AA",X"A8",X"80",X"00",X"A8",X"00",X"00",X"00",
		X"00",X"00",X"AA",X"A0",X"AA",X"A8",X"00",X"08",X"00",X"08",X"AA",X"A8",X"AA",X"A0",X"00",X"00",
		X"00",X"00",X"A8",X"00",X"AA",X"A0",X"00",X"28",X"02",X"A8",X"AA",X"80",X"A0",X"00",X"00",X"00",
		X"00",X"00",X"AA",X"A0",X"AA",X"A8",X"00",X"08",X"2A",X"A0",X"00",X"08",X"AA",X"A0",X"00",X"00",
		X"00",X"00",X"80",X"08",X"A8",X"A8",X"2A",X"A0",X"0A",X"80",X"A8",X"A8",X"80",X"08",X"00",X"00",
		X"00",X"00",X"A0",X"00",X"A8",X"00",X"0A",X"A8",X"02",X"A8",X"AA",X"00",X"A0",X"00",X"00",X"00",
		X"00",X"00",X"A0",X"28",X"80",X"A8",X"82",X"88",X"8A",X"08",X"A8",X"08",X"A0",X"28",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"C0",X"0F",X"F0",X"2F",X"F8",X"EF",X"FB",X"FE",X"BF",X"3A",X"AC",X"0A",X"A0",X"03",X"80",
		X"0A",X"A0",X"0A",X"AC",X"28",X"2B",X"A0",X"2A",X"A0",X"2A",X"28",X"2B",X"0A",X"AC",X"0A",X"A0",
		X"0F",X"F0",X"3F",X"FC",X"FE",X"BF",X"FA",X"AF",X"FA",X"AF",X"FE",X"BF",X"3F",X"FC",X"0F",X"F0",
		X"09",X"E0",X"25",X"D8",X"96",X"D6",X"5B",X"FF",X"FF",X"E5",X"97",X"96",X"27",X"58",X"0B",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"0C",X"00",X"0C",X"00",X"0C",X"FF",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"E0",X"00",X"E0",X"00",X"E0",X"00",X"E0",X"00",
		X"30",X"00",X"30",X"00",X"30",X"00",X"3F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"FF",X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FC",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",
		X"C0",X"00",X"C0",X"00",X"C0",X"00",X"FF",X"FF",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",
		X"C0",X"00",X"C0",X"00",X"C0",X"00",X"FF",X"FF",X"C0",X"08",X"C0",X"08",X"C0",X"08",X"C0",X"08",
		X"00",X"0C",X"00",X"0C",X"00",X"0C",X"FF",X"FC",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",
		X"30",X"00",X"30",X"00",X"30",X"00",X"3F",X"FF",X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00",
		X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00",
		X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",
		X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",
		X"05",X"50",X"15",X"00",X"75",X"40",X"5D",X"55",X"5D",X"55",X"75",X"40",X"15",X"00",X"05",X"50",
		X"00",X"00",X"05",X"05",X"51",X"05",X"15",X"50",X"15",X"50",X"51",X"05",X"05",X"05",X"00",X"00",
		X"55",X"50",X"05",X"45",X"1F",X"54",X"73",X"D5",X"73",X"D5",X"1F",X"54",X"05",X"45",X"55",X"50",
		X"51",X"14",X"44",X"05",X"51",X"14",X"15",X"50",X"15",X"50",X"51",X"14",X"44",X"05",X"51",X"14",
		X"EA",X"AA",X"A5",X"5A",X"95",X"D6",X"9F",X"D6",X"97",X"F6",X"97",X"56",X"A5",X"5A",X"AA",X"AB",
		X"EA",X"AA",X"AA",X"AA",X"AD",X"FA",X"AF",X"DA",X"A7",X"FA",X"AF",X"7A",X"AA",X"AA",X"AA",X"AB",
		X"00",X"00",X"00",X"00",X"3D",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"00",X"10",X"00",X"10",X"00",X"10",X"00",X"30",X"00",X"30",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3D",X"54",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E8",X"2B",X"B8",X"2E",X"A0",X"0A",X"03",X"C0",X"03",X"C0",X"A0",X"0A",X"B8",X"2E",X"E8",X"2B",
		X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"03",X"00",X"03",X"00",X"00",X"00",
		X"AA",X"EA",X"AB",X"EA",X"A7",X"EA",X"A9",X"6A",X"A6",X"FA",X"A6",X"FA",X"AB",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3D",X"54",X"00",X"00",
		X"00",X"00",X"10",X"00",X"10",X"00",X"10",X"00",X"10",X"00",X"30",X"00",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"33",X"FF",X"FF",X"3F",X"FC",X"BF",X"FE",X"EF",X"FB",X"2F",X"F8",X"EB",X"EB",X"EC",X"3B",
		X"EC",X"3B",X"EB",X"EB",X"2F",X"F8",X"EF",X"FB",X"BF",X"FE",X"3F",X"FC",X"FF",X"FF",X"CC",X"33",
		X"03",X"CA",X"83",X"D6",X"A3",X"CA",X"E0",X"0B",X"FC",X"3F",X"EE",X"BB",X"AA",X"BA",X"AA",X"AA",
		X"AA",X"AA",X"AE",X"AA",X"EE",X"BB",X"FC",X"3F",X"E0",X"0B",X"A3",X"CA",X"97",X"C2",X"A3",X"C0",
		X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"3F",X"F0",
		X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"3F",X"F0",
		X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"3F",X"F0",
		X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"3F",X"F0",
		X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"3F",X"F0",
		X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"3F",X"F0",
		X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"3F",X"F0",
		X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"3F",X"F0",
		X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"3F",X"F0",
		X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"3F",X"F0",
		X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"3F",X"F0",
		X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"3F",X"F0",
		X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"3F",X"F0",
		X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"3F",X"F0",
		X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"3F",X"F0",
		X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"3F",X"F0",
		X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"3F",X"F0",
		X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"3F",X"F0",
		X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"00",X"00",
		X"3D",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"03",X"00",X"03",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",
		X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"AA",X"AA",X"02",X"00",X"02",X"00",X"02",X"00",
		X"00",X"00",X"2A",X"A8",X"2A",X"A8",X"20",X"80",X"20",X"A0",X"2A",X"28",X"08",X"08",X"00",X"00",
		X"00",X"00",X"2A",X"A8",X"2A",X"A8",X"20",X"80",X"20",X"80",X"2A",X"A8",X"0A",X"A8",X"00",X"00",
		X"00",X"00",X"0A",X"A0",X"2A",X"A8",X"20",X"08",X"20",X"08",X"28",X"28",X"08",X"20",X"00",X"00",
		X"00",X"00",X"2A",X"A8",X"2A",X"A8",X"02",X"00",X"02",X"80",X"08",X"A8",X"20",X"28",X"00",X"00",
		X"28",X"00",X"82",X"00",X"2A",X"80",X"2A",X"A2",X"2A",X"AA",X"2A",X"A2",X"82",X"80",X"2A",X"00",
		X"94",X"B9",X"16",X"10",X"96",X"9F",X"24",X"D8",X"84",X"FF",X"67",X"89",X"86",X"09",X"37",X"0C",
		X"95",X"BB",X"36",X"B1",X"9E",X"85",X"35",X"DD",X"D7",X"9E",X"86",X"99",X"DE",X"4F",X"D3",X"9B",
		X"35",X"D4",X"A1",X"B3",X"B6",X"8D",X"D6",X"9C",X"73",X"A7",X"8E",X"8F",X"00",X"D5",X"FD",X"89",
		X"77",X"3A",X"CE",X"99",X"FF",X"DF",X"3D",X"99",X"B7",X"BD",X"BB",X"99",X"5C",X"89",X"CA",X"8D",
		X"00",X"CE",X"5F",X"98",X"AF",X"94",X"96",X"9D",X"0F",X"9C",X"7D",X"D8",X"9E",X"8D",X"14",X"9B",
		X"16",X"75",X"17",X"B1",X"E6",X"FD",X"92",X"90",X"86",X"D5",X"77",X"DC",X"3E",X"85",X"83",X"89",
		X"76",X"EC",X"C7",X"98",X"C6",X"3C",X"86",X"89",X"B5",X"FC",X"13",X"BC",X"92",X"C1",X"C4",X"B9",
		X"A6",X"9F",X"17",X"08",X"DE",X"C9",X"02",X"AD",X"37",X"00",X"57",X"98",X"FE",X"F5",X"04",X"8A",
		X"46",X"63",X"E6",X"BC",X"66",X"EB",X"F6",X"31",X"66",X"23",X"2B",X"22",X"2E",X"7D",X"E3",X"CD",
		X"64",X"40",X"E2",X"3E",X"36",X"0D",X"60",X"73",X"E6",X"2B",X"64",X"42",X"EE",X"7F",X"46",X"D9",
		X"44",X"EC",X"64",X"17",X"6F",X"7B",X"C4",X"E3",X"6C",X"2B",X"62",X"36",X"62",X"D4",X"E3",X"FF",
		X"0E",X"54",X"6E",X"1C",X"6E",X"6F",X"ED",X"23",X"40",X"62",X"37",X"68",X"CE",X"2E",X"F6",X"28",
		X"E6",X"D2",X"27",X"FA",X"12",X"5B",X"0E",X"B1",X"46",X"46",X"46",X"EC",X"AC",X"83",X"EA",X"D3",
		X"E6",X"44",X"77",X"D0",X"6A",X"DB",X"2C",X"F3",X"64",X"D8",X"E3",X"08",X"EE",X"7E",X"7B",X"F3",
		X"26",X"73",X"32",X"CE",X"26",X"1F",X"F4",X"EB",X"8C",X"0E",X"E6",X"8A",X"E2",X"79",X"C3",X"79",
		X"EE",X"2A",X"47",X"A8",X"32",X"4C",X"06",X"EC",X"66",X"2E",X"66",X"48",X"0E",X"03",X"E6",X"F3",
		X"44",X"CF",X"54",X"33",X"66",X"3D",X"48",X"FC",X"EE",X"63",X"46",X"F1",X"E4",X"8F",X"C2",X"F5",
		X"E6",X"E4",X"4C",X"A0",X"A6",X"EB",X"2A",X"0F",X"36",X"6E",X"66",X"10",X"FF",X"63",X"42",X"BB",
		X"A6",X"70",X"00",X"09",X"4A",X"5F",X"78",X"79",X"CE",X"83",X"75",X"F4",X"63",X"41",X"4E",X"0F",
		X"34",X"DE",X"26",X"1B",X"36",X"C8",X"C4",X"33",X"64",X"20",X"6E",X"F2",X"3E",X"CB",X"4C",X"30",
		X"44",X"0C",X"72",X"A8",X"66",X"49",X"72",X"37",X"2E",X"F4",X"47",X"3C",X"EE",X"F1",X"30",X"0F",
		X"6E",X"03",X"76",X"3A",X"34",X"6F",X"0F",X"ED",X"68",X"F2",X"66",X"A0",X"46",X"B5",X"76",X"B2",
		X"46",X"06",X"67",X"39",X"23",X"04",X"5A",X"FF",X"C6",X"2D",X"64",X"08",X"E7",X"03",X"EE",X"1B",
		X"66",X"82",X"03",X"CC",X"67",X"51",X"F4",X"0C",X"66",X"C6",X"E2",X"28",X"EE",X"C3",X"60",X"49");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
