`define BUILD_DATE "181125"
`define BUILD_TIME "152519"
