library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ttag_bg_bits_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ttag_bg_bits_1 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"50",X"15",X"01",X"50",X"15",X"01",X"50",X"15",X"50",X"54",X"05",X"40",X"54",X"05",X"40",X"54",
		X"51",X"50",X"15",X"01",X"50",X"15",X"01",X"50",X"55",X"40",X"54",X"05",X"40",X"54",X"05",X"40",
		X"55",X"01",X"50",X"15",X"01",X"50",X"15",X"00",X"54",X"05",X"40",X"54",X"05",X"40",X"54",X"00",
		X"50",X"15",X"01",X"50",X"15",X"01",X"50",X"00",X"50",X"54",X"05",X"40",X"54",X"05",X"40",X"00",
		X"51",X"50",X"15",X"01",X"50",X"15",X"00",X"00",X"55",X"40",X"54",X"05",X"40",X"54",X"00",X"00",
		X"55",X"01",X"50",X"15",X"01",X"50",X"00",X"00",X"54",X"05",X"40",X"54",X"05",X"40",X"00",X"00",
		X"50",X"15",X"01",X"50",X"15",X"00",X"00",X"00",X"50",X"54",X"05",X"40",X"54",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"01",X"55",X"01",X"50",X"15",X"01",X"50",X"15",X"01",X"54",X"05",X"40",X"54",X"05",X"40",X"54",
		X"00",X"54",X"15",X"01",X"50",X"15",X"01",X"50",X"00",X"14",X"54",X"05",X"40",X"54",X"05",X"40",
		X"00",X"15",X"50",X"15",X"01",X"50",X"15",X"00",X"00",X"05",X"40",X"54",X"05",X"40",X"54",X"00",
		X"00",X"01",X"41",X"50",X"15",X"01",X"50",X"00",X"00",X"01",X"55",X"40",X"54",X"05",X"40",X"00",
		X"00",X"00",X"55",X"01",X"50",X"15",X"00",X"00",X"00",X"00",X"14",X"05",X"40",X"54",X"00",X"00",
		X"00",X"00",X"15",X"15",X"01",X"50",X"00",X"00",X"00",X"00",X"05",X"54",X"05",X"40",X"00",X"00",
		X"00",X"00",X"01",X"50",X"15",X"00",X"00",X"00",X"00",X"00",X"01",X"50",X"54",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"55",X"40",X"54",X"05",X"40",X"54",X"05",X"00",X"55",X"01",X"50",X"15",X"01",X"50",X"15",
		X"00",X"15",X"05",X"40",X"54",X"05",X"40",X"55",X"00",X"05",X"15",X"01",X"50",X"15",X"01",X"55",
		X"00",X"05",X"54",X"05",X"40",X"54",X"05",X"45",X"00",X"01",X"50",X"15",X"01",X"50",X"15",X"05",
		X"00",X"00",X"50",X"54",X"05",X"40",X"54",X"05",X"00",X"00",X"55",X"50",X"15",X"01",X"50",X"15",
		X"00",X"00",X"15",X"40",X"54",X"05",X"40",X"55",X"00",X"00",X"05",X"01",X"50",X"15",X"01",X"55",
		X"00",X"00",X"05",X"45",X"40",X"54",X"05",X"45",X"00",X"00",X"01",X"55",X"01",X"50",X"15",X"05",
		X"00",X"00",X"00",X"54",X"05",X"40",X"54",X"05",X"00",X"00",X"00",X"54",X"15",X"01",X"50",X"15",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"41",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"50",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"6A",X"AA",X"75",X"D7",X"5D",X"75",X"AA",X"A9",X"6A",X"82",X"5D",X"75",X"D7",X"5D",X"AA",X"09",
		X"6A",X"AA",X"57",X"5D",X"75",X"D5",X"AA",X"09",X"6A",X"82",X"75",X"D7",X"5D",X"75",X"AA",X"09",
		X"6A",X"82",X"5D",X"75",X"D7",X"5D",X"AA",X"A9",X"6A",X"82",X"55",X"55",X"55",X"55",X"AA",X"A9",
		X"AA",X"AA",X"55",X"55",X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"55",X"55",X"55",X"55",X"AA",X"AA",
		X"AA",X"AA",X"55",X"55",X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"55",X"55",X"55",X"55",X"AA",X"AA",
		X"A0",X"2A",X"55",X"55",X"55",X"55",X"AA",X"0A",X"A0",X"0A",X"55",X"55",X"55",X"55",X"A8",X"0A",
		X"AA",X"AA",X"55",X"55",X"55",X"55",X"AA",X"AA",X"AA",X"02",X"55",X"55",X"55",X"55",X"AA",X"80",
		X"AA",X"02",X"55",X"55",X"55",X"55",X"AA",X"80",X"AA",X"AA",X"55",X"55",X"55",X"55",X"AA",X"AA",
		X"51",X"50",X"15",X"01",X"50",X"00",X"00",X"00",X"55",X"40",X"54",X"05",X"40",X"00",X"00",X"00",
		X"55",X"01",X"50",X"15",X"00",X"00",X"00",X"00",X"54",X"05",X"40",X"54",X"00",X"00",X"00",X"00",
		X"50",X"15",X"01",X"50",X"00",X"00",X"00",X"00",X"50",X"54",X"05",X"40",X"00",X"00",X"00",X"00",
		X"51",X"50",X"15",X"00",X"00",X"00",X"00",X"00",X"55",X"40",X"54",X"00",X"00",X"00",X"00",X"00",
		X"55",X"01",X"50",X"00",X"00",X"00",X"00",X"00",X"54",X"05",X"40",X"00",X"00",X"00",X"00",X"00",
		X"50",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"54",X"00",X"00",X"00",X"00",X"00",X"00",
		X"51",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"55",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"15",X"54",X"05",X"40",X"55",X"00",X"00",X"00",X"05",X"50",X"15",X"01",X"55",
		X"00",X"00",X"00",X"05",X"40",X"54",X"05",X"45",X"00",X"00",X"00",X"15",X"01",X"50",X"15",X"05",
		X"00",X"00",X"00",X"54",X"05",X"40",X"54",X"05",X"00",X"00",X"01",X"50",X"15",X"01",X"50",X"15",
		X"00",X"00",X"05",X"40",X"54",X"05",X"40",X"55",X"00",X"00",X"15",X"01",X"50",X"15",X"01",X"55",
		X"00",X"00",X"54",X"05",X"40",X"54",X"05",X"45",X"00",X"01",X"50",X"15",X"01",X"50",X"15",X"05",
		X"00",X"05",X"40",X"54",X"05",X"40",X"54",X"05",X"00",X"15",X"01",X"50",X"15",X"01",X"50",X"15",
		X"00",X"54",X"05",X"40",X"54",X"05",X"40",X"55",X"01",X"50",X"15",X"01",X"50",X"15",X"01",X"55",
		X"05",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"A8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"95",X"58",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"A8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"95",X"58",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"A8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"95",X"58",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"A8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"95",X"58",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"A8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"95",X"58",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"A8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"95",X"58",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"A8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"57",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"75",X"55",X"55",X"55",X"55",
		X"55",X"55",X"57",X"5D",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"D7",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"75",X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"5D",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"D7",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"75",X"55",X"55",X"55",X"55",
		X"55",X"55",X"57",X"5D",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"D7",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"75",X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"5D",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"D7",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"75",X"55",X"55",X"55",X"55",
		X"55",X"55",X"57",X"5D",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"D7",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"54",X"50",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"40",X"00",X"00",X"00",X"00",X"00",
		X"01",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"50",X"00",X"00",X"00",X"00",X"00",
		X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"01",X"50",X"15",X"01",X"50",X"15",X"00",X"55",X"40",X"54",X"05",X"40",X"54",X"14",X"00",
		X"51",X"50",X"15",X"01",X"50",X"15",X"54",X"00",X"50",X"54",X"05",X"40",X"54",X"05",X"50",X"00",
		X"50",X"15",X"01",X"50",X"15",X"01",X"40",X"00",X"54",X"05",X"40",X"54",X"05",X"45",X"40",X"00",
		X"55",X"01",X"50",X"15",X"01",X"55",X"00",X"00",X"55",X"40",X"54",X"05",X"40",X"54",X"00",X"00",
		X"51",X"50",X"15",X"01",X"50",X"54",X"00",X"00",X"50",X"54",X"05",X"40",X"55",X"50",X"00",X"00",
		X"50",X"15",X"01",X"50",X"15",X"40",X"00",X"00",X"54",X"05",X"40",X"54",X"05",X"40",X"00",X"00",
		X"55",X"01",X"50",X"15",X"15",X"00",X"00",X"00",X"55",X"40",X"54",X"05",X"54",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"54",X"05",X"40",X"54",X"05",X"40",X"15",X"00",X"15",X"01",X"50",X"15",X"01",X"50",X"14",X"00",
		X"05",X"40",X"54",X"05",X"40",X"54",X"54",X"00",X"01",X"50",X"15",X"01",X"50",X"15",X"50",X"00",
		X"00",X"54",X"05",X"40",X"54",X"05",X"40",X"00",X"00",X"15",X"01",X"50",X"15",X"15",X"40",X"00",
		X"00",X"05",X"40",X"54",X"05",X"55",X"00",X"00",X"00",X"01",X"50",X"15",X"01",X"54",X"00",X"00",
		X"00",X"00",X"54",X"05",X"40",X"54",X"00",X"00",X"00",X"00",X"15",X"01",X"51",X"50",X"00",X"00",
		X"00",X"00",X"05",X"40",X"55",X"40",X"00",X"00",X"00",X"00",X"01",X"50",X"15",X"40",X"00",X"00",
		X"00",X"00",X"00",X"54",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"14",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"54",X"05",X"40",X"54",X"05",X"40",X"54",X"05",X"15",X"01",X"50",X"15",X"01",X"50",X"15",X"05",
		X"05",X"40",X"54",X"05",X"40",X"54",X"05",X"45",X"01",X"50",X"15",X"01",X"50",X"15",X"01",X"55",
		X"00",X"54",X"05",X"40",X"54",X"05",X"40",X"55",X"00",X"15",X"01",X"50",X"15",X"01",X"50",X"15",
		X"00",X"05",X"40",X"54",X"05",X"40",X"54",X"05",X"00",X"01",X"50",X"15",X"01",X"50",X"15",X"05",
		X"00",X"00",X"54",X"05",X"40",X"54",X"05",X"45",X"00",X"00",X"15",X"01",X"50",X"15",X"01",X"55",
		X"00",X"00",X"05",X"40",X"54",X"05",X"40",X"55",X"00",X"00",X"01",X"50",X"15",X"01",X"50",X"15",
		X"00",X"00",X"00",X"54",X"05",X"40",X"54",X"05",X"00",X"00",X"00",X"15",X"01",X"50",X"15",X"05",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"AA",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0A",X"66",X"80",X"00",X"00",X"00",X"00",X"00",X"2A",X"AA",X"A0",X"00",X"00",
		X"00",X"00",X"00",X"26",X"66",X"60",X"00",X"00",X"00",X"00",X"00",X"2A",X"AA",X"A0",X"00",X"00",
		X"00",X"00",X"00",X"26",X"66",X"60",X"00",X"00",X"00",X"00",X"00",X"2A",X"AA",X"A0",X"00",X"00",
		X"00",X"00",X"00",X"26",X"66",X"60",X"00",X"00",X"00",X"00",X"00",X"2A",X"AA",X"A0",X"00",X"00",
		X"00",X"00",X"00",X"0A",X"66",X"80",X"00",X"00",X"00",X"00",X"00",X"02",X"AA",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"51",X"50",X"15",X"01",X"54",X"00",X"00",X"00",X"50",X"54",X"05",X"40",X"54",X"00",X"00",X"00",
		X"50",X"15",X"01",X"50",X"15",X"00",X"00",X"00",X"54",X"05",X"40",X"54",X"05",X"40",X"00",X"00",
		X"55",X"01",X"50",X"15",X"01",X"50",X"00",X"00",X"55",X"40",X"54",X"05",X"40",X"54",X"00",X"00",
		X"51",X"50",X"15",X"01",X"50",X"15",X"00",X"00",X"50",X"54",X"05",X"40",X"54",X"05",X"40",X"00",
		X"50",X"15",X"01",X"50",X"15",X"01",X"50",X"00",X"54",X"05",X"40",X"54",X"05",X"40",X"54",X"00",
		X"55",X"01",X"50",X"15",X"01",X"50",X"15",X"00",X"55",X"40",X"54",X"05",X"40",X"54",X"05",X"40",
		X"51",X"50",X"15",X"01",X"50",X"15",X"01",X"50",X"50",X"54",X"05",X"40",X"54",X"05",X"40",X"54",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"05",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"50",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"05",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"50",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"05",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"50",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"50",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"15",
		X"00",X"00",X"00",X"05",X"40",X"54",X"05",X"45",X"00",X"00",X"00",X"01",X"50",X"15",X"01",X"55",
		X"00",X"00",X"00",X"00",X"54",X"05",X"40",X"55",X"00",X"00",X"00",X"00",X"15",X"01",X"50",X"15",
		X"00",X"00",X"00",X"00",X"05",X"40",X"54",X"05",X"00",X"00",X"00",X"00",X"01",X"50",X"15",X"05",
		X"00",X"00",X"00",X"00",X"00",X"54",X"05",X"45",X"00",X"00",X"00",X"00",X"00",X"15",X"01",X"55",
		X"00",X"00",X"00",X"00",X"00",X"05",X"40",X"55",X"00",X"00",X"00",X"00",X"00",X"01",X"50",X"15",
		X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"45",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"15",
		X"AA",X"AA",X"A5",X"44",X"44",X"44",X"44",X"44",X"AA",X"AA",X"A5",X"55",X"11",X"11",X"11",X"11",
		X"82",X"AA",X"A4",X"44",X"44",X"44",X"44",X"44",X"82",X"AA",X"A5",X"11",X"15",X"11",X"11",X"15",
		X"82",X"AA",X"A5",X"54",X"45",X"45",X"44",X"55",X"82",X"AA",X"A5",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"80",X"2A",X"A0",X"2A",X"AA",X"A0",X"2A",X"AA",
		X"80",X"2A",X"A0",X"2A",X"AA",X"A0",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"02",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"02",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"2A",X"AA",X"AA",X"AA",X"A0",X"2A",
		X"AA",X"A0",X"2A",X"AA",X"AA",X"AA",X"A0",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"40",X"00",X"00",X"00",X"0F",X"00",X"04",X"11",X"10",X"00",X"00",X"03",X"FA",
		X"00",X"04",X"44",X"10",X"00",X"00",X"FE",X"AA",X"00",X"04",X"55",X"10",X"00",X"3F",X"AA",X"AA",
		X"00",X"01",X"00",X"40",X"0F",X"EA",X"AA",X"AA",X"00",X"00",X"55",X"03",X"FA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"FE",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"3F",X"AA",X"AA",X"AA",X"AA",X"BF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"AC",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"AB",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"0E",X"AB",X"0F",X"C0",X"00",X"00",X"03",X"FB",X"0E",X"AB",X"0E",X"BF",X"00",
		X"00",X"FE",X"AB",X"0E",X"AB",X"0E",X"AB",X"00",X"3F",X"AA",X"AB",X"0E",X"AB",X"0E",X"AB",X"00",
		X"EA",X"AA",X"AB",X"0E",X"AB",X"0E",X"AB",X"00",X"AA",X"AA",X"AB",X"0E",X"AB",X"0E",X"AB",X"00",
		X"AA",X"AA",X"AB",X"0E",X"AB",X"0E",X"AB",X"00",X"AA",X"AA",X"AB",X"0E",X"AB",X"0E",X"AB",X"00",
		X"AA",X"AA",X"AB",X"0E",X"AB",X"0E",X"AB",X"00",X"AB",X"FA",X"AB",X"0E",X"AB",X"0E",X"AB",X"00",
		X"FC",X"0E",X"AB",X"0E",X"AB",X"0E",X"AB",X"00",X"00",X"0E",X"AB",X"0E",X"AB",X"0E",X"AB",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EB",X"F0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"EA",X"AF",X"C0",X"00",X"00",X"00",X"00",X"00",X"EA",X"AA",X"BF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"2A",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"25",X"56",X"00",X"00",X"00",X"00",X"00",X"00",
		X"25",X"56",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",
		X"25",X"56",X"00",X"00",X"00",X"00",X"00",X"00",X"25",X"56",X"00",X"00",X"00",X"00",X"00",X"00",
		X"2A",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"25",X"56",X"00",X"00",X"00",X"00",X"00",X"00",
		X"25",X"56",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",
		X"25",X"56",X"00",X"00",X"00",X"00",X"00",X"00",X"25",X"56",X"00",X"00",X"00",X"00",X"00",X"00",
		X"2A",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"A8",X"0A",X"80",X"A8",X"0A",X"80",X"A8",X"0A",X"2A",X"02",X"A0",X"2A",X"02",X"A0",X"2A",X"0A",
		X"0A",X"80",X"A8",X"0A",X"80",X"A8",X"0A",X"8A",X"02",X"A0",X"2A",X"02",X"A0",X"2A",X"02",X"AA",
		X"00",X"A8",X"0A",X"80",X"A8",X"0A",X"80",X"AA",X"00",X"2A",X"02",X"A0",X"2A",X"02",X"A0",X"2A",
		X"00",X"0A",X"80",X"A8",X"0A",X"80",X"A8",X"0A",X"00",X"02",X"A0",X"2A",X"02",X"A0",X"2A",X"0A",
		X"00",X"00",X"A8",X"0A",X"80",X"A8",X"0A",X"8A",X"00",X"00",X"2A",X"02",X"A0",X"2A",X"02",X"AA",
		X"00",X"00",X"0A",X"80",X"A8",X"0A",X"80",X"AA",X"00",X"00",X"02",X"A0",X"2A",X"02",X"A0",X"2A",
		X"00",X"00",X"00",X"A8",X"0A",X"80",X"A8",X"0A",X"00",X"00",X"00",X"2A",X"02",X"A0",X"2A",X"0A",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"A0",X"2A",X"02",X"A0",X"2A",X"02",X"A0",X"2A",X"A0",X"A8",X"0A",X"80",X"A8",X"0A",X"80",X"A8",
		X"A2",X"A0",X"2A",X"02",X"A0",X"2A",X"02",X"A0",X"AA",X"80",X"A8",X"0A",X"80",X"A8",X"0A",X"80",
		X"AA",X"02",X"A0",X"2A",X"02",X"A0",X"2A",X"00",X"A8",X"0A",X"80",X"A8",X"0A",X"80",X"A8",X"00",
		X"A0",X"2A",X"02",X"A0",X"2A",X"02",X"A0",X"00",X"A0",X"A8",X"0A",X"80",X"A8",X"0A",X"80",X"00",
		X"A2",X"A0",X"2A",X"02",X"A0",X"2A",X"00",X"00",X"AA",X"80",X"A8",X"0A",X"80",X"A8",X"00",X"00",
		X"AA",X"02",X"A0",X"2A",X"02",X"A0",X"00",X"00",X"A8",X"0A",X"80",X"A8",X"0A",X"80",X"00",X"00",
		X"A0",X"2A",X"02",X"A0",X"2A",X"00",X"00",X"00",X"A0",X"A8",X"0A",X"80",X"A8",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FC",X"0F",X"C0",X"FC",X"0F",X"C0",X"FC",X"0F",X"3F",X"03",X"F0",X"3F",X"03",X"F0",X"3F",X"0F",
		X"0F",X"C0",X"FC",X"0F",X"C0",X"FC",X"0F",X"CF",X"03",X"F0",X"3F",X"03",X"F0",X"3F",X"03",X"FF",
		X"00",X"FC",X"0F",X"C0",X"FC",X"0F",X"C0",X"FF",X"00",X"3F",X"03",X"F0",X"3F",X"03",X"F0",X"3F",
		X"00",X"0F",X"C0",X"FC",X"0F",X"C0",X"FC",X"0F",X"00",X"03",X"F0",X"3F",X"03",X"F0",X"3F",X"0F",
		X"00",X"00",X"FC",X"0F",X"C0",X"FC",X"0F",X"CF",X"00",X"00",X"3F",X"03",X"F0",X"3F",X"03",X"FF",
		X"00",X"00",X"0F",X"C0",X"FC",X"0F",X"C0",X"FF",X"00",X"00",X"03",X"F0",X"3F",X"03",X"F0",X"3F",
		X"00",X"00",X"00",X"FC",X"0F",X"C0",X"FC",X"0F",X"00",X"00",X"00",X"3F",X"03",X"F0",X"3F",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"3F",X"03",X"F0",X"3F",X"03",X"F0",X"3F",X"F0",X"FC",X"0F",X"C0",X"FC",X"0F",X"C0",X"FC",
		X"F3",X"F0",X"3F",X"03",X"F0",X"3F",X"03",X"F0",X"FF",X"C0",X"FC",X"0F",X"C0",X"FC",X"0F",X"C0",
		X"FF",X"03",X"F0",X"3F",X"03",X"F0",X"3F",X"00",X"FC",X"0F",X"C0",X"FC",X"0F",X"C0",X"FC",X"00",
		X"F0",X"3F",X"03",X"F0",X"3F",X"03",X"F0",X"00",X"F0",X"FC",X"0F",X"C0",X"FC",X"0F",X"C0",X"00",
		X"F3",X"F0",X"3F",X"03",X"F0",X"3F",X"00",X"00",X"FF",X"C0",X"FC",X"0F",X"C0",X"FC",X"00",X"00",
		X"FF",X"03",X"F0",X"3F",X"03",X"F0",X"00",X"00",X"FC",X"0F",X"C0",X"FC",X"0F",X"C0",X"00",X"00",
		X"F0",X"3F",X"03",X"F0",X"3F",X"00",X"00",X"00",X"F0",X"FC",X"0F",X"C0",X"FC",X"00",X"00",X"00",
		X"03",X"F0",X"EA",X"AA",X"AA",X"AA",X"AF",X"C0",X"FE",X"B0",X"EA",X"AA",X"AA",X"AB",X"F0",X"00",
		X"EA",X"B0",X"EA",X"AA",X"AA",X"FC",X"00",X"00",X"EA",X"B0",X"EA",X"AA",X"BF",X"00",X"00",X"00",
		X"EA",X"B0",X"EA",X"AF",X"C0",X"00",X"00",X"00",X"EA",X"B0",X"EA",X"B0",X"00",X"00",X"00",X"00",
		X"EA",X"B0",X"EA",X"B0",X"00",X"00",X"00",X"00",X"EA",X"B0",X"EA",X"B0",X"00",X"00",X"00",X"00",
		X"EA",X"B0",X"EA",X"B0",X"00",X"00",X"00",X"00",X"EA",X"B0",X"EA",X"B0",X"00",X"00",X"00",X"0F",
		X"EA",X"B0",X"EA",X"B0",X"00",X"00",X"0F",X"FA",X"EA",X"B0",X"EA",X"B0",X"00",X"0F",X"FA",X"AA",
		X"EA",X"B0",X"EA",X"B0",X"0F",X"FA",X"AA",X"AA",X"EA",X"B0",X"EA",X"AF",X"FA",X"AA",X"AA",X"AA",
		X"EA",X"B0",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"B0",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"0E",X"AB",X"0E",X"AB",X"0E",X"AB",X"00",X"00",X"0E",X"AB",X"0E",X"AB",X"0E",X"AB",X"00",
		X"00",X"0E",X"AB",X"0E",X"AB",X"0E",X"AB",X"00",X"00",X"0E",X"AB",X"0E",X"AB",X"0E",X"AB",X"00",
		X"00",X"0E",X"AB",X"0E",X"AB",X"0E",X"AB",X"00",X"00",X"0E",X"AB",X"0E",X"AB",X"0E",X"AB",X"00",
		X"00",X"0E",X"AB",X"0E",X"AB",X"0E",X"AB",X"00",X"00",X"0E",X"AB",X"0E",X"AB",X"0E",X"AB",X"00",
		X"0F",X"FA",X"AB",X"0E",X"AB",X"0E",X"AB",X"00",X"FA",X"AA",X"AB",X"0E",X"AB",X"0E",X"AB",X"00",
		X"AA",X"AA",X"AB",X"0E",X"AB",X"0E",X"AB",X"00",X"AA",X"AA",X"AB",X"0E",X"AB",X"0E",X"AB",X"00",
		X"AA",X"AA",X"AB",X"0E",X"AB",X"0E",X"AB",X"00",X"AA",X"AA",X"AF",X"0E",X"AB",X"0E",X"AB",X"00",
		X"AA",X"AF",X"F0",X"0E",X"AB",X"0E",X"AB",X"00",X"AF",X"F0",X"00",X"0E",X"AB",X"0E",X"AB",X"00",
		X"00",X"00",X"EA",X"AA",X"AA",X"FC",X"00",X"00",X"00",X"00",X"EA",X"AA",X"AA",X"AB",X"F0",X"00",
		X"00",X"00",X"EA",X"AA",X"AA",X"AA",X"B0",X"00",X"00",X"00",X"EA",X"AA",X"AA",X"AA",X"B0",X"00",
		X"00",X"00",X"EA",X"AF",X"EA",X"AA",X"B0",X"00",X"00",X"00",X"EA",X"B0",X"3E",X"AA",X"B0",X"00",
		X"00",X"00",X"EA",X"B0",X"03",X"AA",X"B0",X"00",X"00",X"00",X"EA",X"B0",X"03",X"AA",X"B0",X"00",
		X"00",X"00",X"EA",X"B0",X"03",X"AA",X"B0",X"00",X"00",X"00",X"EA",X"B0",X"03",X"AA",X"B0",X"00",
		X"00",X"00",X"EA",X"B0",X"03",X"AA",X"B0",X"00",X"00",X"00",X"EB",X"F0",X"03",X"AA",X"B0",X"00",
		X"00",X"00",X"FC",X"00",X"03",X"AA",X"B0",X"00",X"00",X"00",X"00",X"00",X"FE",X"AA",X"B0",X"00",
		X"00",X"00",X"00",X"FF",X"AA",X"AA",X"B0",X"00",X"00",X"00",X"FF",X"AA",X"AA",X"AA",X"B0",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"0A",X"80",X"A8",X"0A",X"8A",X"00",X"00",X"00",X"02",X"A0",X"2A",X"02",X"AA",
		X"00",X"00",X"00",X"00",X"A8",X"0A",X"80",X"AA",X"00",X"00",X"00",X"00",X"2A",X"02",X"A0",X"2A",
		X"00",X"00",X"00",X"00",X"0A",X"80",X"A8",X"0A",X"00",X"00",X"00",X"00",X"02",X"A0",X"2A",X"0A",
		X"00",X"00",X"00",X"00",X"00",X"A8",X"0A",X"8A",X"00",X"00",X"00",X"00",X"00",X"2A",X"02",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"80",X"AA",X"00",X"00",X"00",X"00",X"00",X"02",X"A0",X"2A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"A8",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",X"0A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"8A",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",
		X"A2",X"A0",X"2A",X"02",X"A0",X"00",X"00",X"00",X"AA",X"80",X"A8",X"0A",X"80",X"00",X"00",X"00",
		X"AA",X"02",X"A0",X"2A",X"00",X"00",X"00",X"00",X"A8",X"0A",X"80",X"A8",X"00",X"00",X"00",X"00",
		X"A0",X"2A",X"02",X"A0",X"00",X"00",X"00",X"00",X"A0",X"A8",X"0A",X"80",X"00",X"00",X"00",X"00",
		X"A2",X"A0",X"2A",X"00",X"00",X"00",X"00",X"00",X"AA",X"80",X"A8",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"02",X"A0",X"00",X"00",X"00",X"00",X"00",X"A8",X"0A",X"80",X"00",X"00",X"00",X"00",X"00",
		X"A0",X"2A",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"A8",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A2",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"C0",X"FC",X"0F",X"CF",X"00",X"00",X"00",X"03",X"F0",X"3F",X"03",X"FF",
		X"00",X"00",X"00",X"00",X"FC",X"0F",X"C0",X"FF",X"00",X"00",X"00",X"00",X"3F",X"03",X"F0",X"3F",
		X"00",X"00",X"00",X"00",X"0F",X"C0",X"FC",X"0F",X"00",X"00",X"00",X"00",X"03",X"F0",X"3F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"FC",X"0F",X"CF",X"00",X"00",X"00",X"00",X"00",X"3F",X"03",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"C0",X"FF",X"00",X"00",X"00",X"00",X"00",X"03",X"F0",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"CF",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"F3",X"F0",X"3F",X"03",X"F0",X"00",X"00",X"00",X"FF",X"C0",X"FC",X"0F",X"C0",X"00",X"00",X"00",
		X"FF",X"03",X"F0",X"3F",X"00",X"00",X"00",X"00",X"FC",X"0F",X"C0",X"FC",X"00",X"00",X"00",X"00",
		X"F0",X"3F",X"03",X"F0",X"00",X"00",X"00",X"00",X"F0",X"FC",X"0F",X"C0",X"00",X"00",X"00",X"00",
		X"F3",X"F0",X"3F",X"00",X"00",X"00",X"00",X"00",X"FF",X"C0",X"FC",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"03",X"F0",X"00",X"00",X"00",X"00",X"00",X"FC",X"0F",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F3",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EA",X"B0",X"EA",X"AA",X"AA",X"AA",X"AA",X"AF",X"EA",X"B0",X"EA",X"AA",X"AA",X"AA",X"AF",X"F0",
		X"EA",X"B0",X"EA",X"AA",X"AA",X"AF",X"F0",X"00",X"EA",X"B0",X"EA",X"AA",X"AF",X"F0",X"00",X"03",
		X"EA",X"B0",X"EA",X"AF",X"F0",X"00",X"00",X"0E",X"EA",X"B0",X"EF",X"F0",X"00",X"0F",X"C0",X"3A",
		X"EA",X"B0",X"F0",X"00",X"0F",X"FA",X"B0",X"EA",X"EA",X"B0",X"00",X"0F",X"FA",X"AA",X"AC",X"EA",
		X"EA",X"B0",X"0F",X"FA",X"AA",X"AA",X"AB",X"AA",X"EA",X"B0",X"FA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"EA",X"B0",X"EA",X"AA",X"AA",X"AA",X"AA",X"AB",X"EA",X"B0",X"EA",X"AA",X"AA",X"AA",X"AA",X"AC",
		X"EA",X"B0",X"EA",X"AA",X"AA",X"AF",X"AA",X"B0",X"EA",X"B0",X"EA",X"AA",X"AF",X"F0",X"EA",X"B0",
		X"EA",X"B0",X"EA",X"AF",X"F0",X"00",X"EA",X"B0",X"EA",X"B0",X"EA",X"B0",X"00",X"00",X"EA",X"B0",
		X"F0",X"00",X"0F",X"0E",X"AB",X"0E",X"AB",X"00",X"00",X"0F",X"FB",X"0E",X"AB",X"0E",X"AB",X"00",
		X"0F",X"FA",X"AB",X"0E",X"AB",X"0E",X"AA",X"FF",X"FA",X"AA",X"AB",X"0E",X"AB",X"0E",X"AA",X"AA",
		X"AA",X"AA",X"AB",X"0E",X"AB",X"0E",X"AA",X"AA",X"AA",X"AA",X"AB",X"0E",X"AB",X"0E",X"AA",X"AA",
		X"AA",X"AA",X"AB",X"0E",X"AB",X"0E",X"AA",X"AA",X"AA",X"AA",X"AB",X"0E",X"AB",X"0E",X"AA",X"AA",
		X"AA",X"AA",X"AB",X"0E",X"AB",X"0E",X"AA",X"AA",X"AB",X"FA",X"AB",X"0E",X"AB",X"0E",X"AA",X"FF",
		X"FC",X"0E",X"AB",X"0E",X"AB",X"0E",X"FF",X"00",X"00",X"0E",X"AB",X"0E",X"AB",X"0F",X"00",X"00",
		X"00",X"0E",X"AB",X"0E",X"AB",X"00",X"00",X"FF",X"00",X"0E",X"AB",X"0E",X"AB",X"00",X"FF",X"AA",
		X"00",X"0E",X"AB",X"0E",X"AB",X"0F",X"AA",X"AA",X"00",X"0E",X"AB",X"0E",X"AB",X"0E",X"AA",X"AA",
		X"00",X"FF",X"AA",X"AA",X"AA",X"AA",X"B0",X"00",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"B0",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"F0",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"FF",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"FF",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"FF",X"00",X"00",X"F0",X"00",
		X"AA",X"AA",X"FF",X"00",X"00",X"FF",X"B0",X"00",X"AA",X"FF",X"00",X"00",X"FF",X"AA",X"B0",X"00",
		X"FF",X"00",X"00",X"FF",X"AA",X"AA",X"B0",X"00",X"00",X"00",X"FF",X"AA",X"AA",X"AA",X"B0",X"00",
		X"00",X"FF",X"AA",X"AA",X"AA",X"AA",X"B0",X"00",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"B0",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"F0",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"FF",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"FF",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",
		X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"2A",X"00",X"00",X"00",X"00",X"00",X"02",X"AA",
		X"0A",X"80",X"00",X"00",X"00",X"00",X"0A",X"8A",X"02",X"A0",X"00",X"00",X"00",X"00",X"0A",X"AA",
		X"00",X"A8",X"00",X"00",X"00",X"00",X"2A",X"AA",X"00",X"2A",X"00",X"00",X"00",X"00",X"A8",X"2A",
		X"00",X"0A",X"80",X"00",X"00",X"00",X"A8",X"0A",X"00",X"02",X"A0",X"00",X"00",X"02",X"AA",X"0A",
		X"00",X"00",X"A8",X"00",X"00",X"0A",X"8A",X"8A",X"00",X"00",X"2A",X"00",X"00",X"0A",X"02",X"AA",
		X"00",X"00",X"0A",X"80",X"00",X"2A",X"80",X"AA",X"00",X"00",X"02",X"A0",X"00",X"AA",X"A0",X"2A",
		X"00",X"00",X"00",X"A8",X"00",X"A0",X"A8",X"0A",X"00",X"00",X"00",X"2A",X"02",X"A0",X"2A",X"0A",
		X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",
		X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",X"AA",X"80",X"00",X"00",X"00",X"00",X"00",X"A8",
		X"A2",X"A0",X"00",X"00",X"00",X"00",X"02",X"A0",X"AA",X"A0",X"00",X"00",X"00",X"00",X"0A",X"80",
		X"AA",X"A8",X"00",X"00",X"00",X"00",X"2A",X"00",X"A8",X"2A",X"00",X"00",X"00",X"00",X"A8",X"00",
		X"A0",X"2A",X"00",X"00",X"00",X"02",X"A0",X"00",X"A0",X"AA",X"80",X"00",X"00",X"0A",X"80",X"00",
		X"A2",X"A2",X"A0",X"00",X"00",X"2A",X"00",X"00",X"AA",X"80",X"A0",X"00",X"00",X"A8",X"00",X"00",
		X"AA",X"02",X"A8",X"00",X"02",X"A0",X"00",X"00",X"A8",X"0A",X"AA",X"00",X"0A",X"80",X"00",X"00",
		X"A0",X"2A",X"0A",X"00",X"2A",X"00",X"00",X"00",X"A0",X"A8",X"0A",X"80",X"A8",X"00",X"00",X"00",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"3F",X"00",X"00",X"00",X"00",X"00",X"03",X"FF",
		X"0F",X"C0",X"00",X"00",X"00",X"00",X"0F",X"CF",X"03",X"F0",X"00",X"00",X"00",X"00",X"0F",X"FF",
		X"00",X"FC",X"00",X"00",X"00",X"00",X"3F",X"FF",X"00",X"3F",X"00",X"00",X"00",X"00",X"FC",X"3F",
		X"00",X"0F",X"C0",X"00",X"00",X"00",X"FC",X"0F",X"00",X"03",X"F0",X"00",X"00",X"03",X"FF",X"0F",
		X"00",X"00",X"FC",X"00",X"00",X"0F",X"CF",X"CF",X"00",X"00",X"3F",X"00",X"00",X"0F",X"03",X"FF",
		X"00",X"00",X"0F",X"C0",X"00",X"3F",X"C0",X"FF",X"00",X"00",X"03",X"F0",X"00",X"FF",X"F0",X"3F",
		X"00",X"00",X"00",X"FC",X"00",X"F0",X"FC",X"0F",X"00",X"00",X"00",X"3F",X"03",X"F0",X"3F",X"0F",
		X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"FF",X"C0",X"00",X"00",X"00",X"00",X"00",X"FC",
		X"F3",X"F0",X"00",X"00",X"00",X"00",X"03",X"F0",X"FF",X"F0",X"00",X"00",X"00",X"00",X"0F",X"C0",
		X"FF",X"FC",X"00",X"00",X"00",X"00",X"3F",X"00",X"FC",X"3F",X"00",X"00",X"00",X"00",X"FC",X"00",
		X"F0",X"3F",X"00",X"00",X"00",X"03",X"F0",X"00",X"F0",X"FF",X"C0",X"00",X"00",X"0F",X"C0",X"00",
		X"F3",X"F3",X"F0",X"00",X"00",X"3F",X"00",X"00",X"FF",X"C0",X"F0",X"00",X"00",X"FC",X"00",X"00",
		X"FF",X"03",X"FC",X"00",X"03",X"F0",X"00",X"00",X"FC",X"0F",X"FF",X"00",X"0F",X"C0",X"00",X"00",
		X"F0",X"3F",X"0F",X"00",X"3F",X"00",X"00",X"00",X"F0",X"FC",X"0F",X"C0",X"FC",X"00",X"00",X"00",
		X"EA",X"B0",X"EA",X"B0",X"00",X"00",X"EA",X"B0",X"EA",X"B0",X"EA",X"B0",X"00",X"00",X"EA",X"B0",
		X"EA",X"B0",X"EA",X"B0",X"00",X"00",X"EA",X"B0",X"EA",X"B0",X"EA",X"B0",X"00",X"00",X"EA",X"B0",
		X"EA",X"B0",X"EA",X"AF",X"FF",X"FF",X"AA",X"AF",X"EA",X"B0",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"EA",X"B0",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"B0",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"EA",X"B0",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"B0",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"EA",X"B0",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"B0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EA",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"EA",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EA",X"B0",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"EA",X"B0",X"EA",X"AA",X"AA",X"AA",X"C0",X"00",
		X"00",X"0E",X"AB",X"0E",X"AB",X"0E",X"AA",X"AA",X"00",X"0E",X"AB",X"0E",X"AB",X"0E",X"AA",X"AA",
		X"00",X"0E",X"AB",X"0E",X"AB",X"0E",X"AA",X"AA",X"00",X"0E",X"AB",X"0E",X"AB",X"0E",X"AA",X"BF",
		X"FF",X"FE",X"AB",X"0E",X"AB",X"0E",X"AA",X"C0",X"AA",X"AA",X"AB",X"0E",X"AB",X"0E",X"AA",X"C0",
		X"AA",X"AA",X"AB",X"0E",X"AB",X"0E",X"AA",X"C0",X"AA",X"AA",X"AB",X"0E",X"AB",X"0E",X"AA",X"C0",
		X"AA",X"AA",X"AB",X"0E",X"AB",X"0E",X"AA",X"C0",X"AA",X"AA",X"AB",X"0E",X"AB",X"0E",X"AA",X"C0",
		X"AA",X"AA",X"AB",X"0E",X"AB",X"0E",X"AA",X"BF",X"FF",X"FF",X"FF",X"0E",X"AB",X"0E",X"AA",X"AA",
		X"00",X"00",X"00",X"0E",X"AB",X"0E",X"AA",X"AA",X"00",X"00",X"00",X"0E",X"AB",X"0E",X"AA",X"AA",
		X"00",X"00",X"0F",X"0E",X"AB",X"0E",X"AA",X"AA",X"00",X"0F",X"FB",X"0E",X"AB",X"0F",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"B0",X"00",X"00",X"00",X"00",X"AA",X"FF",X"EA",X"B0",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"EA",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"EA",X"B0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"EA",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"EA",X"B0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"EA",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"EA",X"B0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"EA",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"EA",X"B0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"EA",X"B0",X"00",X"00",X"00",X"00",X"FF",X"00",X"EA",X"B0",X"00",X"00",X"00",X"00",
		X"AA",X"FF",X"EA",X"B0",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"B0",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AF",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"FF",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"0A",X"8A",X"A8",X"0A",X"8A",X"00",X"00",X"00",X"02",X"AA",X"2A",X"02",X"AA",
		X"00",X"00",X"00",X"00",X"AA",X"0A",X"80",X"AA",X"00",X"00",X"00",X"00",X"2A",X"02",X"A0",X"2A",
		X"00",X"00",X"00",X"00",X"0A",X"80",X"A8",X"0A",X"00",X"00",X"00",X"00",X"02",X"A0",X"2A",X"0A",
		X"00",X"00",X"00",X"00",X"00",X"A8",X"0A",X"8A",X"00",X"00",X"00",X"00",X"00",X"2A",X"02",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"80",X"AA",X"00",X"00",X"00",X"00",X"00",X"02",X"A0",X"2A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"A8",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",X"0A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"8A",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",
		X"A2",X"A0",X"2A",X"A2",X"A0",X"00",X"00",X"00",X"AA",X"80",X"A8",X"AA",X"80",X"00",X"00",X"00",
		X"AA",X"02",X"A0",X"AA",X"00",X"00",X"00",X"00",X"A8",X"0A",X"80",X"A8",X"00",X"00",X"00",X"00",
		X"A0",X"2A",X"02",X"A0",X"00",X"00",X"00",X"00",X"A0",X"A8",X"0A",X"80",X"00",X"00",X"00",X"00",
		X"A2",X"A0",X"2A",X"00",X"00",X"00",X"00",X"00",X"AA",X"80",X"A8",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"02",X"A0",X"00",X"00",X"00",X"00",X"00",X"A8",X"0A",X"80",X"00",X"00",X"00",X"00",X"00",
		X"A0",X"2A",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"A8",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A2",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"CF",X"FC",X"0F",X"CF",X"00",X"00",X"00",X"03",X"FF",X"3F",X"03",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"0F",X"C0",X"FF",X"00",X"00",X"00",X"00",X"3F",X"03",X"F0",X"3F",
		X"00",X"00",X"00",X"00",X"0F",X"C0",X"FC",X"0F",X"00",X"00",X"00",X"00",X"03",X"F0",X"3F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"FC",X"0F",X"CF",X"00",X"00",X"00",X"00",X"00",X"3F",X"03",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"C0",X"FF",X"00",X"00",X"00",X"00",X"00",X"03",X"F0",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"CF",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",
		X"F3",X"F0",X"3F",X"F3",X"F0",X"00",X"00",X"00",X"FF",X"C0",X"FC",X"FF",X"C0",X"00",X"00",X"00",
		X"FF",X"03",X"F0",X"FF",X"00",X"00",X"00",X"00",X"FC",X"0F",X"C0",X"FC",X"00",X"00",X"00",X"00",
		X"F0",X"3F",X"03",X"F0",X"00",X"00",X"00",X"00",X"F0",X"FC",X"0F",X"C0",X"00",X"00",X"00",X"00",
		X"F3",X"F0",X"3F",X"00",X"00",X"00",X"00",X"00",X"FF",X"C0",X"FC",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"03",X"F0",X"00",X"00",X"00",X"00",X"00",X"FC",X"0F",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F3",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EA",X"B0",X"EA",X"AA",X"AA",X"AA",X"B0",X"00",X"EA",X"B0",X"EA",X"AA",X"AA",X"AA",X"AC",X"0F",
		X"EA",X"B0",X"EA",X"AA",X"AA",X"AA",X"AB",X"FA",X"EA",X"B0",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"EA",X"B0",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"B0",X"EA",X"AF",X"FF",X"FA",X"AA",X"AA",
		X"EA",X"B0",X"EA",X"B0",X"00",X"0E",X"AA",X"AA",X"EA",X"B0",X"EA",X"B0",X"00",X"03",X"AA",X"AA",
		X"EA",X"B0",X"EA",X"B0",X"00",X"00",X"EA",X"AF",X"EA",X"B0",X"EA",X"B0",X"00",X"00",X"EA",X"B0",
		X"EA",X"B0",X"EA",X"B0",X"00",X"00",X"EA",X"B0",X"EA",X"B0",X"EA",X"B0",X"00",X"00",X"EA",X"B0",
		X"EA",X"B0",X"EA",X"B0",X"00",X"00",X"EA",X"B0",X"EA",X"B0",X"EA",X"B0",X"00",X"00",X"EA",X"B0",
		X"EA",X"B0",X"EA",X"B0",X"00",X"00",X"EA",X"B0",X"EA",X"B0",X"EA",X"AF",X"FF",X"FF",X"AA",X"AF",
		X"0F",X"FA",X"AB",X"0E",X"AB",X"00",X"FF",X"AA",X"FA",X"AA",X"AB",X"0E",X"AB",X"00",X"00",X"FF",
		X"AA",X"AA",X"AB",X"0E",X"AA",X"FF",X"00",X"00",X"AA",X"AA",X"AB",X"0E",X"AA",X"AA",X"FF",X"00",
		X"AA",X"AA",X"AB",X"0E",X"AA",X"AA",X"AA",X"FF",X"AA",X"AA",X"AF",X"0E",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AF",X"F0",X"0E",X"AA",X"AA",X"AA",X"AA",X"AF",X"F0",X"00",X"0E",X"AA",X"AA",X"AA",X"AA",
		X"F0",X"00",X"00",X"0E",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"0E",X"AA",X"FF",X"AA",X"AA",
		X"00",X"00",X"00",X"0E",X"AB",X"00",X"FF",X"AA",X"00",X"00",X"00",X"0E",X"AB",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"0E",X"AB",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"AB",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0E",X"AB",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"0E",X"AB",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"FF",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"F0",X"00",
		X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"B0",X"00",X"00",X"FF",X"AA",X"AA",X"AA",X"AA",X"B0",X"00",
		X"00",X"00",X"FF",X"AA",X"AA",X"AA",X"B0",X"00",X"FF",X"00",X"00",X"FF",X"AA",X"AA",X"B0",X"00",
		X"AA",X"FF",X"00",X"00",X"FF",X"AA",X"B0",X"00",X"AA",X"AA",X"FF",X"00",X"00",X"FF",X"B0",X"00",
		X"AA",X"AA",X"AA",X"FF",X"00",X"00",X"F0",X"00",X"AA",X"AA",X"AA",X"AA",X"FF",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"FF",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"F0",X"00",
		X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"B0",X"00",X"00",X"FF",X"AA",X"AA",X"AA",X"AA",X"B0",X"00",
		X"00",X"00",X"FF",X"AA",X"AA",X"AA",X"B0",X"00",X"00",X"00",X"00",X"FF",X"AA",X"AA",X"B0",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",
		X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"02",X"AA",
		X"AA",X"80",X"00",X"00",X"00",X"00",X"02",X"8A",X"A2",X"A0",X"00",X"00",X"00",X"00",X"0A",X"AA",
		X"A0",X"A8",X"00",X"00",X"00",X"00",X"2A",X"AA",X"A0",X"2A",X"00",X"00",X"00",X"00",X"28",X"2A",
		X"A8",X"0A",X"80",X"00",X"00",X"00",X"A8",X"0A",X"AA",X"02",X"A0",X"00",X"00",X"02",X"AA",X"0A",
		X"AA",X"80",X"A8",X"00",X"00",X"02",X"8A",X"8A",X"A2",X"A0",X"2A",X"00",X"00",X"0A",X"82",X"AA",
		X"A0",X"A8",X"0A",X"80",X"00",X"2A",X"80",X"AA",X"A0",X"2A",X"02",X"A0",X"00",X"2A",X"A0",X"2A",
		X"A8",X"0A",X"80",X"A8",X"00",X"A8",X"A8",X"0A",X"AA",X"02",X"A0",X"2A",X"02",X"A0",X"2A",X"0A",
		X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",
		X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",X"AA",X"80",X"00",X"00",X"00",X"00",X"00",X"AA",
		X"A2",X"80",X"00",X"00",X"00",X"00",X"02",X"AA",X"AA",X"A0",X"00",X"00",X"00",X"00",X"0A",X"8A",
		X"AA",X"A8",X"00",X"00",X"00",X"00",X"2A",X"0A",X"A8",X"28",X"00",X"00",X"00",X"00",X"A8",X"0A",
		X"A0",X"2A",X"00",X"00",X"00",X"02",X"A0",X"2A",X"A0",X"AA",X"80",X"00",X"00",X"0A",X"80",X"AA",
		X"A2",X"A2",X"80",X"00",X"00",X"2A",X"02",X"AA",X"AA",X"82",X"A0",X"00",X"00",X"A8",X"0A",X"8A",
		X"AA",X"02",X"A8",X"00",X"02",X"A0",X"2A",X"0A",X"A8",X"0A",X"A8",X"00",X"0A",X"80",X"A8",X"0A",
		X"A0",X"2A",X"2A",X"00",X"2A",X"02",X"A0",X"2A",X"A0",X"A8",X"0A",X"80",X"A8",X"0A",X"80",X"AA",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",
		X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"03",X"FF",
		X"FF",X"C0",X"00",X"00",X"00",X"00",X"03",X"CF",X"F3",X"F0",X"00",X"00",X"00",X"00",X"0F",X"FF",
		X"F0",X"FC",X"00",X"00",X"00",X"00",X"3F",X"FF",X"F0",X"3F",X"00",X"00",X"00",X"00",X"3C",X"3F",
		X"FC",X"0F",X"C0",X"00",X"00",X"00",X"FC",X"0F",X"FF",X"03",X"F0",X"00",X"00",X"03",X"FF",X"0F",
		X"FF",X"C0",X"FC",X"00",X"00",X"03",X"CF",X"CF",X"F3",X"F0",X"3F",X"00",X"00",X"0F",X"C3",X"FF",
		X"F0",X"FC",X"0F",X"C0",X"00",X"3F",X"C0",X"FF",X"F0",X"3F",X"03",X"F0",X"00",X"3F",X"F0",X"3F",
		X"FC",X"0F",X"C0",X"FC",X"00",X"FC",X"FC",X"0F",X"FF",X"03",X"F0",X"3F",X"03",X"F0",X"3F",X"0F",
		X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"FF",X"C0",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"F3",X"C0",X"00",X"00",X"00",X"00",X"03",X"FF",X"FF",X"F0",X"00",X"00",X"00",X"00",X"0F",X"CF",
		X"FF",X"FC",X"00",X"00",X"00",X"00",X"3F",X"0F",X"FC",X"3C",X"00",X"00",X"00",X"00",X"FC",X"0F",
		X"F0",X"3F",X"00",X"00",X"00",X"03",X"F0",X"3F",X"F0",X"FF",X"C0",X"00",X"00",X"0F",X"C0",X"FF",
		X"F3",X"F3",X"D0",X"00",X"00",X"3F",X"03",X"FF",X"FF",X"C3",X"F0",X"00",X"00",X"FC",X"0F",X"CF",
		X"FF",X"03",X"FC",X"00",X"03",X"F0",X"3F",X"0F",X"FC",X"0F",X"FC",X"00",X"0F",X"C0",X"FC",X"0F",
		X"F0",X"3F",X"3F",X"00",X"3F",X"03",X"F0",X"3F",X"F0",X"FC",X"0F",X"C0",X"FC",X"0F",X"C0",X"FF",
		X"EA",X"B0",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"B0",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"EA",X"B0",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"B0",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"EA",X"B0",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"B0",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"EA",X"B0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EA",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EA",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"EA",X"B0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EA",X"B0",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"B0",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"EA",X"B0",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"B0",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"EA",X"B0",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"B0",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AB",X"0E",X"AB",X"00",X"00",X"00",X"AA",X"AA",X"AB",X"0E",X"AB",X"00",X"00",X"00",
		X"AA",X"AA",X"AB",X"0E",X"AB",X"00",X"00",X"00",X"AA",X"AA",X"AB",X"0E",X"AB",X"00",X"00",X"00",
		X"AA",X"AA",X"AB",X"0E",X"AB",X"00",X"00",X"00",X"AA",X"AA",X"AB",X"0E",X"AB",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"0E",X"AB",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"AB",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0E",X"AB",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"0E",X"AB",X"00",X"00",X"00",
		X"AA",X"AA",X"AB",X"0E",X"AB",X"00",X"00",X"00",X"AA",X"AA",X"AB",X"0E",X"AB",X"00",X"00",X"00",
		X"AA",X"AA",X"AB",X"0E",X"AB",X"00",X"00",X"00",X"AA",X"AA",X"AB",X"0E",X"AB",X"00",X"00",X"00",
		X"AA",X"AA",X"AB",X"0F",X"EB",X"00",X"00",X"00",X"AA",X"AA",X"AB",X"00",X"3F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"AA",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"B0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"80",X"A8",X"0A",X"82",X"A8",X"0A",X"8A",X"A2",X"A0",X"2A",X"02",X"AA",X"AA",X"02",X"AA",
		X"A0",X"A8",X"0A",X"80",X"AA",X"0A",X"80",X"AA",X"A0",X"2A",X"02",X"A0",X"2A",X"02",X"A0",X"2A",
		X"A8",X"0A",X"80",X"A8",X"0A",X"80",X"A8",X"0A",X"AA",X"02",X"A0",X"2A",X"02",X"A0",X"2A",X"0A",
		X"AA",X"80",X"A8",X"0A",X"80",X"A8",X"0A",X"8A",X"A2",X"A0",X"2A",X"02",X"A0",X"2A",X"02",X"AA",
		X"A0",X"A8",X"0A",X"80",X"A8",X"0A",X"80",X"AA",X"A0",X"2A",X"02",X"A0",X"2A",X"02",X"A0",X"2A",
		X"A8",X"0A",X"80",X"A8",X"0A",X"80",X"A8",X"0A",X"AA",X"02",X"A0",X"2A",X"02",X"A0",X"2A",X"0A",
		X"AA",X"80",X"A8",X"0A",X"80",X"A8",X"0A",X"8A",X"A2",X"A0",X"2A",X"02",X"A0",X"2A",X"02",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"A2",X"A0",X"2A",X"82",X"A0",X"2A",X"02",X"AA",X"AA",X"80",X"AA",X"AA",X"80",X"A8",X"0A",X"8A",
		X"AA",X"02",X"A0",X"AA",X"02",X"A0",X"2A",X"0A",X"A8",X"0A",X"80",X"A8",X"0A",X"80",X"A8",X"0A",
		X"A0",X"2A",X"02",X"A0",X"2A",X"02",X"A0",X"2A",X"A0",X"A8",X"0A",X"80",X"A8",X"0A",X"80",X"AA",
		X"A2",X"A0",X"2A",X"02",X"A0",X"2A",X"02",X"AA",X"AA",X"80",X"A8",X"0A",X"80",X"A8",X"0A",X"8A",
		X"AA",X"02",X"A0",X"2A",X"02",X"A0",X"2A",X"0A",X"A8",X"0A",X"80",X"A8",X"0A",X"80",X"A8",X"0A",
		X"A0",X"2A",X"02",X"A0",X"2A",X"02",X"A0",X"2A",X"A0",X"A8",X"0A",X"80",X"A8",X"0A",X"80",X"AA",
		X"A2",X"A0",X"2A",X"02",X"A0",X"2A",X"02",X"AA",X"AA",X"80",X"A8",X"0A",X"80",X"A8",X"0A",X"8A",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"C0",X"FC",X"0F",X"C3",X"FC",X"0F",X"CF",X"F3",X"F0",X"3F",X"03",X"FF",X"FF",X"03",X"FF",
		X"F0",X"FC",X"0F",X"C0",X"FF",X"0F",X"C0",X"FF",X"F0",X"3F",X"03",X"F0",X"3F",X"03",X"F0",X"3F",
		X"FC",X"0F",X"C0",X"FC",X"0F",X"C0",X"FC",X"0F",X"FF",X"03",X"F0",X"3F",X"03",X"F0",X"3F",X"0F",
		X"FF",X"C0",X"FC",X"0F",X"C0",X"FC",X"0F",X"CF",X"F3",X"F0",X"3F",X"03",X"F0",X"3F",X"03",X"FF",
		X"F0",X"FC",X"0F",X"C0",X"FC",X"0F",X"C0",X"FF",X"F0",X"3F",X"03",X"F0",X"3F",X"03",X"F0",X"3F",
		X"FC",X"0F",X"C0",X"FC",X"0F",X"C0",X"FC",X"0F",X"FF",X"03",X"F0",X"3F",X"03",X"F0",X"3F",X"0F",
		X"FF",X"C0",X"FC",X"0F",X"C0",X"FC",X"0F",X"CF",X"F3",X"F0",X"3F",X"03",X"F0",X"3F",X"03",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F3",X"F0",X"3F",X"C3",X"F0",X"3F",X"03",X"FF",X"FF",X"C0",X"FF",X"FF",X"C0",X"FC",X"0F",X"CF",
		X"FF",X"03",X"F0",X"FF",X"03",X"F0",X"3F",X"0F",X"FC",X"0F",X"C0",X"FC",X"0F",X"C0",X"FC",X"0F",
		X"F0",X"3F",X"03",X"F0",X"3F",X"03",X"F0",X"3F",X"F0",X"FC",X"0F",X"C0",X"FC",X"0F",X"C0",X"FF",
		X"F3",X"F0",X"3F",X"03",X"F0",X"3F",X"03",X"FF",X"FF",X"C0",X"FC",X"0F",X"C0",X"FC",X"0F",X"CF",
		X"FF",X"03",X"F0",X"3F",X"03",X"F0",X"3F",X"0F",X"FC",X"0F",X"C0",X"FC",X"0F",X"C0",X"FC",X"0F",
		X"F0",X"3F",X"03",X"F0",X"3F",X"03",X"F0",X"3F",X"F0",X"FC",X"0F",X"C0",X"FC",X"0F",X"C0",X"FF",
		X"F3",X"F0",X"3F",X"03",X"F0",X"3F",X"03",X"FF",X"FF",X"C0",X"FC",X"0F",X"C0",X"FC",X"0F",X"CF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EA",X"B0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EA",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EA",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"EA",X"B0",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"EA",X"B0",X"EF",X"F0",X"00",X"00",X"00",X"00",X"EA",X"B0",X"EA",X"AF",X"F0",X"00",X"00",X"00",
		X"EA",X"B0",X"EA",X"AA",X"AF",X"F0",X"00",X"00",X"EA",X"B0",X"EA",X"AA",X"AA",X"AF",X"F0",X"00",
		X"EA",X"B0",X"EA",X"AA",X"AA",X"AA",X"AF",X"F0",X"EA",X"B0",X"EA",X"AA",X"AA",X"AA",X"AA",X"AF",
		X"EA",X"B0",X"FA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"B0",X"0F",X"FA",X"AA",X"AA",X"AA",X"AA",
		X"EA",X"B0",X"00",X"0F",X"FA",X"AA",X"AA",X"AA",X"EA",X"AF",X"F0",X"00",X"0F",X"FA",X"AA",X"AA",
		X"EA",X"AA",X"AF",X"F0",X"00",X"0F",X"FA",X"AA",X"EA",X"AA",X"AA",X"AF",X"F0",X"00",X"0F",X"FA",
		X"FF",X"FE",X"AB",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"AB",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"AB",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"AB",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"AB",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"AB",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"AB",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"AB",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"AB",X"00",X"00",X"00",X"00",X"00",X"F0",X"0E",X"AB",X"00",X"00",X"00",X"00",X"00",
		X"AF",X"FA",X"AB",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AB",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AB",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AB",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AB",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AB",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"55",X"00",X"55",X"55",X"55",X"55",X"55",X"00",X"00",
		X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"00",X"55",X"00",X"00",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"00",X"00",X"55",X"55",X"00",X"55",X"55",X"55",X"55",X"00",X"00",X"55",
		X"00",X"00",X"55",X"55",X"55",X"55",X"00",X"00",X"55",X"00",X"00",X"55",X"55",X"55",X"55",X"00",
		X"55",X"55",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"01",X"55",
		X"55",X"55",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"55",X"55",X"55",X"00",X"00",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"00",X"00",X"FF",X"FF",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"3F",
		X"00",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"00",
		X"55",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"55",X"00",X"55",X"55",X"55",X"55",X"55",X"00",X"00",
		X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"00",X"55",X"00",X"00",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"F0",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"F0",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"55",X"00",X"00",X"FF",X"FF",X"FF",X"F0",X"00",
		X"55",X"55",X"00",X"00",X"FF",X"FF",X"F0",X"00",X"55",X"55",X"55",X"00",X"00",X"FF",X"F0",X"00",
		X"55",X"55",X"55",X"54",X"00",X"00",X"F0",X"00",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"00",
		X"00",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"50",X"00",
		X"55",X"00",X"00",X"55",X"55",X"55",X"50",X"00",X"55",X"55",X"00",X"00",X"55",X"55",X"50",X"00",
		X"55",X"55",X"55",X"55",X"55",X"5A",X"AA",X"AA",X"55",X"55",X"55",X"55",X"55",X"5A",X"AA",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"5A",X"AA",X"82",X"55",X"55",X"55",X"55",X"55",X"5A",X"AA",X"82",
		X"55",X"55",X"55",X"55",X"55",X"5A",X"A0",X"82",X"55",X"55",X"55",X"55",X"55",X"5A",X"A0",X"AA",
		X"55",X"55",X"55",X"55",X"AA",X"AA",X"A0",X"AA",X"55",X"55",X"55",X"55",X"8A",X"AA",X"AA",X"AA",
		X"55",X"55",X"55",X"55",X"8A",X"A8",X"AA",X"AA",X"55",X"55",X"55",X"55",X"AA",X"AA",X"AA",X"AA",
		X"55",X"55",X"55",X"55",X"AA",X"AA",X"AA",X"82",X"55",X"55",X"55",X"55",X"AA",X"AA",X"AA",X"82",
		X"55",X"55",X"55",X"55",X"AA",X"AA",X"AA",X"82",X"55",X"55",X"55",X"55",X"AA",X"A8",X"0A",X"A2",
		X"55",X"55",X"55",X"55",X"AA",X"A8",X"0A",X"AA",X"55",X"55",X"55",X"55",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EA",X"AA",X"AA",X"AA",X"AF",X"F0",X"00",X"0F",X"EA",X"AA",X"AA",X"AA",X"AA",X"AF",X"F0",X"00",
		X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AF",X"F0",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AF",
		X"EA",X"AF",X"FA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"B0",X"0F",X"FA",X"AA",X"AA",X"AA",X"AA",
		X"EA",X"B0",X"00",X"0F",X"FA",X"AA",X"AA",X"AA",X"EA",X"B0",X"00",X"00",X"0F",X"FA",X"AA",X"AA",
		X"EA",X"B0",X"FF",X"00",X"00",X"0F",X"FA",X"AA",X"EA",X"B0",X"FF",X"FF",X"00",X"00",X"0F",X"FA",
		X"EA",X"B0",X"FF",X"FF",X"FF",X"00",X"00",X"0F",X"EA",X"B0",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"EA",X"B0",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"EA",X"B0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EA",X"B0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EA",X"B0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FA",X"AA",X"AB",X"00",X"00",X"00",X"00",X"00",X"0F",X"FA",X"AB",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"FB",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"AF",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AF",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AF",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AB",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AB",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AB",X"00",X"00",X"00",X"00",X"00",
		X"FA",X"AA",X"AB",X"00",X"00",X"00",X"00",X"00",X"0F",X"FA",X"AB",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"FB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"A8",X"25",X"55",X"55",X"55",X"55",X"55",X"AA",X"A8",X"25",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"A8",X"25",X"55",X"55",X"55",X"55",X"55",X"AA",X"AA",X"A5",X"55",X"55",X"55",X"55",X"55",
		X"82",X"AA",X"A5",X"55",X"55",X"55",X"55",X"55",X"82",X"AA",X"A5",X"55",X"55",X"55",X"55",X"55",
		X"82",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"2A",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"A0",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"A2",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"82",X"AA",X"02",X"AA",X"02",X"AA",X"02",
		X"82",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"8A",X"A0",X"2A",X"AA",X"AA",X"A0",X"2A",X"AA",
		X"AA",X"A0",X"2A",X"AA",X"AA",X"A0",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"5A",X"AA",X"AA",X"55",X"55",X"55",X"55",X"55",X"5A",X"AA",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"5A",X"AA",X"AA",X"55",X"55",X"55",X"55",X"55",X"5A",X"A0",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"5A",X"A0",X"AA",X"55",X"55",X"55",X"55",X"55",X"5A",X"A0",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"2A",X"A0",X"2A",X"A2",X"AA",X"AA",
		X"AA",X"A0",X"2A",X"A0",X"2A",X"A0",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"82",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"02",X"AA",X"82",X"AA",X"AA",X"AA",X"AA",X"AA",X"02",X"AA",X"82",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"82",X"AA",X"AA",X"A0",X"2A",X"AA",X"AA",X"AA",X"A2",
		X"AA",X"AA",X"A0",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"5D",X"FF",X"00",X"00",X"77",X"C0",X"00",X"00",X"57",X"FF",X"00",X"00",X"5F",X"C0",X"00",X"00",
		X"5D",X"FF",X"00",X"00",X"77",X"C0",X"00",X"00",X"57",X"FF",X"00",X"00",X"5F",X"C0",X"00",X"00",
		X"5D",X"FF",X"00",X"00",X"77",X"C0",X"00",X"00",X"57",X"FF",X"00",X"00",X"5F",X"C0",X"00",X"00",
		X"5D",X"FF",X"00",X"00",X"77",X"C0",X"00",X"00",X"57",X"FF",X"00",X"00",X"5F",X"C0",X"00",X"00",
		X"5D",X"FF",X"00",X"00",X"77",X"C0",X"00",X"00",X"57",X"FF",X"00",X"00",X"5F",X"C0",X"00",X"00",
		X"5D",X"FF",X"00",X"00",X"77",X"C0",X"00",X"00",X"57",X"FF",X"00",X"00",X"5F",X"7F",X"FF",X"FF",
		X"5D",X"FF",X"00",X"00",X"75",X"FF",X"FF",X"FF",X"57",X"FF",X"00",X"00",X"5D",X"DD",X"DD",X"DD",
		X"5D",X"FF",X"00",X"00",X"77",X"77",X"77",X"77",X"57",X"FF",X"00",X"00",X"55",X"55",X"55",X"55",
		X"00",X"00",X"03",X"F5",X"00",X"00",X"FF",X"D5",X"00",X"00",X"03",X"DD",X"00",X"00",X"FF",X"75",
		X"00",X"00",X"03",X"F5",X"00",X"00",X"FF",X"D5",X"00",X"00",X"03",X"DD",X"00",X"00",X"FF",X"75",
		X"00",X"00",X"03",X"F5",X"00",X"00",X"FF",X"D5",X"00",X"00",X"03",X"DD",X"00",X"00",X"FF",X"75",
		X"00",X"00",X"03",X"F5",X"00",X"00",X"FF",X"D5",X"00",X"00",X"03",X"DD",X"00",X"00",X"FF",X"75",
		X"00",X"00",X"03",X"F5",X"00",X"00",X"FF",X"D5",X"00",X"00",X"03",X"DD",X"00",X"00",X"FF",X"75",
		X"00",X"00",X"03",X"F5",X"00",X"00",X"FF",X"D5",X"FF",X"FF",X"FD",X"DD",X"00",X"00",X"FF",X"75",
		X"FF",X"FF",X"FF",X"75",X"00",X"00",X"FF",X"D5",X"DD",X"DD",X"DD",X"DD",X"00",X"00",X"FF",X"75",
		X"77",X"77",X"77",X"75",X"00",X"00",X"FF",X"D5",X"55",X"55",X"55",X"55",X"00",X"00",X"FF",X"75",
		X"AA",X"AA",X"A4",X"44",X"00",X"00",X"00",X"00",X"AA",X"AA",X"A5",X"11",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"A4",X"44",X"00",X"00",X"00",X"00",X"AA",X"0A",X"A5",X"14",X"00",X"00",X"00",X"00",
		X"AA",X"0A",X"A4",X"44",X"00",X"00",X"00",X"00",X"AA",X"0A",X"A5",X"55",X"00",X"00",X"00",X"00",
		X"AA",X"0A",X"AA",X"AA",X"00",X"00",X"00",X"00",X"AA",X"AA",X"A0",X"2A",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"A0",X"2A",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",
		X"82",X"AA",X"AA",X"02",X"00",X"00",X"00",X"00",X"82",X"AA",X"AA",X"02",X"00",X"00",X"00",X"00",
		X"82",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",X"8A",X"A0",X"2A",X"AA",X"00",X"00",X"00",X"00",
		X"AA",X"A0",X"2A",X"AA",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",
		X"EA",X"B0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EA",X"B0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EA",X"B0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EA",X"B0",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EA",X"B0",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"EA",X"B0",X"FF",X"00",X"00",X"FF",X"FF",X"FF",
		X"EA",X"B0",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"EA",X"B0",X"FF",X"FF",X"FF",X"00",X"00",X"FF",
		X"EA",X"B0",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"EA",X"B0",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"EA",X"B0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"B0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"03",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"00",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"03",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",
		X"AA",X"AA",X"A5",X"55",X"55",X"55",X"55",X"55",X"AA",X"A8",X"25",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"A8",X"25",X"55",X"55",X"55",X"55",X"55",X"AA",X"A8",X"25",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"A5",X"55",X"55",X"55",X"55",X"55",X"AA",X"AA",X"A5",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"A5",X"55",X"55",X"55",X"55",X"55",X"AA",X"AA",X"A5",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"A5",X"55",X"55",X"55",X"55",X"55",X"82",X"A8",X"25",X"55",X"55",X"55",X"55",X"55",
		X"82",X"A8",X"25",X"55",X"55",X"55",X"55",X"55",X"82",X"A8",X"25",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"A5",X"55",X"55",X"55",X"55",X"55",X"AA",X"AA",X"A5",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"A5",X"55",X"55",X"55",X"55",X"55",X"AA",X"AA",X"A5",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"5D",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"57",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"5D",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"57",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"5D",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"57",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"5D",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"57",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"5D",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"57",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"5D",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"57",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"5D",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"57",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"5D",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"57",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"D5",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"75",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"D5",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"75",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"D5",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"75",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"D5",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"75",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"D5",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"75",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"D5",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"75",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"D5",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"75",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"D5",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"75",
		X"6A",X"AA",X"00",X"00",X"00",X"00",X"AA",X"A9",X"6A",X"82",X"0C",X"30",X"C3",X"0C",X"AA",X"09",
		X"6A",X"82",X"30",X"C3",X"0C",X"30",X"AA",X"09",X"6A",X"82",X"03",X"0C",X"30",X"C0",X"AA",X"09",
		X"6A",X"AA",X"0C",X"30",X"C3",X"0C",X"AA",X"A9",X"6A",X"AA",X"30",X"C3",X"0C",X"30",X"AA",X"A9",
		X"A0",X"AA",X"00",X"00",X"00",X"00",X"AA",X"AA",X"A0",X"AA",X"11",X"11",X"11",X"11",X"AA",X"AA",
		X"A0",X"AA",X"44",X"44",X"44",X"44",X"AA",X"AA",X"AA",X"AA",X"11",X"11",X"11",X"11",X"AA",X"AA",
		X"AA",X"AA",X"44",X"44",X"44",X"44",X"AA",X"AA",X"AA",X"AA",X"11",X"11",X"11",X"11",X"82",X"AA",
		X"AA",X"AA",X"44",X"44",X"54",X"44",X"82",X"AA",X"AA",X"AA",X"15",X"11",X"51",X"15",X"8A",X"AA",
		X"AA",X"AA",X"45",X"55",X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"55",X"55",X"55",X"55",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"00",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"03",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"03",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"55",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"55",X"55",X"55",X"00",X"00",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"00",X"00",X"FF",X"FF",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"FF",
		X"01",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"01",X"55",X"55",X"55",X"55",X"55",X"00",
		X"55",X"00",X"01",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"01",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"00",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"03",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"00",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"03",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"03",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"55",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"F0",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"F0",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"F0",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"F0",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",
		X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"00",X"03",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",
		X"FF",X"00",X"03",X"FF",X"FF",X"FF",X"F0",X"00",X"FF",X"FF",X"00",X"03",X"FF",X"FF",X"F0",X"00",
		X"55",X"55",X"55",X"55",X"55",X"5A",X"AA",X"AA",X"55",X"55",X"55",X"55",X"55",X"58",X"2A",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"58",X"2A",X"AA",X"55",X"55",X"55",X"55",X"55",X"58",X"2A",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"5A",X"AA",X"AA",X"55",X"55",X"55",X"55",X"55",X"5A",X"AA",X"82",
		X"55",X"55",X"55",X"55",X"55",X"5A",X"AA",X"82",X"55",X"55",X"55",X"55",X"55",X"5A",X"AA",X"82",
		X"55",X"55",X"55",X"55",X"55",X"5A",X"AA",X"AA",X"55",X"55",X"55",X"55",X"55",X"5A",X"AA",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"5A",X"AA",X"AA",X"55",X"55",X"55",X"55",X"55",X"5A",X"A0",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"5A",X"A0",X"AA",X"55",X"55",X"55",X"55",X"55",X"5A",X"A0",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"5A",X"AA",X"AA",X"55",X"55",X"55",X"55",X"55",X"5A",X"AA",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"2A",X"AA",X"AA",X"AA",X"A8",X"0A",X"AA",
		X"A0",X"2A",X"AA",X"AA",X"AA",X"A8",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"80",X"AA",X"80",X"AA",X"AA",X"AA",X"AA",X"AA",X"80",X"AA",X"80",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"2A",X"AA",X"AA",X"AA",X"A8",X"0A",
		X"AA",X"A0",X"2A",X"AA",X"AA",X"AA",X"A8",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"5D",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"57",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"5D",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"57",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"5D",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"57",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"5D",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"57",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"5D",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"57",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"5D",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"57",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"5D",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"57",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"D5",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"75",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"D5",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"75",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"D5",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"75",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"D5",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"75",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"D5",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"75",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"D5",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"75",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"D5",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"75",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",X"A8",X"0A",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"A8",X"0A",X"AA",X"A2",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"82",
		X"00",X"00",X"00",X"00",X"80",X"AA",X"82",X"82",X"00",X"00",X"00",X"00",X"80",X"AA",X"8A",X"82",
		X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"15",X"5A",X"A0",X"AA",X"00",X"00",X"00",X"00",X"04",X"5A",X"A0",X"AA",
		X"00",X"00",X"00",X"00",X"11",X"5A",X"A0",X"AA",X"00",X"00",X"00",X"00",X"04",X"5A",X"A0",X"AA",
		X"00",X"00",X"00",X"00",X"51",X"1A",X"AA",X"AA",X"00",X"00",X"00",X"00",X"14",X"5A",X"AA",X"AA",
		X"AA",X"AA",X"A4",X"54",X"04",X"44",X"44",X"00",X"AA",X"AA",X"A5",X"11",X"11",X"11",X"15",X"11",
		X"AA",X"AA",X"A4",X"44",X"44",X"44",X"44",X"44",X"AA",X"AA",X"A5",X"11",X"11",X"11",X"11",X"11",
		X"AA",X"AA",X"A4",X"44",X"54",X"44",X"44",X"54",X"AA",X"AA",X"A5",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"82",X"AA",X"AA",X"AA",X"A8",X"02",X"AA",X"AA",
		X"82",X"AA",X"AA",X"AA",X"A8",X"02",X"AA",X"AA",X"82",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"80",X"AA",X"AA",X"AA",X"A0",X"2A",X"AA",X"AA",X"80",X"AA",X"AA",X"AA",X"A0",X"2A",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"0A",X"AA",X"AA",X"A8",X"02",X"AA",X"AA",
		X"A0",X"0A",X"AA",X"AA",X"A8",X"02",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"40",X"14",X"04",X"40",X"44",X"5A",X"AA",X"AA",X"11",X"11",X"11",X"11",X"11",X"1A",X"AA",X"AA",
		X"54",X"54",X"44",X"45",X"45",X"5A",X"AA",X"AA",X"11",X"11",X"11",X"11",X"11",X"1A",X"AA",X"82",
		X"44",X"44",X"44",X"44",X"44",X"5A",X"AA",X"82",X"55",X"55",X"55",X"55",X"55",X"5A",X"A0",X"82",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"AA",X"AA",X"AA",X"02",X"AA",X"02",X"AA",X"A0",X"AA",
		X"AA",X"AA",X"02",X"AA",X"02",X"AA",X"A0",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"AA",
		X"AA",X"A0",X"2A",X"AA",X"AA",X"AA",X"A8",X"AA",X"AA",X"A0",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"02",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"02",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"A5",X"10",X"00",X"00",X"00",X"00",X"AA",X"A8",X"24",X"44",X"00",X"00",X"00",X"00",
		X"AA",X"A8",X"25",X"10",X"00",X"00",X"00",X"00",X"AA",X"A8",X"24",X"44",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"A5",X"15",X"00",X"00",X"00",X"00",X"82",X"AA",X"A4",X"44",X"00",X"00",X"00",X"00",
		X"82",X"AA",X"A5",X"10",X"00",X"00",X"00",X"00",X"82",X"AA",X"A4",X"44",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"A5",X"11",X"00",X"00",X"00",X"00",X"AA",X"AA",X"A4",X"44",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"A5",X"51",X"00",X"00",X"00",X"00",X"AA",X"0A",X"A4",X"44",X"00",X"00",X"00",X"00",
		X"AA",X"0A",X"A5",X"15",X"00",X"00",X"00",X"00",X"AA",X"0A",X"A4",X"44",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"A5",X"11",X"00",X"00",X"00",X"00",X"AA",X"AA",X"A4",X"44",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"1A",X"AA",X"AA",X"00",X"00",X"00",X"00",X"44",X"58",X"2A",X"AA",
		X"00",X"00",X"00",X"00",X"11",X"18",X"2A",X"AA",X"00",X"00",X"00",X"00",X"45",X"58",X"2A",X"AA",
		X"00",X"00",X"00",X"00",X"11",X"1A",X"AA",X"AA",X"00",X"00",X"00",X"00",X"04",X"5A",X"AA",X"82",
		X"00",X"00",X"00",X"00",X"11",X"5A",X"AA",X"82",X"00",X"00",X"00",X"00",X"44",X"5A",X"A0",X"82",
		X"00",X"00",X"00",X"00",X"11",X"1A",X"A0",X"AA",X"00",X"00",X"00",X"00",X"44",X"5A",X"A0",X"AA",
		X"00",X"00",X"00",X"00",X"11",X"1A",X"AA",X"AA",X"00",X"00",X"00",X"00",X"44",X"5A",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"15",X"1A",X"AA",X"AA",X"00",X"00",X"00",X"00",X"44",X"58",X"2A",X"AA",
		X"00",X"00",X"00",X"00",X"11",X"18",X"2A",X"AA",X"00",X"00",X"00",X"00",X"04",X"58",X"2A",X"AA",
		X"50",X"01",X"11",X"01",X"00",X"11",X"10",X"04",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"51",X"11",X"15",X"11",X"11",X"11",X"11",X"51",X"44",X"54",X"44",X"44",X"44",X"54",X"44",X"44",
		X"51",X"11",X"51",X"11",X"51",X"11",X"15",X"11",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"0A",X"A8",X"0A",X"AA",
		X"AA",X"AA",X"AA",X"A8",X"0A",X"A8",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"02",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"02",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"0A",X"A8",X"0A",X"A8",X"0A",
		X"AA",X"AA",X"A0",X"0A",X"A8",X"0A",X"A8",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"01",X"11",X"11",X"00",X"00",X"00",X"00",X"0C",X"30",X"44",X"45",
		X"00",X"00",X"00",X"00",X"03",X"0D",X"11",X"15",X"00",X"00",X"00",X"00",X"00",X"C0",X"44",X"45",
		X"00",X"00",X"00",X"00",X"0C",X"31",X"11",X"11",X"00",X"00",X"00",X"00",X"03",X"0C",X"44",X"55",
		X"00",X"00",X"00",X"00",X"00",X"C1",X"11",X"15",X"00",X"00",X"00",X"00",X"0C",X"30",X"44",X"45",
		X"00",X"00",X"00",X"00",X"03",X"0D",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"C0",X"44",X"45",
		X"00",X"00",X"00",X"00",X"0C",X"31",X"11",X"15",X"00",X"00",X"00",X"00",X"03",X"0C",X"44",X"55",
		X"00",X"00",X"00",X"00",X"00",X"C1",X"11",X"15",X"00",X"00",X"00",X"00",X"0C",X"30",X"44",X"55",
		X"00",X"00",X"00",X"00",X"03",X"0D",X"11",X"51",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"45",
		X"55",X"11",X"10",X"00",X"00",X"00",X"00",X"00",X"54",X"44",X"47",X"0C",X"00",X"00",X"00",X"00",
		X"51",X"11",X"10",X"C3",X"00",X"00",X"00",X"00",X"54",X"44",X"44",X"30",X"00",X"00",X"00",X"00",
		X"51",X"11",X"13",X"0C",X"00",X"00",X"00",X"00",X"44",X"44",X"44",X"C3",X"00",X"00",X"00",X"00",
		X"55",X"11",X"10",X"30",X"00",X"00",X"00",X"00",X"54",X"44",X"47",X"0C",X"00",X"00",X"00",X"00",
		X"55",X"11",X"10",X"C3",X"00",X"00",X"00",X"00",X"44",X"44",X"44",X"30",X"00",X"00",X"00",X"00",
		X"51",X"11",X"13",X"0C",X"00",X"00",X"00",X"00",X"44",X"44",X"44",X"C3",X"00",X"00",X"00",X"00",
		X"51",X"11",X"10",X"30",X"00",X"00",X"00",X"00",X"54",X"44",X"47",X"0C",X"00",X"00",X"00",X"00",
		X"51",X"11",X"10",X"C3",X"00",X"00",X"00",X"00",X"44",X"44",X"44",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
