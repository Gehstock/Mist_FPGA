library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity HJ7 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of HJ7 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"3C",X"7E",X"7E",X"7E",X"7E",X"3C",X"18",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"3C",X"7E",X"7E",X"7E",X"7E",X"3C",X"18",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"3C",X"7E",X"7E",X"7E",X"7E",X"3C",X"18",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"3C",X"7E",X"7E",X"7E",X"7E",X"3C",X"18",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"38",X"7C",X"FE",X"FE",X"FE",X"7C",X"38",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"38",X"7C",X"FE",X"FE",X"FE",X"7C",X"38",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"78",X"FC",X"FE",X"FE",X"FC",X"78",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"78",X"FC",X"FE",X"FE",X"FC",X"78",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"0C",X"00",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"70",X"F8",X"FC",X"F8",X"70",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"70",X"F8",X"FC",X"F8",X"70",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"70",X"F8",X"FC",X"F8",X"70",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"70",X"F8",X"FC",X"F8",X"70",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"86",X"70",X"80",X"70",X"00",X"40",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"06",X"60",X"90",X"20",X"40",X"80",X"40",X"00",X"00",X"00",X"00",
		X"22",X"77",X"EA",X"7C",X"3E",X"7F",X"BE",X"7C",X"3E",X"7F",X"BE",X"7C",X"1E",X"7F",X"EA",X"44",
		X"5C",X"EC",X"7E",X"FF",X"7E",X"EC",X"5E",X"3B",X"3B",X"5E",X"EC",X"7E",X"FF",X"7E",X"EC",X"5C",
		X"00",X"24",X"76",X"2C",X"3C",X"14",X"2E",X"5F",X"73",X"3E",X"04",X"3C",X"2C",X"76",X"24",X"00",
		X"00",X"00",X"00",X"00",X"18",X"08",X"2C",X"12",X"24",X"1A",X"01",X"0C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"18",X"1C",X"1C",X"0C",X"3C",X"3C",X"18",X"2C",X"18",X"34",X"2C",X"1C",X"3C",X"38",X"18",
		X"00",X"06",X"07",X"07",X"0F",X"0F",X"0F",X"04",X"0D",X"0B",X"07",X"0F",X"0F",X"0F",X"0E",X"06",
		X"00",X"00",X"00",X"00",X"02",X"03",X"00",X"03",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"03",X"00",X"03",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"4A",X"00",X"42",X"01",X"80",X"02",X"89",X"52",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"9D",X"B4",X"49",X"A6",X"C2",X"A1",X"6A",X"45",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FE",X"7F",X"E7",X"67",X"FE",X"7F",X"2A",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"FC",X"26",X"22",X"26",X"FC",X"F8",X"00",
		X"FE",X"FE",X"92",X"92",X"92",X"FE",X"6C",X"00",X"38",X"7C",X"C6",X"82",X"82",X"C6",X"44",X"00",
		X"FE",X"FE",X"82",X"82",X"C6",X"7C",X"38",X"00",X"FE",X"FE",X"92",X"92",X"92",X"82",X"80",X"00",
		X"FE",X"FE",X"12",X"12",X"12",X"12",X"02",X"00",X"38",X"7C",X"C6",X"82",X"92",X"F2",X"F2",X"00",
		X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",X"82",X"82",X"FE",X"FE",X"82",X"82",X"00",X"00",
		X"40",X"C0",X"80",X"80",X"80",X"FE",X"7E",X"00",X"FE",X"FE",X"30",X"78",X"EC",X"C6",X"82",X"00",
		X"FE",X"FE",X"80",X"80",X"80",X"80",X"80",X"00",X"FE",X"FE",X"1C",X"38",X"1C",X"FE",X"FE",X"00",
		X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",X"00",
		X"FE",X"FE",X"22",X"22",X"22",X"3E",X"1C",X"00",X"7C",X"FE",X"82",X"A2",X"E2",X"7E",X"BC",X"00",
		X"FE",X"FE",X"22",X"62",X"F2",X"DE",X"8C",X"00",X"4C",X"DE",X"92",X"92",X"96",X"F4",X"60",X"00",
		X"02",X"02",X"FE",X"FE",X"02",X"02",X"00",X"00",X"7E",X"FE",X"80",X"80",X"80",X"FE",X"7E",X"00",
		X"1E",X"3E",X"70",X"E0",X"70",X"3E",X"1E",X"00",X"FE",X"FE",X"70",X"38",X"70",X"FE",X"FE",X"00",
		X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",X"0E",X"1E",X"F0",X"F0",X"1E",X"0E",X"00",X"00",
		X"C2",X"E2",X"F2",X"BA",X"9E",X"8E",X"86",X"00",X"3C",X"42",X"BD",X"C3",X"C3",X"A5",X"42",X"3C",
		X"3C",X"42",X"FD",X"93",X"93",X"8D",X"42",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"2E",X"10",X"08",X"94",X"CA",X"A8",X"90",X"00",X"18",X"3C",X"FE",X"FF",X"FE",X"3C",X"18",X"00",
		X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",X"00",X"80",X"84",X"FE",X"FE",X"80",X"80",X"00",X"00",
		X"C4",X"E6",X"F2",X"B2",X"BA",X"9E",X"8C",X"00",X"40",X"C2",X"92",X"9A",X"9E",X"F6",X"62",X"00",
		X"30",X"38",X"2C",X"26",X"FE",X"FE",X"20",X"00",X"4E",X"CE",X"8A",X"8A",X"8A",X"FA",X"70",X"00",
		X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",X"00",X"06",X"06",X"E2",X"F2",X"1A",X"0E",X"06",X"00",
		X"6C",X"9E",X"9A",X"B2",X"B2",X"EC",X"60",X"00",X"0C",X"9E",X"92",X"92",X"D2",X"7E",X"3C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"0E",X"02",X"0E",X"06",X"0C",X"00",X"00",X"0C",X"0E",X"0E",X"0E",X"0E",X"0C",X"00",
		X"00",X"0C",X"0E",X"6E",X"2E",X"0E",X"0C",X"00",X"00",X"0C",X"0E",X"6E",X"6E",X"0E",X"0C",X"00",
		X"0C",X"02",X"01",X"01",X"01",X"01",X"02",X"0C",X"1C",X"02",X"31",X"01",X"11",X"01",X"12",X"0C",
		X"1C",X"02",X"31",X"11",X"11",X"31",X"12",X"1C",X"1C",X"12",X"F1",X"91",X"91",X"F1",X"12",X"1C",
		X"00",X"00",X"00",X"00",X"3C",X"7E",X"7E",X"7E",X"7E",X"3C",X"18",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"3C",X"7E",X"7E",X"7E",X"7E",X"3C",X"18",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"3C",X"7E",X"7E",X"7E",X"7E",X"3C",X"18",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"3C",X"7E",X"7E",X"7E",X"7E",X"3C",X"18",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"38",X"7C",X"FE",X"FE",X"FE",X"7C",X"38",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"38",X"7C",X"FE",X"FE",X"FE",X"7C",X"38",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"78",X"FC",X"FE",X"FE",X"FC",X"78",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"78",X"FC",X"FE",X"FE",X"FC",X"78",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"70",X"F8",X"FC",X"F8",X"70",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"70",X"F8",X"FC",X"F8",X"70",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"70",X"F8",X"FC",X"F8",X"70",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"70",X"F8",X"FC",X"F8",X"70",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"C6",X"20",X"90",X"40",X"20",X"80",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"06",X"70",X"80",X"30",X"C0",X"00",X"C0",X"00",X"00",X"00",X"00",
		X"3C",X"7E",X"F7",X"7E",X"3C",X"1C",X"3E",X"7F",X"F7",X"7E",X"3C",X"3C",X"7E",X"F7",X"7E",X"3C",
		X"28",X"7E",X"FE",X"37",X"EA",X"74",X"5F",X"6E",X"6E",X"5F",X"74",X"EA",X"37",X"FE",X"7E",X"14",
		X"00",X"00",X"18",X"18",X"34",X"52",X"34",X"4A",X"52",X"2C",X"4A",X"2C",X"18",X"18",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"38",X"30",X"28",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"0E",X"06",X"1E",X"1E",X"1E",X"08",X"0C",X"1A",X"16",X"0E",X"1E",X"1E",X"1C",X"0C",
		X"00",X"30",X"38",X"38",X"58",X"78",X"58",X"50",X"58",X"38",X"78",X"70",X"68",X"18",X"78",X"30",
		X"00",X"00",X"00",X"00",X"02",X"03",X"00",X"03",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"03",X"00",X"03",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"54",X"CB",X"50",X"A2",X"05",X"B2",X"4B",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"7E",X"7D",X"E6",X"63",X"67",X"FB",X"6E",X"2A",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"18",X"BC",X"7F",X"EF",X"7E",X"FD",X"14",X"A0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
