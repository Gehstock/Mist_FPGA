library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity guzzler_tile_bit2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of guzzler_tile_bit2 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7E",X"D8",X"8F",X"88",X"8F",X"88",X"DF",X"70",X"7F",X"DD",X"88",X"88",X"88",X"88",X"DD",X"77",
		X"FF",X"DD",X"88",X"88",X"88",X"88",X"DD",X"77",X"FE",X"D8",X"8F",X"88",X"8F",X"88",X"DF",X"70",
		X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"03",X"01",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"03",X"01",
		X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"03",X"01",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"03",X"01",
		X"04",X"26",X"73",X"31",X"6E",X"71",X"23",X"02",X"00",X"22",X"77",X"33",X"66",X"77",X"22",X"00",
		X"00",X"22",X"77",X"33",X"66",X"77",X"22",X"00",X"04",X"26",X"73",X"31",X"6E",X"71",X"23",X"02",
		X"00",X"00",X"00",X"07",X"07",X"E3",X"1C",X"F8",X"00",X"00",X"00",X"E0",X"90",X"90",X"F0",X"08",
		X"F7",X"37",X"7B",X"00",X"00",X"00",X"00",X"00",X"E8",X"90",X"90",X"F0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"EB",X"17",X"F7",X"00",X"00",X"00",X"00",X"F0",X"90",X"90",X"E8",
		X"F8",X"3C",X"73",X"07",X"07",X"00",X"00",X"00",X"08",X"F0",X"90",X"90",X"E0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"06",X"03",X"FF",X"3F",X"FF",X"00",X"00",X"00",X"00",X"C0",X"F0",X"F8",X"F8",
		X"FF",X"63",X"07",X"00",X"00",X"00",X"00",X"00",X"F0",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"81",X"81",X"81",X"81",X"81",X"81",X"FF",X"FF",X"FF",X"FF",X"81",X"81",X"81",X"81",X"81",X"81",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"03",X"1B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"01",X"03",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"06",X"07",X"23",X"33",X"31",X"19",X"00",X"00",X"08",X"8C",X"8E",X"CE",X"CE",X"E6",
		X"18",X"BC",X"EC",X"C8",X"E0",X"60",X"20",X"00",X"E6",X"F2",X"70",X"78",X"78",X"38",X"18",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3C",X"5A",X"99",X"BD",X"BD",X"99",X"42",X"3C",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"07",X"00",X"00",X"00",X"00",X"C0",X"C0",X"A0",X"80",
		X"03",X"01",X"00",X"02",X"01",X"00",X"00",X"00",X"C0",X"E0",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"06",X"05",X"0A",X"00",X"00",X"07",X"0C",X"13",X"14",X"2B",X"2A",
		X"0A",X"05",X"06",X"01",X"00",X"00",X"00",X"00",X"2A",X"2B",X"14",X"13",X"0C",X"03",X"00",X"00",
		X"00",X"00",X"03",X"04",X"03",X"00",X"03",X"04",X"00",X"00",X"E0",X"10",X"E0",X"00",X"E0",X"10",
		X"03",X"00",X"00",X"04",X"04",X"07",X"00",X"00",X"E0",X"00",X"60",X"90",X"90",X"A0",X"00",X"00",
		X"00",X"00",X"03",X"04",X"03",X"00",X"03",X"04",X"00",X"00",X"C0",X"20",X"C0",X"00",X"C0",X"20",
		X"03",X"00",X"02",X"05",X"05",X"02",X"00",X"00",X"C0",X"00",X"C0",X"20",X"20",X"C0",X"00",X"00",
		X"03",X"04",X"03",X"00",X"03",X"04",X"03",X"00",X"C0",X"20",X"C0",X"00",X"C0",X"20",X"C0",X"00",
		X"03",X"04",X"03",X"00",X"00",X"07",X"02",X"00",X"C0",X"20",X"C0",X"00",X"20",X"E0",X"20",X"00",
		X"03",X"04",X"03",X"00",X"03",X"04",X"03",X"00",X"C0",X"20",X"C0",X"00",X"C0",X"20",X"C0",X"00",
		X"03",X"04",X"03",X"00",X"03",X"04",X"04",X"02",X"C0",X"20",X"C0",X"00",X"20",X"A0",X"A0",X"60",
		X"03",X"04",X"03",X"00",X"03",X"04",X"03",X"00",X"C0",X"20",X"C0",X"00",X"C0",X"20",X"C0",X"00",
		X"03",X"04",X"03",X"00",X"06",X"05",X"05",X"04",X"C0",X"20",X"C0",X"00",X"C0",X"20",X"20",X"40",
		X"03",X"04",X"03",X"00",X"03",X"04",X"03",X"00",X"C0",X"20",X"C0",X"00",X"C0",X"20",X"C0",X"00",
		X"03",X"04",X"03",X"00",X"00",X"07",X"04",X"03",X"C0",X"20",X"C0",X"00",X"40",X"E0",X"40",X"C0",
		X"03",X"04",X"03",X"00",X"03",X"04",X"03",X"00",X"C0",X"20",X"C0",X"00",X"C0",X"20",X"C0",X"00",
		X"03",X"04",X"03",X"00",X"00",X"05",X"05",X"07",X"C0",X"20",X"C0",X"00",X"C0",X"20",X"20",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"06",X"05",X"05",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BF",X"73",X"61",X"40",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"04",X"07",X"13",X"17",
		X"80",X"C0",X"80",X"80",X"40",X"60",X"B1",X"DF",X"0D",X"09",X"08",X"04",X"04",X"04",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"08",X"1F",X"1E",X"00",X"00",X"00",X"00",X"40",X"CC",X"C5",X"E7",
		X"0C",X"0E",X"06",X"06",X"00",X"00",X"00",X"00",X"67",X"27",X"23",X"32",X"30",X"10",X"10",X"00",
		X"0C",X"0D",X"0F",X"0E",X"0C",X"0C",X"08",X"08",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"7F",X"C3",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",
		X"FF",X"D1",X"D1",X"91",X"95",X"95",X"B5",X"B5",X"FF",X"83",X"83",X"81",X"F9",X"F9",X"FD",X"FD",
		X"B5",X"BD",X"BD",X"99",X"81",X"C3",X"C3",X"FF",X"FD",X"FD",X"F9",X"F9",X"81",X"83",X"83",X"FF",
		X"FF",X"BD",X"BD",X"9D",X"9D",X"8D",X"8D",X"A5",X"FF",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",
		X"A5",X"B1",X"B1",X"B9",X"B9",X"BD",X"BD",X"FF",X"FD",X"FD",X"FD",X"FD",X"81",X"81",X"81",X"FF",
		X"FF",X"BD",X"BD",X"BD",X"BD",X"AD",X"AD",X"AD",X"FF",X"CD",X"CD",X"85",X"85",X"B1",X"B1",X"B1",
		X"AD",X"AD",X"AD",X"AD",X"81",X"81",X"81",X"FF",X"B7",X"B7",X"B7",X"B7",X"81",X"81",X"81",X"FF",
		X"5C",X"DD",X"DF",X"7E",X"3C",X"3C",X"18",X"18",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",
		X"50",X"D0",X"D0",X"70",X"30",X"30",X"10",X"10",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0C",X"00",X"04",X"05",X"05",X"05",X"05",X"05",X"05",
		X"00",X"00",X"00",X"00",X"40",X"40",X"44",X"5C",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"00",X"00",X"00",X"00",X"40",X"40",X"40",X"50",X"5C",X"00",X"00",X"00",X"00",X"00",X"00",X"5C",
		X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"3F",X"3F",X"3F",X"1F",X"0F",X"07",
		X"0F",X"67",X"CF",X"FF",X"FF",X"7F",X"3F",X"1F",X"3F",X"7F",X"7F",X"3F",X"3F",X"7F",X"7F",X"7F",
		X"1E",X"21",X"1E",X"00",X"1E",X"21",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"21",X"1E",X"00",X"06",X"29",X"29",X"3A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"1A",X"0F",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"05",X"05",X"05",X"00",X"08",X"0D",X"07",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"00",
		X"FF",X"FF",X"C1",X"01",X"03",X"03",X"07",X"07",X"FF",X"81",X"81",X"81",X"81",X"81",X"81",X"FF",
		X"C3",X"C3",X"C3",X"C3",X"CB",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5D",X"5F",X"5F",X"5F",X"7F",X"7F",X"7F",X"5F",X"5F",X"5F",
		X"5F",X"7F",X"DF",X"FF",X"FF",X"7F",X"7F",X"5F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"00",X"00",X"1E",X"21",X"1E",X"00",X"1E",X"21",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"00",X"19",X"25",X"25",X"13",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"1E",X"21",X"1E",X"00",X"1E",X"21",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"00",X"06",X"29",X"29",X"3A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"1E",X"21",X"1E",X"00",X"1E",X"21",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"00",X"16",X"29",X"29",X"16",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"21",X"1E",X"00",X"1E",X"21",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"21",X"1E",X"00",X"01",X"3F",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"21",X"1E",X"00",X"1E",X"21",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"21",X"1E",X"00",X"19",X"25",X"25",X"13",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"21",X"1E",X"00",X"1E",X"21",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"21",X"1E",X"00",X"36",X"29",X"29",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"21",X"1E",X"00",X"1E",X"21",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"21",X"1E",X"00",X"02",X"3F",X"22",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"F3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"07",X"07",X"03",X"03",X"03",X"01",X"07",X"07",X"07",X"3F",X"3F",X"3F",X"1F",X"0F",X"07",
		X"0F",X"67",X"CF",X"FF",X"FF",X"7F",X"3F",X"1F",X"3F",X"7F",X"7F",X"3F",X"3F",X"7F",X"7F",X"7F",
		X"5F",X"07",X"07",X"03",X"03",X"03",X"01",X"5F",X"5F",X"07",X"3F",X"3F",X"3F",X"1F",X"0F",X"5F",
		X"5F",X"67",X"CF",X"FF",X"FF",X"7F",X"3F",X"5F",X"7F",X"7F",X"7F",X"3F",X"3F",X"7F",X"7F",X"7F",
		X"00",X"00",X"00",X"30",X"38",X"3C",X"3C",X"3E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3C",X"3C",X"38",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"30",X"78",X"70",X"3A",X"7A",X"7A",X"FA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FA",X"7A",X"3A",X"70",X"70",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"0C",X"18",X"00",X"07",X"18",X"20",X"07",X"E0",X"30",X"18",X"00",X"E0",X"18",X"04",X"E0",
		X"18",X"20",X"00",X"0F",X"1F",X"1F",X"0F",X"07",X"18",X"04",X"00",X"F0",X"F8",X"F8",X"F0",X"E0",
		X"00",X"00",X"00",X"01",X"03",X"03",X"07",X"3C",X"00",X"00",X"00",X"F0",X"FC",X"FF",X"FF",X"FF",
		X"38",X"00",X"00",X"03",X"01",X"00",X"00",X"00",X"7F",X"7F",X"FF",X"FC",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"3F",X"1F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"0F",X"19",X"03",X"02",X"00",X"00",X"00",
		X"00",X"00",X"03",X"04",X"03",X"00",X"03",X"04",X"00",X"00",X"C0",X"20",X"C0",X"00",X"C0",X"20",
		X"03",X"00",X"03",X"04",X"04",X"02",X"00",X"00",X"C0",X"00",X"20",X"A0",X"A0",X"60",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"0F",X"1F",X"3E",X"7C",X"7C",X"7F",X"7F",X"40",X"E0",X"F0",X"3E",X"7E",X"FE",X"FE",X"F2",
		X"7C",X"3B",X"7B",X"7C",X"3B",X"0C",X"00",X"00",X"30",X"DC",X"DC",X"3C",X"DC",X"18",X"18",X"00",
		X"00",X"0F",X"1F",X"3E",X"7C",X"7C",X"7F",X"7F",X"00",X"E0",X"70",X"78",X"70",X"FE",X"FE",X"FE",
		X"7C",X"38",X"78",X"7C",X"38",X"0C",X"00",X"00",X"3E",X"D2",X"D0",X"30",X"C0",X"20",X"00",X"00",
		X"00",X"0F",X"1F",X"3E",X"7C",X"7C",X"7F",X"7F",X"00",X"E0",X"FC",X"3C",X"1C",X"9C",X"F4",X"F0",
		X"7C",X"3B",X"7B",X"7C",X"3B",X"0C",X"00",X"00",X"7E",X"DE",X"DE",X"3E",X"D2",X"20",X"00",X"00",
		X"00",X"04",X"1C",X"3F",X"38",X"77",X"77",X"38",X"30",X"30",X"F8",X"F8",X"78",X"B8",X"B8",X"70",
		X"38",X"77",X"77",X"39",X"3F",X"1C",X"04",X"00",X"70",X"BE",X"FE",X"FE",X"3E",X"32",X"20",X"00",
		X"00",X"04",X"1C",X"3F",X"39",X"71",X"71",X"38",X"00",X"20",X"32",X"3E",X"FE",X"FE",X"BE",X"70",
		X"38",X"71",X"71",X"38",X"3F",X"1C",X"04",X"00",X"70",X"B8",X"B8",X"78",X"F8",X"F8",X"30",X"30",
		X"01",X"0F",X"1F",X"3E",X"7C",X"7C",X"7F",X"7F",X"40",X"C0",X"C0",X"06",X"06",X"06",X"06",X"02",
		X"7C",X"3B",X"7B",X"7C",X"3B",X"0C",X"00",X"00",X"00",X"CC",X"CC",X"0C",X"DC",X"18",X"18",X"00",
		X"00",X"0F",X"1F",X"3E",X"7C",X"7C",X"7F",X"7F",X"00",X"20",X"70",X"78",X"20",X"06",X"06",X"06",
		X"7C",X"38",X"78",X"7C",X"38",X"0C",X"00",X"00",X"06",X"C2",X"C0",X"00",X"C0",X"00",X"00",X"00",
		X"00",X"0F",X"1F",X"3E",X"7C",X"7C",X"7F",X"7F",X"00",X"00",X"0C",X"0C",X"0C",X"0C",X"E4",X"60",
		X"7C",X"3B",X"7B",X"7C",X"3B",X"0C",X"00",X"00",X"46",X"C6",X"C6",X"06",X"C2",X"00",X"00",X"00",
		X"02",X"0F",X"1F",X"3C",X"7C",X"7C",X"7F",X"7F",X"BE",X"BC",X"80",X"00",X"00",X"00",X"00",X"00",
		X"7C",X"3B",X"7B",X"7C",X"7B",X"3C",X"37",X"77",X"00",X"C6",X"C6",X"06",X"C6",X"1A",X"B8",X"B8",
		X"00",X"04",X"1C",X"3F",X"38",X"77",X"77",X"38",X"30",X"30",X"28",X"98",X"18",X"98",X"98",X"00",
		X"38",X"77",X"77",X"39",X"3F",X"1C",X"04",X"00",X"00",X"86",X"C6",X"C6",X"06",X"02",X"00",X"00",
		X"00",X"04",X"1C",X"3F",X"38",X"77",X"F7",X"F8",X"30",X"30",X"22",X"86",X"06",X"86",X"86",X"00",
		X"F8",X"F7",X"77",X"38",X"3F",X"1C",X"04",X"00",X"00",X"86",X"86",X"06",X"86",X"A2",X"30",X"30",
		X"00",X"04",X"1C",X"3F",X"39",X"71",X"71",X"38",X"00",X"00",X"02",X"06",X"C6",X"C6",X"86",X"00",
		X"38",X"71",X"71",X"38",X"3F",X"1C",X"04",X"00",X"00",X"98",X"98",X"18",X"98",X"A8",X"30",X"30",
		X"00",X"04",X"1C",X"3F",X"38",X"77",X"77",X"38",X"30",X"30",X"23",X"87",X"07",X"86",X"87",X"0F",
		X"38",X"77",X"77",X"38",X"3F",X"1C",X"04",X"00",X"0F",X"87",X"86",X"07",X"87",X"A3",X"30",X"30",
		X"01",X"0B",X"19",X"38",X"78",X"78",X"78",X"78",X"40",X"C0",X"C0",X"06",X"06",X"06",X"06",X"02",
		X"78",X"30",X"6E",X"6E",X"30",X"0E",X"00",X"00",X"00",X"0C",X"0C",X"0C",X"1C",X"18",X"18",X"00",
		X"00",X"08",X"18",X"38",X"78",X"78",X"78",X"78",X"00",X"20",X"70",X"78",X"20",X"06",X"06",X"06",
		X"78",X"30",X"66",X"66",X"30",X"06",X"00",X"00",X"06",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"18",X"38",X"78",X"78",X"78",X"78",X"00",X"00",X"0C",X"0C",X"0C",X"0C",X"E4",X"60",
		X"78",X"30",X"6E",X"6E",X"30",X"0E",X"00",X"00",X"46",X"06",X"06",X"06",X"02",X"00",X"00",X"00",
		X"02",X"0F",X"1B",X"38",X"78",X"78",X"78",X"78",X"BE",X"BC",X"80",X"00",X"00",X"00",X"00",X"00",
		X"78",X"30",X"6E",X"6E",X"70",X"2E",X"31",X"77",X"80",X"86",X"86",X"86",X"86",X"BA",X"B8",X"B8",
		X"00",X"00",X"18",X"38",X"38",X"76",X"76",X"38",X"30",X"30",X"28",X"18",X"98",X"98",X"98",X"80",
		X"38",X"76",X"76",X"38",X"39",X"18",X"00",X"00",X"80",X"86",X"A6",X"E6",X"E6",X"02",X"00",X"00",
		X"00",X"00",X"18",X"38",X"30",X"6E",X"EE",X"F0",X"30",X"30",X"22",X"06",X"C6",X"C6",X"C6",X"C0",
		X"F0",X"EE",X"6E",X"30",X"38",X"18",X"00",X"00",X"C0",X"C6",X"C6",X"C6",X"06",X"22",X"30",X"30",
		X"00",X"00",X"18",X"39",X"30",X"6E",X"6E",X"30",X"00",X"00",X"02",X"E6",X"E6",X"E6",X"C6",X"C0",
		X"30",X"6E",X"6E",X"30",X"38",X"18",X"00",X"00",X"C0",X"CC",X"CC",X"CC",X"0C",X"24",X"30",X"30",
		X"00",X"00",X"18",X"38",X"30",X"6E",X"6E",X"30",X"30",X"30",X"23",X"07",X"C7",X"C6",X"C7",X"C7",
		X"30",X"6E",X"6E",X"30",X"38",X"18",X"00",X"00",X"C7",X"C7",X"C6",X"C7",X"07",X"23",X"30",X"30",
		X"01",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"40",X"C0",X"C0",X"06",X"06",X"06",X"06",X"02",
		X"00",X"00",X"0E",X"0E",X"00",X"0E",X"00",X"00",X"00",X"0C",X"0C",X"0C",X"1C",X"18",X"18",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"70",X"78",X"20",X"06",X"06",X"06",
		X"00",X"00",X"06",X"06",X"00",X"06",X"00",X"00",X"06",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0C",X"0C",X"0C",X"E4",X"60",
		X"00",X"00",X"0E",X"0E",X"00",X"0E",X"00",X"00",X"46",X"06",X"06",X"06",X"02",X"00",X"00",X"00",
		X"02",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"BE",X"BC",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0E",X"0E",X"40",X"2E",X"31",X"77",X"80",X"86",X"86",X"86",X"86",X"9A",X"B8",X"B8",
		X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"30",X"30",X"28",X"18",X"98",X"98",X"98",X"80",
		X"00",X"06",X"06",X"00",X"01",X"00",X"00",X"00",X"80",X"86",X"A6",X"E6",X"E6",X"02",X"00",X"00",
		X"00",X"80",X"00",X"00",X"00",X"0E",X"8E",X"C0",X"30",X"30",X"22",X"06",X"C6",X"C6",X"C6",X"C0",
		X"C0",X"8E",X"0E",X"00",X"00",X"00",X"80",X"00",X"C0",X"C6",X"C6",X"C6",X"06",X"22",X"30",X"30",
		X"00",X"00",X"00",X"01",X"00",X"0E",X"0E",X"00",X"00",X"00",X"02",X"E6",X"E6",X"E6",X"C6",X"C0",
		X"00",X"0E",X"0E",X"00",X"00",X"00",X"00",X"00",X"C0",X"CC",X"CC",X"CC",X"0C",X"24",X"30",X"30",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"0E",X"00",X"30",X"30",X"23",X"07",X"C7",X"C6",X"C7",X"C7",
		X"00",X"0E",X"0E",X"00",X"00",X"00",X"00",X"00",X"C7",X"C7",X"C6",X"C7",X"07",X"23",X"30",X"30",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"B8",X"B8",X"B8",X"B8",X"B8",X"B8",X"B8",X"B8",
		X"77",X"77",X"77",X"23",X"00",X"00",X"00",X"00",X"B8",X"B8",X"B8",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"54",X"77",X"23",X"00",X"00",X"00",X"00",X"00",X"A8",X"B8",X"10",X"00",X"00",X"00",X"00",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"B8",X"B8",X"B8",X"B8",X"B8",X"B8",X"B8",X"B8",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"B8",X"B8",X"B8",X"B8",X"B8",X"B8",X"B8",X"B8",
		X"00",X"00",X"00",X"00",X"77",X"77",X"77",X"77",X"00",X"00",X"00",X"00",X"B8",X"B8",X"B8",X"B8",
		X"77",X"77",X"77",X"23",X"00",X"00",X"00",X"00",X"B8",X"B8",X"B8",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"77",X"77",X"23",X"00",X"00",X"00",X"00",X"B8",X"B8",X"B8",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"54",X"77",X"77",X"77",X"77",X"77",X"77",X"00",X"A8",X"B8",X"B8",X"B8",X"B8",X"B8",X"B8",
		X"00",X"07",X"0F",X"07",X"00",X"07",X"0F",X"0F",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",
		X"07",X"00",X"07",X"0F",X"07",X"00",X"00",X"00",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"00",X"06",X"0C",X"06",X"00",X"06",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"00",X"06",X"0C",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",
		X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"00",X"07",X"0F",X"07",X"00",X"07",X"0F",X"0F",X"00",X"F0",X"F0",X"F0",X"00",X"F0",X"F0",X"F0",
		X"07",X"00",X"07",X"0F",X"07",X"00",X"00",X"00",X"F0",X"00",X"F0",X"F0",X"F0",X"00",X"00",X"00",
		X"00",X"07",X"0F",X"07",X"00",X"07",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"00",X"07",X"0F",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FE",X"FC",X"FE",X"00",X"FE",X"FC",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"00",X"FE",X"FC",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"1E",X"1C",X"18",X"0F",X"00",X"00",X"00",X"1C",X"3C",X"38",X"10",X"0F",X"18",X"1C",X"0E",
		X"0C",X"0E",X"06",X"03",X"CF",X"06",X"0E",X"0C",X"04",X"66",X"73",X"31",X"6E",X"71",X"23",X"02",
		X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"FE",X"00",X"00",X"00",X"00",X"00",X"FF",X"C3",X"7C",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"6C",X"74",X"7C",X"60",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"03",X"02",X"05",X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"BD",
		X"03",X"1F",X"1F",X"07",X"03",X"03",X"01",X"00",X"DD",X"ED",X"DD",X"BD",X"DD",X"ED",X"FF",X"00",
		X"00",X"00",X"00",X"01",X"7F",X"7F",X"1E",X"3C",X"00",X"00",X"00",X"F8",X"FC",X"FC",X"7E",X"3E",
		X"7C",X"1E",X"7E",X"CF",X"1F",X"3F",X"03",X"07",X"3E",X"1C",X"18",X"38",X"F8",X"F0",X"C0",X"00",
		X"00",X"01",X"1C",X"3C",X"3C",X"78",X"71",X"7F",X"00",X"80",X"E0",X"F0",X"F8",X"F8",X"FC",X"FC",
		X"7F",X"3F",X"1B",X"11",X"00",X"00",X"00",X"00",X"FC",X"FC",X"F8",X"78",X"30",X"20",X"00",X"00",
		X"00",X"00",X"19",X"39",X"39",X"78",X"7C",X"7F",X"00",X"80",X"C0",X"C0",X"C8",X"DC",X"7C",X"FC",
		X"7F",X"3F",X"3F",X"15",X"00",X"00",X"00",X"00",X"FC",X"F8",X"F8",X"50",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0E",X"1E",X"3E",X"3C",X"71",X"7F",X"00",X"C0",X"60",X"60",X"60",X"E4",X"CC",X"9C",
		X"7F",X"7F",X"3F",X"3D",X"18",X"08",X"00",X"00",X"FC",X"F8",X"B0",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"00",X"03",X"0F",X"07",X"00",X"00",X"F0",X"F8",X"30",X"18",X"88",X"C8",
		X"0F",X"3F",X"3F",X"1E",X"07",X"01",X"00",X"00",X"C8",X"88",X"18",X"30",X"F8",X"F0",X"00",X"00",
		X"00",X"00",X"01",X"07",X"1E",X"3F",X"3F",X"0F",X"00",X"00",X"F0",X"F8",X"7C",X"3C",X"9E",X"DE",
		X"07",X"0F",X"03",X"00",X"03",X"00",X"00",X"00",X"DE",X"9E",X"3C",X"7C",X"F8",X"F0",X"00",X"00",
		X"01",X"00",X"00",X"1C",X"3C",X"79",X"E3",X"FF",X"C0",X"C0",X"C0",X"E0",X"F0",X"F0",X"F8",X"F8",
		X"FF",X"BF",X"3F",X"7F",X"5F",X"10",X"00",X"00",X"F8",X"F8",X"F0",X"E0",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"1C",X"3C",X"38",X"71",X"77",X"00",X"00",X"C0",X"E0",X"F0",X"F8",X"F8",X"F8",
		X"FF",X"DF",X"9F",X"3F",X"67",X"4C",X"08",X"00",X"F8",X"F8",X"F8",X"F0",X"E0",X"00",X"00",X"00",
		X"00",X"00",X"04",X"1C",X"38",X"71",X"F7",X"FF",X"00",X"00",X"E0",X"E0",X"F0",X"F0",X"F8",X"F8",
		X"9F",X"3F",X"7F",X"4F",X"0B",X"01",X"00",X"00",X"F8",X"F8",X"F8",X"F0",X"E0",X"80",X"C0",X"00",
		X"00",X"00",X"00",X"03",X"0F",X"04",X"3E",X"9F",X"18",X"38",X"70",X"F0",X"F8",X"78",X"3C",X"3C",
		X"FF",X"FF",X"7E",X"7C",X"3F",X"0F",X"00",X"00",X"3C",X"3C",X"3C",X"78",X"F8",X"F0",X"70",X"00",
		X"00",X"00",X"0F",X"1F",X"3C",X"7E",X"3F",X"FF",X"00",X"70",X"F0",X"F8",X"78",X"3C",X"3C",X"3C",
		X"7F",X"3E",X"7C",X"0F",X"03",X"00",X"00",X"00",X"3C",X"3C",X"78",X"F8",X"F0",X"70",X"38",X"18",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"38",X"1C",X"0E",X"DE",X"DC",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"DC",X"DE",X"0E",X"1C",X"38",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"3C",X"0E",X"06",X"0A",X"0A",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0A",X"0A",X"06",X"0E",X"3C",X"38",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"C8",X"C8",X"F8",X"70",X"00",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C8",X"C8",X"F8",X"70",X"00",X"00",X"00",X"00",
		X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"C0",X"90",X"00",X"78",X"00",
		X"00",X"00",X"01",X"03",X"00",X"00",X"00",X"00",X"10",X"C0",X"E0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"06",X"0C",X"30",X"00",X"00",X"00",X"F8",X"0C",X"02",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3E",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"7F",X"7C",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"7F",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"3E",X"FE",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"7C",
		X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"60",X"60",X"70",X"30",X"3C",X"1F",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"07",X"1F",X"3C",X"30",X"70",X"60",X"60",X"10",X"00",X"00",X"00",X"80",X"C0",X"71",X"10",
		X"10",X"00",X"00",X"00",X"00",X"00",X"F1",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
