library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity sound_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of sound_rom is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"86",X"FF",X"1F",X"8A",X"8E",X"00",X"00",X"CC",X"00",X"00",X"ED",X"81",X"8C",X"07",X"FF",X"23",
		X"F9",X"10",X"CE",X"08",X"00",X"BD",X"E0",X"76",X"1C",X"AF",X"20",X"FE",X"34",X"FF",X"0C",X"00",
		X"BD",X"E0",X"2F",X"BD",X"E1",X"3F",X"BD",X"F2",X"5D",X"BD",X"E0",X"40",X"35",X"FF",X"3B",X"96",
		X"01",X"26",X"01",X"39",X"0F",X"01",X"CE",X"E6",X"78",X"96",X"02",X"84",X"1F",X"48",X"6E",X"D6",
		X"5F",X"CE",X"01",X"00",X"4F",X"74",X"01",X"1A",X"49",X"74",X"01",X"19",X"49",X"74",X"01",X"18",
		X"49",X"74",X"01",X"14",X"49",X"74",X"01",X"13",X"49",X"74",X"01",X"12",X"49",X"8B",X"C0",X"C6",
		X"07",X"F7",X"20",X"00",X"B7",X"20",X"01",X"39",X"34",X"7E",X"B6",X"A0",X"00",X"97",X"02",X"86",
		X"FF",X"97",X"01",X"35",X"7E",X"3B",X"CE",X"02",X"00",X"86",X"20",X"C6",X"1B",X"6F",X"C4",X"33",
		X"C6",X"5A",X"26",X"F9",X"39",X"0B",X"3C",X"0A",X"9B",X"0A",X"02",X"09",X"73",X"08",X"EB",X"08",
		X"6B",X"07",X"F2",X"07",X"80",X"07",X"14",X"06",X"AE",X"06",X"4E",X"05",X"F4",X"05",X"9E",X"05",
		X"4D",X"05",X"01",X"04",X"B9",X"04",X"75",X"04",X"35",X"03",X"F9",X"03",X"C0",X"03",X"8A",X"03",
		X"57",X"03",X"27",X"02",X"FA",X"02",X"CF",X"02",X"A7",X"02",X"81",X"02",X"5D",X"02",X"3B",X"02",
		X"1B",X"01",X"FC",X"01",X"E0",X"01",X"C5",X"01",X"A5",X"01",X"94",X"01",X"7D",X"01",X"68",X"01",
		X"53",X"01",X"40",X"01",X"2E",X"01",X"1D",X"01",X"0D",X"00",X"FE",X"00",X"F0",X"00",X"E2",X"00",
		X"D6",X"00",X"CA",X"00",X"BE",X"00",X"B4",X"00",X"AA",X"00",X"A0",X"00",X"97",X"00",X"8F",X"00",
		X"87",X"00",X"7F",X"00",X"78",X"00",X"71",X"00",X"6B",X"00",X"65",X"00",X"5F",X"00",X"5A",X"00",
		X"55",X"00",X"50",X"00",X"4C",X"00",X"47",X"00",X"43",X"00",X"40",X"00",X"3C",X"00",X"39",X"00",
		X"35",X"00",X"32",X"00",X"30",X"00",X"2D",X"00",X"2A",X"00",X"28",X"00",X"26",X"00",X"24",X"00",
		X"22",X"00",X"20",X"00",X"1E",X"00",X"1C",X"00",X"1B",X"00",X"19",X"00",X"18",X"00",X"16",X"00",
		X"15",X"00",X"14",X"00",X"13",X"00",X"12",X"00",X"11",X"00",X"10",X"00",X"0F",X"00",X"0E",X"BD",
		X"E1",X"46",X"BD",X"E1",X"6B",X"39",X"8E",X"02",X"00",X"0F",X"0F",X"0F",X"04",X"A6",X"84",X"27",
		X"0B",X"9B",X"0F",X"BD",X"E1",X"9E",X"96",X"0F",X"81",X"03",X"24",X"0E",X"0C",X"04",X"96",X"04",
		X"81",X"0F",X"27",X"06",X"86",X"20",X"30",X"86",X"20",X"E3",X"39",X"8E",X"04",X"60",X"C6",X"60",
		X"A6",X"84",X"26",X"08",X"8E",X"04",X"00",X"A6",X"84",X"26",X"12",X"39",X"BD",X"EE",X"5B",X"86",
		X"20",X"30",X"86",X"BD",X"EE",X"5B",X"86",X"20",X"30",X"86",X"7E",X"EE",X"5B",X"BD",X"EE",X"5B",
		X"86",X"20",X"30",X"86",X"BD",X"EE",X"5B",X"86",X"20",X"30",X"86",X"7E",X"EE",X"60",X"CE",X"E1",
		X"A6",X"96",X"04",X"48",X"6E",X"D6",X"E1",X"C4",X"E2",X"07",X"E2",X"2F",X"E2",X"E5",X"E3",X"BC",
		X"E3",X"BD",X"E4",X"24",X"E4",X"75",X"E4",X"88",X"E4",X"C6",X"E4",X"FB",X"E5",X"2F",X"E5",X"C6",
		X"E5",X"C7",X"E6",X"10",X"6A",X"0D",X"27",X"1B",X"A6",X"0D",X"44",X"CE",X"E1",X"D3",X"A6",X"C6",
		X"A7",X"07",X"39",X"01",X"02",X"03",X"05",X"07",X"09",X"0A",X"0B",X"0C",X"0D",X"0D",X"0D",X"0C",
		X"0A",X"08",X"06",X"A6",X"0C",X"6C",X"0C",X"81",X"05",X"27",X"19",X"CE",X"E1",X"FF",X"A6",X"C6",
		X"CE",X"E0",X"E5",X"48",X"EC",X"C6",X"A7",X"02",X"E7",X"01",X"86",X"1F",X"A7",X"0D",X"39",X"07",
		X"0C",X"10",X"13",X"13",X"6F",X"84",X"39",X"6A",X"0D",X"27",X"01",X"39",X"6C",X"0C",X"A6",X"0C",
		X"81",X"03",X"27",X"18",X"C6",X"3C",X"E7",X"0D",X"81",X"01",X"27",X"08",X"CC",X"00",X"26",X"A7",
		X"02",X"E7",X"01",X"39",X"CC",X"00",X"2A",X"A7",X"02",X"E7",X"01",X"39",X"6F",X"84",X"39",X"A6",
		X"88",X"12",X"26",X"45",X"6A",X"88",X"13",X"27",X"01",X"39",X"6C",X"88",X"12",X"CC",X"00",X"18",
		X"A7",X"02",X"E7",X"01",X"CC",X"00",X"20",X"A7",X"04",X"E7",X"03",X"CC",X"00",X"28",X"A7",X"06",
		X"E7",X"05",X"86",X"00",X"A7",X"0C",X"86",X"0F",X"A7",X"0D",X"86",X"07",X"A7",X"07",X"86",X"01",
		X"A7",X"0E",X"86",X"10",X"A7",X"0F",X"86",X"03",X"A7",X"08",X"86",X"01",X"A7",X"88",X"10",X"86",
		X"10",X"A7",X"88",X"11",X"86",X"0D",X"A7",X"09",X"39",X"BD",X"E2",X"83",X"BD",X"E2",X"A1",X"BD",
		X"E2",X"BF",X"39",X"A6",X"0C",X"84",X"01",X"27",X"0C",X"6A",X"07",X"27",X"01",X"39",X"6A",X"0D",
		X"27",X"50",X"6C",X"0C",X"39",X"6C",X"07",X"A6",X"07",X"A1",X"0D",X"27",X"01",X"39",X"6C",X"0C",
		X"39",X"A6",X"0E",X"84",X"01",X"27",X"0C",X"6A",X"08",X"27",X"01",X"39",X"6A",X"0F",X"27",X"32",
		X"6C",X"0E",X"39",X"6C",X"08",X"A6",X"08",X"A1",X"0F",X"27",X"01",X"39",X"6C",X"0E",X"39",X"A6",
		X"88",X"10",X"84",X"01",X"27",X"0E",X"6A",X"09",X"27",X"01",X"39",X"6A",X"88",X"11",X"27",X"12",
		X"6C",X"88",X"10",X"39",X"6C",X"09",X"A6",X"09",X"A1",X"88",X"11",X"27",X"01",X"39",X"6C",X"88",
		X"10",X"39",X"6F",X"84",X"39",X"A6",X"0D",X"27",X"03",X"6A",X"0D",X"39",X"A6",X"88",X"10",X"6C",
		X"88",X"10",X"81",X"10",X"27",X"21",X"E6",X"0F",X"E7",X"0D",X"CE",X"E3",X"06",X"A6",X"C6",X"A7",
		X"07",X"A7",X"08",X"A7",X"09",X"39",X"09",X"0A",X"0B",X"0C",X"0D",X"0C",X"0B",X"0A",X"09",X"08",
		X"07",X"06",X"05",X"04",X"03",X"02",X"01",X"6F",X"88",X"10",X"A6",X"0C",X"6C",X"0C",X"48",X"48",
		X"CE",X"E3",X"88",X"33",X"C6",X"A6",X"C4",X"81",X"FF",X"27",X"5A",X"A7",X"0F",X"A7",X"0D",X"86",
		X"09",X"A7",X"07",X"A7",X"08",X"A7",X"09",X"A6",X"41",X"BD",X"E3",X"53",X"A7",X"02",X"E7",X"01",
		X"A6",X"42",X"BD",X"E3",X"53",X"A7",X"04",X"E7",X"03",X"A6",X"43",X"BD",X"E3",X"53",X"A7",X"06",
		X"E7",X"05",X"39",X"10",X"8E",X"E3",X"5F",X"48",X"31",X"A6",X"A6",X"A4",X"E6",X"21",X"39",X"00",
		X"00",X"00",X"D6",X"00",X"CA",X"00",X"BE",X"00",X"B4",X"00",X"AA",X"00",X"A0",X"00",X"97",X"00",
		X"8F",X"00",X"87",X"00",X"7F",X"00",X"78",X"00",X"71",X"00",X"6B",X"00",X"65",X"00",X"5F",X"00",
		X"5A",X"00",X"55",X"00",X"50",X"6F",X"84",X"39",X"04",X"01",X"05",X"08",X"02",X"00",X"00",X"00",
		X"02",X"01",X"05",X"08",X"02",X"01",X"05",X"08",X"02",X"01",X"05",X"08",X"02",X"03",X"06",X"0A",
		X"02",X"00",X"00",X"00",X"02",X"03",X"06",X"0A",X"02",X"00",X"00",X"00",X"02",X"03",X"06",X"0C",
		X"02",X"00",X"00",X"00",X"0C",X"05",X"08",X"0D",X"FF",X"FF",X"FF",X"FF",X"39",X"A6",X"0D",X"27",
		X"2E",X"6A",X"0D",X"A6",X"0E",X"27",X"0D",X"81",X"02",X"27",X"15",X"A6",X"0D",X"81",X"20",X"27",
		X"00",X"6C",X"0E",X"39",X"6C",X"07",X"A6",X"07",X"81",X"0D",X"27",X"01",X"39",X"6C",X"0E",X"39",
		X"A6",X"07",X"27",X"0A",X"96",X"00",X"84",X"03",X"27",X"01",X"39",X"6A",X"07",X"39",X"39",X"6F",
		X"0E",X"C6",X"30",X"A6",X"0C",X"6C",X"0C",X"CE",X"E4",X"18",X"A6",X"C6",X"81",X"FF",X"27",X"15",
		X"48",X"24",X"02",X"C6",X"90",X"E7",X"0D",X"CE",X"E0",X"9D",X"EC",X"C6",X"A7",X"02",X"E7",X"01",
		X"86",X"06",X"A7",X"07",X"39",X"6F",X"84",X"39",X"18",X"97",X"18",X"9A",X"15",X"91",X"0E",X"8C",
		X"09",X"85",X"02",X"FF",X"A6",X"0D",X"6C",X"0D",X"CE",X"E4",X"4C",X"A6",X"C6",X"81",X"FF",X"27",
		X"18",X"81",X"FE",X"26",X"07",X"86",X"42",X"A7",X"01",X"8B",X"08",X"39",X"A7",X"07",X"96",X"00",
		X"84",X"01",X"27",X"04",X"6A",X"01",X"6A",X"03",X"39",X"6F",X"84",X"39",X"04",X"05",X"06",X"07",
		X"08",X"09",X"08",X"07",X"06",X"05",X"04",X"03",X"02",X"01",X"FE",X"03",X"04",X"05",X"06",X"07",
		X"08",X"07",X"06",X"05",X"04",X"03",X"04",X"05",X"06",X"07",X"08",X"09",X"08",X"07",X"06",X"05",
		X"04",X"03",X"02",X"01",X"FF",X"E6",X"01",X"A6",X"02",X"83",X"00",X"1E",X"81",X"F0",X"24",X"05",
		X"A7",X"02",X"E7",X"01",X"39",X"6F",X"84",X"39",X"A6",X"0C",X"27",X"1E",X"81",X"02",X"27",X"0C",
		X"6A",X"0D",X"27",X"01",X"39",X"6C",X"0C",X"86",X"10",X"A7",X"0E",X"39",X"6A",X"0E",X"27",X"01",
		X"39",X"6A",X"07",X"27",X"1E",X"86",X"0E",X"A7",X"0E",X"39",X"6C",X"0E",X"A6",X"0E",X"84",X"01",
		X"27",X"01",X"39",X"6C",X"07",X"A6",X"07",X"81",X"0B",X"27",X"01",X"39",X"6C",X"0C",X"86",X"48",
		X"A7",X"0D",X"39",X"6F",X"84",X"39",X"A6",X"0D",X"27",X"09",X"6A",X"0D",X"A6",X"0E",X"A7",X"07",
		X"A7",X"08",X"39",X"A6",X"0C",X"27",X"10",X"6A",X"0E",X"A6",X"0E",X"81",X"02",X"27",X"05",X"86",
		X"05",X"A7",X"0D",X"39",X"6F",X"84",X"39",X"6C",X"0E",X"A6",X"0E",X"81",X"0A",X"27",X"05",X"86",
		X"02",X"A7",X"0D",X"39",X"6C",X"0C",X"86",X"05",X"A7",X"0D",X"39",X"A6",X"0D",X"27",X"12",X"6A",
		X"0D",X"CE",X"E5",X"09",X"A6",X"C6",X"A7",X"07",X"39",X"0B",X"0B",X"0C",X"0C",X"0D",X"0B",X"09",
		X"06",X"E6",X"01",X"5A",X"6C",X"0C",X"A6",X"0C",X"84",X"01",X"27",X"01",X"5A",X"A6",X"0C",X"84",
		X"03",X"26",X"02",X"6A",X"07",X"E7",X"01",X"C1",X"80",X"23",X"01",X"39",X"6F",X"84",X"39",X"96",
		X"00",X"84",X"01",X"27",X"F9",X"6A",X"0D",X"27",X"1A",X"A6",X"0D",X"CE",X"E5",X"43",X"A6",X"C6",
		X"A7",X"07",X"39",X"03",X"04",X"05",X"06",X"07",X"08",X"09",X"09",X"0A",X"0A",X"09",X"09",X"08",
		X"08",X"07",X"06",X"A6",X"0C",X"6C",X"0C",X"81",X"0C",X"27",X"14",X"CE",X"E5",X"BA",X"A6",X"C6",
		X"CE",X"E5",X"8A",X"48",X"EC",X"C6",X"A7",X"02",X"E7",X"01",X"86",X"0C",X"A7",X"0D",X"39",X"6F",
		X"84",X"39",X"03",X"57",X"03",X"27",X"02",X"FA",X"02",X"CF",X"02",X"A7",X"02",X"81",X"02",X"5D",
		X"02",X"3B",X"02",X"1B",X"01",X"FC",X"01",X"E0",X"01",X"C5",X"01",X"A5",X"01",X"94",X"01",X"7D",
		X"01",X"68",X"01",X"53",X"01",X"40",X"01",X"2E",X"01",X"1D",X"01",X"0D",X"00",X"FE",X"00",X"F0",
		X"00",X"E2",X"00",X"D6",X"00",X"CA",X"00",X"BE",X"00",X"B4",X"00",X"AA",X"00",X"A0",X"00",X"97",
		X"00",X"8F",X"00",X"87",X"00",X"7F",X"00",X"78",X"00",X"71",X"00",X"02",X"04",X"05",X"00",X"02",
		X"04",X"05",X"00",X"02",X"04",X"05",X"39",X"A6",X"0D",X"6C",X"0D",X"CE",X"E5",X"EC",X"A6",X"C6",
		X"81",X"FF",X"27",X"03",X"A7",X"07",X"39",X"6C",X"0C",X"A6",X"0C",X"81",X"05",X"27",X"2E",X"C6",
		X"2E",X"85",X"01",X"26",X"02",X"C6",X"34",X"E7",X"01",X"6F",X"0D",X"39",X"04",X"05",X"06",X"07",
		X"08",X"09",X"0A",X"0B",X"0C",X"0D",X"0E",X"0F",X"0F",X"0E",X"0D",X"0C",X"0B",X"0A",X"09",X"09",
		X"08",X"08",X"07",X"07",X"06",X"06",X"05",X"04",X"03",X"02",X"01",X"00",X"FF",X"6F",X"84",X"39",
		X"A6",X"0D",X"27",X"38",X"6A",X"0D",X"A6",X"0E",X"27",X"20",X"81",X"02",X"27",X"0E",X"A6",X"0D",
		X"81",X"20",X"23",X"01",X"39",X"6C",X"0E",X"86",X"02",X"A7",X"0F",X"39",X"6A",X"0F",X"27",X"01",
		X"39",X"6A",X"07",X"6A",X"08",X"86",X"06",X"A7",X"0F",X"39",X"6C",X"07",X"6C",X"08",X"A6",X"07",
		X"81",X"0C",X"27",X"01",X"39",X"6C",X"0E",X"86",X"40",X"A7",X"0F",X"39",X"A6",X"0C",X"6C",X"0C",
		X"CE",X"E6",X"6E",X"A6",X"C6",X"81",X"FF",X"27",X"1C",X"48",X"CE",X"E1",X"15",X"EC",X"C6",X"A7",
		X"02",X"E7",X"01",X"86",X"06",X"A7",X"07",X"6F",X"0E",X"C6",X"30",X"E7",X"0D",X"39",X"00",X"07",
		X"04",X"07",X"0C",X"FF",X"FF",X"6F",X"84",X"39",X"E6",X"FD",X"E7",X"5C",X"E7",X"6E",X"E7",X"91",
		X"EB",X"51",X"E7",X"C2",X"E7",X"C2",X"E7",X"D2",X"E7",X"E9",X"E8",X"04",X"E8",X"2A",X"E8",X"50",
		X"E8",X"6D",X"E8",X"7F",X"E8",X"80",X"E8",X"94",X"E9",X"ED",X"EB",X"D8",X"E6",X"F9",X"ED",X"38",
		X"EC",X"90",X"E6",X"BC",X"F0",X"FA",X"E8",X"A4",X"F1",X"71",X"E6",X"BD",X"E6",X"C1",X"E6",X"C5",
		X"E6",X"C9",X"E6",X"CD",X"E6",X"D1",X"E6",X"D5",X"E6",X"D9",X"E6",X"DD",X"39",X"86",X"07",X"20",
		X"20",X"86",X"08",X"20",X"1C",X"86",X"09",X"20",X"18",X"86",X"0A",X"20",X"14",X"86",X"0B",X"20",
		X"10",X"86",X"0C",X"20",X"0C",X"86",X"0D",X"20",X"08",X"86",X"0E",X"20",X"04",X"86",X"0F",X"20",
		X"00",X"8E",X"04",X"00",X"A7",X"88",X"17",X"A7",X"88",X"37",X"A7",X"88",X"57",X"A7",X"88",X"77",
		X"A7",X"89",X"00",X"97",X"A7",X"89",X"00",X"B7",X"39",X"7F",X"04",X"60",X"39",X"CE",X"02",X"00",
		X"6F",X"C4",X"6F",X"C8",X"20",X"6F",X"C8",X"40",X"6F",X"C8",X"60",X"6F",X"C9",X"00",X"80",X"6F",
		X"C9",X"00",X"A0",X"6F",X"C9",X"00",X"C0",X"6F",X"C9",X"00",X"E0",X"6F",X"C9",X"01",X"00",X"6F",
		X"C9",X"01",X"20",X"6F",X"C9",X"01",X"40",X"6F",X"C9",X"01",X"60",X"6F",X"C9",X"01",X"80",X"6F",
		X"C9",X"01",X"A0",X"6F",X"C9",X"01",X"C0",X"6F",X"C9",X"01",X"E0",X"6F",X"C9",X"02",X"00",X"6F",
		X"C9",X"02",X"20",X"6F",X"C9",X"02",X"40",X"6F",X"C9",X"02",X"C0",X"6F",X"C9",X"02",X"E0",X"6F",
		X"C9",X"03",X"00",X"6F",X"C9",X"03",X"20",X"6F",X"C9",X"03",X"40",X"39",X"8E",X"02",X"00",X"86",
		X"01",X"A7",X"84",X"86",X"FE",X"A7",X"0A",X"86",X"01",X"A7",X"0D",X"6F",X"0C",X"39",X"8E",X"02",
		X"20",X"A6",X"84",X"26",X"1B",X"86",X"01",X"A7",X"84",X"CC",X"00",X"47",X"A7",X"02",X"E7",X"01",
		X"86",X"FE",X"A7",X"0A",X"86",X"0A",X"A7",X"07",X"86",X"00",X"A7",X"0C",X"86",X"3C",X"A7",X"0D",
		X"39",X"8E",X"02",X"40",X"86",X"03",X"A7",X"84",X"CC",X"00",X"50",X"A7",X"02",X"E7",X"01",X"CC",
		X"00",X"58",X"A7",X"04",X"E6",X"03",X"CC",X"00",X"60",X"A7",X"06",X"E7",X"05",X"86",X"F8",X"A7",
		X"0A",X"86",X"09",X"A7",X"07",X"A7",X"08",X"A7",X"09",X"6F",X"88",X"12",X"86",X"30",X"A7",X"88",
		X"13",X"39",X"8E",X"02",X"A0",X"86",X"01",X"A7",X"84",X"86",X"FE",X"A7",X"0A",X"6F",X"0C",X"6F",
		X"0D",X"39",X"8E",X"02",X"C0",X"CC",X"00",X"4C",X"A7",X"02",X"E7",X"01",X"86",X"01",X"A7",X"84",
		X"86",X"F8",X"A7",X"0A",X"6F",X"0C",X"6F",X"0D",X"39",X"8E",X"02",X"E0",X"86",X"01",X"A7",X"84",
		X"CC",X"03",X"FF",X"A7",X"02",X"E7",X"01",X"86",X"08",X"A7",X"07",X"86",X"FE",X"A7",X"0A",X"86",
		X"00",X"A7",X"0C",X"39",X"8E",X"03",X"00",X"86",X"02",X"A7",X"84",X"CC",X"0E",X"80",X"A7",X"02",
		X"E7",X"01",X"CC",X"0E",X"70",X"A7",X"04",X"E7",X"03",X"86",X"04",X"A7",X"07",X"A7",X"08",X"86",
		X"E4",X"A7",X"0A",X"86",X"0E",X"A7",X"0B",X"6F",X"0C",X"39",X"8E",X"03",X"20",X"86",X"02",X"A7",
		X"84",X"CC",X"00",X"24",X"A7",X"02",X"E7",X"01",X"CC",X"00",X"26",X"A7",X"04",X"E7",X"03",X"86",
		X"FC",X"A7",X"0A",X"86",X"00",X"A7",X"0C",X"86",X"04",X"A7",X"0D",X"86",X"08",X"A7",X"0E",X"39",
		X"8E",X"03",X"40",X"86",X"01",X"A7",X"84",X"CC",X"00",X"A2",X"A7",X"02",X"E7",X"01",X"86",X"09",
		X"A7",X"07",X"86",X"FE",X"A7",X"0A",X"6F",X"0C",X"86",X"08",X"A7",X"0D",X"39",X"8E",X"03",X"60",
		X"86",X"01",X"A7",X"84",X"86",X"FE",X"A7",X"0A",X"6F",X"0C",X"86",X"01",X"A7",X"0D",X"39",X"39",
		X"8E",X"03",X"A0",X"86",X"01",X"A7",X"84",X"6F",X"01",X"6F",X"02",X"86",X"FE",X"A7",X"0A",X"6F",
		X"0C",X"6F",X"0D",X"39",X"8E",X"03",X"C0",X"86",X"01",X"A7",X"84",X"86",X"FC",X"A7",X"0A",X"6F",
		X"0C",X"6F",X"0D",X"39",X"8E",X"04",X"60",X"86",X"01",X"A7",X"84",X"86",X"FE",X"A7",X"0A",X"CC",
		X"E8",X"FA",X"ED",X"0C",X"ED",X"88",X"18",X"6F",X"88",X"12",X"86",X"04",X"A7",X"88",X"11",X"8E",
		X"04",X"80",X"86",X"01",X"A7",X"84",X"86",X"FE",X"A7",X"0A",X"CC",X"E9",X"50",X"ED",X"0C",X"ED",
		X"88",X"18",X"6F",X"88",X"12",X"86",X"04",X"A7",X"88",X"11",X"8E",X"04",X"A0",X"86",X"01",X"A7",
		X"84",X"86",X"FE",X"A7",X"0A",X"86",X"17",X"A7",X"0B",X"CC",X"E9",X"97",X"ED",X"0C",X"ED",X"88",
		X"18",X"6F",X"88",X"12",X"86",X"04",X"A7",X"88",X"11",X"39",X"5F",X"0B",X"3F",X"06",X"1F",X"23",
		X"75",X"76",X"95",X"B2",X"B1",X"B4",X"75",X"76",X"95",X"B2",X"B1",X"B4",X"76",X"78",X"99",X"B9",
		X"B8",X"B9",X"BB",X"B9",X"B8",X"B6",X"94",X"98",X"99",X"B4",X"98",X"B9",X"94",X"98",X"99",X"B4",
		X"98",X"B9",X"96",X"99",X"9D",X"B6",X"99",X"BD",X"9D",X"9D",X"99",X"BB",X"99",X"98",X"96",X"94",
		X"98",X"99",X"9B",X"99",X"B8",X"94",X"94",X"98",X"99",X"9B",X"99",X"B8",X"94",X"9E",X"9D",X"9B",
		X"99",X"98",X"99",X"9D",X"9B",X"9B",X"9A",X"9B",X"9A",X"9B",X"99",X"98",X"96",X"7F",X"E9",X"16",
		X"5F",X"0B",X"3F",X"06",X"1F",X"23",X"E0",X"E0",X"E0",X"B2",X"B2",X"B4",X"B2",X"91",X"91",X"91",
		X"B1",X"91",X"B1",X"91",X"91",X"91",X"B1",X"91",X"B1",X"92",X"92",X"92",X"B2",X"92",X"B2",X"92",
		X"92",X"92",X"B2",X"92",X"92",X"92",X"91",X"91",X"91",X"91",X"91",X"B1",X"91",X"91",X"91",X"91",
		X"91",X"91",X"B1",X"91",X"99",X"98",X"96",X"94",X"92",X"94",X"98",X"94",X"96",X"96",X"96",X"96",
		X"96",X"94",X"92",X"91",X"7F",X"E9",X"5D",X"5F",X"0B",X"3F",X"06",X"1F",X"23",X"A5",X"81",X"81",
		X"A8",X"A1",X"A5",X"81",X"81",X"A8",X"A1",X"A6",X"83",X"83",X"A8",X"A6",X"86",X"86",X"83",X"83",
		X"88",X"88",X"86",X"86",X"81",X"81",X"81",X"A1",X"81",X"A1",X"88",X"88",X"88",X"A8",X"88",X"A8",
		X"8A",X"8A",X"8A",X"AA",X"8A",X"AA",X"83",X"83",X"83",X"A3",X"83",X"83",X"83",X"88",X"88",X"88",
		X"88",X"88",X"A8",X"88",X"83",X"83",X"83",X"83",X"83",X"A3",X"83",X"85",X"85",X"85",X"85",X"85",
		X"A5",X"85",X"86",X"88",X"86",X"88",X"83",X"83",X"83",X"83",X"7F",X"E9",X"B4",X"8E",X"04",X"00",
		X"86",X"01",X"A7",X"84",X"86",X"FE",X"A7",X"0A",X"CC",X"EA",X"C5",X"ED",X"0C",X"ED",X"88",X"18",
		X"6F",X"88",X"12",X"86",X"04",X"A7",X"88",X"11",X"8E",X"04",X"20",X"86",X"01",X"A7",X"84",X"86",
		X"FE",X"A7",X"0A",X"CC",X"EA",X"50",X"ED",X"0C",X"ED",X"88",X"18",X"6F",X"88",X"12",X"86",X"04",
		X"A7",X"88",X"11",X"8E",X"04",X"40",X"86",X"01",X"A7",X"84",X"86",X"F6",X"A7",X"0A",X"86",X"17",
		X"A7",X"0B",X"CC",X"EA",X"43",X"ED",X"0C",X"ED",X"88",X"18",X"6F",X"88",X"12",X"86",X"04",X"A7",
		X"88",X"11",X"39",X"5F",X"0B",X"3F",X"06",X"1F",X"23",X"8C",X"6C",X"6C",X"7F",X"EA",X"49",X"FF",
		X"5F",X"0A",X"3F",X"06",X"1F",X"23",X"C0",X"C0",X"C0",X"9F",X"A0",X"80",X"83",X"C5",X"80",X"83",
		X"85",X"88",X"DF",X"8C",X"6C",X"8A",X"88",X"DF",X"8C",X"6C",X"8A",X"88",X"DF",X"8A",X"6A",X"88",
		X"8A",X"A5",X"A5",X"BF",X"01",X"80",X"83",X"85",X"63",X"65",X"C8",X"80",X"8A",X"88",X"8A",X"AC",
		X"8F",X"6C",X"6F",X"DF",X"B1",X"8F",X"AC",X"8A",X"88",X"DF",X"8A",X"6A",X"88",X"8A",X"A5",X"A5",
		X"1F",X"2F",X"5F",X"0D",X"B1",X"AF",X"8C",X"8F",X"AA",X"88",X"8A",X"A5",X"A3",X"A5",X"A3",X"85",
		X"88",X"AA",X"88",X"8A",X"AC",X"8F",X"6C",X"6F",X"D1",X"C0",X"74",X"74",X"71",X"71",X"6F",X"6F",
		X"6C",X"6C",X"6F",X"6F",X"6C",X"6C",X"6A",X"6A",X"68",X"68",X"1F",X"23",X"85",X"80",X"A0",X"5F",
		X"0A",X"7F",X"EA",X"59",X"FF",X"5F",X"0A",X"3F",X"06",X"1F",X"0B",X"B1",X"8C",X"8F",X"DF",X"91",
		X"71",X"8C",X"8F",X"B1",X"8C",X"8F",X"9F",X"DF",X"91",X"71",X"8C",X"8F",X"B1",X"8C",X"8F",X"DF",
		X"91",X"71",X"8C",X"8F",X"B4",X"8F",X"91",X"DF",X"94",X"74",X"8F",X"91",X"DF",X"96",X"76",X"91",
		X"94",X"B1",X"8C",X"8F",X"BF",X"01",X"DF",X"91",X"71",X"8C",X"8F",X"B4",X"8F",X"91",X"DF",X"94",
		X"74",X"8F",X"91",X"B4",X"8F",X"91",X"B1",X"8C",X"8F",X"DF",X"91",X"71",X"8C",X"8F",X"DF",X"96",
		X"76",X"91",X"94",X"DF",X"91",X"71",X"8C",X"8F",X"1F",X"2F",X"5F",X"0D",X"AC",X"AA",X"87",X"8A",
		X"A5",X"83",X"85",X"1F",X"23",X"AC",X"AA",X"AC",X"AA",X"8C",X"1F",X"2F",X"83",X"A5",X"83",X"85",
		X"A7",X"8A",X"67",X"6A",X"CC",X"C0",X"6F",X"6F",X"6C",X"6C",X"6A",X"6A",X"68",X"68",X"6A",X"6A",
		X"68",X"68",X"65",X"65",X"63",X"63",X"1F",X"0B",X"5F",X"0A",X"B1",X"8C",X"8F",X"7F",X"EA",X"D6",
		X"FF",X"8E",X"04",X"60",X"A6",X"84",X"26",X"52",X"86",X"01",X"A7",X"84",X"86",X"FE",X"A7",X"0A",
		X"CC",X"EB",X"AB",X"ED",X"0C",X"ED",X"88",X"18",X"6F",X"88",X"12",X"86",X"04",X"A7",X"88",X"11",
		X"8E",X"04",X"80",X"86",X"01",X"A7",X"84",X"86",X"FE",X"A7",X"0A",X"CC",X"EB",X"BA",X"ED",X"0C",
		X"ED",X"88",X"18",X"6F",X"88",X"12",X"86",X"04",X"A7",X"88",X"11",X"8E",X"04",X"A0",X"86",X"01",
		X"A7",X"84",X"86",X"FE",X"A7",X"0A",X"86",X"17",X"A7",X"0B",X"CC",X"EB",X"C9",X"ED",X"0C",X"ED",
		X"88",X"18",X"6F",X"88",X"12",X"86",X"04",X"A7",X"88",X"11",X"39",X"5F",X"0B",X"3F",X"03",X"1F",
		X"2F",X"A1",X"81",X"81",X"81",X"A3",X"A1",X"A1",X"E3",X"FF",X"5F",X"0B",X"3F",X"03",X"1F",X"2F",
		X"A5",X"85",X"85",X"85",X"A6",X"A6",X"A6",X"E8",X"FF",X"5F",X"0B",X"3F",X"03",X"1F",X"2F",X"A8",
		X"88",X"88",X"88",X"AA",X"AA",X"AC",X"ED",X"FF",X"8E",X"04",X"60",X"86",X"01",X"A7",X"84",X"86",
		X"FE",X"A7",X"0A",X"CC",X"EC",X"2E",X"ED",X"0C",X"ED",X"88",X"18",X"6F",X"88",X"12",X"86",X"04",
		X"A7",X"88",X"11",X"8E",X"04",X"80",X"86",X"01",X"A7",X"84",X"86",X"FE",X"A7",X"0A",X"CC",X"EC",
		X"4A",X"ED",X"0C",X"ED",X"88",X"18",X"6F",X"88",X"12",X"86",X"04",X"A7",X"88",X"11",X"8E",X"04",
		X"A0",X"86",X"01",X"A7",X"84",X"86",X"FE",X"A7",X"0A",X"86",X"17",X"A7",X"0B",X"CC",X"EC",X"66",
		X"ED",X"0C",X"ED",X"88",X"18",X"6F",X"88",X"12",X"86",X"04",X"A7",X"88",X"11",X"39",X"5F",X"0B",
		X"3F",X"05",X"1F",X"23",X"E0",X"E0",X"80",X"94",X"80",X"95",X"80",X"96",X"80",X"97",X"80",X"96",
		X"80",X"97",X"80",X"98",X"80",X"99",X"7F",X"EC",X"34",X"FF",X"5F",X"0B",X"3F",X"05",X"1F",X"23",
		X"E0",X"E0",X"80",X"8E",X"80",X"8F",X"80",X"90",X"80",X"91",X"80",X"90",X"80",X"91",X"80",X"92",
		X"80",X"93",X"7F",X"EC",X"50",X"FF",X"5F",X"0B",X"3F",X"05",X"1F",X"23",X"86",X"87",X"87",X"87",
		X"87",X"87",X"87",X"87",X"86",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"85",X"80",X"86",X"80",
		X"87",X"80",X"88",X"80",X"87",X"80",X"88",X"80",X"89",X"80",X"8A",X"80",X"7F",X"EC",X"6C",X"FF",
		X"7F",X"04",X"00",X"8E",X"04",X"60",X"86",X"01",X"A7",X"84",X"86",X"FE",X"A7",X"0A",X"CC",X"EC",
		X"E9",X"ED",X"0C",X"ED",X"88",X"18",X"6F",X"88",X"12",X"86",X"04",X"A7",X"88",X"11",X"8E",X"04",
		X"80",X"86",X"01",X"A7",X"84",X"86",X"FE",X"A7",X"0A",X"CC",X"ED",X"0F",X"ED",X"0C",X"ED",X"88",
		X"18",X"6F",X"88",X"12",X"86",X"04",X"A7",X"88",X"11",X"8E",X"04",X"A0",X"86",X"01",X"A7",X"84",
		X"86",X"FE",X"A7",X"0A",X"86",X"17",X"A7",X"0B",X"CC",X"ED",X"29",X"ED",X"0C",X"ED",X"88",X"18",
		X"6F",X"88",X"12",X"86",X"04",X"A7",X"88",X"11",X"39",X"5F",X"0B",X"3F",X"07",X"1F",X"23",X"DF",
		X"6F",X"51",X"DF",X"74",X"98",X"54",X"91",X"DF",X"6E",X"51",X"DF",X"74",X"98",X"54",X"91",X"DF",
		X"6D",X"51",X"DF",X"74",X"98",X"54",X"76",X"60",X"94",X"80",X"A0",X"FF",X"7F",X"EC",X"EF",X"5F",
		X"0B",X"3F",X"07",X"1F",X"23",X"A8",X"A8",X"A8",X"A8",X"A5",X"85",X"67",X"60",X"88",X"80",X"1F",
		X"17",X"88",X"1F",X"23",X"80",X"FF",X"7F",X"ED",X"15",X"5F",X"0B",X"3F",X"07",X"1F",X"23",X"A3",
		X"A3",X"A2",X"A2",X"A1",X"81",X"80",X"C0",X"FF",X"8E",X"04",X"60",X"86",X"01",X"A7",X"84",X"86",
		X"FE",X"A7",X"0A",X"CC",X"ED",X"8E",X"ED",X"0C",X"ED",X"88",X"18",X"6F",X"88",X"12",X"86",X"04",
		X"A7",X"88",X"11",X"8E",X"04",X"80",X"86",X"01",X"A7",X"84",X"86",X"FE",X"A7",X"0A",X"CC",X"ED",
		X"CD",X"ED",X"0C",X"ED",X"88",X"18",X"6F",X"88",X"12",X"86",X"04",X"A7",X"88",X"11",X"8E",X"04",
		X"A0",X"86",X"01",X"A7",X"84",X"86",X"FE",X"A7",X"0A",X"86",X"17",X"A7",X"0B",X"CC",X"EE",X"0C",
		X"ED",X"0C",X"ED",X"88",X"18",X"6F",X"88",X"12",X"86",X"04",X"A7",X"88",X"11",X"39",X"5F",X"09",
		X"3F",X"06",X"1F",X"23",X"9F",X"DF",X"B9",X"7B",X"79",X"96",X"99",X"94",X"96",X"DF",X"D1",X"8F",
		X"8D",X"8F",X"92",X"96",X"99",X"80",X"92",X"96",X"99",X"BD",X"BB",X"B9",X"B8",X"BF",X"01",X"9F",
		X"DF",X"B6",X"78",X"76",X"93",X"96",X"91",X"93",X"DF",X"CE",X"8C",X"8A",X"8C",X"8F",X"93",X"96",
		X"80",X"8F",X"93",X"96",X"BA",X"B8",X"B6",X"B8",X"BF",X"01",X"7F",X"ED",X"94",X"5F",X"09",X"3F",
		X"06",X"1F",X"23",X"9F",X"DF",X"B4",X"76",X"74",X"91",X"94",X"8F",X"91",X"DF",X"CC",X"8A",X"88",
		X"8A",X"8D",X"91",X"94",X"80",X"8D",X"91",X"94",X"B4",X"B2",X"B1",X"AF",X"BF",X"01",X"9F",X"DF",
		X"B1",X"73",X"71",X"8E",X"91",X"8C",X"8E",X"DF",X"C9",X"87",X"85",X"87",X"8A",X"8E",X"91",X"80",
		X"8A",X"8E",X"91",X"B1",X"AF",X"AE",X"AC",X"BF",X"01",X"7F",X"ED",X"D3",X"5F",X"09",X"3F",X"06",
		X"1F",X"17",X"9F",X"8D",X"8D",X"94",X"8D",X"8D",X"8D",X"94",X"8D",X"8D",X"8D",X"94",X"8D",X"8D",
		X"8D",X"94",X"8D",X"86",X"86",X"8D",X"86",X"86",X"86",X"8D",X"86",X"88",X"88",X"8F",X"88",X"88",
		X"88",X"8F",X"88",X"BF",X"01",X"9F",X"8A",X"8A",X"91",X"8A",X"8A",X"8A",X"91",X"8A",X"8A",X"8A",
		X"91",X"8A",X"8A",X"8A",X"91",X"8A",X"83",X"83",X"8A",X"83",X"83",X"83",X"8A",X"83",X"85",X"85",
		X"8C",X"85",X"85",X"85",X"8C",X"85",X"BF",X"01",X"7F",X"EE",X"12",X"A6",X"84",X"26",X"4A",X"39",
		X"BD",X"EE",X"8A",X"BD",X"EE",X"67",X"39",X"6C",X"88",X"1E",X"A6",X"88",X"1E",X"84",X"03",X"27",
		X"01",X"39",X"A6",X"07",X"81",X"05",X"27",X"07",X"A6",X"07",X"27",X"02",X"6A",X"07",X"39",X"86",
		X"F6",X"A7",X"0A",X"86",X"03",X"A7",X"0B",X"6A",X"07",X"39",X"A6",X"88",X"12",X"27",X"46",X"6A",
		X"88",X"1A",X"26",X"37",X"6A",X"88",X"12",X"27",X"3C",X"A6",X"88",X"17",X"A7",X"88",X"1A",X"39",
		X"86",X"FE",X"A7",X"0A",X"6F",X"88",X"1E",X"20",X"2C",X"A6",X"88",X"12",X"27",X"27",X"6A",X"88",
		X"1A",X"26",X"18",X"6A",X"88",X"12",X"27",X"1D",X"A6",X"88",X"17",X"A7",X"88",X"1A",X"A6",X"07",
		X"E6",X"88",X"1B",X"A3",X"88",X"1C",X"A7",X"07",X"E7",X"88",X"1B",X"39",X"A6",X"88",X"15",X"A7",
		X"07",X"39",X"6F",X"07",X"39",X"BD",X"F0",X"4F",X"84",X"1F",X"27",X"7A",X"81",X"1F",X"10",X"27",
		X"00",X"C1",X"BD",X"EE",X"EC",X"BD",X"EF",X"5C",X"BD",X"EE",X"CC",X"39",X"10",X"AE",X"88",X"13",
		X"48",X"31",X"A6",X"EC",X"A4",X"A7",X"02",X"E7",X"01",X"39",X"35",X"40",X"BD",X"F0",X"4F",X"84",
		X"1F",X"27",X"08",X"BD",X"EE",X"EC",X"BD",X"EF",X"0F",X"20",X"C1",X"6F",X"02",X"6F",X"01",X"E6",
		X"88",X"16",X"59",X"59",X"59",X"59",X"C4",X"07",X"E7",X"88",X"1F",X"CE",X"EF",X"3E",X"A6",X"C5",
		X"A7",X"88",X"12",X"A6",X"88",X"17",X"A7",X"88",X"1A",X"A6",X"88",X"15",X"A7",X"07",X"6F",X"88",
		X"1B",X"A6",X"88",X"1F",X"48",X"CE",X"EF",X"46",X"EC",X"C6",X"ED",X"88",X"1C",X"39",X"01",X"03",
		X"06",X"0C",X"18",X"30",X"60",X"C0",X"07",X"00",X"03",X"81",X"01",X"C2",X"00",X"E4",X"00",X"78",
		X"00",X"48",X"00",X"3C",X"00",X"4E",X"6F",X"02",X"6F",X"01",X"20",X"89",X"E6",X"88",X"16",X"59",
		X"59",X"59",X"59",X"C4",X"07",X"E7",X"88",X"1F",X"CE",X"EF",X"8B",X"A6",X"C5",X"A7",X"88",X"12",
		X"A6",X"88",X"17",X"A7",X"88",X"1A",X"A6",X"88",X"15",X"A7",X"07",X"6F",X"88",X"1B",X"CE",X"EF",
		X"93",X"A6",X"88",X"1F",X"48",X"EC",X"C6",X"ED",X"88",X"1C",X"39",X"01",X"02",X"04",X"08",X"10",
		X"20",X"40",X"80",X"07",X"00",X"03",X"80",X"01",X"C0",X"00",X"E0",X"00",X"70",X"00",X"38",X"00",
		X"1C",X"00",X"0E",X"BD",X"EF",X"A9",X"16",X"FF",X"2C",X"E6",X"88",X"16",X"59",X"59",X"59",X"59",
		X"C4",X"07",X"58",X"CE",X"EF",X"B8",X"6E",X"D5",X"EF",X"C8",X"EF",X"D5",X"EF",X"DF",X"EF",X"E6",
		X"EF",X"F4",X"EF",X"FC",X"EE",X"FA",X"F0",X"4A",X"BD",X"F0",X"4F",X"CE",X"E0",X"85",X"48",X"33",
		X"C6",X"EF",X"88",X"13",X"39",X"BD",X"F0",X"4F",X"A7",X"88",X"17",X"A7",X"88",X"1A",X"39",X"BD",
		X"F0",X"4F",X"A7",X"88",X"15",X"39",X"BD",X"F0",X"4F",X"E6",X"88",X"16",X"BD",X"F0",X"4F",X"A7",
		X"0D",X"E7",X"0C",X"39",X"EC",X"0C",X"ED",X"0E",X"6F",X"88",X"10",X"39",X"96",X"02",X"81",X"15",
		X"10",X"27",X"00",X"5C",X"BD",X"F0",X"4F",X"6C",X"88",X"10",X"A6",X"88",X"10",X"A1",X"88",X"16",
		X"23",X"01",X"39",X"EC",X"0E",X"ED",X"0C",X"39",X"39",X"BD",X"F0",X"4F",X"6C",X"88",X"10",X"A6",
		X"88",X"10",X"A1",X"88",X"16",X"27",X"07",X"BD",X"F0",X"4F",X"BD",X"F0",X"4F",X"39",X"BD",X"F0",
		X"4F",X"E6",X"88",X"16",X"BD",X"F0",X"4F",X"A7",X"0D",X"E7",X"0C",X"39",X"BD",X"F0",X"4F",X"6C",
		X"88",X"10",X"A1",X"88",X"16",X"27",X"E7",X"7E",X"F0",X"13",X"35",X"40",X"6F",X"84",X"39",X"EE",
		X"0C",X"A6",X"C4",X"A7",X"88",X"16",X"86",X"01",X"33",X"C6",X"EF",X"0C",X"A6",X"88",X"16",X"39",
		X"8E",X"04",X"60",X"86",X"01",X"A7",X"84",X"86",X"FE",X"A7",X"0A",X"CC",X"F0",X"B6",X"ED",X"0C",
		X"ED",X"88",X"18",X"6F",X"88",X"12",X"86",X"04",X"A7",X"88",X"11",X"8E",X"04",X"80",X"86",X"01",
		X"A7",X"84",X"86",X"FE",X"A7",X"0A",X"CC",X"F0",X"CE",X"ED",X"0C",X"ED",X"88",X"18",X"6F",X"88",
		X"12",X"86",X"04",X"A7",X"88",X"11",X"8E",X"04",X"A0",X"86",X"01",X"A7",X"84",X"86",X"FE",X"A7",
		X"0A",X"86",X"17",X"A7",X"0B",X"CC",X"F0",X"E6",X"ED",X"0C",X"ED",X"88",X"18",X"6F",X"88",X"12",
		X"86",X"04",X"A7",X"88",X"11",X"39",X"5F",X"09",X"3F",X"07",X"1F",X"23",X"DF",X"B9",X"79",X"79",
		X"DF",X"B9",X"79",X"79",X"92",X"60",X"76",X"B9",X"95",X"60",X"79",X"BC",X"FD",X"FF",X"5F",X"09",
		X"3F",X"07",X"1F",X"23",X"DF",X"B4",X"74",X"74",X"DF",X"B4",X"74",X"74",X"8D",X"60",X"72",X"B6",
		X"90",X"60",X"75",X"B9",X"F9",X"FF",X"5F",X"09",X"3F",X"07",X"1F",X"17",X"AD",X"AC",X"AA",X"A8",
		X"8A",X"60",X"6B",X"B2",X"8D",X"60",X"70",X"B5",X"F4",X"FF",X"8E",X"04",X"60",X"86",X"01",X"A7",
		X"84",X"86",X"FE",X"A7",X"0A",X"CC",X"F1",X"4D",X"ED",X"0C",X"ED",X"88",X"18",X"6F",X"88",X"12",
		X"86",X"04",X"A7",X"88",X"11",X"8E",X"04",X"80",X"86",X"01",X"A7",X"84",X"86",X"FE",X"A7",X"0A",
		X"CC",X"F1",X"5F",X"ED",X"0C",X"ED",X"88",X"18",X"6F",X"88",X"12",X"86",X"04",X"A7",X"88",X"11",
		X"8E",X"04",X"A0",X"6F",X"01",X"6F",X"02",X"86",X"FE",X"A7",X"0A",X"39",X"CC",X"F1",X"70",X"ED",
		X"0C",X"ED",X"88",X"18",X"6F",X"88",X"12",X"86",X"04",X"A7",X"88",X"11",X"39",X"5F",X"0A",X"3F",
		X"09",X"1F",X"23",X"7E",X"7E",X"7E",X"7E",X"9B",X"99",X"9B",X"7B",X"7B",X"DB",X"A0",X"FF",X"5F",
		X"0A",X"3F",X"09",X"1F",X"23",X"79",X"79",X"79",X"79",X"96",X"94",X"96",X"76",X"76",X"D6",X"A0",
		X"FF",X"8E",X"04",X"60",X"86",X"01",X"A7",X"84",X"86",X"FE",X"A7",X"0A",X"CC",X"F1",X"C7",X"ED",
		X"0C",X"ED",X"88",X"18",X"6F",X"88",X"12",X"86",X"04",X"A7",X"88",X"11",X"8E",X"04",X"80",X"86",
		X"01",X"A7",X"84",X"86",X"FE",X"A7",X"0A",X"CC",X"F1",X"F9",X"ED",X"0C",X"ED",X"88",X"18",X"6F",
		X"88",X"12",X"86",X"04",X"A7",X"88",X"11",X"8E",X"04",X"A0",X"86",X"01",X"A7",X"84",X"86",X"FE",
		X"A7",X"0A",X"86",X"17",X"A7",X"0B",X"CC",X"F2",X"2B",X"ED",X"0C",X"ED",X"88",X"18",X"6F",X"88",
		X"12",X"86",X"04",X"A7",X"88",X"11",X"39",X"5F",X"0B",X"3F",X"07",X"1F",X"23",X"94",X"76",X"71",
		X"74",X"74",X"76",X"71",X"94",X"76",X"71",X"74",X"74",X"76",X"71",X"76",X"79",X"60",X"76",X"79",
		X"60",X"76",X"79",X"6F",X"6F",X"71",X"71",X"72",X"72",X"74",X"74",X"72",X"72",X"76",X"79",X"74",
		X"74",X"78",X"7B",X"79",X"99",X"99",X"7B",X"9D",X"FF",X"5F",X"0B",X"3F",X"07",X"1F",X"23",X"8D",
		X"6D",X"6D",X"6D",X"6D",X"6D",X"6D",X"8E",X"6E",X"6E",X"6E",X"6E",X"6E",X"6E",X"72",X"6F",X"60",
		X"72",X"6F",X"60",X"73",X"6F",X"6A",X"6A",X"6C",X"6C",X"6D",X"6D",X"6E",X"6E",X"6D",X"6D",X"72",
		X"72",X"6F",X"6F",X"74",X"74",X"71",X"91",X"91",X"72",X"94",X"FF",X"5F",X"0B",X"3F",X"07",X"1F",
		X"23",X"81",X"68",X"65",X"61",X"61",X"68",X"65",X"82",X"68",X"65",X"62",X"62",X"68",X"65",X"66",
		X"63",X"60",X"66",X"63",X"60",X"67",X"63",X"69",X"69",X"6B",X"6B",X"6C",X"6C",X"6D",X"6D",X"66",
		X"66",X"6D",X"6A",X"68",X"68",X"6F",X"6C",X"61",X"81",X"81",X"68",X"8D",X"FF",X"86",X"FF",X"B7",
		X"01",X"12",X"B7",X"01",X"13",X"B7",X"01",X"14",X"B7",X"01",X"18",X"B7",X"01",X"19",X"B7",X"01",
		X"1A",X"BD",X"F3",X"14",X"7E",X"F2",X"78",X"39",X"8E",X"04",X"60",X"A6",X"84",X"26",X"12",X"8E",
		X"04",X"00",X"A6",X"84",X"26",X"0B",X"C6",X"07",X"F7",X"40",X"00",X"86",X"FF",X"B7",X"40",X"01",
		X"39",X"5F",X"F7",X"40",X"00",X"A6",X"01",X"B7",X"40",X"01",X"5C",X"F7",X"40",X"00",X"A6",X"02",
		X"B7",X"40",X"01",X"5C",X"F7",X"40",X"00",X"A6",X"88",X"21",X"B7",X"40",X"01",X"5C",X"F7",X"40",
		X"00",X"A6",X"88",X"22",X"B7",X"40",X"01",X"5C",X"F7",X"40",X"00",X"A6",X"88",X"41",X"B7",X"40",
		X"01",X"5C",X"F7",X"40",X"00",X"A6",X"88",X"42",X"B7",X"40",X"01",X"5C",X"F7",X"40",X"00",X"A6",
		X"88",X"4B",X"B7",X"40",X"01",X"C6",X"FF",X"A6",X"0A",X"44",X"56",X"A6",X"88",X"2A",X"44",X"56",
		X"A6",X"88",X"4A",X"44",X"56",X"56",X"56",X"44",X"44",X"44",X"56",X"56",X"56",X"86",X"07",X"B7",
		X"40",X"00",X"F7",X"40",X"01",X"C6",X"08",X"F7",X"40",X"00",X"A6",X"07",X"B7",X"40",X"01",X"5C",
		X"F7",X"40",X"00",X"A6",X"88",X"27",X"B7",X"40",X"01",X"5C",X"F7",X"40",X"00",X"A6",X"88",X"47",
		X"B7",X"40",X"01",X"39",X"8E",X"02",X"00",X"86",X"0F",X"97",X"03",X"0F",X"05",X"A6",X"84",X"27",
		X"03",X"BD",X"F3",X"35",X"96",X"05",X"81",X"03",X"27",X"0A",X"0A",X"03",X"27",X"06",X"86",X"20",
		X"30",X"86",X"20",X"E9",X"39",X"A6",X"84",X"81",X"01",X"27",X"07",X"81",X"02",X"27",X"48",X"16",
		X"00",X"B0",X"D6",X"05",X"58",X"F7",X"20",X"00",X"A6",X"01",X"B7",X"20",X"01",X"5C",X"F7",X"20",
		X"00",X"A6",X"02",X"B7",X"20",X"01",X"96",X"05",X"8B",X"08",X"B7",X"20",X"00",X"A6",X"07",X"B7",
		X"20",X"01",X"A6",X"0B",X"27",X"08",X"C6",X"06",X"F7",X"20",X"00",X"B7",X"20",X"01",X"96",X"05",
		X"10",X"8E",X"01",X"12",X"31",X"A6",X"A6",X"0A",X"44",X"69",X"A4",X"C6",X"06",X"31",X"A5",X"44",
		X"44",X"44",X"69",X"A4",X"0C",X"05",X"39",X"D6",X"05",X"C1",X"02",X"27",X"B5",X"58",X"F7",X"20",
		X"00",X"A6",X"01",X"B7",X"20",X"01",X"5C",X"F7",X"20",X"00",X"A6",X"02",X"B7",X"20",X"01",X"5C",
		X"F7",X"20",X"00",X"A6",X"03",X"B7",X"20",X"01",X"5C",X"F7",X"20",X"00",X"A6",X"04",X"B7",X"20",
		X"01",X"D6",X"05",X"CB",X"08",X"F7",X"20",X"00",X"A6",X"07",X"B7",X"20",X"01",X"5C",X"F7",X"20",
		X"00",X"A6",X"08",X"B7",X"20",X"01",X"A6",X"0B",X"27",X"08",X"C6",X"06",X"F7",X"20",X"00",X"B7",
		X"20",X"01",X"96",X"05",X"10",X"8E",X"01",X"12",X"31",X"A6",X"A6",X"0A",X"46",X"69",X"A4",X"46",
		X"69",X"21",X"C6",X"06",X"31",X"A5",X"46",X"46",X"69",X"A4",X"46",X"69",X"21",X"0C",X"05",X"0C",
		X"05",X"39",X"D6",X"05",X"C1",X"02",X"10",X"27",X"FF",X"48",X"C1",X"01",X"27",X"89",X"58",X"F7",
		X"20",X"00",X"A6",X"01",X"B7",X"20",X"01",X"5C",X"F7",X"20",X"00",X"A6",X"02",X"B7",X"20",X"01",
		X"5C",X"F7",X"20",X"00",X"A6",X"03",X"B7",X"20",X"01",X"5C",X"F7",X"20",X"00",X"A6",X"04",X"B7",
		X"20",X"01",X"5C",X"F7",X"20",X"00",X"A6",X"05",X"B7",X"20",X"01",X"5C",X"F7",X"20",X"00",X"A6",
		X"06",X"B7",X"20",X"01",X"D6",X"05",X"CB",X"08",X"F7",X"20",X"00",X"A6",X"07",X"B7",X"20",X"01",
		X"5C",X"F7",X"20",X"00",X"A6",X"08",X"B7",X"20",X"01",X"5C",X"F7",X"20",X"00",X"A6",X"08",X"B7",
		X"20",X"01",X"A6",X"0B",X"27",X"08",X"C6",X"06",X"F7",X"20",X"00",X"B7",X"20",X"01",X"96",X"05",
		X"10",X"8E",X"01",X"12",X"31",X"A6",X"A6",X"0A",X"46",X"69",X"A4",X"46",X"69",X"21",X"46",X"69",
		X"22",X"C6",X"06",X"31",X"A5",X"46",X"69",X"A0",X"46",X"69",X"A0",X"46",X"69",X"A4",X"0C",X"05",
		X"0C",X"05",X"0C",X"05",X"39",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E0",X"68",X"E0",X"1C",X"FF",X"FF",X"FF",X"FF",X"E0",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
