library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity rom_cpu1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of rom_cpu1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"31",X"00",X"6C",X"C3",X"70",X"02",X"C7",X"C7",X"5E",X"23",X"56",X"23",X"EB",X"C9",X"C7",X"C7",
		X"77",X"23",X"10",X"FC",X"0D",X"20",X"F9",X"C9",X"D1",X"5F",X"CB",X"23",X"16",X"00",X"19",X"5E",
		X"23",X"56",X"EB",X"E9",X"C7",X"C7",X"C7",X"C7",X"21",X"01",X"90",X"C3",X"AD",X"01",X"C7",X"C7",
		X"73",X"CB",X"D4",X"72",X"CB",X"94",X"C9",X"C7",X"F5",X"E5",X"21",X"01",X"60",X"3A",X"00",X"90",
		X"17",X"38",X"05",X"36",X"0A",X"C3",X"A9",X"00",X"7E",X"A7",X"C2",X"A9",X"00",X"C3",X"93",X"00",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"F5",X"E5",X"21",X"01",X"60",X"3A",X"00",X"90",X"17",X"38",
		X"04",X"36",X"0A",X"18",X"1A",X"7E",X"A7",X"20",X"16",X"3A",X"03",X"60",X"A7",X"20",X"10",X"3E",
		X"55",X"32",X"06",X"60",X"32",X"16",X"6B",X"32",X"38",X"6E",X"3E",X"03",X"32",X"03",X"60",X"E1",
		X"F1",X"ED",X"45",X"3A",X"02",X"60",X"A7",X"20",X"10",X"3E",X"55",X"32",X"05",X"60",X"32",X"09",
		X"6B",X"32",X"25",X"6E",X"3E",X"03",X"32",X"02",X"60",X"3A",X"00",X"80",X"E1",X"F1",X"FB",X"C9",
		X"06",X"00",X"4F",X"21",X"6D",X"01",X"09",X"EB",X"7E",X"DD",X"BE",X"00",X"C2",X"57",X"01",X"FD",
		X"BE",X"00",X"C2",X"57",X"01",X"34",X"DD",X"34",X"00",X"FD",X"34",X"00",X"7E",X"DD",X"BE",X"00",
		X"C2",X"57",X"01",X"FD",X"BE",X"00",X"C2",X"57",X"01",X"1A",X"BE",X"28",X"04",X"D0",X"C3",X"57",
		X"01",X"36",X"00",X"DD",X"36",X"00",X"00",X"FD",X"36",X"00",X"00",X"13",X"3A",X"04",X"60",X"21",
		X"5B",X"6B",X"BE",X"C2",X"62",X"01",X"21",X"91",X"6E",X"BE",X"C2",X"62",X"01",X"21",X"04",X"60",
		X"1A",X"86",X"FE",X"63",X"38",X"02",X"3E",X"63",X"77",X"21",X"5B",X"6B",X"1A",X"86",X"FE",X"63",
		X"38",X"02",X"3E",X"63",X"77",X"21",X"91",X"6E",X"1A",X"86",X"FE",X"63",X"38",X"02",X"3E",X"63",
		X"77",X"3A",X"04",X"60",X"21",X"5B",X"6B",X"BE",X"C2",X"62",X"01",X"21",X"91",X"6E",X"BE",X"C2",
		X"62",X"01",X"3A",X"00",X"60",X"CB",X"47",X"20",X"03",X"CD",X"33",X"1E",X"3E",X"00",X"CD",X"86",
		X"0F",X"3E",X"40",X"CD",X"98",X"3B",X"3A",X"00",X"60",X"CB",X"7F",X"C0",X"21",X"DB",X"61",X"36",
		X"80",X"3E",X"FF",X"32",X"0B",X"60",X"C9",X"36",X"00",X"DD",X"36",X"00",X"00",X"FD",X"36",X"00",
		X"00",X"C9",X"AF",X"32",X"04",X"60",X"32",X"5B",X"6B",X"32",X"91",X"6E",X"C9",X"01",X"01",X"01",
		X"02",X"01",X"03",X"01",X"04",X"01",X"05",X"02",X"01",X"02",X"02",X"02",X"03",X"03",X"01",X"03",
		X"02",X"04",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"02",X"01",X"03",X"01",X"04",X"01",X"05",X"02",X"01",X"02",X"02",X"02",X"03",X"03",X"01",X"03",
		X"02",X"04",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"CB",X"7E",X"20",
		X"FC",X"CB",X"7E",X"28",X"FC",X"21",X"01",X"60",X"3A",X"00",X"90",X"17",X"38",X"03",X"36",X"0A",
		X"C9",X"7E",X"A7",X"CA",X"C8",X"01",X"35",X"C9",X"21",X"03",X"60",X"7E",X"A7",X"CA",X"11",X"02",
		X"35",X"C2",X"11",X"02",X"3E",X"55",X"21",X"06",X"60",X"BE",X"20",X"2B",X"21",X"16",X"6B",X"BE",
		X"20",X"25",X"21",X"38",X"6E",X"BE",X"20",X"1F",X"3A",X"03",X"90",X"2F",X"E6",X"F0",X"0F",X"0F",
		X"0F",X"DD",X"E5",X"FD",X"E5",X"11",X"08",X"60",X"DD",X"21",X"3E",X"6B",X"FD",X"21",X"6C",X"6E",
		X"CD",X"B0",X"00",X"FD",X"E1",X"DD",X"E1",X"AF",X"32",X"06",X"60",X"32",X"16",X"6B",X"32",X"38",
		X"6E",X"21",X"02",X"60",X"7E",X"A7",X"C8",X"35",X"C0",X"3E",X"55",X"21",X"05",X"60",X"BE",X"20",
		X"44",X"21",X"09",X"6B",X"BE",X"20",X"3E",X"21",X"25",X"6E",X"BE",X"20",X"38",X"DD",X"E5",X"FD",
		X"E5",X"11",X"07",X"60",X"DD",X"21",X"27",X"6B",X"FD",X"21",X"4F",X"6E",X"3A",X"03",X"90",X"67",
		X"CB",X"0F",X"CB",X"0F",X"CB",X"0F",X"CB",X"0F",X"AC",X"20",X"0B",X"11",X"08",X"60",X"DD",X"21",
		X"3E",X"6B",X"FD",X"21",X"6C",X"6E",X"7C",X"2F",X"E6",X"0F",X"CB",X"27",X"C6",X"20",X"CD",X"B0",
		X"00",X"FD",X"E1",X"DD",X"E1",X"AF",X"32",X"05",X"60",X"32",X"09",X"6B",X"32",X"25",X"6E",X"C9",
		X"3A",X"00",X"90",X"E6",X"60",X"CA",X"80",X"5D",X"21",X"00",X"60",X"01",X"10",X"00",X"AF",X"77",
		X"23",X"10",X"FC",X"0D",X"20",X"F9",X"EF",X"21",X"00",X"70",X"01",X"04",X"00",X"AF",X"D7",X"21",
		X"E5",X"02",X"E5",X"11",X"94",X"6A",X"01",X"03",X"00",X"ED",X"B0",X"E1",X"06",X"05",X"11",X"94",
		X"6A",X"C5",X"E5",X"01",X"03",X"00",X"ED",X"B0",X"E1",X"C1",X"10",X"F5",X"21",X"AE",X"1D",X"11",
		X"A3",X"6A",X"06",X"05",X"C5",X"E5",X"01",X"0A",X"00",X"ED",X"B0",X"E1",X"C1",X"10",X"F5",X"21",
		X"00",X"A0",X"36",X"00",X"21",X"50",X"50",X"22",X"15",X"60",X"21",X"CE",X"61",X"36",X"80",X"CD",
		X"8C",X"3B",X"ED",X"56",X"21",X"00",X"80",X"36",X"00",X"FB",X"AF",X"32",X"0A",X"60",X"AF",X"CD",
		X"98",X"3B",X"C3",X"E8",X"02",X"01",X"00",X"00",X"EF",X"3A",X"0A",X"60",X"CB",X"47",X"20",X"07",
		X"11",X"3C",X"03",X"06",X"0C",X"18",X"05",X"11",X"6C",X"03",X"06",X"11",X"C5",X"EB",X"5E",X"23",
		X"56",X"23",X"EB",X"E5",X"DD",X"E1",X"CB",X"7E",X"20",X"04",X"13",X"13",X"18",X"1E",X"CB",X"76",
		X"28",X"0D",X"23",X"7E",X"A7",X"28",X"05",X"35",X"13",X"13",X"18",X"10",X"2B",X"CB",X"B6",X"EB",
		X"5E",X"23",X"56",X"23",X"EB",X"D5",X"01",X"2B",X"03",X"C5",X"E9",X"D1",X"C1",X"10",X"CD",X"21",
		X"0A",X"60",X"34",X"CD",X"73",X"3B",X"CD",X"13",X"1F",X"C3",X"E8",X"02",X"DF",X"61",X"8A",X"07",
		X"CE",X"61",X"B0",X"03",X"D5",X"61",X"74",X"04",X"DB",X"61",X"71",X"05",X"DD",X"61",X"48",X"06",
		X"E2",X"61",X"68",X"09",X"E8",X"61",X"47",X"24",X"00",X"62",X"6B",X"33",X"D6",X"62",X"F5",X"0F",
		X"EC",X"62",X"F5",X"0F",X"02",X"63",X"58",X"11",X"9C",X"62",X"6E",X"2A",X"28",X"62",X"6E",X"2A",
		X"45",X"62",X"6E",X"2A",X"62",X"62",X"6E",X"2A",X"7F",X"62",X"6E",X"2A",X"20",X"63",X"57",X"12",
		X"47",X"63",X"15",X"15",X"58",X"63",X"15",X"15",X"69",X"63",X"54",X"16",X"7B",X"63",X"54",X"16",
		X"8D",X"63",X"DE",X"17",X"9B",X"63",X"DE",X"17",X"A9",X"63",X"25",X"19",X"BE",X"63",X"25",X"19",
		X"D3",X"63",X"25",X"19",X"11",X"63",X"58",X"11",X"B9",X"62",X"6E",X"2A",X"C5",X"69",X"9D",X"3B",
		X"DD",X"CB",X"00",X"6E",X"28",X"0B",X"DD",X"7E",X"02",X"21",X"BD",X"03",X"DF",X"EF",X"03",X"69",
		X"04",X"DD",X"CB",X"00",X"EE",X"DD",X"36",X"02",X"00",X"AF",X"32",X"00",X"60",X"32",X"00",X"A0",
		X"CD",X"8C",X"3B",X"3E",X"00",X"CD",X"A0",X"1B",X"21",X"66",X"1D",X"CD",X"39",X"1D",X"DD",X"36",
		X"03",X"00",X"DD",X"36",X"04",X"08",X"DD",X"36",X"05",X"10",X"DD",X"36",X"06",X"60",X"C9",X"DD",
		X"7E",X"03",X"FE",X"C0",X"38",X"0C",X"DD",X"36",X"01",X"78",X"DD",X"CB",X"00",X"F6",X"DD",X"34",
		X"02",X"C9",X"DD",X"7E",X"05",X"A7",X"28",X"40",X"DD",X"7E",X"04",X"D6",X"08",X"38",X"39",X"DD",
		X"77",X"04",X"DD",X"7E",X"06",X"16",X"00",X"DD",X"5E",X"03",X"CB",X"3B",X"CB",X"3B",X"CB",X"3B",
		X"21",X"C0",X"D1",X"19",X"77",X"3E",X"6F",X"DD",X"86",X"05",X"21",X"FF",X"D1",X"A7",X"ED",X"52",
		X"77",X"DD",X"7E",X"06",X"C6",X"20",X"21",X"00",X"D2",X"19",X"77",X"C6",X"10",X"21",X"20",X"D2",
		X"19",X"77",X"DD",X"34",X"06",X"DD",X"35",X"05",X"DD",X"7E",X"04",X"C6",X"03",X"DD",X"77",X"04",
		X"DD",X"7E",X"03",X"C6",X"03",X"DD",X"77",X"03",X"32",X"43",X"D0",X"32",X"04",X"D0",X"32",X"24",
		X"D0",X"47",X"3E",X"00",X"90",X"32",X"63",X"D0",X"C9",X"06",X"07",X"CD",X"8D",X"1B",X"21",X"D5",
		X"61",X"36",X"80",X"C9",X"DD",X"7E",X"02",X"21",X"7B",X"04",X"DF",X"83",X"04",X"AF",X"04",X"26",
		X"05",X"50",X"05",X"21",X"17",X"60",X"11",X"FD",X"69",X"CD",X"95",X"1B",X"DD",X"36",X"00",X"80",
		X"DD",X"36",X"02",X"01",X"CD",X"A9",X"05",X"3E",X"02",X"CD",X"A0",X"1B",X"3E",X"80",X"32",X"00",
		X"60",X"CD",X"DF",X"1C",X"3E",X"01",X"32",X"00",X"60",X"21",X"E2",X"61",X"36",X"80",X"C9",X"21",
		X"E8",X"61",X"CB",X"6E",X"CA",X"D0",X"04",X"3A",X"15",X"60",X"E6",X"07",X"87",X"5F",X"16",X"00",
		X"21",X"61",X"05",X"19",X"7E",X"DD",X"77",X"03",X"23",X"7E",X"DD",X"77",X"01",X"C3",X"21",X"05",
		X"3A",X"EA",X"61",X"FE",X"01",X"20",X"05",X"21",X"EF",X"61",X"18",X"03",X"21",X"30",X"60",X"3A",
		X"07",X"62",X"BE",X"28",X"04",X"38",X"06",X"18",X"08",X"06",X"00",X"18",X"06",X"06",X"08",X"18",
		X"02",X"06",X"02",X"DD",X"7E",X"05",X"A7",X"28",X"05",X"DD",X"35",X"05",X"18",X"18",X"3A",X"15",
		X"60",X"E6",X"0F",X"DD",X"77",X"05",X"3A",X"16",X"60",X"E6",X"03",X"5F",X"16",X"00",X"21",X"5B",
		X"05",X"19",X"7E",X"DD",X"77",X"04",X"DD",X"7E",X"04",X"B0",X"DD",X"77",X"03",X"DD",X"36",X"01",
		X"03",X"DD",X"CB",X"00",X"F6",X"C9",X"21",X"17",X"60",X"11",X"FD",X"69",X"CD",X"95",X"1B",X"DD",
		X"36",X"02",X"03",X"DD",X"36",X"00",X"E0",X"DD",X"36",X"01",X"78",X"CD",X"B2",X"1B",X"CD",X"C9",
		X"1B",X"CD",X"B5",X"0D",X"3E",X"01",X"CD",X"E1",X"1B",X"CD",X"DF",X"1C",X"CD",X"5D",X"22",X"C9",
		X"06",X"06",X"CD",X"8D",X"1B",X"21",X"CE",X"61",X"36",X"80",X"C9",X"04",X"00",X"04",X"04",X"00",
		X"00",X"04",X"10",X"01",X"14",X"0C",X"0C",X"09",X"08",X"03",X"06",X"06",X"04",X"08",X"08",X"02",
		X"04",X"DD",X"CB",X"00",X"6E",X"C2",X"CE",X"05",X"AF",X"32",X"0B",X"60",X"21",X"17",X"60",X"11",
		X"FD",X"69",X"CD",X"95",X"1B",X"DD",X"36",X"00",X"A0",X"AF",X"32",X"00",X"60",X"3E",X"02",X"CD",
		X"A0",X"1B",X"3E",X"80",X"32",X"00",X"60",X"CD",X"10",X"1E",X"21",X"73",X"1D",X"CD",X"39",X"1D",
		X"CD",X"39",X"1D",X"CD",X"A9",X"05",X"C3",X"E5",X"05",X"3A",X"02",X"90",X"07",X"07",X"E6",X"03",
		X"5F",X"16",X"00",X"21",X"44",X"06",X"19",X"7E",X"32",X"17",X"60",X"32",X"18",X"60",X"3E",X"01",
		X"32",X"59",X"60",X"32",X"97",X"61",X"AF",X"32",X"28",X"60",X"32",X"29",X"60",X"C9",X"3A",X"04",
		X"60",X"FE",X"02",X"38",X"10",X"DD",X"CB",X"00",X"66",X"20",X"0A",X"DD",X"CB",X"00",X"E6",X"21",
		X"98",X"1D",X"CD",X"39",X"1D",X"3A",X"04",X"60",X"21",X"00",X"90",X"4E",X"CB",X"69",X"28",X"0C",
		X"FE",X"02",X"DA",X"43",X"06",X"CB",X"71",X"28",X"08",X"C3",X"43",X"06",X"01",X"01",X"81",X"18",
		X"03",X"01",X"02",X"C1",X"21",X"00",X"60",X"70",X"3A",X"04",X"60",X"91",X"32",X"04",X"60",X"3A",
		X"5B",X"6B",X"91",X"32",X"5B",X"6B",X"3A",X"91",X"6E",X"91",X"32",X"91",X"6E",X"21",X"0C",X"60",
		X"11",X"12",X"60",X"CD",X"95",X"1B",X"CD",X"DF",X"1C",X"CD",X"33",X"1E",X"06",X"1E",X"CD",X"76",
		X"0F",X"DD",X"36",X"00",X"00",X"21",X"E2",X"61",X"36",X"80",X"23",X"23",X"36",X"00",X"3E",X"15",
		X"CD",X"86",X"0F",X"C9",X"02",X"05",X"04",X"03",X"CD",X"8C",X"3B",X"21",X"DF",X"61",X"11",X"FD",
		X"69",X"CD",X"95",X"1B",X"21",X"17",X"60",X"3A",X"00",X"60",X"CB",X"6F",X"28",X"01",X"23",X"7E",
		X"D6",X"01",X"27",X"77",X"A7",X"28",X"0B",X"3A",X"00",X"60",X"CB",X"77",X"CA",X"CD",X"06",X"C3",
		X"98",X"06",X"21",X"00",X"60",X"CB",X"76",X"CA",X"00",X"07",X"CB",X"6E",X"20",X"04",X"CB",X"D6",
		X"18",X"02",X"CB",X"CE",X"7E",X"E6",X"06",X"FE",X"06",X"CA",X"00",X"07",X"CD",X"45",X"07",X"CD",
		X"60",X"07",X"CD",X"8F",X"1F",X"CD",X"EE",X"3F",X"21",X"00",X"60",X"CB",X"6E",X"20",X"08",X"CB",
		X"4E",X"20",X"2A",X"CB",X"EE",X"18",X"06",X"CB",X"56",X"20",X"22",X"CB",X"AE",X"DD",X"E5",X"21",
		X"52",X"60",X"11",X"90",X"60",X"DD",X"21",X"90",X"61",X"7E",X"DD",X"46",X"00",X"DD",X"77",X"00",
		X"70",X"23",X"DD",X"23",X"E5",X"AF",X"ED",X"52",X"E1",X"20",X"EE",X"DD",X"E1",X"CD",X"B2",X"1B",
		X"CD",X"C9",X"1B",X"3A",X"00",X"60",X"06",X"00",X"CB",X"6F",X"28",X"08",X"3A",X"02",X"90",X"CB",
		X"5F",X"28",X"01",X"05",X"21",X"00",X"A0",X"70",X"21",X"28",X"60",X"3A",X"00",X"60",X"CB",X"6F",
		X"28",X"03",X"21",X"29",X"60",X"7E",X"21",X"E2",X"61",X"36",X"80",X"23",X"23",X"77",X"18",X"40",
		X"CD",X"45",X"07",X"CD",X"60",X"07",X"21",X"00",X"60",X"CB",X"BE",X"CD",X"8F",X"1F",X"CD",X"EE",
		X"3F",X"1E",X"17",X"CD",X"91",X"0F",X"3A",X"0B",X"60",X"A7",X"C2",X"2B",X"07",X"3A",X"1D",X"6C",
		X"A7",X"28",X"08",X"06",X"0A",X"CD",X"76",X"0F",X"C3",X"16",X"07",X"AF",X"32",X"00",X"A0",X"32",
		X"00",X"60",X"21",X"CE",X"61",X"3A",X"04",X"60",X"A7",X"28",X"03",X"21",X"DB",X"61",X"36",X"80",
		X"DD",X"36",X"00",X"00",X"C9",X"21",X"0C",X"60",X"11",X"00",X"6F",X"01",X"06",X"00",X"ED",X"B0",
		X"3E",X"30",X"21",X"00",X"60",X"CB",X"6E",X"CA",X"5C",X"07",X"3E",X"31",X"CD",X"98",X"3B",X"C9",
		X"CD",X"B2",X"1B",X"CD",X"B5",X"0D",X"CD",X"C9",X"1B",X"3E",X"03",X"CD",X"E1",X"1B",X"21",X"B8",
		X"1D",X"CD",X"39",X"1D",X"21",X"C4",X"1D",X"3A",X"00",X"60",X"CB",X"6F",X"28",X"03",X"21",X"CF",
		X"1D",X"CD",X"39",X"1D",X"06",X"3C",X"CD",X"76",X"0F",X"C9",X"FD",X"21",X"E8",X"63",X"DD",X"36",
		X"02",X"0D",X"21",X"75",X"64",X"11",X"80",X"70",X"E5",X"D5",X"FD",X"7E",X"00",X"A7",X"28",X"07",
		X"87",X"87",X"4F",X"06",X"00",X"ED",X"B0",X"AF",X"12",X"FD",X"7E",X"00",X"FE",X"08",X"30",X"08",
		X"D1",X"D5",X"21",X"20",X"00",X"19",X"36",X"00",X"D1",X"E1",X"01",X"40",X"00",X"09",X"EB",X"09",
		X"EB",X"FD",X"23",X"DD",X"35",X"02",X"20",X"D0",X"AF",X"21",X"E8",X"63",X"01",X"01",X"0D",X"D7",
		X"C9",X"E5",X"3A",X"00",X"60",X"CB",X"6F",X"28",X"08",X"3A",X"02",X"90",X"CB",X"5F",X"C2",X"19",
		X"08",X"3E",X"FF",X"DD",X"96",X"07",X"CD",X"2B",X"09",X"E1",X"DD",X"5E",X"08",X"CB",X"23",X"16",
		X"00",X"19",X"CF",X"7C",X"E6",X"30",X"F6",X"C0",X"FD",X"86",X"00",X"FD",X"77",X"00",X"DD",X"7E",
		X"05",X"D6",X"07",X"FD",X"77",X"03",X"CB",X"24",X"CB",X"24",X"CB",X"24",X"CB",X"24",X"DD",X"7E",
		X"09",X"84",X"FD",X"75",X"01",X"FD",X"77",X"02",X"C9",X"DD",X"7E",X"07",X"CD",X"2B",X"09",X"E1",
		X"DD",X"5E",X"08",X"CB",X"23",X"16",X"00",X"19",X"CF",X"7C",X"EE",X"30",X"E6",X"30",X"F6",X"C0",
		X"FD",X"86",X"00",X"FD",X"77",X"00",X"3E",X"F9",X"DD",X"96",X"05",X"FD",X"77",X"03",X"18",X"C6",
		X"3A",X"00",X"60",X"CB",X"6F",X"28",X"07",X"3A",X"02",X"90",X"CB",X"5F",X"20",X"15",X"3E",X"FF",
		X"93",X"CD",X"2B",X"09",X"FD",X"CB",X"00",X"FE",X"FD",X"CB",X"00",X"F6",X"7A",X"D6",X"07",X"FD",
		X"77",X"03",X"C9",X"7B",X"CD",X"2B",X"09",X"FD",X"CB",X"00",X"FE",X"FD",X"CB",X"00",X"F6",X"3E",
		X"F9",X"92",X"FD",X"77",X"03",X"C9",X"3A",X"00",X"60",X"CB",X"6F",X"28",X"07",X"3A",X"02",X"90",
		X"CB",X"5F",X"20",X"15",X"3E",X"FB",X"93",X"CD",X"2B",X"09",X"FD",X"CB",X"00",X"FE",X"FD",X"CB",
		X"00",X"B6",X"7A",X"D6",X"03",X"FD",X"77",X"03",X"C9",X"7B",X"D6",X"04",X"CD",X"2B",X"09",X"FD",
		X"CB",X"00",X"FE",X"FD",X"CB",X"00",X"B6",X"3E",X"FD",X"92",X"FD",X"77",X"03",X"C9",X"7E",X"FD",
		X"77",X"01",X"23",X"7E",X"23",X"07",X"07",X"07",X"07",X"FD",X"77",X"02",X"7E",X"E6",X"0F",X"FD",
		X"86",X"02",X"FD",X"77",X"02",X"3A",X"00",X"60",X"CB",X"6F",X"28",X"07",X"3A",X"02",X"90",X"CB",
		X"5F",X"20",X"05",X"7E",X"E6",X"30",X"18",X"04",X"7E",X"2F",X"E6",X"30",X"FD",X"86",X"00",X"FD",
		X"77",X"00",X"23",X"C9",X"7A",X"D6",X"08",X"57",X"D5",X"E5",X"CD",X"40",X"08",X"E1",X"CD",X"AE",
		X"08",X"D1",X"7A",X"C6",X"10",X"57",X"30",X"05",X"23",X"23",X"23",X"18",X"0A",X"D5",X"E5",X"CD",
		X"40",X"08",X"E1",X"CD",X"AE",X"08",X"D1",X"7A",X"D6",X"08",X"57",X"C9",X"7B",X"C6",X"08",X"5F",
		X"CD",X"E4",X"08",X"7B",X"D6",X"10",X"5F",X"CD",X"E4",X"08",X"C9",X"CD",X"0C",X"09",X"7A",X"D6",
		X"10",X"57",X"E5",X"CD",X"40",X"08",X"E1",X"CD",X"AE",X"08",X"C9",X"D5",X"4F",X"E6",X"F0",X"0F",
		X"0F",X"0F",X"0F",X"47",X"21",X"F5",X"63",X"11",X"40",X"00",X"19",X"10",X"FD",X"D6",X"02",X"E5",
		X"5F",X"16",X"00",X"21",X"E8",X"63",X"19",X"7E",X"FE",X"10",X"38",X"08",X"E1",X"21",X"F5",X"63",
		X"0E",X"00",X"18",X"0C",X"34",X"87",X"87",X"5F",X"16",X"00",X"E1",X"19",X"79",X"E6",X"0F",X"4F",
		X"E5",X"FD",X"E1",X"FD",X"71",X"00",X"D1",X"C9",X"21",X"6F",X"09",X"DD",X"7E",X"02",X"DF",X"75",
		X"09",X"29",X"0A",X"EE",X"0A",X"21",X"2C",X"60",X"3A",X"00",X"60",X"CB",X"6F",X"28",X"03",X"21",
		X"2E",X"60",X"AF",X"01",X"01",X"04",X"D7",X"21",X"52",X"60",X"01",X"01",X"07",X"D7",X"CD",X"15",
		X"0E",X"CD",X"3C",X"0E",X"CD",X"E8",X"0E",X"3A",X"60",X"60",X"CB",X"7F",X"28",X"03",X"CD",X"F0",
		X"0E",X"3E",X"03",X"CD",X"A0",X"1B",X"CD",X"9F",X"3A",X"CD",X"EF",X"3A",X"CD",X"74",X"3F",X"CD",
		X"BA",X"3F",X"CD",X"4D",X"1E",X"CD",X"26",X"0F",X"CD",X"D6",X"32",X"CD",X"5E",X"29",X"DD",X"CB",
		X"00",X"C6",X"DD",X"36",X"04",X"80",X"21",X"00",X"02",X"22",X"52",X"60",X"EF",X"CD",X"FC",X"0A",
		X"3A",X"00",X"60",X"CB",X"7F",X"20",X"05",X"3A",X"0B",X"60",X"A7",X"C0",X"DD",X"E5",X"CD",X"73",
		X"3B",X"CD",X"53",X"1B",X"DD",X"E1",X"DD",X"35",X"04",X"20",X"E1",X"DD",X"CB",X"00",X"86",X"CD",
		X"51",X"1E",X"CD",X"7C",X"1B",X"EF",X"DD",X"E5",X"DD",X"21",X"DF",X"61",X"DD",X"36",X"00",X"80",
		X"CD",X"8A",X"07",X"DD",X"E1",X"06",X"01",X"CD",X"76",X"0F",X"3A",X"1B",X"6C",X"A7",X"20",X"F5",
		X"DD",X"36",X"02",X"02",X"CD",X"9D",X"23",X"21",X"00",X"02",X"22",X"52",X"60",X"21",X"80",X"80",
		X"22",X"30",X"60",X"3E",X"14",X"CD",X"86",X"0F",X"C9",X"3E",X"03",X"CD",X"A0",X"1B",X"CD",X"4D",
		X"1E",X"CD",X"26",X"0F",X"CD",X"9F",X"3A",X"CD",X"EF",X"3A",X"CD",X"74",X"3F",X"CD",X"BA",X"3F",
		X"DD",X"CB",X"00",X"C6",X"DD",X"36",X"04",X"80",X"21",X"00",X"02",X"22",X"52",X"60",X"EF",X"DD",
		X"E5",X"DD",X"21",X"DF",X"61",X"CD",X"8A",X"07",X"CD",X"73",X"3B",X"CD",X"53",X"1B",X"DD",X"E1",
		X"CD",X"FC",X"0A",X"DD",X"E5",X"DD",X"21",X"A9",X"63",X"DD",X"CB",X"00",X"7E",X"28",X"03",X"CD",
		X"25",X"19",X"DD",X"21",X"BE",X"63",X"DD",X"CB",X"00",X"7E",X"28",X"03",X"CD",X"25",X"19",X"DD",
		X"21",X"D3",X"63",X"DD",X"CB",X"00",X"7E",X"28",X"03",X"CD",X"25",X"19",X"DD",X"21",X"8D",X"63",
		X"DD",X"CB",X"00",X"7E",X"28",X"03",X"CD",X"DE",X"17",X"DD",X"E1",X"DD",X"35",X"04",X"20",X"AE",
		X"DD",X"CB",X"00",X"86",X"CD",X"7C",X"1B",X"06",X"5A",X"CD",X"76",X"0F",X"21",X"DF",X"61",X"36",
		X"80",X"CD",X"D6",X"32",X"CD",X"5E",X"29",X"21",X"00",X"02",X"22",X"52",X"60",X"CD",X"51",X"1E",
		X"CD",X"3A",X"33",X"3A",X"60",X"60",X"E6",X"0F",X"FE",X"0F",X"28",X"03",X"CD",X"9D",X"23",X"EF",
		X"DD",X"E5",X"DD",X"21",X"DF",X"61",X"DD",X"36",X"00",X"80",X"CD",X"8A",X"07",X"DD",X"E1",X"06",
		X"5A",X"CD",X"76",X"0F",X"DD",X"36",X"02",X"02",X"3E",X"14",X"CD",X"86",X"0F",X"C9",X"CD",X"6A",
		X"0F",X"C3",X"CA",X"0B",X"21",X"E8",X"61",X"CB",X"6E",X"C2",X"CA",X"0B",X"FD",X"21",X"59",X"60",
		X"2A",X"52",X"60",X"EB",X"2A",X"54",X"60",X"19",X"22",X"54",X"60",X"D5",X"CD",X"BD",X"0D",X"D1",
		X"2A",X"56",X"60",X"19",X"11",X"00",X"08",X"E5",X"AF",X"ED",X"52",X"30",X"07",X"E1",X"22",X"56",
		X"60",X"C3",X"CA",X"0B",X"D1",X"22",X"56",X"60",X"FD",X"7E",X"08",X"FD",X"BE",X"35",X"38",X"1B",
		X"CD",X"15",X"23",X"3A",X"60",X"60",X"E6",X"0F",X"FE",X"0F",X"20",X"12",X"DD",X"E5",X"DD",X"21",
		X"E8",X"61",X"06",X"18",X"CD",X"8D",X"1B",X"DD",X"E1",X"18",X"03",X"FD",X"34",X"08",X"CD",X"17",
		X"0C",X"CD",X"B2",X"23",X"CD",X"DD",X"29",X"21",X"69",X"60",X"7E",X"E6",X"0F",X"CA",X"CA",X"0B",
		X"7E",X"E6",X"F0",X"0F",X"0F",X"0F",X"5F",X"16",X"00",X"23",X"19",X"3A",X"61",X"60",X"BE",X"20",
		X"59",X"23",X"7E",X"47",X"E6",X"F0",X"0F",X"0F",X"0F",X"5F",X"16",X"00",X"21",X"E0",X"0B",X"19",
		X"CF",X"CF",X"3E",X"FF",X"BD",X"28",X"3B",X"CB",X"7E",X"28",X"03",X"EB",X"18",X"F3",X"78",X"E6",
		X"F0",X"FE",X"60",X"CA",X"B8",X"0B",X"DD",X"CB",X"00",X"46",X"20",X"2F",X"FE",X"20",X"20",X"18",
		X"E5",X"21",X"35",X"60",X"3A",X"00",X"60",X"CB",X"6F",X"28",X"03",X"21",X"43",X"60",X"34",X"5E",
		X"16",X"00",X"19",X"7E",X"A7",X"E1",X"28",X"0A",X"CB",X"FE",X"11",X"03",X"00",X"19",X"78",X"E6",
		X"0F",X"77",X"21",X"69",X"60",X"7E",X"3D",X"C6",X"10",X"77",X"C9",X"78",X"E6",X"F0",X"FE",X"70",
		X"C2",X"C2",X"0B",X"06",X"03",X"C3",X"B8",X"0B",X"00",X"02",X"80",X"00",X"03",X"00",X"FD",X"FF",
		X"00",X"00",X"F2",X"0B",X"F7",X"0B",X"FC",X"0B",X"FF",X"0B",X"04",X"0C",X"09",X"0C",X"0E",X"0C",
		X"15",X"0C",X"D6",X"62",X"EC",X"62",X"FF",X"02",X"63",X"11",X"63",X"FF",X"20",X"63",X"FF",X"47",
		X"63",X"58",X"63",X"FF",X"69",X"63",X"7B",X"63",X"FF",X"8D",X"63",X"9B",X"63",X"FF",X"A9",X"63",
		X"BE",X"63",X"D3",X"63",X"FF",X"FF",X"FF",X"FD",X"21",X"59",X"60",X"3A",X"55",X"60",X"CB",X"3F",
		X"CB",X"3F",X"CB",X"3F",X"5F",X"16",X"00",X"21",X"00",X"D3",X"19",X"CD",X"26",X"23",X"01",X"E0",
		X"FF",X"09",X"FD",X"36",X"FF",X"10",X"FD",X"7E",X"21",X"FE",X"13",X"28",X"08",X"1E",X"FD",X"CD",
		X"9F",X"0D",X"57",X"F7",X"09",X"E5",X"FD",X"6E",X"27",X"FD",X"66",X"28",X"7E",X"23",X"FD",X"75",
		X"27",X"FD",X"74",X"28",X"E1",X"47",X"CB",X"38",X"CB",X"38",X"CB",X"38",X"CB",X"38",X"28",X"0C",
		X"F7",X"C5",X"01",X"E0",X"FF",X"09",X"C1",X"FD",X"35",X"FF",X"10",X"F4",X"E6",X"0F",X"28",X"27",
		X"47",X"FD",X"5E",X"22",X"FD",X"56",X"23",X"CD",X"9F",X"0D",X"D5",X"CB",X"22",X"CB",X"22",X"CB",
		X"22",X"82",X"57",X"F7",X"C5",X"01",X"E0",X"FF",X"09",X"C1",X"FD",X"35",X"FF",X"D1",X"13",X"10",
		X"E6",X"FD",X"73",X"22",X"FD",X"72",X"23",X"E5",X"21",X"90",X"60",X"3A",X"8F",X"60",X"5F",X"16",
		X"00",X"19",X"EB",X"FD",X"6E",X"24",X"FD",X"66",X"25",X"01",X"04",X"00",X"ED",X"B0",X"FD",X"75",
		X"24",X"FD",X"74",X"25",X"E1",X"FD",X"35",X"26",X"20",X"08",X"E5",X"FD",X"35",X"1E",X"C4",X"E8",
		X"0E",X"E1",X"FD",X"CB",X"07",X"7E",X"20",X"23",X"1E",X"24",X"FD",X"56",X"01",X"01",X"E0",X"FF",
		X"F7",X"09",X"FD",X"35",X"FF",X"20",X"F9",X"21",X"10",X"61",X"3A",X"8F",X"60",X"5F",X"16",X"00",
		X"19",X"AF",X"06",X"04",X"77",X"23",X"10",X"FC",X"C3",X"8E",X"0D",X"E5",X"FD",X"6E",X"33",X"FD",
		X"66",X"34",X"7E",X"23",X"FD",X"75",X"33",X"FD",X"74",X"34",X"E1",X"47",X"CB",X"38",X"CB",X"38",
		X"CB",X"38",X"CB",X"38",X"E6",X"0F",X"4F",X"80",X"FD",X"96",X"FF",X"ED",X"44",X"C5",X"47",X"1E",
		X"24",X"CD",X"9F",X"0D",X"57",X"F7",X"C5",X"01",X"E0",X"FF",X"09",X"C1",X"FD",X"35",X"FF",X"10",
		X"F0",X"C1",X"78",X"A7",X"28",X"28",X"C5",X"FD",X"5E",X"2E",X"FD",X"56",X"2F",X"CD",X"9F",X"0D",
		X"D5",X"CB",X"22",X"CB",X"22",X"CB",X"22",X"82",X"57",X"F7",X"C5",X"01",X"E0",X"FF",X"09",X"C1",
		X"FD",X"35",X"FF",X"D1",X"13",X"10",X"E6",X"FD",X"73",X"2E",X"FD",X"72",X"2F",X"C1",X"79",X"A7",
		X"28",X"15",X"41",X"1E",X"FE",X"CD",X"9F",X"0D",X"57",X"F7",X"C5",X"01",X"E0",X"FF",X"09",X"C1",
		X"FD",X"35",X"FF",X"28",X"02",X"10",X"F2",X"21",X"10",X"61",X"3A",X"8F",X"60",X"5F",X"16",X"00",
		X"19",X"EB",X"FD",X"6E",X"30",X"FD",X"66",X"31",X"01",X"04",X"00",X"ED",X"B0",X"FD",X"75",X"30",
		X"FD",X"74",X"31",X"FD",X"35",X"32",X"20",X"06",X"FD",X"35",X"2A",X"C4",X"F0",X"0E",X"3A",X"8F",
		X"60",X"C6",X"04",X"FE",X"80",X"38",X"01",X"AF",X"32",X"8F",X"60",X"32",X"8F",X"60",X"C9",X"FD",
		X"7E",X"21",X"FE",X"10",X"28",X"08",X"FE",X"13",X"28",X"08",X"FD",X"7E",X"01",X"C9",X"FD",X"7E",
		X"03",X"C9",X"3E",X"03",X"C9",X"AF",X"06",X"18",X"21",X"E5",X"0D",X"18",X"20",X"06",X"13",X"3A",
		X"00",X"60",X"CB",X"6F",X"28",X"07",X"3A",X"02",X"90",X"CB",X"5F",X"20",X"08",X"21",X"E9",X"0D",
		X"3A",X"55",X"60",X"18",X"08",X"21",X"E9",X"0D",X"3A",X"55",X"60",X"ED",X"44",X"5E",X"23",X"56",
		X"23",X"12",X"10",X"F9",X"C9",X"01",X"D0",X"21",X"D0",X"41",X"D0",X"61",X"D0",X"02",X"D0",X"22",
		X"D0",X"42",X"D0",X"62",X"D0",X"03",X"D0",X"23",X"D0",X"43",X"D0",X"63",X"D0",X"04",X"D0",X"24",
		X"D0",X"44",X"D0",X"64",X"D0",X"05",X"D0",X"25",X"D0",X"45",X"D0",X"65",X"D0",X"06",X"D0",X"26",
		X"D0",X"46",X"D0",X"66",X"D0",X"FD",X"E5",X"FD",X"21",X"59",X"60",X"FD",X"5E",X"00",X"1D",X"CB",
		X"23",X"16",X"00",X"21",X"40",X"50",X"19",X"CF",X"11",X"5A",X"60",X"01",X"04",X"00",X"ED",X"B0",
		X"FD",X"75",X"05",X"FD",X"74",X"06",X"FD",X"E1",X"CD",X"07",X"11",X"C9",X"FD",X"E5",X"FD",X"21",
		X"59",X"60",X"FD",X"6E",X"05",X"FD",X"66",X"06",X"7E",X"FD",X"77",X"07",X"23",X"06",X"3F",X"CB",
		X"6F",X"28",X"02",X"06",X"1F",X"E6",X"0F",X"FE",X"0F",X"20",X"02",X"06",X"A0",X"FD",X"70",X"35",
		X"FD",X"36",X"08",X"00",X"7E",X"FD",X"77",X"1D",X"23",X"7E",X"FD",X"77",X"29",X"23",X"7E",X"FD",
		X"77",X"10",X"23",X"A7",X"28",X"09",X"87",X"4F",X"06",X"00",X"11",X"6A",X"60",X"ED",X"B0",X"FD",
		X"75",X"05",X"FD",X"74",X"06",X"FD",X"5E",X"1D",X"CB",X"23",X"16",X"00",X"21",X"6A",X"53",X"19",
		X"CF",X"FD",X"CB",X"07",X"6E",X"28",X"26",X"23",X"11",X"62",X"60",X"01",X"03",X"00",X"ED",X"B0",
		X"7E",X"FD",X"77",X"1E",X"23",X"FD",X"75",X"1F",X"FD",X"74",X"20",X"5F",X"16",X"00",X"19",X"7E",
		X"FD",X"77",X"2A",X"23",X"FD",X"75",X"2B",X"FD",X"74",X"2C",X"C3",X"E5",X"0E",X"7E",X"FD",X"77",
		X"1E",X"23",X"FD",X"75",X"1F",X"FD",X"74",X"20",X"FD",X"CB",X"07",X"7E",X"28",X"17",X"FD",X"5E",
		X"29",X"CB",X"23",X"16",X"00",X"21",X"6A",X"53",X"19",X"CF",X"7E",X"FD",X"77",X"2A",X"23",X"FD",
		X"75",X"2B",X"FD",X"74",X"2C",X"FD",X"E1",X"C9",X"FD",X"E5",X"FD",X"21",X"59",X"60",X"18",X"06",
		X"FD",X"E5",X"FD",X"21",X"65",X"60",X"FD",X"6E",X"1F",X"FD",X"66",X"20",X"7E",X"FD",X"77",X"21",
		X"23",X"FD",X"75",X"1F",X"FD",X"74",X"20",X"87",X"5F",X"16",X"00",X"21",X"72",X"54",X"19",X"CF",
		X"11",X"22",X"00",X"FD",X"19",X"FD",X"E5",X"D1",X"01",X"05",X"00",X"ED",X"B0",X"FD",X"75",X"05",
		X"FD",X"74",X"06",X"FD",X"E1",X"C9",X"3E",X"FF",X"21",X"C0",X"D0",X"01",X"01",X"20",X"D7",X"C9",
		X"00",X"CD",X"47",X"0F",X"21",X"90",X"60",X"19",X"7E",X"C6",X"48",X"C9",X"CD",X"47",X"0F",X"21",
		X"10",X"61",X"19",X"3E",X"C8",X"96",X"C9",X"5F",X"E6",X"F8",X"57",X"3A",X"55",X"60",X"E6",X"F8",
		X"82",X"CB",X"3F",X"57",X"7B",X"E6",X"07",X"CB",X"3F",X"82",X"CB",X"BF",X"5F",X"16",X"00",X"C9",
		X"21",X"52",X"60",X"5E",X"23",X"56",X"CD",X"4B",X"1F",X"C9",X"21",X"E2",X"61",X"CB",X"66",X"C0",
		X"E1",X"23",X"23",X"23",X"E5",X"C9",X"DD",X"E5",X"C5",X"EF",X"CD",X"73",X"3B",X"CD",X"B5",X"01",
		X"C1",X"10",X"F5",X"DD",X"E1",X"C9",X"5F",X"FE",X"00",X"28",X"06",X"3A",X"00",X"60",X"CB",X"7F",
		X"C8",X"16",X"00",X"21",X"06",X"6C",X"19",X"7B",X"FE",X"14",X"CA",X"B0",X"0F",X"FE",X"10",X"30",
		X"03",X"36",X"01",X"C9",X"D6",X"10",X"E5",X"5F",X"21",X"B6",X"0F",X"19",X"7E",X"E1",X"77",X"C9",
		X"36",X"01",X"CD",X"C8",X"0F",X"C9",X"C1",X"91",X"81",X"C1",X"A1",X"B1",X"A1",X"31",X"5F",X"16",
		X"00",X"21",X"06",X"6C",X"19",X"CB",X"D6",X"C9",X"2A",X"52",X"60",X"CB",X"25",X"CB",X"14",X"CB",
		X"25",X"CB",X"14",X"7C",X"FE",X"09",X"38",X"02",X"3E",X"08",X"6F",X"26",X"00",X"11",X"EB",X"0F",
		X"19",X"3A",X"1A",X"6C",X"E6",X"0F",X"86",X"32",X"1A",X"6C",X"C9",X"70",X"80",X"90",X"A0",X"B0",
		X"C0",X"D0",X"E0",X"F0",X"85",X"DD",X"CB",X"00",X"6E",X"C2",X"4A",X"10",X"DD",X"CB",X"00",X"EE",
		X"DD",X"36",X"01",X"3C",X"DD",X"36",X"02",X"01",X"DD",X"7E",X"03",X"E6",X"03",X"DD",X"77",X"03",
		X"87",X"4F",X"87",X"81",X"4F",X"06",X"00",X"11",X"04",X"00",X"DD",X"E5",X"E1",X"19",X"EB",X"21",
		X"E3",X"10",X"ED",X"B0",X"3A",X"59",X"60",X"3D",X"DD",X"77",X"08",X"DD",X"77",X"0E",X"DD",X"77",
		X"14",X"5F",X"16",X"00",X"21",X"01",X"11",X"19",X"7E",X"DD",X"77",X"09",X"DD",X"77",X"0F",X"DD",
		X"77",X"15",X"3E",X"0A",X"CD",X"86",X"0F",X"C3",X"CC",X"10",X"CD",X"6A",X"0F",X"C3",X"CC",X"10",
		X"DD",X"7E",X"01",X"A7",X"28",X"03",X"DD",X"35",X"01",X"21",X"00",X"02",X"C3",X"7A",X"10",X"DD",
		X"7E",X"02",X"A7",X"20",X"08",X"2A",X"52",X"60",X"CD",X"43",X"1F",X"18",X"0D",X"21",X"40",X"00",
		X"FE",X"02",X"20",X"03",X"21",X"80",X"FF",X"CD",X"F9",X"22",X"EB",X"DD",X"6E",X"04",X"DD",X"66",
		X"05",X"19",X"DD",X"7E",X"01",X"A7",X"20",X"0F",X"7C",X"FE",X"08",X"38",X"04",X"FE",X"F8",X"38",
		X"06",X"06",X"16",X"CD",X"8D",X"1B",X"C9",X"DD",X"75",X"04",X"DD",X"74",X"05",X"DD",X"46",X"03",
		X"05",X"28",X"0F",X"DD",X"75",X"0A",X"DD",X"74",X"0B",X"05",X"28",X"06",X"DD",X"75",X"10",X"DD",
		X"74",X"11",X"CD",X"46",X"33",X"FE",X"10",X"30",X"13",X"3E",X"C4",X"DD",X"46",X"03",X"D6",X"10",
		X"10",X"FC",X"47",X"3A",X"07",X"62",X"B8",X"38",X"03",X"CD",X"60",X"33",X"DD",X"E5",X"DD",X"46",
		X"03",X"C5",X"21",X"F5",X"10",X"CD",X"D1",X"07",X"11",X"06",X"00",X"DD",X"19",X"C1",X"10",X"F1",
		X"DD",X"E1",X"C9",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",
		X"00",X"00",X"A0",X"00",X"00",X"E0",X"01",X"E4",X"01",X"E8",X"01",X"EC",X"01",X"F0",X"01",X"F4",
		X"01",X"09",X"04",X"04",X"05",X"05",X"05",X"21",X"35",X"60",X"3A",X"00",X"60",X"CB",X"6F",X"28",
		X"03",X"21",X"43",X"60",X"01",X"01",X"0E",X"AF",X"D7",X"21",X"4C",X"11",X"3A",X"59",X"60",X"3D",
		X"87",X"5F",X"16",X"00",X"19",X"4E",X"23",X"46",X"11",X"36",X"60",X"3A",X"00",X"60",X"CB",X"6F",
		X"28",X"03",X"11",X"44",X"60",X"CD",X"13",X"1F",X"7D",X"E6",X"0F",X"91",X"30",X"FD",X"81",X"26",
		X"00",X"6F",X"19",X"7E",X"A7",X"20",X"EE",X"36",X"FF",X"10",X"EA",X"C9",X"02",X"01",X"06",X"03",
		X"04",X"02",X"0C",X"06",X"08",X"04",X"0D",X"07",X"DD",X"CB",X"00",X"6E",X"C2",X"96",X"11",X"DD",
		X"CB",X"00",X"EE",X"DD",X"E5",X"E1",X"11",X"04",X"00",X"19",X"EB",X"21",X"03",X"12",X"DD",X"7E",
		X"03",X"87",X"87",X"87",X"DD",X"86",X"03",X"4F",X"06",X"00",X"09",X"01",X"09",X"00",X"ED",X"B0",
		X"DD",X"36",X"0D",X"04",X"DD",X"36",X"0E",X"00",X"3E",X"02",X"CD",X"86",X"0F",X"DD",X"CB",X"00",
		X"F6",X"DD",X"36",X"01",X"2D",X"C9",X"DD",X"35",X"0C",X"20",X"06",X"06",X"0F",X"CD",X"8D",X"1B",
		X"C9",X"CD",X"46",X"33",X"FE",X"0E",X"30",X"0A",X"CD",X"53",X"33",X"FE",X"0E",X"30",X"03",X"CD",
		X"60",X"33",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"DD",X"5E",X"08",X"DD",X"56",X"09",X"19",X"DD",
		X"75",X"04",X"DD",X"74",X"05",X"DD",X"6E",X"06",X"DD",X"66",X"07",X"DD",X"5E",X"0A",X"DD",X"56",
		X"0B",X"19",X"DD",X"75",X"06",X"DD",X"74",X"07",X"DD",X"35",X"0D",X"20",X"07",X"DD",X"36",X"0D",
		X"04",X"DD",X"34",X"0E",X"21",X"27",X"12",X"11",X"0C",X"00",X"DD",X"CB",X"03",X"46",X"28",X"02",
		X"19",X"19",X"DD",X"CB",X"0E",X"46",X"28",X"01",X"19",X"DD",X"56",X"05",X"DD",X"5E",X"07",X"CD",
		X"0C",X"09",X"C9",X"00",X"F8",X"00",X"78",X"00",X"FC",X"00",X"00",X"3C",X"00",X"08",X"00",X"8A",
		X"00",X"04",X"00",X"00",X"3C",X"00",X"F8",X"00",X"C8",X"00",X"FC",X"00",X"FE",X"3C",X"00",X"08",
		X"00",X"C8",X"00",X"04",X"00",X"FE",X"3C",X"C0",X"01",X"01",X"C4",X"01",X"01",X"C8",X"01",X"01",
		X"CC",X"01",X"01",X"D0",X"01",X"01",X"D4",X"01",X"01",X"D8",X"01",X"01",X"DC",X"01",X"01",X"C4",
		X"01",X"21",X"C0",X"01",X"21",X"CC",X"01",X"21",X"C8",X"01",X"21",X"D4",X"01",X"21",X"D0",X"01",
		X"21",X"DC",X"01",X"21",X"D8",X"01",X"21",X"DD",X"CB",X"00",X"6E",X"C2",X"CB",X"12",X"DD",X"36",
		X"00",X"A0",X"21",X"80",X"01",X"DD",X"CB",X"03",X"56",X"28",X"07",X"DD",X"CB",X"00",X"E6",X"21",
		X"00",X"04",X"DD",X"75",X"11",X"DD",X"74",X"12",X"3E",X"01",X"DD",X"CB",X"03",X"46",X"28",X"01",
		X"3C",X"DD",X"77",X"02",X"3A",X"16",X"60",X"E6",X"07",X"5F",X"16",X"00",X"21",X"8E",X"14",X"19",
		X"7E",X"DD",X"77",X"0B",X"DD",X"36",X"0A",X"00",X"DD",X"46",X"02",X"0E",X"10",X"DD",X"CB",X"00",
		X"66",X"20",X"07",X"3E",X"FE",X"81",X"10",X"FD",X"18",X"02",X"3E",X"02",X"DD",X"77",X"05",X"DD",
		X"36",X"04",X"00",X"CD",X"31",X"0F",X"DD",X"86",X"0B",X"C6",X"08",X"DD",X"77",X"07",X"DD",X"36",
		X"08",X"01",X"DD",X"36",X"09",X"0C",X"3E",X"0C",X"CD",X"86",X"0F",X"CD",X"6A",X"0F",X"C3",X"4E",
		X"13",X"DD",X"4E",X"11",X"DD",X"46",X"12",X"DD",X"CB",X"00",X"66",X"28",X"07",X"C5",X"E1",X"CD",
		X"F9",X"22",X"18",X"03",X"CD",X"60",X"0F",X"DD",X"75",X"13",X"DD",X"74",X"14",X"DD",X"CB",X"00",
		X"66",X"20",X"03",X"CD",X"43",X"1F",X"DD",X"5E",X"04",X"DD",X"56",X"05",X"19",X"DD",X"75",X"04",
		X"DD",X"74",X"05",X"7C",X"DD",X"CB",X"00",X"5E",X"20",X"18",X"DD",X"CB",X"00",X"66",X"20",X"0A",
		X"FE",X"80",X"30",X"0E",X"FE",X"70",X"38",X"0A",X"18",X"04",X"FE",X"80",X"38",X"04",X"DD",X"CB",
		X"00",X"DE",X"3A",X"07",X"62",X"DD",X"BE",X"07",X"38",X"0C",X"DD",X"7E",X"07",X"FE",X"A0",X"30",
		X"0F",X"DD",X"34",X"0B",X"18",X"0A",X"DD",X"7E",X"0B",X"FE",X"20",X"38",X"03",X"DD",X"35",X"0B",
		X"DD",X"7E",X"05",X"CD",X"31",X"0F",X"DD",X"86",X"0B",X"C6",X"08",X"DD",X"77",X"07",X"DD",X"7E",
		X"02",X"DD",X"77",X"15",X"DD",X"36",X"16",X"00",X"DD",X"7E",X"05",X"CD",X"A6",X"14",X"C3",X"BE",
		X"13",X"DD",X"34",X"16",X"21",X"96",X"14",X"CD",X"D1",X"07",X"DD",X"56",X"05",X"DD",X"5E",X"07",
		X"DD",X"7E",X"0B",X"CD",X"D4",X"14",X"D5",X"DD",X"6E",X"0C",X"DD",X"66",X"0D",X"ED",X"5B",X"52",
		X"60",X"19",X"E5",X"11",X"00",X"08",X"AF",X"ED",X"52",X"E1",X"38",X"06",X"21",X"00",X"00",X"DD",
		X"34",X"0E",X"DD",X"75",X"0C",X"DD",X"74",X"0D",X"21",X"9A",X"14",X"DD",X"CB",X"0E",X"46",X"20",
		X"03",X"21",X"9D",X"14",X"D1",X"E5",X"CD",X"40",X"08",X"E1",X"CD",X"AE",X"08",X"CD",X"46",X"33",
		X"FE",X"0C",X"30",X"0A",X"CD",X"53",X"33",X"FE",X"0C",X"30",X"03",X"CD",X"60",X"33",X"DD",X"7E",
		X"05",X"DD",X"77",X"17",X"DD",X"E5",X"E1",X"11",X"19",X"00",X"19",X"DD",X"75",X"25",X"DD",X"74",
		X"26",X"DD",X"7E",X"17",X"D6",X"10",X"DD",X"77",X"17",X"CD",X"A6",X"14",X"C3",X"68",X"14",X"DD",
		X"34",X"16",X"DD",X"7E",X"17",X"CD",X"31",X"0F",X"DD",X"86",X"0B",X"C6",X"08",X"DD",X"77",X"18",
		X"DD",X"56",X"17",X"5F",X"CD",X"40",X"08",X"21",X"A3",X"14",X"CD",X"AE",X"08",X"DD",X"56",X"17",
		X"DD",X"5E",X"18",X"DD",X"7E",X"0B",X"CD",X"D4",X"14",X"D5",X"DD",X"6E",X"25",X"DD",X"66",X"26",
		X"E5",X"FD",X"E1",X"FD",X"6E",X"00",X"FD",X"66",X"01",X"ED",X"5B",X"52",X"60",X"19",X"E5",X"11",
		X"00",X"08",X"AF",X"ED",X"52",X"E1",X"38",X"06",X"21",X"00",X"00",X"FD",X"34",X"02",X"FD",X"75",
		X"00",X"FD",X"74",X"01",X"21",X"9A",X"14",X"FD",X"CB",X"02",X"46",X"28",X"03",X"21",X"9D",X"14",
		X"D1",X"E5",X"CD",X"40",X"08",X"E1",X"CD",X"AE",X"08",X"3A",X"05",X"62",X"DD",X"96",X"17",X"30",
		X"02",X"ED",X"44",X"FE",X"0C",X"30",X"11",X"3A",X"07",X"62",X"DD",X"96",X"18",X"30",X"02",X"ED",
		X"44",X"FE",X"0C",X"30",X"03",X"CD",X"60",X"33",X"DD",X"6E",X"25",X"DD",X"66",X"26",X"11",X"03",
		X"00",X"19",X"DD",X"75",X"25",X"DD",X"74",X"26",X"DD",X"35",X"15",X"C2",X"D1",X"13",X"DD",X"7E",
		X"16",X"A7",X"C0",X"06",X"27",X"CD",X"8D",X"1B",X"3E",X"0C",X"CD",X"BE",X"0F",X"C9",X"24",X"28",
		X"2C",X"30",X"34",X"38",X"3C",X"40",X"D0",X"00",X"D0",X"00",X"D8",X"00",X"06",X"DC",X"00",X"06",
		X"D4",X"00",X"06",X"D4",X"00",X"06",X"DD",X"CB",X"00",X"66",X"20",X"12",X"DD",X"CB",X"00",X"5E",
		X"20",X"06",X"FE",X"40",X"30",X"18",X"18",X"1B",X"FE",X"C0",X"38",X"12",X"18",X"15",X"DD",X"CB",
		X"00",X"5E",X"20",X"06",X"FE",X"C0",X"38",X"06",X"18",X"09",X"FE",X"40",X"38",X"05",X"E1",X"23",
		X"23",X"23",X"E5",X"C9",X"CD",X"C8",X"32",X"7B",X"D6",X"10",X"5F",X"78",X"A7",X"28",X"16",X"05",
		X"28",X"13",X"C5",X"D5",X"CD",X"40",X"08",X"21",X"86",X"32",X"CD",X"AE",X"08",X"D1",X"7B",X"D6",
		X"10",X"5F",X"C1",X"10",X"ED",X"79",X"A7",X"28",X"1B",X"D5",X"C5",X"3D",X"4F",X"87",X"81",X"4F",
		X"06",X"00",X"21",X"59",X"32",X"09",X"E5",X"CD",X"40",X"08",X"E1",X"CD",X"AE",X"08",X"C1",X"D1",
		X"7B",X"91",X"5F",X"14",X"C9",X"DD",X"CB",X"00",X"6E",X"C2",X"6B",X"15",X"DD",X"36",X"00",X"A0",
		X"DD",X"36",X"04",X"00",X"3E",X"F8",X"DD",X"77",X"05",X"CD",X"31",X"0F",X"C6",X"08",X"DD",X"77",
		X"07",X"DD",X"36",X"06",X"00",X"DD",X"36",X"08",X"00",X"DD",X"36",X"09",X"07",X"DD",X"7E",X"03",
		X"87",X"87",X"5F",X"16",X"00",X"21",X"3C",X"16",X"19",X"DD",X"E5",X"06",X"04",X"7E",X"DD",X"77",
		X"0A",X"23",X"DD",X"23",X"10",X"F7",X"DD",X"E1",X"DD",X"7E",X"0A",X"DD",X"77",X"0E",X"DD",X"7E",
		X"0B",X"DD",X"77",X"0F",X"DD",X"36",X"10",X"03",X"C3",X"0F",X"16",X"01",X"20",X"01",X"CD",X"60",
		X"0F",X"CD",X"43",X"1F",X"EB",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"19",X"DD",X"75",X"04",X"DD",
		X"74",X"05",X"7C",X"FE",X"08",X"30",X"06",X"06",X"11",X"CD",X"8D",X"1B",X"C9",X"DD",X"6E",X"0E",
		X"DD",X"66",X"0F",X"DD",X"5E",X"0C",X"DD",X"56",X"0D",X"DD",X"CB",X"00",X"66",X"C2",X"D0",X"15",
		X"AF",X"ED",X"52",X"38",X"1C",X"DD",X"75",X"0E",X"DD",X"74",X"0F",X"EB",X"DD",X"6E",X"06",X"DD",
		X"66",X"07",X"19",X"7C",X"FE",X"C0",X"30",X"09",X"DD",X"75",X"06",X"DD",X"74",X"07",X"C3",X"0F",
		X"16",X"DD",X"CB",X"00",X"E6",X"DD",X"36",X"0E",X"00",X"DD",X"36",X"0F",X"00",X"C3",X"0F",X"16",
		X"19",X"DD",X"75",X"0E",X"DD",X"74",X"0F",X"CD",X"43",X"1F",X"EB",X"DD",X"6E",X"06",X"DD",X"66",
		X"07",X"19",X"E5",X"DD",X"7E",X"05",X"CD",X"31",X"0F",X"E1",X"C6",X"08",X"BC",X"38",X"1A",X"67",
		X"2E",X"00",X"DD",X"CB",X"00",X"A6",X"E5",X"3E",X"0B",X"CD",X"86",X"0F",X"E1",X"DD",X"7E",X"0A",
		X"DD",X"77",X"0E",X"DD",X"7E",X"0B",X"DD",X"77",X"0F",X"DD",X"75",X"06",X"DD",X"74",X"07",X"CD",
		X"46",X"33",X"FE",X"0C",X"30",X"0A",X"CD",X"53",X"33",X"FE",X"0C",X"30",X"03",X"CD",X"60",X"33",
		X"DD",X"35",X"10",X"20",X"10",X"DD",X"36",X"10",X"03",X"DD",X"7E",X"08",X"3C",X"FE",X"08",X"38",
		X"01",X"AF",X"DD",X"77",X"08",X"21",X"44",X"16",X"CD",X"D1",X"07",X"C9",X"00",X"07",X"60",X"00",
		X"00",X"05",X"60",X"00",X"E0",X"00",X"E4",X"00",X"E0",X"20",X"F0",X"00",X"E0",X"00",X"E4",X"00",
		X"E0",X"20",X"F0",X"00",X"DD",X"CB",X"00",X"6E",X"C2",X"CF",X"16",X"DD",X"36",X"00",X"A0",X"DD",
		X"7E",X"03",X"E6",X"03",X"87",X"5F",X"16",X"00",X"21",X"B4",X"17",X"19",X"7E",X"DD",X"77",X"0A",
		X"23",X"7E",X"DD",X"77",X"0B",X"3E",X"F8",X"CD",X"31",X"0F",X"C6",X"18",X"DD",X"77",X"07",X"DD",
		X"36",X"06",X"00",X"DD",X"36",X"04",X"00",X"DD",X"36",X"05",X"F8",X"DD",X"36",X"08",X"00",X"DD",
		X"36",X"10",X"00",X"DD",X"36",X"11",X"00",X"DD",X"7E",X"03",X"E6",X"0C",X"CB",X"5F",X"20",X"04",
		X"DD",X"CB",X"00",X"E6",X"0F",X"0F",X"5F",X"16",X"00",X"21",X"BA",X"17",X"19",X"7E",X"DD",X"77",
		X"0E",X"DD",X"77",X"0F",X"3E",X"11",X"CD",X"86",X"0F",X"DD",X"56",X"05",X"DD",X"5E",X"07",X"21",
		X"C6",X"17",X"DD",X"CB",X"08",X"46",X"28",X"03",X"21",X"D2",X"17",X"CD",X"0C",X"09",X"C9",X"CD",
		X"6A",X"0F",X"C3",X"B9",X"16",X"DD",X"4E",X"0A",X"DD",X"46",X"0B",X"CD",X"60",X"0F",X"DD",X"75",
		X"0C",X"DD",X"74",X"0D",X"CD",X"43",X"1F",X"DD",X"5E",X"04",X"DD",X"56",X"05",X"19",X"DD",X"75",
		X"04",X"DD",X"74",X"05",X"7C",X"FE",X"08",X"30",X"13",X"06",X"12",X"CD",X"8D",X"1B",X"3A",X"69",
		X"63",X"21",X"7B",X"63",X"B6",X"C0",X"3E",X"11",X"CD",X"BE",X"0F",X"C9",X"DD",X"CB",X"00",X"66",
		X"28",X"1D",X"DD",X"35",X"0F",X"20",X"4C",X"DD",X"7E",X"0E",X"DD",X"77",X"0F",X"3A",X"07",X"62",
		X"DD",X"BE",X"07",X"30",X"05",X"DD",X"34",X"07",X"18",X"03",X"DD",X"35",X"07",X"18",X"34",X"21",
		X"00",X"01",X"DD",X"CB",X"00",X"56",X"28",X"03",X"CD",X"43",X"1F",X"DD",X"5E",X"06",X"DD",X"56",
		X"07",X"19",X"DD",X"75",X"06",X"DD",X"74",X"07",X"DD",X"35",X"0F",X"20",X"16",X"DD",X"7E",X"0E",
		X"DD",X"77",X"0F",X"DD",X"7E",X"00",X"DD",X"CB",X"00",X"96",X"2F",X"E6",X"04",X"DD",X"86",X"00",
		X"DD",X"77",X"00",X"DD",X"7E",X"07",X"FE",X"98",X"38",X"04",X"DD",X"36",X"07",X"98",X"DD",X"7E",
		X"05",X"CD",X"31",X"0F",X"C6",X"18",X"DD",X"BE",X"07",X"38",X"07",X"FE",X"98",X"30",X"03",X"DD",
		X"77",X"07",X"CD",X"46",X"33",X"FE",X"12",X"30",X"0A",X"CD",X"53",X"33",X"FE",X"12",X"30",X"03",
		X"CD",X"60",X"33",X"DD",X"6E",X"10",X"DD",X"66",X"11",X"DD",X"5E",X"0C",X"DD",X"56",X"0D",X"19",
		X"7C",X"FE",X"08",X"38",X"06",X"D6",X"08",X"67",X"DD",X"34",X"08",X"DD",X"75",X"10",X"DD",X"74",
		X"11",X"C3",X"B9",X"16",X"40",X"01",X"00",X"01",X"C0",X"00",X"0C",X"06",X"08",X"18",X"71",X"74",
		X"77",X"7A",X"7D",X"81",X"84",X"87",X"00",X"01",X"0B",X"04",X"01",X"0B",X"08",X"01",X"0B",X"0C",
		X"01",X"0B",X"10",X"01",X"0B",X"14",X"01",X"0B",X"18",X"01",X"0B",X"1C",X"01",X"0B",X"DD",X"CB",
		X"00",X"6E",X"20",X"23",X"DD",X"36",X"00",X"A0",X"DD",X"36",X"04",X"00",X"DD",X"36",X"05",X"20",
		X"DD",X"36",X"06",X"00",X"DD",X"36",X"07",X"58",X"DD",X"36",X"02",X"00",X"DD",X"36",X"0D",X"50",
		X"DD",X"36",X"08",X"01",X"C3",X"14",X"18",X"DD",X"7E",X"02",X"21",X"0E",X"18",X"DF",X"14",X"18",
		X"14",X"18",X"14",X"18",X"CD",X"6A",X"0F",X"C3",X"5C",X"18",X"DD",X"6E",X"04",X"DD",X"66",X"05",
		X"ED",X"5B",X"52",X"60",X"AF",X"ED",X"52",X"DD",X"75",X"04",X"DD",X"74",X"05",X"7C",X"FE",X"80",
		X"38",X"07",X"DD",X"CB",X"00",X"C6",X"C3",X"4B",X"18",X"DD",X"CB",X"00",X"46",X"CA",X"4B",X"18",
		X"FE",X"08",X"D2",X"4B",X"18",X"06",X"0E",X"CD",X"8D",X"1B",X"C9",X"CD",X"46",X"33",X"FE",X"14",
		X"30",X"0A",X"CD",X"53",X"33",X"FE",X"14",X"30",X"03",X"CD",X"60",X"33",X"DD",X"7E",X"09",X"A7",
		X"28",X"05",X"DD",X"35",X"09",X"18",X"2C",X"DD",X"34",X"08",X"21",X"E3",X"18",X"DD",X"7E",X"08",
		X"FE",X"04",X"38",X"04",X"AF",X"DD",X"77",X"08",X"5F",X"16",X"00",X"21",X"19",X"19",X"19",X"7E",
		X"DD",X"77",X"09",X"C3",X"A9",X"18",X"CB",X"23",X"21",X"1D",X"19",X"19",X"CF",X"DD",X"75",X"0A",
		X"DD",X"74",X"0B",X"C3",X"A9",X"18",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"DD",X"5E",X"0A",X"DD",
		X"56",X"0B",X"19",X"DD",X"75",X"04",X"DD",X"74",X"05",X"DD",X"CB",X"00",X"46",X"28",X"18",X"DD",
		X"7E",X"08",X"07",X"07",X"5F",X"07",X"83",X"5F",X"16",X"00",X"21",X"E3",X"18",X"19",X"DD",X"56",
		X"05",X"DD",X"5E",X"07",X"CD",X"0C",X"09",X"DD",X"7E",X"05",X"DD",X"CB",X"00",X"46",X"28",X"03",
		X"FE",X"28",X"D8",X"D6",X"20",X"DD",X"77",X"0C",X"57",X"DD",X"5E",X"0D",X"21",X"13",X"19",X"CD",
		X"E4",X"08",X"C9",X"24",X"01",X"2E",X"20",X"01",X"2E",X"2C",X"01",X"2E",X"28",X"01",X"2E",X"34",
		X"01",X"2E",X"30",X"01",X"2E",X"3C",X"01",X"2E",X"38",X"01",X"2E",X"44",X"01",X"2E",X"40",X"01",
		X"2E",X"4C",X"01",X"2E",X"48",X"01",X"2E",X"34",X"01",X"2E",X"30",X"01",X"2E",X"3C",X"01",X"2E",
		X"38",X"01",X"2E",X"50",X"01",X"00",X"54",X"01",X"00",X"04",X"04",X"04",X"04",X"C0",X"FF",X"00",
		X"00",X"40",X"00",X"00",X"00",X"DD",X"CB",X"00",X"6E",X"C2",X"8D",X"19",X"DD",X"CB",X"00",X"EE",
		X"DD",X"36",X"02",X"00",X"3A",X"18",X"6C",X"A7",X"20",X"05",X"3E",X"12",X"CD",X"86",X"0F",X"DD",
		X"E5",X"21",X"0A",X"1B",X"06",X"0C",X"7E",X"DD",X"77",X"04",X"23",X"DD",X"23",X"10",X"F7",X"DD",
		X"E1",X"DD",X"7E",X"03",X"E6",X"03",X"FE",X"03",X"20",X"07",X"DD",X"36",X"02",X"04",X"C3",X"40",
		X"1A",X"5F",X"16",X"00",X"21",X"18",X"1B",X"19",X"7E",X"DD",X"77",X"10",X"87",X"DD",X"77",X"12",
		X"DD",X"7E",X"03",X"E6",X"0C",X"0F",X"0F",X"5F",X"16",X"00",X"21",X"1A",X"1B",X"19",X"7E",X"DD",
		X"77",X"11",X"DD",X"36",X"13",X"00",X"DD",X"36",X"14",X"00",X"C3",X"BE",X"19",X"DD",X"7E",X"02",
		X"FE",X"05",X"CA",X"1C",X"1B",X"CD",X"6A",X"0F",X"C3",X"40",X"1A",X"DD",X"CB",X"00",X"66",X"C2",
		X"BE",X"19",X"21",X"A9",X"19",X"DD",X"7E",X"02",X"DF",X"B5",X"19",X"70",X"1A",X"B7",X"1A",X"C3",
		X"1A",X"BE",X"19",X"1C",X"1B",X"DD",X"35",X"12",X"20",X"04",X"DD",X"36",X"02",X"01",X"21",X"E8",
		X"61",X"CB",X"6E",X"C2",X"40",X"1A",X"2A",X"52",X"60",X"CD",X"43",X"1F",X"EB",X"DD",X"6E",X"04",
		X"DD",X"66",X"05",X"19",X"DD",X"75",X"04",X"DD",X"74",X"05",X"DD",X"CB",X"00",X"5E",X"20",X"09",
		X"7C",X"FE",X"80",X"30",X"04",X"DD",X"CB",X"00",X"DE",X"DD",X"6E",X"0A",X"DD",X"66",X"0B",X"19",
		X"DD",X"75",X"0A",X"DD",X"74",X"0B",X"DD",X"CB",X"00",X"5E",X"28",X"1C",X"7C",X"FE",X"10",X"30",
		X"17",X"06",X"15",X"CD",X"8D",X"1B",X"3A",X"A9",X"63",X"21",X"BE",X"63",X"B6",X"21",X"D3",X"63",
		X"B6",X"C0",X"3E",X"12",X"CD",X"BE",X"0F",X"C9",X"DD",X"7E",X"0B",X"DD",X"96",X"05",X"FE",X"20",
		X"38",X"1E",X"3A",X"05",X"62",X"47",X"DD",X"7E",X"05",X"C6",X"10",X"B8",X"30",X"12",X"DD",X"7E",
		X"0B",X"D6",X"10",X"B8",X"38",X"0A",X"21",X"00",X"62",X"CB",X"EE",X"21",X"03",X"62",X"36",X"09",
		X"DD",X"CB",X"00",X"5E",X"28",X"07",X"DD",X"7E",X"05",X"FE",X"E0",X"30",X"06",X"21",X"16",X"1B",
		X"CD",X"D1",X"07",X"DD",X"CB",X"00",X"5E",X"20",X"07",X"DD",X"7E",X"0B",X"FE",X"20",X"38",X"0F",
		X"DD",X"E5",X"11",X"06",X"00",X"DD",X"19",X"21",X"16",X"1B",X"CD",X"D1",X"07",X"DD",X"E1",X"C9",
		X"DD",X"6E",X"13",X"DD",X"66",X"14",X"E5",X"11",X"00",X"10",X"AF",X"ED",X"52",X"E1",X"38",X"0D",
		X"DD",X"36",X"02",X"02",X"DD",X"7E",X"11",X"DD",X"77",X"12",X"C3",X"BE",X"19",X"11",X"80",X"00",
		X"19",X"DD",X"75",X"13",X"DD",X"74",X"14",X"DD",X"6E",X"0A",X"DD",X"66",X"0B",X"19",X"DD",X"75",
		X"0A",X"DD",X"74",X"0B",X"11",X"80",X"FF",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"19",X"DD",X"75",
		X"04",X"DD",X"74",X"05",X"C3",X"BE",X"19",X"DD",X"35",X"12",X"20",X"04",X"DD",X"36",X"02",X"03",
		X"C3",X"BE",X"19",X"DD",X"7E",X"14",X"A7",X"28",X"04",X"CB",X"7F",X"28",X"0D",X"DD",X"36",X"02",
		X"00",X"DD",X"7E",X"10",X"DD",X"77",X"12",X"C3",X"BE",X"19",X"11",X"80",X"00",X"DD",X"6E",X"04",
		X"DD",X"66",X"05",X"19",X"DD",X"75",X"04",X"DD",X"74",X"05",X"11",X"80",X"FF",X"DD",X"6E",X"0A",
		X"DD",X"66",X"0B",X"19",X"DD",X"75",X"0A",X"DD",X"74",X"0B",X"DD",X"6E",X"13",X"DD",X"66",X"14",
		X"19",X"DD",X"75",X"13",X"DD",X"74",X"14",X"C3",X"BE",X"19",X"00",X"F7",X"00",X"63",X"00",X"08",
		X"00",X"07",X"00",X"63",X"00",X"08",X"EC",X"00",X"05",X"0F",X"03",X"05",X"DD",X"5E",X"13",X"DD",
		X"56",X"14",X"7A",X"A7",X"CA",X"48",X"1B",X"CB",X"7F",X"C2",X"48",X"1B",X"DD",X"6E",X"04",X"DD",
		X"66",X"05",X"19",X"DD",X"75",X"04",X"DD",X"74",X"05",X"DD",X"6E",X"0A",X"DD",X"66",X"0B",X"AF",
		X"ED",X"52",X"DD",X"75",X"0A",X"DD",X"74",X"0B",X"DD",X"CB",X"00",X"E6",X"DD",X"36",X"02",X"04",
		X"C3",X"40",X"1A",X"3A",X"D5",X"61",X"CB",X"7F",X"C0",X"21",X"19",X"60",X"34",X"4E",X"21",X"51",
		X"1D",X"3A",X"00",X"60",X"CB",X"6F",X"28",X"03",X"21",X"57",X"1D",X"CB",X"51",X"20",X"05",X"CD",
		X"39",X"1D",X"18",X"07",X"CF",X"3E",X"24",X"01",X"01",X"03",X"D7",X"C9",X"21",X"51",X"1D",X"3A",
		X"00",X"60",X"CB",X"6F",X"28",X"03",X"21",X"57",X"1D",X"CD",X"39",X"1D",X"C9",X"DD",X"E5",X"E1",
		X"0E",X"01",X"AF",X"D7",X"C9",X"AF",X"77",X"23",X"E5",X"ED",X"52",X"E1",X"C8",X"38",X"F6",X"C9",
		X"F5",X"CD",X"B2",X"1B",X"CD",X"C9",X"1B",X"CD",X"B5",X"0D",X"F1",X"CD",X"E1",X"1B",X"CD",X"DF",
		X"1C",X"C9",X"21",X"E8",X"63",X"01",X"05",X"0C",X"AF",X"D7",X"EF",X"06",X"00",X"11",X"04",X"00",
		X"21",X"00",X"70",X"AF",X"77",X"19",X"10",X"FC",X"C9",X"21",X"80",X"D0",X"01",X"03",X"00",X"3E",
		X"24",X"D7",X"21",X"80",X"D4",X"01",X"00",X"03",X"CB",X"9E",X"23",X"0B",X"78",X"B1",X"20",X"F8",
		X"C9",X"87",X"5F",X"16",X"00",X"21",X"FC",X"1B",X"19",X"CF",X"11",X"80",X"D4",X"7E",X"A7",X"C8",
		X"47",X"23",X"4E",X"23",X"EB",X"71",X"23",X"10",X"FC",X"EB",X"18",X"F1",X"06",X"1C",X"25",X"1C",
		X"5E",X"1C",X"81",X"1C",X"9C",X"1C",X"13",X"00",X"04",X"02",X"09",X"03",X"03",X"01",X"07",X"00",
		X"09",X"01",X"04",X"02",X"09",X"03",X"80",X"02",X"80",X"02",X"A0",X"02",X"A0",X"03",X"08",X"01",
		X"18",X"03",X"60",X"00",X"00",X"13",X"00",X"04",X"02",X"09",X"03",X"03",X"01",X"07",X"00",X"09",
		X"01",X"04",X"02",X"09",X"03",X"40",X"00",X"08",X"00",X"08",X"03",X"30",X"00",X"08",X"02",X"08",
		X"03",X"30",X"02",X"08",X"04",X"08",X"03",X"30",X"04",X"08",X"05",X"08",X"03",X"30",X"05",X"08",
		X"06",X"08",X"03",X"30",X"06",X"C0",X"00",X"08",X"01",X"18",X"03",X"60",X"00",X"00",X"13",X"00",
		X"04",X"02",X"09",X"03",X"03",X"01",X"07",X"00",X"09",X"01",X"04",X"02",X"09",X"03",X"C0",X"05",
		X"80",X"00",X"80",X"02",X"12",X"05",X"0E",X"03",X"60",X"00",X"08",X"01",X"18",X"03",X"60",X"00",
		X"00",X"13",X"00",X"04",X"02",X"09",X"03",X"03",X"01",X"07",X"00",X"09",X"01",X"04",X"02",X"09",
		X"03",X"20",X"06",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"60",X"03",X"00",X"13",X"00",X"04",X"02",
		X"09",X"03",X"03",X"01",X"07",X"00",X"09",X"01",X"04",X"02",X"09",X"03",X"40",X"00",X"08",X"00",
		X"08",X"03",X"30",X"00",X"08",X"02",X"08",X"03",X"30",X"02",X"08",X"04",X"08",X"03",X"30",X"04",
		X"08",X"05",X"08",X"03",X"30",X"05",X"08",X"06",X"08",X"03",X"30",X"06",X"3C",X"00",X"04",X"01",
		X"3C",X"00",X"04",X"01",X"3C",X"00",X"04",X"01",X"3C",X"00",X"04",X"03",X"40",X"00",X"00",X"21",
		X"46",X"1D",X"CD",X"39",X"1D",X"CD",X"39",X"1D",X"DD",X"E5",X"DD",X"21",X"94",X"6A",X"06",X"06",
		X"21",X"AB",X"D0",X"CD",X"95",X"1E",X"DD",X"21",X"0C",X"60",X"06",X"06",X"21",X"97",X"D0",X"CD",
		X"95",X"1E",X"CD",X"4D",X"1E",X"3A",X"00",X"60",X"CB",X"7F",X"20",X"11",X"21",X"5D",X"1D",X"CD",
		X"39",X"1D",X"CD",X"33",X"1E",X"21",X"A9",X"1D",X"CD",X"39",X"1D",X"18",X"07",X"3A",X"00",X"60",
		X"CB",X"77",X"28",X"12",X"21",X"57",X"1D",X"CD",X"39",X"1D",X"DD",X"21",X"0F",X"60",X"06",X"06",
		X"21",X"B7",X"D0",X"CD",X"95",X"1E",X"DD",X"E1",X"C9",X"5E",X"23",X"56",X"23",X"46",X"23",X"7E",
		X"12",X"13",X"23",X"10",X"FA",X"C9",X"8A",X"D0",X"08",X"11",X"12",X"2D",X"1C",X"0C",X"18",X"1B",
		X"0E",X"93",X"D0",X"03",X"01",X"1C",X"1D",X"B3",X"D0",X"03",X"02",X"17",X"0D",X"02",X"D3",X"06",
		X"0C",X"1B",X"0E",X"0D",X"12",X"1D",X"46",X"D1",X"0A",X"15",X"0E",X"1D",X"3B",X"1C",X"24",X"19",
		X"15",X"0A",X"22",X"E7",X"D1",X"11",X"19",X"1E",X"1C",X"11",X"24",X"1C",X"1D",X"0A",X"1B",X"1D",
		X"24",X"0B",X"1E",X"1D",X"1D",X"18",X"17",X"48",X"D2",X"0E",X"24",X"18",X"17",X"15",X"22",X"24",
		X"01",X"24",X"19",X"15",X"0A",X"22",X"0E",X"1B",X"48",X"D2",X"0E",X"01",X"24",X"18",X"1B",X"24",
		X"02",X"24",X"19",X"15",X"0A",X"22",X"0E",X"1B",X"1C",X"4A",X"D3",X"0B",X"3A",X"24",X"1E",X"17",
		X"12",X"1F",X"0E",X"1B",X"1C",X"0A",X"15",X"24",X"6A",X"D1",X"09",X"10",X"0A",X"16",X"0E",X"24",
		X"18",X"1F",X"0E",X"1B",X"CB",X"D1",X"08",X"19",X"15",X"0A",X"22",X"0E",X"1B",X"24",X"01",X"CB",
		X"D1",X"08",X"19",X"15",X"0A",X"22",X"0E",X"1B",X"24",X"02",X"CB",X"D1",X"0F",X"0B",X"18",X"17",
		X"1E",X"1C",X"24",X"0C",X"11",X"0A",X"1B",X"0A",X"17",X"10",X"0E",X"28",X"0C",X"D2",X"0B",X"19",
		X"1E",X"1C",X"11",X"24",X"0B",X"1E",X"1D",X"1D",X"18",X"17",X"79",X"D2",X"03",X"19",X"1D",X"1C",
		X"EF",X"D1",X"08",X"17",X"18",X"24",X"0B",X"18",X"17",X"1E",X"1C",X"11",X"0B",X"D1",X"18",X"03",
		X"11",X"28",X"D1",X"3E",X"60",X"01",X"04",X"10",X"D5",X"12",X"D5",X"EB",X"11",X"00",X"04",X"19",
		X"36",X"02",X"D1",X"3C",X"13",X"10",X"F2",X"06",X"10",X"D1",X"21",X"20",X"00",X"19",X"EB",X"0D",
		X"20",X"E6",X"C9",X"3A",X"04",X"60",X"CD",X"27",X"1F",X"32",X"09",X"60",X"DD",X"E5",X"DD",X"21",
		X"09",X"60",X"06",X"02",X"21",X"09",X"D3",X"CD",X"95",X"1E",X"DD",X"E1",X"C9",X"06",X"00",X"18",
		X"02",X"06",X"01",X"21",X"17",X"60",X"3A",X"00",X"60",X"CB",X"6F",X"28",X"01",X"23",X"E5",X"7E",
		X"90",X"38",X"21",X"FE",X"06",X"38",X"02",X"3E",X"06",X"47",X"3E",X"06",X"90",X"4F",X"21",X"A3",
		X"D0",X"78",X"A7",X"28",X"05",X"36",X"3C",X"23",X"10",X"FB",X"79",X"A7",X"28",X"06",X"47",X"36",
		X"24",X"23",X"10",X"FB",X"E1",X"DD",X"E5",X"E5",X"DD",X"E1",X"06",X"02",X"21",X"A1",X"D0",X"CD",
		X"95",X"1E",X"DD",X"E1",X"C9",X"0E",X"00",X"DD",X"7E",X"00",X"CB",X"40",X"20",X"08",X"E6",X"F0",
		X"0F",X"0F",X"0F",X"0F",X"18",X"04",X"E6",X"0F",X"DD",X"23",X"A7",X"28",X"04",X"0E",X"FF",X"18",
		X"0E",X"CB",X"41",X"20",X"0A",X"78",X"FE",X"01",X"28",X"04",X"3E",X"24",X"18",X"01",X"AF",X"77",
		X"23",X"10",X"D4",X"C9",X"DD",X"E5",X"FD",X"E5",X"FD",X"21",X"00",X"60",X"FD",X"CB",X"00",X"7E",
		X"CA",X"02",X"1F",X"21",X"14",X"60",X"11",X"0E",X"60",X"FD",X"CB",X"00",X"6E",X"28",X"03",X"11",
		X"11",X"60",X"CD",X"07",X"1F",X"06",X"06",X"DD",X"21",X"0C",X"60",X"21",X"97",X"D0",X"FD",X"CB",
		X"00",X"6E",X"28",X"07",X"DD",X"21",X"0F",X"60",X"21",X"B7",X"D0",X"DD",X"E5",X"CD",X"95",X"1E",
		X"DD",X"E1",X"FD",X"E1",X"DD",X"E1",X"C9",X"AF",X"06",X"03",X"1A",X"8E",X"27",X"12",X"2B",X"1B",
		X"10",X"F8",X"C9",X"2A",X"15",X"60",X"7C",X"CB",X"25",X"CB",X"14",X"CB",X"BC",X"E6",X"60",X"E2",
		X"23",X"1F",X"23",X"22",X"15",X"60",X"C9",X"FE",X"64",X"38",X"04",X"D6",X"64",X"18",X"F8",X"01",
		X"00",X"0A",X"90",X"38",X"03",X"0C",X"18",X"FA",X"80",X"CB",X"21",X"CB",X"21",X"CB",X"21",X"CB",
		X"21",X"81",X"C9",X"7C",X"2F",X"67",X"7D",X"2F",X"6F",X"23",X"C9",X"D5",X"21",X"00",X"00",X"78",
		X"A7",X"28",X"0A",X"CB",X"18",X"30",X"01",X"19",X"EB",X"29",X"EB",X"18",X"F2",X"D1",X"CB",X"3A",
		X"CB",X"1B",X"79",X"A7",X"C8",X"CB",X"11",X"30",X"F5",X"19",X"18",X"F2",X"FD",X"21",X"00",X"00",
		X"11",X"00",X"01",X"78",X"B1",X"C8",X"AF",X"ED",X"42",X"38",X"04",X"FD",X"19",X"18",X"F7",X"09",
		X"CB",X"38",X"CB",X"19",X"78",X"B1",X"C8",X"CB",X"3A",X"CB",X"1B",X"D8",X"18",X"E8",X"C3",X"21",
		X"89",X"6A",X"01",X"01",X"0A",X"3E",X"24",X"D7",X"DD",X"E5",X"FD",X"E5",X"FD",X"21",X"94",X"6A",
		X"DD",X"21",X"0C",X"60",X"3A",X"00",X"60",X"CB",X"6F",X"28",X"04",X"DD",X"21",X"0F",X"60",X"01",
		X"00",X"05",X"DD",X"56",X"00",X"DD",X"5E",X"01",X"FD",X"66",X"00",X"FD",X"6E",X"01",X"AF",X"ED",
		X"52",X"20",X"08",X"FD",X"7E",X"02",X"DD",X"96",X"02",X"28",X"0E",X"38",X"0C",X"FD",X"23",X"FD",
		X"23",X"FD",X"23",X"0C",X"10",X"E2",X"C3",X"94",X"21",X"DD",X"7E",X"02",X"DD",X"21",X"80",X"6A",
		X"DD",X"72",X"06",X"DD",X"73",X"07",X"DD",X"77",X"08",X"DD",X"71",X"00",X"DD",X"56",X"06",X"DD",
		X"5E",X"07",X"DD",X"7E",X"08",X"08",X"FD",X"66",X"00",X"FD",X"6E",X"01",X"FD",X"7E",X"02",X"DD");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
