library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity GFX1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of GFX1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"88",X"CC",X"22",X"22",X"66",X"CC",X"88",X"00",X"33",X"77",X"CC",X"88",X"88",X"77",X"33",X"00",
		X"22",X"22",X"EE",X"EE",X"22",X"22",X"00",X"00",X"00",X"00",X"FF",X"FF",X"44",X"00",X"00",X"00",
		X"22",X"22",X"AA",X"AA",X"EE",X"EE",X"66",X"00",X"66",X"FF",X"BB",X"99",X"99",X"CC",X"44",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"88",X"DD",X"FF",X"BB",X"99",X"88",X"00",X"00",
		X"88",X"EE",X"EE",X"88",X"88",X"88",X"88",X"00",X"00",X"FF",X"FF",X"CC",X"66",X"33",X"11",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"11",X"BB",X"AA",X"AA",X"AA",X"EE",X"EE",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",X"00",X"99",X"99",X"99",X"DD",X"77",X"33",X"00",
		X"00",X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"CC",X"EE",X"BB",X"99",X"88",X"CC",X"CC",X"00",
		X"CC",X"EE",X"AA",X"AA",X"22",X"22",X"CC",X"00",X"00",X"66",X"99",X"99",X"BB",X"FF",X"66",X"00",
		X"88",X"CC",X"66",X"22",X"22",X"22",X"00",X"00",X"77",X"FF",X"99",X"99",X"99",X"FF",X"66",X"00",
		X"31",X"73",X"F7",X"FF",X"FE",X"FE",X"FE",X"FE",X"8E",X"8E",X"8E",X"9E",X"BD",X"BD",X"BD",X"BD",
		X"80",X"E8",X"FE",X"FF",X"FA",X"FB",X"FA",X"F3",X"F0",X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",X"FC",
		X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"FE",X"FF",X"FF",X"F1",X"F6",X"73",X"F7",X"F7",X"BD",X"BD",X"BD",X"BD",X"9E",X"8E",X"8E",X"8E",
		X"F8",X"FF",X"FC",X"FD",X"F4",X"FB",X"FC",X"FD",X"F1",X"FF",X"FF",X"F1",X"FE",X"FF",X"BB",X"BB",
		X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"F7",X"F7",X"F7",X"73",X"F7",X"FF",X"FD",X"D0",X"0C",X"0C",X"0C",X"0C",X"0C",X"1C",X"3D",X"1C",
		X"FC",X"75",X"75",X"75",X"FC",X"C8",X"80",X"00",X"FF",X"FF",X"EE",X"BB",X"BB",X"FF",X"FE",X"E0",
		X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"0F",X"0F",X"8F",X"CF",X"CF",X"CF",X"01",X"00",
		X"F8",X"FF",X"FC",X"FD",X"F4",X"FB",X"FC",X"FD",X"F1",X"FF",X"FF",X"F1",X"FE",X"FF",X"FF",X"DD",
		X"FC",X"76",X"76",X"76",X"FC",X"C8",X"80",X"00",X"FF",X"FF",X"EE",X"FF",X"DD",X"FF",X"FE",X"E0",
		X"0D",X"0D",X"0D",X"0D",X"0D",X"0D",X"0D",X"0D",X"0F",X"07",X"03",X"03",X"03",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"10",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"00",X"00",X"00",X"10",X"70",X"B7",X"BF",X"BF",X"00",X"00",X"00",X"00",X"30",X"F0",X"93",X"13",
		X"C3",X"C3",X"03",X"0B",X"0F",X"8F",X"8F",X"0F",X"00",X"50",X"F0",X"8F",X"FF",X"FF",X"FF",X"FF",
		X"70",X"40",X"E0",X"60",X"C0",X"80",X"00",X"80",X"0C",X"0C",X"0C",X"0C",X"0C",X"1C",X"1C",X"0C",
		X"BF",X"BF",X"CF",X"FF",X"7F",X"3F",X"DF",X"FF",X"03",X"01",X"01",X"01",X"00",X"01",X"13",X"13",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"FF",X"EF",X"1F",X"FF",X"FF",X"FF",X"FF",
		X"70",X"10",X"10",X"00",X"00",X"00",X"0F",X"0F",X"0C",X"0C",X"0C",X"0C",X"0C",X"0E",X"0F",X"0F",
		X"DF",X"1F",X"1F",X"CF",X"EF",X"EF",X"0F",X"0F",X"13",X"01",X"C0",X"41",X"21",X"01",X"0F",X"0F",
		X"8F",X"8F",X"8F",X"8F",X"0B",X"07",X"0F",X"0F",X"F3",X"B3",X"FF",X"FF",X"F7",X"07",X"03",X"0F",
		X"00",X"00",X"00",X"10",X"70",X"B7",X"BF",X"BF",X"00",X"00",X"00",X"00",X"30",X"F0",X"93",X"13",
		X"C3",X"C3",X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"00",X"50",X"0F",X"FF",X"FF",X"FF",X"FF",X"EF",
		X"FF",X"7F",X"3F",X"DF",X"FF",X"DF",X"1F",X"1F",X"01",X"00",X"01",X"13",X"13",X"13",X"01",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"8F",X"8F",X"8F",X"1F",X"FF",X"FF",X"FF",X"FF",X"73",X"33",X"FF",
		X"CF",X"EF",X"EF",X"1F",X"00",X"80",X"69",X"3C",X"01",X"01",X"C1",X"40",X"20",X"10",X"0F",X"0F",
		X"8F",X"0B",X"03",X"03",X"4B",X"87",X"0F",X"0F",X"FF",X"7F",X"07",X"03",X"00",X"00",X"B4",X"4B",
		X"0F",X"0F",X"00",X"10",X"30",X"30",X"30",X"10",X"07",X"0F",X"0E",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"0F",X"0F",X"00",X"00",X"C0",X"C0",X"E0",X"E0",X"0F",X"0F",X"00",X"00",X"E0",X"F0",X"F0",X"F0",
		X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"08",X"0F",X"0F",X"00",X"00",X"22",X"EE",X"BB",X"FF",
		X"0F",X"0F",X"00",X"00",X"00",X"00",X"80",X"80",X"0F",X"0F",X"00",X"E0",X"F0",X"F0",X"70",X"F0",
		X"10",X"10",X"10",X"00",X"00",X"40",X"E0",X"F0",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"1C",
		X"E0",X"E0",X"C0",X"81",X"83",X"07",X"07",X"06",X"F0",X"F0",X"F0",X"70",X"70",X"70",X"20",X"80",
		X"C0",X"E0",X"F0",X"F0",X"F0",X"C0",X"80",X"00",X"F0",X"30",X"1C",X"0E",X"1C",X"38",X"70",X"70",
		X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"60",X"64",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"70",X"20",X"00",X"1C",X"1C",X"1C",X"1C",X"0C",X"0C",X"0C",X"0C",
		X"06",X"04",X"FF",X"FF",X"20",X"70",X"F0",X"F0",X"C0",X"F1",X"F1",X"E0",X"E0",X"C0",X"90",X"30",
		X"00",X"80",X"B3",X"F3",X"F1",X"E0",X"F0",X"70",X"70",X"60",X"10",X"FE",X"FE",X"76",X"D4",X"C4",
		X"00",X"00",X"88",X"EE",X"77",X"33",X"CC",X"FF",X"66",X"FF",X"BB",X"CC",X"CC",X"77",X"33",X"CC",
		X"03",X"03",X"47",X"CF",X"CF",X"8B",X"03",X"47",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"CC",
		X"F0",X"F0",X"F0",X"A0",X"00",X"00",X"0F",X"0F",X"30",X"70",X"70",X"70",X"30",X"00",X"0F",X"0F",
		X"F0",X"F1",X"F1",X"F0",X"F0",X"E0",X"C3",X"0F",X"80",X"90",X"30",X"30",X"30",X"10",X"0F",X"0F",
		X"33",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"CC",X"88",X"00",X"60",X"E0",X"60",X"0F",X"0F",
		X"CF",X"CF",X"CF",X"47",X"03",X"07",X"0F",X"0F",X"FF",X"33",X"00",X"00",X"00",X"00",X"0F",X"0F",
		X"E0",X"E0",X"C0",X"E6",X"A2",X"11",X"11",X"00",X"F0",X"F0",X"F0",X"70",X"70",X"70",X"20",X"80",
		X"C0",X"E0",X"F0",X"70",X"60",X"C0",X"80",X"00",X"F0",X"14",X"0E",X"0F",X"0F",X"0E",X"1C",X"38",
		X"CC",X"EE",X"AA",X"AA",X"22",X"22",X"CC",X"00",X"00",X"66",X"99",X"99",X"BB",X"FF",X"66",X"00",
		X"88",X"CC",X"66",X"22",X"22",X"22",X"00",X"00",X"77",X"FF",X"99",X"99",X"99",X"FF",X"66",X"00",
		X"00",X"00",X"00",X"00",X"88",X"44",X"22",X"00",X"88",X"44",X"22",X"11",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"0F",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"0F",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",
		X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"0F",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"0F",
		X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"88",X"88",X"88",X"EE",X"EE",X"00",X"33",X"77",X"CC",X"88",X"CC",X"77",X"33",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"EE",X"00",X"66",X"FF",X"99",X"99",X"99",X"FF",X"FF",X"00",
		X"44",X"66",X"22",X"22",X"66",X"CC",X"88",X"00",X"44",X"CC",X"88",X"88",X"CC",X"77",X"33",X"00",
		X"88",X"CC",X"66",X"22",X"22",X"EE",X"EE",X"00",X"33",X"77",X"CC",X"88",X"88",X"FF",X"FF",X"00",
		X"22",X"22",X"22",X"22",X"EE",X"EE",X"00",X"00",X"88",X"99",X"99",X"99",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"00",X"88",X"99",X"99",X"99",X"99",X"FF",X"FF",X"00",
		X"EE",X"EE",X"22",X"22",X"66",X"CC",X"88",X"00",X"99",X"99",X"99",X"88",X"CC",X"77",X"33",X"00",
		X"EE",X"EE",X"00",X"00",X"00",X"EE",X"EE",X"00",X"FF",X"FF",X"11",X"11",X"11",X"FF",X"FF",X"00",
		X"22",X"22",X"EE",X"EE",X"22",X"22",X"00",X"00",X"88",X"88",X"FF",X"FF",X"88",X"88",X"00",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"66",X"EE",X"CC",X"88",X"EE",X"EE",X"00",X"88",X"CC",X"66",X"33",X"11",X"FF",X"FF",X"00",
		X"22",X"22",X"22",X"22",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"EE",X"EE",X"00",X"88",X"00",X"EE",X"EE",X"00",X"FF",X"FF",X"77",X"33",X"77",X"FF",X"FF",X"00",
		X"EE",X"EE",X"CC",X"88",X"00",X"EE",X"EE",X"00",X"FF",X"FF",X"11",X"33",X"77",X"FF",X"FF",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",X"77",X"FF",X"88",X"88",X"88",X"FF",X"77",X"00",
		X"00",X"88",X"88",X"88",X"88",X"EE",X"EE",X"00",X"77",X"FF",X"88",X"88",X"88",X"FF",X"FF",X"00",
		X"AA",X"CC",X"EE",X"AA",X"22",X"EE",X"CC",X"00",X"77",X"FF",X"88",X"88",X"88",X"FF",X"77",X"00",
		X"22",X"66",X"EE",X"CC",X"88",X"EE",X"EE",X"00",X"77",X"FF",X"99",X"88",X"88",X"FF",X"FF",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"00",X"55",X"DD",X"99",X"99",X"FF",X"66",X"00",
		X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"00",X"88",X"88",X"FF",X"FF",X"88",X"88",X"00",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"88",X"CC",X"EE",X"CC",X"88",X"00",X"00",X"FF",X"FF",X"11",X"00",X"11",X"FF",X"FF",X"00",
		X"EE",X"EE",X"CC",X"88",X"CC",X"EE",X"EE",X"00",X"FF",X"FF",X"11",X"33",X"11",X"FF",X"FF",X"00",
		X"66",X"EE",X"CC",X"88",X"CC",X"EE",X"66",X"00",X"CC",X"EE",X"77",X"33",X"77",X"EE",X"CC",X"00",
		X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"00",X"EE",X"FF",X"11",X"11",X"FF",X"EE",X"00",X"00",
		X"22",X"22",X"22",X"AA",X"EE",X"EE",X"66",X"00",X"CC",X"EE",X"FF",X"BB",X"99",X"88",X"88",X"00",
		X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0B",X"0B",X"07",X"0F",X"0F",X"0F",X"00",X"00",X"01",X"00",X"00",X"01",X"0F",X"0F",
		X"00",X"00",X"C0",X"C0",X"30",X"F8",X"F4",X"F3",X"00",X"00",X"3C",X"3C",X"2C",X"E0",X"D0",X"D0",
		X"00",X"00",X"00",X"00",X"00",X"88",X"C0",X"E0",X"00",X"00",X"00",X"00",X"E0",X"F0",X"F1",X"FE",
		X"F0",X"30",X"00",X"00",X"00",X"0F",X"0F",X"1F",X"10",X"30",X"20",X"20",X"20",X"20",X"21",X"21",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F1",X"0F",X"0F",X"0F",X"03",X"00",X"C0",X"E0",X"FF",
		X"F7",X"F6",X"F3",X"B7",X"79",X"F0",X"70",X"10",X"F0",X"F0",X"F0",X"D0",X"D0",X"C0",X"E0",X"F0",
		X"E0",X"F0",X"F8",X"F8",X"E0",X"E8",X"C4",X"00",X"FF",X"F3",X"F1",X"FF",X"FF",X"F0",X"F0",X"F0",
		X"FF",X"BB",X"BF",X"33",X"33",X"00",X"80",X"C0",X"21",X"21",X"21",X"20",X"20",X"30",X"10",X"00",
		X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"FF",X"EE",X"CC",X"00",X"00",X"03",X"0E",
		X"C0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"06",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"F0",X"F0",X"F0",X"F0",X"3C",X"0F",X"0F",X"0F",X"02",X"01",X"09",X"0F",X"07",X"03",X"03",X"03",
		X"F0",X"78",X"B4",X"F3",X"FE",X"F6",X"F3",X"B3",X"F0",X"F0",X"F0",X"F0",X"D2",X"D2",X"1E",X"1E",
		X"00",X"88",X"C0",X"E0",X"E0",X"F0",X"F8",X"F8",X"E0",X"F0",X"F1",X"FE",X"FF",X"F3",X"F1",X"FF",
		X"0F",X"0F",X"0F",X"07",X"07",X"00",X"F0",X"F0",X"03",X"01",X"06",X"0F",X"0F",X"0F",X"F0",X"F0",
		X"F9",X"F0",X"70",X"10",X"C0",X"F0",X"F0",X"F0",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"F0",X"F0",
		X"E0",X"E8",X"C4",X"00",X"00",X"00",X"F0",X"F0",X"FF",X"F0",X"F0",X"F0",X"00",X"00",X"F0",X"F0",
		X"00",X"00",X"C0",X"C0",X"31",X"F0",X"F0",X"F3",X"00",X"00",X"3C",X"3C",X"2C",X"E0",X"D0",X"D0",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"00",X"00",X"00",X"00",X"E0",X"F8",X"F0",X"FE",
		X"FF",X"F7",X"F3",X"F3",X"F1",X"F0",X"70",X"60",X"F0",X"F1",X"F0",X"D0",X"D0",X"C0",X"E0",X"F0",
		X"E0",X"F0",X"FA",X"FC",X"E0",X"E0",X"C0",X"00",X"FB",X"FB",X"F3",X"F7",X"FF",X"F8",X"F4",X"F2",
		X"F0",X"F0",X"F0",X"F3",X"FF",X"F7",X"F3",X"F3",X"F0",X"F0",X"F0",X"F0",X"D2",X"D3",X"1E",X"1E",
		X"00",X"80",X"C0",X"E0",X"E0",X"F0",X"F2",X"FC",X"E0",X"F8",X"F4",X"FE",X"FB",X"FB",X"F7",X"F7",
		X"F1",X"F0",X"70",X"10",X"C0",X"F0",X"F0",X"F0",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"F0",X"F0",
		X"E0",X"E0",X"C0",X"00",X"00",X"00",X"F0",X"F0",X"FF",X"F8",X"F4",X"F2",X"00",X"00",X"F0",X"F0",
		X"C0",X"00",X"40",X"20",X"10",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"D2",X"D2",X"1E",X"1E",X"1E",
		X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"20",X"00",X"00",
		X"10",X"20",X"40",X"00",X"C0",X"F0",X"F0",X"F0",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"F0",X"F0",
		X"00",X"00",X"80",X"00",X"00",X"00",X"F0",X"F0",X"20",X"10",X"00",X"00",X"00",X"00",X"F0",X"F0",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"30",X"40",X"F0",X"F0",X"F0",X"D2",X"D2",X"1E",X"1E",X"1E",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"40",X"30",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"F0",X"F0",X"F0",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"80",X"80",X"40",X"00",X"00",X"00",X"F0",X"F0",
		X"F0",X"30",X"00",X"00",X"0F",X"0F",X"3F",X"FF",X"10",X"30",X"20",X"20",X"21",X"21",X"21",X"31",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"E0",X"0F",X"0F",X"0F",X"03",X"10",X"C0",X"EE",X"FF",
		X"11",X"11",X"3B",X"33",X"33",X"00",X"80",X"C0",X"21",X"21",X"20",X"20",X"20",X"30",X"10",X"00",
		X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"55",X"11",X"33",X"00",X"00",X"00",X"03",X"0E",
		X"13",X"11",X"33",X"33",X"33",X"00",X"80",X"C0",X"21",X"21",X"20",X"20",X"20",X"30",X"10",X"00",
		X"0F",X"0F",X"00",X"00",X"00",X"30",X"F1",X"F7",X"0F",X"0F",X"0E",X"0C",X"0C",X"0C",X"0C",X"1C",
		X"87",X"87",X"00",X"F0",X"F0",X"00",X"00",X"00",X"3C",X"78",X"70",X"30",X"10",X"C0",X"EC",X"FE",
		X"0F",X"0F",X"00",X"F0",X"F0",X"70",X"F0",X"FE",X"0F",X"0F",X"00",X"F0",X"F0",X"00",X"30",X"73",
		X"0F",X"0F",X"00",X"00",X"00",X"00",X"E0",X"EC",X"0F",X"0F",X"00",X"C0",X"E0",X"F0",X"F6",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3C",X"79",X"3C",X"1C",X"1C",X"1C",X"1C",X"1C",
		X"80",X"B0",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FF",X"FF",X"FF",X"F7",X"F7",X"FE",X"F8",X"FE",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FF",X"F8",X"FF",X"F3",X"F3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EC",X"EC",X"EC",X"E4",X"E4",X"E4",X"E4",X"E0",X"FF",X"FF",X"FF",X"FF",X"F7",X"F0",X"F0",X"FF",
		X"FF",X"F7",X"FF",X"FF",X"FF",X"F7",X"73",X"30",X"1C",X"0C",X"1C",X"79",X"78",X"0C",X"0C",X"0C",
		X"FB",X"FB",X"F8",X"80",X"80",X"00",X"00",X"00",X"FF",X"F7",X"F7",X"FF",X"FE",X"FC",X"E0",X"80",
		X"FF",X"FF",X"FF",X"F0",X"00",X"00",X"00",X"00",X"FF",X"FF",X"F3",X"F0",X"00",X"00",X"00",X"00",
		X"E4",X"E4",X"E4",X"E4",X"E0",X"00",X"00",X"00",X"FF",X"FF",X"F0",X"80",X"00",X"00",X"00",X"00",
		X"0F",X"78",X"F0",X"80",X"80",X"C0",X"00",X"00",X"0F",X"0F",X"10",X"30",X"30",X"D0",X"EC",X"FE",
		X"0F",X"0F",X"00",X"F0",X"70",X"70",X"F0",X"FE",X"0F",X"C3",X"E0",X"30",X"00",X"00",X"30",X"73",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"00",X"70",X"F2",X"FF",X"F7",X"72",X"0F",X"0F",X"0E",X"0C",X"1C",X"3D",X"1C",X"0C",
		X"0F",X"0F",X"00",X"E0",X"FE",X"FE",X"F1",X"1E",X"0F",X"0F",X"00",X"70",X"F1",X"FD",X"FE",X"F2",
		X"0F",X"87",X"90",X"90",X"90",X"90",X"F0",X"FF",X"0F",X"F0",X"F7",X"F3",X"73",X"73",X"F3",X"FF",
		X"0F",X"0F",X"C0",X"C8",X"C8",X"C0",X"80",X"80",X"0F",X"0F",X"F0",X"FF",X"FF",X"F3",X"F3",X"FB",
		X"F6",X"F6",X"F6",X"F7",X"F7",X"F6",X"F6",X"F6",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"D2",X"96",X"D2",X"96",X"D2",X"96",X"D2",X"1E",X"7A",X"73",X"F3",X"FF",X"FF",X"F3",X"72",X"7A",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"80",X"80",X"00",X"00",X"00",X"E0",X"E8",X"EC",X"FF",X"FE",X"FE",X"FE",X"FE",X"FC",X"FD",X"FF",
		X"72",X"F7",X"FF",X"F4",X"E0",X"00",X"00",X"00",X"0C",X"0C",X"3C",X"3C",X"0C",X"0C",X"0C",X"0C",
		X"F0",X"FF",X"FE",X"E0",X"80",X"00",X"00",X"00",X"F2",X"FF",X"FD",X"FD",X"F0",X"00",X"00",X"00",
		X"FC",X"F0",X"10",X"90",X"80",X"80",X"80",X"00",X"FF",X"F2",X"72",X"72",X"73",X"73",X"70",X"00",
		X"EC",X"EC",X"EC",X"E4",X"E4",X"E4",X"E0",X"00",X"F7",X"F6",X"FE",X"F0",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"80",X"80",X"90",X"90",X"F0",X"FF",X"0F",X"0F",X"00",X"F0",X"F3",X"73",X"F3",X"FF",
		X"0F",X"E1",X"E4",X"E4",X"E4",X"EC",X"EC",X"EC",X"0F",X"0F",X"00",X"00",X"F0",X"FE",X"FE",X"FF",
		X"D0",X"90",X"D0",X"90",X"D0",X"90",X"D0",X"10",X"72",X"72",X"F3",X"FF",X"FF",X"F3",X"72",X"72",
		X"EC",X"E8",X"E0",X"00",X"00",X"80",X"80",X"80",X"FF",X"FD",X"FC",X"FE",X"FE",X"FE",X"FF",X"FB",
		X"FF",X"F0",X"90",X"90",X"90",X"10",X"10",X"10",X"FF",X"F3",X"73",X"73",X"70",X"00",X"00",X"00",
		X"80",X"80",X"C0",X"C8",X"C8",X"C8",X"C0",X"00",X"FB",X"F3",X"F3",X"F3",X"FF",X"FF",X"F0",X"00",
		X"FF",X"FF",X"FF",X"F7",X"FB",X"F3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",
		X"FF",X"DD",X"DD",X"55",X"77",X"77",X"FF",X"FF",X"FF",X"DD",X"DD",X"DD",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"33",X"FF",X"FF",X"FF",X"FF",X"FF",X"88",X"FF",X"EE",X"FF",X"88",X"FF",X"FF",
		X"FF",X"F7",X"7B",X"3D",X"7B",X"7B",X"F7",X"FF",X"FF",X"FF",X"FC",X"CB",X"CB",X"ED",X"FE",X"FF",
		X"FF",X"FF",X"FF",X"FB",X"F7",X"7B",X"F3",X"FF",X"FF",X"FF",X"FF",X"FD",X"FB",X"FE",X"EE",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F4",X"F6",X"F4",X"FF",X"FF",X"FF",X"FF",X"FF",X"F2",X"FB",X"F2",
		X"F4",X"FD",X"F4",X"FF",X"FF",X"FF",X"FF",X"FF",X"F2",X"F6",X"F2",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F5",X"F1",X"FF",X"F5",X"F1",X"FF",X"F5",X"F1",
		X"F8",X"FA",X"FF",X"F8",X"FA",X"FF",X"F8",X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"F1",X"F6",X"F8",X"F8",X"FC",X"FC",X"FF",
		X"FF",X"F8",X"F6",X"F1",X"F1",X"F3",X"F3",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"F1",X"F1",X"F7",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"FA",X"FA",X"F9",
		X"FF",X"F7",X"F1",X"F1",X"FF",X"FF",X"FF",X"FF",X"F9",X"FA",X"FA",X"FC",X"FE",X"FF",X"FF",X"FF",
		X"FF",X"F3",X"F3",X"F1",X"F1",X"F6",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",X"FF",X"FC",X"FC",X"F8",X"F8",X"F6",X"F1",X"FF",
		X"F9",X"F5",X"F5",X"F3",X"F7",X"FF",X"FF",X"FF",X"FF",X"FE",X"F8",X"F8",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"F7",X"F3",X"F5",X"F5",X"F9",X"FF",X"FF",X"FF",X"FF",X"F8",X"F8",X"FE",X"FF",
		X"FF",X"FF",X"FF",X"77",X"33",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CC",X"DD",X"EE",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"33",X"BB",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"CC",X"FF",X"FF",X"FF",
		X"F8",X"FA",X"FF",X"F8",X"FA",X"F4",X"F0",X"F2",X"FF",X"FF",X"FF",X"FF",X"FF",X"F2",X"FB",X"F2",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F4",X"F6",X"F4",X"F5",X"F1",X"FF",X"F5",X"F1",X"F2",X"F9",X"F0",
		X"F0",X"F9",X"F4",X"F8",X"FA",X"FF",X"F8",X"FA",X"F2",X"F6",X"F2",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F4",X"FD",X"F4",X"FF",X"FF",X"FF",X"FF",X"FF",X"F4",X"F0",X"F2",X"F5",X"F1",X"FF",X"F5",X"F1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"CC",X"88",X"88",X"00",X"00",X"00",X"00",
		X"FF",X"33",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"CC",X"FF",
		X"00",X"00",X"00",X"00",X"11",X"11",X"33",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"C8",X"EC",X"FE",X"00",X"00",X"C0",X"FC",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"EC",X"8C",X"80",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FC",X"C0",X"00",X"00",
		X"00",X"70",X"F7",X"FF",X"FF",X"3F",X"37",X"FF",X"00",X"00",X"00",X"10",X"10",X"21",X"21",X"37",
		X"FF",X"37",X"3F",X"FF",X"FF",X"F7",X"70",X"00",X"73",X"21",X"21",X"10",X"10",X"00",X"00",X"00",
		X"00",X"08",X"0C",X"04",X"04",X"02",X"02",X"02",X"00",X"00",X"01",X"01",X"01",X"02",X"02",X"02",
		X"02",X"02",X"02",X"04",X"04",X"0C",X"08",X"00",X"02",X"02",X"02",X"01",X"01",X"01",X"00",X"00",
		X"FE",X"E8",X"EC",X"FE",X"FA",X"E4",X"C4",X"C4",X"FF",X"FF",X"FF",X"FF",X"F6",X"73",X"30",X"31",
		X"00",X"00",X"00",X"80",X"C8",X"EC",X"EC",X"FE",X"80",X"E8",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"7F",X"F3",X"30",X"00",X"00",X"00",X"00",X"43",X"21",X"10",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"1F",X"3F",X"1F",X"0F",X"3F",X"1F",X"7F",X"10",X"21",X"43",X"87",X"87",X"87",X"87",X"87",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"CF",X"EF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"EF",X"EF",X"CF",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"79",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"2F",X"0F",X"0F",X"0F",X"0F",X"4F",X"0F",X"0F",X"8F",X"0F",X"0F",X"1F",X"8F",X"0F",X"0F",X"2F",
		X"BF",X"1F",X"6F",X"0F",X"6F",X"1F",X"1F",X"BF",X"CF",X"BF",X"9F",X"0F",X"6F",X"2F",X"0F",X"CF",
		X"FF",X"FF",X"BF",X"FF",X"3F",X"DF",X"7F",X"FF",X"FF",X"AF",X"BF",X"EF",X"EF",X"BF",X"9F",X"FF",
		X"FF",X"FF",X"FF",X"7F",X"FF",X"BF",X"FF",X"FF",X"FF",X"BF",X"EF",X"EF",X"FF",X"DF",X"FF",X"FF",
		X"F2",X"F1",X"F2",X"F1",X"F2",X"F1",X"F2",X"F1",X"F8",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",
		X"F2",X"F1",X"F2",X"F1",X"F2",X"F1",X"F2",X"F1",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",
		X"F1",X"F1",X"F1",X"F1",X"F0",X"F0",X"F0",X"F0",X"F4",X"F8",X"F4",X"F8",X"F4",X"F8",X"F4",X"F8",
		X"F0",X"F0",X"F0",X"F0",X"F1",X"F1",X"F1",X"F1",X"F4",X"F8",X"F4",X"F8",X"F4",X"F8",X"F4",X"F8",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FA",X"F5",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"FA",X"F5",
		X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"FA",X"F5",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FA",X"F5",
		X"F5",X"FA",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F5",X"FA",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",
		X"F5",X"FA",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"F5",X"FA",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"30",X"30",X"30",X"30",X"30",X"F0",X"F0",X"FF",X"C0",X"C0",X"C0",X"C0",X"C0",X"F0",X"F0",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"F0",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"F0",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"FF",X"C0",X"C0",X"C0",X"C0",X"C0",X"F0",X"F0",X"FF",
		X"30",X"30",X"30",X"30",X"30",X"F0",X"F0",X"FF",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"FF",
		X"FF",X"F0",X"F0",X"30",X"30",X"30",X"30",X"30",X"FF",X"F0",X"F0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"0F",X"F0",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"F0",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"FF",X"F0",X"F0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"FF",X"F0",X"F0",X"30",X"30",X"30",X"30",X"30",X"FF",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"71",X"71",X"71",X"71",X"71",X"71",X"F1",X"F1",X"C0",X"C0",X"C0",X"C0",X"C0",X"E0",X"F0",X"F8",
		X"E9",X"E9",X"E9",X"E9",X"E9",X"E9",X"E9",X"E9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F1",X"F1",X"71",X"71",X"71",X"71",X"71",X"71",X"F8",X"F0",X"E0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"71",X"71",X"71",X"71",X"71",X"71",X"F1",X"F1",X"C0",X"C0",X"C0",X"C0",X"C0",X"E0",X"F0",X"F8",
		X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"F8",X"E8",X"E8",X"E8",X"E8",X"E8",X"E8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"68",X"68",X"68",X"68",X"68",X"68",X"68",X"68",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"68",X"68",X"68",X"68",X"68",X"68",X"78",X"78",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"F0",X"E0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"F1",X"F0",X"70",X"30",X"30",X"30",X"30",X"30",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"C0",X"C0",X"C0",X"C0",X"C0",X"E0",X"F0",X"F8",
		X"30",X"30",X"30",X"30",X"30",X"70",X"F0",X"F1",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",
		X"F1",X"F0",X"70",X"30",X"30",X"30",X"30",X"30",X"F8",X"F0",X"E0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"30",X"30",X"30",X"30",X"30",X"70",X"F0",X"F1",X"C0",X"C0",X"C0",X"C0",X"C0",X"E0",X"F0",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",
		X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"F3",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"EE",X"66",X"33",X"DD",X"55",X"DD",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"33",X"33",X"66",X"55",X"55",X"55",X"66",X"FF",X"88",X"00",X"55",X"88",X"00",X"88",X"FF",
		X"66",X"EE",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"88",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"77",X"44",X"44",X"77",X"00",X"00",X"00",X"00",X"FF",X"11",X"11",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"44",X"44",X"77",X"00",X"00",X"00",X"00",X"FF",X"99",X"99",X"99",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"77",X"44",X"44",X"77",X"00",X"77",X"44",X"00",X"FF",X"11",X"11",X"FF",X"00",X"FF",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"77",X"00",X"77",X"44",X"00",X"00",X"00",X"11",X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"77",X"44",X"44",X"77",X"00",X"77",X"44",X"00",X"FF",X"11",X"11",X"FF",X"00",X"FF",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"77",X"00",X"77",X"44",X"44",X"00",X"00",X"11",X"FF",X"00",X"99",X"99",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"77",X"44",X"44",X"77",X"00",X"77",X"44",X"00",X"FF",X"11",X"11",X"FF",X"00",X"FF",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"77",X"00",X"77",X"00",X"00",X"77",X"00",X"11",X"FF",X"00",X"FF",X"88",X"88",X"88",X"00",
		X"F0",X"F0",X"F0",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FE",X"F9",X"F7",X"F7",X"F3",X"F3",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F1",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F7",X"F9",X"FE",X"FE",X"FC",X"FC",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F1",X"F3",X"F5",X"F5",X"F6",
		X"F0",X"F0",X"F0",X"F0",X"FE",X"FE",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F8",X"FE",X"FE",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F6",X"F5",X"F5",X"F3",X"F1",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"77",X"44",X"44",X"77",X"00",X"77",X"44",X"00",X"FF",X"11",X"11",X"FF",X"00",X"FF",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"77",X"00",X"77",X"44",X"44",X"77",X"00",X"11",X"FF",X"00",X"FF",X"99",X"99",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"44",X"44",X"77",X"00",X"77",X"44",X"44",X"FF",X"11",X"11",X"FF",X"00",X"FF",X"11",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"00",X"44",X"44",X"44",X"77",X"00",X"77",X"FF",X"00",X"FF",X"99",X"99",X"FF",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"44",X"77",X"00",X"77",X"44",X"77",X"00",X"FF",X"11",X"FF",X"00",X"FF",X"11",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"44",X"44",X"00",X"77",X"44",X"44",X"00",X"99",X"99",X"FF",X"00",X"FF",X"99",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"44",X"77",X"00",X"77",X"44",X"77",X"00",X"FF",X"11",X"FF",X"00",X"FF",X"11",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"00",X"77",X"00",X"44",X"44",X"77",X"00",X"FF",X"44",X"44",X"00",X"FF",X"99",X"FF",X"00",
		X"80",X"80",X"80",X"C0",X"C0",X"80",X"00",X"00",X"10",X"10",X"10",X"30",X"30",X"10",X"00",X"00",
		X"70",X"43",X"0F",X"2F",X"4F",X"97",X"C3",X"70",X"E0",X"3C",X"0F",X"4F",X"2F",X"9E",X"3C",X"E0",
		X"00",X"80",X"80",X"00",X"80",X"80",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"30",X"30",
		X"A1",X"E1",X"43",X"43",X"C3",X"C3",X"F0",X"C0",X"48",X"78",X"3C",X"2C",X"3C",X"3C",X"E0",X"00",
		X"00",X"00",X"00",X"C0",X"C0",X"E0",X"4C",X"4C",X"00",X"00",X"10",X"F0",X"43",X"C3",X"97",X"87",
		X"00",X"00",X"80",X"C0",X"68",X"BC",X"1E",X"5E",X"00",X"00",X"00",X"60",X"60",X"70",X"C3",X"0F",
		X"2C",X"2C",X"F0",X"F0",X"30",X"30",X"00",X"00",X"87",X"97",X"C3",X"43",X"F0",X"10",X"00",X"00",
		X"5E",X"1E",X"BC",X"68",X"C0",X"80",X"00",X"00",X"0F",X"C3",X"70",X"C0",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"01",X"01",X"11",
		X"00",X"10",X"11",X"11",X"11",X"11",X"11",X"11",X"00",X"00",X"00",X"10",X"11",X"11",X"11",X"11",
		X"00",X"10",X"10",X"10",X"10",X"00",X"00",X"00",X"11",X"01",X"01",X"10",X"10",X"00",X"00",X"00",
		X"11",X"11",X"11",X"11",X"11",X"11",X"10",X"00",X"11",X"11",X"11",X"11",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"80",X"88",X"88",X"00",X"00",X"00",X"10",X"10",X"01",X"01",X"11",
		X"00",X"10",X"91",X"91",X"91",X"19",X"19",X"99",X"00",X"80",X"80",X"98",X"99",X"99",X"99",X"99",
		X"88",X"98",X"98",X"90",X"10",X"00",X"00",X"00",X"11",X"01",X"01",X"10",X"10",X"00",X"00",X"00",
		X"99",X"19",X"19",X"99",X"99",X"91",X"10",X"00",X"99",X"99",X"99",X"99",X"98",X"80",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"44",X"77",X"00",X"77",X"44",X"77",X"00",X"FF",X"11",X"FF",X"00",X"FF",X"11",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"44",X"77",X"00",X"77",X"44",X"77",X"00",X"FF",X"11",X"FF",X"00",X"FF",X"88",X"88",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"77",X"44",X"77",X"00",X"77",X"44",X"77",X"00",X"FF",X"11",X"FF",X"00",X"FF",X"11",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"77",X"44",X"77",X"00",X"00",X"77",X"00",X"00",X"FF",X"11",X"FF",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"01",X"01",X"01",X"00",X"10",X"30",
		X"02",X"2F",X"EF",X"BB",X"FF",X"5B",X"E1",X"F0",X"00",X"00",X"00",X"08",X"8C",X"CE",X"EF",X"7F",
		X"01",X"00",X"00",X"00",X"04",X"04",X"01",X"03",X"70",X"F0",X"F0",X"F0",X"F0",X"E0",X"C0",X"00",
		X"E1",X"E1",X"D3",X"93",X"13",X"13",X"01",X"00",X"7F",X"EF",X"CE",X"CE",X"8D",X"8C",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",
		X"04",X"4E",X"EF",X"BB",X"FF",X"5F",X"34",X"70",X"00",X"00",X"00",X"80",X"8C",X"CE",X"6F",X"B7",
		X"08",X"00",X"00",X"00",X"04",X"04",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"E1",X"D3",X"93",X"01",X"00",X"B7",X"6F",X"4E",X"CF",X"8C",X"8C",X"08",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"99",X"11",X"11",X"FF",X"FF",X"FF",X"FF",X"FF",X"CC",X"CE",X"89",
		X"FF",X"EE",X"CC",X"CC",X"CC",X"44",X"00",X"00",X"FF",X"00",X"00",X"00",X"11",X"77",X"77",X"00",
		X"11",X"11",X"99",X"FF",X"FF",X"FF",X"FF",X"FF",X"89",X"CE",X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"44",X"44",X"CC",X"CC",X"CC",X"EE",X"FF",X"00",X"77",X"77",X"11",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"31",X"31",X"10",X"00",
		X"00",X"00",X"10",X"21",X"EA",X"FB",X"F7",X"F7",X"40",X"E4",X"FE",X"76",X"46",X"EF",X"FE",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"20",
		X"F7",X"F6",X"F4",X"F5",X"F1",X"71",X"30",X"C0",X"F0",X"E4",X"ED",X"EC",X"EF",X"EC",X"E1",X"00",
		X"00",X"20",X"10",X"20",X"90",X"D0",X"E0",X"ED",X"00",X"00",X"00",X"10",X"10",X"00",X"10",X"31",
		X"00",X"00",X"C0",X"EC",X"FC",X"F3",X"FF",X"77",X"00",X"00",X"00",X"00",X"F0",X"FF",X"FC",X"F9",
		X"EC",X"EC",X"E8",X"A0",X"00",X"00",X"00",X"00",X"62",X"F7",X"73",X"30",X"00",X"00",X"00",X"00",
		X"77",X"FF",X"EF",X"34",X"00",X"00",X"00",X"00",X"F3",X"F7",X"F0",X"82",X"00",X"00",X"00",X"00",
		X"F0",X"70",X"B0",X"B0",X"70",X"F0",X"B0",X"70",X"F0",X"E0",X"D0",X"D0",X"E0",X"F0",X"D0",X"E0",
		X"E0",X"72",X"B0",X"B0",X"30",X"B0",X"30",X"B0",X"70",X"E4",X"D0",X"D0",X"C0",X"D0",X"C0",X"D0",
		X"F0",X"F0",X"B0",X"70",X"B0",X"F0",X"F0",X"F0",X"F0",X"F0",X"D0",X"E0",X"D0",X"F0",X"F0",X"F0",
		X"30",X"70",X"70",X"70",X"90",X"E0",X"70",X"00",X"C0",X"E0",X"E0",X"E0",X"90",X"30",X"70",X"70",
		X"F0",X"F0",X"70",X"F0",X"F0",X"70",X"30",X"80",X"F0",X"F0",X"C0",X"B0",X"B0",X"C0",X"F4",X"70",
		X"F0",X"F0",X"D0",X"60",X"50",X"00",X"F0",X"F0",X"F0",X"F0",X"D0",X"E0",X"00",X"70",X"F0",X"F0",
		X"A0",X"60",X"60",X"C0",X"F0",X"70",X"F0",X"F0",X"70",X"F4",X"C0",X"B0",X"B0",X"C0",X"F0",X"F0",
		X"F0",X"F0",X"00",X"50",X"60",X"D0",X"F0",X"F0",X"F0",X"F0",X"70",X"00",X"E0",X"D0",X"F0",X"F0",
		X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"FF",X"7F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"80",X"80",X"C0",X"80",X"40",X"00",X"00",X"00",X"00",X"10",X"10",X"30",X"30",
		X"00",X"10",X"60",X"F0",X"F0",X"F3",X"F7",X"74",X"00",X"C0",X"F0",X"70",X"FC",X"FE",X"FE",X"F6",
		X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"20",X"10",X"30",X"10",X"10",X"00",X"00",X"00",
		X"F6",X"F7",X"F7",X"F3",X"E0",X"F0",X"30",X"00",X"E2",X"FE",X"FC",X"F0",X"F0",X"60",X"80",X"00",
		X"00",X"00",X"00",X"80",X"00",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"10",X"10",X"30",X"30",
		X"00",X"10",X"70",X"F0",X"70",X"B3",X"F7",X"96",X"00",X"C0",X"F0",X"F0",X"FC",X"EE",X"96",X"96",
		X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"30",X"30",X"30",X"10",X"00",X"00",X"00",X"00",
		X"96",X"96",X"F7",X"73",X"F0",X"F0",X"30",X"00",X"96",X"FC",X"DC",X"E0",X"F0",X"E0",X"80",X"00",
		X"F0",X"F0",X"F0",X"70",X"70",X"30",X"30",X"30",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"C0",X"C0",
		X"F0",X"E0",X"80",X"00",X"00",X"30",X"70",X"70",X"F0",X"30",X"00",X"00",X"C0",X"E0",X"A4",X"68",
		X"30",X"30",X"70",X"70",X"F0",X"F0",X"F0",X"F0",X"C0",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F0",
		X"61",X"52",X"70",X"30",X"00",X"00",X"C0",X"F0",X"E0",X"E0",X"C0",X"00",X"00",X"10",X"20",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"B7",X"B7",X"B7",X"B7",X"B7",X"B7",X"B7",X"B7",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"B7",X"B7",X"B7",X"B7",X"B7",X"B7",X"B7",X"B7",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"A0",X"50",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"A0",X"50",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",
		X"A0",X"50",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"A0",X"50",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"D0",X"E0",X"D0",X"E0",X"D0",X"E0",X"D0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"70",X"70",X"70",X"F0",X"F0",X"F0",X"F0",
		X"D0",X"E0",X"D0",X"E0",X"D0",X"E0",X"D0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"70",X"70",X"70",X"70",
		X"00",X"80",X"80",X"80",X"88",X"CC",X"88",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"11",X"10",
		X"00",X"11",X"73",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"98",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F7",X"33",X"77",X"F7",X"F7",X"F3",X"00",X"00",X"FE",X"FC",X"FE",X"EE",X"EE",X"CC",X"80",X"40",
		X"00",X"00",X"00",X"00",X"00",X"88",X"DC",X"EC",X"00",X"00",X"00",X"70",X"71",X"31",X"33",X"77",
		X"00",X"00",X"44",X"EE",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"60",X"FB",X"FF",X"FF",
		X"CC",X"CC",X"C8",X"C0",X"00",X"00",X"00",X"00",X"77",X"33",X"31",X"11",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"44",X"00",X"00",X"FF",X"FF",X"BB",X"90",X"80",X"00",X"00",X"00",
		X"FF",X"77",X"77",X"33",X"33",X"33",X"77",X"99",X"FF",X"EE",X"EE",X"CC",X"CC",X"CC",X"EE",X"FF",
		X"EE",X"88",X"60",X"62",X"00",X"22",X"55",X"00",X"77",X"11",X"66",X"62",X"00",X"AA",X"44",X"00",
		X"11",X"33",X"FF",X"77",X"77",X"11",X"11",X"FF",X"FF",X"FF",X"CC",X"99",X"FF",X"88",X"99",X"FF",
		X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"33",X"00",X"00",X"00",X"00",X"00",X"22",X"77",
		X"FF",X"99",X"99",X"11",X"33",X"77",X"33",X"11",X"FF",X"FF",X"EE",X"88",X"CC",X"B9",X"B8",X"00",
		X"FF",X"EE",X"22",X"11",X"00",X"44",X"22",X"44",X"FF",X"77",X"33",X"22",X"88",X"88",X"00",X"00",
		X"11",X"33",X"33",X"33",X"BB",X"99",X"99",X"FF",X"00",X"B9",X"B8",X"CC",X"88",X"EE",X"FF",X"FF",
		X"22",X"44",X"22",X"00",X"11",X"33",X"FF",X"FF",X"00",X"00",X"88",X"88",X"DD",X"CC",X"EE",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"31",X"71",X"73",X"F3",X"F3",X"70",
		X"80",X"C0",X"E8",X"FC",X"FE",X"FC",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"00",X"00",X"80",X"80",X"00",X"00",X"10",X"30",X"71",X"F3",X"F3",X"71",X"30",
		X"60",X"F0",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"80",X"C0",X"F8",X"FE",X"FE",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F3",X"72",X"70",X"20",X"00",X"00",X"00",X"00",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"E8",X"E8",X"00",X"00",X"40",X"60",X"00",X"10",X"70",X"31",
		X"20",X"E0",X"F3",X"F3",X"F3",X"F7",X"FF",X"FF",X"00",X"80",X"C0",X"E8",X"FC",X"FE",X"FF",X"FF",
		X"C0",X"80",X"80",X"C0",X"C0",X"80",X"00",X"00",X"31",X"71",X"70",X"30",X"10",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"F7",X"FF",X"10",X"00",X"00",X"BF",X"3F",X"FF",X"FB",X"F8",X"C0",X"00",X"00",
		X"00",X"80",X"E0",X"C0",X"00",X"E0",X"FC",X"FE",X"00",X"00",X"00",X"10",X"C0",X"C4",X"80",X"10",
		X"60",X"F0",X"F7",X"FF",X"F7",X"F7",X"F7",X"F7",X"00",X"80",X"D0",X"E8",X"FC",X"FE",X"FF",X"FF",
		X"FE",X"7E",X"7E",X"7C",X"EC",X"E0",X"40",X"00",X"30",X"71",X"F3",X"F7",X"F3",X"71",X"30",X"10",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"E8",X"C0",X"FF",X"FF",X"EF",X"C7",X"F3",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"80",X"C8",X"EC",X"EC",X"EC",X"00",X"00",X"00",X"10",X"31",X"73",X"73",X"73",
		X"00",X"10",X"71",X"97",X"BD",X"9F",X"FF",X"FF",X"00",X"80",X"E8",X"9E",X"DB",X"9F",X"FF",X"FF",
		X"C8",X"C8",X"80",X"80",X"00",X"00",X"00",X"00",X"31",X"31",X"10",X"10",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"F7",X"73",X"F6",X"E0",X"FF",X"FF",X"FF",X"FF",X"FC",X"C8",X"80",X"00",
		X"00",X"00",X"00",X"00",X"80",X"80",X"C8",X"EC",X"00",X"00",X"00",X"10",X"10",X"21",X"21",X"73",
		X"00",X"70",X"F7",X"FF",X"FF",X"3F",X"B7",X"FF",X"00",X"00",X"C0",X"FC",X"FF",X"FF",X"FF",X"FF",
		X"EC",X"FE",X"FA",X"B0",X"10",X"00",X"00",X"00",X"73",X"21",X"21",X"10",X"10",X"00",X"00",X"00",
		X"FF",X"B7",X"3F",X"FF",X"FF",X"F7",X"70",X"00",X"FF",X"FF",X"FF",X"FF",X"FC",X"C0",X"00",X"00",
		X"F0",X"F0",X"F0",X"78",X"3C",X"1E",X"1E",X"1E",X"F0",X"F0",X"F0",X"E1",X"C3",X"87",X"87",X"87",
		X"F0",X"E1",X"87",X"0F",X"0F",X"2D",X"0F",X"0F",X"F0",X"78",X"1E",X"0F",X"0F",X"B4",X"0F",X"0F",
		X"3C",X"3C",X"78",X"78",X"F0",X"F0",X"F0",X"F0",X"C3",X"C3",X"E1",X"E1",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"C3",X"87",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"3C",X"78",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"78",X"78",X"3C",X"1E",X"F0",X"F0",X"F0",X"E1",X"E1",X"C3",X"C3",X"87",
		X"F0",X"87",X"0F",X"0F",X"0F",X"0F",X"4B",X"0F",X"F0",X"F0",X"3C",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"1E",X"1E",X"5A",X"78",X"F0",X"F0",X"F0",X"F0",X"87",X"C3",X"C3",X"E1",X"E1",X"F0",X"F0",X"F0",
		X"0F",X"4B",X"0F",X"0F",X"0F",X"0F",X"87",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"3C",X"F0",X"F0",
		X"80",X"48",X"2C",X"1E",X"1E",X"1E",X"E5",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"21",X"43",X"43",X"63",X"F7",X"F7",X"F0",X"0F",X"0F",X"0F",X"0F",X"8F",X"AF",X"EF",
		X"FE",X"EC",X"EC",X"C8",X"80",X"00",X"00",X"00",X"10",X"31",X"F3",X"72",X"F1",X"10",X"30",X"10",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"F9",X"A0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"E8",X"80",
		X"00",X"00",X"80",X"48",X"48",X"48",X"EC",X"EC",X"00",X"00",X"00",X"10",X"10",X"10",X"00",X"00",
		X"30",X"43",X"87",X"0F",X"0F",X"2F",X"F7",X"F7",X"E0",X"1E",X"0F",X"0F",X"0F",X"9F",X"AF",X"FF",
		X"FE",X"EC",X"EC",X"C8",X"80",X"C8",X"80",X"40",X"10",X"31",X"73",X"72",X"B1",X"10",X"31",X"10",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"F9",X"90",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F5",X"50",
		X"00",X"00",X"00",X"80",X"C8",X"EC",X"EC",X"FE",X"10",X"21",X"43",X"87",X"87",X"87",X"87",X"87",
		X"F0",X"1F",X"3F",X"1F",X"0F",X"3F",X"1F",X"7F",X"80",X"E8",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"F9",X"FD",X"FE",X"FA",X"F5",X"C8",X"C8",X"43",X"21",X"10",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"7F",X"F3",X"30",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"F6",X"73",X"30",X"31",
		X"00",X"00",X"50",X"E4",X"FE",X"EC",X"FE",X"EC",X"00",X"00",X"10",X"21",X"43",X"87",X"87",X"87",
		X"00",X"30",X"F3",X"3F",X"5F",X"3F",X"1F",X"7F",X"80",X"E8",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"E8",X"EC",X"FE",X"FA",X"A0",X"00",X"80",X"87",X"87",X"43",X"21",X"10",X"00",X"00",X"00",
		X"3F",X"7F",X"3F",X"3C",X"C0",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"F6",X"73",X"30",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
