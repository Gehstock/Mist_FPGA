library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity tn03 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of tn03 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"0F",X"21",X"74",X"20",X"7E",X"FE",X"30",X"DC",X"22",X"10",X"FE",X"E8",X"D4",X"2A",X"10",X"2B",
		X"7E",X"FE",X"18",X"DA",X"31",X"10",X"21",X"71",X"20",X"CD",X"A1",X"0D",X"2A",X"73",X"20",X"C3",
		X"2B",X"0F",X"F5",X"E5",X"2A",X"73",X"20",X"C3",X"4B",X"0F",X"E5",X"2A",X"73",X"20",X"C3",X"57",
		X"0F",X"2A",X"73",X"20",X"CD",X"3E",X"0F",X"21",X"6E",X"46",X"11",X"6E",X"20",X"C3",X"67",X"0F",
		X"21",X"11",X"20",X"AF",X"BE",X"C8",X"36",X"00",X"21",X"14",X"20",X"34",X"21",X"00",X"00",X"22",
		X"16",X"20",X"2A",X"1A",X"20",X"CD",X"C3",X"08",X"21",X"60",X"20",X"AF",X"BE",X"CA",X"B0",X"10",
		X"21",X"65",X"20",X"CD",X"8F",X"10",X"D4",X"6C",X"10",X"C3",X"B0",X"10",X"CD",X"96",X"10",X"DA",
		X"73",X"10",X"C9",X"CD",X"9D",X"10",X"D2",X"7A",X"10",X"C9",X"CD",X"A9",X"10",X"DA",X"81",X"10",
		X"C9",X"E1",X"2A",X"65",X"20",X"22",X"93",X"20",X"21",X"91",X"20",X"34",X"C3",X"5E",X"0F",X"3A",
		X"1A",X"20",X"C6",X"08",X"BE",X"C9",X"F5",X"3E",X"10",X"86",X"C3",X"A5",X"10",X"3A",X"1B",X"20",
		X"23",X"F5",X"7E",X"D6",X"08",X"47",X"F1",X"B8",X"C9",X"F5",X"3E",X"10",X"86",X"C3",X"A5",X"10",
		X"21",X"67",X"20",X"AF",X"BE",X"CA",X"E7",X"10",X"21",X"6C",X"20",X"CD",X"8F",X"10",X"D4",X"C4",
		X"10",X"C3",X"E7",X"10",X"CD",X"96",X"10",X"DA",X"CB",X"10",X"C9",X"CD",X"9D",X"10",X"D2",X"D2",
		X"10",X"C9",X"CD",X"A9",X"10",X"DA",X"D9",X"10",X"C9",X"E1",X"2A",X"6C",X"20",X"22",X"93",X"20",
		X"21",X"91",X"20",X"34",X"C3",X"CB",X"0F",X"21",X"6E",X"20",X"AF",X"BE",X"CA",X"1E",X"11",X"21",
		X"73",X"20",X"CD",X"8F",X"10",X"D4",X"FB",X"10",X"C3",X"1E",X"11",X"CD",X"96",X"10",X"DA",X"02",
		X"11",X"C9",X"CD",X"9D",X"10",X"D2",X"09",X"11",X"C9",X"CD",X"A9",X"10",X"DA",X"10",X"11",X"C9",
		X"E1",X"2A",X"73",X"20",X"22",X"93",X"20",X"21",X"91",X"20",X"34",X"C3",X"31",X"10",X"21",X"38",
		X"20",X"22",X"75",X"20",X"0E",X"06",X"7E",X"A7",X"CA",X"33",X"11",X"23",X"23",X"CD",X"8F",X"10",
		X"D4",X"44",X"11",X"2A",X"75",X"20",X"11",X"04",X"00",X"19",X"22",X"75",X"20",X"0D",X"C2",X"26",
		X"11",X"C3",X"71",X"11",X"CD",X"96",X"10",X"DA",X"4B",X"11",X"C9",X"CD",X"9D",X"10",X"D2",X"52",
		X"11",X"C9",X"CD",X"A9",X"10",X"DA",X"59",X"11",X"C9",X"F1",X"2B",X"2B",X"2B",X"36",X"00",X"CD",
		X"6A",X"11",X"22",X"29",X"20",X"21",X"27",X"20",X"34",X"C9",X"23",X"23",X"5E",X"23",X"56",X"EB",
		X"C9",X"CD",X"07",X"13",X"22",X"77",X"20",X"0E",X"06",X"E5",X"21",X"1F",X"20",X"34",X"E1",X"7E",
		X"07",X"DC",X"9D",X"11",X"2A",X"77",X"20",X"11",X"04",X"00",X"19",X"22",X"77",X"20",X"0D",X"C2",
		X"79",X"11",X"21",X"1F",X"20",X"36",X"00",X"CD",X"E2",X"14",X"C3",X"7D",X"15",X"CD",X"6A",X"11",
		X"7C",X"FE",X"3C",X"D0",X"C5",X"CD",X"49",X"0D",X"22",X"79",X"20",X"C1",X"21",X"79",X"20",X"3A",
		X"1A",X"20",X"C6",X"0A",X"BE",X"D2",X"B9",X"11",X"C9",X"F5",X"3E",X"20",X"86",X"47",X"F1",X"B8",
		X"DA",X"C4",X"11",X"C9",X"3A",X"1B",X"20",X"23",X"F5",X"7E",X"D6",X"08",X"47",X"F1",X"B8",X"D2",
		X"D3",X"11",X"C9",X"F5",X"3E",X"23",X"86",X"47",X"F1",X"B8",X"DA",X"DE",X"11",X"C9",X"F1",X"E5",
		X"21",X"1D",X"20",X"34",X"2A",X"1A",X"20",X"01",X"00",X"F6",X"09",X"22",X"22",X"20",X"2A",X"77",
		X"20",X"7E",X"E6",X"0F",X"77",X"CD",X"6A",X"11",X"CD",X"89",X"08",X"E1",X"2B",X"3E",X"05",X"86",
		X"47",X"3A",X"1A",X"20",X"B8",X"D2",X"0E",X"12",X"CD",X"67",X"1A",X"C3",X"0C",X"13",X"21",X"24",
		X"20",X"34",X"CD",X"5F",X"1A",X"C3",X"0C",X"13",X"2E",X"24",X"CD",X"52",X"1A",X"7E",X"FE",X"06",
		X"D2",X"24",X"12",X"C9",X"E5",X"3A",X"1D",X"20",X"A7",X"D3",X"06",X"C2",X"25",X"12",X"E1",X"36",
		X"00",X"CD",X"0D",X"19",X"CD",X"4C",X"00",X"21",X"7B",X"20",X"34",X"21",X"00",X"46",X"11",X"00",
		X"20",X"06",X"31",X"CD",X"8B",X"03",X"21",X"35",X"46",X"11",X"35",X"20",X"06",X"46",X"CD",X"8B",
		X"03",X"21",X"81",X"46",X"11",X"81",X"20",X"06",X"3F",X"CD",X"8B",X"03",X"21",X"14",X"20",X"34",
		X"CD",X"1E",X"14",X"CD",X"52",X"1A",X"2E",X"26",X"34",X"7E",X"47",X"0F",X"DA",X"71",X"12",X"2B",
		X"34",X"78",X"FE",X"08",X"CC",X"13",X"13",X"FE",X"0F",X"CC",X"13",X"13",X"CD",X"AD",X"12",X"CD",
		X"07",X"13",X"23",X"23",X"5E",X"23",X"56",X"21",X"09",X"20",X"73",X"23",X"72",X"3E",X"30",X"CD",
		X"D5",X"14",X"21",X"05",X"20",X"34",X"7E",X"A7",X"D3",X"06",X"C2",X"96",X"12",X"21",X"7B",X"20",
		X"36",X"00",X"2E",X"2F",X"34",X"2E",X"14",X"36",X"00",X"CD",X"78",X"1A",X"C9",X"CD",X"52",X"1A",
		X"2E",X"25",X"7E",X"FE",X"0B",X"DA",X"BB",X"12",X"3E",X"03",X"77",X"47",X"FE",X"07",X"DA",X"C3",
		X"12",X"06",X"06",X"3E",X"18",X"D6",X"03",X"05",X"C2",X"C5",X"12",X"4F",X"CD",X"07",X"13",X"23",
		X"23",X"EB",X"69",X"26",X"27",X"CD",X"00",X"03",X"2E",X"25",X"CD",X"52",X"1A",X"7E",X"0F",X"0F",
		X"11",X"E8",X"44",X"DA",X"E9",X"12",X"11",X"F8",X"44",X"CD",X"07",X"13",X"CD",X"EF",X"02",X"CD",
		X"07",X"13",X"7E",X"0F",X"0F",X"01",X"20",X"00",X"DA",X"FE",X"12",X"01",X"E0",X"FF",X"21",X"28",
		X"21",X"71",X"23",X"70",X"C3",X"BC",X"00",X"2E",X"04",X"C3",X"52",X"1A",X"2E",X"24",X"CD",X"52",
		X"1A",X"34",X"C9",X"F5",X"3E",X"FF",X"CD",X"04",X"02",X"3E",X"04",X"CD",X"FB",X"01",X"CD",X"C1",
		X"00",X"3E",X"20",X"CD",X"FB",X"01",X"CD",X"83",X"1A",X"CD",X"BC",X"00",X"CD",X"69",X"13",X"3E",
		X"04",X"CD",X"04",X"02",X"2E",X"26",X"CD",X"52",X"1A",X"7E",X"0F",X"DA",X"49",X"13",X"21",X"12",
		X"30",X"11",X"14",X"40",X"06",X"04",X"C3",X"51",X"13",X"21",X"12",X"2D",X"11",X"18",X"40",X"06",
		X"0A",X"CD",X"60",X"02",X"CD",X"B6",X"00",X"CD",X"4C",X"00",X"3E",X"80",X"CD",X"D5",X"14",X"CD",
		X"92",X"13",X"21",X"30",X"20",X"36",X"00",X"F1",X"C9",X"21",X"03",X"24",X"22",X"2D",X"21",X"21",
		X"1C",X"40",X"22",X"2F",X"21",X"0E",X"71",X"C5",X"2A",X"2D",X"21",X"CD",X"BB",X"13",X"22",X"2D",
		X"21",X"2A",X"2F",X"21",X"CD",X"CF",X"13",X"22",X"2F",X"21",X"C1",X"0D",X"C2",X"77",X"13",X"CD",
		X"FC",X"00",X"0E",X"79",X"21",X"1C",X"33",X"22",X"2D",X"21",X"21",X"03",X"32",X"22",X"2F",X"21",
		X"C5",X"AF",X"2A",X"2D",X"21",X"CD",X"D1",X"13",X"22",X"2D",X"21",X"AF",X"2A",X"2F",X"21",X"CD",
		X"BD",X"13",X"22",X"2F",X"21",X"C1",X"0D",X"C2",X"A0",X"13",X"C9",X"3E",X"FF",X"06",X"1A",X"E5",
		X"77",X"23",X"CD",X"E3",X"13",X"05",X"C2",X"C0",X"13",X"E1",X"11",X"20",X"00",X"19",X"C9",X"3E",
		X"FF",X"06",X"1A",X"E5",X"77",X"2B",X"CD",X"E3",X"13",X"05",X"C2",X"D4",X"13",X"E1",X"11",X"E0",
		X"FF",X"19",X"C9",X"1E",X"20",X"D3",X"06",X"1D",X"C2",X"E5",X"13",X"C9",X"DB",X"02",X"E6",X"04",
		X"C8",X"3A",X"03",X"20",X"A7",X"C0",X"31",X"00",X"24",X"06",X"04",X"C5",X"CD",X"1E",X"14",X"C1",
		X"05",X"C2",X"FB",X"13",X"3E",X"01",X"32",X"03",X"20",X"CD",X"B6",X"00",X"FB",X"11",X"22",X"40",
		X"21",X"16",X"30",X"06",X"04",X"CD",X"60",X"02",X"CD",X"C1",X"00",X"C3",X"18",X"00",X"21",X"03",
		X"24",X"01",X"DF",X"1A",X"C5",X"E5",X"36",X"00",X"23",X"05",X"C2",X"26",X"14",X"E1",X"11",X"20",
		X"00",X"19",X"C1",X"0D",X"C2",X"24",X"14",X"C9",X"CD",X"50",X"0C",X"E6",X"10",X"CA",X"4D",X"14",
		X"21",X"14",X"20",X"AF",X"BE",X"C0",X"23",X"BE",X"C0",X"34",X"23",X"34",X"C9",X"21",X"15",X"20",
		X"36",X"00",X"C9",X"21",X"16",X"20",X"AF",X"BE",X"C8",X"23",X"BE",X"C2",X"69",X"14",X"34",X"2A",
		X"33",X"20",X"01",X"10",X"05",X"09",X"22",X"1A",X"20",X"2A",X"1A",X"20",X"CD",X"C3",X"08",X"2A",
		X"1A",X"20",X"3A",X"54",X"20",X"A7",X"7D",X"C2",X"88",X"14",X"FE",X"E0",X"D2",X"8D",X"14",X"C6",
		X"03",X"6F",X"22",X"1A",X"20",X"C3",X"CB",X"08",X"FE",X"C0",X"C3",X"7C",X"14",X"2A",X"1A",X"20",
		X"22",X"BD",X"20",X"21",X"BB",X"20",X"34",X"21",X"16",X"46",X"11",X"16",X"20",X"06",X"07",X"C3",
		X"8B",X"03",X"21",X"BB",X"20",X"AF",X"BE",X"C8",X"23",X"BE",X"C2",X"BD",X"14",X"34",X"2A",X"BD",
		X"20",X"11",X"CD",X"14",X"01",X"08",X"01",X"CD",X"76",X"03",X"C3",X"D5",X"01",X"AF",X"77",X"2B",
		X"77",X"2A",X"BD",X"20",X"01",X"08",X"01",X"CD",X"76",X"03",X"C3",X"8C",X"08",X"A9",X"5C",X"BE",
		X"7F",X"FE",X"7F",X"7E",X"95",X"32",X"00",X"20",X"3A",X"00",X"20",X"A7",X"D3",X"06",X"C2",X"D8",
		X"14",X"C9",X"21",X"82",X"20",X"AF",X"BE",X"C8",X"3A",X"1A",X"20",X"D6",X"08",X"21",X"83",X"20",
		X"BE",X"D0",X"C6",X"12",X"BE",X"D8",X"3A",X"1B",X"20",X"23",X"D6",X"03",X"BE",X"D0",X"C6",X"09",
		X"BE",X"D8",X"2A",X"83",X"20",X"22",X"8D",X"20",X"CD",X"5B",X"0A",X"21",X"82",X"20",X"36",X"00",
		X"21",X"8B",X"20",X"34",X"C9",X"21",X"82",X"20",X"AF",X"BE",X"C8",X"23",X"5E",X"23",X"56",X"EB",
		X"E5",X"CD",X"5B",X"0A",X"E1",X"11",X"F9",X"FF",X"19",X"22",X"83",X"20",X"7D",X"FE",X"18",X"D2",
		X"42",X"0A",X"22",X"87",X"20",X"21",X"85",X"20",X"36",X"FF",X"21",X"82",X"20",X"36",X"00",X"C9",
		X"21",X"85",X"20",X"AF",X"BE",X"C8",X"23",X"34",X"7E",X"FE",X"01",X"CA",X"83",X"15",X"FE",X"04",
		X"C2",X"59",X"15",X"11",X"24",X"44",X"C3",X"86",X"15",X"FE",X"07",X"D8",X"11",X"3C",X"44",X"CD",
		X"86",X"15",X"21",X"00",X"00",X"22",X"81",X"20",X"22",X"85",X"20",X"CD",X"E0",X"15",X"21",X"88",
		X"20",X"D2",X"7A",X"15",X"CD",X"E7",X"15",X"C3",X"7D",X"15",X"CD",X"07",X"16",X"21",X"14",X"20",
		X"36",X"00",X"C9",X"11",X"0C",X"44",X"2A",X"87",X"20",X"CD",X"76",X"03",X"01",X"0C",X"02",X"C3",
		X"D5",X"01",X"21",X"8B",X"20",X"AF",X"BE",X"C8",X"23",X"34",X"7E",X"FE",X"01",X"CA",X"CE",X"15",
		X"FE",X"04",X"C2",X"AB",X"15",X"11",X"B4",X"44",X"C3",X"D1",X"15",X"FE",X"07",X"D8",X"2A",X"8D",
		X"20",X"CD",X"76",X"03",X"01",X"10",X"02",X"CD",X"8C",X"08",X"21",X"00",X"00",X"22",X"8B",X"20",
		X"21",X"81",X"20",X"36",X"00",X"CD",X"6F",X"1A",X"CD",X"D7",X"15",X"C3",X"7D",X"15",X"11",X"94",
		X"44",X"2A",X"8D",X"20",X"C3",X"89",X"15",X"CD",X"E0",X"15",X"DA",X"ED",X"15",X"C3",X"0D",X"16",
		X"CD",X"07",X"13",X"7E",X"0F",X"0F",X"C9",X"AF",X"3A",X"34",X"20",X"BE",X"D0",X"21",X"80",X"20",
		X"34",X"7E",X"FE",X"03",X"DA",X"FF",X"15",X"36",X"00",X"3E",X"E8",X"2B",X"86",X"77",X"C9",X"FE",
		X"02",X"3E",X"F0",X"DA",X"FB",X"15",X"C9",X"AF",X"3A",X"34",X"20",X"BE",X"D8",X"21",X"7E",X"20",
		X"34",X"7E",X"FE",X"03",X"DA",X"1F",X"16",X"36",X"00",X"3E",X"15",X"2B",X"86",X"77",X"C9",X"FE",
		X"02",X"3E",X"0D",X"DA",X"1B",X"16",X"C9",X"21",X"91",X"20",X"AF",X"BE",X"C8",X"23",X"34",X"7E",
		X"FE",X"01",X"CA",X"BA",X"16",X"FE",X"04",X"CA",X"C9",X"16",X"FE",X"07",X"D8",X"CD",X"CF",X"16",
		X"21",X"00",X"00",X"22",X"91",X"20",X"CD",X"5F",X"1A",X"21",X"95",X"20",X"34",X"7E",X"FE",X"03",
		X"D2",X"5E",X"16",X"3E",X"50",X"32",X"C2",X"20",X"CD",X"8C",X"02",X"C3",X"7D",X"15",X"CD",X"88",
		X"16",X"21",X"C1",X"20",X"70",X"78",X"C6",X"20",X"CD",X"2E",X"03",X"2A",X"93",X"20",X"CD",X"76",
		X"03",X"CD",X"45",X"03",X"11",X"34",X"04",X"CD",X"45",X"03",X"11",X"34",X"04",X"CD",X"45",X"03",
		X"21",X"96",X"20",X"34",X"23",X"36",X"0A",X"C9",X"3A",X"01",X"20",X"0F",X"0F",X"06",X"03",X"0F",
		X"D8",X"06",X"05",X"0F",X"D8",X"06",X"07",X"0F",X"D8",X"06",X"09",X"C9",X"21",X"96",X"20",X"AF",
		X"BE",X"C8",X"23",X"BE",X"CA",X"A9",X"16",X"35",X"C9",X"CD",X"8C",X"02",X"01",X"18",X"01",X"CD",
		X"D2",X"16",X"21",X"96",X"20",X"36",X"00",X"C3",X"7D",X"15",X"11",X"94",X"44",X"2A",X"93",X"20",
		X"CD",X"76",X"03",X"01",X"10",X"02",X"C3",X"D5",X"01",X"11",X"B4",X"44",X"C3",X"BD",X"16",X"01",
		X"10",X"02",X"2A",X"93",X"20",X"CD",X"76",X"03",X"C3",X"8C",X"08",X"21",X"81",X"20",X"AF",X"BE",
		X"C0",X"CD",X"07",X"13",X"E5",X"7E",X"FE",X"FF",X"C2",X"ED",X"16",X"E1",X"C9",X"07",X"DA",X"F9",
		X"16",X"E1",X"23",X"23",X"23",X"23",X"C3",X"E4",X"16",X"E1",X"E5",X"CD",X"40",X"0D",X"4D",X"44",
		X"CD",X"E0",X"15",X"21",X"7F",X"20",X"DA",X"2F",X"17",X"2E",X"7D",X"7E",X"B8",X"D2",X"F1",X"16",
		X"C6",X"04",X"B8",X"DA",X"F1",X"16",X"21",X"83",X"20",X"71",X"23",X"78",X"FE",X"30",X"DA",X"F1",
		X"16",X"FE",X"F0",X"D2",X"F1",X"16",X"70",X"21",X"FF",X"FF",X"22",X"81",X"20",X"E1",X"C9",X"7E",
		X"B8",X"D2",X"F1",X"16",X"C6",X"06",X"B8",X"DA",X"F1",X"16",X"C3",X"16",X"17",X"3A",X"AA",X"20",
		X"A7",X"C8",X"21",X"A2",X"20",X"CD",X"F0",X"0D",X"CD",X"5D",X"17",X"21",X"AE",X"20",X"35",X"7E",
		X"A7",X"C2",X"57",X"17",X"C3",X"82",X"17",X"21",X"A0",X"20",X"C3",X"A1",X"0D",X"7D",X"E6",X"07",
		X"D3",X"02",X"CD",X"76",X"03",X"C5",X"E5",X"1A",X"D3",X"04",X"DB",X"03",X"B6",X"77",X"23",X"13",
		X"AF",X"D3",X"04",X"DB",X"03",X"B6",X"77",X"E1",X"01",X"20",X"00",X"09",X"C1",X"05",X"C2",X"65",
		X"17",X"C9",X"2A",X"A8",X"20",X"EB",X"1A",X"2A",X"AF",X"20",X"2D",X"CA",X"BA",X"17",X"22",X"AF",
		X"20",X"32",X"AE",X"20",X"13",X"1A",X"E6",X"0F",X"07",X"01",X"BF",X"17",X"26",X"00",X"6F",X"09",
		X"E5",X"C1",X"21",X"A0",X"20",X"0A",X"77",X"03",X"23",X"0A",X"77",X"13",X"1A",X"6F",X"13",X"1A",
		X"67",X"22",X"A2",X"20",X"EB",X"23",X"22",X"A8",X"20",X"C9",X"AF",X"32",X"AA",X"20",X"C9",X"00",
		X"02",X"02",X"02",X"02",X"00",X"02",X"FE",X"00",X"FE",X"FE",X"FE",X"FE",X"00",X"FE",X"02",X"01",
		X"02",X"02",X"01",X"02",X"FF",X"01",X"FE",X"FF",X"FE",X"FE",X"FF",X"FE",X"01",X"FF",X"02",X"FF",
		X"FF",X"24",X"06",X"D7",X"30",X"10",X"00",X"D7",X"30",X"04",X"07",X"D7",X"50",X"0A",X"06",X"CF",
		X"58",X"04",X"05",X"BC",X"58",X"04",X"07",X"B4",X"50",X"0A",X"06",X"AC",X"58",X"04",X"05",X"98");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
