library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity MRDONIGHTMARE_1K is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of MRDONIGHTMARE_1K is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",X"00",X"02",X"02",X"FE",X"FE",X"42",X"02",X"00",X"00",
		X"62",X"F2",X"BA",X"9A",X"9E",X"CE",X"46",X"00",X"8C",X"DE",X"F2",X"B2",X"92",X"86",X"04",X"00",
		X"08",X"FE",X"FE",X"C8",X"68",X"38",X"18",X"00",X"1C",X"BE",X"A2",X"A2",X"A2",X"E6",X"E4",X"00",
		X"0C",X"9E",X"92",X"92",X"D2",X"7E",X"3C",X"00",X"C0",X"E0",X"B0",X"9E",X"8E",X"C0",X"C0",X"00",
		X"0C",X"6E",X"9A",X"9A",X"B2",X"F2",X"6C",X"00",X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",X"00",
		X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",
		X"44",X"C6",X"82",X"82",X"C6",X"7C",X"38",X"00",X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",
		X"82",X"92",X"92",X"92",X"FE",X"FE",X"00",X"00",X"80",X"90",X"90",X"90",X"90",X"FE",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",
		X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",X"44",X"C6",X"82",X"82",X"C6",X"7C",X"38",X"00",
		X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",X"82",X"92",X"92",X"92",X"FE",X"FE",X"00",X"00",
		X"80",X"90",X"90",X"90",X"90",X"FE",X"FE",X"00",X"9E",X"9E",X"92",X"82",X"C6",X"7C",X"38",X"00",
		X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",X"82",X"82",X"FE",X"FE",X"82",X"82",X"00",X"00",
		X"FC",X"FE",X"02",X"02",X"02",X"06",X"04",X"00",X"82",X"C6",X"6E",X"3C",X"18",X"FE",X"FE",X"00",
		X"02",X"02",X"02",X"02",X"FE",X"FE",X"00",X"00",X"FE",X"FE",X"70",X"38",X"70",X"FE",X"FE",X"00",
		X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",X"00",
		X"70",X"F8",X"88",X"88",X"88",X"FE",X"FE",X"00",X"7A",X"FC",X"8E",X"8A",X"82",X"FE",X"7C",X"00",
		X"72",X"F6",X"9E",X"8C",X"88",X"FE",X"FE",X"00",X"0C",X"5E",X"D2",X"92",X"92",X"F6",X"64",X"00",
		X"80",X"80",X"FE",X"FE",X"80",X"80",X"00",X"00",X"FC",X"FE",X"02",X"02",X"02",X"FE",X"FC",X"00",
		X"F0",X"F8",X"1C",X"0E",X"1C",X"F8",X"F0",X"00",X"F8",X"FE",X"1C",X"38",X"1C",X"FE",X"F8",X"00",
		X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",X"C0",X"F0",X"1E",X"1E",X"F0",X"C0",X"00",X"00",
		X"C2",X"E2",X"F2",X"BA",X"9E",X"8E",X"86",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"30",X"42",X"23",X"03",X"42",X"60",X"42",X"40",X"08",X"20",X"80",X"00",X"08",X"84",X"00",
		X"20",X"41",X"22",X"40",X"42",X"23",X"18",X"05",X"82",X"84",X"88",X"00",X"80",X"E0",X"08",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"3C",X"7E",X"66",X"5A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"7E",X"7E",X"7E",X"3C",X"18",X"00",X"00",
		X"00",X"00",X"00",X"02",X"07",X"17",X"0B",X"88",X"00",X"00",X"18",X"0C",X"46",X"6E",X"6E",X"06",
		X"F8",X"08",X"10",X"00",X"00",X"00",X"00",X"00",X"0E",X"1E",X"06",X"0E",X"0C",X"18",X"00",X"00",
		X"00",X"00",X"00",X"03",X"05",X"05",X"1A",X"1C",X"00",X"00",X"00",X"00",X"80",X"C0",X"60",X"30",
		X"0B",X"0D",X"12",X"0A",X"03",X"02",X"00",X"00",X"C0",X"A0",X"40",X"80",X"00",X"00",X"00",X"00",
		X"03",X"07",X"3F",X"7F",X"4F",X"4F",X"3F",X"1F",X"FE",X"FF",X"9F",X"DE",X"DC",X"9C",X"BE",X"BF",
		X"1F",X"3F",X"4F",X"4F",X"7F",X"3F",X"07",X"03",X"BF",X"BE",X"9C",X"DC",X"DE",X"9F",X"FF",X"FE",
		X"FF",X"FF",X"FF",X"7F",X"4F",X"AB",X"05",X"02",X"A0",X"D8",X"FA",X"FC",X"FE",X"FE",X"FE",X"BE",
		X"00",X"00",X"60",X"28",X"64",X"7A",X"7E",X"7F",X"4F",X"27",X"0B",X"02",X"00",X"00",X"80",X"00",
		X"00",X"FF",X"F7",X"BF",X"FF",X"00",X"FF",X"FE",X"00",X"FF",X"F3",X"5F",X"FF",X"00",X"FF",X"FF",
		X"D7",X"FF",X"00",X"FF",X"FB",X"9E",X"FF",X"00",X"DB",X"FF",X"00",X"FF",X"DF",X"FD",X"FF",X"00",
		X"80",X"80",X"C0",X"C0",X"80",X"80",X"80",X"40",X"03",X"02",X"02",X"02",X"06",X"02",X"02",X"02",
		X"60",X"60",X"40",X"40",X"40",X"70",X"40",X"C0",X"06",X"06",X"02",X"03",X"01",X"01",X"01",X"01",
		X"00",X"02",X"00",X"00",X"04",X"03",X"2B",X"07",X"00",X"DE",X"18",X"80",X"08",X"40",X"90",X"80",
		X"0F",X"29",X"0F",X"06",X"00",X"00",X"00",X"00",X"94",X"00",X"22",X"02",X"02",X"32",X"00",X"00",
		X"00",X"10",X"00",X"00",X"08",X"23",X"0B",X"07",X"00",X"00",X"00",X"00",X"00",X"44",X"94",X"80",
		X"2F",X"09",X"0F",X"06",X"00",X"00",X"00",X"00",X"88",X"22",X"02",X"12",X"02",X"30",X"00",X"00",
		X"00",X"20",X"00",X"00",X"08",X"03",X"2B",X"07",X"00",X"30",X"00",X"20",X"00",X"12",X"82",X"A2",
		X"2F",X"09",X"0F",X"06",X"00",X"00",X"00",X"00",X"8A",X"22",X"08",X"48",X"08",X"C8",X"00",X"00",
		X"00",X"3C",X"01",X"00",X"21",X"24",X"00",X"01",X"00",X"02",X"02",X"16",X"46",X"00",X"22",X"CA",
		X"07",X"0D",X"0D",X"07",X"00",X"02",X"00",X"00",X"E0",X"E2",X"90",X"40",X"00",X"40",X"00",X"00",
		X"00",X"1E",X"00",X"01",X"28",X"22",X"00",X"01",X"00",X"00",X"60",X"00",X"40",X"00",X"40",X"C0",
		X"07",X"0D",X"0D",X"07",X"00",X"01",X"00",X"00",X"E0",X"E0",X"80",X"50",X"02",X"20",X"00",X"00",
		X"00",X"03",X"00",X"3D",X"00",X"02",X"28",X"21",X"00",X"E0",X"00",X"00",X"22",X"8A",X"00",X"C0",
		X"07",X"0D",X"0D",X"07",X"00",X"01",X"00",X"00",X"E0",X"E0",X"80",X"50",X"00",X"42",X"00",X"00",
		X"00",X"E0",X"60",X"E0",X"C0",X"00",X"E0",X"60",X"00",X"07",X"03",X"05",X"07",X"00",X"03",X"05",
		X"E0",X"E0",X"00",X"E0",X"A0",X"E0",X"C0",X"00",X"07",X"07",X"00",X"07",X"06",X"03",X"03",X"00",
		X"00",X"00",X"00",X"04",X"0E",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"0E",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"07",X"02",X"00",X"00",X"00",X"00",X"30",X"08",X"04",X"00",X"00",
		X"00",X"00",X"04",X"0E",X"04",X"00",X"00",X"00",X"00",X"04",X"08",X"10",X"20",X"00",X"00",X"00",
		X"00",X"00",X"1A",X"36",X"36",X"3E",X"1E",X"0E",X"00",X"00",X"38",X"3C",X"38",X"30",X"38",X"3C",
		X"1E",X"36",X"36",X"3F",X"1B",X"01",X"00",X"00",X"3C",X"38",X"30",X"78",X"FC",X"F8",X"00",X"00",
		X"00",X"00",X"34",X"4C",X"4C",X"7C",X"3C",X"1C",X"00",X"00",X"0E",X"0C",X"08",X"0E",X"0C",X"08",
		X"3C",X"4C",X"4C",X"7E",X"37",X"03",X"00",X"00",X"08",X"0C",X"0E",X"18",X"FC",X"FE",X"00",X"00",
		X"43",X"30",X"0C",X"03",X"00",X"00",X"00",X"00",X"8C",X"43",X"20",X"43",X"8C",X"90",X"90",X"8C",
		X"17",X"10",X"30",X"40",X"83",X"8C",X"90",X"90",X"14",X"12",X"09",X"09",X"13",X"14",X"14",X"14",
		X"90",X"90",X"88",X"47",X"20",X"11",X"12",X"14",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"44",X"88",X"90",X"90",X"90",X"90",X"90",X"90",X"00",X"00",X"01",X"02",X"04",X"08",X"11",X"22",
		X"00",X"00",X"11",X"3B",X"3F",X"3F",X"00",X"00",X"00",X"00",X"88",X"DC",X"FC",X"FC",X"1C",X"0C",
		X"00",X"3F",X"1F",X"27",X"3E",X"1C",X"00",X"00",X"1C",X"F8",X"F0",X"98",X"F8",X"70",X"00",X"00",
		X"00",X"24",X"36",X"3F",X"00",X"00",X"00",X"00",X"00",X"24",X"6C",X"FC",X"1C",X"0C",X"0C",X"0C",
		X"00",X"00",X"3F",X"1F",X"27",X"26",X"1C",X"00",X"0C",X"1C",X"F8",X"F0",X"98",X"98",X"70",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"0F",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",
		X"0F",X"0F",X"07",X"03",X"00",X"00",X"00",X"00",X"E0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"03",X"00",X"38",X"7C",X"72",X"7E",X"7E",X"72",X"02",X"02",X"02",X"02",X"94",X"00",X"A0",X"00",
		X"7C",X"38",X"02",X"00",X"20",X"09",X"00",X"09",X"A0",X"00",X"20",X"0C",X"04",X"84",X"04",X"00",
		X"00",X"00",X"00",X"01",X"0B",X"03",X"2B",X"03",X"00",X"78",X"00",X"C0",X"E0",X"90",X"F0",X"F4",
		X"0B",X"23",X"09",X"00",X"04",X"00",X"00",X"0F",X"94",X"E0",X"C0",X"00",X"28",X"08",X"00",X"80",
		X"1F",X"38",X"20",X"08",X"00",X"05",X"00",X"01",X"0C",X"00",X"04",X"00",X"38",X"7C",X"72",X"7E",
		X"44",X"51",X"44",X"60",X"20",X"20",X"00",X"00",X"7E",X"72",X"7C",X"38",X"00",X"08",X"00",X"0C",
		X"03",X"00",X"00",X"00",X"00",X"70",X"51",X"50",X"CC",X"00",X"04",X"80",X"38",X"7C",X"72",X"7E",
		X"51",X"50",X"71",X"00",X"00",X"00",X"00",X"03",X"7E",X"72",X"7C",X"38",X"00",X"88",X"00",X"CC",
		X"3C",X"7E",X"FE",X"7E",X"FE",X"FC",X"FE",X"F6",X"48",X"50",X"50",X"49",X"26",X"10",X"0C",X"03",
		X"00",X"00",X"00",X"00",X"03",X"0C",X"10",X"27",X"7E",X"FE",X"FE",X"EC",X"FE",X"FE",X"7C",X"00",
		X"00",X"E0",X"18",X"06",X"C1",X"30",X"0C",X"03",X"00",X"00",X"C0",X"00",X"01",X"06",X"08",X"06",
		X"FE",X"06",X"18",X"E0",X"01",X"06",X"08",X"06",X"20",X"40",X"40",X"20",X"1F",X"00",X"00",X"00",
		X"1F",X"20",X"C0",X"00",X"00",X"C1",X"21",X"21",X"40",X"40",X"3F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"07",X"18",X"30",X"20",X"40",X"90",X"90",X"88",X"04",X"02",X"3C",X"C0",X"00",
		X"90",X"A0",X"A1",X"A1",X"A1",X"A1",X"A1",X"A0",X"C7",X"20",X"E0",X"00",X"03",X"04",X"08",X"90",
		X"A1",X"A1",X"A1",X"A0",X"20",X"20",X"10",X"08",X"0F",X"10",X"20",X"47",X"88",X"90",X"A0",X"A0",
		X"88",X"48",X"48",X"48",X"C8",X"08",X"10",X"E0",X"88",X"48",X"48",X"48",X"88",X"10",X"20",X"10",
		X"C8",X"48",X"48",X"48",X"88",X"10",X"20",X"10",X"E0",X"04",X"0F",X"08",X"C8",X"48",X"48",X"48",
		X"F8",X"04",X"02",X"02",X"E2",X"12",X"11",X"10",X"04",X"04",X"FC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"E0",X"10",X"08",X"04",X"04",X"7C",X"00",X"00",X"00",X"00",X"01",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"80",X"82",X"82",X"01",X"01",X"01",X"01",X"01",X"01",X"21",X"A1",
		X"82",X"83",X"80",X"80",X"80",X"80",X"80",X"FF",X"A1",X"E1",X"01",X"01",X"01",X"01",X"01",X"FF",
		X"80",X"80",X"80",X"80",X"80",X"80",X"83",X"80",X"01",X"01",X"01",X"01",X"01",X"01",X"61",X"81",
		X"80",X"83",X"80",X"80",X"80",X"80",X"80",X"80",X"81",X"61",X"01",X"01",X"01",X"01",X"01",X"01",
		X"80",X"80",X"80",X"80",X"80",X"80",X"82",X"82",X"F0",X"08",X"04",X"E2",X"11",X"09",X"05",X"05",
		X"83",X"82",X"82",X"80",X"80",X"80",X"80",X"80",X"E1",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"80",X"80",X"80",X"80",X"80",X"80",X"81",X"82",X"01",X"01",X"01",X"01",X"01",X"01",X"21",X"A1",
		X"82",X"83",X"80",X"80",X"80",X"80",X"80",X"80",X"C1",X"E1",X"01",X"01",X"01",X"01",X"01",X"01",
		X"FF",X"80",X"80",X"80",X"80",X"80",X"81",X"82",X"FF",X"01",X"01",X"01",X"01",X"01",X"E1",X"81",
		X"82",X"81",X"80",X"80",X"80",X"80",X"80",X"80",X"81",X"E1",X"01",X"01",X"01",X"01",X"01",X"01",
		X"80",X"80",X"80",X"80",X"80",X"80",X"82",X"82",X"01",X"01",X"01",X"01",X"01",X"01",X"21",X"A1",
		X"82",X"83",X"80",X"80",X"80",X"80",X"80",X"FF",X"A1",X"E1",X"01",X"01",X"01",X"01",X"01",X"FF",
		X"80",X"80",X"80",X"80",X"80",X"80",X"83",X"80",X"01",X"01",X"01",X"01",X"01",X"01",X"61",X"81",
		X"80",X"83",X"80",X"80",X"80",X"80",X"80",X"80",X"81",X"61",X"01",X"01",X"01",X"01",X"01",X"01",
		X"80",X"80",X"80",X"80",X"80",X"80",X"82",X"82",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"83",X"82",X"82",X"80",X"80",X"80",X"80",X"80",X"E1",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"80",X"80",X"80",X"80",X"80",X"80",X"81",X"82",X"01",X"01",X"01",X"01",X"01",X"01",X"21",X"A1",
		X"82",X"83",X"80",X"80",X"80",X"80",X"80",X"80",X"C1",X"E1",X"01",X"01",X"01",X"01",X"01",X"01",
		X"FF",X"80",X"80",X"80",X"80",X"80",X"81",X"82",X"FF",X"01",X"01",X"01",X"01",X"01",X"E1",X"81",
		X"82",X"81",X"80",X"80",X"80",X"80",X"80",X"80",X"81",X"E1",X"01",X"01",X"01",X"01",X"01",X"01",
		X"00",X"0F",X"38",X"70",X"70",X"60",X"60",X"70",X"00",X"E0",X"31",X"19",X"0B",X"0E",X"0C",X"08",
		X"70",X"60",X"60",X"70",X"70",X"38",X"0F",X"00",X"08",X"0C",X"0E",X"0B",X"19",X"31",X"E0",X"00",
		X"00",X"0F",X"38",X"70",X"70",X"43",X"47",X"74",X"00",X"E4",X"34",X"1C",X"0C",X"0C",X"8C",X"D8",
		X"74",X"46",X"42",X"70",X"70",X"38",X"0F",X"00",X"D8",X"0C",X"0E",X"0B",X"19",X"31",X"E0",X"00",
		X"00",X"0F",X"38",X"70",X"60",X"63",X"67",X"74",X"00",X"E0",X"31",X"19",X"0B",X"0E",X"8C",X"D8",
		X"74",X"66",X"62",X"60",X"70",X"38",X"0F",X"00",X"D8",X"0C",X"0C",X"0C",X"1C",X"34",X"E4",X"00",
		X"7C",X"82",X"01",X"01",X"01",X"01",X"01",X"82",X"E0",X"00",X"38",X"C7",X"00",X"00",X"00",X"00",
		X"23",X"24",X"24",X"C4",X"05",X"05",X"09",X"11",X"CF",X"30",X"00",X"8F",X"90",X"A0",X"A0",X"A0",
		X"02",X"04",X"F8",X"00",X"00",X"00",X"00",X"00",X"09",X"09",X"09",X"09",X"09",X"09",X"11",X"E1",
		X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"12",X"09",X"09",X"09",X"09",X"09",X"09",X"09",
		X"0A",X"12",X"14",X"24",X"48",X"88",X"C4",X"22",X"0A",X"09",X"09",X"05",X"05",X"05",X"09",X"09",
		X"E2",X"04",X"08",X"10",X"C8",X"24",X"14",X"12",X"05",X"85",X"85",X"85",X"05",X"05",X"09",X"11",
		X"09",X"30",X"42",X"23",X"02",X"40",X"63",X"40",X"48",X"04",X"02",X"E2",X"00",X"02",X"E0",X"02",
		X"23",X"40",X"23",X"40",X"42",X"23",X"18",X"05",X"62",X"80",X"62",X"02",X"A0",X"E2",X"00",X"24",
		X"00",X"10",X"70",X"E0",X"E0",X"C0",X"C0",X"E0",X"00",X"08",X"09",X"05",X"05",X"07",X"06",X"04",
		X"E0",X"C0",X"C0",X"E0",X"E0",X"70",X"10",X"00",X"04",X"06",X"07",X"05",X"05",X"09",X"08",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
