library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity obj_7m is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of obj_7m is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0D",X"00",X"0F",X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",X"1F",X"1F",X"0F",X"07",X"07",X"0F",X"06",X"0D",
		X"00",X"00",X"00",X"07",X"0F",X"0F",X"0F",X"4F",X"EF",X"FF",X"7F",X"3F",X"07",X"0F",X"06",X"0D",
		X"00",X"00",X"1E",X"1F",X"1F",X"1F",X"1F",X"3F",X"7F",X"7F",X"3F",X"0A",X"07",X"0F",X"06",X"0D",
		X"00",X"00",X"3C",X"3F",X"1F",X"4F",X"EF",X"EF",X"FF",X"7F",X"3F",X"0F",X"07",X"0F",X"07",X"0E",
		X"00",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"07",X"17",X"3F",X"3F",X"3F",X"1F",X"07",X"07",X"03",X"07",X"03",X"06",X"06",
		X"00",X"00",X"0C",X"0F",X"07",X"07",X"07",X"07",X"07",X"07",X"03",X"03",X"07",X"03",X"06",X"06",
		X"00",X"00",X"00",X"1F",X"1F",X"4F",X"FF",X"FF",X"7F",X"0F",X"1D",X"1B",X"00",X"0F",X"07",X"00",
		X"34",X"06",X"3F",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"06",X"0F",X"0F",X"07",X"0F",X"4F",X"EF",X"FF",X"7F",X"3F",X"1F",X"3F",X"1A",X"37",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"2D",X"6F",X"63",X"FD",X"FF",X"FD",X"F9",X"2D",X"2D",X"2D",X"0D",X"04",X"01",X"01",X"01",
		X"35",X"04",X"3F",X"1F",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"27",X"EF",X"FF",X"EF",X"FF",X"FF",X"7F",X"3F",X"1F",X"3F",X"1A",X"37",
		X"00",X"00",X"00",X"03",X"27",X"EF",X"FF",X"EF",X"FF",X"FF",X"7F",X"3F",X"1F",X"3F",X"1A",X"37",
		X"00",X"00",X"00",X"03",X"27",X"EF",X"FF",X"EF",X"EF",X"FF",X"7F",X"3F",X"1F",X"3F",X"1A",X"37",
		X"00",X"3C",X"3F",X"3F",X"1F",X"DF",X"FE",X"FF",X"7F",X"0F",X"06",X"0D",X"0D",X"00",X"0F",X"07",
		X"00",X"3F",X"3F",X"DF",X"FE",X"FF",X"3F",X"0F",X"1D",X"1B",X"00",X"0F",X"07",X"00",X"00",X"00",
		X"0F",X"0F",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"07",X"1F",X"1F",X"3D",X"3F",X"3F",X"0F",X"0B",X"1F",X"1C",X"39",X"F9",X"ED",X"24",X"04",
		X"03",X"07",X"1F",X"1F",X"3D",X"BF",X"FF",X"EF",X"7B",X"7F",X"3C",X"19",X"09",X"0D",X"04",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"EE",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"00",X"1F",X"3F",X"3F",X"3F",X"1F",X"1F",X"4F",X"FF",X"FF",X"FF",X"03",X"03",
		X"06",X"06",X"06",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",X"7F",X"FF",X"FF",X"6F",X"06",X"0D",
		X"00",X"00",X"02",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"03",X"07",X"03",X"06",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0E",X"1D",X"3F",X"33",X"60",X"60",X"60",X"60",X"60",X"60",X"30",X"38",X"1C",X"0F",X"07",
		X"6B",X"DE",X"0B",X"12",X"43",X"07",X"07",X"05",X"17",X"06",X"0D",X"0B",X"0B",X"1B",X"17",X"0F",
		X"0D",X"0F",X"1F",X"3F",X"31",X"60",X"60",X"60",X"60",X"60",X"60",X"30",X"38",X"1C",X"0F",X"07",
		X"FC",X"75",X"22",X"17",X"07",X"27",X"86",X"0D",X"0B",X"0B",X"0B",X"17",X"17",X"0F",X"0F",X"0E",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",X"00",X"00",X"00",
		X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",X"FE",X"7E",X"7E",X"3E",X"1E",X"06",X"00",X"00",X"00",X"00",
		X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",X"FE",X"7E",X"7E",X"3E",X"1E",X"06",X"00",X"00",X"00",X"00",
		X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",X"FE",X"7E",X"7E",X"3E",X"1E",X"06",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"FC",X"FC",X"FC",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FC",X"FC",X"FC",
		X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",X"FE",X"7E",X"3E",X"7E",X"FE",X"FE",X"FC",X"FC",X"FC",X"FC",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",X"FE",X"7E",X"7E",X"3E",X"1E",X"06",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"00",X"00",X"00",X"00",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"00",X"00",X"00",X"00",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"4E",X"0E",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"00",X"00",X"40",X"40",X"4E",X"0E",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"00",X"00",X"40",X"40",X"4E",X"0E",X"0E",
		X"00",X"00",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"4E",X"0E",X"0E",
		X"00",X"00",X"02",X"02",X"00",X"00",X"00",X"02",X"02",X"00",X"00",X"40",X"40",X"4E",X"0E",X"0E",
		X"00",X"00",X"02",X"02",X"00",X"40",X"40",X"4E",X"0E",X"00",X"00",X"40",X"40",X"4E",X"0E",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FE",X"FE",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"4E",X"4E",X"4E",X"4E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"4F",X"4F",X"4F",X"4F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"00",X"00",X"00",X"00",X"06",X"1E",X"3E",X"7E",X"7E",X"FE",X"FE",X"FE",X"FC",X"FC",X"FC",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"AA",X"AA",X"AA",X"AA",X"44",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"31",X"4A",X"4A",X"4A",X"4A",X"31",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"31",X"4A",X"4A",X"4A",X"4A",X"31",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"31",X"4A",X"4A",X"4A",X"4A",X"31",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"31",X"4A",X"4A",X"4A",X"4A",X"31",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"55",X"55",X"55",X"55",X"22",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"55",X"55",X"55",X"55",X"22",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"AA",X"AA",X"AA",X"AA",X"44",X"00",X"00",
		X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"13",X"17",X"3F",X"3F",X"FF",X"3C",X"3B",X"0C",X"0F",X"0F",X"08",X"03",X"D3",X"DD",X"4F",X"07",
		X"13",X"17",X"3F",X"3F",X"FF",X"BC",X"FB",X"C4",X"0F",X"0F",X"08",X"03",X"03",X"1D",X"0F",X"07",
		X"07",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"04",X"44",X"9F",X"BF",X"BF",X"7F",X"1B",X"11",X"41",X"C1",X"C1",X"C1",X"03",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",
		X"01",X"01",X"01",X"01",X"03",X"03",X"0F",X"FE",X"F8",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"07",X"0F",X"1F",X"1F",X"3F",X"BF",X"7F",X"3F",X"7F",X"7F",X"F3",X"E7",X"4F",X"0E",X"06",X"00",
		X"07",X"0F",X"1F",X"1F",X"3F",X"3F",X"7F",X"BF",X"3F",X"3F",X"33",X"73",X"71",X"21",X"00",X"00",
		X"E0",X"7F",X"7F",X"FF",X"7F",X"FF",X"7F",X"3F",X"3F",X"1F",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"70",X"61",X"7F",X"7F",X"FF",X"7F",X"FF",X"7F",X"3F",X"3F",X"1F",X"0E",X"00",X"00",X"00",X"00",
		X"E3",X"7F",X"7F",X"FF",X"7F",X"FF",X"7F",X"3F",X"3F",X"1F",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"38",X"7F",X"7F",X"FF",X"7F",X"FF",X"7F",X"3F",X"3F",X"1F",X"0E",X"00",X"00",X"00",X"00",
		X"38",X"7F",X"7F",X"FF",X"FF",X"FF",X"7F",X"3F",X"3F",X"1F",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"1C",X"41",X"21",X"00",X"03",X"07",X"0E",X"0D",X"03",X"03",X"03",X"03",X"01",X"01",X"00",
		X"01",X"0D",X"0E",X"23",X"40",X"03",X"07",X"0E",X"0D",X"03",X"03",X"03",X"03",X"01",X"01",X"00",
		X"0E",X"1C",X"00",X"10",X"21",X"03",X"07",X"06",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",
		X"F4",X"72",X"30",X"00",X"00",X"00",X"CB",X"CB",X"7B",X"37",X"03",X"03",X"03",X"01",X"01",X"00",
		X"03",X"03",X"02",X"00",X"00",X"00",X"06",X"1D",X"3D",X"7B",X"F7",X"E7",X"67",X"26",X"02",X"01",
		X"01",X"07",X"0F",X"1F",X"1F",X"1F",X"0F",X"0F",X"03",X"3D",X"0F",X"07",X"34",X"7E",X"3F",X"0F",
		X"01",X"07",X"0F",X"1F",X"1F",X"1F",X"1F",X"0F",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"0F",X"1F",X"1F",X"3F",X"3F",X"3F",X"3F",X"7F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"0F",X"1F",X"1F",X"3F",X"3F",X"7F",X"3F",X"7F",X"7F",X"37",X"00",X"00",X"00",X"00",X"00",
		X"07",X"0F",X"1F",X"1F",X"3F",X"BF",X"7F",X"3F",X"7F",X"7F",X"73",X"27",X"01",X"00",X"00",X"00",
		X"01",X"03",X"0B",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"03",X"03",X"07",X"07",X"07",X"0F",X"0F",X"07",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"07",X"03",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"1F",X"1F",X"1F",X"1F",X"0F",X"03",X"01",
		X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"1F",X"1F",X"1F",X"1F",X"0F",X"03",X"01",X"00",X"00",
		X"00",X"00",X"01",X"07",X"0F",X"1F",X"1F",X"1F",X"1F",X"0F",X"03",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"44",X"62",X"61",X"30",X"32",X"14",X"18",X"1A",X"0A",X"03",X"03",X"01",X"01",
		X"20",X"11",X"0A",X"44",X"62",X"61",X"20",X"32",X"15",X"1B",X"1A",X"0A",X"02",X"02",X"01",X"01",
		X"20",X"30",X"58",X"48",X"62",X"61",X"20",X"30",X"10",X"00",X"10",X"08",X"00",X"02",X"01",X"01",
		X"00",X"30",X"08",X"00",X"42",X"40",X"40",X"70",X"00",X"00",X"00",X"42",X"62",X"03",X"08",X"00",
		X"20",X"20",X"08",X"00",X"00",X"80",X"40",X"00",X"00",X"00",X"00",X"80",X"40",X"00",X"02",X"11",
		X"4C",X"08",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"30",X"0C",X"03",X"01",X"07",X"7F",X"FF",X"3F",X"0F",X"03",X"00",
		X"00",X"00",X"00",X"00",X"80",X"40",X"20",X"F8",X"F7",X"F0",X"F0",X"F0",X"70",X"31",X"1B",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"01",X"03",X"07",X"0F",X"1F",X"3F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"80",X"60",X"10",X"0F",X"80",X"E0",X"F8",X"FF",X"7F",X"1F",X"07",
		X"00",X"00",X"00",X"00",X"00",X"80",X"60",X"18",X"07",X"80",X"E0",X"F8",X"FF",X"7F",X"1F",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"60",X"C0",X"80",X"FF",X"FF",X"7F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"EE",X"EE",X"EE",X"EE",X"0E",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"EE",X"EE",X"EE",X"EE",X"EE",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"0E",X"EE",X"EE",X"EE",X"EE",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"22",X"66",X"76",X"7F",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"22",X"66",X"76",X"7F",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"66",X"EE",X"FF",X"FF",X"FF",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"08",X"05",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"40",X"21",X"19",X"8B",X"6D",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"B1",X"69",X"16",X"36",X"30",X"27",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"81",X"63",X"9E",X"6D",X"21",X"74",X"86",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"30",X"0C",X"03",X"30",X"3C",X"7C",X"FC",X"3C",X"0E",X"03",X"00",
		X"00",X"00",X"00",X"00",X"80",X"40",X"20",X"98",X"C7",X"C0",X"C0",X"C3",X"63",X"23",X"1F",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"3C",X"3C",X"3C",X"7E",X"FF",
		X"00",X"03",X"0F",X"1F",X"1D",X"39",X"35",X"34",X"36",X"37",X"37",X"1B",X"1C",X"0F",X"03",X"00",
		X"00",X"00",X"00",X"01",X"03",X"03",X"23",X"37",X"3E",X"1E",X"1C",X"0F",X"07",X"03",X"00",X"00",
		X"00",X"03",X"0F",X"0C",X"19",X"1B",X"1B",X"1C",X"0F",X"03",X"00",X"00",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"0E",X"0E",X"1B",X"19",X"1A",X"1A",X"0C",X"0F",X"07",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"0B",X"0F",X"06",X"03",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"07",X"06",X"06",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"07",X"07",X"06",X"03",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"04",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"04",X"03",X"00",X"00",X"00",X"00",
		X"00",X"02",X"04",X"04",X"08",X"08",X"00",X"00",X"00",X"04",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"02",X"02",X"02",X"00",X"00",X"00",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"30",X"30",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"54",X"54",X"50",X"43",X"37",X"07",X"17",X"27",X"72",X"56",X"56",X"46",X"26",X"00",X"00",X"00",
		X"A4",X"A4",X"90",X"43",X"37",X"07",X"37",X"67",X"E2",X"A6",X"86",X"C6",X"06",X"00",X"00",X"00",
		X"04",X"A8",X"A8",X"50",X"43",X"17",X"07",X"37",X"27",X"72",X"2E",X"26",X"16",X"0E",X"00",X"00",
		X"A8",X"A8",X"9D",X"4D",X"35",X"25",X"57",X"E7",X"F7",X"52",X"56",X"05",X"37",X"07",X"04",X"08",
		X"54",X"54",X"2D",X"1D",X"05",X"05",X"37",X"67",X"C7",X"E2",X"F6",X"D5",X"57",X"67",X"34",X"18",
		X"24",X"48",X"4D",X"0D",X"35",X"05",X"77",X"C7",X"E7",X"F2",X"56",X"55",X"27",X"37",X"04",X"08",
		X"0E",X"20",X"4E",X"7E",X"E3",X"C7",X"57",X"67",X"0F",X"37",X"48",X"90",X"20",X"00",X"00",X"00",
		X"0E",X"20",X"4E",X"7E",X"E3",X"C7",X"57",X"67",X"0F",X"17",X"08",X"28",X"24",X"20",X"10",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F1",X"FF",X"7F",X"FF",X"7F",X"7F",X"7F",X"3F",X"3F",X"1F",X"0F",X"0E",X"00",X"00",X"00",X"00",
		X"CF",X"67",X"3F",X"7F",X"3F",X"3F",X"1F",X"1F",X"0F",X"0F",X"0E",X"05",X"01",X"00",X"00",X"00",
		X"38",X"1C",X"3C",X"1C",X"1C",X"1F",X"3F",X"7F",X"7F",X"7F",X"7B",X"31",X"39",X"18",X"00",X"00",
		X"38",X"1C",X"18",X"1F",X"0F",X"4F",X"CF",X"FF",X"FF",X"FF",X"EE",X"C6",X"66",X"64",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",
		X"00",X"00",X"0C",X"0C",X"00",X"0C",X"0E",X"06",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"18",X"18",X"18",X"7F",X"04",X"08",X"00",X"00",X"0F",X"08",X"00",X"08",X"04",X"03",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"00",X"00",X"00",X"F0",X"F8",X"1C",X"0F",X"00",
		X"00",X"00",X"0C",X"0C",X"00",X"0C",X"0E",X"06",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0F",X"00",X"18",X"18",X"18",X"7F",
		X"00",X"18",X"18",X"18",X"7F",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"00",X"00",X"01",X"02",X"04",X"09",X"10",X"01",X"04",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"07",X"78",X"C7",X"00",X"00",X"00",X"00",X"C7",X"FF",X"78",X"00",X"03",
		X"FF",X"FF",X"FF",X"FF",X"F0",X"07",X"F8",X"00",X"00",X"00",X"00",X"F8",X"FF",X"0F",X"00",X"E0",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"00",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"00",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"88",X"6D",X"1D",X"0D",X"3D",X"27",X"73",X"77",X"FA",X"5E",X"4F",X"4F",X"27",X"24",X"18",
		X"04",X"08",X"08",X"0B",X"03",X"02",X"01",X"01",X"01",X"03",X"07",X"06",X"06",X"06",X"06",X"02",
		X"05",X"09",X"08",X"03",X"03",X"03",X"1B",X"33",X"63",X"F1",X"FB",X"5B",X"4A",X"2A",X"20",X"10",
		X"04",X"08",X"08",X"0B",X"03",X"02",X"01",X"01",X"01",X"03",X"07",X"06",X"06",X"06",X"06",X"02",
		X"00",X"03",X"04",X"04",X"0F",X"1A",X"1A",X"0E",X"03",X"01",X"05",X"19",X"37",X"0E",X"3E",X"1C",
		X"00",X"03",X"04",X"04",X"0F",X"1A",X"1A",X"0E",X"13",X"71",X"F5",X"F1",X"E3",X"40",X"00",X"00",
		X"00",X"03",X"04",X"04",X"0F",X"3A",X"9A",X"CE",X"F3",X"71",X"05",X"01",X"03",X"00",X"00",X"00",
		X"07",X"08",X"8F",X"D7",X"79",X"2C",X"03",X"11",X"05",X"01",X"03",X"00",X"00",X"00",X"00",X"00",
		X"41",X"E5",X"F1",X"13",X"0E",X"1A",X"1A",X"0F",X"08",X"04",X"03",X"00",X"00",X"00",X"00",X"00",
		X"41",X"E5",X"F1",X"13",X"0E",X"1A",X"1A",X"0F",X"08",X"04",X"03",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"40",X"40",X"60",X"60",X"30",X"30",X"10",X"10",X"1F",X"0B",X"03",X"03",X"01",X"01",
		X"00",X"00",X"40",X"40",X"60",X"60",X"3F",X"3C",X"1C",X"1C",X"1F",X"0B",X"03",X"03",X"01",X"01",
		X"00",X"00",X"40",X"7F",X"7A",X"7D",X"3F",X"3C",X"1C",X"1C",X"1F",X"0B",X"03",X"03",X"01",X"01",
		X"3F",X"60",X"7F",X"7A",X"7D",X"7F",X"3F",X"3C",X"1C",X"1C",X"1F",X"0B",X"03",X"03",X"01",X"01",
		X"3F",X"60",X"7F",X"7F",X"7A",X"7D",X"3F",X"3C",X"1C",X"1C",X"1F",X"0B",X"03",X"03",X"01",X"01",
		X"00",X"00",X"40",X"40",X"60",X"60",X"30",X"30",X"10",X"10",X"1A",X"0A",X"03",X"03",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"08",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"08",X"00",
		X"00",X"0C",X"0C",X"0C",X"0C",X"4C",X"4C",X"4C",X"4C",X"4C",X"4C",X"4C",X"0C",X"0C",X"0C",X"00",
		X"02",X"06",X"06",X"26",X"26",X"66",X"66",X"66",X"66",X"66",X"66",X"26",X"26",X"06",X"06",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"04",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"04",X"03",X"00",X"00",X"00",
		X"00",X"00",X"02",X"04",X"04",X"08",X"08",X"00",X"00",X"00",X"04",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"02",X"02",X"02",X"00",X"00",X"00",X"02",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"04",X"05",X"05",X"05",X"05",X"05",X"04",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"0F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"07",X"0E",X"0D",X"FF",X"0D",X"0E",X"07",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"0F",X"1C",X"19",X"1B",X"FF",X"1B",X"19",X"1C",X"0F",X"07",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"07",X"07",X"07",X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"00",X"01",X"03",X"23",X"03",X"01",X"00",X"00",X"08",X"00",X"00",X"00",
		X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"05",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"03",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"03",X"01",X"00",X"00",X"01",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"02",X"04",X"04",X"04",X"0C",X"0C",X"0C",X"0C",X"14",
		X"00",X"00",X"00",X"00",X"20",X"22",X"72",X"22",X"24",X"04",X"04",X"0C",X"0C",X"0C",X"0C",X"14",
		X"20",X"20",X"20",X"20",X"20",X"22",X"FA",X"22",X"24",X"24",X"24",X"2C",X"2C",X"2C",X"0C",X"14",
		X"07",X"0F",X"1F",X"1F",X"3F",X"3F",X"7F",X"BF",X"7F",X"3F",X"33",X"73",X"71",X"21",X"00",X"00",
		X"31",X"07",X"3F",X"3F",X"3F",X"7F",X"7F",X"27",X"1F",X"3F",X"38",X"13",X"07",X"07",X"07",X"03",
		X"00",X"00",X"00",X"06",X"0F",X"07",X"03",X"31",X"7B",X"F3",X"FF",X"CF",X"EF",X"66",X"04",X"00",
		X"00",X"03",X"1B",X"1B",X"3D",X"3C",X"14",X"B3",X"FF",X"FF",X"7F",X"37",X"03",X"01",X"01",X"00",
		X"00",X"06",X"01",X"1F",X"1E",X"0F",X"0F",X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"03",
		X"00",X"00",X"06",X"1F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"3F",X"7C",X"9C",X"0E",X"0E",X"04",
		X"07",X"25",X"57",X"57",X"F3",X"E7",X"DF",X"77",X"07",X"1B",X"2C",X"48",X"90",X"00",X"00",X"00",
		X"0C",X"10",X"2C",X"78",X"60",X"3F",X"07",X"1F",X"07",X"2B",X"09",X"00",X"03",X"00",X"00",X"01",
		X"01",X"00",X"00",X"03",X"00",X"08",X"2B",X"07",X"1F",X"07",X"1F",X"23",X"7C",X"70",X"3C",X"10",
		X"00",X"00",X"00",X"10",X"92",X"4A",X"14",X"0F",X"6F",X"DF",X"EF",X"67",X"3F",X"CF",X"6A",X"0E",
		X"00",X"20",X"32",X"6A",X"24",X"A5",X"8F",X"0F",X"3F",X"7F",X"5F",X"77",X"2F",X"0B",X"0E",X"06",
		X"06",X"0F",X"0D",X"37",X"7A",X"6F",X"3F",X"3F",X"0F",X"2F",X"47",X"27",X"EA",X"FA",X"78",X"30",
		X"01",X"05",X"01",X"13",X"4E",X"FA",X"FA",X"CF",X"08",X"04",X"03",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"1F",X"19",X"17",X"03",X"03",X"05",X"04",X"02",X"02",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"02",X"04",X"05",X"03",X"03",X"0F",X"1D",X"19",X"0A",
		X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"04",X"47",X"DD",X"ED",X"7F",X"39",X"00",X"02",X"00",
		X"00",X"30",X"78",X"18",X"4B",X"7C",X"3A",X"17",X"1D",X"2B",X"0E",X"1D",X"27",X"0B",X"00",X"00",
		X"00",X"00",X"0B",X"27",X"1D",X"0E",X"2B",X"1D",X"17",X"3A",X"3C",X"2B",X"2C",X"34",X"18",X"00",
		X"1B",X"09",X"0D",X"05",X"07",X"07",X"02",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"27",X"32",X"12",X"1A",X"1E",X"0A",X"0B",X"0D",X"07",X"07",X"07",X"07",X"05",X"01",X"01",X"01",
		X"12",X"09",X"0D",X"05",X"07",X"07",X"03",X"03",X"03",X"03",X"0A",X"25",X"1F",X"3F",X"1F",X"0E",
		X"32",X"0B",X"05",X"07",X"03",X"03",X"03",X"02",X"40",X"00",X"80",X"C0",X"60",X"7A",X"30",X"00",
		X"0E",X"03",X"81",X"00",X"00",X"02",X"00",X"20",X"30",X"18",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"00",X"00",X"08",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"35",X"53",X"55",X"57",X"60",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"08",X"0E",X"02",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"07",X"0C",X"09",X"09",X"09",X"0C",X"0F",X"08",X"0F",X"0C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"07",X"08",X"08",X"09",X"09",X"09",X"09",X"08",X"0F",X"0C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"07",X"0D",X"0D",X"0D",X"0D",X"0D",X"0D",X"0D",X"07",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"1E",X"3E",X"7E",X"7E",X"FE",X"FE",X"FE",X"FC",X"FC",X"FC",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FE",X"FE",
		X"7F",X"80",X"80",X"00",X"D9",X"FB",X"AA",X"AA",X"AA",X"AA",X"AA",X"A9",X"00",X"80",X"80",X"7F",
		X"00",X"00",X"00",X"7F",X"80",X"80",X"00",X"D9",X"FA",X"AA",X"AA",X"A9",X"00",X"80",X"80",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"80",X"80",X"FB",X"AA",X"AB",X"80",X"80",X"7F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
