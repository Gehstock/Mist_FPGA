library IEEE;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity rom_bas is
	port (
		clk: in std_logic;
		addr: in std_logic_vector(12 downto 0);
		data: out std_logic_vector(7 downto 0)
	);
end entity;

architecture Behavioral of rom_bas is
	type romDef is array(0 to 8191) of std_logic_vector(7 downto 0);
	constant romData: romDef := (
x"4C", x"A3", x"DE", x"4C", x"7F", x"C2", x"FE", x"CE",
x"D1", x"D0", x"5D", x"C6", x"5B", x"C5", x"FF", x"CA",
x"66", x"C7", x"BB", x"C9", x"D9", x"CD", x"EF", x"C9",
x"13", x"C8", x"13", x"C7", x"EB", x"C6", x"96", x"C7",
x"30", x"C6", x"F6", x"C6", x"40", x"C7", x"A9", x"C7",
x"5B", x"C6", x"B9", x"C7", x"02", x"F0", x"6B", x"D5",
x"14", x"F0", x"9E", x"C6", x"F0", x"D0", x"62", x"D5",
x"A8", x"C8", x"84", x"C6", x"BB", x"C4", x"80", x"C4",
x"FF", x"EF", x"64", x"C4", x"78", x"D9", x"0B", x"DA",
x"97", x"D9", x"03", x"00", x"BD", x"D0", x"DE", x"D0",
x"75", x"DC", x"96", x"DD", x"29", x"D7", x"F1", x"DC",
x"D2", x"DD", x"D9", x"DD", x"22", x"DE", x"B1", x"C3",
x"4C", x"D5", x"BA", x"D4", x"A3", x"D1", x"EB", x"D4",
x"C9", x"D4", x"2A", x"D4", x"3E", x"D4", x"6A", x"D4",
x"75", x"D4", x"79", x"A8", x"D5", x"79", x"91", x"D5",
x"7B", x"69", x"D7", x"7B", x"50", x"D8", x"7F", x"7E",
x"DC", x"50", x"41", x"CD", x"46", x"3E", x"CD", x"7D",
x"B7", x"DC", x"5A", x"9B", x"CC", x"64", x"6E", x"CD",
x"45", x"4E", x"C4", x"46", x"4F", x"D2", x"4E", x"45",
x"58", x"D4", x"44", x"41", x"54", x"C1", x"49", x"4E",
x"50", x"55", x"D4", x"44", x"49", x"CD", x"52", x"45",
x"41", x"C4", x"44", x"44", x"D4", x"47", x"4F", x"54",
x"CF", x"52", x"55", x"CE", x"49", x"C6", x"52", x"45",
x"53", x"54", x"4F", x"52", x"C5", x"47", x"4F", x"53",
x"55", x"C2", x"52", x"45", x"54", x"55", x"52", x"CE",
x"52", x"45", x"CD", x"53", x"54", x"4F", x"D0", x"4F",
x"CE", x"44", x"52", x"41", x"D7", x"57", x"41", x"49",
x"D4", x"4C", x"4F", x"41", x"C4", x"53", x"41", x"56",
x"C5", x"44", x"45", x"C6", x"50", x"4F", x"4B", x"C5",
x"50", x"52", x"49", x"4E", x"D4", x"43", x"4F", x"4E",
x"D4", x"4C", x"49", x"53", x"D4", x"43", x"4C", x"45",
x"41", x"D2", x"47", x"45", x"D4", x"4E", x"45", x"D7",
x"54", x"41", x"42", x"A8", x"54", x"CF", x"46", x"CE",
x"53", x"50", x"43", x"A8", x"54", x"48", x"45", x"CE",
x"4E", x"4F", x"D4", x"53", x"54", x"45", x"D0", x"AB",
x"AD", x"AA", x"AF", x"E0", x"41", x"4E", x"C4", x"4F",
x"D2", x"BE", x"BD", x"BC", x"53", x"47", x"CE", x"49",
x"4E", x"D4", x"41", x"42", x"D3", x"55", x"53", x"D2",
x"46", x"52", x"C5", x"50", x"4F", x"D3", x"53", x"51",
x"D2", x"52", x"4E", x"C4", x"4C", x"4F", x"C7", x"45",
x"58", x"D0", x"43", x"4F", x"D3", x"53", x"49", x"CE",
x"54", x"41", x"CE", x"41", x"54", x"CE", x"50", x"45",
x"45", x"CB", x"4C", x"45", x"CE", x"53", x"54", x"52",
x"A4", x"56", x"41", x"CC", x"41", x"53", x"C3", x"43",
x"48", x"52", x"A4", x"4C", x"45", x"46", x"54", x"A4",
x"52", x"49", x"47", x"48", x"54", x"A4", x"4D", x"49",
x"44", x"A4", x"47", x"CF", x"00", x"4E", x"46", x"53",
x"4E", x"52", x"47", x"4F", x"44", x"46", x"43", x"4F",
x"56", x"4F", x"4D", x"55", x"53", x"42", x"53", x"44",
x"44", x"2F", x"30", x"49", x"44", x"54", x"4D", x"4C",
x"53", x"53", x"54", x"43", x"4E", x"55", x"46", x"20",
x"45", x"52", x"52", x"4F", x"52", x"00", x"20", x"49",
x"4E", x"20", x"00", x"0D", x"0A", x"20", x"42", x"52",
x"45", x"41", x"4B", x"00", x"BA", x"E8", x"E8", x"E8",
x"E8", x"BD", x"01", x"01", x"C9", x"81", x"D0", x"21",
x"A5", x"92", x"D0", x"0A", x"BD", x"02", x"01", x"85",
x"91", x"BD", x"03", x"01", x"85", x"92", x"DD", x"03",
x"01", x"D0", x"07", x"A5", x"91", x"DD", x"02", x"01",
x"F0", x"07", x"8A", x"18", x"69", x"12", x"AA", x"D0",
x"D8", x"60", x"20", x"2A", x"C2", x"85", x"79", x"84",
x"7A", x"38", x"A5", x"A2", x"E5", x"A7", x"85", x"6A",
x"A8", x"A5", x"A3", x"E5", x"A8", x"AA", x"E8", x"98",
x"F0", x"23", x"A5", x"A2", x"38", x"E5", x"6A", x"85",
x"A2", x"B0", x"03", x"C6", x"A3", x"38", x"A5", x"A0",
x"E5", x"6A", x"85", x"A0", x"B0", x"08", x"C6", x"A1",
x"90", x"04", x"B1", x"A2", x"91", x"A0", x"88", x"D0",
x"F9", x"B1", x"A2", x"91", x"A0", x"C6", x"A3", x"C6",
x"A1", x"CA", x"D0", x"F2", x"60", x"0A", x"69", x"44",
x"B0", x"35", x"85", x"6A", x"BA", x"E4", x"6A", x"90",
x"2E", x"60", x"C4", x"7C", x"90", x"28", x"D0", x"04",
x"C5", x"7B", x"90", x"22", x"48", x"A2", x"09", x"98",
x"48", x"B5", x"9F", x"CA", x"10", x"FA", x"20", x"64",
x"D2", x"A2", x"F7", x"68", x"95", x"A9", x"E8", x"30",
x"FA", x"68", x"A8", x"68", x"C4", x"7C", x"90", x"06",
x"D0", x"05", x"C5", x"7B", x"B0", x"01", x"60", x"A2",
x"0C", x"46", x"10", x"20", x"00", x"C9", x"20", x"6A",
x"C9", x"BD", x"75", x"C1", x"20", x"6C", x"C9", x"BD",
x"76", x"C1", x"20", x"6C", x"C9", x"20", x"9A", x"C4",
x"A9", x"97", x"A0", x"C1", x"20", x"4A", x"C9", x"A4",
x"82", x"C8", x"F0", x"03", x"20", x"1E", x"F0", x"46",
x"10", x"20", x"00", x"00", x"20", x"65", x"C3", x"86",
x"C6", x"84", x"C7", x"20", x"BF", x"00", x"AA", x"F0",
x"F3", x"A2", x"FF", x"86", x"82", x"90", x"06", x"20",
x"AE", x"C3", x"4C", x"F8", x"C5", x"20", x"DA", x"C7",
x"20", x"AE", x"C3", x"84", x"08", x"20", x"36", x"C4",
x"90", x"44", x"A0", x"01", x"B1", x"A7", x"85", x"6B",
x"A5", x"75", x"85", x"6A", x"A5", x"A8", x"85", x"6D",
x"A5", x"A7", x"88", x"F1", x"A7", x"18", x"65", x"75",
x"85", x"75", x"85", x"6C", x"A5", x"76", x"69", x"FF",
x"85", x"76", x"E5", x"A8", x"AA", x"38", x"A5", x"A7",
x"E5", x"75", x"A8", x"B0", x"03", x"E8", x"C6", x"6D",
x"18", x"65", x"6A", x"90", x"03", x"C6", x"6B", x"18",
x"B1", x"6A", x"91", x"6C", x"C8", x"D0", x"F9", x"E6",
x"6B", x"E6", x"6D", x"CA", x"D0", x"F2", x"20", x"7C",
x"C4", x"20", x"29", x"C3", x"A5", x"16", x"F0", x"8C",
x"18", x"A5", x"75", x"85", x"A2", x"65", x"08", x"85",
x"A0", x"A4", x"76", x"84", x"A3", x"90", x"01", x"C8",
x"84", x"A1", x"20", x"DA", x"C1", x"A5", x"79", x"A4",
x"7A", x"85", x"75", x"84", x"76", x"A4", x"08", x"88",
x"B9", x"12", x"00", x"91", x"A7", x"88", x"10", x"F8",
x"20", x"7C", x"C4", x"20", x"29", x"C3", x"4C", x"84",
x"C2", x"A5", x"73", x"A4", x"74", x"85", x"6A", x"84",
x"6B", x"18", x"A0", x"01", x"B1", x"6A", x"F0", x"1D",
x"A0", x"04", x"C8", x"B1", x"6A", x"D0", x"FB", x"C8",
x"98", x"65", x"6A", x"AA", x"A0", x"00", x"91", x"6A",
x"A5", x"6B", x"69", x"00", x"C8", x"91", x"6A", x"86",
x"6A", x"85", x"6B", x"90", x"DD", x"60", x"CA", x"30",
x"09", x"EA", x"EA", x"EA", x"4C", x"67", x"C3", x"20",
x"6C", x"C9", x"20", x"00", x"C9", x"A2", x"00", x"20",
x"9E", x"C3", x"C9", x"1A", x"D0", x"06", x"20", x"18",
x"F0", x"4C", x"65", x"C3", x"C9", x"03", x"F0", x"14",
x"C9", x"0D", x"F0", x"1F", x"C9", x"08", x"F0", x"D6",
x"C9", x"18", x"F0", x"DB", x"C9", x"20", x"90", x"0E",
x"C9", x"80", x"B0", x"DB", x"E0", x"47", x"B0", x"04",
x"95", x"16", x"E8", x"2C", x"A9", x"07", x"20", x"2A",
x"F0", x"D0", x"CC", x"4C", x"FA", x"C8", x"20", x"AB",
x"C6", x"C9", x"0F", x"D0", x"08", x"48", x"A5", x"10",
x"49", x"FF", x"85", x"10", x"68", x"60", x"4C", x"36",
x"F0", x"A5", x"AE", x"48", x"10", x"03", x"20", x"E1",
x"C3", x"A5", x"A9", x"48", x"C9", x"81", x"90", x"07",
x"A9", x"FB", x"A0", x"D6", x"20", x"4E", x"D8", x"A9",
x"EC", x"A0", x"C3", x"20", x"5A", x"DD", x"68", x"C9",
x"81", x"90", x"07", x"A9", x"4E", x"A0", x"DE", x"20",
x"8F", x"D5", x"68", x"10", x"03", x"4C", x"E1", x"C3",
x"60", x"A5", x"A9", x"F0", x"06", x"A5", x"AE", x"49",
x"FF", x"85", x"AE", x"60", x"0C", x"76", x"B3", x"83",
x"BD", x"D3", x"79", x"1E", x"F4", x"A6", x"F5", x"7B",
x"83", x"FC", x"B0", x"10", x"7C", x"0C", x"1F", x"67",
x"CA", x"7C", x"DE", x"53", x"CB", x"C1", x"7D", x"14",
x"64", x"70", x"4C", x"7D", x"B7", x"EA", x"51", x"7A",
x"7D", x"63", x"30", x"88", x"7E", x"7E", x"92", x"44",
x"99", x"3A", x"7E", x"4C", x"CC", x"91", x"C7", x"7F",
x"AA", x"AA", x"AA", x"13", x"81", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"A5", x"73",
x"A6", x"74", x"A0", x"01", x"85", x"A7", x"86", x"A8",
x"B1", x"A7", x"F0", x"1F", x"C8", x"C8", x"A5", x"15",
x"D1", x"A7", x"90", x"18", x"F0", x"03", x"88", x"D0",
x"09", x"A5", x"14", x"88", x"D1", x"A7", x"90", x"0C",
x"F0", x"0A", x"88", x"B1", x"A7", x"AA", x"88", x"B1",
x"A7", x"B0", x"D7", x"18", x"60", x"D0", x"FD", x"A9",
x"00", x"A8", x"91", x"73", x"C8", x"91", x"73", x"A5",
x"73", x"18", x"69", x"02", x"85", x"75", x"A5", x"74",
x"69", x"00", x"85", x"76", x"20", x"AE", x"C4", x"A9",
x"00", x"D0", x"2A", x"A5", x"7F", x"A4", x"80", x"85",
x"7B", x"84", x"7C", x"A5", x"75", x"A4", x"76", x"85",
x"77", x"84", x"78", x"85", x"79", x"84", x"7A", x"20",
x"31", x"C6", x"A2", x"61", x"86", x"5E", x"68", x"A8",
x"68", x"A2", x"FD", x"9A", x"48", x"98", x"48", x"A9",
x"00", x"85", x"86", x"85", x"0D", x"60", x"18", x"A5",
x"73", x"69", x"FF", x"85", x"C6", x"A5", x"74", x"69",
x"FF", x"85", x"C7", x"60", x"48", x"A9", x"00", x"85",
x"0E", x"68", x"08", x"20", x"DA", x"C7", x"20", x"36",
x"C4", x"28", x"F0", x"14", x"20", x"C5", x"00", x"F0",
x"15", x"C9", x"A5", x"D0", x"8F", x"20", x"BF", x"00",
x"F0", x"06", x"20", x"DA", x"C7", x"F0", x"07", x"60",
x"A9", x"FF", x"85", x"14", x"85", x"15", x"68", x"68",
x"A0", x"01", x"B1", x"A7", x"F0", x"39", x"20", x"40",
x"C6", x"20", x"00", x"C9", x"C8", x"B1", x"A7", x"AA",
x"C8", x"B1", x"A7", x"C5", x"15", x"D0", x"04", x"E4",
x"14", x"F0", x"02", x"B0", x"22", x"84", x"91", x"20",
x"0C", x"DB", x"A9", x"20", x"A4", x"91", x"29", x"7F",
x"20", x"6C", x"C9", x"C8", x"F0", x"11", x"B1", x"A7",
x"D0", x"22", x"A8", x"B1", x"A7", x"AA", x"C8", x"B1",
x"A7", x"86", x"A7", x"85", x"A8", x"D0", x"C1", x"A5",
x"0E", x"F0", x"0E", x"20", x"00", x"C9", x"20", x"00",
x"C9", x"A9", x"1A", x"20", x"6C", x"C9", x"20", x"1B",
x"F0", x"4C", x"7F", x"C2", x"10", x"D2", x"4C", x"39",
x"F0", x"AA", x"84", x"91", x"A0", x"FF", x"CA", x"F0",
x"08", x"C8", x"B9", x"90", x"C0", x"10", x"FA", x"30",
x"F5", x"C8", x"B9", x"90", x"C0", x"30", x"B5", x"20",
x"6C", x"C9", x"D0", x"F5", x"A9", x"80", x"85", x"0D",
x"20", x"14", x"C8", x"20", x"AC", x"C1", x"D0", x"05",
x"8A", x"69", x"0F", x"AA", x"9A", x"68", x"68", x"A9",
x"09", x"20", x"1D", x"C2", x"20", x"75", x"C7", x"18",
x"98", x"65", x"C6", x"48", x"A5", x"C7", x"69", x"00",
x"48", x"A5", x"82", x"48", x"A5", x"81", x"48", x"A9",
x"9E", x"20", x"C7", x"CC", x"20", x"6E", x"CB", x"20",
x"6B", x"CB", x"A5", x"AE", x"09", x"7F", x"25", x"AA",
x"85", x"AA", x"A9", x"A5", x"A0", x"C5", x"85", x"6A",
x"84", x"6B", x"4C", x"24", x"CC", x"A9", x"FB", x"A0",
x"D6", x"20", x"E1", x"D8", x"20", x"C5", x"00", x"C9",
x"A3", x"D0", x"06", x"20", x"BF", x"00", x"20", x"6B",
x"CB", x"20", x"6A", x"D9", x"20", x"19", x"CC", x"A5",
x"92", x"48", x"A5", x"91", x"48", x"A9", x"81", x"48",
x"20", x"40", x"C6", x"A5", x"C6", x"A4", x"C7", x"F0",
x"06", x"85", x"85", x"84", x"86", x"A0", x"00", x"B1",
x"C6", x"D0", x"40", x"A0", x"02", x"B1", x"C6", x"18",
x"D0", x"03", x"4C", x"75", x"C6", x"C8", x"B1", x"C6",
x"85", x"81", x"C8", x"B1", x"C6", x"85", x"82", x"98",
x"65", x"C6", x"85", x"C6", x"90", x"02", x"E6", x"C7",
x"20", x"BF", x"00", x"20", x"01", x"C6", x"4C", x"C8",
x"C5", x"4C", x"33", x"F0", x"EA", x"90", x"11", x"C9",
x"1D", x"B0", x"17", x"0A", x"A8", x"B9", x"0B", x"C0",
x"48", x"B9", x"0A", x"C0", x"48", x"4C", x"BF", x"00",
x"4C", x"14", x"C8", x"C9", x"3A", x"F0", x"D9", x"4C",
x"D0", x"CC", x"C9", x"45", x"D0", x"F9", x"20", x"BF",
x"00", x"A9", x"9E", x"20", x"C7", x"CC", x"4C", x"14",
x"C7", x"38", x"A5", x"73", x"E9", x"01", x"A4", x"74",
x"B0", x"01", x"88", x"85", x"89", x"84", x"8A", x"60",
x"AD", x"FD", x"87", x"29", x"30", x"C9", x"10", x"38",
x"D0", x"F5", x"AD", x"7F", x"87", x"29", x"30", x"C9",
x"10", x"38", x"D0", x"EB", x"20", x"30", x"F0", x"EA",
x"A9", x"03", x"C9", x"03", x"B0", x"01", x"18", x"D0",
x"3D", x"A5", x"C6", x"A4", x"C7", x"F0", x"0C", x"85",
x"85", x"84", x"86", x"A5", x"81", x"A4", x"82", x"85",
x"83", x"84", x"84", x"68", x"68", x"A9", x"A3", x"A0",
x"C1", x"A2", x"00", x"86", x"10", x"90", x"03", x"4C",
x"74", x"C2", x"4C", x"7F", x"C2", x"D0", x"17", x"A2",
x"1E", x"A4", x"86", x"D0", x"03", x"4C", x"59", x"C2",
x"A5", x"85", x"85", x"C6", x"84", x"C7", x"A5", x"83",
x"A4", x"84", x"85", x"81", x"84", x"82", x"60", x"48",
x"20", x"12", x"F0", x"20", x"67", x"C9", x"A9", x"FF",
x"4C", x"BF", x"C4", x"AD", x"40", x"02", x"20", x"D8",
x"C6", x"D0", x"03", x"4C", x"0F", x"F0", x"4C", x"24",
x"F0", x"48", x"AD", x"41", x"02", x"20", x"D8", x"C6",
x"D0", x"04", x"68", x"4C", x"0C", x"F0", x"68", x"C9",
x"0A", x"EA", x"EA", x"C9", x"0D", x"F0", x"03", x"4C",
x"27", x"F0", x"20", x"27", x"F0", x"A9", x"0D", x"60",
x"C9", x"54", x"F0", x"06", x"C9", x"44", x"F0", x"02",
x"C9", x"FF", x"60", x"20", x"B0", x"E5", x"EA", x"90",
x"EF", x"EA", x"EA", x"60", x"D0", x"03", x"4C", x"7C",
x"C4", x"20", x"83", x"C4", x"4C", x"0B", x"C7", x"A9",
x"03", x"20", x"1D", x"C2", x"A5", x"C7", x"48", x"A5",
x"C6", x"48", x"A5", x"82", x"48", x"A5", x"81", x"48",
x"A9", x"8C", x"48", x"20", x"C5", x"00", x"20", x"14",
x"C7", x"4C", x"C8", x"C5", x"20", x"DA", x"C7", x"20",
x"78", x"C7", x"A5", x"82", x"C5", x"15", x"B0", x"0B",
x"98", x"38", x"65", x"C6", x"A6", x"C7", x"90", x"07",
x"E8", x"B0", x"04", x"A5", x"73", x"A6", x"74", x"20",
x"3A", x"C4", x"90", x"1E", x"A5", x"A7", x"E9", x"01",
x"85", x"C6", x"A5", x"A8", x"E9", x"00", x"85", x"C7",
x"60", x"D0", x"FD", x"A9", x"FF", x"85", x"92", x"20",
x"AC", x"C1", x"9A", x"C9", x"8C", x"F0", x"0B", x"A2",
x"04", x"2C", x"A2", x"0E", x"4C", x"59", x"C2", x"4C",
x"D0", x"CC", x"68", x"68", x"85", x"81", x"68", x"85",
x"82", x"68", x"85", x"C6", x"68", x"85", x"C7", x"20",
x"75", x"C7", x"98", x"18", x"65", x"C6", x"85", x"C6",
x"90", x"02", x"E6", x"C7", x"60", x"A2", x"3A", x"2C",
x"A2", x"00", x"86", x"06", x"A0", x"00", x"84", x"07",
x"A5", x"07", x"A6", x"06", x"85", x"06", x"86", x"07",
x"B1", x"C6", x"F0", x"E8", x"C5", x"07", x"F0", x"E4",
x"C8", x"C9", x"22", x"D0", x"F3", x"F0", x"E9", x"20",
x"7F", x"CB", x"20", x"C5", x"00", x"C9", x"88", x"F0",
x"05", x"A9", x"A1", x"20", x"C7", x"CC", x"A5", x"A9",
x"D0", x"05", x"20", x"78", x"C7", x"F0", x"BB", x"20",
x"C5", x"00", x"B0", x"03", x"4C", x"14", x"C7", x"4C",
x"01", x"C6", x"20", x"DC", x"D4", x"48", x"C9", x"8C",
x"F0", x"04", x"C9", x"88", x"D0", x"91", x"C6", x"AD",
x"D0", x"04", x"68", x"4C", x"21", x"F0", x"20", x"BF",
x"00", x"20", x"DA", x"C7", x"C9", x"2C", x"F0", x"EE",
x"68", x"60", x"A2", x"00", x"86", x"14", x"86", x"15",
x"B0", x"F7", x"E9", x"2F", x"85", x"06", x"A5", x"15",
x"85", x"6A", x"C9", x"19", x"B0", x"D4", x"A5", x"14",
x"0A", x"26", x"6A", x"0A", x"26", x"6A", x"65", x"14",
x"85", x"14", x"A5", x"6A", x"65", x"15", x"85", x"15",
x"06", x"14", x"26", x"15", x"A5", x"14", x"65", x"06",
x"85", x"14", x"90", x"02", x"E6", x"15", x"20", x"BF",
x"00", x"4C", x"E0", x"C7", x"20", x"E4", x"CD", x"85",
x"91", x"84", x"92", x"A9", x"AC", x"20", x"C7", x"CC",
x"A5", x"0B", x"48", x"A5", x"0A", x"48", x"20", x"4B",
x"F0", x"68", x"2A", x"20", x"71", x"CB", x"D0", x"18",
x"68", x"10", x"12", x"20", x"5A", x"D9", x"20", x"FE",
x"CE", x"A0", x"00", x"A5", x"AC", x"91", x"91", x"C8",
x"A5", x"AD", x"91", x"91", x"60", x"4C", x"0F", x"D9",
x"68", x"A0", x"02", x"B1", x"AC", x"C5", x"7C", x"90",
x"17", x"D0", x"07", x"88", x"B1", x"AC", x"C5", x"7B",
x"90", x"0E", x"A4", x"AD", x"C4", x"76", x"90", x"08",
x"D0", x"0D", x"A5", x"AC", x"C5", x"75", x"B0", x"07",
x"A5", x"AC", x"A4", x"AD", x"4C", x"85", x"C8", x"A0",
x"00", x"B1", x"AC", x"20", x"B3", x"D1", x"A5", x"98",
x"A4", x"99", x"85", x"B7", x"84", x"B8", x"20", x"B8",
x"D3", x"A9", x"A9", x"A0", x"00", x"85", x"98", x"84",
x"99", x"20", x"19", x"D4", x"A0", x"00", x"B1", x"98",
x"91", x"91", x"C8", x"B1", x"98", x"91", x"91", x"C8",
x"B1", x"98", x"91", x"91", x"60", x"C9", x"21", x"D0",
x"FB", x"A9", x"FF", x"8D", x"10", x"02", x"4C", x"BF",
x"00", x"AD", x"10", x"02", x"85", x"BE", x"20", x"BA",
x"C8", x"A5", x"BE", x"8D", x"10", x"02", x"60", x"20",
x"4D", x"C9", x"20", x"C5", x"00", x"F0", x"41", x"F0",
x"51", x"20", x"9D", x"C8", x"F0", x"4C", x"C9", x"9D",
x"F0", x"60", x"C9", x"A0", x"18", x"F0", x"5B", x"C9",
x"2C", x"F0", x"40", x"C9", x"3B", x"F0", x"68", x"20",
x"7F", x"CB", x"24", x"0A", x"30", x"D9", x"20", x"1C",
x"DB", x"20", x"C5", x"D1", x"A0", x"00", x"B1", x"AC",
x"18", x"65", x"11", x"C5", x"12", x"90", x"03", x"20",
x"00", x"C9", x"20", x"4D", x"C9", x"20", x"67", x"C9",
x"D0", x"C0", x"A0", x"00", x"94", x"16", x"A2", x"15",
x"A9", x"0D", x"85", x"11", x"20", x"6C", x"C9", x"A9",
x"0A", x"20", x"6C", x"C9", x"A9", x"00", x"85", x"11",
x"49", x"FF", x"60", x"A5", x"11", x"C5", x"13", x"90",
x"06", x"20", x"00", x"C9", x"4C", x"3F", x"C9", x"38",
x"E9", x"0A", x"B0", x"FC", x"49", x"FF", x"69", x"01",
x"D0", x"10", x"08", x"20", x"D9", x"D4", x"C9", x"29",
x"D0", x"68", x"28", x"90", x"06", x"8A", x"E5", x"11",
x"90", x"05", x"AA", x"E8", x"CA", x"D0", x"06", x"20",
x"BF", x"00", x"4C", x"BF", x"C8", x"20", x"67", x"C9",
x"D0", x"F2", x"20", x"C5", x"D1", x"20", x"E4", x"D3",
x"AA", x"A0", x"00", x"E8", x"CA", x"F0", x"BB", x"B1",
x"6A", x"20", x"6C", x"C9", x"C8", x"C9", x"0D", x"D0",
x"F3", x"20", x"0C", x"C9", x"4C", x"54", x"C9", x"A9",
x"20", x"2C", x"A9", x"3F", x"24", x"10", x"30", x"15",
x"48", x"C9", x"20", x"90", x"0C", x"A5", x"11", x"C5",
x"12", x"D0", x"04", x"A9", x"00", x"85", x"11", x"E6",
x"11", x"68", x"20", x"B9", x"C6", x"29", x"FF", x"60",
x"A5", x"0E", x"F0", x"11", x"30", x"04", x"A0", x"FF",
x"D0", x"04", x"A5", x"87", x"A4", x"88", x"85", x"81",
x"84", x"82", x"4C", x"D0", x"CC", x"A9", x"ED", x"A0",
x"CA", x"20", x"4A", x"C9", x"A5", x"85", x"A4", x"86",
x"85", x"C6", x"84", x"C7", x"60", x"20", x"E4", x"D0",
x"A2", x"17", x"A0", x"00", x"84", x"17", x"A9", x"40",
x"20", x"F6", x"C9", x"60", x"46", x"10", x"AD", x"10",
x"02", x"85", x"BE", x"20", x"FA", x"DF", x"C9", x"22",
x"D0", x"0B", x"20", x"85", x"CC", x"A9", x"3B", x"20",
x"C7", x"CC", x"20", x"4D", x"C9", x"20", x"E4", x"D0",
x"A9", x"2C", x"85", x"15", x"20", x"E7", x"C9", x"A5",
x"16", x"20", x"5D", x"DF", x"4C", x"F5", x"C9", x"20",
x"6A", x"C9", x"20", x"67", x"C9", x"4C", x"65", x"C3",
x"A6", x"89", x"A4", x"8A", x"A9", x"98", x"85", x"0E",
x"86", x"8B", x"84", x"8C", x"20", x"E4", x"CD", x"85",
x"91", x"84", x"92", x"A5", x"C6", x"A4", x"C7", x"85",
x"93", x"84", x"94", x"A6", x"8B", x"A4", x"8C", x"86",
x"C6", x"84", x"C7", x"20", x"C5", x"00", x"D0", x"1B",
x"24", x"0E", x"50", x"0B", x"20", x"E3", x"C6", x"85",
x"16", x"A2", x"15", x"A0", x"00", x"F0", x"08", x"30",
x"71", x"20", x"6A", x"C9", x"20", x"E7", x"C9", x"86",
x"C6", x"84", x"C7", x"20", x"BF", x"00", x"24", x"0A",
x"10", x"31", x"24", x"0E", x"50", x"09", x"E8", x"86",
x"C6", x"A9", x"00", x"85", x"06", x"F0", x"0C", x"85",
x"06", x"C9", x"22", x"F0", x"07", x"A9", x"3A", x"85",
x"06", x"A9", x"2C", x"18", x"85", x"07", x"A5", x"C6",
x"A4", x"C7", x"69", x"00", x"90", x"01", x"C8", x"20",
x"CB", x"D1", x"20", x"21", x"D5", x"20", x"49", x"C8",
x"4C", x"73", x"CA", x"20", x"32", x"DA", x"A5", x"0B",
x"20", x"31", x"C8", x"20", x"C5", x"00", x"F0", x"07",
x"C9", x"2C", x"F0", x"03", x"4C", x"88", x"C9", x"A5",
x"C6", x"A4", x"C7", x"85", x"8B", x"84", x"8C", x"A5",
x"93", x"A4", x"94", x"85", x"C6", x"84", x"C7", x"20",
x"C5", x"00", x"F0", x"2C", x"20", x"C5", x"CC", x"4C",
x"FC", x"C9", x"20", x"75", x"C7", x"C8", x"AA", x"D0",
x"12", x"A2", x"06", x"C8", x"B1", x"C6", x"F0", x"6C",
x"C8", x"B1", x"C6", x"85", x"87", x"C8", x"B1", x"C6",
x"C8", x"85", x"88", x"B1", x"C6", x"AA", x"20", x"6A",
x"C7", x"E0", x"83", x"D0", x"DD", x"4C", x"33", x"CA",
x"A5", x"8B", x"A4", x"8C", x"A6", x"0E", x"10", x"03",
x"4C", x"3B", x"C6", x"A0", x"00", x"20", x"B1", x"C8",
x"B1", x"8B", x"F0", x"07", x"A9", x"DC", x"A0", x"CA",
x"4C", x"4A", x"C9", x"60", x"3F", x"45", x"58", x"54",
x"52", x"41", x"20", x"49", x"47", x"4E", x"4F", x"52",
x"45", x"44", x"0D", x"0A", x"00", x"3F", x"52", x"45",
x"44", x"4F", x"20", x"46", x"52", x"4F", x"4D", x"20",
x"53", x"54", x"41", x"52", x"54", x"0D", x"0A", x"00",
x"D0", x"04", x"A0", x"00", x"F0", x"03", x"20", x"E4",
x"CD", x"85", x"91", x"84", x"92", x"20", x"AC", x"C1",
x"F0", x"04", x"A2", x"00", x"F0", x"66", x"9A", x"8A",
x"18", x"69", x"04", x"48", x"69", x"06", x"85", x"6C",
x"68", x"A0", x"01", x"20", x"E1", x"D8", x"BA", x"BD",
x"09", x"01", x"85", x"AE", x"A5", x"91", x"A4", x"92",
x"20", x"A6", x"D5", x"20", x"0F", x"D9", x"A0", x"01",
x"20", x"9C", x"D9", x"BA", x"38", x"FD", x"09", x"01",
x"F0", x"17", x"BD", x"0F", x"01", x"85", x"81", x"BD",
x"10", x"01", x"85", x"82", x"BD", x"12", x"01", x"85",
x"C6", x"BD", x"11", x"01", x"85", x"C7", x"4C", x"C8",
x"C5", x"8A", x"69", x"11", x"AA", x"9A", x"20", x"C5",
x"00", x"C9", x"2C", x"D0", x"F1", x"20", x"BF", x"00",
x"20", x"06", x"CB", x"20", x"7F", x"CB", x"18", x"24",
x"38", x"24", x"0A", x"30", x"03", x"B0", x"03", x"60",
x"B0", x"FD", x"A2", x"18", x"4C", x"59", x"C2", x"A6",
x"C6", x"D0", x"02", x"C6", x"C7", x"C6", x"C6", x"A2",
x"00", x"24", x"48", x"8A", x"48", x"A9", x"01", x"20",
x"1D", x"C2", x"20", x"64", x"CC", x"A9", x"00", x"85",
x"95", x"20", x"C5", x"00", x"38", x"E9", x"AB", x"90",
x"17", x"C9", x"03", x"B0", x"13", x"C9", x"01", x"2A",
x"49", x"01", x"45", x"95", x"C5", x"95", x"90", x"61",
x"85", x"95", x"20", x"BF", x"00", x"4C", x"9C", x"CB",
x"A6", x"95", x"D0", x"2C", x"B0", x"7B", x"69", x"07",
x"90", x"77", x"65", x"0A", x"D0", x"03", x"4C", x"7B",
x"D3", x"69", x"FF", x"85", x"6A", x"0A", x"65", x"6A",
x"A8", x"68", x"D9", x"72", x"C0", x"B0", x"67", x"20",
x"6E", x"CB", x"48", x"20", x"01", x"CC", x"68", x"A4",
x"93", x"10", x"17", x"AA", x"F0", x"56", x"D0", x"5F",
x"46", x"0A", x"8A", x"2A", x"A6", x"C6", x"D0", x"02",
x"C6", x"C7", x"C6", x"C6", x"A0", x"1B", x"85", x"95",
x"D0", x"D7", x"D9", x"72", x"C0", x"B0", x"48", x"90",
x"D9", x"B9", x"74", x"C0", x"48", x"B9", x"73", x"C0",
x"48", x"20", x"14", x"CC", x"A5", x"95", x"4C", x"8A",
x"CB", x"4C", x"D0", x"CC", x"A5", x"AE", x"BE", x"72",
x"C0", x"A8", x"68", x"85", x"6A", x"E6", x"6A", x"68",
x"85", x"6B", x"98", x"48", x"20", x"5A", x"D9", x"A5",
x"AD", x"48", x"A5", x"AC", x"48", x"A5", x"AB", x"48",
x"A5", x"AA", x"48", x"A5", x"A9", x"48", x"6C", x"6A",
x"00", x"A0", x"FF", x"68", x"F0", x"23", x"C9", x"64",
x"F0", x"03", x"20", x"6E", x"CB", x"84", x"93", x"68",
x"4A", x"85", x"0F", x"68", x"85", x"B1", x"68", x"85",
x"B2", x"68", x"85", x"B3", x"68", x"85", x"B4", x"68",
x"85", x"B5", x"68", x"85", x"B6", x"45", x"AE", x"85",
x"B7", x"A5", x"A9", x"60", x"A9", x"00", x"85", x"0A",
x"20", x"BF", x"00", x"B0", x"03", x"4C", x"32", x"DA",
x"20", x"6E", x"CE", x"B0", x"67", x"C9", x"2E", x"F0",
x"F4", x"C9", x"A5", x"F0", x"58", x"C9", x"A4", x"F0",
x"E7", x"C9", x"22", x"D0", x"0F", x"A5", x"C6", x"A4",
x"C7", x"69", x"00", x"90", x"01", x"C8", x"20", x"C5",
x"D1", x"4C", x"21", x"D5", x"C9", x"A2", x"D0", x"13",
x"A0", x"18", x"D0", x"3B", x"20", x"FE", x"CE", x"A5",
x"AD", x"49", x"FF", x"A8", x"A5", x"AC", x"49", x"FF",
x"4C", x"D1", x"D0", x"C9", x"9F", x"D0", x"03", x"4C",
x"32", x"D1", x"C9", x"AE", x"90", x"03", x"4C", x"00",
x"CD", x"20", x"C2", x"CC", x"20", x"7F", x"CB", x"A9",
x"29", x"2C", x"A9", x"28", x"2C", x"A9", x"2C", x"A0",
x"00", x"D1", x"C6", x"D0", x"03", x"4C", x"BF", x"00",
x"A2", x"02", x"4C", x"59", x"C2", x"A0", x"15", x"68",
x"68", x"4C", x"DB", x"CB", x"20", x"E4", x"CD", x"85",
x"AC", x"84", x"AD", x"A6", x"0A", x"F0", x"05", x"A2",
x"00", x"86", x"B8", x"60", x"A6", x"0B", x"10", x"0D",
x"A0", x"00", x"B1", x"AC", x"AA", x"C8", x"B1", x"AC",
x"A8", x"8A", x"4C", x"D1", x"D0", x"4C", x"E1", x"D8",
x"0A", x"48", x"AA", x"20", x"BF", x"00", x"E0", x"83",
x"90", x"20", x"20", x"C2", x"CC", x"20", x"7F", x"CB",
x"20", x"C5", x"CC", x"20", x"70", x"CB", x"68", x"AA",
x"A5", x"AD", x"48", x"A5", x"AC", x"48", x"8A", x"48",
x"20", x"DC", x"D4", x"68", x"A8", x"8A", x"48", x"4C",
x"2F", x"CD", x"20", x"B9", x"CC", x"68", x"A8", x"B9",
x"E8", x"BF", x"85", x"9D", x"B9", x"E9", x"BF", x"85",
x"9E", x"20", x"9C", x"00", x"4C", x"6E", x"CB", x"A0",
x"FF", x"2C", x"A0", x"00", x"84", x"08", x"20", x"FE",
x"CE", x"A5", x"AC", x"45", x"08", x"85", x"06", x"A5",
x"AD", x"45", x"08", x"85", x"07", x"20", x"3B", x"D9",
x"20", x"FE", x"CE", x"A5", x"AD", x"45", x"08", x"25",
x"07", x"45", x"08", x"A8", x"A5", x"AC", x"45", x"08",
x"25", x"06", x"45", x"08", x"4C", x"D1", x"D0", x"20",
x"71", x"CB", x"B0", x"13", x"A5", x"B6", x"09", x"7F",
x"25", x"B2", x"85", x"B2", x"A9", x"B1", x"A0", x"00",
x"20", x"9A", x"D9", x"AA", x"4C", x"BA", x"CD", x"A9",
x"00", x"85", x"0A", x"C6", x"95", x"20", x"E4", x"D3",
x"85", x"A9", x"86", x"AA", x"84", x"AB", x"A5", x"B4",
x"A4", x"B5", x"20", x"E8", x"D3", x"86", x"B4", x"84",
x"B5", x"AA", x"38", x"E5", x"A9", x"F0", x"08", x"A9",
x"01", x"90", x"04", x"A6", x"A9", x"A9", x"FF", x"85",
x"AE", x"A0", x"FF", x"E8", x"C8", x"CA", x"D0", x"07",
x"A6", x"AE", x"30", x"0F", x"18", x"90", x"0C", x"B1",
x"B4", x"D1", x"AA", x"F0", x"EF", x"A2", x"FF", x"B0",
x"02", x"A2", x"01", x"E8", x"8A", x"2A", x"25", x"0F",
x"F0", x"02", x"A9", x"FF", x"4C", x"7B", x"D9", x"20",
x"C5", x"CC", x"AA", x"20", x"E9", x"CD", x"20", x"C5",
x"00", x"D0", x"F4", x"60", x"A2", x"00", x"20", x"C5",
x"00", x"86", x"09", x"85", x"8D", x"20", x"C5", x"00",
x"20", x"6E", x"CE", x"B0", x"03", x"4C", x"D0", x"CC",
x"A2", x"00", x"86", x"0A", x"86", x"0B", x"20", x"BF",
x"00", x"90", x"05", x"20", x"6E", x"CE", x"90", x"0B",
x"AA", x"20", x"BF", x"00", x"90", x"FB", x"20", x"6E",
x"CE", x"B0", x"F6", x"C9", x"24", x"D0", x"06", x"A9",
x"FF", x"85", x"0A", x"D0", x"10", x"C9", x"25", x"D0",
x"13", x"A5", x"0D", x"D0", x"D0", x"A9", x"80", x"85",
x"0B", x"05", x"8D", x"85", x"8D", x"8A", x"09", x"80",
x"AA", x"20", x"BF", x"00", x"86", x"8E", x"38", x"05",
x"0D", x"E9", x"28", x"D0", x"03", x"4C", x"10", x"CF",
x"A9", x"00", x"85", x"0D", x"A5", x"75", x"A6", x"76",
x"A0", x"00", x"86", x"A8", x"85", x"A7", x"E4", x"78",
x"D0", x"04", x"C5", x"77", x"F0", x"22", x"A5", x"8D",
x"D1", x"A7", x"D0", x"08", x"A5", x"8E", x"C8", x"D1",
x"A7", x"F0", x"6A", x"88", x"18", x"A5", x"A7", x"69",
x"07", x"90", x"E1", x"E8", x"D0", x"DC", x"C9", x"41",
x"90", x"05", x"4C", x"3C", x"F0", x"EA", x"EA", x"60",
x"68", x"48", x"C9", x"DE", x"D0", x"0D", x"BA", x"BD",
x"02", x"01", x"C9", x"CC", x"D0", x"05", x"A9", x"4E",
x"A0", x"DC", x"60", x"A5", x"77", x"A4", x"78", x"85",
x"A7", x"84", x"A8", x"A5", x"79", x"A4", x"7A", x"85",
x"A2", x"84", x"A3", x"18", x"69", x"07", x"90", x"01",
x"C8", x"85", x"A0", x"84", x"A1", x"20", x"DA", x"C1",
x"A5", x"A0", x"A4", x"A1", x"C8", x"85", x"77", x"84",
x"78", x"A0", x"00", x"A5", x"8D", x"91", x"A7", x"C8",
x"A5", x"8E", x"91", x"A7", x"A9", x"00", x"C8", x"91",
x"A7", x"C8", x"91", x"A7", x"C8", x"91", x"A7", x"C8",
x"91", x"A7", x"C8", x"91", x"A7", x"A5", x"A7", x"18",
x"69", x"02", x"A4", x"A8", x"90", x"01", x"C8", x"85",
x"8F", x"84", x"90", x"60", x"A5", x"08", x"0A", x"69",
x"05", x"65", x"A7", x"A4", x"A8", x"90", x"01", x"C8",
x"85", x"A0", x"84", x"A1", x"60", x"90", x"80", x"00",
x"00", x"20", x"BF", x"00", x"20", x"7F", x"CB", x"20",
x"6E", x"CB", x"A5", x"AE", x"30", x"0D", x"A5", x"A9",
x"C9", x"90", x"90", x"09", x"A9", x"ED", x"A0", x"CE",
x"20", x"9A", x"D9", x"D0", x"7A", x"4C", x"DA", x"D9",
x"A5", x"09", x"05", x"0B", x"48", x"A5", x"0A", x"48",
x"A0", x"00", x"98", x"48", x"A5", x"8E", x"48", x"A5",
x"8D", x"48", x"20", x"F1", x"CE", x"68", x"85", x"8D",
x"68", x"85", x"8E", x"68", x"A8", x"BA", x"BD", x"02",
x"01", x"48", x"BD", x"01", x"01", x"48", x"A5", x"AC",
x"9D", x"02", x"01", x"A5", x"AD", x"9D", x"01", x"01",
x"C8", x"20", x"C5", x"00", x"C9", x"2C", x"F0", x"D2",
x"84", x"08", x"20", x"BF", x"CC", x"68", x"85", x"0A",
x"68", x"85", x"0B", x"29", x"7F", x"85", x"09", x"A6",
x"77", x"A5", x"78", x"86", x"A7", x"85", x"A8", x"C5",
x"7A", x"D0", x"04", x"E4", x"79", x"F0", x"39", x"A0",
x"00", x"B1", x"A7", x"C8", x"C5", x"8D", x"D0", x"06",
x"A5", x"8E", x"D1", x"A7", x"F0", x"16", x"C8", x"B1",
x"A7", x"18", x"65", x"A7", x"AA", x"C8", x"B1", x"A7",
x"65", x"A8", x"90", x"D7", x"A2", x"10", x"2C", x"A2",
x"08", x"4C", x"59", x"C2", x"A2", x"12", x"A5", x"09",
x"D0", x"F7", x"20", x"DC", x"CE", x"A5", x"08", x"A0",
x"04", x"D1", x"A7", x"D0", x"E7", x"4C", x"2A", x"D0",
x"20", x"DC", x"CE", x"20", x"2A", x"C2", x"A9", x"00",
x"A8", x"85", x"BA", x"A2", x"05", x"A5", x"8D", x"91",
x"A7", x"10", x"01", x"CA", x"C8", x"A5", x"8E", x"91",
x"A7", x"10", x"02", x"CA", x"CA", x"86", x"B9", x"A5",
x"08", x"C8", x"C8", x"C8", x"91", x"A7", x"A2", x"0B",
x"A9", x"00", x"24", x"09", x"50", x"08", x"68", x"18",
x"69", x"01", x"AA", x"68", x"69", x"00", x"C8", x"91",
x"A7", x"C8", x"8A", x"91", x"A7", x"20", x"8C", x"D0",
x"86", x"B9", x"85", x"BA", x"A4", x"6A", x"C6", x"08",
x"D0", x"DC", x"65", x"A1", x"B0", x"5D", x"85", x"A1",
x"A8", x"8A", x"65", x"A0", x"90", x"03", x"C8", x"F0",
x"52", x"20", x"2A", x"C2", x"85", x"79", x"84", x"7A",
x"A9", x"00", x"E6", x"BA", x"A4", x"B9", x"F0", x"05",
x"88", x"91", x"A0", x"D0", x"FB", x"C6", x"A1", x"C6",
x"BA", x"D0", x"F5", x"E6", x"A1", x"38", x"A5", x"79",
x"E5", x"A7", x"A0", x"02", x"91", x"A7", x"A5", x"7A",
x"C8", x"E5", x"A8", x"91", x"A7", x"A5", x"09", x"D0",
x"62", x"C8", x"B1", x"A7", x"85", x"08", x"A9", x"00",
x"85", x"B9", x"85", x"BA", x"C8", x"68", x"AA", x"85",
x"AC", x"68", x"85", x"AD", x"D1", x"A7", x"90", x"0E",
x"D0", x"06", x"C8", x"8A", x"D1", x"A7", x"90", x"07",
x"4C", x"84", x"CF", x"4C", x"57", x"C2", x"C8", x"A5",
x"BA", x"05", x"B9", x"18", x"F0", x"0A", x"20", x"8C",
x"D0", x"8A", x"65", x"AC", x"AA", x"98", x"A4", x"6A",
x"65", x"AD", x"86", x"B9", x"C6", x"08", x"D0", x"CA",
x"85", x"BA", x"A2", x"05", x"A5", x"8D", x"10", x"01",
x"CA", x"A5", x"8E", x"10", x"02", x"CA", x"CA", x"86",
x"70", x"A9", x"00", x"20", x"95", x"D0", x"8A", x"65",
x"A0", x"85", x"8F", x"98", x"65", x"A1", x"85", x"90",
x"A8", x"A5", x"8F", x"60", x"84", x"6A", x"B1", x"A7",
x"85", x"70", x"88", x"B1", x"A7", x"85", x"71", x"A9",
x"10", x"85", x"A5", x"A2", x"00", x"A0", x"00", x"8A",
x"0A", x"AA", x"98", x"2A", x"A8", x"B0", x"A4", x"06",
x"B9", x"26", x"BA", x"90", x"0B", x"18", x"8A", x"65",
x"70", x"AA", x"98", x"65", x"71", x"A8", x"B0", x"93",
x"C6", x"A5", x"D0", x"E3", x"60", x"A5", x"0A", x"F0",
x"03", x"20", x"E4", x"D3", x"20", x"64", x"D2", x"38",
x"A5", x"7B", x"E5", x"79", x"A8", x"A5", x"7C", x"E5",
x"7A", x"A2", x"00", x"86", x"0A", x"85", x"AA", x"84",
x"AB", x"A2", x"90", x"4C", x"83", x"D9", x"A4", x"11",
x"A9", x"00", x"F0", x"ED", x"A6", x"82", x"E8", x"D0",
x"A2", x"A2", x"16", x"2C", x"A2", x"20", x"4C", x"59",
x"C2", x"20", x"1F", x"D1", x"20", x"E4", x"D0", x"20",
x"C2", x"CC", x"A9", x"80", x"85", x"0D", x"20", x"E4",
x"CD", x"20", x"6E", x"CB", x"20", x"BF", x"CC", x"A9",
x"AC", x"20", x"C7", x"CC", x"48", x"A5", x"90", x"48",
x"A5", x"8F", x"48", x"A5", x"C7", x"48", x"A5", x"C6",
x"48", x"20", x"67", x"C7", x"4C", x"8D", x"D1", x"A9",
x"9F", x"20", x"C7", x"CC", x"09", x"80", x"85", x"0D",
x"20", x"EB", x"CD", x"85", x"96", x"84", x"97", x"4C",
x"6E", x"CB", x"20", x"1F", x"D1", x"A5", x"97", x"48",
x"A5", x"96", x"48", x"20", x"B9", x"CC", x"20", x"6E",
x"CB", x"68", x"85", x"96", x"68", x"85", x"97", x"A0",
x"02", x"B1", x"96", x"85", x"8F", x"AA", x"C8", x"B1",
x"96", x"F0", x"99", x"85", x"90", x"C8", x"B1", x"8F",
x"48", x"88", x"10", x"FA", x"A4", x"90", x"20", x"13",
x"D9", x"A5", x"C7", x"48", x"A5", x"C6", x"48", x"B1",
x"96", x"85", x"C6", x"C8", x"B1", x"96", x"85", x"C7",
x"A5", x"90", x"48", x"A5", x"8F", x"48", x"20", x"6B",
x"CB", x"68", x"85", x"96", x"68", x"85", x"97", x"20",
x"C5", x"00", x"F0", x"03", x"4C", x"D0", x"CC", x"68",
x"85", x"C6", x"68", x"85", x"C7", x"A0", x"00", x"68",
x"91", x"96", x"68", x"C8", x"91", x"96", x"68", x"C8",
x"91", x"96", x"68", x"C8", x"91", x"96", x"68", x"C8",
x"91", x"96", x"60", x"20", x"6E", x"CB", x"A0", x"00",
x"20", x"1E", x"DB", x"68", x"68", x"A9", x"FF", x"A0",
x"03", x"D0", x"12", x"A6", x"AC", x"A4", x"AD", x"86",
x"98", x"84", x"99", x"20", x"32", x"D2", x"86", x"AA",
x"84", x"AB", x"85", x"A9", x"60", x"A2", x"22", x"86",
x"06", x"86", x"07", x"85", x"B7", x"84", x"B8", x"85",
x"AA", x"84", x"AB", x"A0", x"FF", x"C8", x"B1", x"B7",
x"F0", x"0C", x"C5", x"06", x"F0", x"04", x"C5", x"07",
x"D0", x"F3", x"C9", x"22", x"F0", x"01", x"18", x"84",
x"A9", x"98", x"65", x"B7", x"85", x"B9", x"A6", x"B8",
x"90", x"01", x"E8", x"86", x"BA", x"A5", x"B8", x"F0",
x"04", x"C9", x"03", x"D0", x"0B", x"98", x"20", x"B3",
x"D1", x"A6", x"B7", x"A4", x"B8", x"20", x"C6", x"D3",
x"A6", x"5E", x"E0", x"6A", x"D0", x"05", x"A2", x"1C",
x"4C", x"59", x"C2", x"A5", x"A9", x"95", x"00", x"A5",
x"AA", x"95", x"01", x"A5", x"AB", x"95", x"02", x"A0",
x"00", x"86", x"AC", x"84", x"AD", x"84", x"B8", x"88",
x"84", x"0A", x"86", x"5F", x"E8", x"E8", x"E8", x"86",
x"5E", x"60", x"46", x"0C", x"48", x"49", x"FF", x"38",
x"65", x"7B", x"A4", x"7C", x"B0", x"01", x"88", x"C4",
x"7A", x"90", x"11", x"D0", x"04", x"C5", x"79", x"90",
x"0B", x"85", x"7B", x"84", x"7C", x"85", x"7D", x"84",
x"7E", x"AA", x"68", x"60", x"A2", x"0C", x"A5", x"0C",
x"30", x"B6", x"20", x"64", x"D2", x"A9", x"80", x"85",
x"0C", x"68", x"D0", x"D0", x"A6", x"7F", x"A5", x"80",
x"86", x"7B", x"85", x"7C", x"A0", x"00", x"84", x"97",
x"84", x"96", x"A5", x"79", x"A6", x"7A", x"85", x"A7",
x"86", x"A8", x"A9", x"61", x"A2", x"00", x"85", x"6A",
x"86", x"6B", x"C5", x"5E", x"F0", x"05", x"20", x"05",
x"D3", x"F0", x"F7", x"A9", x"07", x"85", x"9B", x"A5",
x"75", x"A6", x"76", x"85", x"6A", x"86", x"6B", x"E4",
x"78", x"D0", x"04", x"C5", x"77", x"F0", x"05", x"20",
x"FB", x"D2", x"F0", x"F3", x"85", x"A0", x"86", x"A1",
x"A9", x"03", x"85", x"9B", x"A5", x"A0", x"A6", x"A1",
x"E4", x"7A", x"D0", x"07", x"C5", x"79", x"D0", x"03",
x"4C", x"44", x"D3", x"85", x"6A", x"86", x"6B", x"A0",
x"00", x"B1", x"6A", x"AA", x"C8", x"B1", x"6A", x"08",
x"C8", x"B1", x"6A", x"65", x"A0", x"85", x"A0", x"C8",
x"B1", x"6A", x"65", x"A1", x"85", x"A1", x"28", x"10",
x"D3", x"8A", x"30", x"D0", x"C8", x"B1", x"6A", x"A0",
x"00", x"0A", x"69", x"05", x"65", x"6A", x"85", x"6A",
x"90", x"02", x"E6", x"6B", x"A6", x"6B", x"E4", x"A1",
x"D0", x"04", x"C5", x"A0", x"F0", x"BA", x"20", x"05",
x"D3", x"F0", x"F3", x"B1", x"6A", x"30", x"35", x"C8",
x"B1", x"6A", x"10", x"30", x"C8", x"B1", x"6A", x"F0",
x"2B", x"C8", x"B1", x"6A", x"AA", x"C8", x"B1", x"6A",
x"C5", x"7C", x"90", x"06", x"D0", x"1E", x"E4", x"7B",
x"B0", x"1A", x"C5", x"A8", x"90", x"16", x"D0", x"04",
x"E4", x"A7", x"90", x"10", x"86", x"A7", x"85", x"A8",
x"A5", x"6A", x"A6", x"6B", x"85", x"96", x"86", x"97",
x"A5", x"9B", x"85", x"9D", x"A5", x"9B", x"18", x"65",
x"6A", x"85", x"6A", x"90", x"02", x"E6", x"6B", x"A6",
x"6B", x"A0", x"00", x"60", x"A5", x"97", x"05", x"96",
x"F0", x"F5", x"A5", x"9D", x"29", x"04", x"4A", x"A8",
x"85", x"9D", x"B1", x"96", x"65", x"A7", x"85", x"A2",
x"A5", x"A8", x"69", x"00", x"85", x"A3", x"A5", x"7B",
x"A6", x"7C", x"85", x"A0", x"86", x"A1", x"20", x"E1",
x"C1", x"A4", x"9D", x"C8", x"A5", x"A0", x"91", x"96",
x"AA", x"E6", x"A1", x"A5", x"A1", x"C8", x"91", x"96",
x"4C", x"68", x"D2", x"A5", x"AD", x"48", x"A5", x"AC",
x"48", x"20", x"64", x"CC", x"20", x"70", x"CB", x"68",
x"85", x"B7", x"68", x"85", x"B8", x"A0", x"00", x"B1",
x"B7", x"18", x"71", x"AC", x"90", x"05", x"A2", x"1A",
x"4C", x"59", x"C2", x"20", x"B3", x"D1", x"20", x"B8",
x"D3", x"A5", x"98", x"A4", x"99", x"20", x"E8", x"D3",
x"20", x"CA", x"D3", x"A5", x"B7", x"A4", x"B8", x"20",
x"E8", x"D3", x"20", x"08", x"D2", x"4C", x"99", x"CB",
x"A0", x"00", x"B1", x"B7", x"48", x"C8", x"B1", x"B7",
x"AA", x"C8", x"B1", x"B7", x"A8", x"68", x"86", x"6A",
x"84", x"6B", x"A8", x"F0", x"0A", x"48", x"88", x"B1",
x"6A", x"91", x"7D", x"98", x"D0", x"F8", x"68", x"18",
x"65", x"7D", x"85", x"7D", x"90", x"02", x"E6", x"7E",
x"60", x"20", x"70", x"CB", x"A5", x"AC", x"A4", x"AD",
x"85", x"6A", x"84", x"6B", x"20", x"19", x"D4", x"08",
x"A0", x"00", x"B1", x"6A", x"48", x"C8", x"B1", x"6A",
x"AA", x"C8", x"B1", x"6A", x"A8", x"68", x"28", x"D0",
x"13", x"C4", x"7C", x"D0", x"0F", x"E4", x"7B", x"D0",
x"0B", x"48", x"18", x"65", x"7B", x"85", x"7B", x"90",
x"02", x"E6", x"7C", x"68", x"86", x"6A", x"84", x"6B",
x"60", x"C4", x"60", x"D0", x"0C", x"C5", x"5F", x"D0",
x"08", x"85", x"5E", x"E9", x"03", x"85", x"5F", x"A0",
x"00", x"60", x"20", x"DF", x"D4", x"8A", x"48", x"A9",
x"01", x"20", x"BB", x"D1", x"68", x"A0", x"00", x"91",
x"AA", x"68", x"68", x"4C", x"08", x"D2", x"20", x"9F",
x"D4", x"D1", x"98", x"98", x"90", x"04", x"B1", x"98",
x"AA", x"98", x"48", x"8A", x"48", x"20", x"BB", x"D1",
x"A5", x"98", x"A4", x"99", x"20", x"E8", x"D3", x"68",
x"A8", x"68", x"18", x"65", x"6A", x"85", x"6A", x"90",
x"02", x"E6", x"6B", x"98", x"20", x"CA", x"D3", x"4C",
x"08", x"D2", x"20", x"9F", x"D4", x"18", x"F1", x"98",
x"49", x"FF", x"4C", x"44", x"D4", x"A9", x"FF", x"85",
x"AD", x"20", x"C5", x"00", x"C9", x"29", x"F0", x"06",
x"20", x"C5", x"CC", x"20", x"DC", x"D4", x"20", x"9F",
x"D4", x"F0", x"4B", x"CA", x"8A", x"48", x"18", x"A2",
x"00", x"F1", x"98", x"B0", x"B6", x"49", x"FF", x"C5",
x"AD", x"90", x"B1", x"A5", x"AD", x"B0", x"AD", x"20",
x"BF", x"CC", x"68", x"A8", x"68", x"85", x"9D", x"68",
x"68", x"68", x"AA", x"68", x"85", x"98", x"68", x"85",
x"99", x"A5", x"9D", x"48", x"98", x"48", x"A0", x"00",
x"8A", x"60", x"20", x"C0", x"D4", x"4C", x"E0", x"D0",
x"20", x"E1", x"D3", x"A2", x"00", x"86", x"0A", x"A8",
x"60", x"20", x"C0", x"D4", x"F0", x"08", x"A0", x"00",
x"B1", x"6A", x"A8", x"4C", x"E0", x"D0", x"4C", x"87",
x"CF", x"20", x"BF", x"00", x"20", x"6B", x"CB", x"20",
x"F7", x"CE", x"A6", x"AC", x"D0", x"F0", x"A6", x"AD",
x"4C", x"C5", x"00", x"20", x"C0", x"D4", x"D0", x"03",
x"4C", x"36", x"D6", x"A6", x"C6", x"A4", x"C7", x"86",
x"B9", x"84", x"BA", x"A6", x"6A", x"86", x"C6", x"18",
x"65", x"6A", x"85", x"6C", x"A6", x"6B", x"86", x"C7",
x"90", x"01", x"E8", x"86", x"6D", x"A0", x"00", x"B1",
x"6C", x"48", x"A9", x"00", x"91", x"6C", x"20", x"C5",
x"00", x"20", x"32", x"DA", x"68", x"A0", x"00", x"91",
x"6C", x"A6", x"B9", x"A4", x"BA", x"86", x"C6", x"84",
x"C7", x"60", x"20", x"6B", x"CB", x"20", x"36", x"D5",
x"20", x"C5", x"CC", x"4C", x"DC", x"D4", x"A5", x"AE",
x"30", x"9C", x"A5", x"A9", x"C9", x"91", x"B0", x"96",
x"20", x"DA", x"D9", x"A5", x"AC", x"A4", x"AD", x"84",
x"14", x"85", x"15", x"60", x"A5", x"15", x"48", x"A5",
x"14", x"48", x"20", x"36", x"D5", x"A0", x"00", x"B1",
x"14", x"A8", x"68", x"85", x"14", x"68", x"85", x"15",
x"4C", x"E0", x"D0", x"20", x"2A", x"D5", x"8A", x"A0",
x"00", x"91", x"14", x"60", x"20", x"2A", x"D5", x"86",
x"91", x"A2", x"00", x"20", x"C5", x"00", x"F0", x"03",
x"20", x"30", x"D5", x"86", x"92", x"A0", x"00", x"B1",
x"14", x"45", x"92", x"25", x"91", x"F0", x"F8", x"60",
x"A9", x"4C", x"A0", x"DC", x"4C", x"A6", x"D5", x"20",
x"CB", x"D7", x"A5", x"AE", x"49", x"FF", x"85", x"AE",
x"45", x"B6", x"85", x"B7", x"A5", x"A9", x"4C", x"A9",
x"D5", x"20", x"D8", x"D6", x"90", x"3C", x"20", x"CB",
x"D7", x"D0", x"03", x"4C", x"3B", x"D9", x"A6", x"B8",
x"86", x"9E", x"A2", x"B1", x"A5", x"B1", x"A8", x"F0",
x"CE", x"38", x"E5", x"A9", x"F0", x"24", x"90", x"12",
x"84", x"A9", x"A4", x"B6", x"84", x"AE", x"49", x"FF",
x"69", x"00", x"A0", x"00", x"84", x"9E", x"A2", x"A9",
x"D0", x"04", x"A0", x"00", x"84", x"B8", x"C9", x"F9",
x"30", x"C7", x"A8", x"A5", x"B8", x"56", x"01", x"20",
x"EF", x"D6", x"24", x"B7", x"10", x"57", x"A0", x"A9",
x"E0", x"B1", x"F0", x"02", x"A0", x"B1", x"38", x"49",
x"FF", x"65", x"9E", x"85", x"B8", x"B9", x"04", x"00",
x"F5", x"04", x"85", x"AD", x"B9", x"03", x"00", x"F5",
x"03", x"85", x"AC", x"B9", x"02", x"00", x"F5", x"02",
x"85", x"AB", x"B9", x"01", x"00", x"F5", x"01", x"85",
x"AA", x"B0", x"03", x"20", x"86", x"D6", x"A0", x"00",
x"98", x"18", x"A6", x"AA", x"D0", x"4A", x"A6", x"AB",
x"86", x"AA", x"A6", x"AC", x"86", x"AB", x"A6", x"AD",
x"86", x"AC", x"A6", x"B8", x"86", x"AD", x"84", x"B8",
x"69", x"08", x"C9", x"20", x"D0", x"E4", x"A9", x"00",
x"85", x"A9", x"85", x"AE", x"60", x"65", x"9E", x"85",
x"B8", x"A5", x"AD", x"65", x"B5", x"85", x"AD", x"A5",
x"AC", x"65", x"B4", x"85", x"AC", x"A5", x"AB", x"65",
x"B3", x"85", x"AB", x"A5", x"AA", x"65", x"B2", x"85",
x"AA", x"4C", x"75", x"D6", x"69", x"01", x"06", x"B8",
x"26", x"AD", x"26", x"AC", x"26", x"AB", x"26", x"AA",
x"10", x"F2", x"38", x"E5", x"A9", x"B0", x"C7", x"49",
x"FF", x"69", x"01", x"85", x"A9", x"90", x"0E", x"E6",
x"A9", x"F0", x"42", x"66", x"AA", x"66", x"AB", x"66",
x"AC", x"66", x"AD", x"66", x"B8", x"60", x"A5", x"AE",
x"49", x"FF", x"85", x"AE", x"A5", x"AA", x"49", x"FF",
x"85", x"AA", x"A5", x"AB", x"49", x"FF", x"85", x"AB",
x"A5", x"AC", x"49", x"FF", x"85", x"AC", x"A5", x"AD",
x"49", x"FF", x"85", x"AD", x"A5", x"B8", x"49", x"FF",
x"85", x"B8", x"E6", x"B8", x"D0", x"0E", x"E6", x"AD",
x"D0", x"0A", x"E6", x"AC", x"D0", x"06", x"E6", x"AB",
x"D0", x"02", x"E6", x"AA", x"60", x"A2", x"0A", x"4C",
x"59", x"C2", x"A2", x"6D", x"B4", x"04", x"84", x"B8",
x"B4", x"03", x"94", x"04", x"B4", x"02", x"94", x"03",
x"B4", x"01", x"94", x"02", x"A4", x"B0", x"94", x"01",
x"69", x"08", x"30", x"E8", x"F0", x"E6", x"E9", x"08",
x"A8", x"A5", x"B8", x"B0", x"14", x"16", x"01", x"90",
x"02", x"F6", x"01", x"76", x"01", x"76", x"01", x"76",
x"02", x"76", x"03", x"76", x"04", x"6A", x"C8", x"D0",
x"EC", x"18", x"60", x"81", x"00", x"00", x"00", x"00",
x"03", x"7F", x"5E", x"56", x"CB", x"79", x"80", x"13",
x"9B", x"0B", x"64", x"80", x"76", x"38", x"93", x"16",
x"82", x"38", x"AA", x"3B", x"20", x"80", x"35", x"04",
x"F3", x"34", x"81", x"35", x"04", x"F3", x"34", x"80",
x"80", x"00", x"00", x"00", x"80", x"31", x"72", x"17",
x"F8", x"20", x"6A", x"D9", x"F0", x"02", x"10", x"03",
x"4C", x"87", x"CF", x"A5", x"A9", x"E9", x"7F", x"48",
x"A9", x"80", x"85", x"A9", x"A9", x"15", x"A0", x"D7",
x"20", x"A6", x"D5", x"A9", x"1A", x"A0", x"D7", x"20",
x"4E", x"D8", x"A9", x"FB", x"A0", x"D6", x"20", x"8F",
x"D5", x"A9", x"00", x"A0", x"D7", x"20", x"44", x"DD",
x"A9", x"1F", x"A0", x"D7", x"20", x"A6", x"D5", x"68",
x"20", x"BD", x"DA", x"A9", x"24", x"A0", x"D7", x"20",
x"CB", x"D7", x"D0", x"03", x"4C", x"CA", x"D7", x"20",
x"F6", x"D7", x"A9", x"00", x"85", x"6E", x"85", x"6F",
x"85", x"70", x"85", x"71", x"A5", x"B8", x"20", x"98",
x"D7", x"A5", x"AD", x"20", x"98", x"D7", x"A5", x"AC",
x"20", x"98", x"D7", x"A5", x"AB", x"20", x"98", x"D7",
x"A5", x"AA", x"20", x"9D", x"D7", x"4C", x"CE", x"D8",
x"D0", x"03", x"4C", x"C2", x"D6", x"4A", x"09", x"80",
x"A8", x"90", x"19", x"18", x"A5", x"71", x"65", x"B5",
x"85", x"71", x"A5", x"70", x"65", x"B4", x"85", x"70",
x"A5", x"6F", x"65", x"B3", x"85", x"6F", x"A5", x"6E",
x"65", x"B2", x"85", x"6E", x"66", x"6E", x"66", x"6F",
x"66", x"70", x"66", x"71", x"66", x"B8", x"98", x"4A",
x"D0", x"D6", x"60", x"85", x"6A", x"84", x"6B", x"A0",
x"04", x"B1", x"6A", x"85", x"B5", x"88", x"B1", x"6A",
x"85", x"B4", x"88", x"B1", x"6A", x"85", x"B3", x"88",
x"B1", x"6A", x"85", x"B6", x"45", x"AE", x"85", x"B7",
x"A5", x"B6", x"09", x"80", x"85", x"B2", x"88", x"B1",
x"6A", x"85", x"B1", x"A5", x"A9", x"60", x"A5", x"B1",
x"F0", x"1F", x"18", x"65", x"A9", x"90", x"04", x"30",
x"1D", x"18", x"2C", x"10", x"14", x"69", x"80", x"85",
x"A9", x"D0", x"03", x"4C", x"3A", x"D6", x"A5", x"B7",
x"85", x"AE", x"60", x"A5", x"AE", x"49", x"FF", x"30",
x"05", x"68", x"68", x"4C", x"36", x"D6", x"4C", x"BD",
x"D6", x"20", x"4B", x"D9", x"AA", x"F0", x"10", x"18",
x"69", x"02", x"B0", x"F2", x"A2", x"00", x"86", x"B7",
x"20", x"B6", x"D5", x"E6", x"A9", x"F0", x"E7", x"60",
x"84", x"20", x"00", x"00", x"00", x"20", x"4B", x"D9",
x"A9", x"38", x"A0", x"D8", x"A2", x"00", x"86", x"B7",
x"20", x"E1", x"D8", x"4C", x"51", x"D8", x"20", x"CB",
x"D7", x"F0", x"76", x"20", x"5A", x"D9", x"A9", x"00",
x"38", x"E5", x"A9", x"85", x"A9", x"20", x"F6", x"D7",
x"E6", x"A9", x"F0", x"BA", x"A2", x"FC", x"A9", x"01",
x"A4", x"B2", x"C4", x"AA", x"D0", x"10", x"A4", x"B3",
x"C4", x"AB", x"D0", x"0A", x"A4", x"B4", x"C4", x"AC",
x"D0", x"04", x"A4", x"B5", x"C4", x"AD", x"08", x"2A",
x"90", x"09", x"E8", x"95", x"71", x"F0", x"32", x"10",
x"34", x"A9", x"01", x"28", x"B0", x"0E", x"06", x"B5",
x"26", x"B4", x"26", x"B3", x"26", x"B2", x"B0", x"E6",
x"30", x"CE", x"10", x"E2", x"A8", x"A5", x"B5", x"E5",
x"AD", x"85", x"B5", x"A5", x"B4", x"E5", x"AC", x"85",
x"B4", x"A5", x"B3", x"E5", x"AB", x"85", x"B3", x"A5",
x"B2", x"E5", x"AA", x"85", x"B2", x"98", x"4C", x"8E",
x"D8", x"A9", x"40", x"D0", x"CE", x"0A", x"0A", x"0A",
x"0A", x"0A", x"0A", x"85", x"B8", x"28", x"4C", x"CE",
x"D8", x"A2", x"14", x"4C", x"59", x"C2", x"A5", x"6E",
x"85", x"AA", x"A5", x"6F", x"85", x"AB", x"A5", x"70",
x"85", x"AC", x"A5", x"71", x"85", x"AD", x"4C", x"16",
x"D6", x"85", x"6A", x"84", x"6B", x"A0", x"04", x"B1",
x"6A", x"85", x"AD", x"88", x"B1", x"6A", x"85", x"AC",
x"88", x"B1", x"6A", x"85", x"AB", x"88", x"B1", x"6A",
x"85", x"AE", x"09", x"80", x"85", x"AA", x"88", x"B1",
x"6A", x"85", x"A9", x"84", x"B8", x"60", x"A2", x"A4",
x"2C", x"A2", x"9F", x"A0", x"00", x"F0", x"04", x"A6",
x"91", x"A4", x"92", x"20", x"5A", x"D9", x"86", x"6A",
x"84", x"6B", x"A0", x"04", x"A5", x"AD", x"91", x"6A",
x"88", x"A5", x"AC", x"91", x"6A", x"88", x"A5", x"AB",
x"91", x"6A", x"88", x"A5", x"AE", x"09", x"7F", x"25",
x"AA", x"91", x"6A", x"88", x"A5", x"A9", x"91", x"6A",
x"84", x"B8", x"60", x"A5", x"B6", x"85", x"AE", x"A2",
x"05", x"B5", x"B0", x"95", x"A8", x"CA", x"D0", x"F9",
x"86", x"B8", x"60", x"20", x"5A", x"D9", x"A2", x"06",
x"B5", x"A8", x"95", x"B0", x"CA", x"D0", x"F9", x"86",
x"B8", x"60", x"A5", x"A9", x"F0", x"FB", x"06", x"B8",
x"90", x"F7", x"20", x"AE", x"D6", x"D0", x"F2", x"4C",
x"77", x"D6", x"A5", x"A9", x"F0", x"09", x"A5", x"AE",
x"2A", x"A9", x"FF", x"B0", x"02", x"A9", x"01", x"60",
x"20", x"6A", x"D9", x"85", x"AA", x"A9", x"00", x"85",
x"AB", x"A2", x"88", x"A5", x"AA", x"49", x"FF", x"2A",
x"A9", x"00", x"85", x"AD", x"85", x"AC", x"86", x"A9",
x"85", x"B8", x"85", x"AE", x"4C", x"11", x"D6", x"46",
x"AE", x"60", x"85", x"6C", x"84", x"6D", x"A0", x"00",
x"B1", x"6C", x"C8", x"AA", x"F0", x"C4", x"B1", x"6C",
x"45", x"AE", x"30", x"C2", x"E4", x"A9", x"D0", x"21",
x"B1", x"6C", x"09", x"80", x"C5", x"AA", x"D0", x"19",
x"C8", x"B1", x"6C", x"C5", x"AB", x"D0", x"12", x"C8",
x"B1", x"6C", x"C5", x"AC", x"D0", x"0B", x"C8", x"A9",
x"7F", x"C5", x"B8", x"B1", x"6C", x"E5", x"AD", x"F0",
x"28", x"A5", x"AE", x"90", x"02", x"49", x"FF", x"4C",
x"70", x"D9", x"A5", x"A9", x"F0", x"4A", x"38", x"E9",
x"A0", x"24", x"AE", x"10", x"09", x"AA", x"A9", x"FF",
x"85", x"B0", x"20", x"8C", x"D6", x"8A", x"A2", x"A9",
x"C9", x"F9", x"10", x"06", x"20", x"D8", x"D6", x"84",
x"B0", x"60", x"A8", x"A5", x"AE", x"29", x"80", x"46",
x"AA", x"05", x"AA", x"85", x"AA", x"20", x"EF", x"D6",
x"84", x"B0", x"60", x"A5", x"A9", x"C9", x"A0", x"B0",
x"20", x"20", x"DA", x"D9", x"84", x"B8", x"A5", x"AE",
x"84", x"AE", x"49", x"80", x"2A", x"A9", x"A0", x"85",
x"A9", x"A5", x"AD", x"85", x"06", x"4C", x"11", x"D6",
x"85", x"AA", x"85", x"AB", x"85", x"AC", x"85", x"AD",
x"A8", x"60", x"A0", x"00", x"A2", x"0A", x"94", x"A5",
x"CA", x"10", x"FB", x"90", x"0F", x"C9", x"2D", x"D0",
x"04", x"86", x"AF", x"F0", x"04", x"C9", x"2B", x"D0",
x"05", x"20", x"BF", x"00", x"90", x"5B", x"C9", x"2E",
x"F0", x"2E", x"C9", x"45", x"D0", x"30", x"20", x"BF",
x"00", x"90", x"17", x"C9", x"A5", x"F0", x"0E", x"C9",
x"2D", x"F0", x"0A", x"C9", x"A4", x"F0", x"08", x"C9",
x"2B", x"F0", x"04", x"D0", x"07", x"66", x"A8", x"20",
x"BF", x"00", x"90", x"5C", x"24", x"A8", x"10", x"0E",
x"A9", x"00", x"38", x"E5", x"A6", x"4C", x"88", x"DA",
x"66", x"A7", x"24", x"A7", x"50", x"C3", x"A5", x"A6",
x"38", x"E5", x"A5", x"85", x"A6", x"F0", x"12", x"10",
x"09", x"20", x"3D", x"D8", x"E6", x"A6", x"D0", x"F9",
x"F0", x"07", x"20", x"21", x"D8", x"C6", x"A6", x"D0",
x"F9", x"A5", x"AF", x"30", x"01", x"60", x"4C", x"B8",
x"DC", x"48", x"24", x"A7", x"10", x"02", x"E6", x"A5",
x"20", x"21", x"D8", x"68", x"38", x"E9", x"30", x"20",
x"BD", x"DA", x"4C", x"49", x"DA", x"48", x"20", x"4B",
x"D9", x"68", x"20", x"7B", x"D9", x"A5", x"B6", x"45",
x"AE", x"85", x"B7", x"A6", x"A9", x"4C", x"A9", x"D5",
x"A5", x"A6", x"C9", x"0A", x"90", x"09", x"A9", x"64",
x"24", x"A8", x"30", x"11", x"4C", x"BD", x"D6", x"0A",
x"0A", x"18", x"65", x"A6", x"0A", x"18", x"A0", x"00",
x"71", x"C6", x"38", x"E9", x"30", x"85", x"A6", x"4C",
x"6F", x"DA", x"9B", x"3E", x"BC", x"1F", x"FD", x"9E",
x"6E", x"6B", x"27", x"FD", x"9E", x"6E", x"6B", x"28",
x"00", x"A9", x"9E", x"A0", x"C1", x"20", x"19", x"DB",
x"A5", x"82", x"A6", x"81", x"85", x"AA", x"86", x"AB",
x"A2", x"90", x"38", x"20", x"88", x"D9", x"20", x"1C",
x"DB", x"4C", x"4A", x"C9", x"A0", x"01", x"A9", x"20",
x"24", x"AE", x"10", x"02", x"A9", x"2D", x"99", x"FF",
x"03", x"85", x"AE", x"84", x"B9", x"C8", x"A9", x"30",
x"A6", x"A9", x"D0", x"03", x"4C", x"3F", x"DC", x"A9",
x"00", x"E0", x"80", x"F0", x"02", x"B0", x"09", x"A9",
x"FC", x"A0", x"DA", x"20", x"67", x"D7", x"A9", x"F7",
x"85", x"A5", x"A9", x"F7", x"A0", x"DA", x"20", x"9A",
x"D9", x"F0", x"1E", x"10", x"12", x"A9", x"F2", x"A0",
x"DA", x"20", x"9A", x"D9", x"F0", x"02", x"10", x"0E",
x"20", x"21", x"D8", x"C6", x"A5", x"D0", x"EE", x"20",
x"3D", x"D8", x"E6", x"A5", x"D0", x"DC", x"20", x"88",
x"D5", x"20", x"DA", x"D9", x"A2", x"01", x"A5", x"A5",
x"18", x"69", x"0A", x"30", x"09", x"C9", x"0B", x"B0",
x"06", x"69", x"FF", x"AA", x"A9", x"02", x"38", x"E9",
x"02", x"85", x"A6", x"86", x"A5", x"8A", x"F0", x"02",
x"10", x"13", x"A4", x"B9", x"A9", x"2E", x"C8", x"99",
x"FF", x"03", x"8A", x"F0", x"06", x"A9", x"30", x"C8",
x"99", x"FF", x"03", x"84", x"B9", x"A0", x"00", x"A2",
x"80", x"A5", x"AD", x"18", x"79", x"54", x"DC", x"85",
x"AD", x"A5", x"AC", x"79", x"53", x"DC", x"85", x"AC",
x"A5", x"AB", x"79", x"52", x"DC", x"85", x"AB", x"A5",
x"AA", x"79", x"51", x"DC", x"85", x"AA", x"E8", x"B0",
x"04", x"10", x"DE", x"30", x"02", x"30", x"DA", x"8A",
x"90", x"04", x"49", x"FF", x"69", x"0A", x"69", x"2F",
x"C8", x"C8", x"C8", x"C8", x"84", x"8F", x"A4", x"B9",
x"C8", x"AA", x"29", x"7F", x"99", x"FF", x"03", x"C6",
x"A5", x"D0", x"06", x"A9", x"2E", x"C8", x"99", x"FF",
x"03", x"84", x"B9", x"A4", x"8F", x"8A", x"49", x"FF",
x"29", x"80", x"AA", x"C0", x"24", x"D0", x"AA", x"A4",
x"B9", x"B9", x"FF", x"03", x"88", x"C9", x"30", x"F0",
x"F8", x"C9", x"2E", x"F0", x"01", x"C8", x"A9", x"2B",
x"A6", x"A6", x"F0", x"2E", x"10", x"08", x"A9", x"00",
x"38", x"E5", x"A6", x"AA", x"A9", x"2D", x"99", x"01",
x"04", x"A9", x"45", x"99", x"00", x"04", x"8A", x"A2",
x"2F", x"38", x"E8", x"E9", x"0A", x"B0", x"FB", x"69",
x"3A", x"99", x"03", x"04", x"8A", x"99", x"02", x"04",
x"A9", x"00", x"99", x"04", x"04", x"F0", x"08", x"99",
x"FF", x"03", x"A9", x"00", x"99", x"00", x"04", x"A9",
x"00", x"A0", x"04", x"60", x"80", x"00", x"00", x"00",
x"00", x"FA", x"0A", x"1F", x"00", x"00", x"98", x"96",
x"80", x"FF", x"F0", x"BD", x"C0", x"00", x"01", x"86",
x"A0", x"FF", x"FF", x"D8", x"F0", x"00", x"00", x"03",
x"E8", x"FF", x"FF", x"FF", x"9C", x"00", x"00", x"00",
x"0A", x"FF", x"FF", x"FF", x"FF", x"20", x"4B", x"D9",
x"A9", x"4C", x"A0", x"DC", x"20", x"E1", x"D8", x"F0",
x"70", x"A5", x"B1", x"D0", x"03", x"4C", x"38", x"D6",
x"A2", x"96", x"A0", x"00", x"20", x"13", x"D9", x"A5",
x"B6", x"10", x"0F", x"20", x"0B", x"DA", x"A9", x"96",
x"A0", x"00", x"20", x"9A", x"D9", x"D0", x"03", x"98",
x"A4", x"06", x"20", x"3D", x"D9", x"98", x"48", x"20",
x"29", x"D7", x"A9", x"96", x"A0", x"00", x"20", x"67",
x"D7", x"20", x"F1", x"DC", x"68", x"4A", x"90", x"0A",
x"A5", x"A9", x"F0", x"06", x"A5", x"AE", x"49", x"FF",
x"85", x"AE", x"60", x"81", x"38", x"AA", x"3B", x"29",
x"07", x"71", x"34", x"58", x"3E", x"56", x"74", x"16",
x"7E", x"B3", x"1B", x"77", x"2F", x"EE", x"E3", x"85",
x"7A", x"1D", x"84", x"1C", x"2A", x"7C", x"63", x"59",
x"58", x"0A", x"7E", x"75", x"FD", x"E7", x"C6", x"80",
x"31", x"72", x"18", x"10", x"81", x"00", x"00", x"00",
x"00", x"A9", x"C3", x"A0", x"DC", x"20", x"67", x"D7",
x"A5", x"B8", x"69", x"50", x"90", x"03", x"20", x"62",
x"D9", x"85", x"9E", x"20", x"4E", x"D9", x"A5", x"A9",
x"C9", x"88", x"90", x"03", x"20", x"13", x"D8", x"20",
x"0B", x"DA", x"A5", x"06", x"18", x"69", x"81", x"F0",
x"F3", x"38", x"E9", x"01", x"48", x"A2", x"05", x"B5",
x"B1", x"B4", x"A9", x"95", x"A9", x"94", x"B1", x"CA",
x"10", x"F5", x"A5", x"9E", x"85", x"B8", x"20", x"92",
x"D5", x"20", x"B8", x"DC", x"A9", x"C8", x"A0", x"DC",
x"20", x"5A", x"DD", x"A9", x"00", x"85", x"B7", x"68",
x"20", x"F8", x"D7", x"60", x"85", x"B9", x"84", x"BA",
x"20", x"09", x"D9", x"A9", x"9F", x"20", x"67", x"D7",
x"20", x"5E", x"DD", x"A9", x"9F", x"A0", x"00", x"4C",
x"67", x"D7", x"85", x"B9", x"84", x"BA", x"20", x"06",
x"D9", x"B1", x"B9", x"85", x"AF", x"A4", x"B9", x"C8",
x"98", x"D0", x"02", x"E6", x"BA", x"85", x"B9", x"A4",
x"BA", x"20", x"67", x"D7", x"A5", x"B9", x"A4", x"BA",
x"18", x"69", x"05", x"90", x"01", x"C8", x"85", x"B9",
x"84", x"BA", x"20", x"A6", x"D5", x"A9", x"A4", x"A0",
x"00", x"C6", x"AF", x"D0", x"E4", x"60", x"98", x"35",
x"44", x"7A", x"68", x"28", x"B1", x"46", x"20", x"6A",
x"D9", x"AA", x"30", x"18", x"A9", x"D7", x"A0", x"00",
x"20", x"E1", x"D8", x"8A", x"F0", x"E7", x"A9", x"8E",
x"A0", x"DD", x"20", x"67", x"D7", x"A9", x"92", x"A0",
x"DD", x"20", x"A6", x"D5", x"A6", x"AD", x"A5", x"AA",
x"85", x"AD", x"86", x"AA", x"A9", x"00", x"85", x"AE",
x"A5", x"A9", x"85", x"B8", x"A9", x"80", x"85", x"A9",
x"20", x"16", x"D6", x"A2", x"D7", x"A0", x"00", x"4C",
x"13", x"D9", x"A9", x"4E", x"A0", x"DE", x"20", x"A6",
x"D5", x"20", x"4B", x"D9", x"A9", x"53", x"A0", x"DE",
x"A6", x"B6", x"20", x"46", x"D8", x"20", x"4B", x"D9",
x"20", x"0B", x"DA", x"A9", x"00", x"85", x"B7", x"20",
x"92", x"D5", x"A9", x"58", x"A0", x"DE", x"20", x"8F",
x"D5", x"A5", x"AE", x"48", x"10", x"0D", x"20", x"88",
x"D5", x"A5", x"AE", x"30", x"09", x"A5", x"0F", x"49",
x"FF", x"85", x"0F", x"20", x"B8", x"DC", x"A9", x"58",
x"A0", x"DE", x"20", x"A6", x"D5", x"68", x"10", x"03",
x"20", x"B8", x"DC", x"A9", x"5D", x"A0", x"DE", x"4C",
x"44", x"DD", x"20", x"09", x"D9", x"A9", x"00", x"85",
x"0F", x"20", x"D9", x"DD", x"A2", x"96", x"A0", x"00",
x"20", x"CF", x"DD", x"A9", x"9F", x"A0", x"00", x"20",
x"E1", x"D8", x"A9", x"00", x"85", x"AE", x"A5", x"0F",
x"20", x"4A", x"DE", x"A9", x"96", x"A0", x"00", x"4C",
x"4E", x"D8", x"48", x"4C", x"0B", x"DE", x"81", x"49",
x"0F", x"DA", x"A2", x"83", x"49", x"0F", x"DA", x"A2",
x"7F", x"00", x"00", x"00", x"00", x"05", x"84", x"E6",
x"1A", x"2D", x"1B", x"86", x"28", x"07", x"FB", x"F8",
x"87", x"99", x"68", x"89", x"01", x"87", x"23", x"35",
x"DF", x"E1", x"86", x"A5", x"5D", x"E7", x"28", x"83",
x"49", x"0F", x"DA", x"A2", x"A1", x"54", x"46", x"8F",
x"13", x"8F", x"52", x"43", x"89", x"CD", x"E6", x"C6",
x"D0", x"02", x"E6", x"C7", x"AD", x"60", x"EA", x"C9",
x"3A", x"B0", x"0A", x"C9", x"20", x"F0", x"EF", x"38",
x"E9", x"30", x"38", x"E9", x"D0", x"60", x"80", x"4F",
x"C7", x"52", x"58", x"A2", x"FF", x"86", x"82", x"A2",
x"FE", x"9A", x"A9", x"A3", x"A0", x"DE", x"85", x"01",
x"84", x"02", x"A9", x"4C", x"85", x"00", x"85", x"9C",
x"85", x"BB", x"85", x"03", x"20", x"43", x"DF", x"EA",
x"A9", x"87", x"A0", x"CF", x"85", x"04", x"84", x"05",
x"A9", x"20", x"85", x"12", x"A9", x"1E", x"85", x"13",
x"A2", x"1C", x"BD", x"85", x"DE", x"95", x"BE", x"CA",
x"D0", x"F8", x"A9", x"03", x"85", x"9B", x"8A", x"85",
x"B0", x"85", x"60", x"48", x"85", x"10", x"20", x"00",
x"C9", x"A2", x"61", x"86", x"5E", x"A9", x"AF", x"A0",
x"DF", x"20", x"4A", x"C9", x"20", x"E7", x"C9", x"86",
x"C6", x"84", x"C7", x"20", x"BF", x"00", x"A8", x"D0",
x"2B", x"A9", x"11", x"A0", x"04", x"85", x"73", x"84",
x"74", x"85", x"14", x"84", x"15", x"A0", x"00", x"E6",
x"14", x"D0", x"08", x"E6", x"15", x"A5", x"15", x"C5",
x"BC", x"F0", x"1D", x"A9", x"55", x"91", x"14", x"D1",
x"14", x"D0", x"15", x"0A", x"91", x"14", x"D1", x"14",
x"D0", x"0E", x"F0", x"E3", x"20", x"C5", x"00", x"20",
x"DA", x"C7", x"A8", x"F0", x"03", x"4C", x"D0", x"CC",
x"A5", x"14", x"A4", x"15", x"85", x"7F", x"84", x"80",
x"4C", x"70", x"DF", x"A9", x"60", x"85", x"BC", x"A2",
x"42", x"A0", x"40", x"BD", x"00", x"B0", x"5D", x"00",
x"B0", x"CA", x"CA", x"CA", x"D0", x"F8", x"C9", x"4C",
x"D0", x"02", x"84", x"BC", x"60", x"C9", x"03", x"D0",
x"FB", x"A9", x"00", x"85", x"C7", x"4C", x"58", x"C6",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"A2", x"11", x"A0", x"04", x"86", x"73", x"84", x"74",
x"A0", x"00", x"98", x"91", x"73", x"E6", x"73", x"D0",
x"02", x"E6", x"74", x"20", x"67", x"C4", x"A5", x"73",
x"A4", x"74", x"20", x"2A", x"C2", x"20", x"00", x"C9",
x"A5", x"7F", x"38", x"E5", x"73", x"AA", x"A5", x"80",
x"E5", x"74", x"20", x"0C", x"DB", x"A9", x"EB", x"A0",
x"DF", x"20", x"4A", x"C9", x"A9", x"00", x"A0", x"C9",
x"85", x"01", x"84", x"02", x"4C", x"7F", x"C2", x"0C",
x"20", x"20", x"3E", x"45", x"41", x"47", x"4C", x"45",
x"3C", x"20", x"45", x"58", x"54", x"45", x"4E", x"44",
x"45", x"44", x"20", x"42", x"41", x"53", x"49", x"43",
x"0D", x"0A", x"0A", x"20", x"20", x"20", x"20", x"20",
x"56", x"20", x"31", x"2E", x"30", x"20", x"28", x"43",
x"29", x"20", x"38", x"35", x"0D", x"0A", x"0A", x"0A",
x"4D", x"45", x"4D", x"20", x"53", x"49", x"5A", x"45",
x"20", x"20", x"00", x"20", x"42", x"59", x"54", x"45",
x"53", x"20", x"46", x"52", x"45", x"45", x"0D", x"0A",
x"0A", x"00", x"20", x"C5", x"00", x"4C", x"9D", x"C8"
	);
begin
	process(clk)
	begin
		if rising_edge(clk) then
			data <= romData(conv_integer(addr));
		end if;
	end process;
end architecture;

