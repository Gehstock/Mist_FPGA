library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity pickin_tile_bit1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of pickin_tile_bit1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"3E",X"41",X"41",X"41",X"41",X"41",X"3E",X"00",X"00",X"00",X"7F",X"20",X"10",X"00",X"00",
		X"00",X"31",X"49",X"49",X"49",X"49",X"49",X"27",X"00",X"46",X"69",X"59",X"49",X"41",X"41",X"41",
		X"00",X"04",X"7F",X"44",X"44",X"24",X"14",X"0C",X"00",X"46",X"49",X"49",X"49",X"49",X"49",X"79",
		X"00",X"46",X"49",X"49",X"49",X"49",X"49",X"3E",X"00",X"60",X"50",X"48",X"47",X"40",X"40",X"40",
		X"00",X"36",X"49",X"49",X"49",X"49",X"49",X"36",X"00",X"3E",X"49",X"49",X"49",X"49",X"49",X"31",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"48",X"48",X"48",X"48",X"48",X"3F",
		X"00",X"36",X"49",X"49",X"49",X"49",X"49",X"7F",X"00",X"41",X"41",X"41",X"41",X"41",X"41",X"3E",
		X"00",X"3E",X"41",X"41",X"41",X"41",X"41",X"7F",X"00",X"41",X"41",X"49",X"49",X"49",X"49",X"7F",
		X"00",X"40",X"40",X"48",X"48",X"48",X"48",X"7F",X"00",X"4F",X"49",X"49",X"41",X"41",X"41",X"3E",
		X"00",X"7F",X"08",X"08",X"08",X"08",X"08",X"7F",X"00",X"00",X"00",X"00",X"7F",X"00",X"00",X"00",
		X"00",X"7E",X"01",X"01",X"01",X"01",X"01",X"06",X"00",X"41",X"22",X"14",X"08",X"04",X"02",X"7F",
		X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"7F",X"00",X"7F",X"20",X"10",X"08",X"10",X"20",X"7F",
		X"00",X"7F",X"02",X"04",X"08",X"10",X"20",X"7F",X"00",X"3E",X"41",X"41",X"41",X"41",X"41",X"3E",
		X"00",X"30",X"48",X"48",X"48",X"48",X"48",X"7F",X"00",X"3D",X"42",X"45",X"41",X"41",X"41",X"3E",
		X"00",X"31",X"4A",X"4C",X"48",X"48",X"48",X"7F",X"00",X"46",X"49",X"49",X"49",X"49",X"49",X"31",
		X"00",X"40",X"40",X"40",X"7F",X"40",X"40",X"40",X"00",X"7E",X"01",X"01",X"01",X"01",X"01",X"7E",
		X"00",X"78",X"04",X"02",X"01",X"02",X"04",X"78",X"00",X"7C",X"02",X"01",X"06",X"01",X"02",X"7C",
		X"00",X"41",X"22",X"14",X"08",X"14",X"22",X"41",X"00",X"40",X"20",X"10",X"0F",X"10",X"20",X"40",
		X"00",X"41",X"61",X"51",X"49",X"45",X"43",X"41",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"60",X"10",X"00",X"00",X"00",X"00",X"00",X"60",X"10",X"00",X"60",X"10",
		X"00",X"10",X"60",X"00",X"10",X"60",X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"08",X"08",X"00",
		X"00",X"40",X"20",X"10",X"08",X"04",X"02",X"01",X"00",X"08",X"08",X"08",X"7F",X"08",X"08",X"08",
		X"00",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"00",X"08",X"08",X"08",X"2A",X"08",X"08",X"08",
		X"00",X"00",X"7D",X"00",X"00",X"7D",X"00",X"00",X"7E",X"C3",X"A5",X"A5",X"A5",X"BD",X"C3",X"7E",
		X"F6",X"F6",X"00",X"00",X"F6",X"F6",X"00",X"00",X"FA",X"FA",X"00",X"00",X"FA",X"FA",X"00",X"00",
		X"00",X"00",X"00",X"F6",X"F6",X"00",X"00",X"00",X"00",X"00",X"00",X"FA",X"FA",X"00",X"00",X"00",
		X"00",X"00",X"00",X"E0",X"C0",X"00",X"00",X"00",X"00",X"E0",X"C0",X"00",X"E0",X"C0",X"00",X"00",
		X"00",X"60",X"E0",X"00",X"60",X"E0",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"38",X"10",X"00",X"40",X"02",X"07",X"D7",X"D0",X"D7",X"80",X"0F",X"20",X"3F",X"00",
		X"02",X"20",X"70",X"21",X"00",X"04",X"0E",X"04",X"07",X"0C",X"1F",X"39",X"2C",X"18",X"1F",X"0F",
		X"00",X"00",X"00",X"10",X"38",X"10",X"00",X"40",X"D7",X"D0",X"D7",X"80",X"0F",X"10",X"1F",X"00",
		X"04",X"0E",X"04",X"00",X"20",X"70",X"21",X"00",X"07",X"0C",X"1F",X"39",X"2C",X"18",X"1F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D7",X"D0",X"D7",X"80",X"0F",X"10",X"1F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"0C",X"1F",X"39",X"2C",X"18",X"1F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D7",X"D0",X"D7",X"80",X"0F",X"00",X"3F",X"D0",
		X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"FF",X"A0",X"AE",X"12",X"0A",X"0A",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"06",X"1F",X"00",X"00",X"00",X"11",X"17",X"97",X"07",X"05",
		X"1D",X"1D",X"01",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"D5",X"54",X"54",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"36",X"FF",X"00",X"00",X"00",X"00",X"09",X"2B",X"2B",X"AB",
		X"EA",X"EA",X"46",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"28",X"44",X"82",X"44",X"28",X"10",
		X"00",X"03",X"01",X"00",X"01",X"00",X"03",X"00",X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",
		X"81",X"01",X"01",X"01",X"01",X"01",X"02",X"FC",X"3F",X"40",X"80",X"80",X"80",X"80",X"80",X"81",
		X"FC",X"02",X"01",X"01",X"01",X"01",X"01",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"FF",
		X"FF",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"80",X"80",X"80",X"80",X"80",X"40",X"3F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",X"FF",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"00",X"00",X"00",X"00",X"00",X"18",X"6C",X"FE",X"00",X"00",X"78",X"B8",X"90",X"D0",X"50",X"50",
		X"D7",X"C5",X"8D",X"01",X"00",X"00",X"01",X"00",X"50",X"50",X"50",X"50",X"50",X"90",X"B8",X"3C",
		X"04",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"04",X"08",X"10",X"3E",X"00",X"1A",
		X"24",X"24",X"24",X"3E",X"00",X"3E",X"02",X"02",X"02",X"3E",X"00",X"20",X"20",X"3E",X"20",X"20",
		X"00",X"22",X"2A",X"2A",X"2A",X"3E",X"00",X"1A",X"24",X"24",X"24",X"3E",X"00",X"00",X"00",X"00",
		X"00",X"02",X"02",X"02",X"02",X"3E",X"00",X"3E",X"02",X"02",X"02",X"3E",X"00",X"22",X"22",X"22",
		X"22",X"3E",X"00",X"22",X"2A",X"2A",X"2A",X"3E",X"00",X"1A",X"24",X"24",X"24",X"3E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"22",X"2A",X"2A",X"2A",X"3E",X"00",X"2E",X"2A",X"2A",X"2A",X"3A",
		X"00",X"1E",X"24",X"24",X"24",X"1E",X"00",X"1A",X"24",X"24",X"24",X"3E",X"00",X"22",X"2A",X"2A",
		X"2A",X"3E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",
		X"20",X"3E",X"20",X"20",X"00",X"3E",X"04",X"08",X"10",X"3E",X"00",X"22",X"2A",X"2A",X"2A",X"3E",
		X"00",X"3E",X"10",X"08",X"10",X"3E",X"00",X"22",X"2A",X"2A",X"2A",X"3E",X"00",X"22",X"22",X"22",
		X"22",X"3E",X"00",X"1E",X"24",X"24",X"24",X"1E",X"00",X"20",X"28",X"28",X"28",X"3E",X"00",X"20",
		X"28",X"28",X"28",X"3E",X"00",X"22",X"2A",X"2A",X"2A",X"3E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"2A",X"2A",X"2A",X"3E",X"00",X"22",X"22",X"22",X"22",
		X"3E",X"00",X"3E",X"04",X"08",X"10",X"3E",X"00",X"1E",X"24",X"24",X"24",X"1E",X"00",X"38",X"04",
		X"02",X"04",X"38",X"00",X"1C",X"22",X"22",X"22",X"3E",X"00",X"1E",X"24",X"24",X"24",X"1E",X"00",
		X"00",X"00",X"00",X"00",X"22",X"2A",X"2A",X"2A",X"3E",X"00",X"22",X"22",X"22",X"22",X"3E",X"00",
		X"3E",X"04",X"08",X"10",X"3E",X"00",X"1E",X"24",X"24",X"24",X"1E",X"00",X"38",X"04",X"02",X"04",
		X"38",X"00",X"1E",X"24",X"24",X"24",X"1A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"2A",
		X"2A",X"2A",X"3E",X"00",X"1A",X"24",X"24",X"24",X"3E",X"00",X"3E",X"02",X"02",X"02",X"3E",X"00",
		X"20",X"20",X"3E",X"20",X"20",X"00",X"3E",X"00",X"00",X"1A",X"24",X"24",X"24",X"3E",X"00",X"22",
		X"22",X"22",X"22",X"3E",X"00",X"20",X"2A",X"2A",X"2A",X"3E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"2A",X"2A",X"2A",X"3E",X"00",X"20",X"20",X"3E",
		X"20",X"20",X"00",X"3E",X"00",X"1A",X"24",X"24",X"24",X"3E",X"00",X"38",X"04",X"02",X"3C",X"02",
		X"08",X"08",X"08",X"08",X"08",X"0C",X"06",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"08",X"08",X"08",X"08",X"08",X"18",X"30",X"E0",X"E0",X"30",X"18",X"08",X"08",X"08",X"08",X"08",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"06",X"0C",X"08",X"08",X"08",X"08",X"08",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"20",X"20",X"20",X"60",X"60",X"41",X"E3",X"E3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"E0",X"E0",X"E0",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"0F",X"3F",X"FF",X"FF",X"FF",X"E7",X"87",X"07",X"07",X"07",X"07",X"87",X"E7",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"03",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"E0",X"E0",X"20",X"00",X"00",X"00",
		X"3F",X"0F",X"07",X"07",X"07",X"07",X"07",X"07",X"00",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"80",
		X"07",X"3F",X"3F",X"3F",X"1F",X"1F",X"1F",X"0F",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"E0",
		X"0F",X"0F",X"07",X"07",X"07",X"07",X"07",X"3F",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"80",X"00",X"00",X"00",
		X"3F",X"07",X"07",X"07",X"07",X"C7",X"F7",X"FF",X"FF",X"7F",X"1F",X"07",X"01",X"00",X"00",X"00",
		X"00",X"01",X"07",X"1F",X"7F",X"FF",X"FC",X"F8",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"07",X"07",X"07",X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"07",X"07",X"07",X"04",X"00",X"00",X"00",X"00",X"00",
		X"07",X"02",X"02",X"02",X"02",X"02",X"02",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",
		X"BF",X"3F",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"3F",X"BF",
		X"FD",X"FC",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FC",X"FD",
		X"00",X"00",X"F8",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"F8",X"00",X"00",
		X"00",X"00",X"1F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",X"00",X"00",
		X"3F",X"41",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"41",X"3F",
		X"3F",X"40",X"80",X"80",X"80",X"80",X"80",X"FF",X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",
		X"81",X"81",X"81",X"81",X"81",X"81",X"82",X"FC",X"FC",X"82",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"82",X"FC",X"FC",X"02",X"01",X"01",X"01",X"01",X"01",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"02",X"FC",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"FF",
		X"81",X"01",X"01",X"01",X"01",X"01",X"02",X"FC",X"FF",X"80",X"80",X"80",X"80",X"80",X"40",X"3F",
		X"FC",X"02",X"01",X"01",X"01",X"01",X"01",X"81",X"3F",X"40",X"80",X"80",X"80",X"80",X"80",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"80",X"80",X"80",X"80",X"80",X"40",X"3F",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",
		X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",
		X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",
		X"01",X"01",X"01",X"03",X"03",X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"7C",X"3C",X"1C",X"06",X"02",X"00",X"00",X"00",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"FC",X"FC",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"FC",X"FE",X"FB",X"F1",
		X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"03",X"1F",X"3F",X"7E",X"FE",X"FC",X"FC",
		X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"18",X"1E",X"0F",X"07",
		X"E0",X"70",X"38",X"1C",X"0E",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"00",X"F8",X"FF",X"0F",X"03",X"01",X"00",X"00",X"1F",X"0F",X"07",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"30",X"3C",X"1E",X"0F",X"07",X"03",X"01",X"00",X"00",X"00",X"00",
		X"C0",X"E0",X"F0",X"FC",X"7E",X"3F",X"3F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"3C",X"1E",X"1E",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",
		X"00",X"60",X"78",X"3C",X"3E",X"1C",X"00",X"00",X"0F",X"07",X"07",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"7F",X"3F",X"3F",X"1F",X"1F",X"1F",X"0F",X"03",X"03",X"03",X"03",X"03",X"C3",X"C3",X"E7",
		X"07",X"07",X"03",X"03",X"03",X"03",X"03",X"03",X"3C",X"3C",X"1E",X"1E",X"0F",X"0F",X"07",X"07",
		X"0F",X"07",X"03",X"C1",X"E0",X"F0",X"F8",X"78",X"00",X"00",X"00",X"18",X"1C",X"1E",X"1F",X"0F",
		X"07",X"07",X"03",X"01",X"01",X"00",X"00",X"00",X"7E",X"7F",X"3F",X"3F",X"3F",X"1E",X"1F",X"0F",
		X"07",X"03",X"00",X"00",X"00",X"00",X"70",X"7C",X"E0",X"F0",X"F8",X"FC",X"FE",X"7F",X"3F",X"1F",
		X"0C",X"0C",X"04",X"06",X"02",X"03",X"81",X"C0",X"00",X"00",X"00",X"00",X"0F",X"1F",X"1F",X"1E",
		X"1F",X"0F",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"18",X"1E",X"1F",
		X"06",X"07",X"07",X"03",X"01",X"00",X"00",X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"04",
		X"0C",X"1E",X"1F",X"1F",X"0F",X"0F",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DC",X"8F",X"07",X"01",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"C0",X"C0",X"E0",X"F0",X"F8",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"E0",X"F0",X"F8",X"FC",X"7F",X"1F",X"07",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"E0",X"E0",X"F0",X"F8",X"7F",X"1F",
		X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"E0",X"F0",X"F9",X"3F",X"0F",X"01",X"00",X"00",
		X"40",X"61",X"31",X"1B",X"0F",X"0F",X"87",X"C3",X"70",X"30",X"18",X"08",X"04",X"02",X"81",X"81",
		X"07",X"03",X"01",X"00",X"00",X"80",X"C0",X"E0",X"80",X"C0",X"C0",X"E0",X"F0",X"FF",X"7F",X"1F",
		X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"83",X"C1",X"E0",X"F0",X"F9",X"3F",X"1F",
		X"0F",X"87",X"C3",X"60",X"70",X"38",X"1C",X"0E",X"00",X"00",X"00",X"80",X"C0",X"E0",X"F0",X"1C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"F0",X"F8",X"FC",X"3C",X"0E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1C",X"1C",X"3C",X"7C",X"FC",X"FC",X"F8",X"C0",X"C0",X"80",X"40",X"60",X"30",X"38",X"38",X"18",
		X"1C",X"1C",X"1C",X"1C",X"3C",X"78",X"F8",X"E0",X"40",X"60",X"30",X"30",X"38",X"18",X"18",X"1C",
		X"C0",X"E0",X"F0",X"F8",X"FC",X"80",X"00",X"80",X"FC",X"F8",X"F0",X"E0",X"80",X"00",X"00",X"80",
		X"18",X"08",X"0C",X"0C",X"0E",X"1E",X"1E",X"3E",X"80",X"00",X"00",X"80",X"40",X"40",X"20",X"10",
		X"38",X"38",X"3C",X"7C",X"FC",X"F8",X"F8",X"F0",X"C0",X"80",X"80",X"80",X"40",X"60",X"20",X"30",
		X"00",X"80",X"C0",X"E0",X"F0",X"F8",X"F8",X"F0",X"FC",X"FC",X"FC",X"FC",X"38",X"00",X"00",X"00",
		X"00",X"80",X"40",X"60",X"20",X"30",X"38",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"F0",X"F8",X"FC",X"3C",X"0E",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"55",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"AA",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"AA",
		X"55",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"55",X"03",X"07",X"0F",X"1F",X"3F",X"7F",X"FF",
		X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"AA",X"FF",X"7F",X"3F",X"1F",X"0F",X"07",X"03",X"AB",
		X"55",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"55",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"AA",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"AA",
		X"FF",X"FF",X"3F",X"9F",X"0F",X"87",X"03",X"81",X"FF",X"FE",X"FD",X"F8",X"F1",X"E0",X"C1",X"80",
		X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"AA",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"55",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"01",X"83",X"07",X"8F",X"1F",X"BF",X"7F",X"FF",X"81",X"C0",X"E1",X"F0",X"F9",X"FC",X"FF",X"FF",
		X"55",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"55",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"AA",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"AA",
		X"D5",X"C0",X"E0",X"F0",X"F8",X"FC",X"FE",X"FF",X"55",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"FF",X"FE",X"FC",X"F8",X"F0",X"E0",X"C0",X"AA",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"AA",
		X"55",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"55",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"AA",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"01",X"03",X"07",X"2F",X"1F",X"00",X"00",X"98",X"C4",X"E8",X"F0",X"F8",X"FC",
		X"1F",X"1F",X"2F",X"07",X"03",X"01",X"00",X"00",X"FE",X"FC",X"F8",X"F0",X"E6",X"C1",X"86",X"00",
		X"00",X"00",X"00",X"01",X"03",X"07",X"2F",X"1F",X"00",X"00",X"86",X"C1",X"E6",X"F0",X"F8",X"FC",
		X"1F",X"1F",X"2F",X"07",X"03",X"01",X"00",X"00",X"FE",X"FC",X"F8",X"F0",X"E8",X"C4",X"98",X"00",
		X"00",X"00",X"00",X"11",X"2B",X"27",X"0F",X"1F",X"00",X"04",X"8A",X"CA",X"E0",X"F0",X"F8",X"FC",
		X"3F",X"1F",X"07",X"07",X"03",X"01",X"02",X"00",X"FE",X"FC",X"F0",X"F0",X"E0",X"C0",X"20",X"00",
		X"00",X"10",X"28",X"29",X"03",X"07",X"0F",X"1F",X"00",X"00",X"80",X"C4",X"EA",X"F2",X"F8",X"FC",
		X"1F",X"1F",X"07",X"07",X"03",X"01",X"02",X"00",X"FE",X"FC",X"F0",X"F0",X"E0",X"C0",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"01",X"01",X"00",X"01",X"03",X"0F",X"00",X"00",X"00",X"80",X"80",X"80",X"C0",X"D8",
		X"1B",X"03",X"01",X"01",X"01",X"00",X"00",X"00",X"F0",X"C0",X"80",X"00",X"80",X"80",X"00",X"00",
		X"00",X"00",X"01",X"01",X"00",X"03",X"03",X"0F",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"D8",
		X"1B",X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"F0",X"C0",X"C0",X"00",X"80",X"80",X"00",X"00",
		X"00",X"00",X"00",X"01",X"04",X"07",X"03",X"0F",X"00",X"00",X"00",X"80",X"A0",X"E0",X"C0",X"D0",
		X"0B",X"03",X"07",X"05",X"01",X"00",X"00",X"00",X"F0",X"C0",X"E0",X"20",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"0C",X"07",X"03",X"07",X"00",X"00",X"00",X"10",X"B0",X"E0",X"C0",X"C0",
		X"03",X"03",X"07",X"0D",X"08",X"00",X"00",X"00",X"E0",X"C0",X"E0",X"30",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"0C",X"07",X"03",X"03",X"00",X"00",X"00",X"10",X"30",X"E0",X"C0",X"C0",
		X"03",X"03",X"07",X"0C",X"08",X"00",X"00",X"00",X"C0",X"C0",X"E0",X"30",X"10",X"00",X"00",X"00",
		X"00",X"00",X"03",X"07",X"0E",X"0F",X"1E",X"19",X"00",X"00",X"C0",X"E0",X"70",X"F0",X"38",X"98",
		X"11",X"18",X"0C",X"0E",X"07",X"03",X"00",X"00",X"88",X"18",X"30",X"70",X"E0",X"C0",X"00",X"00",
		X"00",X"00",X"03",X"07",X"0E",X"0C",X"18",X"18",X"00",X"00",X"C0",X"E0",X"70",X"30",X"18",X"98",
		X"19",X"18",X"0C",X"0E",X"07",X"03",X"00",X"00",X"98",X"18",X"30",X"70",X"E0",X"C0",X"00",X"00",
		X"00",X"00",X"1F",X"3F",X"3F",X"3F",X"3F",X"3F",X"00",X"00",X"F8",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",X"00",X"00",X"FC",X"FC",X"FC",X"FC",X"FC",X"F8",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"0B",X"1F",X"9F",X"00",X"00",X"00",X"E0",X"F0",X"F8",X"FC",X"FA",
		X"5F",X"3F",X"1F",X"0F",X"07",X"00",X"00",X"00",X"F9",X"F8",X"D0",X"C0",X"80",X"00",X"00",X"00",
		X"00",X"00",X"01",X"03",X"07",X"07",X"07",X"1F",X"00",X"00",X"FC",X"F0",X"E0",X"E0",X"F0",X"F8",
		X"1F",X"0F",X"07",X"07",X"0F",X"3F",X"00",X"00",X"F8",X"E0",X"E0",X"E0",X"C0",X"80",X"00",X"00",
		X"00",X"01",X"02",X"07",X"0F",X"1F",X"1F",X"1F",X"00",X"00",X"00",X"C0",X"E0",X"C0",X"F8",X"F8",
		X"1F",X"1F",X"03",X"07",X"03",X"00",X"00",X"01",X"F8",X"F8",X"F8",X"F0",X"E0",X"40",X"80",X"00",
		X"00",X"00",X"20",X"21",X"33",X"3F",X"3F",X"3F",X"00",X"00",X"00",X"80",X"80",X"E0",X"F0",X"F8",
		X"1F",X"0F",X"07",X"01",X"01",X"00",X"00",X"00",X"FC",X"FC",X"FC",X"CC",X"84",X"04",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"07",X"2E",X"1C",X"00",X"00",X"98",X"C4",X"E8",X"70",X"38",X"1C",
		X"18",X"1C",X"2E",X"07",X"03",X"01",X"00",X"00",X"0E",X"1C",X"38",X"70",X"E6",X"C1",X"86",X"00",
		X"00",X"00",X"00",X"01",X"03",X"07",X"2E",X"1C",X"00",X"00",X"86",X"C1",X"E6",X"70",X"38",X"1C",
		X"18",X"1C",X"2E",X"07",X"03",X"01",X"00",X"00",X"0E",X"1C",X"38",X"70",X"E8",X"C4",X"98",X"00",
		X"00",X"00",X"00",X"11",X"2B",X"27",X"0E",X"1C",X"00",X"04",X"8A",X"CA",X"E0",X"70",X"38",X"1C",
		X"38",X"1C",X"06",X"07",X"03",X"01",X"02",X"00",X"06",X"0C",X"10",X"30",X"60",X"C0",X"20",X"00",
		X"00",X"10",X"28",X"29",X"03",X"07",X"0E",X"1C",X"00",X"00",X"80",X"C4",X"EA",X"72",X"38",X"1C",
		X"38",X"1C",X"06",X"07",X"03",X"01",X"02",X"00",X"0E",X"1C",X"30",X"70",X"E0",X"C0",X"20",X"00",
		X"00",X"01",X"02",X"04",X"08",X"10",X"20",X"40",X"00",X"00",X"80",X"40",X"20",X"10",X"08",X"04",
		X"80",X"40",X"20",X"10",X"08",X"04",X"02",X"01",X"02",X"04",X"08",X"10",X"20",X"40",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"80",
		X"01",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"80",
		X"01",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"80",
		X"01",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"80",
		X"01",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"3E",X"41",X"41",X"41",X"41",X"41",X"3E",X"00",X"00",X"00",X"7F",X"20",X"10",X"00",X"00",
		X"00",X"31",X"49",X"49",X"49",X"49",X"49",X"27",X"00",X"46",X"69",X"59",X"49",X"41",X"41",X"41",
		X"00",X"04",X"7F",X"44",X"44",X"24",X"14",X"0C",X"00",X"46",X"49",X"49",X"49",X"49",X"49",X"79",
		X"00",X"46",X"49",X"49",X"49",X"49",X"49",X"3E",X"00",X"60",X"50",X"48",X"47",X"40",X"40",X"40",
		X"00",X"36",X"49",X"49",X"49",X"49",X"49",X"36",X"00",X"3E",X"49",X"49",X"49",X"49",X"49",X"31",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"48",X"48",X"48",X"48",X"48",X"3F",
		X"00",X"36",X"49",X"49",X"49",X"49",X"49",X"7F",X"00",X"41",X"41",X"41",X"41",X"41",X"41",X"3E",
		X"00",X"3E",X"41",X"41",X"41",X"41",X"41",X"7F",X"00",X"41",X"41",X"49",X"49",X"49",X"49",X"7F",
		X"00",X"40",X"40",X"48",X"48",X"48",X"48",X"7F",X"00",X"4F",X"49",X"49",X"41",X"41",X"41",X"3E",
		X"00",X"7F",X"08",X"08",X"08",X"08",X"08",X"7F",X"00",X"00",X"00",X"00",X"7F",X"00",X"00",X"00",
		X"00",X"7E",X"01",X"01",X"01",X"01",X"01",X"06",X"00",X"41",X"22",X"14",X"08",X"04",X"02",X"7F",
		X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"7F",X"00",X"7F",X"20",X"10",X"08",X"10",X"20",X"7F",
		X"00",X"7F",X"02",X"04",X"08",X"10",X"20",X"7F",X"00",X"3E",X"41",X"41",X"41",X"41",X"41",X"3E",
		X"00",X"30",X"48",X"48",X"48",X"48",X"48",X"7F",X"00",X"3D",X"42",X"45",X"41",X"41",X"41",X"3E",
		X"00",X"31",X"4A",X"4C",X"48",X"48",X"48",X"7F",X"00",X"46",X"49",X"49",X"49",X"49",X"49",X"31",
		X"00",X"40",X"40",X"40",X"7F",X"40",X"40",X"40",X"00",X"7E",X"01",X"01",X"01",X"01",X"01",X"7E",
		X"00",X"78",X"04",X"02",X"01",X"02",X"04",X"78",X"00",X"7C",X"02",X"01",X"06",X"01",X"02",X"7C",
		X"00",X"41",X"22",X"14",X"08",X"14",X"22",X"41",X"00",X"40",X"20",X"10",X"0F",X"10",X"20",X"40",
		X"00",X"41",X"61",X"51",X"49",X"45",X"43",X"41",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"60",X"10",X"00",X"00",X"00",X"00",X"00",X"60",X"10",X"00",X"60",X"10",
		X"00",X"10",X"60",X"00",X"10",X"60",X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"08",X"08",X"00",
		X"00",X"40",X"20",X"10",X"08",X"04",X"02",X"01",X"00",X"08",X"08",X"08",X"7F",X"08",X"08",X"08",
		X"00",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"00",X"08",X"08",X"08",X"2A",X"08",X"08",X"08",
		X"00",X"00",X"7D",X"00",X"00",X"7D",X"00",X"00",X"7E",X"C3",X"A5",X"A5",X"A5",X"BD",X"C3",X"7E",
		X"F6",X"F6",X"00",X"00",X"F6",X"F6",X"00",X"00",X"FA",X"FA",X"00",X"00",X"FA",X"FA",X"00",X"00",
		X"00",X"00",X"00",X"F6",X"F6",X"00",X"00",X"00",X"00",X"00",X"00",X"FA",X"FA",X"00",X"00",X"00",
		X"00",X"00",X"00",X"E0",X"C0",X"00",X"00",X"00",X"00",X"E0",X"C0",X"00",X"E0",X"C0",X"00",X"00",
		X"00",X"60",X"E0",X"00",X"60",X"E0",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"C0",X"80",X"C0",X"80",X"C0",X"80",X"C0",X"80",X"03",X"01",X"03",X"01",X"03",X"01",X"03",X"01",
		X"E0",X"C0",X"E0",X"C0",X"E0",X"C0",X"E0",X"C0",X"07",X"03",X"07",X"03",X"07",X"03",X"07",X"03",
		X"F0",X"E0",X"F0",X"E0",X"F0",X"E0",X"F0",X"E0",X"0F",X"07",X"0F",X"07",X"0F",X"07",X"0F",X"07",
		X"F8",X"F0",X"F8",X"F0",X"F8",X"F0",X"F8",X"F0",X"1F",X"0F",X"1F",X"0F",X"1F",X"0F",X"1F",X"0F",
		X"FC",X"F8",X"FC",X"F8",X"FC",X"F8",X"FC",X"F8",X"3F",X"1F",X"3F",X"1F",X"3F",X"1F",X"3F",X"1F",
		X"FE",X"FC",X"FE",X"FC",X"FE",X"FC",X"FE",X"FC",X"7F",X"3F",X"7F",X"3F",X"7F",X"3F",X"7F",X"3F",
		X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"7F",X"FF",X"7F",X"FF",X"7F",X"FF",X"7F",
		X"00",X"10",X"38",X"10",X"00",X"40",X"02",X"07",X"3F",X"3F",X"3F",X"07",X"0F",X"1F",X"07",X"0F",
		X"02",X"20",X"70",X"21",X"00",X"04",X"0E",X"04",X"07",X"03",X"00",X"06",X"03",X"07",X"1F",X"0F",
		X"00",X"00",X"00",X"10",X"38",X"10",X"00",X"40",X"3F",X"3F",X"3F",X"07",X"0F",X"0F",X"03",X"0F",
		X"04",X"04",X"00",X"20",X"70",X"21",X"00",X"80",X"07",X"03",X"00",X"06",X"03",X"07",X"1F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"3F",X"3F",X"07",X"0F",X"0F",X"03",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"03",X"00",X"06",X"03",X"07",X"1F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"3F",X"3F",X"07",X"0F",X"0F",X"0F",X"8F",
		X"01",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"8F",X"FF",X"FF",X"EF",X"FF",X"0F",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0C",X"00",X"00",X"00",X"18",X"3C",X"3C",X"3C",X"3F",
		X"07",X"07",X"06",X"07",X"00",X"00",X"00",X"00",X"FF",X"FF",X"7F",X"7E",X"7C",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"60",X"00",X"00",X"00",X"00",X"18",X"3C",X"7C",X"FC",
		X"2B",X"2B",X"79",X"3E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"C1",X"00",X"00",X"00",X"00",X"38",X"78",X"F8",X"F0",
		X"E9",X"FB",X"F3",X"7D",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F8",X"F8",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"F8",X"F8",X"E0",X"C0",X"80",
		X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"18",X"3C",X"7E",X"FF",
		X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",
		X"FF",X"7E",X"3C",X"18",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",
		X"01",X"03",X"07",X"1F",X"1F",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"71",X"89",X"89",X"89",X"89",X"89",X"67",X"00",X"6E",X"91",X"91",X"91",X"91",X"91",X"6E",X"00",
		X"7E",X"91",X"91",X"91",X"91",X"91",X"61",X"00",X"FF",X"40",X"20",X"00",X"00",X"00",X"00",X"00",
		X"7E",X"C3",X"A5",X"A5",X"A5",X"BD",X"C3",X"7E",X"00",X"40",X"40",X"40",X"7F",X"40",X"40",X"40",
		X"00",X"7F",X"02",X"04",X"08",X"10",X"20",X"7F",X"00",X"46",X"49",X"49",X"49",X"49",X"49",X"31",
		X"00",X"41",X"41",X"49",X"49",X"49",X"49",X"7F",X"00",X"31",X"4A",X"4C",X"48",X"48",X"48",X"7F",
		X"00",X"30",X"48",X"48",X"48",X"48",X"48",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"8F",X"2F",X"EF",X"EF",X"EF",X"EF",X"8F",X"3F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"3F",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"F8",X"E3",
		X"8F",X"3F",X"FF",X"FF",X"FF",X"E7",X"87",X"37",X"77",X"77",X"37",X"87",X"E7",X"FF",X"FF",X"FF",
		X"FF",X"FE",X"F8",X"F3",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F3",X"F8",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"EF",X"EF",X"EF",X"2F",X"0F",X"7F",X"7F",
		X"3F",X"8F",X"E7",X"F7",X"F7",X"F7",X"F7",X"F7",X"0F",X"EF",X"EF",X"EF",X"CF",X"DF",X"DF",X"9F",
		X"87",X"BF",X"BF",X"BF",X"9F",X"DF",X"DF",X"CF",X"BF",X"BF",X"3F",X"7F",X"7F",X"0F",X"0F",X"EF",
		X"EF",X"EF",X"E7",X"F7",X"F7",X"F7",X"87",X"BF",X"EF",X"0F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"1F",X"CF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"8F",X"1F",X"7F",X"FF",
		X"BF",X"87",X"F7",X"77",X"17",X"C7",X"F7",X"FF",X"FF",X"7F",X"1F",X"C7",X"F1",X"FC",X"FE",X"FE",
		X"FC",X"F1",X"C7",X"1F",X"7F",X"FF",X"FC",X"F9",X"C7",X"1F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"F1",X"F4",X"F7",X"F7",X"F7",X"F7",X"F1",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FC",X"F1",X"F7",X"F7",X"F7",X"F7",X"F4",X"F1",X"FF",X"FF",X"FF",X"FF",
		X"EF",X"EF",X"E7",X"F7",X"F7",X"F7",X"87",X"BF",X"EF",X"0F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"1F",X"CF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"8F",X"1F",X"7F",X"FF",
		X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"00",X"F8",X"04",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"04",X"F8",X"00",
		X"00",X"1F",X"20",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"20",X"1F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"02",X"02",X"02",X"01",X"01",X"01",
		X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"02",X"02",X"02",X"04",X"04",X"04",X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"02",
		X"82",X"42",X"22",X"19",X"05",X"03",X"01",X"00",X"04",X"04",X"04",X"04",X"04",X"04",X"02",X"02",
		X"09",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"04",X"02",X"01",X"04",X"0A",
		X"04",X"04",X"04",X"08",X"08",X"08",X"08",X"08",X"03",X"1C",X"20",X"40",X"81",X"01",X"02",X"02",
		X"08",X"04",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"48",X"26",X"21",X"10",X"08",
		X"10",X"88",X"44",X"22",X"11",X"08",X"04",X"02",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"20",
		X"F8",X"07",X"00",X"F0",X"0C",X"02",X"01",X"00",X"20",X"10",X"08",X"07",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"30",X"4C",X"42",X"21",X"10",X"08",X"04",X"02",X"01",X"00",X"00",X"00",
		X"20",X"10",X"0C",X"02",X"81",X"40",X"40",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",
		X"42",X"21",X"21",X"11",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"78",X"44",
		X"60",X"98",X"84",X"42",X"41",X"23",X"1D",X"00",X"10",X"08",X"08",X"07",X"00",X"00",X"00",X"00",
		X"00",X"80",X"40",X"40",X"20",X"20",X"20",X"10",X"44",X"44",X"44",X"44",X"C4",X"24",X"24",X"18",
		X"08",X"08",X"04",X"04",X"04",X"04",X"04",X"04",X"42",X"42",X"21",X"21",X"10",X"10",X"08",X"08",
		X"10",X"08",X"C4",X"22",X"11",X"08",X"04",X"84",X"00",X"80",X"B8",X"24",X"22",X"21",X"20",X"10",
		X"08",X"08",X"04",X"02",X"02",X"01",X"00",X"00",X"81",X"80",X"40",X"40",X"40",X"21",X"20",X"10",
		X"08",X"04",X"03",X"00",X"00",X"70",X"8C",X"82",X"10",X"08",X"04",X"02",X"01",X"80",X"40",X"20",
		X"12",X"12",X"0A",X"09",X"05",X"84",X"42",X"21",X"00",X"00",X"00",X"0F",X"10",X"20",X"20",X"21",
		X"20",X"10",X"08",X"04",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"30",X"28",X"26",X"21",X"20",
		X"09",X"08",X"08",X"04",X"02",X"01",X"00",X"00",X"04",X"02",X"01",X"00",X"00",X"00",X"0C",X"0A",
		X"12",X"21",X"20",X"20",X"10",X"10",X"08",X"04",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",
		X"23",X"50",X"88",X"06",X"01",X"00",X"00",X"00",X"20",X"20",X"20",X"20",X"20",X"10",X"08",X"04",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"40",X"40",X"20",X"20",X"20",X"20",X"20",X"20",
		X"07",X"00",X"00",X"00",X"80",X"80",X"40",X"40",X"20",X"10",X"08",X"04",X"03",X"80",X"60",X"18",
		X"10",X"0F",X"00",X"00",X"00",X"00",X"80",X"40",X"40",X"20",X"10",X"10",X"08",X"07",X"80",X"60",
		X"80",X"80",X"40",X"40",X"C0",X"00",X"80",X"80",X"12",X"09",X"06",X"C0",X"30",X"0E",X"01",X"01",
		X"A1",X"92",X"4A",X"24",X"10",X"90",X"48",X"24",X"88",X"48",X"24",X"14",X"0A",X"85",X"42",X"42",
		X"18",X"04",X"02",X"01",X"80",X"40",X"20",X"10",X"40",X"20",X"20",X"10",X"0F",X"00",X"80",X"60",
		X"18",X"06",X"01",X"01",X"00",X"00",X"00",X"80",X"88",X"44",X"22",X"11",X"09",X"06",X"C0",X"20",
		X"90",X"48",X"24",X"93",X"88",X"44",X"22",X"11",X"01",X"01",X"80",X"40",X"20",X"10",X"0C",X"E3",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"06",X"03",X"60",X"10",X"08",X"04",X"02",X"C2",X"31",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"22",X"42",X"82",X"02",X"02",X"04",X"38",X"20",X"40",X"A0",X"90",X"48",X"44",X"44",X"24",
		X"22",X"22",X"22",X"22",X"42",X"84",X"04",X"18",X"A0",X"90",X"48",X"48",X"44",X"24",X"24",X"22",
		X"20",X"10",X"08",X"04",X"02",X"7C",X"80",X"40",X"02",X"04",X"08",X"10",X"60",X"80",X"80",X"40",
		X"24",X"14",X"12",X"12",X"11",X"21",X"21",X"C1",X"70",X"80",X"80",X"40",X"A0",X"A0",X"50",X"28",
		X"44",X"44",X"42",X"82",X"02",X"04",X"04",X"08",X"38",X"40",X"40",X"40",X"A0",X"90",X"50",X"48",
		X"80",X"40",X"20",X"10",X"08",X"04",X"04",X"0C",X"02",X"02",X"02",X"02",X"C4",X"38",X"00",X"00",
		X"80",X"40",X"A0",X"90",X"50",X"48",X"44",X"84",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"10",X"08",X"04",X"02",X"C2",X"31",X"0E",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"FF",X"7F",X"3F",X"1F",X"0F",X"07",X"03",X"01",
		X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"AA",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"AA",
		X"55",X"83",X"07",X"8F",X"1F",X"BF",X"7F",X"FF",X"FF",X"FC",X"F9",X"F0",X"E1",X"C0",X"81",X"00",
		X"FF",X"FF",X"3F",X"9F",X"0F",X"87",X"03",X"AB",X"01",X"80",X"C1",X"E0",X"F1",X"F8",X"FD",X"FE",
		X"55",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"55",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"AA",X"01",X"03",X"07",X"0F",X"1F",X"3F",X"7F",X"FF",
		X"55",X"80",X"C0",X"E0",X"F0",X"F8",X"FC",X"FE",X"55",X"01",X"03",X"07",X"0F",X"1F",X"3F",X"7F",
		X"FF",X"FF",X"3F",X"9F",X"0F",X"87",X"03",X"AB",X"FF",X"FE",X"FD",X"F8",X"F1",X"E0",X"C1",X"AA",
		X"55",X"83",X"07",X"8F",X"1F",X"BF",X"7F",X"FF",X"D5",X"C0",X"E1",X"F0",X"F9",X"FC",X"FF",X"FF",
		X"FF",X"FF",X"3F",X"9F",X"0F",X"87",X"03",X"AB",X"FF",X"FE",X"FD",X"F8",X"F1",X"E0",X"C1",X"AA",
		X"55",X"83",X"07",X"8F",X"1F",X"BF",X"7F",X"FF",X"D5",X"C0",X"E1",X"F0",X"F9",X"FC",X"FF",X"FF",
		X"FE",X"FC",X"F8",X"F0",X"E0",X"C0",X"80",X"AA",X"7F",X"3F",X"1F",X"0F",X"07",X"03",X"AA",X"FF",
		X"FF",X"FE",X"FC",X"F8",X"F0",X"E0",X"C0",X"80",X"55",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"AA",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"AA",
		X"7F",X"BF",X"1F",X"8F",X"07",X"83",X"01",X"80",X"D5",X"C0",X"E1",X"F0",X"F9",X"FC",X"FF",X"FF",
		X"00",X"81",X"03",X"87",X"0F",X"9F",X"3F",X"FF",X"FF",X"FE",X"FB",X"F8",X"F1",X"E0",X"C1",X"AA",
		X"55",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"55",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"80",X"C0",X"E0",X"F0",X"F8",X"FC",X"FE",X"FF",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"19",X"06",X"05",X"2A",X"15",X"00",X"00",X"80",X"58",X"B0",X"50",X"A8",X"54",
		X"0A",X"15",X"2A",X"05",X"06",X"09",X"00",X"00",X"AA",X"54",X"A8",X"50",X"B0",X"4E",X"80",X"00",
		X"00",X"00",X"00",X"09",X"06",X"05",X"2A",X"15",X"00",X"00",X"80",X"4E",X"B0",X"50",X"A8",X"54",
		X"0A",X"15",X"2A",X"05",X"06",X"19",X"00",X"00",X"AA",X"54",X"A8",X"50",X"B0",X"58",X"80",X"00",
		X"00",X"00",X"00",X"01",X"12",X"1D",X"0A",X"15",X"00",X"00",X"84",X"44",X"A4",X"58",X"A8",X"54",
		X"2A",X"15",X"0A",X"15",X"12",X"01",X"02",X"00",X"AA",X"54",X"A8",X"54",X"A0",X"40",X"20",X"00",
		X"00",X"00",X"10",X"11",X"12",X"0D",X"0A",X"15",X"00",X"00",X"80",X"40",X"A4",X"5C",X"A8",X"54",
		X"2A",X"15",X"0A",X"15",X"02",X"01",X"02",X"00",X"A8",X"54",X"A8",X"54",X"A4",X"40",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"04",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"20",
		X"04",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"20",X"40",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"07",X"08",X"11",X"12",X"14",X"00",X"00",X"00",X"E0",X"10",X"88",X"48",X"28",
		X"14",X"12",X"11",X"08",X"07",X"00",X"00",X"00",X"28",X"48",X"88",X"10",X"E0",X"00",X"00",X"00",
		X"00",X"1F",X"20",X"47",X"48",X"51",X"52",X"54",X"00",X"F8",X"04",X"E2",X"12",X"8A",X"4A",X"2A",
		X"54",X"52",X"51",X"48",X"47",X"20",X"1F",X"00",X"2A",X"4A",X"8A",X"12",X"E2",X"04",X"F8",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"01",X"00",X"00",X"00",X"00",X"03",X"21",X"00",X"80",X"00",X"00",X"00",X"00",X"C0",X"84",
		X"21",X"03",X"00",X"00",X"00",X"00",X"01",X"00",X"84",X"C0",X"00",X"00",X"00",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"40",X"C0",X"80",
		X"01",X"03",X"02",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"06",X"03",X"01",X"00",X"00",X"00",X"00",X"20",X"60",X"C0",X"80",
		X"01",X"03",X"06",X"04",X"00",X"00",X"00",X"00",X"80",X"C0",X"60",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"0C",X"06",X"03",X"01",X"00",X"00",X"00",X"10",X"30",X"60",X"C0",X"80",
		X"01",X"03",X"06",X"0C",X"08",X"00",X"00",X"00",X"80",X"C0",X"60",X"30",X"10",X"00",X"00",X"00",
		X"00",X"00",X"18",X"08",X"0C",X"06",X"03",X"01",X"00",X"00",X"18",X"10",X"30",X"60",X"C0",X"80",
		X"01",X"03",X"06",X"0C",X"08",X"18",X"00",X"00",X"80",X"C0",X"60",X"30",X"10",X"18",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"0F",X"00",X"00",X"00",X"00",X"80",X"C0",X"70",X"F0",
		X"0F",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"07",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"E0",
		X"07",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"E0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"1F",X"20",X"40",X"40",X"40",X"40",X"40",X"00",X"F8",X"04",X"02",X"02",X"02",X"02",X"02",
		X"40",X"40",X"40",X"40",X"40",X"20",X"1F",X"00",X"02",X"02",X"02",X"02",X"02",X"04",X"F8",X"00",
		X"00",X"00",X"00",X"00",X"04",X"07",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"F0",
		X"0F",X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"E0",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"1F",X"0F",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"F0",
		X"0F",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"F0",X"F8",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"07",X"00",X"00",X"00",X"00",X"C0",X"F0",X"F0",X"F0",
		X"0F",X"0F",X"0F",X"03",X"00",X"00",X"00",X"00",X"E0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"03",X"07",X"07",X"00",X"00",X"00",X"40",X"E0",X"C0",X"E0",X"E0",
		X"07",X"07",X"03",X"07",X"02",X"00",X"00",X"00",X"E0",X"E0",X"C0",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"19",X"06",X"05",X"2A",X"14",X"00",X"00",X"80",X"58",X"B0",X"50",X"28",X"14",
		X"08",X"14",X"2A",X"05",X"06",X"09",X"00",X"00",X"0A",X"14",X"28",X"50",X"B0",X"4E",X"80",X"00",
		X"00",X"00",X"00",X"09",X"06",X"05",X"2A",X"14",X"00",X"00",X"80",X"4E",X"B0",X"50",X"28",X"14",
		X"08",X"14",X"2A",X"05",X"06",X"19",X"00",X"00",X"0A",X"14",X"28",X"50",X"B0",X"58",X"80",X"00",
		X"00",X"00",X"00",X"01",X"12",X"1D",X"0A",X"14",X"00",X"00",X"84",X"44",X"A4",X"58",X"28",X"14",
		X"28",X"14",X"0A",X"15",X"12",X"01",X"02",X"00",X"0A",X"14",X"28",X"54",X"A0",X"40",X"20",X"00",
		X"00",X"00",X"10",X"11",X"12",X"0D",X"0A",X"14",X"00",X"00",X"80",X"40",X"A4",X"5C",X"28",X"14",
		X"28",X"14",X"0A",X"15",X"02",X"01",X"02",X"00",X"0A",X"14",X"28",X"54",X"A4",X"40",X"20",X"00",
		X"00",X"00",X"01",X"02",X"04",X"08",X"10",X"20",X"00",X"00",X"00",X"80",X"40",X"20",X"10",X"08",
		X"40",X"20",X"10",X"08",X"04",X"02",X"01",X"00",X"04",X"08",X"10",X"20",X"40",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"1D",X"FF",X"00",X"00",X"00",X"00",X"00",X"C0",X"B8",X"FE",
		X"7F",X"1D",X"03",X"00",X"00",X"00",X"00",X"00",X"FF",X"B8",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"1F",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"F0",
		X"0F",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"F8",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"07",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"E0",
		X"07",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"E0",X"80",X"80",X"80",X"80",X"00",X"00",X"00",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"C0",
		X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"C0",X"80",X"80",X"80",X"80",X"80",X"80",X"80");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
