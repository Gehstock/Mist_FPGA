library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity fg1_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of fg1_rom is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"99",X"99",X"AA",X"AA",X"99",X"99",X"AA",X"AA",X"99",X"99",X"AA",X"AA",X"99",X"99",
		X"55",X"55",X"EE",X"EE",X"58",X"88",X"8B",X"BB",X"99",X"9B",X"97",X"78",X"99",X"AA",X"AA",X"AA",
		X"55",X"55",X"EE",X"55",X"88",X"88",X"88",X"BB",X"9B",X"BB",X"99",X"AA",X"9A",X"A9",X"99",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"11",X"11",X"11",X"21",X"21",X"12",X"12",
		X"21",X"21",X"22",X"22",X"32",X"32",X"23",X"23",X"32",X"32",X"33",X"33",X"43",X"43",X"34",X"34",
		X"43",X"43",X"34",X"34",X"54",X"54",X"45",X"45",X"54",X"54",X"45",X"45",X"65",X"65",X"56",X"56",
		X"65",X"65",X"56",X"56",X"76",X"76",X"67",X"67",X"76",X"76",X"67",X"67",X"87",X"87",X"78",X"78",
		X"87",X"87",X"78",X"78",X"98",X"98",X"89",X"89",X"98",X"98",X"89",X"89",X"A9",X"A9",X"9A",X"9A",
		X"A9",X"A9",X"9A",X"9A",X"BA",X"BA",X"AB",X"AB",X"BA",X"BA",X"AB",X"AB",X"CB",X"CB",X"BC",X"BC",
		X"CB",X"CB",X"BC",X"BC",X"DC",X"DC",X"CD",X"CD",X"DC",X"DC",X"CD",X"CD",X"ED",X"ED",X"DE",X"DE",
		X"ED",X"ED",X"DE",X"DE",X"FE",X"FE",X"EF",X"EF",X"FE",X"FE",X"EF",X"EF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"40",
		X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"4A",X"00",X"AA",X"00",X"DA",X"04",X"AA",X"00",X"AA",
		X"4A",X"A4",X"4A",X"AA",X"AA",X"AA",X"AA",X"AD",X"AA",X"AA",X"AD",X"AA",X"AA",X"AA",X"AA",X"AD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"44",X"00",X"4A",X"00",X"A4",X"00",X"AA",X"04",X"AA",X"44",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"41",X"00",X"11",X"40",X"11",X"44",X"11",
		X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"44",
		X"44",X"44",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"00",X"11",X"44",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"44",X"44",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"44",X"44",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"44",X"44",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"00",X"00",X"40",X"00",X"14",X"00",X"14",X"00",X"14",X"00",X"14",X"00",X"14",X"00",X"14",X"00",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"40",X"11",X"14",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"DA",X"AA",X"AA",X"AA",X"AA",X"DA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"A4",X"11",X"AA",X"33",X"AA",X"44",X"44",X"AA",X"4A",X"44",X"AA",X"33",X"A4",X"33",X"44",X"44",
		X"AA",X"DA",X"AA",X"AA",X"AA",X"A4",X"4A",X"4F",X"E4",X"A4",X"E4",X"44",X"5E",X"04",X"5E",X"04",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"44",X"44",X"00",X"DD",X"00",X"DD",X"00",X"DD",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"44",X"44",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"44",X"44",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"44",X"44",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"44",X"44",X"DD",X"DD",X"DD",X"4D",X"DD",X"4D",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"44",X"44",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"44",X"44",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"44",X"44",X"DD",X"D4",X"DD",X"D4",X"DD",X"D4",
		X"FF",X"5E",X"FF",X"5E",X"FF",X"5E",X"FF",X"E5",X"44",X"E5",X"34",X"E5",X"34",X"56",X"34",X"56",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"44",X"44",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"44",X"44",
		X"66",X"88",X"66",X"57",X"66",X"58",X"66",X"55",X"66",X"22",X"66",X"99",X"66",X"BB",X"65",X"99",
		X"88",X"88",X"77",X"77",X"58",X"88",X"35",X"55",X"32",X"22",X"39",X"99",X"39",X"BB",X"39",X"99",
		X"5E",X"04",X"65",X"04",X"65",X"04",X"65",X"04",X"66",X"44",X"66",X"44",X"66",X"44",X"44",X"E4",
		X"00",X"DD",X"00",X"DD",X"00",X"54",X"00",X"C4",X"00",X"C4",X"00",X"C4",X"00",X"C4",X"00",X"C4",
		X"00",X"E4",X"00",X"E4",X"00",X"4E",X"00",X"4E",X"00",X"4E",X"00",X"4C",X"00",X"4C",X"00",X"4C",
		X"00",X"C4",X"00",X"C4",X"00",X"C4",X"04",X"44",X"49",X"99",X"04",X"BB",X"00",X"55",X"00",X"54",
		X"DD",X"DD",X"DD",X"DD",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"DD",X"4D",X"DD",X"4D",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"64",X"44",X"76",X"48",X"88",X"99",X"99",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"43",X"44",X"43",X"44",X"99",X"99",X"44",X"44",X"44",X"44",X"44",X"44",
		X"DD",X"D4",X"DD",X"D4",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"3C",X"56",X"35",X"66",X"35",X"66",X"35",X"66",X"5E",X"66",X"5E",X"66",X"5E",X"66",X"E5",X"66",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"99",X"99",X"BB",X"44",X"44",X"44",X"44",X"44",
		X"E5",X"55",X"E5",X"B9",X"55",X"B9",X"55",X"B9",X"55",X"B9",X"35",X"22",X"35",X"55",X"35",X"88",
		X"65",X"9B",X"53",X"9B",X"53",X"9B",X"B3",X"9B",X"B3",X"9B",X"B3",X"9B",X"B3",X"9B",X"B3",X"9B",
		X"39",X"B9",X"39",X"B9",X"39",X"B9",X"39",X"B9",X"39",X"B9",X"39",X"B9",X"39",X"B9",X"39",X"B9",
		X"B3",X"9B",X"B3",X"9B",X"B3",X"9B",X"B3",X"9B",X"B3",X"9B",X"23",X"22",X"53",X"55",X"53",X"88",
		X"39",X"B9",X"39",X"B9",X"39",X"B9",X"39",X"B9",X"39",X"B9",X"32",X"22",X"35",X"55",X"35",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"09",X"00",X"9D",X"00",X"9D",
		X"00",X"00",X"00",X"00",X"99",X"99",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"00",X"9D",X"00",X"9D",X"00",X"9D",X"00",X"9D",X"00",X"09",X"00",X"09",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"90",
		X"DD",X"90",X"DD",X"90",X"DD",X"90",X"DD",X"90",X"DD",X"90",X"DD",X"90",X"DD",X"90",X"DD",X"90",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"99",X"99",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"99",X"DD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"BB",X"09",X"BB",X"9B",X"BB",X"9B",X"BB",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"D9",X"99",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"9B",X"BB",X"9B",X"BB",X"9B",X"BB",X"09",X"BB",X"09",X"BB",X"00",X"BB",X"00",X"9B",X"00",X"09",
		X"00",X"DD",X"00",X"DD",X"00",X"DD",X"99",X"DD",X"BB",X"99",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"99",X"DD",X"BB",X"99",X"BB",X"BB",
		X"90",X"00",X"90",X"00",X"90",X"00",X"90",X"00",X"90",X"00",X"90",X"00",X"90",X"00",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"99",X"00",X"BB",X"99",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"B9",X"09",X"B9",X"09",X"B9",X"09",X"B9",X"9D",
		X"DD",X"90",X"DD",X"90",X"DD",X"90",X"DD",X"90",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",
		X"00",X"00",X"00",X"09",X"00",X"9D",X"00",X"9D",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",
		X"99",X"99",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"99",X"BB",X"9D",X"9B",X"9D",X"D9",X"D9",X"DD",X"D9",X"DD",X"D9",X"DD",X"D9",X"DD",X"D9",X"99",
		X"BB",X"BB",X"BB",X"BB",X"99",X"BB",X"DD",X"99",X"DD",X"90",X"DD",X"00",X"99",X"99",X"DD",X"DD",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"99",X"99",X"00",X"00",X"09",X"00",X"09",X"90",X"09",
		X"B9",X"9D",X"90",X"DD",X"99",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"D9",X"00",X"D9",X"00",X"9D",X"90",
		X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",
		X"D9",X"DD",X"D9",X"DD",X"D9",X"DD",X"D9",X"DD",X"D9",X"DD",X"D9",X"DD",X"D9",X"DD",X"D9",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"D9",X"DD",X"9B",X"DD",X"9B",X"DD",X"9B",
		X"90",X"00",X"90",X"00",X"99",X"00",X"BB",X"99",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"DD",X"DD",X"DD",X"DD",X"99",X"DD",X"BB",X"99",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"9B",X"BB",
		X"DD",X"D9",X"DD",X"9D",X"99",X"DD",X"DD",X"DD",X"9D",X"DD",X"99",X"DD",X"B9",X"DD",X"BB",X"DD",
		X"DD",X"D9",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"09",X"DD",X"09",X"DD",X"09",X"DD",X"09",X"DD",
		X"D9",X"DD",X"D9",X"DD",X"D9",X"DD",X"90",X"DD",X"90",X"DD",X"90",X"DD",X"90",X"DD",X"90",X"DD",
		X"DD",X"9B",X"DD",X"9B",X"DD",X"9B",X"DD",X"D9",X"DD",X"D9",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"9B",X"BB",X"D9",X"BB",
		X"9B",X"BB",X"B9",X"BB",X"B9",X"BB",X"B9",X"BB",X"B9",X"BB",X"9B",X"BB",X"99",X"BB",X"DD",X"BB",
		X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",X"B9",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"09",X"DD",X"09",X"DD",X"09",X"DD",X"09",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"9D",X"00",X"09",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"99",X"99",X"00",
		X"90",X"DD",X"90",X"DD",X"90",X"DD",X"00",X"9D",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"99",X"DD",X"00",X"99",
		X"DD",X"99",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"99",X"99",
		X"DD",X"99",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"99",X"99",
		X"9D",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"99",X"99",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"D9",X"DD",X"90",X"DD",X"00",X"99",X"00",
		X"00",X"99",X"09",X"DD",X"09",X"DD",X"9D",X"DD",X"9D",X"DD",X"9D",X"DD",X"9D",X"DD",X"9D",X"DD",
		X"99",X"90",X"DD",X"D9",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"99",X"09",X"DD",X"9D",X"DD",X"9D",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"00",X"00",X"99",X"99",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"9D",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"D9",X"DD",X"9B",
		X"00",X"00",X"99",X"99",X"DD",X"D9",X"DD",X"9B",X"D9",X"BB",X"9B",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"00",X"00",X"99",X"99",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"B9",X"00",X"B9",X"00",X"BB",X"00",X"BB",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"9D",X"DD",X"9D",X"DD",X"09",X"DD",X"00",X"99",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"D9",X"99",X"9B",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"D9",X"DD",X"9B",X"D9",X"BB",X"9B",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"D9",X"BB",X"9B",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"B9",X"BB",X"90",X"B9",X"00",X"90",X"00",
		X"BB",X"00",X"B9",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"9D",X"00",X"DD",X"00",X"DD",X"09",X"DD",X"09",X"DD",X"09",X"D9",X"09",X"9B",
		X"99",X"99",X"DD",X"DD",X"DD",X"D9",X"DD",X"9B",X"D9",X"BB",X"9B",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"99",X"BB",X"9B",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"B9",X"BB",X"9D",X"B9",X"DD",X"9D",X"DD",
		X"BB",X"B9",X"BB",X"9D",X"B9",X"DD",X"9D",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"99",X"99",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"99",X"00",X"DD",X"90",X"DD",X"D9",X"DD",X"D9",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"09",X"BB",X"09",X"BB",X"09",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"B9",X"BB",X"9D",X"B9",X"DD",X"99",X"99",
		X"BB",X"B9",X"BB",X"9D",X"B9",X"DD",X"9D",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"99",X"99",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"99",X"99",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"D9",X"DD",X"D9",X"DD",X"90",X"99",X"00",
		X"00",X"9B",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"09",X"00",X"9D",X"00",X"9D",X"00",X"9D",
		X"BB",X"B9",X"BB",X"9D",X"99",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"D9",X"DD",X"9B",X"DD",X"BB",X"D9",X"BB",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"99",X"DD",X"BB",X"9D",X"BB",X"B9",X"BB",X"BB",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"90",X"00",X"D9",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",
		X"00",X"9D",X"00",X"9D",X"00",X"9D",X"00",X"9D",X"00",X"9D",X"00",X"9D",X"00",X"9D",X"00",X"9D",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"D9",X"99",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"9B",X"BB",X"9B",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"9B",X"BB",X"9B",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"DD",X"DD",X"DD",X"DD",X"9D",X"DD",X"9D",X"DD",X"99",X"99",X"9D",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",
		X"00",X"9D",X"00",X"9D",X"00",X"9D",X"00",X"09",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"9D",X"DD",X"09",X"99",
		X"D9",X"BB",X"DD",X"BB",X"DD",X"9B",X"DD",X"D9",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"99",X"99",
		X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"D9",X"00",X"90",X"00",X"00",X"00",
		X"00",X"9D",X"00",X"9D",X"00",X"9D",X"00",X"9D",X"00",X"9D",X"00",X"9D",X"00",X"9D",X"00",X"9D",
		X"BB",X"BB",X"BB",X"B9",X"BB",X"9D",X"99",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"99",X"99",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"99",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"DD",X"00",X"DD",X"09",X"DD",
		X"00",X"00",X"00",X"00",X"99",X"00",X"DD",X"90",X"DD",X"D9",X"DD",X"D9",X"DD",X"DD",X"DD",X"DD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"9D",X"00",X"DD",X"00",X"DD",X"00",X"DD",
		X"9D",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"D9",X"DD",X"D9",X"DD",X"90",X"DD",X"00",X"DD",X"00",
		X"00",X"DD",X"09",X"DD",X"09",X"DD",X"09",X"DD",X"09",X"DD",X"09",X"DD",X"09",X"DD",X"09",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"D9",X"00",X"90",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",
		X"09",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"9D",
		X"90",X"00",X"D9",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"90",X"DD",X"D9",X"DD",X"D9",X"DD",X"DD",
		X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DD",X"DD",X"DD",X"D9",X"DD",X"9D",X"9D",X"DD",X"09",X"DD",X"9D",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"DD",X"9D",X"DD",X"D9",X"DD",X"DD",X"DD",X"DD",X"99",X"DD",X"D9",X"DD",X"D9",X"DD",X"D9",
		X"00",X"00",X"00",X"09",X"00",X"09",X"00",X"9D",X"00",X"9D",X"00",X"DD",X"00",X"DD",X"00",X"DD",
		X"DD",X"D9",X"DD",X"D9",X"DD",X"D9",X"DD",X"90",X"DD",X"90",X"DD",X"00",X"DD",X"99",X"DD",X"DD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",
		X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"09",X"DD",X"09",X"DD",X"09",X"DD",X"09",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"D9",X"DD",X"9D",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"D9",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"90",X"DD",X"90",X"DD",X"D9",X"DD",X"D9",
		X"09",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"99",X"00",X"00",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"D9",X"DD",X"90",X"DD",X"90",X"DD",X"00",X"99",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"D9",X"DD",X"D9",X"99",X"90",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"99",X"99",
		X"98",X"99",X"88",X"88",X"88",X"98",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"98",X"88",X"88",
		X"88",X"98",X"88",X"88",X"99",X"89",X"88",X"88",X"99",X"88",X"88",X"88",X"88",X"89",X"88",X"88",
		X"88",X"89",X"88",X"88",X"88",X"89",X"88",X"88",X"88",X"98",X"89",X"88",X"89",X"88",X"88",X"89",
		X"88",X"98",X"88",X"88",X"88",X"98",X"88",X"88",X"98",X"98",X"98",X"98",X"98",X"98",X"99",X"88",
		X"98",X"00",X"98",X"00",X"98",X"09",X"98",X"98",X"98",X"88",X"88",X"88",X"98",X"98",X"98",X"98",
		X"09",X"98",X"09",X"98",X"99",X"99",X"88",X"88",X"99",X"89",X"99",X"89",X"88",X"89",X"98",X"89",
		X"98",X"98",X"98",X"88",X"98",X"88",X"98",X"88",X"88",X"98",X"88",X"88",X"98",X"89",X"09",X"90",
		X"98",X"89",X"98",X"88",X"98",X"88",X"98",X"88",X"88",X"88",X"88",X"99",X"98",X"09",X"09",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"9D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"9D",X"90",X"99",X"99",
		X"00",X"D0",X"00",X"D0",X"00",X"90",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"9D",X"99",X"9D",X"99",X"D0",X"9D",X"00",X"D0",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"99",X"95",X"55",X"95",X"99",X"95",X"99",X"95",X"55",X"95",X"99",X"95",X"99",X"95",X"55",
		X"99",X"99",X"55",X"55",X"99",X"55",X"99",X"55",X"55",X"55",X"99",X"55",X"99",X"55",X"55",X"55",
		X"09",X"99",X"09",X"55",X"09",X"59",X"09",X"55",X"09",X"59",X"09",X"55",X"09",X"59",X"09",X"55",
		X"99",X"99",X"55",X"55",X"99",X"55",X"55",X"55",X"99",X"55",X"55",X"55",X"99",X"55",X"55",X"55",
		X"99",X"99",X"55",X"59",X"55",X"59",X"55",X"95",X"55",X"55",X"55",X"99",X"55",X"55",X"55",X"55",
		X"55",X"90",X"55",X"90",X"59",X"59",X"99",X"55",X"55",X"55",X"55",X"95",X"55",X"55",X"55",X"95",
		X"55",X"55",X"55",X"55",X"55",X"99",X"55",X"00",X"55",X"09",X"55",X"99",X"55",X"95",X"95",X"59",
		X"55",X"95",X"55",X"55",X"55",X"99",X"55",X"00",X"59",X"99",X"99",X"55",X"99",X"55",X"00",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"55",X"05",X"99",X"00",X"95",X"00",X"95",X"00",X"95",X"00",X"95",X"00",X"95",X"00",X"50",
		X"55",X"05",X"99",X"59",X"95",X"95",X"95",X"55",X"95",X"05",X"95",X"05",X"95",X"05",X"50",X"00",
		X"04",X"AA",X"00",X"AD",X"00",X"DA",X"00",X"AA",X"00",X"AA",X"04",X"AA",X"04",X"AA",X"04",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AD",X"AA",X"AA",X"DD",X"AA",X"AA",X"DA",X"AA",X"AA",X"AA",X"AA",X"AD",
		X"4A",X"AA",X"04",X"AD",X"4D",X"AA",X"4A",X"AA",X"04",X"AA",X"04",X"AA",X"4D",X"AA",X"4A",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AD",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A5",X"AA",X"56",X"AA",X"56",
		X"4A",X"AA",X"4A",X"AA",X"04",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"44",X"00",X"00",
		X"DA",X"A5",X"AA",X"55",X"AA",X"88",X"AA",X"88",X"AA",X"58",X"A4",X"48",X"40",X"04",X"00",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"48",X"00",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"00",X"14",X"00",X"11",X"40",X"11",X"14",X"11",X"11",X"11",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"44",X"44",
		X"14",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"14",X"00",X"40",X"00",X"00",X"00",
		X"88",X"88",X"77",X"77",X"58",X"88",X"35",X"55",X"32",X"22",X"39",X"99",X"39",X"BB",X"39",X"99",
		X"44",X"00",X"77",X"00",X"44",X"00",X"34",X"44",X"32",X"22",X"39",X"99",X"39",X"BB",X"39",X"99",
		X"39",X"B9",X"39",X"B9",X"39",X"B9",X"39",X"B9",X"39",X"B9",X"39",X"B9",X"39",X"B9",X"39",X"B9",
		X"39",X"B9",X"39",X"B9",X"39",X"B9",X"39",X"B9",X"39",X"B9",X"39",X"B9",X"39",X"B9",X"39",X"B9",
		X"39",X"B9",X"39",X"B9",X"39",X"B9",X"39",X"B9",X"39",X"B9",X"32",X"22",X"35",X"44",X"35",X"00",
		X"39",X"B9",X"39",X"B9",X"39",X"B9",X"39",X"B9",X"39",X"B9",X"32",X"22",X"34",X"44",X"34",X"00",
		X"44",X"44",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"44",X"44",
		X"44",X"00",X"66",X"44",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"44",X"44",X"00",
		X"00",X"44",X"00",X"66",X"04",X"66",X"46",X"66",X"46",X"66",X"04",X"66",X"00",X"66",X"00",X"44",
		X"00",X"66",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"66",X"44",X"66",X"00",X"64",X"00",X"40",X"00",X"40",X"00",X"64",X"00",X"66",X"00",X"66",X"44",
		X"44",X"44",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"44",X"44",
		X"AA",X"4A",X"99",X"4A",X"AA",X"4A",X"44",X"94",X"AA",X"A4",X"AA",X"44",X"4A",X"A4",X"94",X"AB",
		X"4A",X"77",X"49",X"74",X"A4",X"74",X"A4",X"74",X"A4",X"49",X"A4",X"99",X"AA",X"99",X"AA",X"94",
		X"AA",X"AB",X"99",X"BB",X"AA",X"4B",X"99",X"4B",X"AA",X"A4",X"99",X"94",X"AA",X"AA",X"99",X"99",
		X"AA",X"94",X"AA",X"49",X"AA",X"4A",X"AA",X"49",X"AA",X"AA",X"AA",X"99",X"AA",X"AA",X"AA",X"99",
		X"AA",X"AA",X"44",X"99",X"A4",X"AA",X"99",X"49",X"AA",X"A4",X"99",X"AA",X"AA",X"AA",X"99",X"AA",
		X"AA",X"AA",X"99",X"99",X"AA",X"AA",X"99",X"99",X"AA",X"AA",X"99",X"94",X"AA",X"A4",X"99",X"4B",
		X"AA",X"AA",X"99",X"94",X"AA",X"47",X"99",X"47",X"AA",X"47",X"99",X"77",X"AA",X"77",X"99",X"77",
		X"AA",X"4B",X"99",X"4B",X"AA",X"4B",X"99",X"94",X"AA",X"A4",X"99",X"99",X"AA",X"AA",X"99",X"99",
		X"AA",X"AA",X"99",X"99",X"AA",X"AA",X"44",X"99",X"99",X"AA",X"44",X"99",X"4B",X"4A",X"94",X"49",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"B4",X"99",X"B4",X"AA",X"B4",X"99",X"B4",X"AA",X"44",X"99",X"94",X"AA",X"AA",X"99",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"06",X"00",X"69",X"66",X"97",X"99",X"72",X"77",X"26",X"22",X"61",X"66",X"10",X"11",X"00",
		X"66",X"C0",X"77",X"CC",X"22",X"CC",X"66",X"CC",X"11",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"62",X"00",X"62",X"00",X"62",X"00",X"62",X"00",X"62",X"00",X"62",X"00",X"62",X"00",X"62",
		X"84",X"AC",X"84",X"AC",X"84",X"AC",X"84",X"AC",X"84",X"AC",X"84",X"AC",X"84",X"AC",X"84",X"AC",
		X"00",X"62",X"00",X"62",X"00",X"62",X"00",X"62",X"00",X"62",X"00",X"62",X"00",X"62",X"00",X"62",
		X"84",X"AC",X"84",X"AC",X"84",X"AC",X"84",X"AC",X"84",X"AC",X"84",X"AC",X"84",X"AC",X"84",X"AC",
		X"DB",X"59",X"DB",X"59",X"DB",X"59",X"DB",X"59",X"DB",X"59",X"DB",X"59",X"DB",X"59",X"DB",X"59",
		X"37",X"10",X"37",X"10",X"37",X"10",X"37",X"10",X"37",X"10",X"37",X"10",X"37",X"10",X"37",X"10",
		X"DB",X"59",X"DB",X"59",X"DB",X"59",X"DB",X"59",X"DB",X"59",X"DC",X"C5",X"DC",X"11",X"CC",X"11",
		X"37",X"10",X"37",X"10",X"37",X"61",X"37",X"66",X"13",X"22",X"11",X"1C",X"CC",X"48",X"55",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"02",X"00",X"21",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"01",
		X"00",X"12",X"01",X"21",X"12",X"12",X"21",X"21",X"12",X"02",X"21",X"20",X"12",X"12",X"21",X"21",
		X"00",X"12",X"00",X"21",X"00",X"12",X"00",X"21",X"00",X"12",X"00",X"21",X"00",X"12",X"01",X"21",
		X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",
		X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",
		X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",
		X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",
		X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"00",X"12",X"66",X"20",X"66",X"06",X"66",X"66",X"66",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"01",X"44",X"02",X"44",X"01",X"44",X"02",X"44",X"01",X"44",X"12",X"44",X"21",X"44",X"12",
		X"44",X"44",X"40",X"00",X"06",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"44",X"21",X"44",X"12",X"00",X"21",X"66",X"12",X"66",X"21",X"66",X"12",X"60",X"21",X"60",X"12",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"00",X"00",X"00",X"00",X"40",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"02",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"01",X"44",X"02",X"44",X"01",X"44",X"02",X"44",X"01",X"44",X"02",X"44",X"01",X"44",X"02",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"40",X"44",X"03",X"44",X"33",
		X"44",X"44",X"44",X"44",X"44",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"03",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"33",X"03",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"40",X"44",X"00",X"44",X"00",
		X"44",X"44",X"44",X"44",X"44",X"40",X"44",X"00",X"44",X"00",X"44",X"00",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"03",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"03",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"40",X"44",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"40",X"44",X"40",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"40",X"00",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"40",X"00",X"40",X"00",X"40",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"00",X"44",X"00",X"44",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"00",X"00",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"11",X"11",X"11",X"44",X"14",X"44",X"14",X"44",X"14",X"14",X"14",X"41",X"14",X"44",X"11",X"11",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"00",X"44",X"33",X"00",X"33",X"33",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"00",X"00",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"77",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"77",X"44",
		X"44",X"44",X"44",X"74",X"44",X"77",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"74",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"33",X"44",X"33",X"43",X"43",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"43",X"33",X"44",X"33",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"34",X"44",X"43",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"40",X"44",X"40",X"44",X"00",X"44",X"00",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",
		X"33",X"30",X"33",X"30",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"30",X"00",X"30",X"00",
		X"11",X"11",X"10",X"00",X"10",X"00",X"10",X"00",X"10",X"00",X"10",X"00",X"10",X"00",X"10",X"00",
		X"00",X"44",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"04",X"44",X"00",X"44",X"00",X"44",X"00",X"44",
		X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"00",X"02",X"00",X"29",X"00",X"99",X"00",X"99",X"02",X"99",X"02",X"99",X"29",X"99",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"11",X"11",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"11",X"11",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"94",X"44",X"94",X"44",X"94",X"00",X"94",X"CC",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"04",X"44",X"C0",X"44",
		X"44",X"44",X"44",X"44",X"44",X"42",X"44",X"42",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"42",X"44",X"42",X"44",X"42",X"44",X"22",X"44",X"22",X"44",X"44",X"44",X"44",X"44",X"44",X"24",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"24",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"29",X"99",X"29",X"99",X"99",X"92",X"99",X"90",X"99",X"05",X"92",X"55",X"90",X"55",X"0C",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"CC",X"CC",X"55",X"CC",X"55",X"CC",X"55",X"CC",X"55",X"0C",X"55",X"00",X"C5",X"00",X"00",
		X"0C",X"CC",X"CC",X"CC",X"5C",X"C5",X"5C",X"55",X"CC",X"55",X"CC",X"C5",X"CC",X"C0",X"CC",X"0F",
		X"CC",X"04",X"5C",X"F0",X"50",X"FF",X"00",X"FF",X"F0",X"FF",X"FF",X"F0",X"FF",X"0F",X"FF",X"FF",
		X"CC",X"FF",X"CC",X"FF",X"CC",X"FF",X"C0",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"0F",X"F0",
		X"FF",X"F0",X"F0",X"F0",X"0F",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"00",X"44",X"00",X"44",
		X"14",X"44",X"14",X"44",X"14",X"44",X"14",X"44",X"14",X"44",X"14",X"44",X"14",X"44",X"11",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"44",X"44",X"44",X"44",X"44",X"04",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"F0",X"FF",X"F0",X"FF",X"F0",X"FF",X"F0",X"FF",X"F0",X"FF",X"0F",X"0F",X"0F",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"04",X"44",X"04",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"44",X"44",X"44",X"44",X"44",X"04",X"44",X"04",X"44",X"00",X"44",X"00",X"44",X"00",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"33",X"00",X"33",X"03",X"33",X"33",X"33",
		X"03",X"04",X"33",X"30",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"66",X"66",X"66",X"00",X"66",X"11",X"00",X"00",X"11",X"33",X"00",X"33",X"33",X"33",X"33",X"30",
		X"11",X"33",X"00",X"33",X"33",X"00",X"33",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"00",X"33",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"60",X"66",X"01",X"60",X"11",X"01",X"10",
		X"66",X"60",X"66",X"01",X"66",X"11",X"60",X"11",X"01",X"11",X"11",X"10",X"11",X"03",X"11",X"33",
		X"11",X"03",X"10",X"33",X"00",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"30",X"33",X"00",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"06",X"66",X"60",X"66",X"66",X"66",X"66",
		X"60",X"21",X"00",X"12",X"01",X"21",X"02",X"12",X"21",X"21",X"12",X"12",X"01",X"21",X"60",X"12",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"06",X"66",X"10",X"66",
		X"66",X"01",X"66",X"60",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"21",X"21",X"12",X"10",X"21",X"06",X"12",X"66",X"21",X"66",X"12",X"66",X"21",X"66",X"10",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"20",X"66",X"06",X"66",X"06",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"60",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"40",X"44",X"06",X"44",X"66",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"00",X"40",X"00",
		X"44",X"66",X"44",X"66",X"40",X"66",X"40",X"66",X"00",X"66",X"10",X"66",X"10",X"66",X"11",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"30",X"00",X"33",X"00",X"33",X"00",
		X"01",X"66",X"01",X"66",X"30",X"06",X"33",X"10",X"03",X"11",X"03",X"01",X"00",X"30",X"00",X"33",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"40",X"44",X"03",X"44",X"33",X"44",X"33",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"33",X"44",X"33",X"40",X"33",X"40",X"33",X"40",X"33",X"03",X"33",X"03",X"33",X"03",X"33",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"30",X"33",X"30",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"33",X"00",X"33",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"30",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"30",
		X"11",X"66",X"01",X"06",X"30",X"10",X"33",X"11",X"33",X"11",X"33",X"01",X"33",X"30",X"33",X"33",
		X"66",X"66",X"66",X"60",X"66",X"60",X"66",X"06",X"06",X"06",X"10",X"06",X"11",X"06",X"11",X"00",
		X"03",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"11",X"30",X"00",X"33",X"11",X"33",X"11",X"30",X"11",X"01",X"10",X"11",X"03",X"11",X"33",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"60",X"66",X"00",X"66",X"11",X"00",X"11",
		X"66",X"01",X"66",X"11",X"60",X"11",X"01",X"11",X"11",X"10",X"11",X"03",X"11",X"33",X"10",X"33",
		X"11",X"11",X"11",X"10",X"11",X"03",X"10",X"33",X"03",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"03",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"30",X"33",X"00",
		X"11",X"33",X"00",X"33",X"03",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"30",X"33",X"00",
		X"33",X"00",X"33",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"00",X"33",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"04",X"44",X"30",X"44",X"33",X"44",X"33",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"00",X"33",X"00",X"33",X"00",X"33",X"03",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"03",X"00",X"33",X"00",X"33",X"00",X"33",X"03",X"33",X"33",X"33",X"33",X"33",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"33",X"44",X"33",X"04",X"33",X"04",X"33",X"30",X"33",X"30",X"33",X"30",X"33",X"33",X"33",X"33",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"04",X"44",X"04",X"44",X"04",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"12",X"00",X"21",X"00",X"12",X"00",X"21",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"12",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"21",
		X"00",X"00",X"00",X"21",X"00",X"12",X"01",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",
		X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"77",X"78",X"21",X"21",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"12",X"01",X"21",X"12",X"12",X"21",X"21",
		X"00",X"00",X"00",X"00",X"02",X"00",X"21",X"21",X"12",X"12",X"21",X"01",X"12",X"12",X"21",X"21",
		X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"88",X"12",X"21",X"88",
		X"12",X"12",X"21",X"21",X"12",X"10",X"21",X"20",X"12",X"10",X"21",X"04",X"12",X"04",X"21",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"04",X"44",X"00",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"12",X"10",X"21",X"20",X"12",X"10",X"21",X"20",X"12",X"10",X"21",X"20",X"12",X"10",X"21",X"20",
		X"00",X"12",X"00",X"21",X"00",X"12",X"01",X"21",X"02",X"12",X"21",X"21",X"12",X"12",X"21",X"21",
		X"12",X"10",X"21",X"20",X"12",X"10",X"21",X"20",X"12",X"10",X"21",X"20",X"12",X"12",X"21",X"21",
		X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",
		X"12",X"12",X"21",X"21",X"1A",X"12",X"21",X"77",X"12",X"88",X"21",X"28",X"12",X"12",X"21",X"21",
		X"12",X"12",X"21",X"21",X"12",X"12",X"AA",X"21",X"88",X"A7",X"10",X"7A",X"70",X"08",X"78",X"A1",
		X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",
		X"12",X"12",X"21",X"81",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",
		X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",
		X"12",X"44",X"21",X"44",X"12",X"44",X"21",X"44",X"10",X"44",X"04",X"44",X"44",X"44",X"44",X"44",
		X"12",X"10",X"21",X"04",X"12",X"04",X"21",X"44",X"12",X"44",X"21",X"44",X"12",X"44",X"21",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"42",X"44",X"42",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"42",X"44",X"42",X"44",X"42",X"44",X"22",X"44",X"22",X"44",X"44",X"44",X"44",X"44",X"44",X"24",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"24",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",
		X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",
		X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"20",X"21",X"12",X"12",X"21",X"21",
		X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",
		X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",
		X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",
		X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",
		X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"20",X"12",X"04",X"44",X"44",X"FF",X"44",X"F0",X"44",
		X"12",X"44",X"21",X"44",X"12",X"44",X"21",X"44",X"12",X"44",X"21",X"44",X"12",X"44",X"21",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"12",X"44",X"20",X"44",X"04",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"12",X"02",X"21",X"40",X"12",X"44",X"21",X"44",X"12",X"44",X"21",X"44",X"12",X"40",X"21",X"06",
		X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"02",X"12",X"00",X"21",X"66",X"02",X"66",X"60",
		X"10",X"66",X"06",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"12",X"12",X"21",X"20",X"12",X"10",X"21",X"06",X"12",X"06",X"21",X"66",X"12",X"66",X"00",X"66",
		X"44",X"44",X"44",X"44",X"44",X"44",X"00",X"44",X"66",X"44",X"66",X"04",X"66",X"60",X"66",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"60",X"66",X"01",X"66",X"10",X"60",X"03",
		X"44",X"44",X"44",X"44",X"44",X"24",X"44",X"22",X"44",X"42",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"22",X"44",X"22",X"44",X"22",X"44",X"22",X"44",X"22",X"44",X"42",X"44",X"42",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"04",X"44",X"30",X"44",X"30",X"44",
		X"44",X"44",X"44",X"24",X"44",X"24",X"44",X"42",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"00",X"44",X"21",X"44",X"00",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"40",X"00",X"00",X"12",X"21",X"00",X"22",X"12",X"00",X"21",X"44",X"02",
		X"44",X"44",X"44",X"40",X"44",X"40",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"04",X"40",X"10",X"44",X"21",X"04",X"02",X"10",X"00",X"21",X"44",X"12",X"44",X"02",X"44",X"40");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
