library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity obj_7u is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of obj_7u is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"F0",X"E0",X"00",X"00",X"00",X"40",X"30",X"70",X"60",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"1C",X"1C",X"1C",X"04",X"90",X"6C",X"EC",X"DC",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"38",X"1C",X"14",X"C0",X"F0",X"F8",X"B0",X"40",X"80",X"00",X"00",X"00",X"00",
		X"1E",X"1C",X"00",X"00",X"00",X"00",X"00",X"94",X"66",X"EC",X"E0",X"C0",X"00",X"00",X"00",X"00",
		X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"E0",X"00",X"00",X"00",X"00",X"26",X"9C",X"B8",X"B0",X"60",X"00",X"00",X"00",X"00",X"40",
		X"3C",X"38",X"00",X"00",X"00",X"E0",X"E0",X"C0",X"B8",X"30",X"60",X"00",X"00",X"00",X"00",X"60",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"8C",X"77",X"E6",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",
		X"1C",X"1C",X"1C",X"18",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"86",X"52",X"E2",X"C0",X"90",X"38",X"38",X"1C",X"0C",
		X"10",X"38",X"70",X"60",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"F8",X"F8",X"E8",X"70",X"78",X"38",X"98",X"80",X"C0",X"A0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"1C",X"0E",X"02",X"02",X"00",X"00",X"44",X"36",X"6E",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"88",X"1C",X"0E",X"02",X"02",X"00",X"00",X"44",X"36",X"68",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"08",X"1C",X"0E",X"02",X"02",X"00",X"00",X"44",X"06",X"6E",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"00",X"00",X"00",X"00",X"00",X"54",X"EF",X"DE",X"00",X"00",X"00",X"80",X"C0",X"00",X"00",
		X"1E",X"00",X"00",X"00",X"10",X"EF",X"CE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"08",X"04",X"04",X"23",X"C0",X"20",X"C8",X"C8",X"0C",X"0C",X"0E",X"04",X"60",X"60",X"00",
		X"08",X"08",X"04",X"04",X"23",X"C0",X"20",X"C4",X"CE",X"0E",X"0C",X"08",X"00",X"60",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"60",X"74",X"F4",X"EC",X"00",X"00",X"00",
		X"00",X"60",X"C0",X"E0",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"06",X"03",X"03",X"01",X"00",X"00",X"40",X"38",X"68",X"D0",X"00",X"00",X"00",X"00",
		X"00",X"04",X"06",X"03",X"03",X"01",X"00",X"20",X"9C",X"34",X"68",X"00",X"00",X"00",X"00",X"40",
		X"00",X"00",X"FC",X"FE",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"FE",X"FC",
		X"00",X"00",X"18",X"1C",X"BC",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"F8",X"F0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"18",X"1C",X"7C",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"F8",X"F0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",X"FE",X"7E",X"7E",X"3E",X"1E",X"06",X"00",X"00",X"00",X"00",
		X"7E",X"7E",X"7E",X"7E",X"FE",X"FE",X"FE",X"FC",X"FC",X"F8",X"F0",X"C0",X"00",X"00",X"00",X"00",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"52",X"52",X"52",X"F7",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"7E",X"7E",X"7E",X"7E",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"7E",X"7E",X"7E",X"7E",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"00",X"00",X"00",X"00",X"C0",X"F0",X"F8",X"FC",X"FC",X"FE",X"FE",X"FE",X"7E",X"7E",X"7E",X"7E",
		X"00",X"00",X"00",X"00",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"00",X"00",X"00",X"00",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"00",X"00",X"00",X"00",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"00",X"00",X"00",X"00",X"1E",X"1E",X"1E",X"1E",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"7C",X"3E",X"0E",X"00",X"00",X"00",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"FE",X"FE",X"7E",X"7E",X"7E",X"7C",X"FC",X"EC",X"0C",X"08",X"00",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",X"00",X"00",
		X"F0",X"FC",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7C",X"FC",X"EC",X"0C",X"08",X"00",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",X"00",X"00",
		X"F8",X"FC",X"7E",X"00",X"00",X"F0",X"FC",X"7E",X"7E",X"7E",X"7C",X"FC",X"EC",X"0C",X"08",X"00",
		X"1E",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"52",X"F7",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"FE",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F7",X"F7",X"F7",X"F7",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"F0",X"F8",X"FC",X"FC",X"FE",X"FE",X"FE",X"7E",X"7E",X"7E",X"7E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"E0",X"F8",X"F8",X"BC",X"FC",X"FC",X"F0",X"70",X"F8",X"38",X"9C",X"9F",X"B7",X"24",X"E0",
		X"C0",X"E0",X"F8",X"F8",X"BC",X"FD",X"FF",X"F7",X"7E",X"FE",X"3C",X"98",X"90",X"B0",X"20",X"E0",
		X"0E",X"1C",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"E0",X"F0",X"F0",X"68",X"FA",X"FF",X"FF",X"FF",X"F0",X"F8",X"C0",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"FF",X"FF",X"00",X"FF",X"FF",X"00",X"FF",X"FF",X"00",
		X"B6",X"B6",X"B6",X"B6",X"B6",X"36",X"76",X"66",X"EE",X"CC",X"9C",X"38",X"F8",X"E0",X"80",X"00",
		X"B6",X"B6",X"B6",X"B6",X"B6",X"B6",X"B6",X"B6",X"B6",X"B6",X"B6",X"B6",X"B6",X"B6",X"B6",X"B6",
		X"00",X"00",X"00",X"00",X"A0",X"60",X"20",X"60",X"C0",X"80",X"04",X"0E",X"0E",X"0E",X"2E",X"04",
		X"00",X"00",X"00",X"00",X"A0",X"60",X"20",X"60",X"C2",X"87",X"07",X"17",X"07",X"02",X"00",X"00",
		X"00",X"00",X"80",X"C0",X"40",X"C0",X"40",X"00",X"00",X"00",X"1A",X"38",X"38",X"38",X"38",X"10",
		X"00",X"00",X"1C",X"F8",X"C0",X"40",X"C0",X"40",X"00",X"00",X"1A",X"38",X"38",X"38",X"38",X"10",
		X"30",X"20",X"C0",X"C0",X"40",X"C0",X"40",X"00",X"00",X"1A",X"38",X"38",X"38",X"38",X"10",X"00",
		X"C0",X"80",X"00",X"80",X"C0",X"40",X"C0",X"40",X"00",X"00",X"1A",X"38",X"38",X"38",X"38",X"10",
		X"80",X"00",X"80",X"C0",X"40",X"C0",X"40",X"00",X"00",X"1A",X"38",X"38",X"38",X"38",X"10",X"00",
		X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"08",X"F0",X"F0",X"70",
		X"00",X"00",X"80",X"C0",X"C0",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"08",X"F0",X"F0",X"70",
		X"00",X"00",X"E0",X"C0",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"04",X"78",X"78",X"38",X"00",
		X"00",X"00",X"00",X"C0",X"00",X"80",X"80",X"80",X"00",X"00",X"00",X"08",X"70",X"70",X"70",X"30",
		X"00",X"00",X"E0",X"F0",X"F0",X"F0",X"C0",X"00",X"00",X"01",X"02",X"C0",X"00",X"E0",X"E0",X"E0",
		X"A0",X"10",X"A8",X"48",X"48",X"48",X"A8",X"18",X"B0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A0",X"10",X"A8",X"48",X"48",X"48",X"A8",X"18",X"B0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"A0",X"60",X"20",X"60",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"A0",X"70",X"30",X"70",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"A0",X"64",X"2E",X"6E",X"CE",X"84",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"20",X"C0",X"20",X"10",X"28",X"C0",X"20",X"1C",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"20",X"20",X"5C",X"84",X"48",X"50",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"C4",X"34",X"24",X"48",X"88",X"50",X"60",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"A0",X"10",X"A8",X"48",X"48",X"48",X"A8",X"18",X"B0",X"E0",
		X"00",X"00",X"00",X"20",X"A0",X"10",X"A8",X"48",X"48",X"48",X"A8",X"18",X"B0",X"E0",X"00",X"00",
		X"00",X"20",X"A0",X"10",X"A8",X"48",X"48",X"48",X"A8",X"18",X"B0",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"F8",X"04",X"00",X"00",X"20",X"C0",X"80",X"80",X"80",X"40",X"20",X"00",X"00",X"00",X"00",
		X"00",X"80",X"00",X"08",X"10",X"20",X"D0",X"00",X"80",X"80",X"40",X"20",X"00",X"00",X"00",X"00",
		X"80",X"04",X"08",X"10",X"30",X"60",X"D0",X"88",X"80",X"C0",X"60",X"10",X"00",X"00",X"00",X"00",
		X"00",X"08",X"30",X"00",X"00",X"00",X"00",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"06",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"08",X"00",X"00",X"00",X"00",X"20",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"3E",X"1C",X"08",X"10",X"20",X"40",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"FD",X"FB",X"E0",X"00",X"E0",X"C0",X"80",X"01",X"03",X"07",X"1F",
		X"FF",X"FF",X"FF",X"FF",X"FC",X"F2",X"CC",X"3C",X"18",X"00",X"00",X"00",X"03",X"0F",X"3F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"F8",X"F0",X"01",X"06",X"18",X"E0",X"00",X"01",X"07",X"1F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"01",X"00",X"FE",X"00",X"00",X"01",X"03",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"F8",X"E0",X"01",X"06",X"18",X"E0",X"00",X"01",X"07",X"1F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F1",X"F1",X"10",X"10",X"01",X"01",X"11",X"11",X"1F",X"1F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"1F",X"11",X"11",X"01",X"01",X"11",X"11",X"F1",X"F1",
		X"FF",X"FF",X"FF",X"F1",X"11",X"10",X"00",X"01",X"11",X"11",X"11",X"1F",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"01",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"7E",X"3C",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"FD",X"FB",X"E6",X"00",X"E0",X"C0",X"00",X"01",X"03",X"07",X"1F",
		X"FF",X"FF",X"FF",X"FF",X"FC",X"F2",X"CC",X"3C",X"70",X"00",X"00",X"00",X"03",X"0F",X"3F",X"FF",
		X"E0",X"10",X"88",X"34",X"6C",X"42",X"60",X"B0",X"50",X"48",X"28",X"28",X"50",X"B0",X"60",X"80",
		X"F0",X"98",X"6C",X"94",X"0A",X"0A",X"0A",X"0A",X"0A",X"12",X"34",X"E4",X"C8",X"10",X"E0",X"00",
		X"F0",X"18",X"E8",X"34",X"14",X"0A",X"0A",X"0A",X"8A",X"6A",X"3A",X"B4",X"AC",X"98",X"70",X"C0",
		X"00",X"00",X"80",X"E0",X"90",X"00",X"80",X"40",X"A0",X"A0",X"A0",X"A0",X"40",X"80",X"00",X"00",
		X"00",X"00",X"00",X"F0",X"88",X"68",X"94",X"14",X"14",X"34",X"C8",X"10",X"E0",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"30",X"D0",X"28",X"28",X"28",X"A8",X"58",X"90",X"50",X"E0",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"80",X"40",X"40",X"40",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"60",X"90",X"60",X"A0",X"D0",X"20",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"A0",X"50",X"50",X"90",X"50",X"60",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"10",X"00",X"00",X"08",X"00",X"00",X"10",X"80",X"00",X"00",X"00",X"00",
		X"80",X"02",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"02",X"80",X"00",
		X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"40",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"00",X"20",X"40",X"00",X"00",X"00",X"00",
		X"00",X"20",X"10",X"90",X"48",X"48",X"48",X"48",X"48",X"00",X"10",X"20",X"00",X"00",X"00",X"00",
		X"00",X"E0",X"D0",X"E8",X"E8",X"E8",X"E8",X"E8",X"E8",X"E8",X"D0",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"0C",X"0C",X"00",X"E0",X"1F",X"00",X"A0",X"70",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C4",X"20",X"00",X"00",X"80",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"24",X"00",X"00",X"80",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"C0",X"28",X"00",X"00",X"80",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"80",X"80",X"80",X"80",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"20",
		X"00",X"00",X"80",X"80",X"80",X"80",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"20",
		X"00",X"00",X"80",X"88",X"80",X"80",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"20",
		X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"00",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"44",X"40",X"C0",X"42",X"02",X"00",X"60",X"E0",X"E8",X"E0",X"E0",X"40",
		X"00",X"E0",X"F0",X"FC",X"D8",X"48",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"C0",X"80",X"80",
		X"00",X"C0",X"EE",X"F0",X"70",X"30",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C8",X"FC",X"E2",X"D5",X"48",X"C8",X"B4",X"48",X"40",X"20",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"F0",X"10",X"1F",X"FF",X"F0",X"30",X"30",X"30",X"30",X"10",X"10",X"30",X"30",X"F0",
		X"67",X"63",X"61",X"30",X"18",X"0F",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"00",X"E6",X"F6",X"FE",X"EE",X"E6",X"E6",X"7E",X"E6",X"E6",X"EE",X"FE",X"F6",
		X"00",X"00",X"80",X"E0",X"70",X"38",X"1C",X"8C",X"CC",X"66",X"66",X"66",X"66",X"66",X"E6",X"FE",
		X"66",X"67",X"63",X"31",X"18",X"0C",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"E6",X"FE",X"33",X"33",X"33",X"00",
		X"FE",X"30",X"30",X"30",X"00",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"00",X"00",X"00",X"60",X"C0",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"0C",X"12",X"07",X"E7",
		X"FF",X"FF",X"F0",X"10",X"1F",X"FF",X"F0",X"30",X"30",X"30",X"30",X"10",X"10",X"30",X"30",X"F0",
		X"FF",X"FF",X"70",X"10",X"9F",X"FF",X"70",X"30",X"30",X"30",X"30",X"10",X"10",X"30",X"30",X"70",
		X"FF",X"F0",X"10",X"1F",X"FF",X"F0",X"B0",X"30",X"30",X"30",X"30",X"30",X"10",X"10",X"30",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"80",X"80",X"80",X"00",X"80",X"00",X"00",X"00",X"80",X"00",X"80",X"40",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"9E",X"5C",X"70",X"E0",X"14",X"1C",X"78",X"80",X"00",X"00",X"30",X"F8",X"F8",X"F8",X"70",
		X"00",X"9E",X"5C",X"70",X"E4",X"1C",X"18",X"70",X"90",X"1C",X"1E",X"1E",X"AE",X"1C",X"00",X"00",
		X"3C",X"B8",X"50",X"60",X"E0",X"1C",X"1E",X"7E",X"9E",X"1C",X"00",X"00",X"A0",X"18",X"00",X"00",
		X"CE",X"2C",X"FA",X"D6",X"3C",X"78",X"98",X"18",X"04",X"00",X"A0",X"18",X"00",X"00",X"00",X"00",
		X"03",X"0F",X"1E",X"9C",X"78",X"10",X"10",X"E0",X"30",X"50",X"A0",X"30",X"30",X"10",X"00",X"00",
		X"03",X"0F",X"1E",X"9C",X"78",X"10",X"10",X"E0",X"30",X"4C",X"8E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"F8",X"04",X"00",X"00",X"00",X"00",X"A0",X"A0",X"A0",X"B0",X"D0",X"80",X"80",X"80",X"00",
		X"00",X"F8",X"04",X"00",X"00",X"00",X"FC",X"B8",X"B8",X"B8",X"B0",X"D0",X"80",X"80",X"80",X"00",
		X"00",X"F8",X"04",X"FE",X"AE",X"5C",X"FC",X"B8",X"B8",X"B8",X"B0",X"D0",X"80",X"80",X"80",X"00",
		X"FC",X"FE",X"FE",X"AE",X"5E",X"FC",X"FC",X"B8",X"B8",X"B8",X"B0",X"D0",X"80",X"80",X"80",X"00",
		X"00",X"F8",X"04",X"00",X"00",X"00",X"00",X"A0",X"A0",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"F8",X"04",X"00",X"00",X"00",X"00",X"A0",X"A0",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"80",X"80",X"80",X"80",X"80",
		X"00",X"00",X"40",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"00",X"20",X"40",X"80",X"80",X"80",
		X"00",X"00",X"20",X"10",X"90",X"48",X"48",X"48",X"48",X"48",X"08",X"10",X"20",X"80",X"80",X"80",
		X"00",X"00",X"E0",X"D0",X"E8",X"E8",X"E8",X"E8",X"E8",X"E8",X"E8",X"D0",X"E0",X"80",X"80",X"80",
		X"00",X"00",X"C0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"C0",X"80",X"80",X"80",
		X"00",X"00",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"80",
		X"00",X"00",X"00",X"C0",X"80",X"40",X"40",X"40",X"40",X"40",X"00",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"60",X"10",X"68",X"34",X"14",X"00",X"14",X"34",X"68",X"10",X"60",X"00",X"00",X"00",
		X"70",X"78",X"0C",X"76",X"1B",X"0B",X"0B",X"00",X"0B",X"0B",X"1B",X"76",X"0C",X"78",X"70",X"00",
		X"00",X"F0",X"F8",X"FC",X"1E",X"0E",X"8E",X"CE",X"8E",X"0E",X"1E",X"FC",X"F8",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"E0",X"F8",X"38",X"98",X"D8",X"98",X"38",X"F8",X"F0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"30",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"40",X"40",X"40",X"C0",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"E0",X"E0",X"E0",X"60",X"40",X"40",X"00",X"00",X"40",X"60",X"00",
		X"00",X"00",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"50",X"50",X"50",X"50",X"58",X"58",X"10",
		X"00",X"00",X"40",X"40",X"40",X"40",X"00",X"40",X"40",X"40",X"40",X"50",X"50",X"58",X"58",X"10",
		X"00",X"00",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"50",X"50",X"50",X"58",X"58",X"10",
		X"00",X"00",X"00",X"00",X"A0",X"60",X"20",X"60",X"C0",X"80",X"04",X"14",X"00",X"00",X"00",X"00",
		X"00",X"40",X"80",X"40",X"20",X"20",X"C0",X"00",X"20",X"E0",X"00",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"00",X"18",X"20",X"40",X"A4",X"18",X"A4",X"44",X"48",X"B0",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"0E",X"90",X"60",X"90",X"08",X"90",X"60",X"90",X"08",
		X"00",X"40",X"00",X"00",X"00",X"00",X"80",X"40",X"A0",X"10",X"A8",X"48",X"44",X"B4",X"40",X"00",
		X"00",X"00",X"04",X"84",X"40",X"40",X"42",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"50",X"80",X"80",X"20",X"10",X"10",X"D0",X"20",X"00",X"40",X"40",X"00",X"00",X"00",X"00",
		X"00",X"40",X"20",X"20",X"98",X"64",X"24",X"90",X"50",X"40",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"60",X"D0",X"D0",X"D0",X"84",X"04",X"28",X"00",X"20",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"20",X"E0",X"C0",X"80",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"20",X"A0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"60",X"E0",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"9C",X"7E",X"1F",X"1F",X"E6",X"30",X"50",X"A0",X"30",X"30",X"10",X"00",X"00",
		X"00",X"80",X"C0",X"64",X"38",X"10",X"10",X"88",X"88",X"4C",X"3C",X"DC",X"FC",X"BC",X"98",X"00",
		X"00",X"8C",X"9E",X"5E",X"DE",X"3C",X"4C",X"88",X"88",X"10",X"10",X"38",X"64",X"C0",X"00",X"00",
		X"00",X"00",X"08",X"18",X"18",X"D0",X"28",X"18",X"F3",X"0F",X"0F",X"3E",X"CC",X"80",X"80",X"80",
		X"80",X"80",X"80",X"00",X"00",X"80",X"40",X"40",X"2E",X"AC",X"58",X"40",X"F0",X"F8",X"F8",X"70",
		X"30",X"F8",X"F8",X"F8",X"40",X"50",X"AC",X"2E",X"40",X"40",X"80",X"00",X"00",X"80",X"80",X"80",
		X"E0",X"E0",X"E0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C8",X"D0",X"B0",X"A0",X"40",X"40",X"C0",X"C0",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",
		X"F0",X"E0",X"E0",X"C0",X"C0",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"50",X"00",X"80",X"40",X"20",
		X"F8",X"F0",X"E0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"04",X"00",X"00",X"06",X"0C",X"00",X"00",
		X"80",X"00",X"02",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"07",X"07",X"07",X"7F",X"E7",X"E7",X"E7",X"E7",X"7F",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"FD",X"FF",X"FF",X"FF",X"CF",X"FF",X"FF",X"FF",X"FF",X"07",X"01",X"00",X"00",
		X"01",X"01",X"01",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"01",X"00",X"00",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"FF",X"7C",X"3C",X"30",X"2C",X"2C",X"2C",X"2C",X"70",X"FF",X"00",X"00",X"01",
		X"FF",X"FF",X"FF",X"01",X"00",X"00",X"FF",X"7C",X"30",X"2C",X"2C",X"70",X"FF",X"00",X"00",X"01",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"30",X"2C",X"20",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
