library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity domino_sp_bits_3 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of domino_sp_bits_3 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"91",X"00",X"00",X"99",X"91",
		X"99",X"00",X"91",X"11",X"92",X"99",X"11",X"91",X"52",X"11",X"11",X"91",X"52",X"11",X"11",X"91",
		X"99",X"99",X"11",X"19",X"00",X"00",X"11",X"91",X"00",X"00",X"99",X"19",X"00",X"00",X"00",X"91",
		X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"91",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"9C",X"90",X"00",X"00",X"CC",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"AA",X"99",X"00",X"00",X"A2",X"C9",X"00",X"00",X"99",X"C9",X"00",X"00",X"9C",X"C9",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"00",X"00",
		X"00",X"C9",X"99",X"00",X"00",X"CC",X"44",X"00",X"09",X"99",X"99",X"00",X"99",X"44",X"99",X"00",
		X"94",X"44",X"99",X"00",X"44",X"99",X"99",X"00",X"44",X"44",X"99",X"00",X"99",X"44",X"99",X"00",
		X"44",X"44",X"99",X"00",X"99",X"99",X"99",X"00",X"CC",X"22",X"99",X"00",X"CC",X"29",X"99",X"00",
		X"99",X"92",X"99",X"00",X"00",X"92",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"90",X"99",X"00",
		X"00",X"90",X"99",X"00",X"00",X"90",X"99",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"9C",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"9A",X"99",X"00",X"00",X"92",X"CC",X"00",X"00",X"99",X"9C",X"00",X"00",X"C9",X"CC",X"00",
		X"00",X"49",X"49",X"00",X"00",X"99",X"C9",X"00",X"00",X"99",X"99",X"00",X"00",X"C9",X"90",X"00",
		X"09",X"CC",X"99",X"00",X"99",X"9C",X"49",X"00",X"94",X"99",X"44",X"00",X"94",X"44",X"99",X"00",
		X"94",X"44",X"99",X"00",X"94",X"99",X"99",X"00",X"99",X"44",X"99",X"00",X"9C",X"44",X"99",X"00",
		X"9C",X"44",X"99",X"00",X"99",X"99",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"29",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"9C",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"AA",X"C9",X"00",X"00",X"2A",X"C9",X"00",X"00",X"99",X"C9",X"00",X"00",X"CC",X"99",X"00",
		X"00",X"C9",X"CC",X"00",X"00",X"99",X"CC",X"00",X"00",X"99",X"CC",X"00",X"00",X"99",X"CC",X"00",
		X"00",X"99",X"99",X"00",X"00",X"09",X"44",X"00",X"09",X"99",X"44",X"99",X"9D",X"99",X"44",X"99",
		X"9D",X"99",X"4F",X"99",X"9D",X"99",X"99",X"99",X"9D",X"CC",X"99",X"99",X"9D",X"CC",X"99",X"99",
		X"9D",X"CC",X"99",X"99",X"9D",X"99",X"99",X"99",X"9D",X"99",X"99",X"99",X"9D",X"99",X"99",X"99",
		X"9D",X"9F",X"F9",X"99",X"9D",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"09",X"90",X"22",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"99",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"CC",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"A9",X"99",X"00",X"00",X"29",X"99",X"00",X"00",X"9C",X"99",X"00",X"00",X"CC",X"99",X"00",
		X"00",X"9C",X"CC",X"00",X"00",X"99",X"C9",X"00",X"00",X"99",X"C9",X"00",X"00",X"99",X"C9",X"00",
		X"00",X"99",X"99",X"00",X"00",X"9C",X"99",X"00",X"00",X"99",X"94",X"00",X"99",X"99",X"44",X"90",
		X"D9",X"99",X"44",X"90",X"D9",X"99",X"49",X"90",X"D9",X"99",X"99",X"90",X"D9",X"99",X"99",X"90",
		X"D9",X"99",X"99",X"90",X"D9",X"99",X"99",X"90",X"D9",X"99",X"99",X"90",X"D9",X"99",X"99",X"90",
		X"D9",X"99",X"99",X"90",X"D9",X"F9",X"99",X"90",X"D9",X"99",X"99",X"90",X"99",X"99",X"99",X"90",
		X"00",X"99",X"90",X"00",X"00",X"11",X"90",X"00",X"00",X"11",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"9C",X"00",X"00",X"C9",X"CC",X"00",X"00",X"CC",X"CC",X"00",
		X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"C9",X"00",X"00",X"99",X"99",X"00",
		X"00",X"49",X"49",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"99",X"44",X"00",
		X"00",X"99",X"44",X"00",X"00",X"99",X"44",X"00",X"00",X"99",X"44",X"00",X"00",X"99",X"44",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"92",X"00",X"00",X"99",X"92",X"00",
		X"00",X"91",X"22",X"00",X"00",X"11",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"11",X"99",X"00",
		X"00",X"11",X"91",X"00",X"00",X"11",X"91",X"00",X"00",X"91",X"99",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"C9",X"99",X"00",X"00",X"CC",X"9C",X"00",
		X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"9C",X"CC",X"00",X"00",X"99",X"99",X"00",
		X"00",X"94",X"94",X"00",X"00",X"44",X"44",X"00",X"00",X"99",X"44",X"00",X"00",X"99",X"44",X"00",
		X"00",X"99",X"44",X"90",X"00",X"99",X"44",X"90",X"00",X"99",X"44",X"90",X"00",X"99",X"94",X"90",
		X"00",X"99",X"99",X"90",X"00",X"99",X"22",X"90",X"00",X"99",X"29",X"90",X"00",X"99",X"99",X"90",
		X"00",X"99",X"91",X"90",X"00",X"99",X"11",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"11",X"00",
		X"00",X"99",X"11",X"00",X"00",X"99",X"11",X"00",X"00",X"09",X"91",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"99",X"CC",X"00",X"00",X"99",X"9C",X"00",X"00",X"99",X"9C",X"00",
		X"00",X"09",X"9C",X"00",X"00",X"09",X"9C",X"00",X"00",X"09",X"CC",X"00",X"00",X"09",X"CC",X"00",
		X"00",X"09",X"CC",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",
		X"00",X"99",X"44",X"99",X"00",X"44",X"CC",X"C9",X"99",X"44",X"99",X"C9",X"19",X"44",X"94",X"C9",
		X"11",X"44",X"44",X"C9",X"99",X"99",X"99",X"99",X"92",X"99",X"44",X"00",X"22",X"44",X"94",X"00",
		X"22",X"44",X"99",X"99",X"22",X"99",X"99",X"91",X"92",X"29",X"99",X"91",X"99",X"99",X"00",X"11",
		X"09",X"00",X"00",X"11",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"CC",X"00",X"00",X"99",X"9C",X"00",
		X"00",X"99",X"9C",X"00",X"00",X"99",X"9C",X"00",X"00",X"09",X"9C",X"00",X"00",X"09",X"CC",X"00",
		X"00",X"09",X"CC",X"00",X"00",X"09",X"CC",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"99",X"99",
		X"00",X"00",X"99",X"9C",X"00",X"99",X"44",X"9C",X"00",X"44",X"CC",X"CC",X"00",X"44",X"99",X"C9",
		X"00",X"44",X"94",X"C9",X"00",X"44",X"44",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"00",
		X"00",X"44",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"29",X"00",X"00",
		X"00",X"99",X"00",X"00",X"09",X"92",X"00",X"00",X"99",X"22",X"00",X"00",X"19",X"29",X"00",X"00",
		X"11",X"99",X"00",X"00",X"11",X"99",X"00",X"00",X"99",X"11",X"00",X"00",X"99",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"9C",X"99",X"00",X"00",X"CC",X"99",X"00",X"00",X"CC",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"A9",X"C9",X"00",X"00",X"99",X"C9",X"00",X"00",X"9C",X"C9",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"9F",X"CC",X"00",
		X"00",X"99",X"CC",X"00",X"00",X"9C",X"9C",X"00",X"09",X"99",X"CC",X"00",X"09",X"94",X"CC",X"00",
		X"09",X"94",X"99",X"00",X"09",X"99",X"99",X"00",X"09",X"44",X"49",X"00",X"09",X"44",X"49",X"00",
		X"00",X"44",X"49",X"00",X"00",X"99",X"99",X"00",X"00",X"22",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"92",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"C9",X"00",
		X"00",X"99",X"C9",X"00",X"00",X"99",X"C9",X"00",X"00",X"CC",X"CC",X"00",X"00",X"4C",X"CC",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"9C",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"9C",X"99",X"00",X"00",X"CC",X"C9",X"00",X"00",X"CC",X"CC",X"00",
		X"00",X"99",X"CC",X"00",X"00",X"99",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"99",X"44",X"00",
		X"00",X"44",X"99",X"00",X"00",X"99",X"92",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"91",X"00",
		X"00",X"99",X"11",X"00",X"00",X"92",X"11",X"00",X"00",X"99",X"11",X"00",X"00",X"91",X"99",X"00",
		X"00",X"99",X"11",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"9C",X"00",X"00",X"C9",X"CC",X"00",X"00",X"CC",X"CC",X"00",
		X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"C9",X"C9",X"00",X"00",X"99",X"99",X"00",
		X"00",X"44",X"49",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"94",X"00",X"00",X"44",X"44",X"00",X"00",X"49",X"99",X"00",
		X"00",X"99",X"29",X"00",X"00",X"22",X"22",X"00",X"00",X"99",X"92",X"00",X"00",X"91",X"22",X"00",
		X"00",X"11",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"11",X"99",X"00",X"00",X"11",X"91",X"00",
		X"00",X"11",X"99",X"00",X"00",X"91",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"9C",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"CC",X"00",X"00",X"99",X"CC",X"00",X"00",X"C9",X"CC",X"00",
		X"00",X"CC",X"C9",X"00",X"00",X"CC",X"C9",X"00",X"00",X"99",X"99",X"00",X"00",X"94",X"99",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"49",X"00",X"00",X"44",X"49",X"00",
		X"00",X"99",X"49",X"00",X"00",X"99",X"49",X"00",X"00",X"44",X"49",X"00",X"00",X"99",X"49",X"00",
		X"00",X"22",X"99",X"00",X"00",X"29",X"29",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"99",X"00",
		X"00",X"90",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"DD",X"9C",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"CC",X"00",X"99",X"99",X"9C",X"00",
		X"99",X"99",X"94",X"00",X"99",X"99",X"44",X"00",X"9F",X"9C",X"9C",X"00",X"99",X"99",X"9C",X"00",
		X"99",X"99",X"C9",X"00",X"99",X"49",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"94",X"00",
		X"99",X"94",X"49",X"00",X"DD",X"94",X"44",X"00",X"99",X"99",X"99",X"00",X"99",X"94",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"92",X"00",X"99",X"09",X"22",X"00",X"99",X"09",X"22",X"00",
		X"9F",X"09",X"22",X"00",X"99",X"09",X"92",X"00",X"99",X"09",X"29",X"00",X"99",X"09",X"22",X"00",
		X"99",X"99",X"99",X"00",X"99",X"91",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"99",X"99",X"00",
		X"00",X"00",X"90",X"00",X"00",X"99",X"C9",X"00",X"00",X"99",X"AC",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"DD",X"00",X"00",X"99",X"99",X"00",X"00",X"C9",X"99",X"00",X"00",X"C9",X"F9",X"00",
		X"00",X"99",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"49",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"C9",X"F9",X"00",X"00",X"C9",X"99",X"00",
		X"00",X"CC",X"99",X"00",X"00",X"CC",X"DD",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"99",X"00",
		X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",
		X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"F9",X"00",X"00",X"09",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"11",X"11",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"9C",X"00",X"00",X"C9",X"CC",X"00",X"00",X"CC",X"CC",X"00",
		X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"C9",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"94",X"00",X"00",X"49",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"99",X"44",X"00",X"00",X"99",X"44",X"00",X"00",X"94",X"44",X"00",X"00",X"94",X"44",X"00",
		X"00",X"44",X"99",X"00",X"00",X"99",X"22",X"00",X"00",X"92",X"22",X"00",X"00",X"92",X"92",X"00",
		X"00",X"92",X"22",X"00",X"00",X"92",X"22",X"00",X"00",X"92",X"22",X"00",X"00",X"99",X"22",X"00",
		X"00",X"99",X"22",X"00",X"00",X"19",X"99",X"00",X"00",X"11",X"11",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"CC",X"00",X"00",X"99",X"9C",X"00",X"00",X"99",X"9C",X"00",
		X"00",X"CC",X"97",X"00",X"00",X"9C",X"99",X"00",X"00",X"CC",X"CC",X"00",X"00",X"9C",X"CC",X"00",
		X"00",X"CC",X"C9",X"00",X"00",X"CC",X"94",X"00",X"00",X"CC",X"94",X"00",X"00",X"CC",X"94",X"00",
		X"00",X"C9",X"49",X"00",X"00",X"CC",X"49",X"00",X"00",X"99",X"99",X"00",X"09",X"44",X"90",X"00",
		X"99",X"44",X"00",X"00",X"94",X"44",X"99",X"00",X"49",X"44",X"49",X"00",X"44",X"44",X"44",X"00",
		X"CC",X"44",X"44",X"00",X"C9",X"94",X"49",X"00",X"99",X"99",X"99",X"00",X"00",X"22",X"91",X"00",
		X"00",X"22",X"91",X"00",X"00",X"92",X"91",X"00",X"00",X"99",X"91",X"00",X"00",X"09",X"91",X"00",
		X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"99",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"CC",X"90",X"00",X"00",X"9C",X"99",X"00",X"00",X"CC",X"CC",X"00",X"00",X"9C",X"CC",X"00",
		X"00",X"CC",X"C9",X"00",X"00",X"CC",X"90",X"00",X"00",X"C9",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"C9",X"00",X"90",X"00",X"CC",X"99",X"99",X"00",X"99",X"44",X"CC",X"00",X"44",X"94",X"C9",
		X"00",X"44",X"99",X"99",X"00",X"44",X"99",X"00",X"00",X"44",X"49",X"90",X"00",X"99",X"44",X"90",
		X"00",X"11",X"44",X"90",X"00",X"11",X"49",X"90",X"00",X"11",X"99",X"90",X"99",X"11",X"22",X"90",
		X"CC",X"11",X"22",X"90",X"CC",X"11",X"99",X"90",X"99",X"99",X"00",X"00",X"09",X"11",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"CC",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"C9",X"00",X"00",X"CC",X"C9",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"94",X"00",X"00",X"99",X"99",X"00",X"00",X"94",X"99",X"00",
		X"00",X"94",X"94",X"00",X"00",X"99",X"44",X"00",X"00",X"CC",X"99",X"00",X"00",X"99",X"90",X"00",
		X"00",X"44",X"90",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"49",X"90",X"00",X"99",X"44",X"90",
		X"00",X"11",X"44",X"90",X"00",X"11",X"49",X"90",X"00",X"11",X"99",X"90",X"99",X"11",X"22",X"90",
		X"CC",X"11",X"22",X"90",X"CC",X"11",X"99",X"90",X"99",X"99",X"00",X"00",X"09",X"11",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9F",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9D",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"9F",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9D",X"00",X"00",X"00",
		X"D9",X"00",X"00",X"00",X"D9",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"9F",X"00",X"00",X"99",X"D9",X"00",X"00",X"09",X"9D",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"F9",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"D9",X"00",X"00",X"09",X"9D",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"09",X"99",X"99",X"00",
		X"99",X"9F",X"99",X"00",X"DD",X"DD",X"DD",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"90",X"00",X"00",X"DD",X"D0",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"DD",X"90",X"00",
		X"00",X"9D",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"09",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"D9",X"00",X"00",
		X"09",X"D9",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"D9",X"00",X"00",X"00",X"9D",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"9F",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"9D",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"D9",X"00",X"00",X"00",X"9D",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",
		X"00",X"00",X"99",X"D9",X"00",X"09",X"99",X"99",X"00",X"99",X"DD",X"99",X"00",X"99",X"9D",X"99",
		X"00",X"D9",X"99",X"99",X"00",X"DD",X"99",X"99",X"00",X"9D",X"9D",X"90",X"00",X"99",X"DD",X"00",
		X"00",X"99",X"D9",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"09",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"DD",X"DD",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"F9",X"F9",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"F9",X"F9",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"DD",X"DD",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"F9",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"F9",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"DD",X"DD",X"00",X"00",
		X"99",X"99",X"00",X"00",X"FF",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"9D",X"DD",X"00",X"00",X"99",X"99",X"00",X"00",
		X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"F9",X"00",X"00",X"99",X"99",X"00",X"00",X"DD",X"DD",X"00",X"00",
		X"9F",X"9F",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"DD",X"DD",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"9D",X"DD",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"DD",X"DD",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"C9",X"C9",X"00",
		X"00",X"CC",X"C9",X"00",X"00",X"99",X"9C",X"00",X"00",X"99",X"99",X"00",X"00",X"2A",X"AE",X"00",
		X"00",X"22",X"2E",X"00",X"00",X"CC",X"CC",X"00",X"00",X"C9",X"CC",X"00",X"00",X"CC",X"CC",X"90",
		X"09",X"CC",X"CC",X"90",X"99",X"99",X"CC",X"99",X"99",X"F9",X"9C",X"99",X"99",X"99",X"9C",X"99",
		X"99",X"9F",X"CC",X"99",X"99",X"99",X"C9",X"99",X"99",X"CC",X"C9",X"99",X"99",X"CC",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"C9",X"C9",X"99",X"99",X"CE",X"EC",X"99",X"99",X"EE",
		X"EE",X"94",X"99",X"CC",X"EC",X"94",X"99",X"EE",X"CE",X"94",X"99",X"CC",X"EC",X"99",X"99",X"EC",
		X"EE",X"99",X"99",X"CC",X"EC",X"99",X"99",X"C9",X"CE",X"99",X"99",X"C9",X"EC",X"9C",X"CC",X"99",
		X"EE",X"CC",X"CC",X"90",X"CC",X"99",X"CC",X"90",X"CE",X"CC",X"EC",X"00",X"CC",X"CC",X"CE",X"00",
		X"CC",X"CC",X"99",X"00",X"CC",X"99",X"BB",X"00",X"C9",X"BB",X"BB",X"00",X"C9",X"BB",X"BB",X"00",
		X"C9",X"BB",X"BB",X"00",X"C9",X"BB",X"BB",X"00",X"99",X"BB",X"BB",X"00",X"99",X"BB",X"BB",X"00",
		X"9B",X"BB",X"BB",X"00",X"9B",X"B9",X"BB",X"00",X"99",X"B9",X"BB",X"00",X"09",X"B9",X"BB",X"00",
		X"99",X"B9",X"BB",X"00",X"99",X"99",X"BB",X"00",X"99",X"99",X"BB",X"00",X"97",X"79",X"BB",X"00",
		X"97",X"79",X"BB",X"00",X"97",X"79",X"BB",X"00",X"99",X"99",X"BB",X"00",X"99",X"99",X"BB",X"00",
		X"09",X"90",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"E7",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"90",X"00",X"99",X"00",X"99",X"00",
		X"95",X"99",X"59",X"00",X"55",X"59",X"59",X"00",X"57",X"25",X"59",X"00",X"97",X"9E",X"99",X"00",
		X"99",X"2E",X"90",X"00",X"55",X"E5",X"00",X"00",X"55",X"55",X"99",X"00",X"55",X"55",X"55",X"00",
		X"55",X"95",X"99",X"99",X"55",X"45",X"99",X"59",X"55",X"44",X"99",X"55",X"55",X"44",X"59",X"95",
		X"59",X"45",X"55",X"95",X"99",X"55",X"55",X"95",X"00",X"55",X"55",X"95",X"00",X"55",X"55",X"95",
		X"00",X"55",X"55",X"99",X"00",X"99",X"55",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",
		X"00",X"99",X"95",X"00",X"00",X"97",X"55",X"00",X"00",X"99",X"55",X"00",X"00",X"59",X"59",X"00",
		X"00",X"55",X"99",X"00",X"00",X"55",X"99",X"00",X"00",X"95",X"09",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",
		X"99",X"59",X"00",X"00",X"95",X"25",X"00",X"00",X"57",X"25",X"00",X"99",X"99",X"25",X"00",X"95",
		X"55",X"55",X"00",X"95",X"55",X"59",X"00",X"95",X"55",X"59",X"99",X"95",X"55",X"59",X"55",X"95",
		X"55",X"59",X"55",X"55",X"55",X"59",X"99",X"59",X"55",X"59",X"99",X"99",X"59",X"55",X"99",X"00",
		X"99",X"95",X"59",X"00",X"00",X"55",X"55",X"00",X"00",X"55",X"55",X"99",X"99",X"55",X"55",X"79",
		X"97",X"95",X"55",X"97",X"77",X"99",X"55",X"99",X"99",X"09",X"99",X"59",X"99",X"00",X"00",X"55",
		X"95",X"00",X"00",X"55",X"55",X"00",X"00",X"55",X"59",X"00",X"00",X"55",X"59",X"00",X"00",X"55",
		X"99",X"00",X"00",X"59",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"CC",X"A9",X"00",X"00",X"C9",X"A9",X"00",X"00",X"CC",X"9C",X"00",X"00",X"99",X"CC",X"00",
		X"00",X"CC",X"CC",X"00",X"00",X"44",X"99",X"00",X"00",X"C9",X"99",X"00",X"00",X"CC",X"99",X"00",
		X"00",X"CC",X"90",X"00",X"00",X"9C",X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"99",X"99",X"00",
		X"99",X"49",X"99",X"90",X"9F",X"44",X"99",X"90",X"99",X"44",X"49",X"90",X"99",X"94",X"44",X"90",
		X"99",X"99",X"44",X"90",X"99",X"99",X"99",X"90",X"99",X"22",X"22",X"90",X"99",X"22",X"29",X"90",
		X"9F",X"92",X"29",X"90",X"99",X"99",X"99",X"90",X"99",X"29",X"99",X"90",X"99",X"99",X"99",X"00",
		X"00",X"19",X"99",X"00",X"00",X"19",X"11",X"00",X"00",X"19",X"11",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"C9",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"C9",X"CC",X"00",X"00",X"9C",X"CC",X"00",
		X"00",X"CC",X"C9",X"00",X"00",X"44",X"99",X"00",X"00",X"C9",X"90",X"00",X"00",X"CC",X"90",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"99",X"99",X"99",X"00",X"99",X"49",X"99",X"00",
		X"94",X"44",X"99",X"00",X"44",X"44",X"99",X"00",X"44",X"44",X"49",X"00",X"99",X"44",X"44",X"00",
		X"44",X"44",X"44",X"00",X"99",X"99",X"99",X"90",X"CC",X"99",X"29",X"90",X"CC",X"99",X"22",X"90",
		X"99",X"29",X"22",X"90",X"99",X"22",X"92",X"00",X"99",X"22",X"22",X"00",X"00",X"99",X"92",X"00",
		X"00",X"90",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"99",X"99",X"90",X"00",
		X"C9",X"C9",X"90",X"00",X"C9",X"99",X"99",X"00",X"99",X"C9",X"CC",X"00",X"99",X"9C",X"CC",X"00",
		X"44",X"CC",X"C9",X"00",X"44",X"44",X"99",X"00",X"44",X"C9",X"90",X"00",X"94",X"CC",X"90",X"00",
		X"99",X"CC",X"00",X"00",X"09",X"9C",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"49",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"44",X"90",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"49",X"00",
		X"00",X"44",X"49",X"00",X"00",X"99",X"99",X"90",X"00",X"99",X"29",X"90",X"00",X"99",X"22",X"90",
		X"00",X"29",X"22",X"90",X"00",X"22",X"92",X"00",X"00",X"22",X"22",X"00",X"00",X"99",X"92",X"00",
		X"00",X"90",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"99",X"00",X"00",
		X"05",X"99",X"90",X"00",X"05",X"99",X"99",X"55",X"55",X"99",X"99",X"50",X"50",X"C9",X"C9",X"00",
		X"00",X"CC",X"C9",X"00",X"00",X"9F",X"9C",X"00",X"A0",X"9F",X"F9",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"99",X"99",X"00",X"00",X"CC",X"9C",X"00",
		X"09",X"CC",X"C9",X"00",X"99",X"CC",X"C9",X"90",X"99",X"9C",X"99",X"90",X"99",X"99",X"99",X"99",
		X"99",X"99",X"9C",X"99",X"99",X"CC",X"99",X"99",X"99",X"CC",X"49",X"99",X"99",X"CC",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"CC",X"99",X"99",X"CE",X"EC",X"99",X"99",X"EE",
		X"CC",X"94",X"99",X"CC",X"EC",X"94",X"99",X"EE",X"99",X"94",X"99",X"99",X"09",X"99",X"99",X"09",
		X"00",X"00",X"99",X"90",X"90",X"00",X"00",X"00",X"99",X"09",X"00",X"00",X"00",X"09",X"09",X"90",
		X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"49",X"49",X"00",
		X"00",X"44",X"49",X"00",X"00",X"99",X"94",X"00",X"00",X"9A",X"99",X"00",X"00",X"A9",X"A9",X"00",
		X"00",X"AA",X"AA",X"00",X"00",X"A4",X"AA",X"00",X"00",X"49",X"44",X"00",X"00",X"44",X"49",X"90",
		X"09",X"94",X"99",X"90",X"99",X"99",X"F9",X"99",X"99",X"FF",X"99",X"99",X"99",X"99",X"94",X"99",
		X"99",X"FF",X"44",X"99",X"99",X"9F",X"49",X"99",X"99",X"49",X"49",X"99",X"99",X"44",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"C9",X"C9",X"99",X"99",X"CE",X"EC",X"99",X"99",X"EE",
		X"EE",X"94",X"99",X"CC",X"EC",X"94",X"99",X"EE",X"CE",X"94",X"99",X"CC",X"EC",X"99",X"99",X"EC",
		X"EE",X"99",X"99",X"CC",X"EC",X"99",X"99",X"C9",X"CE",X"99",X"99",X"C9",X"EC",X"9C",X"CC",X"99",
		X"EE",X"CC",X"CC",X"90",X"CC",X"99",X"CC",X"90",X"CC",X"CC",X"EC",X"00",X"CC",X"CC",X"CE",X"00",
		X"CC",X"CC",X"99",X"00",X"CC",X"99",X"4F",X"00",X"C9",X"F4",X"4F",X"00",X"C9",X"FF",X"FF",X"00",
		X"C9",X"4F",X"44",X"00",X"C9",X"49",X"44",X"00",X"99",X"FF",X"FF",X"00",X"F9",X"FF",X"FF",X"00",
		X"99",X"99",X"99",X"00",X"9E",X"EC",X"EE",X"00",X"9C",X"CC",X"CC",X"00",X"99",X"EE",X"CE",X"00",
		X"09",X"CE",X"EE",X"00",X"00",X"EC",X"CC",X"00",X"00",X"CE",X"CE",X"00",X"00",X"EC",X"EC",X"00",
		X"09",X"C9",X"CE",X"90",X"99",X"99",X"EC",X"90",X"B1",X"90",X"9C",X"99",X"BB",X"90",X"99",X"B9",
		X"BB",X"99",X"00",X"99",X"BB",X"B9",X"99",X"1B",X"9B",X"99",X"BB",X"BB",X"99",X"9B",X"BB",X"BB",
		X"99",X"BB",X"BB",X"B9",X"99",X"B9",X"99",X"B9",X"BB",X"99",X"99",X"99",X"99",X"BB",X"BB",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"09",X"77",
		X"00",X"00",X"99",X"77",X"99",X"00",X"9E",X"99",X"9C",X"00",X"EE",X"BB",X"9C",X"00",X"EE",X"BB",
		X"9C",X"99",X"EE",X"BB",X"9C",X"97",X"99",X"99",X"9C",X"99",X"45",X"45",X"9C",X"90",X"45",X"45",
		X"9C",X"00",X"45",X"45",X"99",X"00",X"45",X"45",X"09",X"00",X"45",X"45",X"09",X"00",X"45",X"45",
		X"09",X"00",X"45",X"45",X"09",X"00",X"45",X"45",X"99",X"00",X"45",X"45",X"96",X"00",X"47",X"45",
		X"99",X"00",X"47",X"47",X"9A",X"00",X"47",X"49",X"9A",X"00",X"47",X"99",X"99",X"00",X"99",X"90",
		X"09",X"00",X"95",X"90",X"99",X"00",X"99",X"00",X"9A",X"00",X"99",X"00",X"9A",X"00",X"90",X"99",
		X"9A",X"00",X"99",X"AB",X"99",X"00",X"A9",X"55",X"99",X"00",X"99",X"BB",X"99",X"00",X"90",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"09",X"77",
		X"00",X"00",X"99",X"77",X"99",X"00",X"9E",X"99",X"9C",X"00",X"EE",X"BB",X"9C",X"00",X"EE",X"BB",
		X"9C",X"99",X"99",X"99",X"9C",X"97",X"45",X"45",X"9C",X"99",X"45",X"45",X"9C",X"90",X"45",X"45",
		X"9C",X"00",X"45",X"45",X"99",X"00",X"45",X"45",X"09",X"00",X"45",X"45",X"09",X"00",X"45",X"45",
		X"09",X"00",X"45",X"45",X"09",X"00",X"45",X"45",X"09",X"00",X"47",X"45",X"99",X"00",X"47",X"47",
		X"96",X"00",X"47",X"49",X"99",X"00",X"47",X"99",X"AA",X"00",X"99",X"90",X"9A",X"00",X"95",X"00",
		X"99",X"00",X"99",X"00",X"99",X"99",X"09",X"00",X"29",X"A9",X"99",X"90",X"22",X"A9",X"B9",X"99",
		X"29",X"99",X"5B",X"B9",X"99",X"99",X"5B",X"A9",X"99",X"99",X"A9",X"99",X"99",X"90",X"99",X"90",
		X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"94",X"99",X"00",
		X"00",X"44",X"49",X"00",X"00",X"44",X"CC",X"00",X"00",X"44",X"CC",X"00",X"00",X"44",X"99",X"00",
		X"00",X"4C",X"C9",X"00",X"00",X"4C",X"C9",X"00",X"00",X"49",X"C9",X"00",X"09",X"99",X"99",X"00",
		X"99",X"AA",X"9A",X"90",X"9C",X"AA",X"AA",X"99",X"CC",X"AA",X"AA",X"C9",X"CC",X"99",X"99",X"CC",
		X"CC",X"99",X"99",X"CC",X"CC",X"AA",X"AA",X"CC",X"99",X"AA",X"AA",X"C9",X"00",X"AA",X"AA",X"99",
		X"99",X"AA",X"AA",X"44",X"55",X"22",X"22",X"99",X"55",X"AA",X"AA",X"55",X"55",X"99",X"99",X"55",
		X"45",X"CC",X"CC",X"55",X"45",X"99",X"CC",X"54",X"45",X"90",X"CC",X"54",X"55",X"99",X"CC",X"54",
		X"55",X"29",X"CC",X"55",X"99",X"99",X"99",X"99",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"94",X"99",X"00",
		X"00",X"4A",X"49",X"00",X"00",X"C2",X"44",X"00",X"00",X"CC",X"44",X"00",X"00",X"9C",X"44",X"00",
		X"00",X"C4",X"44",X"00",X"00",X"C9",X"44",X"00",X"09",X"C4",X"44",X"00",X"99",X"9C",X"99",X"90",
		X"9C",X"99",X"AA",X"99",X"CC",X"AA",X"AA",X"C9",X"CC",X"AA",X"AA",X"CC",X"CC",X"AA",X"AA",X"CC",
		X"CC",X"99",X"99",X"CC",X"99",X"AA",X"99",X"C9",X"00",X"AA",X"AA",X"99",X"99",X"AA",X"AA",X"44",
		X"55",X"AA",X"AA",X"99",X"55",X"22",X"22",X"55",X"55",X"AA",X"AA",X"55",X"45",X"99",X"99",X"54",
		X"45",X"C9",X"CC",X"54",X"45",X"C9",X"9C",X"54",X"55",X"C9",X"9C",X"55",X"55",X"C9",X"99",X"55",
		X"99",X"C9",X"22",X"99",X"00",X"99",X"99",X"00",X"00",X"29",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"94",X"99",X"00",
		X"00",X"44",X"49",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"49",X"00",
		X"00",X"94",X"99",X"00",X"09",X"99",X"9A",X"00",X"99",X"99",X"AA",X"00",X"9C",X"A9",X"AA",X"90",
		X"CC",X"AA",X"AA",X"99",X"CC",X"AA",X"AA",X"C9",X"9C",X"AA",X"AA",X"CC",X"CC",X"AA",X"AA",X"99",
		X"CC",X"A9",X"9A",X"CC",X"99",X"99",X"99",X"C9",X"00",X"AA",X"AA",X"99",X"99",X"AA",X"AA",X"00",
		X"55",X"AA",X"AA",X"99",X"55",X"AA",X"AA",X"55",X"55",X"AA",X"AA",X"55",X"45",X"99",X"99",X"55",
		X"45",X"C9",X"CC",X"54",X"45",X"C9",X"9C",X"54",X"55",X"C9",X"9C",X"54",X"55",X"C9",X"99",X"55",
		X"99",X"C9",X"22",X"55",X"00",X"99",X"99",X"99",X"00",X"29",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"55",X"99",X"00",X"00",X"99",X"55",X"00",
		X"00",X"9F",X"95",X"00",X"00",X"FF",X"95",X"00",X"00",X"FF",X"99",X"00",X"00",X"FF",X"F9",X"00",
		X"00",X"FF",X"FF",X"00",X"00",X"99",X"FF",X"00",X"00",X"99",X"FF",X"00",X"00",X"F9",X"FF",X"00",
		X"00",X"FF",X"FF",X"00",X"00",X"FF",X"F9",X"00",X"00",X"FF",X"F9",X"90",X"00",X"FF",X"95",X"90",
		X"00",X"FF",X"95",X"90",X"00",X"9F",X"55",X"90",X"00",X"99",X"59",X"90",X"00",X"55",X"99",X"90",
		X"00",X"99",X"99",X"90",X"00",X"99",X"99",X"90",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"AA",X"00",X"00",X"00",X"D9",X"09",X"00",X"00",X"CC",X"09",X"00",X"00",X"9C",X"09",X"00",
		X"9D",X"99",X"99",X"00",X"9D",X"C4",X"93",X"00",X"90",X"CC",X"33",X"00",X"90",X"9C",X"33",X"00",
		X"99",X"99",X"99",X"00",X"95",X"33",X"29",X"00",X"55",X"93",X"29",X"00",X"55",X"99",X"29",X"00",
		X"55",X"99",X"99",X"00",X"55",X"99",X"96",X"00",X"55",X"99",X"66",X"00",X"99",X"33",X"66",X"90",
		X"66",X"99",X"66",X"99",X"22",X"22",X"22",X"55",X"22",X"22",X"22",X"55",X"22",X"22",X"29",X"59",
		X"29",X"92",X"99",X"99",X"99",X"99",X"97",X"96",X"97",X"79",X"77",X"96",X"97",X"79",X"75",X"96",
		X"97",X"79",X"77",X"99",X"99",X"99",X"97",X"90",X"09",X"90",X"99",X"00",X"00",X"00",X"09",X"00",
		X"00",X"99",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"99",X"00",X"00",X"99",X"94",X"00",
		X"00",X"A9",X"44",X"00",X"00",X"CC",X"99",X"00",X"00",X"9C",X"9C",X"00",X"00",X"99",X"CC",X"00",
		X"9D",X"44",X"C9",X"00",X"9D",X"99",X"9C",X"00",X"90",X"CC",X"99",X"00",X"90",X"CC",X"90",X"00",
		X"90",X"99",X"90",X"00",X"99",X"33",X"99",X"00",X"95",X"93",X"29",X"00",X"55",X"99",X"29",X"00",
		X"55",X"99",X"A9",X"00",X"55",X"99",X"99",X"00",X"55",X"99",X"96",X"00",X"55",X"33",X"66",X"00",
		X"99",X"33",X"66",X"90",X"66",X"99",X"66",X"99",X"22",X"22",X"29",X"55",X"29",X"22",X"99",X"55",
		X"99",X"92",X"97",X"59",X"97",X"92",X"77",X"99",X"97",X"96",X"77",X"96",X"97",X"96",X"77",X"96",
		X"95",X"96",X"77",X"96",X"99",X"99",X"97",X"99",X"09",X"00",X"99",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"99",X"EE",X"00",X"00",X"EE",X"AE",X"00",X"00",X"99",X"EE",X"00",X"00",X"EE",X"EE",X"00",
		X"00",X"EE",X"9E",X"00",X"00",X"EE",X"9E",X"00",X"00",X"EE",X"99",X"00",X"00",X"E9",X"E9",X"00",
		X"09",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"9E",X"90",X"99",X"00",X"99",X"00",X"99",X"00",
		X"09",X"00",X"99",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"99",X"00",X"09",X"99",X"EE",X"00",
		X"09",X"EE",X"AE",X"00",X"00",X"99",X"AE",X"00",X"00",X"9E",X"EE",X"00",X"00",X"EE",X"9E",X"00",
		X"00",X"EE",X"9E",X"00",X"00",X"EE",X"99",X"00",X"00",X"EE",X"E9",X"00",X"00",X"9E",X"99",X"00",
		X"00",X"99",X"09",X"00",X"00",X"EE",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"EA",X"00",X"00",X"00",X"EA",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"E9",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"E9",X"00",X"00",
		X"00",X"E9",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"9E",X"00",X"00",
		X"99",X"99",X"00",X"00",X"9E",X"9E",X"00",X"00",X"9E",X"EE",X"00",X"00",X"99",X"EE",X"00",X"00",
		X"09",X"99",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"00",X"00",X"99",X"94",X"00",X"00",X"09",X"09",X"00",X"00",X"00",X"00",X"90",
		X"00",X"09",X"00",X"99",X"99",X"99",X"90",X"A9",X"9A",X"9D",X"99",X"A9",X"AA",X"99",X"99",X"9A",
		X"AA",X"99",X"92",X"AA",X"99",X"99",X"99",X"99",X"AA",X"95",X"90",X"90",X"AA",X"99",X"90",X"00",
		X"99",X"99",X"90",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"94",X"90",X"00",X"00",X"44",X"99",X"00",X"FF",X"99",X"49",X"00",
		X"00",X"C9",X"C9",X"00",X"00",X"C9",X"99",X"00",X"00",X"CC",X"90",X"00",X"00",X"94",X"90",X"00",
		X"00",X"9C",X"99",X"00",X"00",X"99",X"59",X"00",X"00",X"55",X"55",X"00",X"00",X"55",X"55",X"00",
		X"00",X"99",X"99",X"00",X"00",X"59",X"99",X"00",X"00",X"55",X"99",X"00",X"00",X"55",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"22",X"90",X"00",X"00",X"22",X"90",X"00",
		X"00",X"22",X"90",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"99",X"00",
		X"00",X"09",X"9E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"9E",X"00",
		X"00",X"00",X"9E",X"00",X"00",X"00",X"99",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"94",X"90",X"00",X"00",X"44",X"90",X"00",
		X"00",X"49",X"90",X"00",X"00",X"94",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"95",X"00",X"00",X"79",X"97",X"00",X"00",X"79",X"57",X"00",
		X"00",X"99",X"79",X"00",X"00",X"77",X"79",X"00",X"00",X"77",X"99",X"00",X"00",X"97",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"22",X"90",X"00",X"00",X"22",X"90",X"00",
		X"00",X"22",X"90",X"00",X"00",X"92",X"90",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"92",X"99",X"00",X"00",X"22",X"9E",X"00",
		X"00",X"99",X"9E",X"00",X"00",X"90",X"9E",X"00",X"00",X"90",X"EE",X"00",X"00",X"90",X"99",X"00",
		X"99",X"99",X"00",X"00",X"CC",X"44",X"00",X"00",X"CC",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"9C",X"00",X"00",X"99",X"9C",X"00",X"00",X"29",X"CC",X"00",X"00",X"29",X"99",X"00",X"00",
		X"29",X"CC",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"CC",X"90",X"00",X"99",X"99",X"90",X"00",
		X"99",X"22",X"90",X"00",X"99",X"22",X"90",X"00",X"00",X"22",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"22",X"90",X"00",X"00",X"22",X"90",X"00",X"00",X"22",X"90",X"00",X"00",X"22",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"66",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",
		X"00",X"09",X"90",X"00",X"00",X"99",X"99",X"00",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"90",X"94",X"9C",X"90",X"90",X"94",X"9C",X"90",X"90",X"94",X"99",X"90",X"90",X"99",X"90",X"90",
		X"90",X"99",X"90",X"90",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"00",X"09",X"90",X"00",
		X"00",X"09",X"90",X"00",X"00",X"09",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"92",X"92",X"00",X"00",X"92",X"22",X"00",X"00",X"92",X"29",X"00",X"00",X"92",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"96",X"99",X"09",X"00",X"99",X"99",X"99",X"00",X"99",X"90",X"11",
		X"00",X"66",X"90",X"11",X"00",X"66",X"90",X"19",X"00",X"99",X"00",X"19",X"00",X"99",X"00",X"90",
		X"00",X"19",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"90",X"00",X"09",X"49",X"90",X"00",X"09",X"44",X"90",X"00",X"99",X"44",X"99",
		X"00",X"94",X"44",X"99",X"00",X"94",X"94",X"99",X"00",X"94",X"44",X"99",X"00",X"99",X"99",X"90",
		X"00",X"09",X"9C",X"90",X"00",X"09",X"CC",X"99",X"00",X"99",X"99",X"99",X"00",X"29",X"92",X"99",
		X"00",X"29",X"29",X"99",X"00",X"99",X"22",X"99",X"00",X"92",X"22",X"00",X"00",X"22",X"22",X"00",
		X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"92",X"22",X"00",X"00",X"99",X"29",X"00",
		X"00",X"99",X"99",X"00",X"00",X"96",X"66",X"00",X"00",X"96",X"99",X"00",X"00",X"99",X"66",X"00",
		X"00",X"09",X"69",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"99",X"00",
		X"00",X"99",X"91",X"00",X"00",X"91",X"91",X"00",X"00",X"11",X"99",X"00",X"00",X"99",X"09",X"00",
		X"00",X"99",X"00",X"00",X"00",X"44",X"00",X"00",X"99",X"99",X"99",X"99",X"99",X"C9",X"99",X"99",
		X"00",X"C9",X"90",X"00",X"00",X"C9",X"90",X"00",X"00",X"9C",X"90",X"00",X"00",X"CC",X"90",X"00",
		X"00",X"49",X"90",X"00",X"99",X"9C",X"99",X"99",X"99",X"99",X"99",X"99",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",
		X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"00",X"79",X"00",X"94",X"00",X"79",X"00",X"44",X"90",X"AA",X"00",X"44",X"99",X"AA",X"00",
		X"99",X"99",X"97",X"00",X"EE",X"C9",X"97",X"00",X"EE",X"CC",X"97",X"90",X"C4",X"99",X"99",X"99",
		X"C4",X"00",X"00",X"39",X"CC",X"00",X"99",X"99",X"99",X"00",X"33",X"90",X"55",X"00",X"11",X"00",
		X"55",X"00",X"33",X"00",X"55",X"00",X"99",X"00",X"95",X"90",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"EE",X"00",X"00",X"55",X"CC",X"09",X"99",X"55",X"9C",X"99",X"99",X"55",X"9C",X"77",X"44",
		X"99",X"99",X"77",X"44",X"11",X"00",X"74",X"44",X"11",X"00",X"94",X"44",X"91",X"90",X"99",X"49",
		X"99",X"99",X"09",X"99",X"99",X"11",X"00",X"90",X"19",X"11",X"00",X"00",X"99",X"19",X"00",X"90",
		X"90",X"99",X"00",X"90",X"99",X"99",X"00",X"90",X"99",X"00",X"00",X"90",X"99",X"00",X"00",X"00",
		X"09",X"00",X"00",X"69",X"99",X"00",X"09",X"97",X"94",X"99",X"09",X"77",X"44",X"49",X"09",X"77",
		X"99",X"99",X"09",X"77",X"EE",X"CC",X"09",X"99",X"EE",X"CC",X"09",X"69",X"EC",X"99",X"00",X"69",
		X"CC",X"90",X"00",X"99",X"9C",X"90",X"99",X"09",X"99",X"90",X"33",X"99",X"55",X"00",X"11",X"93",
		X"55",X"00",X"31",X"31",X"95",X"90",X"99",X"99",X"99",X"99",X"00",X"00",X"99",X"EE",X"00",X"90",
		X"55",X"CC",X"99",X"99",X"55",X"9C",X"99",X"99",X"55",X"9C",X"77",X"44",X"99",X"99",X"77",X"44",
		X"11",X"00",X"44",X"44",X"11",X"00",X"94",X"44",X"11",X"00",X"99",X"49",X"99",X"00",X"09",X"99",
		X"19",X"00",X"00",X"90",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"19",X"00",X"00",X"00",
		X"19",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"9C",X"99",X"00",X"00",X"99",X"99",X"00",X"99",X"99",X"CC",X"00",X"9C",X"99",X"9C",X"00",
		X"CC",X"99",X"94",X"00",X"9C",X"99",X"44",X"00",X"99",X"9C",X"9C",X"00",X"00",X"99",X"9C",X"00",
		X"00",X"49",X"C9",X"00",X"00",X"44",X"99",X"00",X"00",X"99",X"94",X"00",X"00",X"99",X"44",X"00",
		X"00",X"99",X"49",X"00",X"00",X"94",X"99",X"00",X"00",X"94",X"44",X"00",X"00",X"94",X"44",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"92",X"00",X"00",X"92",X"22",X"00",X"00",X"92",X"22",X"00",
		X"00",X"22",X"22",X"00",X"00",X"22",X"92",X"00",X"00",X"22",X"29",X"00",X"00",X"92",X"22",X"00",
		X"00",X"99",X"99",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"99",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"94",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"A9",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"C9",X"00",X"00",X"00",X"CC",X"90",X"00",X"00",X"49",X"99",X"00",
		X"00",X"9C",X"79",X"00",X"00",X"99",X"79",X"00",X"00",X"97",X"99",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"99",X"00",X"99",X"CC",X"99",X"00",X"49",X"CC",X"79",X"00",X"00",X"99",X"99",X"00",
		X"00",X"09",X"D9",X"00",X"00",X"09",X"D9",X"00",X"00",X"09",X"D9",X"00",X"00",X"09",X"99",X"00",
		X"00",X"00",X"9D",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"DD",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
