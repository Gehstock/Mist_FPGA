library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity kbe1_IC4 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of kbe1_IC4 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"21",X"FF",X"FF",X"2D",X"20",X"FD",X"25",X"20",X"FA",X"DB",X"00",X"FE",X"F0",X"28",X"FA",X"3E",
		X"10",X"3D",X"20",X"FD",X"DB",X"00",X"FE",X"F0",X"28",X"EF",X"FE",X"F1",X"20",X"25",X"21",X"80",
		X"01",X"01",X"4F",X"06",X"DD",X"21",X"2A",X"00",X"18",X"4C",X"06",X"02",X"21",X"FF",X"FF",X"2D",
		X"20",X"FD",X"25",X"20",X"05",X"05",X"20",X"02",X"18",X"CF",X"DB",X"00",X"FE",X"F1",X"28",X"EF",
		X"C3",X"09",X"00",X"FE",X"F2",X"C2",X"5B",X"00",X"21",X"50",X"06",X"01",X"8F",X"10",X"DD",X"21",
		X"55",X"00",X"C3",X"76",X"00",X"DB",X"00",X"FE",X"F2",X"28",X"FA",X"FE",X"F3",X"C2",X"09",X"00",
		X"21",X"90",X"10",X"01",X"FF",X"17",X"DD",X"21",X"6D",X"00",X"C3",X"76",X"00",X"DB",X"00",X"FE",
		X"F3",X"28",X"FA",X"C3",X"09",X"00",X"50",X"59",X"7E",X"E6",X"F0",X"D3",X"00",X"3E",X"1B",X"3D",
		X"20",X"FD",X"7E",X"E6",X"0F",X"07",X"07",X"07",X"07",X"D3",X"00",X"3E",X"19",X"3D",X"20",X"FD",
		X"23",X"EB",X"ED",X"52",X"EB",X"20",X"DF",X"DD",X"E9",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",
		X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",
		X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",
		X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",
		X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",
		X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",
		X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",
		X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",
		X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",
		X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",
		X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",
		X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",
		X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",
		X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",
		X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",
		X"88",X"89",X"88",X"88",X"88",X"88",X"88",X"98",X"99",X"99",X"88",X"98",X"88",X"88",X"88",X"88",
		X"89",X"99",X"98",X"98",X"88",X"88",X"87",X"88",X"87",X"78",X"9A",X"AA",X"89",X"88",X"98",X"87",
		X"78",X"78",X"77",X"8B",X"CB",X"87",X"88",X"A8",X"87",X"78",X"87",X"78",X"AC",X"C9",X"87",X"89",
		X"88",X"77",X"87",X"68",X"AD",X"C9",X"87",X"89",X"87",X"67",X"76",X"9C",X"CA",X"77",X"89",X"86",
		X"67",X"77",X"AD",X"C9",X"56",X"99",X"96",X"55",X"6E",X"EC",X"85",X"79",X"87",X"67",X"65",X"EE",
		X"C8",X"37",X"9A",X"75",X"76",X"8F",X"CB",X"53",X"88",X"95",X"56",X"4F",X"FA",X"A1",X"89",X"87",
		X"45",X"4D",X"F8",X"B2",X"5B",X"78",X"45",X"5E",X"F7",X"83",X"5C",X"76",X"65",X"5F",X"F8",X"70",
		X"8A",X"94",X"56",X"6F",X"C8",X"50",X"C7",X"83",X"37",X"DF",X"F8",X"05",X"E7",X"71",X"48",X"FF",
		X"63",X"0D",X"8A",X"51",X"3F",X"F6",X"A0",X"89",X"68",X"32",X"EF",X"4C",X"05",X"B5",X"73",X"3B",
		X"FA",X"D2",X"4D",X"4A",X"41",X"BF",X"FD",X"32",X"F4",X"98",X"0D",X"F0",X"F1",X"3D",X"3C",X"51",
		X"FF",X"3D",X"06",X"94",X"F6",X"0F",X"F9",X"A0",X"A5",X"7F",X"36",X"FF",X"F2",X"5B",X"29",X"F0",
		X"FC",X"0F",X"0E",X"24",X"FA",X"3F",X"FC",X"A0",X"D0",X"5F",X"0F",X"F0",X"F0",X"86",X"3A",X"F4",
		X"FF",X"8A",X"0D",X"26",X"D5",X"F8",X"4E",X"0A",X"46",X"A3",X"FA",X"2E",X"3A",X"83",X"E8",X"CF",
		X"0C",X"65",X"C3",X"BA",X"8F",X"07",X"61",X"B8",X"9D",X"6F",X"07",X"80",X"94",X"9E",X"8F",X"14",
		X"A0",X"C3",X"8B",X"5F",X"F6",X"80",X"F5",X"A8",X"0F",X"F6",X"E0",X"D7",X"6F",X"0F",X"F1",X"F0",
		X"A8",X"5C",X"2F",X"F1",X"E0",X"8C",X"6C",X"0F",X"F1",X"C0",X"AC",X"8B",X"0F",X"F4",X"A0",X"8B",
		X"CB",X"0F",X"F3",X"F0",X"98",X"9E",X"0F",X"F0",X"F0",X"BE",X"3D",X"0F",X"F0",X"F0",X"9F",X"27",
		X"2F",X"F0",X"E0",X"CF",X"A4",X"3F",X"F0",X"E0",X"AF",X"67",X"9F",X"F1",X"D0",X"6F",X"64",X"FF",
		X"F4",X"A0",X"BF",X"20",X"FF",X"07",X"42",X"CF",X"70",X"FF",X"0D",X"20",X"EE",X"70",X"FF",X"00",
		X"25",X"FB",X"43",X"FF",X"00",X"07",X"FD",X"31",X"FF",X"09",X"08",X"FB",X"45",X"FF",X"0F",X"00",
		X"F9",X"18",X"FF",X"0F",X"00",X"F2",X"37",X"FF",X"0F",X"06",X"F7",X"0C",X"FF",X"5F",X"0A",X"F4",
		X"0F",X"FF",X"0F",X"0F",X"F4",X"0F",X"FF",X"5D",X"0F",X"E7",X"0F",X"FF",X"2F",X"00",X"F3",X"0F",
		X"FF",X"7F",X"00",X"D0",X"0F",X"F0",X"0E",X"0D",X"F0",X"0F",X"F0",X"0C",X"0F",X"F0",X"0F",X"F0",
		X"0A",X"0F",X"C3",X"0F",X"F0",X"08",X"0F",X"F0",X"0F",X"F0",X"06",X"0F",X"F0",X"3F",X"F0",X"00",
		X"0F",X"A0",X"7F",X"F0",X"00",X"0F",X"F0",X"FF",X"F0",X"00",X"5F",X"60",X"FF",X"F0",X"40",X"0F",
		X"F0",X"FF",X"F0",X"F0",X"EF",X"00",X"FF",X"00",X"F0",X"0F",X"00",X"FF",X"00",X"F0",X"FF",X"05",
		X"FF",X"00",X"40",X"FF",X"07",X"FF",X"00",X"A0",X"FF",X"00",X"FF",X"00",X"01",X"F1",X"0F",X"FF",
		X"00",X"01",X"FF",X"00",X"FF",X"0F",X"06",X"F3",X"0F",X"FF",X"0F",X"00",X"F0",X"0F",X"FF",X"0F",
		X"FB",X"F0",X"0F",X"F0",X"0F",X"00",X"F0",X"0F",X"F0",X"0F",X"0F",X"F0",X"1F",X"F0",X"0D",X"0F",
		X"E0",X"5F",X"F0",X"0F",X"00",X"F0",X"0F",X"F0",X"0F",X"0F",X"F0",X"AF",X"F0",X"0F",X"0F",X"90",
		X"0F",X"F0",X"0E",X"0F",X"A0",X"0F",X"F0",X"0E",X"0F",X"E0",X"0F",X"F0",X"04",X"0F",X"E0",X"FF",
		X"F0",X"0D",X"0E",X"F0",X"BF",X"F0",X"0C",X"2F",X"F0",X"5F",X"F0",X"87",X"1C",X"F0",X"AF",X"F0",
		X"CD",X"2B",X"C0",X"3F",X"F0",X"08",X"AB",X"E2",X"1F",X"F6",X"61",X"1E",X"F2",X"6F",X"B0",X"5A",
		X"4A",X"F1",X"1F",X"F6",X"02",X"DE",X"B4",X"4F",X"FC",X"30",X"4D",X"E4",X"7F",X"F7",X"03",X"8A",
		X"B8",X"48",X"FF",X"00",X"5F",X"C7",X"76",X"FE",X"33",X"49",X"C8",X"74",X"FF",X"60",X"0D",X"DB",
		X"83",X"BF",X"96",X"27",X"7A",X"A6",X"FF",X"50",X"3C",X"BA",X"64",X"9F",X"FC",X"00",X"8F",X"D3",
		X"AE",X"88",X"57",X"68",X"96",X"8D",X"FD",X"10",X"6F",X"B5",X"93",X"9F",X"F0",X"0A",X"F8",X"88",
		X"CF",X"80",X"2B",X"C4",X"88",X"9F",X"F0",X"0C",X"E5",X"75",X"3F",X"F8",X"01",X"AA",X"B8",X"7F",
		X"F1",X"0A",X"C6",X"78",X"6F",X"F7",X"06",X"A8",X"77",X"6A",X"FF",X"30",X"16",X"B9",X"7D",X"FD",
		X"21",X"57",X"88",X"8C",X"FD",X"66",X"26",X"96",X"8A",X"BE",X"E8",X"03",X"88",X"77",X"DF",X"F9",
		X"02",X"55",X"6A",X"BF",X"FD",X"22",X"55",X"58",X"9C",X"FF",X"63",X"44",X"56",X"6C",X"FF",X"74",
		X"66",X"45",X"56",X"FF",X"BA",X"95",X"56",X"33",X"DD",X"9A",X"C9",X"69",X"42",X"BD",X"86",X"AC",
		X"9A",X"75",X"AA",X"64",X"8A",X"8B",X"A5",X"BB",X"85",X"77",X"59",X"A7",X"BD",X"A7",X"89",X"57",
		X"86",X"AA",X"87",X"B9",X"79",X"A7",X"79",X"75",X"98",X"7A",X"A9",X"9A",X"98",X"A7",X"67",X"79",
		X"9A",X"97",X"BA",X"89",X"89",X"88",X"66",X"A8",X"8A",X"AB",X"99",X"75",X"A8",X"68",X"9B",X"AA",
		X"87",X"B8",X"66",X"79",X"8A",X"87",X"BA",X"88",X"99",X"69",X"85",X"99",X"99",X"BC",X"79",X"85",
		X"88",X"86",X"8B",X"9C",X"95",X"88",X"87",X"99",X"6A",X"A8",X"77",X"87",X"AB",X"8A",X"97",X"77",
		X"76",X"8A",X"8C",X"BA",X"77",X"96",X"78",X"69",X"9A",X"A8",X"87",X"99",X"79",X"AA",X"78",X"86",
		X"79",X"88",X"AB",X"89",X"A9",X"97",X"77",X"88",X"78",X"97",X"AB",X"97",X"9B",X"88",X"86",X"67",
		X"88",X"9A",X"99",X"A8",X"89",X"98",X"99",X"79",X"A7",X"68",X"86",X"8A",X"9A",X"CA",X"98",X"86",
		X"78",X"78",X"A9",X"78",X"98",X"AA",X"77",X"A9",X"88",X"87",X"78",X"68",X"BA",X"99",X"87",X"89",
		X"67",X"AA",X"A9",X"87",X"79",X"88",X"A9",X"99",X"77",X"88",X"67",X"AA",X"AA",X"97",X"77",X"66",
		X"8A",X"BB",X"98",X"87",X"67",X"89",X"BB",X"98",X"87",X"67",X"78",X"AB",X"AA",X"A8",X"67",X"67",
		X"99",X"AA",X"A9",X"78",X"67",X"89",X"99",X"A9",X"89",X"77",X"88",X"88",X"A8",X"89",X"88",X"99",
		X"89",X"98",X"79",X"87",X"88",X"9A",X"A8",X"79",X"88",X"88",X"89",X"A8",X"78",X"88",X"99",X"89",
		X"A8",X"89",X"88",X"88",X"89",X"A9",X"89",X"98",X"77",X"78",X"A9",X"89",X"99",X"98",X"78",X"88",
		X"89",X"98",X"98",X"88",X"88",X"89",X"99",X"98",X"89",X"97",X"79",X"99",X"98",X"89",X"88",X"88",
		X"89",X"97",X"88",X"87",X"8A",X"98",X"99",X"88",X"87",X"89",X"98",X"98",X"99",X"87",X"89",X"98",
		X"88",X"88",X"87",X"89",X"A9",X"A9",X"88",X"66",X"69",X"99",X"9A",X"98",X"76",X"69",X"99",X"89",
		X"A8",X"97",X"7A",X"8A",X"78",X"77",X"98",X"89",X"A9",X"9A",X"88",X"98",X"79",X"87",X"88",X"88",
		X"A9",X"87",X"88",X"89",X"99",X"99",X"78",X"78",X"89",X"99",X"A9",X"88",X"87",X"89",X"98",X"99",
		X"88",X"88",X"8A",X"99",X"99",X"88",X"77",X"78",X"89",X"A9",X"89",X"88",X"88",X"88",X"99",X"89",
		X"88",X"88",X"88",X"99",X"88",X"88",X"88",X"88",X"98",X"89",X"98",X"89",X"89",X"99",X"89",X"97",
		X"88",X"89",X"AA",X"9A",X"98",X"88",X"88",X"98",X"89",X"98",X"89",X"88",X"98",X"89",X"98",X"89",
		X"88",X"88",X"89",X"98",X"88",X"77",X"88",X"88",X"98",X"78",X"87",X"88",X"78",X"99",X"89",X"98",
		X"89",X"88",X"99",X"88",X"99",X"99",X"99",X"99",X"88",X"87",X"88",X"88",X"88",X"88",X"88",X"88",
		X"98",X"89",X"88",X"98",X"78",X"88",X"88",X"88",X"77",X"77",X"88",X"79",X"98",X"99",X"99",X"AA",
		X"9A",X"AA",X"AA",X"AA",X"A9",X"99",X"98",X"98",X"88",X"88",X"78",X"87",X"78",X"78",X"88",X"78",
		X"98",X"89",X"99",X"AA",X"AB",X"BA",X"AA",X"AA",X"AA",X"AA",X"A9",X"99",X"88",X"87",X"66",X"54",
		X"45",X"34",X"43",X"34",X"44",X"56",X"67",X"89",X"9A",X"BB",X"BB",X"BB",X"AA",X"AB",X"A9",X"99",
		X"99",X"99",X"89",X"98",X"77",X"88",X"88",X"99",X"AA",X"AA",X"AA",X"AA",X"AA",X"BA",X"AA",X"AA",
		X"A9",X"AA",X"A9",X"99",X"99",X"87",X"78",X"87",X"66",X"66",X"66",X"66",X"66",X"66",X"67",X"78",
		X"88",X"88",X"88",X"99",X"99",X"99",X"99",X"88",X"89",X"88",X"88",X"89",X"88",X"88",X"88",X"99",
		X"9A",X"AA",X"AA",X"AA",X"AA",X"9A",X"A9",X"99",X"98",X"88",X"77",X"77",X"76",X"66",X"66",X"66",
		X"66",X"77",X"77",X"88",X"88",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"99",X"98",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"78",X"87",X"88",X"77",X"77",X"77",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"9A",X"AB",X"A9",X"88",X"78",X"89",X"99",X"98",X"87",X"77",
		X"78",X"88",X"87",X"77",X"77",X"76",X"8C",X"BD",X"C9",X"87",X"67",X"89",X"AA",X"99",X"77",X"77",
		X"89",X"99",X"98",X"88",X"88",X"88",X"88",X"87",X"77",X"77",X"79",X"DD",X"DC",X"87",X"66",X"8A",
		X"AA",X"98",X"87",X"78",X"89",X"99",X"98",X"88",X"88",X"88",X"87",X"77",X"77",X"66",X"9D",X"DC",
		X"C7",X"66",X"69",X"BB",X"A9",X"77",X"67",X"89",X"9A",X"98",X"87",X"77",X"78",X"87",X"66",X"66",
		X"7B",X"FB",X"E8",X"56",X"78",X"CB",X"B9",X"66",X"77",X"9A",X"9A",X"A9",X"87",X"67",X"78",X"87",
		X"55",X"58",X"EF",X"BD",X"66",X"78",X"AB",X"98",X"87",X"98",X"98",X"88",X"A8",X"98",X"77",X"66",
		X"55",X"56",X"8F",X"CB",X"A4",X"7A",X"8D",X"B8",X"86",X"6A",X"88",X"9A",X"89",X"76",X"65",X"66",
		X"65",X"8C",X"F7",X"E4",X"69",X"7C",X"C8",X"98",X"6C",X"7A",X"A6",X"97",X"77",X"55",X"45",X"7B",
		X"F8",X"D5",X"28",X"79",X"E8",X"BA",X"6A",X"87",X"86",X"88",X"66",X"44",X"49",X"FF",X"9D",X"06",
		X"67",X"DA",X"BB",X"8A",X"85",X"93",X"85",X"57",X"36",X"9F",X"FB",X"C1",X"66",X"6D",X"9C",X"A7",
		X"B7",X"78",X"56",X"44",X"46",X"CF",X"CD",X"71",X"85",X"9D",X"DE",X"97",X"63",X"84",X"75",X"35",
		X"5C",X"F8",X"F5",X"5A",X"3B",X"BB",X"E6",X"A4",X"57",X"43",X"12",X"7D",X"F9",X"F4",X"5A",X"4D",
		X"AA",X"C9",X"96",X"75",X"31",X"05",X"BF",X"D9",X"80",X"B5",X"DF",X"8D",X"89",X"45",X"43",X"21",
		X"7F",X"FF",X"F0",X"B5",X"7F",X"4E",X"79",X"93",X"70",X"00",X"4E",X"FF",X"F0",X"84",X"8F",X"4F",
		X"4B",X"64",X"60",X"30",X"9F",X"FF",X"90",X"C0",X"F6",X"BD",X"4C",X"09",X"02",X"46",X"FF",X"F9",
		X"0A",X"0F",X"7E",X"A6",X"70",X"80",X"33",X"CF",X"BF",X"09",X"1B",X"98",X"D6",X"A1",X"52",X"36",
		X"FE",X"FE",X"3A",X"49",X"99",X"D6",X"50",X"11",X"5F",X"FF",X"F9",X"C1",X"82",X"A8",X"79",X"18",
		X"0E",X"9E",X"CC",X"CA",X"86",X"A6",X"62",X"37",X"6E",X"F8",X"F4",X"B5",X"8B",X"6D",X"25",X"16",
		X"CE",X"DF",X"5C",X"2A",X"56",X"72",X"87",X"DF",X"8F",X"0D",X"0E",X"58",X"40",X"A6",X"F7",X"F1",
		X"B3",X"97",X"46",X"0D",X"7F",X"AF",X"17",X"29",X"56",X"53",X"DB",X"F9",X"F0",X"72",X"87",X"45",
		X"6A",X"FE",X"F3",X"80",X"93",X"63",X"AA",X"FF",X"F5",X"52",X"36",X"59",X"9E",X"FE",X"B7",X"61",
		X"31",X"5A",X"FF",X"FC",X"54",X"23",X"33",X"8C",X"FF",X"FA",X"63",X"22",X"25",X"AE",X"FE",X"D6",
		X"71",X"31",X"4A",X"CF",X"EF",X"59",X"04",X"02",X"AA",X"FD",X"F7",X"92",X"10",X"19",X"AF",X"CF",
		X"6B",X"03",X"12",X"A9",X"FC",X"F5",X"90",X"31",X"3A",X"BF",X"DF",X"69",X"12",X"02",X"9B",X"FD",
		X"F7",X"A1",X"30",X"57",X"DF",X"FF",X"8A",X"03",X"05",X"8E",X"FF",X"D9",X"60",X"10",X"78",X"FF",
		X"F9",X"A3",X"20",X"09",X"9F",X"DF",X"5B",X"03",X"02",X"7C",X"06",X"F8",X"90",X"20",X"06",X"EF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
