`define BUILD_DATE "180812"
`define BUILD_TIME "154434"
