library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity tn02 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of tn02 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"AF",X"BE",X"C2",X"0B",X"08",X"78",X"FE",X"3E",X"D2",X"69",X"08",X"78",X"FE",X"3C",X"DA",X"25",
		X"08",X"2A",X"09",X"20",X"01",X"1E",X"02",X"CD",X"8C",X"08",X"21",X"05",X"20",X"36",X"00",X"21",
		X"BF",X"20",X"36",X"00",X"C9",X"2A",X"07",X"20",X"EB",X"2A",X"09",X"20",X"01",X"1E",X"02",X"C3",
		X"D5",X"01",X"36",X"FF",X"21",X"05",X"21",X"CD",X"A0",X"08",X"EB",X"2E",X"06",X"CD",X"52",X"1A",
		X"E5",X"C1",X"0A",X"6F",X"03",X"0A",X"67",X"CD",X"D2",X"01",X"C3",X"25",X"08",X"36",X"FF",X"21",
		X"09",X"21",X"CD",X"A0",X"08",X"EB",X"2E",X"0A",X"C3",X"3D",X"08",X"36",X"FF",X"21",X"0D",X"21",
		X"CD",X"A0",X"08",X"EB",X"2E",X"0E",X"C3",X"3D",X"08",X"36",X"FF",X"21",X"11",X"21",X"CD",X"A0",
		X"08",X"EB",X"2E",X"12",X"C3",X"3D",X"08",X"21",X"06",X"20",X"34",X"7E",X"E6",X"01",X"C2",X"85",
		X"08",X"21",X"72",X"40",X"C9",X"21",X"36",X"40",X"C9",X"01",X"20",X"03",X"AF",X"C5",X"E5",X"77",
		X"23",X"05",X"C2",X"8F",X"08",X"E1",X"01",X"20",X"00",X"09",X"C1",X"0D",X"C2",X"8D",X"08",X"C9",
		X"7E",X"21",X"1D",X"41",X"3D",X"C8",X"11",X"60",X"00",X"19",X"C3",X"A4",X"08",X"AF",X"7C",X"1F",
		X"57",X"7D",X"1F",X"E6",X"F0",X"0F",X"0F",X"0F",X"0F",X"5F",X"7A",X"E6",X"0F",X"07",X"07",X"07",
		X"07",X"B3",X"C9",X"11",X"DD",X"43",X"06",X"02",X"C3",X"AD",X"0E",X"11",X"DD",X"43",X"06",X"02",
		X"C3",X"9A",X"19",X"CD",X"38",X"14",X"CD",X"53",X"14",X"CD",X"40",X"10",X"CD",X"42",X"09",X"CD",
		X"F8",X"08",X"CD",X"65",X"09",X"3A",X"E4",X"20",X"A7",X"CA",X"22",X"05",X"CD",X"89",X"1A",X"CD",
		X"13",X"09",X"CD",X"35",X"1B",X"C3",X"22",X"05",X"21",X"1F",X"20",X"7E",X"A7",X"C8",X"46",X"36",
		X"00",X"21",X"24",X"20",X"7E",X"0F",X"D0",X"36",X"00",X"2A",X"22",X"20",X"EB",X"21",X"38",X"20",
		X"C3",X"0D",X"0A",X"CD",X"52",X"1A",X"2E",X"24",X"7E",X"FE",X"03",X"D8",X"21",X"BF",X"20",X"AF",
		X"BE",X"C0",X"34",X"21",X"35",X"09",X"C3",X"7B",X"1A",X"00",X"00",X"07",X"07",X"01",X"00",X"01",
		X"00",X"06",X"06",X"01",X"00",X"00",X"00",X"04",X"04",X"01",X"00",X"00",X"02",X"00",X"01",X"01",
		X"01",X"00",X"3A",X"E4",X"20",X"A7",X"C8",X"21",X"38",X"20",X"7E",X"FE",X"FF",X"CA",X"60",X"09",
		X"0F",X"D2",X"59",X"09",X"3E",X"10",X"C3",X"0E",X"02",X"23",X"23",X"23",X"23",X"C3",X"4A",X"09",
		X"3E",X"10",X"C3",X"17",X"02",X"21",X"04",X"20",X"34",X"7E",X"E6",X"03",X"77",X"A7",X"CA",X"28",
		X"19",X"FE",X"01",X"CA",X"38",X"19",X"FE",X"02",X"CA",X"66",X"19",X"FE",X"03",X"CA",X"85",X"19",
		X"C9",X"21",X"38",X"20",X"CD",X"21",X"0A",X"21",X"3C",X"20",X"CD",X"21",X"0A",X"11",X"9D",X"20",
		X"CD",X"DF",X"09",X"CD",X"07",X"13",X"CD",X"6A",X"0A",X"C3",X"D9",X"09",X"21",X"40",X"20",X"CD",
		X"21",X"0A",X"21",X"44",X"20",X"CD",X"21",X"0A",X"11",X"9E",X"20",X"CD",X"DF",X"09",X"2E",X"0C",
		X"CD",X"52",X"1A",X"CD",X"6A",X"0A",X"CD",X"D9",X"09",X"C3",X"15",X"15",X"21",X"48",X"20",X"CD",
		X"21",X"0A",X"21",X"4C",X"20",X"CD",X"21",X"0A",X"11",X"9F",X"20",X"CD",X"DF",X"09",X"2E",X"14",
		X"CD",X"52",X"1A",X"CD",X"6A",X"0A",X"C3",X"D9",X"09",X"21",X"9C",X"20",X"36",X"00",X"C9",X"21",
		X"9B",X"20",X"7E",X"A7",X"CA",X"EB",X"09",X"23",X"36",X"00",X"C9",X"EB",X"34",X"7E",X"FE",X"02",
		X"D2",X"F8",X"09",X"EB",X"23",X"36",X"FF",X"C9",X"36",X"00",X"EB",X"23",X"36",X"00",X"C9",X"57",
		X"3A",X"9C",X"20",X"A7",X"7A",X"C2",X"0A",X"0A",X"37",X"C9",X"37",X"3F",X"C9",X"78",X"3D",X"CA",
		X"19",X"0A",X"23",X"23",X"23",X"23",X"C3",X"0E",X"0A",X"36",X"01",X"23",X"23",X"73",X"23",X"72",
		X"C9",X"7E",X"0F",X"D0",X"23",X"23",X"E5",X"CD",X"6C",X"11",X"CD",X"5B",X"0A",X"E1",X"E5",X"CD",
		X"6C",X"11",X"7D",X"FE",X"18",X"DA",X"48",X"0A",X"01",X"F9",X"FF",X"09",X"EB",X"E1",X"73",X"23",
		X"72",X"EB",X"11",X"DA",X"43",X"C3",X"CF",X"0E",X"E1",X"E5",X"CD",X"6C",X"11",X"22",X"B7",X"20",
		X"E1",X"2B",X"AF",X"77",X"2B",X"77",X"21",X"B5",X"20",X"34",X"C9",X"11",X"DA",X"43",X"C3",X"AB",
		X"0E",X"7C",X"B5",X"37",X"C8",X"7B",X"95",X"7A",X"9C",X"C9",X"E5",X"7E",X"47",X"07",X"D2",X"8A",
		X"0A",X"23",X"23",X"CD",X"15",X"0B",X"78",X"0F",X"0F",X"7A",X"D2",X"DA",X"0A",X"FE",X"4B",X"DA",
		X"A1",X"0A",X"36",X"25",X"E1",X"E5",X"3E",X"DF",X"A6",X"77",X"21",X"37",X"20",X"34",X"E1",X"23",
		X"23",X"23",X"23",X"3A",X"37",X"20",X"FE",X"02",X"DA",X"6A",X"0A",X"21",X"37",X"20",X"36",X"00",
		X"C9",X"FE",X"3C",X"D2",X"CC",X"0A",X"78",X"0F",X"E1",X"E5",X"23",X"7E",X"23",X"4E",X"23",X"46",
		X"2B",X"2B",X"DA",X"2F",X"0B",X"CD",X"FF",X"09",X"D2",X"BF",X"0A",X"3D",X"CA",X"23",X"0B",X"77",
		X"CD",X"A1",X"08",X"EB",X"60",X"69",X"CD",X"D2",X"01",X"C3",X"8A",X"0A",X"E1",X"E5",X"CD",X"03",
		X"0B",X"E1",X"E5",X"7E",X"0F",X"0F",X"0F",X"C3",X"8A",X"0A",X"2B",X"2B",X"2B",X"FE",X"25",X"DA",
		X"EE",X"0A",X"FE",X"3C",X"DA",X"FB",X"0A",X"7E",X"0F",X"0F",X"0F",X"C3",X"8A",X"0A",X"CD",X"08",
		X"0B",X"E1",X"E5",X"23",X"23",X"23",X"36",X"48",X"C3",X"8A",X"0A",X"46",X"3E",X"DF",X"A6",X"77",
		X"C3",X"A6",X"0A",X"7E",X"07",X"07",X"07",X"D8",X"3E",X"20",X"B6",X"77",X"23",X"23",X"5E",X"23",
		X"56",X"EB",X"C3",X"89",X"08",X"E5",X"5E",X"23",X"56",X"2A",X"28",X"21",X"19",X"EB",X"E1",X"73",
		X"23",X"72",X"C9",X"36",X"01",X"2B",X"3E",X"01",X"B6",X"77",X"3E",X"01",X"C3",X"C0",X"0A",X"CD",
		X"FF",X"09",X"D2",X"BF",X"0A",X"3C",X"FE",X"08",X"DA",X"BF",X"0A",X"36",X"07",X"2B",X"3E",X"FE",
		X"A6",X"77",X"3E",X"07",X"C3",X"C0",X"0A",X"CD",X"56",X"0B",X"CD",X"AB",X"0B",X"CD",X"D6",X"0B",
		X"CD",X"40",X"15",X"C3",X"27",X"16",X"AF",X"21",X"B5",X"20",X"BE",X"C8",X"23",X"34",X"7E",X"FE",
		X"01",X"CA",X"01",X"0C",X"FE",X"04",X"CA",X"07",X"0C",X"FE",X"07",X"D8",X"11",X"3C",X"44",X"CD",
		X"0A",X"0C",X"CD",X"E0",X"15",X"21",X"B8",X"20",X"D2",X"81",X"0B",X"CD",X"9B",X"0B",X"C3",X"84",
		X"0B",X"CD",X"8B",X"0B",X"21",X"00",X"00",X"22",X"B5",X"20",X"C9",X"AF",X"3A",X"34",X"20",X"BE",
		X"D8",X"7E",X"21",X"7D",X"20",X"BE",X"D8",X"77",X"C3",X"0D",X"16",X"AF",X"3A",X"34",X"20",X"BE",
		X"D0",X"7E",X"21",X"7F",X"20",X"BE",X"D0",X"77",X"C3",X"ED",X"15",X"AF",X"21",X"1D",X"20",X"BE",
		X"C8",X"23",X"34",X"7E",X"FE",X"01",X"CA",X"16",X"0C",X"FE",X"04",X"CA",X"1C",X"0C",X"FE",X"07",
		X"D8",X"2A",X"22",X"20",X"CD",X"76",X"03",X"01",X"10",X"02",X"CD",X"8C",X"08",X"21",X"00",X"00",
		X"22",X"1D",X"20",X"C3",X"7D",X"15",X"AF",X"21",X"27",X"20",X"BE",X"C8",X"23",X"34",X"7E",X"FE",
		X"01",X"CA",X"2B",X"0C",X"FE",X"04",X"CA",X"47",X"0C",X"FE",X"07",X"D8",X"2A",X"2D",X"20",X"01",
		X"10",X"02",X"CD",X"8C",X"08",X"21",X"00",X"00",X"22",X"27",X"20",X"CD",X"6F",X"1A",X"C3",X"7D",
		X"15",X"11",X"0C",X"44",X"C3",X"0A",X"0C",X"11",X"24",X"44",X"2A",X"B7",X"20",X"CD",X"76",X"03",
		X"01",X"0C",X"02",X"C3",X"D5",X"01",X"11",X"54",X"44",X"C3",X"1F",X"0C",X"11",X"74",X"44",X"2A",
		X"22",X"20",X"CD",X"76",X"03",X"01",X"10",X"02",X"C3",X"D5",X"01",X"2A",X"29",X"20",X"11",X"DA",
		X"43",X"CD",X"AD",X"0E",X"2A",X"29",X"20",X"CD",X"76",X"03",X"22",X"2D",X"20",X"11",X"94",X"44",
		X"01",X"10",X"02",X"CD",X"D5",X"01",X"C9",X"2A",X"2D",X"20",X"11",X"B4",X"44",X"C3",X"40",X"0C",
		X"3A",X"E4",X"20",X"A7",X"C8",X"3A",X"DB",X"20",X"0F",X"DB",X"01",X"D0",X"DB",X"02",X"C9",X"21",
		X"2F",X"20",X"AF",X"BE",X"C8",X"23",X"BE",X"C2",X"6E",X"0C",X"34",X"CD",X"E4",X"0C",X"3A",X"E4",
		X"20",X"A7",X"C2",X"9D",X"0C",X"2A",X"E2",X"20",X"3A",X"E1",X"20",X"3C",X"32",X"E1",X"20",X"E6",
		X"0F",X"C2",X"8B",X"0C",X"7D",X"FE",X"13",X"CC",X"9A",X"0C",X"23",X"22",X"E2",X"20",X"7E",X"0F",
		X"DA",X"06",X"0D",X"0F",X"DA",X"23",X"0D",X"C3",X"A9",X"0C",X"2E",X"00",X"C9",X"CD",X"50",X"0C",
		X"07",X"07",X"DA",X"06",X"0D",X"07",X"DA",X"23",X"0D",X"06",X"00",X"21",X"32",X"20",X"70",X"CD",
		X"E4",X"0C",X"21",X"31",X"20",X"CD",X"A1",X"0D",X"2A",X"33",X"20",X"11",X"BE",X"43",X"01",X"02",
		X"0E",X"CD",X"71",X"03",X"C5",X"E5",X"1A",X"A6",X"CA",X"D0",X"0C",X"3E",X"01",X"32",X"35",X"20",
		X"1A",X"AE",X"77",X"23",X"13",X"0D",X"C2",X"C6",X"0C",X"E1",X"01",X"20",X"00",X"09",X"C1",X"05",
		X"C2",X"C4",X"0C",X"C9",X"2A",X"33",X"20",X"11",X"BE",X"43",X"01",X"02",X"0E",X"CD",X"71",X"03",
		X"C5",X"E5",X"1A",X"AE",X"77",X"23",X"13",X"0D",X"C2",X"F2",X"0C",X"E1",X"01",X"20",X"00",X"09",
		X"C1",X"05",X"C2",X"F0",X"0C",X"C9",X"3A",X"34",X"20",X"FE",X"DA",X"D2",X"A9",X"0C",X"2A",X"33",
		X"20",X"01",X"F8",X"0F",X"09",X"CD",X"76",X"03",X"7E",X"FE",X"7F",X"C2",X"A9",X"0C",X"06",X"02",
		X"C3",X"AB",X"0C",X"3A",X"34",X"20",X"FE",X"38",X"DA",X"A9",X"0C",X"2A",X"33",X"20",X"01",X"F8",
		X"FC",X"09",X"CD",X"76",X"03",X"7E",X"FE",X"7F",X"C2",X"A9",X"0C",X"06",X"FE",X"C3",X"AB",X"0C",
		X"23",X"23",X"5E",X"23",X"7E",X"C6",X"02",X"57",X"EB",X"CD",X"AD",X"08",X"57",X"7D",X"E6",X"1F",
		X"07",X"07",X"07",X"5F",X"EB",X"C9",X"21",X"54",X"20",X"AF",X"BE",X"C8",X"23",X"BE",X"C2",X"73",
		X"0D",X"34",X"23",X"BE",X"21",X"00",X"FD",X"22",X"58",X"20",X"21",X"C8",X"D0",X"C4",X"1A",X"0E",
		X"22",X"5A",X"20",X"3A",X"56",X"20",X"A7",X"21",X"5B",X"20",X"7E",X"C2",X"AD",X"0D",X"FE",X"28",
		X"DA",X"C9",X"0D",X"21",X"57",X"20",X"34",X"E6",X"01",X"21",X"AE",X"40",X"CC",X"C1",X"0D",X"22",
		X"5C",X"20",X"21",X"5A",X"20",X"CD",X"F0",X"0D",X"CD",X"02",X"0E",X"CD",X"24",X"0E",X"21",X"58",
		X"20",X"4E",X"23",X"46",X"23",X"79",X"86",X"77",X"23",X"78",X"86",X"77",X"C9",X"FE",X"D0",X"D2",
		X"C9",X"0D",X"21",X"57",X"20",X"34",X"E6",X"01",X"21",X"36",X"40",X"CC",X"C5",X"0D",X"C3",X"8F",
		X"0D",X"21",X"E5",X"40",X"C9",X"21",X"72",X"40",X"C9",X"2A",X"5A",X"20",X"01",X"1B",X"02",X"CD",
		X"76",X"03",X"CD",X"8C",X"08",X"06",X"0C",X"21",X"54",X"46",X"11",X"54",X"20",X"CD",X"8B",X"03",
		X"21",X"13",X"20",X"34",X"7E",X"E6",X"01",X"21",X"56",X"20",X"36",X"01",X"C0",X"36",X"00",X"C9",
		X"E5",X"23",X"23",X"5E",X"23",X"56",X"23",X"4E",X"23",X"46",X"E1",X"D5",X"5E",X"23",X"56",X"EB",
		X"D1",X"C9",X"CD",X"76",X"03",X"C5",X"E5",X"1A",X"77",X"23",X"13",X"0D",X"C2",X"07",X"0E",X"E1",
		X"01",X"20",X"00",X"09",X"C1",X"05",X"C2",X"05",X"0E",X"C9",X"21",X"00",X"03",X"22",X"58",X"20",
		X"21",X"C8",X"28",X"C9",X"3A",X"56",X"20",X"A7",X"C2",X"A1",X"0E",X"CD",X"35",X"0E",X"D6",X"0A",
		X"B8",X"DA",X"3D",X"0E",X"C9",X"2A",X"34",X"20",X"44",X"3A",X"0A",X"20",X"C9",X"21",X"B0",X"20",
		X"AF",X"BE",X"CA",X"47",X"0E",X"35",X"C9",X"E5",X"CD",X"4B",X"1A",X"23",X"7E",X"FE",X"04",X"06",
		X"50",X"D2",X"56",X"0E",X"06",X"60",X"E1",X"70",X"FE",X"0B",X"D2",X"7A",X"0E",X"FE",X"09",X"CD",
		X"52",X"1A",X"2E",X"24",X"7E",X"FE",X"04",X"D2",X"8F",X"0E",X"21",X"60",X"20",X"34",X"2E",X"67",
		X"34",X"2E",X"6E",X"34",X"21",X"95",X"20",X"36",X"00",X"C9",X"21",X"FB",X"03",X"22",X"63",X"20",
		X"21",X"FA",X"02",X"22",X"6A",X"20",X"21",X"FB",X"FA",X"22",X"71",X"20",X"C3",X"6A",X"0E",X"21",
		X"FC",X"02",X"22",X"63",X"20",X"21",X"FB",X"01",X"22",X"6A",X"20",X"21",X"FB",X"FD",X"C3",X"89",
		X"0E",X"CD",X"35",X"0E",X"C6",X"08",X"B8",X"D2",X"3D",X"0E",X"C9",X"06",X"03",X"CD",X"71",X"03",
		X"C5",X"E5",X"1A",X"D3",X"04",X"DB",X"03",X"2F",X"A6",X"77",X"23",X"13",X"AF",X"D3",X"04",X"DB",
		X"03",X"2F",X"A6",X"77",X"E1",X"01",X"20",X"00",X"09",X"C1",X"05",X"C2",X"B0",X"0E",X"C9",X"06",
		X"03",X"CD",X"71",X"03",X"C5",X"E5",X"1A",X"D3",X"04",X"DB",X"03",X"AE",X"77",X"23",X"13",X"AF",
		X"D3",X"04",X"DB",X"03",X"AE",X"77",X"E1",X"01",X"20",X"00",X"09",X"C1",X"05",X"C2",X"D4",X"0E",
		X"C9",X"21",X"60",X"20",X"AF",X"BE",X"C8",X"23",X"BE",X"C2",X"FE",X"0E",X"35",X"C9",X"23",X"BE",
		X"C2",X"0A",X"0F",X"34",X"CD",X"33",X"0F",X"22",X"65",X"20",X"CD",X"3B",X"0F",X"21",X"66",X"20",
		X"7E",X"FE",X"30",X"DC",X"46",X"0F",X"FE",X"E8",X"D4",X"53",X"0F",X"2B",X"7E",X"FE",X"18",X"DA",
		X"5E",X"0F",X"21",X"63",X"20",X"CD",X"A1",X"0D",X"2A",X"65",X"20",X"11",X"DA",X"0F",X"06",X"08",
		X"C3",X"D1",X"0E",X"2A",X"5A",X"20",X"01",X"00",X"08",X"09",X"C9",X"2A",X"65",X"20",X"11",X"DA",
		X"0F",X"06",X"08",X"C3",X"AD",X"0E",X"F5",X"E5",X"2A",X"65",X"20",X"CD",X"3E",X"0F",X"E1",X"36",
		X"E0",X"F1",X"C9",X"E5",X"2A",X"65",X"20",X"CD",X"3E",X"0F",X"E1",X"36",X"34",X"C9",X"CD",X"3B",
		X"0F",X"21",X"60",X"46",X"11",X"60",X"20",X"06",X"07",X"C3",X"8B",X"03",X"21",X"67",X"20",X"AF",
		X"BE",X"C8",X"23",X"BE",X"CA",X"79",X"0F",X"35",X"C9",X"23",X"BE",X"C2",X"85",X"0F",X"34",X"CD",
		X"33",X"0F",X"22",X"6C",X"20",X"2A",X"6C",X"20",X"CD",X"3E",X"0F",X"21",X"6D",X"20",X"7E",X"FE",
		X"30",X"DC",X"BC",X"0F",X"FE",X"E8",X"D4",X"C4",X"0F",X"2B",X"7E",X"47",X"CD",X"52",X"1A",X"2E",
		X"24",X"7E",X"FE",X"05",X"0E",X"13",X"D2",X"AB",X"0F",X"0E",X"18",X"78",X"B9",X"DA",X"CB",X"0F",
		X"21",X"6A",X"20",X"CD",X"A1",X"0D",X"2A",X"6C",X"20",X"C3",X"2B",X"0F",X"F5",X"E5",X"2A",X"6C",
		X"20",X"C3",X"57",X"0F",X"E5",X"2A",X"6C",X"20",X"C3",X"4B",X"0F",X"2A",X"6C",X"20",X"CD",X"3E",
		X"0F",X"21",X"67",X"46",X"11",X"67",X"20",X"C3",X"67",X"0F",X"60",X"F0",X"F0",X"F0",X"F0",X"60",
		X"90",X"90",X"21",X"6E",X"20",X"AF",X"BE",X"C8",X"23",X"BE",X"CA",X"EF",X"0F",X"35",X"C9",X"23",
		X"BE",X"C2",X"FB",X"0F",X"34",X"CD",X"33",X"0F",X"22",X"73",X"20",X"2A",X"73",X"20",X"CD",X"3E");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
